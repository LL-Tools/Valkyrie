

module b20_C_AntiSAT_k_128_8 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, 
        ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, 
        ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, 
        ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, 
        ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, 
        U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, 
        P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, 
        P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, 
        P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, 
        P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, 
        P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, 
        P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, 
        P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, 
        P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, 
        P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, 
        P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, 
        P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, 
        P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, 
        P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, 
        P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, 
        P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, 
        P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, 
        P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, 
        P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, 
        P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, 
        P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, 
        P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, 
        P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, 
        P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, 
        P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, 
        P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, 
        P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, 
        P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, 
        P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, 
        P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, 
        P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, 
        P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, 
        P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, 
        P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, 
        P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, 
        P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, 
        P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, 
        P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, 
        P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, 
        P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, 
        P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, 
        P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, 
        P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, 
        P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, 
        P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, 
        P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, 
        P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, 
        P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, 
        P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, 
        P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, 
        P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, 
        P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, 
        P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, 
        P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, 
        P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, 
        P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, 
        P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, 
        P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, 
        P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, 
        P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, 
        P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, 
        P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, 
        P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, 
        P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, 
        P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, 
        P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, 
        P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, 
        P2_U3893 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339,
         n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349,
         n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359,
         n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369,
         n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379,
         n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389,
         n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399,
         n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409,
         n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419,
         n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429,
         n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439,
         n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449,
         n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459,
         n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469,
         n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479,
         n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489,
         n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499,
         n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509,
         n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519,
         n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529,
         n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539,
         n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549,
         n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559,
         n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569,
         n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579,
         n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589,
         n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599,
         n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609,
         n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619,
         n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
         n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
         n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
         n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
         n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669,
         n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679,
         n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689,
         n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
         n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
         n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719,
         n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729,
         n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739,
         n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749,
         n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759,
         n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769,
         n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779,
         n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789,
         n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799,
         n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809,
         n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819,
         n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829,
         n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839,
         n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849,
         n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859,
         n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869,
         n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879,
         n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889,
         n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899,
         n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909,
         n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919,
         n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929,
         n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939,
         n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949,
         n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959,
         n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969,
         n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979,
         n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989,
         n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999,
         n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009,
         n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019,
         n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029,
         n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039,
         n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049,
         n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059,
         n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069,
         n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079,
         n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089,
         n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099,
         n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109,
         n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119,
         n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129,
         n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139,
         n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149,
         n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159,
         n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169,
         n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179,
         n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189,
         n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199,
         n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209,
         n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219,
         n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229,
         n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239,
         n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249,
         n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259,
         n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269,
         n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279,
         n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289,
         n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299,
         n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309,
         n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319,
         n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329,
         n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339,
         n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349,
         n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359,
         n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369,
         n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379,
         n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389,
         n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399,
         n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409,
         n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419,
         n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429,
         n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439,
         n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449,
         n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459,
         n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469,
         n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479,
         n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489,
         n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499,
         n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509,
         n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519,
         n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529,
         n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539,
         n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549,
         n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559,
         n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569,
         n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579,
         n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589,
         n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599,
         n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609,
         n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619,
         n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629,
         n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639,
         n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649,
         n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659,
         n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669,
         n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679,
         n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689,
         n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699,
         n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709,
         n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719,
         n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729,
         n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739,
         n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749,
         n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759,
         n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769,
         n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779,
         n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789,
         n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799,
         n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809,
         n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819,
         n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829,
         n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839,
         n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849,
         n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859,
         n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869,
         n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879,
         n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889,
         n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899,
         n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909,
         n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919,
         n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929,
         n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939,
         n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949,
         n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959,
         n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969,
         n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979,
         n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989,
         n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999,
         n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009,
         n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019,
         n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029,
         n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039,
         n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049,
         n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059,
         n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069,
         n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079,
         n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089,
         n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099,
         n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109,
         n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119,
         n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129,
         n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139,
         n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149,
         n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159,
         n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169,
         n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179,
         n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189,
         n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199,
         n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209,
         n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219,
         n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229,
         n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239,
         n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249,
         n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259,
         n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269,
         n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279,
         n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289,
         n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299,
         n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309,
         n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319,
         n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329,
         n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339,
         n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349,
         n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359,
         n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369,
         n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379,
         n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389,
         n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399,
         n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409,
         n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419,
         n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429,
         n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439,
         n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449,
         n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459,
         n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469,
         n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479,
         n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489,
         n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499,
         n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509,
         n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519,
         n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529,
         n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539,
         n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549,
         n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559,
         n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569,
         n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579,
         n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589,
         n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599,
         n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609,
         n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619,
         n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629,
         n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639,
         n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649,
         n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659,
         n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669,
         n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679,
         n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689,
         n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699,
         n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709,
         n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719,
         n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729,
         n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739,
         n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749,
         n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759,
         n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769,
         n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779,
         n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789,
         n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799,
         n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809,
         n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819,
         n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829,
         n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839,
         n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849,
         n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859,
         n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869,
         n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879,
         n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889,
         n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899,
         n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909,
         n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919,
         n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929,
         n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939,
         n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949,
         n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959,
         n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969,
         n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979,
         n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989,
         n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999,
         n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009,
         n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019,
         n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029,
         n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039,
         n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049,
         n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059,
         n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069,
         n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079,
         n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089,
         n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099,
         n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109,
         n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119,
         n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129,
         n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139,
         n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149,
         n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159,
         n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169,
         n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179,
         n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189,
         n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199,
         n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209,
         n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219,
         n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229,
         n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239,
         n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249,
         n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259,
         n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269,
         n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279,
         n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289,
         n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299,
         n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309,
         n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319,
         n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329,
         n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339,
         n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349,
         n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359,
         n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369,
         n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379,
         n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389,
         n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399,
         n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409,
         n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419,
         n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429,
         n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439,
         n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449,
         n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459,
         n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469,
         n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479,
         n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489,
         n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499,
         n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509,
         n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519,
         n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529,
         n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539,
         n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549,
         n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559,
         n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569,
         n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579,
         n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589,
         n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599,
         n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609,
         n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619,
         n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629,
         n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639,
         n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649,
         n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659,
         n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669,
         n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679,
         n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689,
         n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699,
         n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709,
         n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719,
         n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729,
         n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739,
         n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749,
         n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759,
         n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769,
         n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779,
         n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789,
         n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799,
         n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809,
         n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819,
         n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829,
         n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839,
         n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849,
         n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859,
         n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869,
         n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879,
         n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889,
         n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899,
         n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909,
         n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919,
         n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929,
         n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939,
         n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949,
         n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959,
         n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969,
         n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979,
         n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989,
         n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999,
         n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009,
         n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019,
         n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029,
         n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039,
         n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049,
         n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059,
         n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069,
         n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079,
         n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089,
         n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099,
         n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109,
         n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119,
         n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129,
         n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139,
         n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149,
         n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159,
         n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169,
         n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179,
         n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189,
         n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199,
         n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209,
         n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219,
         n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229,
         n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239,
         n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249,
         n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259,
         n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269,
         n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279,
         n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289,
         n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299,
         n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309,
         n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319,
         n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329,
         n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339,
         n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349,
         n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359,
         n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369,
         n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379,
         n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389,
         n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399,
         n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409,
         n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419,
         n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429,
         n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439,
         n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449,
         n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459,
         n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469,
         n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479,
         n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489,
         n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499,
         n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509,
         n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519,
         n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529,
         n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539,
         n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549,
         n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559,
         n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569,
         n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579,
         n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589,
         n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599,
         n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609,
         n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619,
         n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629,
         n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639,
         n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649,
         n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659,
         n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669,
         n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679,
         n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689,
         n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699,
         n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709,
         n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719,
         n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729,
         n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739,
         n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749,
         n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759,
         n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769,
         n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779,
         n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789,
         n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799,
         n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809,
         n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819,
         n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829,
         n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839,
         n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849,
         n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859,
         n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869,
         n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879,
         n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889,
         n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899,
         n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909,
         n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919,
         n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929,
         n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939,
         n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949,
         n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959,
         n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969,
         n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979,
         n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989,
         n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999,
         n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009,
         n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019,
         n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029,
         n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039,
         n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049,
         n9050, n9051, n9052, n9054, n9055, n9056, n9057, n9058, n9059, n9060,
         n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070,
         n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080,
         n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090,
         n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100,
         n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110,
         n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120,
         n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130,
         n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140,
         n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150,
         n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160,
         n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170,
         n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180,
         n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190,
         n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200,
         n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210,
         n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220,
         n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230,
         n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240,
         n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250,
         n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260,
         n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270,
         n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280,
         n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290,
         n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300,
         n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310,
         n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320,
         n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330,
         n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340,
         n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350,
         n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360,
         n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370,
         n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380,
         n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390,
         n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400,
         n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410,
         n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420,
         n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430,
         n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440,
         n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450,
         n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460,
         n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470,
         n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480,
         n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490,
         n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500,
         n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510,
         n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520,
         n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530,
         n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540,
         n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550,
         n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560,
         n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570,
         n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580,
         n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590,
         n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600,
         n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610,
         n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620,
         n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630,
         n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640,
         n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650,
         n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660,
         n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670,
         n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680,
         n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690,
         n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700,
         n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710,
         n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720,
         n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730,
         n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740,
         n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750,
         n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760,
         n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770,
         n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780,
         n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790,
         n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800,
         n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810,
         n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820,
         n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830,
         n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840,
         n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850,
         n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860,
         n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870,
         n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880,
         n9881, n9882, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891,
         n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901,
         n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911,
         n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921,
         n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931,
         n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941,
         n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951,
         n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961,
         n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971,
         n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981,
         n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991,
         n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209;

  INV_X2 U4836 ( .A(n8584), .ZN(n8748) );
  INV_X1 U4837 ( .A(n6810), .ZN(n6777) );
  NAND2_X1 U4838 ( .A1(n6303), .A2(n6302), .ZN(n7105) );
  INV_X1 U4839 ( .A(n6285), .ZN(n6216) );
  INV_X1 U4840 ( .A(n8567), .ZN(n8552) );
  BUF_X2 U4841 ( .A(n4997), .Z(n5465) );
  INV_X1 U4842 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n6138) );
  OR2_X1 U4843 ( .A1(n6374), .A2(n5944), .ZN(n5952) );
  CLKBUF_X2 U4844 ( .A(n4995), .Z(n4331) );
  AND2_X1 U4846 ( .A1(n4769), .A2(n4358), .ZN(n8677) );
  AND2_X1 U4847 ( .A1(n6443), .A2(n8358), .ZN(n5967) );
  INV_X1 U4848 ( .A(n8368), .ZN(n6282) );
  INV_X2 U4849 ( .A(n6443), .ZN(n6184) );
  INV_X2 U4851 ( .A(n5874), .ZN(n5886) );
  XNOR2_X1 U4852 ( .A(n9540), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n9548) );
  NAND2_X1 U4853 ( .A1(n5088), .A2(n5087), .ZN(n4825) );
  NOR2_X1 U4854 ( .A1(n8610), .A2(n8972), .ZN(n8425) );
  AOI211_X1 U4856 ( .C1(n9548), .C2(n9915), .A(n9937), .B(n9547), .ZN(n9550)
         );
  NAND2_X1 U4857 ( .A1(n5670), .A2(n9298), .ZN(n5671) );
  NOR2_X1 U4858 ( .A1(n9787), .A2(n9709), .ZN(n9690) );
  INV_X1 U4859 ( .A(n7302), .ZN(n9976) );
  NAND2_X1 U4860 ( .A1(n4825), .A2(n5090), .ZN(n5131) );
  NAND3_X2 U4861 ( .A1(n5951), .A2(n5952), .A3(n6489), .ZN(n6443) );
  AOI211_X1 U4862 ( .C1(n7725), .C2(n7724), .A(n8353), .B(n7819), .ZN(n7726)
         );
  NAND2_X1 U4863 ( .A1(n8223), .A2(n8222), .ZN(n8303) );
  NAND2_X1 U4864 ( .A1(n8294), .A2(n4434), .ZN(n8331) );
  NAND2_X1 U4865 ( .A1(n5307), .A2(n5306), .ZN(n7946) );
  XNOR2_X1 U4866 ( .A(n5131), .B(n5129), .ZN(n6472) );
  INV_X2 U4867 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n6513) );
  INV_X1 U4868 ( .A(n6982), .ZN(n9336) );
  OR2_X1 U4869 ( .A1(n4616), .A2(n8376), .ZN(n4330) );
  NAND2_X2 U4870 ( .A1(n5071), .A2(n5070), .ZN(n5088) );
  AOI21_X2 U4871 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n7346), .A(n7345), .ZN(
        n7347) );
  NOR2_X2 U4872 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5968) );
  BUF_X2 U4873 ( .A(n4995), .Z(n4332) );
  NAND2_X1 U4874 ( .A1(n4539), .A2(n4538), .ZN(n4995) );
  NOR2_X2 U4875 ( .A1(n4925), .A2(n4924), .ZN(n4926) );
  XNOR2_X2 U4876 ( .A(n8219), .B(n8220), .ZN(n8234) );
  NAND2_X2 U4877 ( .A1(n8322), .A2(n8218), .ZN(n8219) );
  AOI21_X2 U4878 ( .B1(P1_REG2_REG_5__SCAN_IN), .B2(n6658), .A(n6652), .ZN(
        n6635) );
  OAI211_X2 U4879 ( .C1(n5052), .C2(n6450), .A(n4976), .B(n4975), .ZN(n6982)
         );
  XNOR2_X1 U4880 ( .A(n6357), .B(P2_IR_REG_27__SCAN_IN), .ZN(n4333) );
  XNOR2_X2 U4881 ( .A(n6357), .B(P2_IR_REG_27__SCAN_IN), .ZN(n6568) );
  AOI21_X1 U4882 ( .B1(n7250), .B2(n8604), .A(n7249), .ZN(n7252) );
  INV_X2 U4883 ( .A(n9723), .ZN(n4334) );
  INV_X1 U4884 ( .A(n7317), .ZN(n9985) );
  INV_X2 U4885 ( .A(n6256), .ZN(n6197) );
  XNOR2_X1 U4886 ( .A(n5933), .B(n5932), .ZN(n8181) );
  INV_X2 U4887 ( .A(n4982), .ZN(n4935) );
  NOR2_X1 U4888 ( .A1(n6137), .A2(n6136), .ZN(n6151) );
  OR2_X1 U4889 ( .A1(n6138), .A2(n5968), .ZN(n5969) );
  NOR2_X1 U4890 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(P1_IR_REG_26__SCAN_IN), .ZN(
        n4927) );
  INV_X2 U4891 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  AND2_X1 U4892 ( .A1(n9574), .A2(n9570), .ZN(n5592) );
  XNOR2_X1 U4893 ( .A(n5662), .B(n9411), .ZN(n8168) );
  NAND2_X1 U4894 ( .A1(n4425), .A2(n4424), .ZN(n6343) );
  NAND2_X1 U4895 ( .A1(n8852), .A2(n4422), .ZN(n8841) );
  NOR2_X1 U4896 ( .A1(n9277), .A2(n4560), .ZN(n4559) );
  AOI21_X1 U4897 ( .B1(n4787), .B2(n8631), .A(n4784), .ZN(n8765) );
  NAND2_X1 U4898 ( .A1(n8882), .A2(n8881), .ZN(n8880) );
  NAND2_X1 U4899 ( .A1(n9192), .A2(n9191), .ZN(n9190) );
  AND2_X1 U4900 ( .A1(n4725), .A2(n5788), .ZN(n9192) );
  OAI21_X1 U4901 ( .B1(n4463), .B2(n4362), .A(n4460), .ZN(n5785) );
  NAND2_X1 U4902 ( .A1(n4649), .A2(n4647), .ZN(n7862) );
  NAND2_X1 U4903 ( .A1(n6334), .A2(n6333), .ZN(n7836) );
  NAND2_X1 U4904 ( .A1(n5380), .A2(n5379), .ZN(n9831) );
  NOR2_X1 U4905 ( .A1(n4445), .A2(n5756), .ZN(n9856) );
  NOR2_X1 U4906 ( .A1(n7535), .A2(n4446), .ZN(n4445) );
  NOR2_X1 U4907 ( .A1(n7536), .A2(n7537), .ZN(n7535) );
  AOI21_X1 U4908 ( .B1(n9400), .B2(n5295), .A(n4383), .ZN(n4721) );
  OAI21_X1 U4909 ( .B1(n7585), .B2(P1_REG2_REG_12__SCAN_IN), .A(n7580), .ZN(
        n7583) );
  OR2_X1 U4910 ( .A1(n5297), .A2(n5296), .ZN(n5302) );
  NAND2_X1 U4911 ( .A1(n7252), .A2(n7251), .ZN(n7465) );
  OR2_X1 U4912 ( .A1(n7338), .A2(n5154), .ZN(n9342) );
  NAND2_X1 U4913 ( .A1(n5242), .A2(n5241), .ZN(n9076) );
  NAND2_X1 U4914 ( .A1(n4889), .A2(n4888), .ZN(n4892) );
  OAI21_X1 U4915 ( .B1(n5236), .B2(n5235), .A(n5234), .ZN(n5252) );
  OAI21_X1 U4916 ( .B1(n6844), .B2(n6843), .A(n6842), .ZN(n6845) );
  NAND2_X2 U4917 ( .A1(n6961), .A2(n8770), .ZN(n8915) );
  OR2_X1 U4918 ( .A1(n7080), .A2(n7079), .ZN(n7397) );
  OAI21_X1 U4919 ( .B1(n5213), .B2(n5212), .A(n5211), .ZN(n5236) );
  AOI21_X1 U4920 ( .B1(n5192), .B2(n5191), .A(n4897), .ZN(n5213) );
  NAND2_X2 U4921 ( .A1(n7034), .A2(n9727), .ZN(n9723) );
  AOI21_X1 U4922 ( .B1(n8626), .B2(n6985), .A(n8627), .ZN(n8633) );
  NAND2_X1 U4923 ( .A1(n8428), .A2(n8431), .ZN(n6298) );
  AND2_X2 U4924 ( .A1(n7645), .A2(n6440), .ZN(P1_U3973) );
  BUF_X2 U4925 ( .A(n5780), .Z(n5853) );
  CLKBUF_X2 U4926 ( .A(n6282), .Z(n8362) );
  INV_X1 U4927 ( .A(n5672), .ZN(n9970) );
  NAND2_X1 U4928 ( .A1(n6098), .A2(n6097), .ZN(n6116) );
  NAND4_X1 U4929 ( .A1(n5966), .A2(n5965), .A3(n5964), .A4(n5963), .ZN(n8608)
         );
  NAND2_X1 U4930 ( .A1(n5967), .A2(n6452), .ZN(n5955) );
  INV_X1 U4931 ( .A(n5967), .ZN(n6022) );
  NAND2_X1 U4932 ( .A1(n6439), .A2(n4766), .ZN(n5724) );
  AND2_X1 U4933 ( .A1(n5544), .A2(n5593), .ZN(n9296) );
  NAND4_X1 U4934 ( .A1(n4965), .A2(n4964), .A3(n4963), .A4(n4962), .ZN(n9468)
         );
  NAND2_X1 U4935 ( .A1(n5020), .A2(n5019), .ZN(n5032) );
  NAND4_X1 U4936 ( .A1(n4854), .A2(n4853), .A3(n4357), .A4(n4851), .ZN(n6695)
         );
  NAND4_X1 U4937 ( .A1(n4988), .A2(n4987), .A3(n4986), .A4(n4985), .ZN(n9467)
         );
  NAND2_X1 U4938 ( .A1(n5608), .A2(n5606), .ZN(n6439) );
  INV_X2 U4939 ( .A(n5013), .ZN(n5345) );
  AND2_X1 U4940 ( .A1(n6391), .A2(n4868), .ZN(n4866) );
  AND2_X2 U4941 ( .A1(n4936), .A2(n9851), .ZN(n4979) );
  XNOR2_X1 U4942 ( .A(n6373), .B(n6372), .ZN(n7816) );
  NAND2_X1 U4943 ( .A1(n9054), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5933) );
  OAI21_X1 U4944 ( .B1(n5604), .B2(n5603), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5605) );
  XNOR2_X1 U4945 ( .A(n4930), .B(n4929), .ZN(n4936) );
  XNOR2_X1 U4946 ( .A(n5547), .B(n5546), .ZN(n9298) );
  NOR2_X2 U4947 ( .A1(n6447), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6448) );
  AND2_X1 U4948 ( .A1(n5925), .A2(n6060), .ZN(n6290) );
  NAND2_X2 U4949 ( .A1(n6447), .A2(P1_U3086), .ZN(n7965) );
  AND2_X1 U4950 ( .A1(n6060), .A2(n6059), .ZN(n6083) );
  XNOR2_X1 U4951 ( .A(n4974), .B(P1_IR_REG_2__SCAN_IN), .ZN(n9891) );
  AND2_X1 U4952 ( .A1(n4723), .A2(n4945), .ZN(n4466) );
  BUF_X1 U4953 ( .A(n6509), .Z(n6540) );
  NAND3_X1 U4954 ( .A1(n4542), .A2(n4541), .A3(n4540), .ZN(n4539) );
  NAND3_X1 U4955 ( .A1(n4822), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n4538) );
  AND2_X1 U4956 ( .A1(n4927), .A2(n5597), .ZN(n4723) );
  INV_X1 U4957 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5340) );
  INV_X1 U4958 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5343) );
  INV_X1 U4959 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4542) );
  INV_X1 U4960 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5602) );
  INV_X1 U4961 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5600) );
  CLKBUF_X1 U4962 ( .A(P1_IR_REG_1__SCAN_IN), .Z(n4998) );
  INV_X1 U4963 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4822) );
  INV_X1 U4964 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5319) );
  NOR2_X1 U4965 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n4834) );
  INV_X1 U4966 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n8144) );
  INV_X1 U4967 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n4896) );
  INV_X1 U4968 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5914) );
  INV_X1 U4969 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5915) );
  NOR2_X1 U4970 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n5917) );
  INV_X1 U4971 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n6082) );
  INV_X1 U4972 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n6135) );
  INV_X1 U4973 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n6134) );
  INV_X1 U4974 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n6133) );
  NOR2_X1 U4975 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n5921) );
  INV_X4 U4976 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  AOI21_X2 U4977 ( .B1(n7573), .B2(n7574), .A(n7467), .ZN(n7470) );
  AOI211_X2 U4978 ( .C1(n9297), .C2(n9296), .A(n9295), .B(n9414), .ZN(n9438)
         );
  AOI21_X2 U4979 ( .B1(n5659), .B2(n9698), .A(n5658), .ZN(n8170) );
  AOI21_X2 U4980 ( .B1(n8880), .B2(n8869), .A(n8870), .ZN(n8868) );
  NAND2_X4 U4981 ( .A1(n5654), .A2(n9878), .ZN(n5013) );
  XNOR2_X2 U4982 ( .A(n4946), .B(n4945), .ZN(n9878) );
  XNOR2_X2 U4983 ( .A(n4943), .B(P1_IR_REG_27__SCAN_IN), .ZN(n5654) );
  INV_X4 U4984 ( .A(n5724), .ZN(n5780) );
  OAI21_X2 U4985 ( .B1(n5577), .B2(n4857), .A(n4855), .ZN(n9652) );
  AND2_X4 U4986 ( .A1(n8181), .A2(n5936), .ZN(n5983) );
  OAI211_X2 U4987 ( .C1(n5052), .C2(n6452), .A(n4951), .B(n4950), .ZN(n5672)
         );
  OR2_X1 U4988 ( .A1(n4984), .A2(n9470), .ZN(n4939) );
  NAND2_X2 U4989 ( .A1(n9848), .A2(n9851), .ZN(n4984) );
  OR2_X1 U4990 ( .A1(n9010), .A2(n8844), .ZN(n8405) );
  NAND2_X1 U4991 ( .A1(n5365), .A2(n5364), .ZN(n5377) );
  XNOR2_X1 U4992 ( .A(n8709), .B(n8728), .ZN(n8703) );
  AND2_X1 U4993 ( .A1(n4572), .A2(n4571), .ZN(n4570) );
  NAND2_X1 U4994 ( .A1(n9228), .A2(n9349), .ZN(n4571) );
  AND2_X1 U4995 ( .A1(n9399), .A2(n9348), .ZN(n4572) );
  NAND2_X1 U4996 ( .A1(n8525), .A2(n8510), .ZN(n4497) );
  NAND2_X1 U4997 ( .A1(n9260), .A2(n9261), .ZN(n4580) );
  NOR2_X1 U4998 ( .A1(n6328), .A2(n4665), .ZN(n4664) );
  INV_X1 U4999 ( .A(n6327), .ZN(n4665) );
  AND2_X1 U5000 ( .A1(n4803), .A2(n4802), .ZN(n4801) );
  NOR2_X1 U5001 ( .A1(n5403), .A2(n4807), .ZN(n4806) );
  INV_X1 U5002 ( .A(n4809), .ZN(n4807) );
  OAI21_X1 U5003 ( .B1(n4831), .B2(n4830), .A(n5296), .ZN(n4828) );
  AND2_X1 U5004 ( .A1(n5188), .A2(n5187), .ZN(n5189) );
  XNOR2_X1 U5005 ( .A(n5158), .B(SI_10_), .ZN(n5157) );
  NAND2_X1 U5006 ( .A1(n5112), .A2(SI_9_), .ZN(n5156) );
  INV_X1 U5007 ( .A(n5090), .ZN(n4824) );
  OR2_X1 U5008 ( .A1(n8780), .A2(n8592), .ZN(n8570) );
  INV_X1 U5009 ( .A(n4645), .ZN(n4644) );
  OAI21_X1 U5010 ( .B1(n8516), .B2(n4646), .A(n6339), .ZN(n4645) );
  NOR2_X1 U5011 ( .A1(n6344), .A2(n4656), .ZN(n4655) );
  INV_X1 U5012 ( .A(n4659), .ZN(n4656) );
  AND2_X1 U5013 ( .A1(n9004), .A2(n8832), .ZN(n6344) );
  AND2_X1 U5014 ( .A1(n8404), .A2(n8827), .ZN(n8406) );
  AND2_X1 U5015 ( .A1(n4399), .A2(n5928), .ZN(n4675) );
  INV_X1 U5016 ( .A(n9080), .ZN(n4736) );
  NOR2_X1 U5017 ( .A1(n9580), .A2(n4714), .ZN(n4713) );
  INV_X1 U5018 ( .A(n5499), .ZN(n4714) );
  NAND2_X1 U5019 ( .A1(n4494), .A2(n4493), .ZN(n4492) );
  INV_X1 U5020 ( .A(n9568), .ZN(n4494) );
  NAND2_X1 U5021 ( .A1(n9696), .A2(n9695), .ZN(n5577) );
  NAND2_X1 U5022 ( .A1(n4385), .A2(n5231), .ZN(n4704) );
  AOI21_X1 U5023 ( .B1(n5559), .B2(n9337), .A(n4835), .ZN(n4839) );
  INV_X1 U5024 ( .A(n5560), .ZN(n4835) );
  OAI21_X1 U5025 ( .B1(n8175), .B2(n8174), .A(n8173), .ZN(n8357) );
  OR2_X1 U5026 ( .A1(n8172), .A2(n8171), .ZN(n8173) );
  XNOR2_X1 U5027 ( .A(n8172), .B(n8171), .ZN(n8175) );
  NAND2_X1 U5028 ( .A1(n5425), .A2(n5424), .ZN(n5440) );
  NAND2_X1 U5029 ( .A1(n4816), .A2(n4817), .ZN(n5363) );
  NAND2_X1 U5030 ( .A1(n4413), .A2(n5333), .ZN(n4817) );
  NAND2_X1 U5031 ( .A1(n5210), .A2(SI_12_), .ZN(n5211) );
  INV_X1 U5032 ( .A(n5208), .ZN(n5212) );
  NOR2_X1 U5033 ( .A1(n7150), .A2(n6846), .ZN(n4888) );
  NAND2_X1 U5034 ( .A1(n8181), .A2(n8188), .ZN(n6256) );
  NAND2_X1 U5035 ( .A1(n6579), .A2(n6578), .ZN(n6776) );
  NOR2_X1 U5036 ( .A1(n7399), .A2(n7384), .ZN(n7521) );
  OR2_X1 U5037 ( .A1(n7504), .A2(n7503), .ZN(n7600) );
  NOR2_X1 U5038 ( .A1(n8675), .A2(n8665), .ZN(n4783) );
  INV_X1 U5039 ( .A(n8541), .ZN(n4618) );
  NAND2_X1 U5040 ( .A1(n7213), .A2(n8462), .ZN(n4632) );
  NAND2_X1 U5041 ( .A1(n8364), .A2(n8363), .ZN(n8575) );
  INV_X1 U5042 ( .A(n8832), .ZN(n8805) );
  NAND2_X1 U5043 ( .A1(n9017), .A2(n8859), .ZN(n4424) );
  NAND2_X1 U5044 ( .A1(n8841), .A2(n6341), .ZN(n4425) );
  OR2_X1 U5045 ( .A1(n8238), .A2(n8859), .ZN(n8826) );
  NAND2_X1 U5046 ( .A1(n6186), .A2(n6185), .ZN(n8954) );
  NAND2_X1 U5047 ( .A1(n7862), .A2(n6337), .ZN(n7913) );
  OR2_X1 U5048 ( .A1(n6397), .A2(n8578), .ZN(n8895) );
  OR2_X1 U5049 ( .A1(n4984), .A2(n4952), .ZN(n4854) );
  OAI21_X1 U5050 ( .B1(n9891), .B2(n7193), .A(n4440), .ZN(n9890) );
  NAND2_X1 U5051 ( .A1(n9891), .A2(n7193), .ZN(n4440) );
  NOR2_X1 U5052 ( .A1(n9741), .A2(n8194), .ZN(n9554) );
  INV_X1 U5053 ( .A(n9407), .ZN(n4715) );
  AND2_X1 U5054 ( .A1(n9324), .A2(n9316), .ZN(n9407) );
  OR2_X1 U5055 ( .A1(n9583), .A2(n9444), .ZN(n4716) );
  INV_X1 U5056 ( .A(n9593), .ZN(n5498) );
  NOR2_X1 U5057 ( .A1(n5456), .A2(n4684), .ZN(n4683) );
  INV_X1 U5058 ( .A(n4685), .ZN(n4684) );
  OR2_X1 U5059 ( .A1(n9624), .A2(n9086), .ZN(n9301) );
  NOR2_X1 U5060 ( .A1(n4706), .A2(n4389), .ZN(n4705) );
  NAND2_X1 U5061 ( .A1(n5467), .A2(n5466), .ZN(n9611) );
  AND4_X1 U5062 ( .A1(n4917), .A2(n4916), .A3(n4915), .A4(n4914), .ZN(n4918)
         );
  XNOR2_X1 U5063 ( .A(n5641), .B(n5640), .ZN(n7963) );
  NAND2_X1 U5064 ( .A1(n5524), .A2(n5523), .ZN(n5641) );
  NAND2_X1 U5065 ( .A1(n4876), .A2(n4877), .ZN(n7929) );
  AOI21_X1 U5066 ( .B1(n4880), .B2(n7724), .A(n4344), .ZN(n4877) );
  NAND2_X1 U5067 ( .A1(n8310), .A2(n8214), .ZN(n8264) );
  INV_X1 U5068 ( .A(n8788), .ZN(n8806) );
  INV_X1 U5069 ( .A(n8450), .ZN(n4521) );
  NAND2_X1 U5070 ( .A1(n4523), .A2(n8469), .ZN(n4518) );
  INV_X1 U5071 ( .A(n8418), .ZN(n4523) );
  NAND2_X1 U5072 ( .A1(n8496), .A2(n4365), .ZN(n4517) );
  AND2_X1 U5073 ( .A1(n4498), .A2(n8504), .ZN(n8525) );
  NAND2_X1 U5074 ( .A1(n8503), .A2(n4499), .ZN(n4498) );
  AOI21_X1 U5075 ( .B1(n4567), .B2(n4569), .A(n4844), .ZN(n4566) );
  INV_X1 U5076 ( .A(n4570), .ZN(n4569) );
  NOR2_X1 U5077 ( .A1(n4532), .A2(n4531), .ZN(n4530) );
  NAND2_X1 U5078 ( .A1(n8531), .A2(n8552), .ZN(n4531) );
  INV_X1 U5079 ( .A(n8827), .ZN(n4532) );
  AND2_X1 U5080 ( .A1(n8535), .A2(n8567), .ZN(n4533) );
  NOR2_X1 U5081 ( .A1(n4526), .A2(n4525), .ZN(n4524) );
  OAI22_X1 U5082 ( .A1(n4343), .A2(n4528), .B1(n4379), .B2(n4527), .ZN(n4526)
         );
  INV_X1 U5083 ( .A(n8536), .ZN(n4525) );
  INV_X1 U5084 ( .A(n4533), .ZN(n4527) );
  NOR2_X1 U5085 ( .A1(n4530), .A2(n4533), .ZN(n4529) );
  INV_X1 U5086 ( .A(n9653), .ZN(n4579) );
  INV_X1 U5087 ( .A(n9324), .ZN(n4562) );
  AOI21_X1 U5088 ( .B1(n4338), .B2(n4577), .A(n4575), .ZN(n4574) );
  NAND2_X1 U5089 ( .A1(n9316), .A2(n9278), .ZN(n4557) );
  INV_X1 U5090 ( .A(n4814), .ZN(n4813) );
  OAI21_X1 U5091 ( .B1(n5511), .B2(n4815), .A(n5640), .ZN(n4814) );
  INV_X1 U5092 ( .A(n5523), .ZN(n4815) );
  INV_X1 U5093 ( .A(n4460), .ZN(n4459) );
  NAND2_X1 U5094 ( .A1(n5457), .A2(n4791), .ZN(n4790) );
  INV_X1 U5095 ( .A(n5439), .ZN(n4791) );
  INV_X1 U5096 ( .A(n4832), .ZN(n4831) );
  OAI21_X1 U5097 ( .B1(n5279), .B2(n4833), .A(n5258), .ZN(n4832) );
  INV_X1 U5098 ( .A(SI_15_), .ZN(n4833) );
  NAND2_X1 U5099 ( .A1(n4587), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n4586) );
  NOR2_X1 U5100 ( .A1(n4781), .A2(n6777), .ZN(n4780) );
  OR2_X1 U5101 ( .A1(n4607), .A2(n4605), .ZN(n4597) );
  NAND2_X1 U5102 ( .A1(n7615), .A2(n7614), .ZN(n7749) );
  INV_X1 U5103 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n6150) );
  INV_X1 U5104 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n6163) );
  OR2_X1 U5105 ( .A1(n8985), .A2(n8551), .ZN(n8253) );
  AOI21_X1 U5106 ( .B1(n4664), .B2(n6326), .A(n4380), .ZN(n4663) );
  OR2_X1 U5107 ( .A1(n6075), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6087) );
  OR2_X1 U5108 ( .A1(n6050), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n6065) );
  NAND2_X1 U5109 ( .A1(n10072), .A2(n8607), .ZN(n8456) );
  NAND2_X1 U5110 ( .A1(n4439), .A2(n4438), .ZN(n8428) );
  INV_X1 U5111 ( .A(n8547), .ZN(n4612) );
  OR2_X1 U5112 ( .A1(n8991), .A2(n8806), .ZN(n8548) );
  OR2_X1 U5113 ( .A1(n8998), .A2(n6346), .ZN(n8545) );
  OR2_X1 U5114 ( .A1(n9020), .A2(n8843), .ZN(n8535) );
  NOR2_X1 U5115 ( .A1(n6200), .A2(n4630), .ZN(n4629) );
  OR2_X1 U5116 ( .A1(n9026), .A2(n8857), .ZN(n8530) );
  OR2_X1 U5117 ( .A1(n9032), .A2(n8268), .ZN(n8408) );
  INV_X1 U5118 ( .A(n8520), .ZN(n4637) );
  OR2_X1 U5119 ( .A1(n8959), .A2(n8298), .ZN(n8521) );
  OR2_X1 U5120 ( .A1(n8289), .A2(n8283), .ZN(n8520) );
  INV_X1 U5121 ( .A(n8513), .ZN(n4638) );
  INV_X1 U5122 ( .A(n4663), .ZN(n4661) );
  OR2_X1 U5123 ( .A1(n8488), .A2(n8597), .ZN(n6330) );
  AND2_X1 U5124 ( .A1(n5927), .A2(n6293), .ZN(n5928) );
  INV_X1 U5125 ( .A(n7238), .ZN(n4734) );
  NOR2_X1 U5126 ( .A1(n4758), .A2(n9175), .ZN(n4757) );
  INV_X1 U5127 ( .A(n4759), .ZN(n4758) );
  XNOR2_X1 U5128 ( .A(n5714), .B(n5874), .ZN(n5716) );
  NAND2_X1 U5129 ( .A1(n4732), .A2(n5744), .ZN(n4730) );
  INV_X1 U5130 ( .A(n9093), .ZN(n4752) );
  AND2_X1 U5131 ( .A1(n4753), .A2(n4752), .ZN(n4751) );
  NAND2_X1 U5132 ( .A1(n7162), .A2(n7167), .ZN(n5733) );
  NAND2_X1 U5133 ( .A1(n7161), .A2(n4363), .ZN(n5734) );
  OR2_X1 U5134 ( .A1(n8164), .A2(n5648), .ZN(n9327) );
  OR2_X1 U5135 ( .A1(n5448), .A2(n9152), .ZN(n5468) );
  NOR2_X1 U5136 ( .A1(n7766), .A2(n4848), .ZN(n4847) );
  INV_X1 U5137 ( .A(n4703), .ZN(n4702) );
  OAI21_X1 U5138 ( .B1(n4704), .B2(n9396), .A(n5251), .ZN(n4703) );
  NOR2_X1 U5139 ( .A1(n7773), .A2(n9076), .ZN(n4488) );
  OR2_X1 U5140 ( .A1(n10017), .A2(n5127), .ZN(n9214) );
  AND2_X1 U5141 ( .A1(n7174), .A2(n9383), .ZN(n4694) );
  INV_X1 U5142 ( .A(n5045), .ZN(n4696) );
  NAND2_X1 U5143 ( .A1(n9376), .A2(n9296), .ZN(n5675) );
  NAND2_X1 U5144 ( .A1(n5502), .A2(n5501), .ZN(n5504) );
  NAND2_X1 U5145 ( .A1(n5512), .A2(n5511), .ZN(n5524) );
  NAND2_X1 U5146 ( .A1(n4800), .A2(n4797), .ZN(n5425) );
  AOI21_X1 U5147 ( .B1(n4799), .B2(n4803), .A(n4798), .ZN(n4797) );
  INV_X1 U5148 ( .A(n5415), .ZN(n4798) );
  NOR2_X1 U5149 ( .A1(n5233), .A2(n8067), .ZN(n5235) );
  INV_X1 U5150 ( .A(n5232), .ZN(n5233) );
  XNOR2_X1 U5151 ( .A(n5209), .B(SI_12_), .ZN(n5208) );
  AND2_X1 U5152 ( .A1(n5184), .A2(n5185), .ZN(n5191) );
  NOR2_X1 U5153 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n4913) );
  NAND2_X1 U5154 ( .A1(n8253), .A2(n8252), .ZN(n8375) );
  INV_X1 U5155 ( .A(n8602), .ZN(n7474) );
  NAND2_X1 U5156 ( .A1(n4879), .A2(n4878), .ZN(n4881) );
  INV_X1 U5157 ( .A(n7725), .ZN(n4879) );
  OR2_X1 U5158 ( .A1(n7715), .A2(n7716), .ZN(n4865) );
  NOR2_X1 U5159 ( .A1(n4893), .A2(n7152), .ZN(n4890) );
  AND2_X1 U5160 ( .A1(n8580), .A2(n4794), .ZN(n4793) );
  NAND2_X1 U5161 ( .A1(n4795), .A2(n4360), .ZN(n4794) );
  INV_X1 U5162 ( .A(n8581), .ZN(n4795) );
  AND2_X1 U5163 ( .A1(n7410), .A2(n7409), .ZN(n8769) );
  NAND2_X1 U5164 ( .A1(n4588), .A2(n6611), .ZN(n4587) );
  INV_X1 U5165 ( .A(n6587), .ZN(n4588) );
  NAND2_X1 U5166 ( .A1(n4601), .A2(n4607), .ZN(n4600) );
  OR2_X1 U5167 ( .A1(n6770), .A2(n10140), .ZN(n6824) );
  NAND2_X1 U5168 ( .A1(n4603), .A2(n4337), .ZN(n4602) );
  NAND2_X1 U5169 ( .A1(n6776), .A2(n6775), .ZN(n4770) );
  NAND2_X1 U5170 ( .A1(n4775), .A2(n4772), .ZN(n4771) );
  NOR2_X1 U5171 ( .A1(n6777), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n4776) );
  OR2_X1 U5172 ( .A1(n4778), .A2(n4777), .ZN(n6819) );
  NAND2_X1 U5173 ( .A1(n4779), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n4778) );
  INV_X1 U5174 ( .A(n6817), .ZN(n4777) );
  AOI21_X1 U5175 ( .B1(P2_REG2_REG_8__SCAN_IN), .B2(n7004), .A(n8633), .ZN(
        n7075) );
  OR2_X1 U5176 ( .A1(n7065), .A2(n7064), .ZN(n7381) );
  OR2_X1 U5177 ( .A1(n7521), .A2(n7520), .ZN(n4768) );
  NAND2_X1 U5178 ( .A1(n4768), .A2(n4767), .ZN(n7615) );
  INV_X1 U5179 ( .A(n7523), .ZN(n4767) );
  XNOR2_X1 U5180 ( .A(n7749), .B(n7616), .ZN(n7617) );
  NOR2_X1 U5181 ( .A1(n7604), .A2(n7617), .ZN(n7752) );
  OR2_X1 U5182 ( .A1(n8653), .A2(n7844), .ZN(n4769) );
  OR2_X1 U5183 ( .A1(n6252), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6262) );
  AND2_X1 U5184 ( .A1(n8544), .A2(n8545), .ZN(n8808) );
  OR2_X1 U5185 ( .A1(n9020), .A2(n8873), .ZN(n4422) );
  OR2_X1 U5186 ( .A1(n6203), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n6211) );
  AOI21_X1 U5187 ( .B1(n4644), .B2(n4646), .A(n4373), .ZN(n4642) );
  NAND2_X1 U5188 ( .A1(n6115), .A2(n6114), .ZN(n6126) );
  INV_X1 U5189 ( .A(n6116), .ZN(n6115) );
  OR2_X1 U5190 ( .A1(n6087), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6099) );
  AND4_X1 U5191 ( .A1(n6071), .A2(n6070), .A3(n6069), .A4(n6068), .ZN(n7717)
         );
  OR2_X1 U5192 ( .A1(n7468), .A2(n7716), .ZN(n8417) );
  NAND2_X1 U5193 ( .A1(n6057), .A2(n6056), .ZN(n7136) );
  AND2_X1 U5194 ( .A1(n8448), .A2(n8445), .ZN(n4631) );
  NAND2_X1 U5195 ( .A1(n7096), .A2(n8459), .ZN(n7213) );
  INV_X1 U5196 ( .A(n8375), .ZN(n8786) );
  NAND2_X1 U5197 ( .A1(n8789), .A2(n8899), .ZN(n4672) );
  AND2_X1 U5198 ( .A1(n8548), .A2(n8547), .ZN(n8794) );
  INV_X1 U5199 ( .A(n4615), .ZN(n4614) );
  OAI21_X1 U5200 ( .B1(n4351), .B2(n4330), .A(n8545), .ZN(n4615) );
  NAND2_X1 U5201 ( .A1(n4655), .A2(n6342), .ZN(n4654) );
  AND2_X1 U5202 ( .A1(n6237), .A2(n8405), .ZN(n8403) );
  OR2_X1 U5203 ( .A1(n6236), .A2(n8826), .ZN(n6237) );
  NAND2_X1 U5204 ( .A1(n9010), .A2(n8816), .ZN(n4659) );
  AOI21_X1 U5205 ( .B1(n4629), .B2(n8904), .A(n4627), .ZN(n4626) );
  INV_X1 U5206 ( .A(n8508), .ZN(n4627) );
  INV_X1 U5207 ( .A(n4629), .ZN(n4628) );
  AND2_X1 U5208 ( .A1(n8530), .A2(n8532), .ZN(n8870) );
  NAND2_X1 U5209 ( .A1(n8903), .A2(n8893), .ZN(n8952) );
  NAND2_X1 U5210 ( .A1(n7913), .A2(n8516), .ZN(n7915) );
  OR2_X1 U5211 ( .A1(n4640), .A2(n4336), .ZN(n7867) );
  OR2_X1 U5212 ( .A1(n7836), .A2(n8501), .ZN(n7834) );
  INV_X1 U5213 ( .A(n8858), .ZN(n8898) );
  OR2_X1 U5214 ( .A1(n6940), .A2(n8588), .ZN(n10116) );
  INV_X1 U5215 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5916) );
  NAND2_X1 U5216 ( .A1(n4734), .A2(n4733), .ZN(n4732) );
  INV_X1 U5217 ( .A(n7239), .ZN(n4733) );
  NAND2_X1 U5218 ( .A1(n4361), .A2(n5734), .ZN(n4731) );
  AOI21_X1 U5219 ( .B1(n9079), .B2(n9167), .A(n4736), .ZN(n4735) );
  NAND2_X1 U5220 ( .A1(n4350), .A2(n5754), .ZN(n4447) );
  NAND2_X1 U5221 ( .A1(n4350), .A2(n4449), .ZN(n4448) );
  INV_X1 U5222 ( .A(n7537), .ZN(n4449) );
  AOI21_X1 U5223 ( .B1(n4757), .B2(n4755), .A(n4754), .ZN(n4753) );
  INV_X1 U5224 ( .A(n9176), .ZN(n4754) );
  INV_X1 U5225 ( .A(n5803), .ZN(n4755) );
  INV_X1 U5226 ( .A(n4757), .ZN(n4756) );
  AND2_X2 U5227 ( .A1(n5675), .A2(n5671), .ZN(n5874) );
  AOI21_X1 U5228 ( .B1(n6695), .B2(n5780), .A(n4902), .ZN(n5689) );
  XOR2_X1 U5229 ( .A(n5869), .B(n5868), .Z(n9115) );
  NAND2_X1 U5230 ( .A1(n5844), .A2(n5845), .ZN(n9143) );
  NAND2_X1 U5231 ( .A1(n9083), .A2(n9143), .ZN(n5859) );
  AND2_X1 U5232 ( .A1(n9115), .A2(n4741), .ZN(n4740) );
  NAND2_X1 U5233 ( .A1(n4742), .A2(n5860), .ZN(n4741) );
  INV_X1 U5234 ( .A(n9144), .ZN(n4742) );
  AND2_X1 U5235 ( .A1(n9282), .A2(n9202), .ZN(n9417) );
  AND2_X1 U5236 ( .A1(n9806), .A2(n9425), .ZN(n9427) );
  INV_X1 U5237 ( .A(n4979), .ZN(n5290) );
  OR2_X1 U5238 ( .A1(n4984), .A2(n7322), .ZN(n5010) );
  AND2_X1 U5239 ( .A1(n4477), .A2(n4476), .ZN(n9905) );
  NAND2_X1 U5240 ( .A1(n8182), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n4476) );
  NOR2_X1 U5241 ( .A1(n9482), .A2(n4415), .ZN(n9506) );
  NAND2_X1 U5242 ( .A1(n4919), .A2(n4765), .ZN(n4764) );
  AND2_X1 U5243 ( .A1(n9926), .A2(n9509), .ZN(n9510) );
  INV_X1 U5244 ( .A(n9411), .ZN(n9277) );
  INV_X1 U5245 ( .A(n4713), .ZN(n4709) );
  AND2_X1 U5246 ( .A1(n9327), .A2(n9366), .ZN(n9411) );
  NAND2_X1 U5247 ( .A1(n9575), .A2(n9315), .ZN(n5639) );
  AOI21_X1 U5248 ( .B1(n4353), .B2(n4683), .A(n4682), .ZN(n4681) );
  INV_X1 U5249 ( .A(n9261), .ZN(n4682) );
  OR2_X1 U5250 ( .A1(n9824), .A2(n9448), .ZN(n4685) );
  NAND2_X1 U5251 ( .A1(n5579), .A2(n4341), .ZN(n9620) );
  NAND2_X1 U5252 ( .A1(n4719), .A2(n4717), .ZN(n9665) );
  AOI21_X1 U5253 ( .B1(n9680), .B2(n5373), .A(n4718), .ZN(n4717) );
  NAND2_X1 U5254 ( .A1(n9690), .A2(n9781), .ZN(n9682) );
  NAND2_X1 U5255 ( .A1(n5577), .A2(n4860), .ZN(n9678) );
  NAND2_X1 U5256 ( .A1(n5575), .A2(n9241), .ZN(n9696) );
  OR2_X1 U5257 ( .A1(n9706), .A2(n9703), .ZN(n5575) );
  OR2_X1 U5258 ( .A1(n9711), .A2(n9793), .ZN(n9709) );
  NAND2_X1 U5259 ( .A1(n9704), .A2(n5328), .ZN(n4707) );
  AND2_X1 U5260 ( .A1(n9239), .A2(n9363), .ZN(n9695) );
  NAND2_X1 U5261 ( .A1(n4842), .A2(n4840), .ZN(n7883) );
  NOR2_X1 U5262 ( .A1(n5294), .A2(n4841), .ZN(n4840) );
  INV_X1 U5263 ( .A(n4843), .ZN(n4841) );
  OR2_X2 U5264 ( .A1(n7691), .A2(n4846), .ZN(n4842) );
  INV_X1 U5265 ( .A(n4847), .ZN(n4846) );
  AOI21_X1 U5266 ( .B1(n4847), .B2(n4845), .A(n4844), .ZN(n4843) );
  NAND2_X1 U5267 ( .A1(n7691), .A2(n9399), .ZN(n7695) );
  AND2_X1 U5268 ( .A1(n9223), .A2(n9221), .ZN(n9394) );
  NAND2_X1 U5269 ( .A1(n9346), .A2(n7334), .ZN(n4849) );
  NOR2_X1 U5270 ( .A1(n7553), .A2(n7979), .ZN(n7633) );
  OR2_X1 U5271 ( .A1(n7444), .A2(n7802), .ZN(n7553) );
  AOI21_X1 U5272 ( .B1(n7334), .B2(n4691), .A(n4382), .ZN(n4690) );
  INV_X1 U5273 ( .A(n5128), .ZN(n4691) );
  INV_X1 U5274 ( .A(n4839), .ZN(n4583) );
  INV_X1 U5275 ( .A(n9338), .ZN(n4837) );
  NAND2_X1 U5276 ( .A1(n5026), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5059) );
  NAND2_X1 U5277 ( .A1(n5550), .A2(n7182), .ZN(n7037) );
  AND2_X1 U5278 ( .A1(n5628), .A2(n9842), .ZN(n5890) );
  NAND2_X1 U5279 ( .A1(n5447), .A2(n5446), .ZN(n9624) );
  INV_X1 U5280 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n4928) );
  INV_X1 U5281 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n4919) );
  XNOR2_X1 U5282 ( .A(n8361), .B(n8360), .ZN(n9199) );
  NAND2_X1 U5283 ( .A1(n9843), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4930) );
  XNOR2_X1 U5284 ( .A(n8357), .B(n8356), .ZN(n8366) );
  XNOR2_X1 U5285 ( .A(n5464), .B(n5463), .ZN(n7798) );
  NAND2_X1 U5286 ( .A1(n5458), .A2(n5457), .ZN(n5481) );
  OAI21_X1 U5287 ( .B1(n5377), .B2(n4805), .A(n4803), .ZN(n5417) );
  NAND2_X1 U5288 ( .A1(n4808), .A2(n4809), .ZN(n5404) );
  NAND2_X1 U5289 ( .A1(n5377), .A2(n4810), .ZN(n4808) );
  NAND2_X1 U5290 ( .A1(n5321), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5341) );
  INV_X1 U5291 ( .A(n5363), .ZN(n5360) );
  NAND2_X1 U5292 ( .A1(n5301), .A2(n5302), .ZN(n5318) );
  NAND2_X1 U5293 ( .A1(n5259), .A2(n5258), .ZN(n5277) );
  XNOR2_X1 U5294 ( .A(n5138), .B(n5137), .ZN(n6480) );
  OAI21_X1 U5295 ( .B1(n5113), .B2(n4507), .A(n4502), .ZN(n4501) );
  AND2_X1 U5296 ( .A1(n4834), .A2(n4973), .ZN(n5014) );
  INV_X1 U5297 ( .A(n4998), .ZN(n4469) );
  AOI21_X1 U5298 ( .B1(n8331), .B2(n8332), .A(n4433), .ZN(n8243) );
  AND2_X1 U5299 ( .A1(n8208), .A2(n8298), .ZN(n4433) );
  INV_X1 U5300 ( .A(n4881), .ZN(n7819) );
  AND2_X1 U5301 ( .A1(n6235), .A2(n6234), .ZN(n8859) );
  AND2_X1 U5302 ( .A1(n8215), .A2(n8857), .ZN(n4432) );
  NAND2_X1 U5303 ( .A1(n8206), .A2(n8283), .ZN(n4434) );
  AOI21_X1 U5304 ( .B1(n4873), .B2(n4875), .A(n4408), .ZN(n4870) );
  AND2_X1 U5305 ( .A1(n7926), .A2(n7927), .ZN(n4431) );
  NAND2_X1 U5306 ( .A1(n6268), .A2(n6267), .ZN(n8788) );
  OAI211_X1 U5307 ( .C1(n7600), .C2(n7751), .A(n4608), .B(n4419), .ZN(n7601)
         );
  NAND2_X1 U5308 ( .A1(n7600), .A2(n4417), .ZN(n4608) );
  INV_X1 U5309 ( .A(n7599), .ZN(n4609) );
  NOR2_X1 U5310 ( .A1(n7601), .A2(n7668), .ZN(n7729) );
  AND2_X1 U5311 ( .A1(n4368), .A2(n4782), .ZN(n8712) );
  INV_X1 U5312 ( .A(n4437), .ZN(n4423) );
  AOI21_X1 U5313 ( .B1(n8782), .B2(n7217), .A(n6365), .ZN(n4437) );
  NAND2_X1 U5314 ( .A1(n6141), .A2(n6140), .ZN(n8966) );
  OR2_X1 U5315 ( .A1(n5013), .A2(n6637), .ZN(n4950) );
  NAND2_X1 U5316 ( .A1(n6426), .A2(n4451), .ZN(n4450) );
  NAND2_X1 U5317 ( .A1(n9147), .A2(n4452), .ZN(n4451) );
  NOR2_X1 U5318 ( .A1(n9115), .A2(n4743), .ZN(n4452) );
  INV_X1 U5319 ( .A(n9186), .ZN(n9863) );
  AND2_X1 U5320 ( .A1(n5899), .A2(n5893), .ZN(n9865) );
  INV_X1 U5321 ( .A(n9183), .ZN(n9861) );
  NOR2_X1 U5322 ( .A1(n9887), .A2(n4359), .ZN(n6680) );
  AND2_X1 U5323 ( .A1(n9884), .A2(n4478), .ZN(n6684) );
  NAND2_X1 U5324 ( .A1(n9891), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n4478) );
  NOR2_X1 U5325 ( .A1(n6655), .A2(n4407), .ZN(n6646) );
  NOR2_X1 U5326 ( .A1(n6801), .A2(n6800), .ZN(n6881) );
  NOR2_X1 U5327 ( .A1(n9555), .A2(n9977), .ZN(n9736) );
  OR2_X1 U5328 ( .A1(n9554), .A2(n8196), .ZN(n9563) );
  NAND2_X1 U5329 ( .A1(n5661), .A2(n5536), .ZN(n9564) );
  NAND2_X1 U5330 ( .A1(n4712), .A2(n4710), .ZN(n5661) );
  NAND2_X1 U5331 ( .A1(n4712), .A2(n4716), .ZN(n5535) );
  INV_X1 U5332 ( .A(n9720), .ZN(n9721) );
  NAND2_X1 U5333 ( .A1(n5526), .A2(n5525), .ZN(n9568) );
  NAND2_X1 U5334 ( .A1(n7963), .A2(n5114), .ZN(n5526) );
  AND2_X1 U5335 ( .A1(n10049), .A2(n9993), .ZN(n9832) );
  NAND2_X1 U5336 ( .A1(n4522), .A2(n4519), .ZN(n8469) );
  NAND2_X1 U5337 ( .A1(n8452), .A2(n4520), .ZN(n4519) );
  NOR2_X1 U5338 ( .A1(n8567), .A2(n4521), .ZN(n4520) );
  NAND2_X1 U5339 ( .A1(n4553), .A2(n4552), .ZN(n4551) );
  AOI21_X1 U5340 ( .B1(n4516), .B2(n8495), .A(n6335), .ZN(n4515) );
  AND2_X1 U5341 ( .A1(n4517), .A2(n8500), .ZN(n4516) );
  AND2_X1 U5342 ( .A1(n8512), .A2(n8552), .ZN(n4499) );
  AOI21_X1 U5343 ( .B1(n4570), .B2(n4568), .A(n4391), .ZN(n4567) );
  INV_X1 U5344 ( .A(n9228), .ZN(n4568) );
  INV_X1 U5345 ( .A(n4530), .ZN(n4528) );
  NAND2_X1 U5346 ( .A1(n4496), .A2(n4495), .ZN(n8527) );
  NAND2_X1 U5347 ( .A1(n8511), .A2(n8552), .ZN(n4495) );
  NAND2_X1 U5348 ( .A1(n4497), .A2(n4367), .ZN(n4496) );
  NOR2_X1 U5349 ( .A1(n9237), .A2(n9236), .ZN(n4549) );
  OAI21_X1 U5350 ( .B1(n8543), .B2(n8542), .A(n8808), .ZN(n4513) );
  NAND2_X1 U5351 ( .A1(n4393), .A2(n4580), .ZN(n4576) );
  NOR2_X1 U5352 ( .A1(n9259), .A2(n9619), .ZN(n4581) );
  NAND2_X1 U5353 ( .A1(n4582), .A2(n4579), .ZN(n4578) );
  NAND2_X1 U5354 ( .A1(n4582), .A2(n4580), .ZN(n4577) );
  INV_X1 U5355 ( .A(n9265), .ZN(n4575) );
  NAND2_X1 U5356 ( .A1(n4512), .A2(n4510), .ZN(n8561) );
  NOR2_X1 U5357 ( .A1(n8558), .A2(n4511), .ZN(n4510) );
  NAND2_X1 U5358 ( .A1(n4513), .A2(n4370), .ZN(n4512) );
  INV_X1 U5359 ( .A(n8549), .ZN(n4511) );
  INV_X1 U5360 ( .A(n5416), .ZN(n4802) );
  NAND2_X1 U5361 ( .A1(n4462), .A2(n4461), .ZN(n4460) );
  INV_X1 U5362 ( .A(n9070), .ZN(n4461) );
  NAND2_X1 U5363 ( .A1(n9275), .A2(n4561), .ZN(n4560) );
  NAND2_X1 U5364 ( .A1(n4562), .A2(n9278), .ZN(n4561) );
  NAND2_X1 U5365 ( .A1(n4564), .A2(n4339), .ZN(n4563) );
  NOR2_X1 U5366 ( .A1(n9268), .A2(n4557), .ZN(n4556) );
  NAND2_X1 U5367 ( .A1(n9269), .A2(n9325), .ZN(n4558) );
  NOR2_X1 U5368 ( .A1(n7890), .A2(n4487), .ZN(n4486) );
  INV_X1 U5369 ( .A(n4488), .ZN(n4487) );
  NAND2_X1 U5370 ( .A1(n4812), .A2(n4811), .ZN(n8172) );
  AOI21_X1 U5371 ( .B1(n4813), .B2(n4815), .A(n4418), .ZN(n4811) );
  AND2_X1 U5372 ( .A1(n4805), .A2(n4802), .ZN(n4799) );
  INV_X1 U5373 ( .A(n5316), .ZN(n4819) );
  AND2_X1 U5374 ( .A1(n4820), .A2(n5333), .ZN(n4818) );
  NAND2_X1 U5375 ( .A1(n5164), .A2(n5163), .ZN(n5185) );
  NAND2_X1 U5376 ( .A1(n5093), .A2(n5092), .ZN(n5133) );
  INV_X1 U5377 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4540) );
  OR2_X1 U5378 ( .A1(n8571), .A2(n8374), .ZN(n8574) );
  NAND2_X1 U5379 ( .A1(n6576), .A2(n6586), .ZN(n6577) );
  NAND2_X1 U5380 ( .A1(n4774), .A2(n4773), .ZN(n4772) );
  NAND2_X1 U5381 ( .A1(n4781), .A2(n6777), .ZN(n4773) );
  OR2_X1 U5382 ( .A1(n4780), .A2(n6778), .ZN(n4774) );
  INV_X1 U5383 ( .A(n6818), .ZN(n4775) );
  NAND2_X1 U5384 ( .A1(n7397), .A2(n7396), .ZN(n7517) );
  INV_X1 U5385 ( .A(n6338), .ZN(n4646) );
  NAND2_X1 U5386 ( .A1(n6064), .A2(n7083), .ZN(n6075) );
  INV_X1 U5387 ( .A(n6065), .ZN(n6064) );
  NAND2_X1 U5388 ( .A1(n6037), .A2(n6036), .ZN(n6050) );
  INV_X1 U5389 ( .A(n6038), .ZN(n6037) );
  NAND2_X1 U5390 ( .A1(n7108), .A2(n6844), .ZN(n8441) );
  NAND2_X1 U5391 ( .A1(n4867), .A2(n4866), .ZN(n6379) );
  AND2_X1 U5392 ( .A1(n8998), .A2(n6346), .ZN(n8376) );
  INV_X1 U5393 ( .A(n8760), .ZN(n6399) );
  INV_X1 U5394 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n6294) );
  INV_X1 U5395 ( .A(n5768), .ZN(n4745) );
  OR2_X1 U5396 ( .A1(n5831), .A2(n5830), .ZN(n5832) );
  AOI21_X1 U5397 ( .B1(n4458), .B2(n4746), .A(n4362), .ZN(n4456) );
  OR2_X1 U5398 ( .A1(n9568), .A2(n9272), .ZN(n9324) );
  NAND2_X1 U5399 ( .A1(n5489), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n5528) );
  INV_X1 U5400 ( .A(n9245), .ZN(n4859) );
  INV_X1 U5401 ( .A(n9247), .ZN(n4856) );
  NOR2_X1 U5402 ( .A1(n9831), .A2(n4484), .ZN(n4483) );
  INV_X1 U5403 ( .A(n5329), .ZN(n4706) );
  AOI21_X1 U5404 ( .B1(n4702), .B2(n4704), .A(n4701), .ZN(n4700) );
  OR2_X1 U5405 ( .A1(n7890), .A2(n5293), .ZN(n9353) );
  INV_X1 U5406 ( .A(n5175), .ZN(n5173) );
  NOR2_X1 U5407 ( .A1(n4688), .A2(n4689), .ZN(n4687) );
  INV_X1 U5408 ( .A(n9391), .ZN(n4689) );
  INV_X1 U5409 ( .A(n7360), .ZN(n7358) );
  NOR2_X1 U5410 ( .A1(n9204), .A2(n9946), .ZN(n7362) );
  AND3_X1 U5411 ( .A1(n7321), .A2(n4480), .A3(n4479), .ZN(n7370) );
  NOR2_X1 U5412 ( .A1(n7179), .A2(n9992), .ZN(n4480) );
  INV_X1 U5413 ( .A(n9337), .ZN(n4838) );
  INV_X1 U5414 ( .A(n9469), .ZN(n4957) );
  NOR2_X1 U5415 ( .A1(n9637), .A2(n9624), .ZN(n5590) );
  NAND2_X1 U5416 ( .A1(n7699), .A2(n4486), .ZN(n7945) );
  OAI22_X1 U5417 ( .A1(n5440), .A2(n4789), .B1(n4348), .B2(n5479), .ZN(n5502)
         );
  NAND2_X1 U5418 ( .A1(n5457), .A2(n5478), .ZN(n4789) );
  INV_X1 U5419 ( .A(n4806), .ZN(n4805) );
  AOI21_X1 U5420 ( .B1(n4804), .B2(n4806), .A(n4412), .ZN(n4803) );
  INV_X1 U5421 ( .A(n4810), .ZN(n4804) );
  NAND2_X1 U5422 ( .A1(n5604), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5548) );
  NAND2_X1 U5423 ( .A1(n5375), .A2(n5376), .ZN(n4809) );
  OR2_X1 U5424 ( .A1(n5375), .A2(n5376), .ZN(n4810) );
  NOR2_X1 U5425 ( .A1(n4764), .A2(P1_IR_REG_16__SCAN_IN), .ZN(n4763) );
  INV_X1 U5426 ( .A(n5317), .ZN(n4820) );
  INV_X1 U5427 ( .A(n4828), .ZN(n4827) );
  NAND2_X1 U5428 ( .A1(n4826), .A2(n4829), .ZN(n5297) );
  AND2_X1 U5429 ( .A1(n5160), .A2(n5159), .ZN(n5187) );
  OR2_X1 U5430 ( .A1(n5157), .A2(n5156), .ZN(n5160) );
  AND2_X1 U5431 ( .A1(n5155), .A2(n5137), .ZN(n5184) );
  NAND2_X1 U5432 ( .A1(n4825), .A2(n4823), .ZN(n5192) );
  AND2_X1 U5433 ( .A1(n5133), .A2(n5132), .ZN(n5155) );
  NAND2_X1 U5434 ( .A1(n4507), .A2(n4503), .ZN(n4502) );
  NAND2_X1 U5435 ( .A1(n4509), .A2(n4505), .ZN(n4503) );
  AOI21_X1 U5436 ( .B1(n4823), .B2(n5086), .A(n4508), .ZN(n4507) );
  INV_X1 U5437 ( .A(n5133), .ZN(n4508) );
  INV_X1 U5438 ( .A(n5113), .ZN(n4505) );
  NAND2_X1 U5439 ( .A1(n4823), .A2(n5113), .ZN(n4500) );
  OR2_X1 U5440 ( .A1(n5096), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n5142) );
  INV_X1 U5441 ( .A(n5066), .ZN(n5067) );
  XNOR2_X1 U5442 ( .A(n5069), .B(SI_6_), .ZN(n5066) );
  OAI21_X1 U5443 ( .B1(n4332), .B2(P1_DATAO_REG_1__SCAN_IN), .A(n4947), .ZN(
        n4968) );
  NAND2_X1 U5444 ( .A1(n4995), .A2(n6451), .ZN(n4947) );
  NOR2_X1 U5445 ( .A1(n8281), .A2(n4886), .ZN(n4885) );
  INV_X1 U5446 ( .A(n4887), .ZN(n4886) );
  INV_X1 U5447 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n6773) );
  NAND2_X1 U5448 ( .A1(n5995), .A2(n6773), .ZN(n6011) );
  INV_X1 U5449 ( .A(n6009), .ZN(n5995) );
  AND2_X1 U5450 ( .A1(n8273), .A2(n4874), .ZN(n4873) );
  OR2_X1 U5451 ( .A1(n8304), .A2(n4875), .ZN(n4874) );
  INV_X1 U5452 ( .A(n8225), .ZN(n4875) );
  AND2_X1 U5453 ( .A1(n7410), .A2(n6289), .ZN(n8592) );
  NAND4_X1 U5454 ( .A1(n5941), .A2(n5940), .A3(n5939), .A4(n5938), .ZN(n6299)
         );
  OR2_X1 U5455 ( .A1(n6285), .A2(n4641), .ZN(n5939) );
  NAND2_X1 U5456 ( .A1(n6577), .A2(n4436), .ZN(n6601) );
  OR2_X1 U5457 ( .A1(n6576), .A2(n6586), .ZN(n4436) );
  NAND2_X1 U5458 ( .A1(n4589), .A2(n6588), .ZN(n6768) );
  NAND2_X1 U5459 ( .A1(n4585), .A2(n6589), .ZN(n6604) );
  INV_X1 U5460 ( .A(n4586), .ZN(n4585) );
  NAND2_X1 U5461 ( .A1(n6776), .A2(n4780), .ZN(n4779) );
  AND2_X1 U5462 ( .A1(n6910), .A2(n6909), .ZN(n6911) );
  NAND2_X1 U5463 ( .A1(n4337), .A2(n4604), .ZN(n4599) );
  OAI21_X1 U5464 ( .B1(n4601), .B2(n4605), .A(n4596), .ZN(n4598) );
  AND2_X1 U5465 ( .A1(n4597), .A2(n4604), .ZN(n4596) );
  NAND2_X1 U5466 ( .A1(n6912), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n8626) );
  NOR2_X1 U5467 ( .A1(n7077), .A2(n7078), .ZN(n7080) );
  XNOR2_X1 U5468 ( .A(n7517), .B(n7398), .ZN(n7399) );
  AND2_X1 U5469 ( .A1(n7381), .A2(n7380), .ZN(n7498) );
  NOR2_X1 U5470 ( .A1(n7753), .A2(n7752), .ZN(n7756) );
  INV_X1 U5471 ( .A(n7749), .ZN(n7750) );
  INV_X1 U5472 ( .A(n8661), .ZN(n4595) );
  NAND2_X1 U5473 ( .A1(n6165), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6167) );
  OR2_X1 U5474 ( .A1(n8687), .A2(n8688), .ZN(n8734) );
  OR2_X1 U5475 ( .A1(n6262), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6273) );
  NAND2_X1 U5476 ( .A1(n6242), .A2(n6241), .ZN(n6252) );
  AND2_X1 U5477 ( .A1(n8826), .A2(n8827), .ZN(n8846) );
  NAND2_X1 U5478 ( .A1(n6210), .A2(n6209), .ZN(n6228) );
  INV_X1 U5479 ( .A(n6211), .ZN(n6210) );
  NAND2_X1 U5480 ( .A1(n6194), .A2(n6193), .ZN(n6203) );
  INV_X1 U5481 ( .A(n6195), .ZN(n6194) );
  NAND2_X1 U5482 ( .A1(n6172), .A2(n6171), .ZN(n6187) );
  INV_X1 U5483 ( .A(n6173), .ZN(n6172) );
  NAND2_X1 U5484 ( .A1(n6143), .A2(n6142), .ZN(n6155) );
  INV_X1 U5485 ( .A(n6144), .ZN(n6143) );
  INV_X1 U5486 ( .A(n6099), .ZN(n6098) );
  NAND2_X1 U5487 ( .A1(n4662), .A2(n4663), .ZN(n7660) );
  AOI21_X1 U5488 ( .B1(n7134), .B2(n4619), .A(n4620), .ZN(n7479) );
  INV_X1 U5489 ( .A(n4621), .ZN(n4619) );
  NAND2_X1 U5490 ( .A1(n4904), .A2(n8417), .ZN(n4621) );
  NAND2_X1 U5491 ( .A1(n5985), .A2(n5984), .ZN(n6009) );
  INV_X1 U5492 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n5984) );
  NAND2_X1 U5493 ( .A1(n8441), .A2(n8456), .ZN(n7104) );
  NAND2_X1 U5494 ( .A1(n6269), .A2(n8548), .ZN(n8785) );
  NAND2_X1 U5495 ( .A1(n4613), .A2(n4611), .ZN(n6269) );
  AOI21_X1 U5496 ( .B1(n4614), .B2(n4330), .A(n4612), .ZN(n4611) );
  NOR2_X1 U5497 ( .A1(n4652), .A2(n4386), .ZN(n4650) );
  AND2_X1 U5498 ( .A1(n4625), .A2(n8530), .ZN(n4624) );
  AOI22_X1 U5499 ( .A1(n8894), .A2(n8904), .B1(n8883), .B2(n8954), .ZN(n8882)
         );
  OAI21_X1 U5500 ( .B1(n7833), .B2(n4635), .A(n4636), .ZN(n6161) );
  NAND2_X1 U5501 ( .A1(n8502), .A2(n8515), .ZN(n4635) );
  AOI21_X1 U5502 ( .B1(n4336), .B2(n8515), .A(n4637), .ZN(n4636) );
  OAI21_X1 U5503 ( .B1(n7654), .B2(n8498), .A(n7650), .ZN(n7833) );
  NOR2_X1 U5504 ( .A1(n6331), .A2(n4352), .ZN(n7651) );
  AND2_X1 U5505 ( .A1(n4662), .A2(n4660), .ZN(n6331) );
  NOR2_X1 U5506 ( .A1(n4661), .A2(n6329), .ZN(n4660) );
  AND2_X1 U5507 ( .A1(n5981), .A2(n4633), .ZN(n10072) );
  INV_X1 U5508 ( .A(n4634), .ZN(n4633) );
  OAI21_X1 U5509 ( .B1(n6022), .B2(n8184), .A(n5980), .ZN(n4634) );
  NAND2_X1 U5510 ( .A1(n4867), .A2(n6391), .ZN(n6461) );
  XNOR2_X1 U5511 ( .A(n5950), .B(n5949), .ZN(n6489) );
  NAND2_X1 U5512 ( .A1(n4355), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5950) );
  NAND2_X1 U5513 ( .A1(n6369), .A2(n6368), .ZN(n6371) );
  INV_X1 U5514 ( .A(n4349), .ZN(n4462) );
  NAND2_X1 U5515 ( .A1(n5429), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n5448) );
  AND2_X1 U5516 ( .A1(n9143), .A2(n5848), .ZN(n9080) );
  AND2_X1 U5517 ( .A1(n5878), .A2(n5877), .ZN(n5896) );
  AND2_X1 U5518 ( .A1(n5077), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5100) );
  NAND2_X1 U5519 ( .A1(n5707), .A2(n9469), .ZN(n5680) );
  XNOR2_X1 U5520 ( .A(n5676), .B(n5874), .ZN(n5684) );
  NAND2_X1 U5521 ( .A1(n5672), .A2(n5703), .ZN(n5673) );
  NAND2_X1 U5522 ( .A1(n9469), .A2(n5780), .ZN(n5674) );
  AND2_X1 U5523 ( .A1(n5860), .A2(n5858), .ZN(n9144) );
  AND2_X1 U5524 ( .A1(n5100), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5121) );
  NAND2_X1 U5525 ( .A1(n4728), .A2(n4727), .ZN(n7486) );
  NAND2_X1 U5526 ( .A1(n4730), .A2(n4729), .ZN(n4727) );
  INV_X1 U5527 ( .A(n5746), .ZN(n4729) );
  INV_X1 U5528 ( .A(n4730), .ZN(n4726) );
  NAND2_X1 U5529 ( .A1(n4750), .A2(n4748), .ZN(n9157) );
  AND2_X1 U5530 ( .A1(n4749), .A2(n9091), .ZN(n4748) );
  INV_X1 U5531 ( .A(n5350), .ZN(n5348) );
  AND2_X1 U5532 ( .A1(n7894), .A2(n7895), .ZN(n5776) );
  INV_X1 U5533 ( .A(n5671), .ZN(n4766) );
  CLKBUF_X1 U5534 ( .A(n7804), .Z(n7805) );
  NAND2_X1 U5535 ( .A1(n5308), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n5324) );
  INV_X1 U5536 ( .A(n5310), .ZN(n5308) );
  OR2_X1 U5537 ( .A1(n5324), .A2(n9182), .ZN(n5350) );
  NOR2_X1 U5538 ( .A1(n5802), .A2(n4374), .ZN(n4759) );
  NAND2_X1 U5539 ( .A1(n9123), .A2(n5803), .ZN(n4760) );
  AND2_X1 U5540 ( .A1(n7645), .A2(n6439), .ZN(n5904) );
  AND2_X1 U5541 ( .A1(n9889), .A2(n9890), .ZN(n9887) );
  OR2_X1 U5542 ( .A1(n6684), .A2(n6683), .ZN(n4477) );
  AOI21_X1 U5543 ( .B1(P1_REG2_REG_3__SCAN_IN), .B2(n8182), .A(n6679), .ZN(
        n9912) );
  NOR2_X1 U5544 ( .A1(n6881), .A2(n4470), .ZN(n6882) );
  NOR2_X1 U5545 ( .A1(n4472), .A2(n4471), .ZN(n4470) );
  INV_X1 U5546 ( .A(n6886), .ZN(n4472) );
  NAND2_X1 U5547 ( .A1(n6882), .A2(n6883), .ZN(n7021) );
  NOR2_X1 U5548 ( .A1(n7341), .A2(n4474), .ZN(n7343) );
  AND2_X1 U5549 ( .A1(n7346), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n4474) );
  NAND2_X1 U5550 ( .A1(n7343), .A2(n7342), .ZN(n7584) );
  NOR2_X1 U5551 ( .A1(n9486), .A2(n4416), .ZN(n9498) );
  NOR2_X1 U5552 ( .A1(n9508), .A2(n9507), .ZN(n9930) );
  OR2_X1 U5553 ( .A1(n9930), .A2(n9929), .ZN(n9926) );
  NOR2_X1 U5554 ( .A1(n8164), .A2(n4490), .ZN(n4489) );
  OR2_X1 U5555 ( .A1(n4492), .A2(n9812), .ZN(n4490) );
  AND2_X1 U5556 ( .A1(n9325), .A2(n9315), .ZN(n9580) );
  NAND2_X1 U5557 ( .A1(n5580), .A2(n9310), .ZN(n9590) );
  NOR2_X1 U5558 ( .A1(n9378), .A2(n4863), .ZN(n4862) );
  INV_X1 U5559 ( .A(n9301), .ZN(n4863) );
  AOI21_X1 U5560 ( .B1(n4678), .B2(n4677), .A(n4384), .ZN(n4676) );
  INV_X1 U5561 ( .A(n4683), .ZN(n4677) );
  NOR2_X1 U5562 ( .A1(n9623), .A2(n9611), .ZN(n9610) );
  NAND2_X1 U5563 ( .A1(n5578), .A2(n9251), .ZN(n9634) );
  NAND2_X1 U5564 ( .A1(n9690), .A2(n4481), .ZN(n9637) );
  AND2_X1 U5565 ( .A1(n4335), .A2(n9638), .ZN(n4481) );
  AND2_X1 U5566 ( .A1(n9253), .A2(n9251), .ZN(n9653) );
  INV_X1 U5567 ( .A(n4858), .ZN(n4857) );
  AOI21_X1 U5568 ( .B1(n4858), .B2(n4861), .A(n4856), .ZN(n4855) );
  NOR2_X1 U5569 ( .A1(n9662), .A2(n4859), .ZN(n4858) );
  NAND2_X1 U5570 ( .A1(n9690), .A2(n4483), .ZN(n4903) );
  NAND2_X1 U5571 ( .A1(n5577), .A2(n9363), .ZN(n9675) );
  OR2_X1 U5572 ( .A1(n5286), .A2(n5285), .ZN(n5310) );
  NAND2_X1 U5573 ( .A1(n4699), .A2(n4702), .ZN(n7777) );
  NAND2_X1 U5574 ( .A1(n7699), .A2(n10040), .ZN(n7772) );
  NAND2_X1 U5575 ( .A1(n5243), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n5266) );
  INV_X1 U5576 ( .A(n5245), .ZN(n5243) );
  OR2_X1 U5577 ( .A1(n5223), .A2(n5222), .ZN(n5245) );
  NAND2_X1 U5578 ( .A1(n7632), .A2(n9396), .ZN(n7631) );
  AND2_X1 U5579 ( .A1(n7633), .A2(n7902), .ZN(n7699) );
  OR2_X1 U5580 ( .A1(n5148), .A2(n5147), .ZN(n5175) );
  NAND2_X1 U5581 ( .A1(n5121), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n5148) );
  OR2_X1 U5582 ( .A1(n7328), .A2(n7334), .ZN(n7435) );
  OR2_X1 U5583 ( .A1(n7495), .A2(n7418), .ZN(n7415) );
  NAND2_X1 U5584 ( .A1(n7321), .A2(n4480), .ZN(n9955) );
  AOI21_X1 U5585 ( .B1(n7174), .B2(n4696), .A(n4381), .ZN(n4695) );
  INV_X1 U5586 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n5058) );
  NOR2_X1 U5587 ( .A1(n5059), .A2(n5058), .ZN(n5077) );
  NOR2_X1 U5588 ( .A1(n7318), .A2(n7317), .ZN(n7321) );
  AND2_X1 U5589 ( .A1(n7321), .A2(n7205), .ZN(n7203) );
  NAND2_X1 U5590 ( .A1(n6974), .A2(n5554), .ZN(n7298) );
  NOR2_X1 U5591 ( .A1(n5672), .A2(n7182), .ZN(n7045) );
  AND2_X1 U5592 ( .A1(n5630), .A2(n9298), .ZN(n9957) );
  AND2_X1 U5593 ( .A1(n5624), .A2(n9841), .ZN(n7032) );
  NAND2_X1 U5594 ( .A1(n5263), .A2(n5262), .ZN(n7773) );
  AND2_X1 U5595 ( .A1(n4919), .A2(n5597), .ZN(n4584) );
  XNOR2_X1 U5596 ( .A(n5502), .B(n5501), .ZN(n7830) );
  XNOR2_X1 U5597 ( .A(n5458), .B(n5457), .ZN(n7761) );
  XNOR2_X1 U5598 ( .A(n5033), .B(SI_4_), .ZN(n5031) );
  NAND2_X1 U5599 ( .A1(n4994), .A2(n4993), .ZN(n5016) );
  XNOR2_X1 U5600 ( .A(n4968), .B(SI_1_), .ZN(n4967) );
  AND2_X1 U5601 ( .A1(n6280), .A2(n6279), .ZN(n8551) );
  NAND2_X1 U5602 ( .A1(n6227), .A2(n6226), .ZN(n8238) );
  NAND2_X1 U5603 ( .A1(n8243), .A2(n8242), .ZN(n8241) );
  NAND2_X1 U5604 ( .A1(n4872), .A2(n8225), .ZN(n8272) );
  NAND2_X1 U5605 ( .A1(n8303), .A2(n8304), .ZN(n4872) );
  NAND2_X1 U5606 ( .A1(n8201), .A2(n4887), .ZN(n8280) );
  OR2_X1 U5607 ( .A1(n6845), .A2(n6846), .ZN(n4895) );
  NAND2_X1 U5608 ( .A1(n7470), .A2(n7469), .ZN(n7714) );
  NAND2_X1 U5609 ( .A1(n8241), .A2(n8211), .ZN(n8312) );
  NAND2_X1 U5610 ( .A1(n4881), .A2(n4880), .ZN(n7904) );
  NAND2_X1 U5611 ( .A1(n4892), .A2(n4891), .ZN(n7151) );
  INV_X1 U5612 ( .A(n4893), .ZN(n4891) );
  INV_X1 U5613 ( .A(n8258), .ZN(n8346) );
  NAND2_X1 U5614 ( .A1(n4792), .A2(n4378), .ZN(n8583) );
  NAND2_X1 U5615 ( .A1(n4796), .A2(n4793), .ZN(n4792) );
  CLKBUF_X1 U5616 ( .A(n6299), .Z(n8609) );
  NAND4_X1 U5617 ( .A1(n5960), .A2(n5959), .A3(n5958), .A4(n5957), .ZN(n8610)
         );
  OR2_X1 U5618 ( .A1(n6285), .A2(n5956), .ZN(n5958) );
  NAND2_X1 U5619 ( .A1(n4587), .A2(n6589), .ZN(n6606) );
  NAND2_X1 U5620 ( .A1(n6817), .A2(n4779), .ZN(n6779) );
  NAND2_X1 U5621 ( .A1(n4602), .A2(n4600), .ZN(n6895) );
  NOR2_X1 U5622 ( .A1(n7061), .A2(n7062), .ZN(n7065) );
  XNOR2_X1 U5623 ( .A(n7498), .B(n7519), .ZN(n7382) );
  INV_X1 U5624 ( .A(n4768), .ZN(n7524) );
  NOR2_X1 U5625 ( .A1(n7729), .A2(n7730), .ZN(n7733) );
  INV_X1 U5626 ( .A(n4594), .ZN(n8659) );
  INV_X1 U5627 ( .A(n4769), .ZN(n8674) );
  OR2_X1 U5628 ( .A1(n8639), .A2(n8640), .ZN(n4594) );
  INV_X1 U5629 ( .A(n8660), .ZN(n4593) );
  NAND2_X1 U5630 ( .A1(n4591), .A2(n4590), .ZN(n8686) );
  NAND2_X1 U5631 ( .A1(n8660), .A2(n4595), .ZN(n4590) );
  OR2_X1 U5632 ( .A1(n8639), .A2(n4592), .ZN(n4591) );
  NAND2_X1 U5633 ( .A1(n4595), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n4592) );
  XNOR2_X1 U5634 ( .A(n8729), .B(n8728), .ZN(n8687) );
  INV_X1 U5635 ( .A(n8734), .ZN(n8727) );
  INV_X1 U5636 ( .A(n4782), .ZN(n8710) );
  AOI21_X1 U5637 ( .B1(n8734), .B2(n8733), .A(n8732), .ZN(n8742) );
  NAND2_X1 U5638 ( .A1(n4786), .A2(n4785), .ZN(n4784) );
  INV_X1 U5639 ( .A(n8762), .ZN(n4785) );
  NAND2_X1 U5640 ( .A1(n8764), .A2(n8763), .ZN(n4786) );
  XNOR2_X1 U5641 ( .A(n4788), .B(n8755), .ZN(n4787) );
  XNOR2_X1 U5642 ( .A(n8573), .B(n8558), .ZN(n8782) );
  OR2_X1 U5643 ( .A1(n8915), .A2(n8790), .ZN(n4668) );
  NAND2_X1 U5644 ( .A1(n4617), .A2(n8540), .ZN(n8809) );
  NAND2_X1 U5645 ( .A1(n6238), .A2(n4351), .ZN(n4617) );
  NAND2_X1 U5646 ( .A1(n7915), .A2(n6338), .ZN(n7956) );
  NAND2_X1 U5647 ( .A1(n6170), .A2(n6169), .ZN(n8959) );
  NAND2_X1 U5648 ( .A1(n6154), .A2(n6153), .ZN(n8289) );
  NAND2_X1 U5649 ( .A1(n7834), .A2(n6336), .ZN(n7863) );
  NAND2_X1 U5650 ( .A1(n6086), .A2(n6085), .ZN(n10131) );
  NAND2_X1 U5651 ( .A1(n6074), .A2(n6073), .ZN(n10124) );
  OAI21_X1 U5652 ( .B1(n7452), .B2(n6326), .A(n6327), .ZN(n7480) );
  NAND2_X1 U5653 ( .A1(n7136), .A2(n8417), .ZN(n7451) );
  NAND2_X1 U5654 ( .A1(n6063), .A2(n6062), .ZN(n7796) );
  NAND2_X1 U5655 ( .A1(n4632), .A2(n8445), .ZN(n7122) );
  INV_X1 U5656 ( .A(n8912), .ZN(n8888) );
  NAND2_X1 U5657 ( .A1(n6284), .A2(n6283), .ZN(n8780) );
  AND2_X1 U5658 ( .A1(n10152), .A2(n10132), .ZN(n8948) );
  INV_X1 U5659 ( .A(n8575), .ZN(n8979) );
  XNOR2_X1 U5660 ( .A(n8785), .B(n8786), .ZN(n8988) );
  NAND2_X1 U5661 ( .A1(n6271), .A2(n6270), .ZN(n8985) );
  AOI21_X1 U5662 ( .B1(n4673), .B2(n8895), .A(n4670), .ZN(n8983) );
  NAND2_X1 U5663 ( .A1(n4672), .A2(n4671), .ZN(n4670) );
  NAND2_X1 U5664 ( .A1(n8788), .A2(n8898), .ZN(n4671) );
  NAND2_X1 U5665 ( .A1(n6261), .A2(n6260), .ZN(n8991) );
  OAI21_X1 U5666 ( .B1(n6238), .B2(n4330), .A(n4614), .ZN(n8793) );
  AND2_X1 U5667 ( .A1(n4651), .A2(n4653), .ZN(n8803) );
  NAND2_X1 U5668 ( .A1(n6238), .A2(n8403), .ZN(n8822) );
  NAND2_X1 U5669 ( .A1(n6240), .A2(n6239), .ZN(n9004) );
  NAND2_X1 U5670 ( .A1(n4657), .A2(n4659), .ZN(n8814) );
  OR2_X1 U5671 ( .A1(n6343), .A2(n6342), .ZN(n4657) );
  INV_X1 U5672 ( .A(n6343), .ZN(n8830) );
  NAND2_X1 U5673 ( .A1(n6208), .A2(n6207), .ZN(n9020) );
  NAND2_X1 U5674 ( .A1(n6202), .A2(n6201), .ZN(n9026) );
  NAND2_X1 U5675 ( .A1(n4623), .A2(n4626), .ZN(n8867) );
  OR2_X1 U5676 ( .A1(n8903), .A2(n4628), .ZN(n4623) );
  NAND2_X1 U5677 ( .A1(n6192), .A2(n6191), .ZN(n9032) );
  NAND2_X1 U5678 ( .A1(n8952), .A2(n8411), .ZN(n8879) );
  OR3_X1 U5679 ( .A1(n8957), .A2(n8956), .A3(n8955), .ZN(n9038) );
  NAND2_X1 U5680 ( .A1(n7867), .A2(n8515), .ZN(n7912) );
  NAND2_X1 U5681 ( .A1(n6125), .A2(n6124), .ZN(n7930) );
  NAND2_X1 U5682 ( .A1(n6113), .A2(n6112), .ZN(n7909) );
  NAND2_X1 U5683 ( .A1(n6096), .A2(n6095), .ZN(n8488) );
  AND2_X1 U5684 ( .A1(n6403), .A2(n6402), .ZN(n10135) );
  INV_X1 U5685 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5930) );
  INV_X1 U5686 ( .A(n5936), .ZN(n8188) );
  INV_X1 U5687 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6454) );
  NAND2_X1 U5688 ( .A1(n4731), .A2(n4732), .ZN(n7241) );
  OR2_X1 U5689 ( .A1(n4350), .A2(n5754), .ZN(n4446) );
  NAND2_X1 U5690 ( .A1(n4747), .A2(n4753), .ZN(n9095) );
  OR2_X1 U5691 ( .A1(n9123), .A2(n4756), .ZN(n4747) );
  NAND2_X1 U5692 ( .A1(n5347), .A2(n5346), .ZN(n9787) );
  NAND2_X1 U5693 ( .A1(n6870), .A2(n5711), .ZN(n6923) );
  NAND2_X1 U5694 ( .A1(n5838), .A2(n9079), .ZN(n9166) );
  NAND2_X1 U5695 ( .A1(n4760), .A2(n4759), .ZN(n9179) );
  INV_X1 U5696 ( .A(n9865), .ZN(n9188) );
  AND2_X1 U5697 ( .A1(n6426), .A2(n6427), .ZN(n6429) );
  NAND2_X1 U5698 ( .A1(n4739), .A2(n4738), .ZN(n9063) );
  AOI21_X1 U5699 ( .B1(n4740), .B2(n4743), .A(n4390), .ZN(n4738) );
  NAND4_X1 U5700 ( .A1(n5030), .A2(n5029), .A3(n5028), .A4(n5027), .ZN(n9465)
         );
  NAND4_X1 U5701 ( .A1(n5012), .A2(n5011), .A3(n5010), .A4(n5009), .ZN(n9466)
         );
  OR2_X1 U5702 ( .A1(n4982), .A2(n4983), .ZN(n4986) );
  NAND2_X1 U5703 ( .A1(n4979), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n4851) );
  OR2_X1 U5704 ( .A1(n4980), .A2(n7190), .ZN(n4853) );
  NAND2_X1 U5705 ( .A1(n9476), .A2(n9475), .ZN(n9474) );
  INV_X1 U5706 ( .A(n4477), .ZN(n6682) );
  NOR2_X1 U5707 ( .A1(n9907), .A2(n4356), .ZN(n6657) );
  NOR2_X1 U5708 ( .A1(n6657), .A2(n6656), .ZN(n6655) );
  NOR2_X1 U5709 ( .A1(n6646), .A2(n6645), .ZN(n6668) );
  AOI21_X1 U5710 ( .B1(P1_REG2_REG_7__SCAN_IN), .B2(n6798), .A(n6793), .ZN(
        n6796) );
  NOR2_X1 U5711 ( .A1(n6797), .A2(n4406), .ZN(n6801) );
  AOI21_X1 U5712 ( .B1(P1_REG2_REG_10__SCAN_IN), .B2(n7266), .A(n7262), .ZN(
        n7264) );
  NOR2_X1 U5713 ( .A1(n7265), .A2(n4475), .ZN(n7269) );
  AND2_X1 U5714 ( .A1(n7266), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n4475) );
  NOR2_X1 U5715 ( .A1(n7269), .A2(n7268), .ZN(n7341) );
  NOR2_X1 U5716 ( .A1(n7681), .A2(n4473), .ZN(n7683) );
  AND2_X1 U5717 ( .A1(n7682), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n4473) );
  NOR2_X1 U5718 ( .A1(n7683), .A2(n7684), .ZN(n9486) );
  XNOR2_X1 U5719 ( .A(n9506), .B(n9505), .ZN(n9485) );
  XNOR2_X1 U5720 ( .A(n9498), .B(n9505), .ZN(n9488) );
  INV_X1 U5721 ( .A(n4764), .ZN(n4762) );
  AND2_X1 U5722 ( .A1(n9521), .A2(n9520), .ZN(n9524) );
  OAI21_X1 U5723 ( .B1(n5500), .B2(n4711), .A(n4708), .ZN(n5662) );
  AOI21_X1 U5724 ( .B1(n4710), .B2(n4709), .A(n4377), .ZN(n4708) );
  NAND2_X1 U5725 ( .A1(n4680), .A2(n4681), .ZN(n9604) );
  NAND2_X1 U5726 ( .A1(n9632), .A2(n4683), .ZN(n4680) );
  NAND2_X1 U5727 ( .A1(n9620), .A2(n9301), .ZN(n9606) );
  OAI21_X1 U5728 ( .B1(n9632), .B2(n4353), .A(n4685), .ZN(n9618) );
  NAND2_X1 U5729 ( .A1(n9678), .A2(n9245), .ZN(n9659) );
  NAND2_X1 U5730 ( .A1(n9780), .A2(n5373), .ZN(n9663) );
  AND2_X1 U5731 ( .A1(n5368), .A2(n5367), .ZN(n9781) );
  OR2_X1 U5732 ( .A1(n9681), .A2(n9680), .ZN(n9780) );
  NAND2_X1 U5733 ( .A1(n4707), .A2(n5329), .ZN(n9689) );
  NAND2_X1 U5734 ( .A1(n5323), .A2(n5322), .ZN(n9793) );
  NAND2_X1 U5735 ( .A1(n9874), .A2(n5295), .ZN(n7939) );
  NAND2_X1 U5736 ( .A1(n4842), .A2(n4843), .ZN(n7881) );
  OR2_X1 U5737 ( .A1(n7885), .A2(n9400), .ZN(n9874) );
  NAND2_X1 U5738 ( .A1(n7695), .A2(n9351), .ZN(n7767) );
  NAND2_X1 U5739 ( .A1(n4722), .A2(n7430), .ZN(n7552) );
  NAND2_X1 U5740 ( .A1(n5172), .A2(n5171), .ZN(n7802) );
  NAND2_X1 U5741 ( .A1(n7420), .A2(n9391), .ZN(n4692) );
  NAND2_X1 U5742 ( .A1(n5119), .A2(n5118), .ZN(n10017) );
  NAND2_X1 U5743 ( .A1(n7199), .A2(n9383), .ZN(n4697) );
  OR2_X1 U5744 ( .A1(n4334), .A2(n9549), .ZN(n9671) );
  OR2_X1 U5745 ( .A1(n5902), .A2(n9292), .ZN(n9727) );
  OR2_X1 U5746 ( .A1(n4334), .A2(n7035), .ZN(n9720) );
  NAND2_X1 U5747 ( .A1(n5220), .A2(n5219), .ZN(n9729) );
  AND2_X1 U5748 ( .A1(n9201), .A2(n9200), .ZN(n9806) );
  NAND2_X1 U5749 ( .A1(n8193), .A2(n8192), .ZN(n9741) );
  NAND2_X1 U5750 ( .A1(n5196), .A2(n5195), .ZN(n7979) );
  AND2_X1 U5751 ( .A1(n4919), .A2(n4928), .ZN(n4465) );
  XNOR2_X1 U5752 ( .A(n5041), .B(P1_IR_REG_5__SCAN_IN), .ZN(n6658) );
  NAND2_X1 U5753 ( .A1(n4430), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4974) );
  NAND3_X1 U5754 ( .A1(n4430), .A2(n4468), .A3(n4467), .ZN(n6637) );
  NAND2_X1 U5755 ( .A1(n4392), .A2(n4998), .ZN(n4467) );
  NAND2_X1 U5756 ( .A1(n4469), .A2(n9844), .ZN(n4468) );
  INV_X1 U5757 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4541) );
  OAI21_X1 U5758 ( .B1(n8983), .B2(n8909), .A(n4666), .ZN(P2_U3205) );
  AOI21_X1 U5759 ( .B1(n4669), .B2(n8906), .A(n4667), .ZN(n4666) );
  NAND2_X1 U5760 ( .A1(n8792), .A2(n4668), .ZN(n4667) );
  INV_X1 U5761 ( .A(n8988), .ZN(n4669) );
  NAND2_X1 U5762 ( .A1(n4450), .A2(n9865), .ZN(n9122) );
  AOI21_X1 U5763 ( .B1(n4429), .B2(n9549), .A(n4428), .ZN(n4427) );
  OR2_X1 U5764 ( .A1(n9551), .A2(n9549), .ZN(n4426) );
  OAI21_X1 U5765 ( .B1(n9553), .B2(n4542), .A(n9552), .ZN(n4428) );
  NAND2_X1 U5766 ( .A1(n9568), .A2(n9777), .ZN(n5631) );
  NAND2_X1 U5767 ( .A1(n9568), .A2(n9832), .ZN(n5636) );
  AND2_X1 U5768 ( .A1(n4483), .A2(n4482), .ZN(n4335) );
  OR2_X1 U5769 ( .A1(n5800), .A2(n9132), .ZN(n5801) );
  INV_X2 U5770 ( .A(n6067), .ZN(n6049) );
  AND2_X1 U5771 ( .A1(n5937), .A2(n8188), .ZN(n5973) );
  AND2_X1 U5772 ( .A1(n9353), .A2(n9357), .ZN(n9400) );
  OR2_X1 U5773 ( .A1(n7866), .A2(n4638), .ZN(n4336) );
  INV_X1 U5774 ( .A(n6285), .ZN(n5972) );
  NAND2_X1 U5775 ( .A1(n4737), .A2(n5839), .ZN(n9082) );
  AND2_X1 U5776 ( .A1(n4607), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n4337) );
  NAND2_X1 U5777 ( .A1(n6219), .A2(n6218), .ZN(n9010) );
  INV_X1 U5778 ( .A(n6823), .ZN(n4607) );
  AND2_X1 U5779 ( .A1(n4576), .A2(n9310), .ZN(n4338) );
  INV_X1 U5780 ( .A(n9662), .ZN(n4718) );
  INV_X1 U5781 ( .A(n9227), .ZN(n4844) );
  AND3_X1 U5782 ( .A1(n9325), .A2(n9324), .A3(n4552), .ZN(n4339) );
  AND2_X1 U5783 ( .A1(n4760), .A2(n5801), .ZN(n9134) );
  AND2_X1 U5784 ( .A1(n8574), .A2(n8552), .ZN(n4340) );
  INV_X1 U5785 ( .A(n7866), .ZN(n4648) );
  AND2_X1 U5786 ( .A1(n4864), .A2(n9300), .ZN(n4341) );
  AND2_X1 U5787 ( .A1(n4403), .A2(n4602), .ZN(n4342) );
  AND2_X1 U5788 ( .A1(n8533), .A2(n8530), .ZN(n4343) );
  AND2_X1 U5789 ( .A1(n7903), .A2(n4882), .ZN(n4344) );
  NAND2_X1 U5790 ( .A1(n6251), .A2(n6250), .ZN(n8998) );
  INV_X1 U5791 ( .A(n8998), .ZN(n4658) );
  NAND2_X1 U5792 ( .A1(n6908), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n4606) );
  AND2_X1 U5793 ( .A1(n4486), .A2(n4485), .ZN(n4345) );
  NOR2_X1 U5794 ( .A1(n9242), .A2(n4552), .ZN(n4346) );
  INV_X1 U5795 ( .A(n4744), .ZN(n4464) );
  AOI21_X1 U5796 ( .B1(n5776), .B2(n4745), .A(n4387), .ZN(n4744) );
  NAND2_X1 U5797 ( .A1(n5411), .A2(n5410), .ZN(n9647) );
  INV_X1 U5798 ( .A(n9647), .ZN(n4482) );
  AND2_X1 U5799 ( .A1(n4457), .A2(n4462), .ZN(n4347) );
  AND2_X1 U5800 ( .A1(n4790), .A2(n5480), .ZN(n4348) );
  INV_X1 U5801 ( .A(n4984), .ZN(n5516) );
  INV_X2 U5802 ( .A(n5052), .ZN(n5114) );
  INV_X1 U5803 ( .A(n5703), .ZN(n5820) );
  INV_X1 U5804 ( .A(n6728), .ZN(n8227) );
  INV_X1 U5805 ( .A(n8227), .ZN(n8254) );
  XOR2_X1 U5806 ( .A(n5781), .B(n5886), .Z(n4349) );
  OAI21_X1 U5807 ( .B1(n5859), .B2(n4743), .A(n4740), .ZN(n6426) );
  XNOR2_X1 U5808 ( .A(n5886), .B(n5755), .ZN(n4350) );
  INV_X1 U5809 ( .A(n6611), .ZN(n6586) );
  NAND2_X1 U5810 ( .A1(n4735), .A2(n4453), .ZN(n9083) );
  NAND2_X1 U5811 ( .A1(n4674), .A2(n5928), .ZN(n6296) );
  NAND2_X1 U5812 ( .A1(n9190), .A2(n5788), .ZN(n9123) );
  NAND2_X1 U5813 ( .A1(n5133), .A2(n5095), .ZN(n5129) );
  AND2_X1 U5814 ( .A1(n8403), .A2(n4618), .ZN(n4351) );
  NOR2_X1 U5815 ( .A1(n8492), .A2(n7662), .ZN(n4352) );
  AND2_X1 U5816 ( .A1(n9824), .A2(n9448), .ZN(n4353) );
  OR2_X1 U5817 ( .A1(n6443), .A2(n5954), .ZN(n4354) );
  AND3_X1 U5818 ( .A1(n4834), .A2(n4913), .A3(n4973), .ZN(n5053) );
  NAND2_X1 U5819 ( .A1(n6290), .A2(n4675), .ZN(n4355) );
  AND2_X1 U5820 ( .A1(n9910), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n4356) );
  OR2_X1 U5821 ( .A1(n4982), .A2(n4852), .ZN(n4357) );
  OR2_X1 U5822 ( .A1(n8673), .A2(n8672), .ZN(n4358) );
  NAND2_X1 U5823 ( .A1(n4871), .A2(n4870), .ZN(n8340) );
  INV_X1 U5824 ( .A(n4606), .ZN(n4605) );
  AND2_X1 U5825 ( .A1(n9891), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n4359) );
  AND4_X1 U5826 ( .A1(n8402), .A2(n8786), .A3(n8401), .A4(n8821), .ZN(n4360)
         );
  AND2_X1 U5827 ( .A1(n4734), .A2(n4899), .ZN(n4361) );
  NAND2_X1 U5828 ( .A1(n8370), .A2(n8369), .ZN(n8571) );
  AND2_X1 U5829 ( .A1(n4349), .A2(n9070), .ZN(n4362) );
  NAND2_X1 U5830 ( .A1(n6259), .A2(n6258), .ZN(n8815) );
  INV_X1 U5831 ( .A(n8815), .ZN(n6346) );
  OR2_X1 U5832 ( .A1(n7162), .A2(n7167), .ZN(n4363) );
  OR3_X1 U5833 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(n4998), .A3(
        P1_IR_REG_0__SCAN_IN), .ZN(n4364) );
  INV_X1 U5834 ( .A(n6775), .ZN(n4781) );
  INV_X1 U5835 ( .A(n7724), .ZN(n4878) );
  INV_X1 U5836 ( .A(n8816), .ZN(n8844) );
  AND2_X1 U5837 ( .A1(n9351), .A2(n9226), .ZN(n9399) );
  INV_X1 U5838 ( .A(n9399), .ZN(n4845) );
  INV_X1 U5839 ( .A(n5086), .ZN(n5087) );
  XNOR2_X1 U5840 ( .A(n5089), .B(SI_7_), .ZN(n5086) );
  NOR2_X1 U5841 ( .A1(n8493), .A2(n8492), .ZN(n4365) );
  OR2_X1 U5842 ( .A1(n9595), .A2(n4492), .ZN(n4366) );
  OR2_X1 U5843 ( .A1(n8954), .A2(n8334), .ZN(n8411) );
  INV_X1 U5844 ( .A(n8411), .ZN(n4630) );
  INV_X1 U5845 ( .A(n8540), .ZN(n4616) );
  INV_X1 U5846 ( .A(n6299), .ZN(n4438) );
  NOR2_X1 U5847 ( .A1(n8509), .A2(n8552), .ZN(n4367) );
  OR2_X1 U5848 ( .A1(n8728), .A2(n8709), .ZN(n4368) );
  INV_X1 U5849 ( .A(n7890), .ZN(n5589) );
  NAND2_X1 U5850 ( .A1(n5284), .A2(n5283), .ZN(n7890) );
  AND2_X1 U5851 ( .A1(n7600), .A2(n7599), .ZN(n4369) );
  INV_X1 U5852 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5546) );
  AND2_X1 U5853 ( .A1(n8794), .A2(n8546), .ZN(n4370) );
  INV_X1 U5854 ( .A(n4861), .ZN(n4860) );
  NAND2_X1 U5855 ( .A1(n9680), .A2(n9363), .ZN(n4861) );
  NAND2_X1 U5856 ( .A1(n5647), .A2(n5646), .ZN(n8164) );
  NAND2_X1 U5857 ( .A1(n9611), .A2(n9446), .ZN(n4371) );
  INV_X1 U5858 ( .A(n4491), .ZN(n9582) );
  NOR2_X1 U5859 ( .A1(n9595), .A2(n9583), .ZN(n4491) );
  AND2_X1 U5860 ( .A1(n5715), .A2(n5711), .ZN(n4372) );
  AND2_X1 U5861 ( .A1(n8959), .A2(n8897), .ZN(n4373) );
  NOR2_X1 U5862 ( .A1(n5806), .A2(n5805), .ZN(n4374) );
  AND2_X1 U5863 ( .A1(n4594), .A2(n4593), .ZN(n4375) );
  AND2_X1 U5864 ( .A1(n5579), .A2(n9300), .ZN(n4376) );
  AND2_X1 U5865 ( .A1(n9568), .A2(n9443), .ZN(n4377) );
  OR2_X1 U5866 ( .A1(n8979), .A2(n8582), .ZN(n4378) );
  AND2_X1 U5867 ( .A1(n8533), .A2(n8532), .ZN(n4379) );
  NOR2_X1 U5868 ( .A1(n10124), .A2(n8599), .ZN(n4380) );
  NOR2_X1 U5869 ( .A1(n7179), .A2(n9464), .ZN(n4381) );
  NOR2_X1 U5870 ( .A1(n7338), .A2(n9460), .ZN(n4382) );
  NOR2_X1 U5871 ( .A1(n7946), .A2(n9453), .ZN(n4383) );
  NOR2_X1 U5872 ( .A1(n9611), .A2(n9446), .ZN(n4384) );
  OR2_X1 U5873 ( .A1(n9076), .A2(n9456), .ZN(n4385) );
  INV_X1 U5874 ( .A(n4823), .ZN(n4509) );
  NOR2_X1 U5875 ( .A1(n5129), .A2(n4824), .ZN(n4823) );
  AND2_X1 U5876 ( .A1(n6346), .A2(n4658), .ZN(n4386) );
  NOR2_X1 U5877 ( .A1(n5779), .A2(n5778), .ZN(n4387) );
  OR2_X1 U5878 ( .A1(n6818), .A2(n4776), .ZN(n4388) );
  AND2_X1 U5879 ( .A1(n9787), .A2(n9451), .ZN(n4389) );
  INV_X1 U5880 ( .A(n4711), .ZN(n4710) );
  NAND2_X1 U5881 ( .A1(n4715), .A2(n4716), .ZN(n4711) );
  NAND2_X1 U5882 ( .A1(n6428), .A2(n6427), .ZN(n4390) );
  INV_X1 U5883 ( .A(n4679), .ZN(n4678) );
  NAND2_X1 U5884 ( .A1(n4681), .A2(n4371), .ZN(n4679) );
  OAI21_X1 U5885 ( .B1(n4621), .B2(n6056), .A(n8473), .ZN(n4620) );
  NAND2_X1 U5886 ( .A1(n9229), .A2(n9351), .ZN(n4391) );
  INV_X1 U5887 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n4765) );
  AND2_X1 U5888 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n4392) );
  INV_X1 U5889 ( .A(n9680), .ZN(n5372) );
  AND2_X1 U5890 ( .A1(n9246), .A2(n9245), .ZN(n9680) );
  INV_X1 U5891 ( .A(n9254), .ZN(n4582) );
  NOR2_X2 U5892 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n4973) );
  INV_X1 U5893 ( .A(n4973), .ZN(n4430) );
  NAND2_X1 U5894 ( .A1(n4581), .A2(n4578), .ZN(n4393) );
  NAND2_X1 U5895 ( .A1(n5488), .A2(n5487), .ZN(n9812) );
  OAI21_X1 U5896 ( .B1(n9632), .B2(n4679), .A(n4676), .ZN(n9593) );
  AND2_X1 U5897 ( .A1(n4626), .A2(n8532), .ZN(n4394) );
  AND3_X1 U5898 ( .A1(n4518), .A2(n8417), .A3(n4904), .ZN(n4395) );
  AND2_X1 U5899 ( .A1(n8513), .A2(n8502), .ZN(n8501) );
  AND2_X1 U5900 ( .A1(n5205), .A2(n7430), .ZN(n4396) );
  AND2_X1 U5901 ( .A1(n4849), .A2(n9218), .ZN(n4397) );
  INV_X1 U5902 ( .A(n4884), .ZN(n4883) );
  NAND2_X1 U5903 ( .A1(n8813), .A2(n8805), .ZN(n4398) );
  AND2_X1 U5904 ( .A1(n4898), .A2(n5929), .ZN(n4399) );
  NOR2_X1 U5905 ( .A1(n4464), .A2(n4459), .ZN(n4458) );
  AND2_X1 U5906 ( .A1(n8212), .A2(n8211), .ZN(n4400) );
  AND2_X1 U5907 ( .A1(n5928), .A2(n6394), .ZN(n4401) );
  NAND2_X1 U5908 ( .A1(n5428), .A2(n5427), .ZN(n9824) );
  NAND2_X1 U5909 ( .A1(n9240), .A2(n9362), .ZN(n4402) );
  AND2_X1 U5910 ( .A1(n4600), .A2(n4606), .ZN(n4403) );
  OR2_X1 U5911 ( .A1(n9583), .A2(n6431), .ZN(n9325) );
  AND2_X1 U5912 ( .A1(n7821), .A2(n4884), .ZN(n4880) );
  INV_X1 U5913 ( .A(n4653), .ZN(n4652) );
  AND2_X1 U5914 ( .A1(n4654), .A2(n4398), .ZN(n4653) );
  INV_X1 U5915 ( .A(n5776), .ZN(n4746) );
  OR2_X1 U5916 ( .A1(n8181), .A2(n8188), .ZN(n6285) );
  INV_X1 U5917 ( .A(n7773), .ZN(n4701) );
  INV_X1 U5918 ( .A(n6909), .ZN(n4604) );
  XNOR2_X1 U5919 ( .A(n5548), .B(P1_IR_REG_21__SCAN_IN), .ZN(n5670) );
  NAND2_X1 U5920 ( .A1(n5515), .A2(n5514), .ZN(n9583) );
  INV_X1 U5921 ( .A(n9583), .ZN(n4493) );
  INV_X1 U5922 ( .A(n5973), .ZN(n6067) );
  NAND2_X1 U5923 ( .A1(n5552), .A2(n9333), .ZN(n7038) );
  INV_X1 U5924 ( .A(n7334), .ZN(n4688) );
  NOR2_X1 U5925 ( .A1(n7833), .A2(n6132), .ZN(n4640) );
  NAND2_X1 U5926 ( .A1(n7804), .A2(n5768), .ZN(n7893) );
  AND2_X1 U5927 ( .A1(n9690), .A2(n4335), .ZN(n4404) );
  AND2_X1 U5928 ( .A1(n7699), .A2(n4488), .ZN(n4405) );
  AND2_X1 U5929 ( .A1(n6798), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n4406) );
  NAND2_X1 U5930 ( .A1(n4761), .A2(n4919), .ZN(n5281) );
  INV_X1 U5931 ( .A(n9619), .ZN(n4864) );
  NAND2_X1 U5932 ( .A1(n7631), .A2(n5231), .ZN(n7697) );
  INV_X1 U5933 ( .A(n5860), .ZN(n4743) );
  INV_X1 U5934 ( .A(n4830), .ZN(n4829) );
  NOR2_X1 U5935 ( .A1(n5278), .A2(SI_15_), .ZN(n4830) );
  XNOR2_X1 U5936 ( .A(n5605), .B(P1_IR_REG_24__SCAN_IN), .ZN(n5608) );
  AND2_X1 U5937 ( .A1(n6658), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n4407) );
  INV_X1 U5938 ( .A(n9351), .ZN(n4848) );
  INV_X1 U5939 ( .A(n9167), .ZN(n5839) );
  INV_X1 U5940 ( .A(n4761), .ZN(n5238) );
  AND2_X1 U5941 ( .A1(n8226), .A2(n8805), .ZN(n4408) );
  AND2_X1 U5942 ( .A1(n4639), .A2(n8513), .ZN(n4409) );
  AND2_X1 U5943 ( .A1(n7893), .A2(n5776), .ZN(n4410) );
  NAND2_X1 U5944 ( .A1(n4761), .A2(n4762), .ZN(n4411) );
  INV_X1 U5945 ( .A(n4457), .ZN(n4463) );
  AND2_X1 U5946 ( .A1(n5402), .A2(SI_21_), .ZN(n4412) );
  OR2_X1 U5947 ( .A1(n5334), .A2(n4819), .ZN(n4413) );
  AND2_X1 U5948 ( .A1(n4463), .A2(n4349), .ZN(n4414) );
  INV_X1 U5949 ( .A(n7946), .ZN(n4485) );
  AND2_X1 U5950 ( .A1(n6379), .A2(n6475), .ZN(n6724) );
  INV_X1 U5951 ( .A(n5707), .ZN(n5782) );
  NAND2_X1 U5952 ( .A1(n5734), .A2(n4899), .ZN(n7228) );
  INV_X1 U5953 ( .A(n5478), .ZN(n5479) );
  NAND2_X1 U5954 ( .A1(n4697), .A2(n5045), .ZN(n7173) );
  NAND2_X1 U5955 ( .A1(n4692), .A2(n5128), .ZN(n7333) );
  INV_X1 U5956 ( .A(n9781), .ZN(n4484) );
  AND2_X1 U5957 ( .A1(n9487), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n4415) );
  AND2_X1 U5958 ( .A1(n9487), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n4416) );
  AND2_X1 U5959 ( .A1(n7751), .A2(n7599), .ZN(n4417) );
  AND2_X1 U5960 ( .A1(n5644), .A2(n5643), .ZN(n4418) );
  NAND2_X1 U5961 ( .A1(n4609), .A2(n7616), .ZN(n4419) );
  AND2_X1 U5962 ( .A1(n8652), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n4420) );
  AND2_X1 U5963 ( .A1(n4895), .A2(n4894), .ZN(n4421) );
  NAND2_X1 U5964 ( .A1(n4770), .A2(n6777), .ZN(n6817) );
  INV_X1 U5965 ( .A(n9278), .ZN(n4552) );
  NAND2_X1 U5966 ( .A1(n5075), .A2(n5074), .ZN(n9954) );
  INV_X1 U5967 ( .A(n9954), .ZN(n4479) );
  NAND2_X1 U5968 ( .A1(n6870), .A2(n4372), .ZN(n6924) );
  INV_X1 U5969 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n4641) );
  NAND4_X1 U5970 ( .A1(n4920), .A2(n4926), .A3(n4465), .A4(n4466), .ZN(n9843)
         );
  INV_X1 U5971 ( .A(n4936), .ZN(n9848) );
  INV_X1 U5972 ( .A(n4934), .ZN(n9851) );
  INV_X1 U5973 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n5985) );
  INV_X1 U5974 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n4852) );
  INV_X1 U5975 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n4471) );
  INV_X2 U5976 ( .A(n9056), .ZN(n8186) );
  NAND3_X1 U5977 ( .A1(n4547), .A2(n9363), .A3(n9246), .ZN(n4546) );
  NAND2_X1 U5978 ( .A1(n4558), .A2(n4556), .ZN(n4555) );
  MUX2_X2 U5979 ( .A(n9281), .B(n9278), .S(n9741), .Z(n9280) );
  OAI21_X2 U5980 ( .B1(n9280), .B2(n9417), .A(n9279), .ZN(n9285) );
  OAI21_X1 U5981 ( .B1(n7311), .B2(n4583), .A(n4836), .ZN(n7175) );
  NAND2_X1 U5982 ( .A1(n4543), .A2(n5551), .ZN(n7040) );
  OAI21_X1 U5983 ( .B1(n9217), .B2(n9216), .A(n9215), .ZN(n9219) );
  NAND2_X1 U5984 ( .A1(n9203), .A2(n9214), .ZN(n4553) );
  AOI21_X1 U5985 ( .B1(n9278), .B2(n9244), .A(n9243), .ZN(n9250) );
  NAND2_X1 U5986 ( .A1(n7883), .A2(n9353), .ZN(n7941) );
  NAND2_X1 U5987 ( .A1(n4850), .A2(n4397), .ZN(n7547) );
  NAND3_X1 U5988 ( .A1(n5666), .A2(n4907), .A3(n5665), .ZN(P1_U3519) );
  NAND2_X1 U5989 ( .A1(n5557), .A2(n5556), .ZN(n7311) );
  NAND2_X1 U5990 ( .A1(n4554), .A2(n9276), .ZN(n9281) );
  NAND2_X1 U5991 ( .A1(n7175), .A2(n5561), .ZN(n7360) );
  INV_X1 U5992 ( .A(n7038), .ZN(n4543) );
  NAND2_X1 U5993 ( .A1(n4724), .A2(n4723), .ZN(n4944) );
  NOR2_X1 U5994 ( .A1(n7417), .A2(n7416), .ZN(n9203) );
  NAND2_X1 U5995 ( .A1(n9264), .A2(n9317), .ZN(n4564) );
  NOR2_X2 U5996 ( .A1(n8712), .A2(n8711), .ZN(n8754) );
  NAND4_X2 U5997 ( .A1(n6513), .A2(n5914), .A3(n4896), .A4(n5915), .ZN(n5991)
         );
  NAND2_X2 U5998 ( .A1(n6006), .A2(n6005), .ZN(n6908) );
  NOR2_X1 U5999 ( .A1(n8628), .A2(n6911), .ZN(n6912) );
  XNOR2_X1 U6000 ( .A(n8672), .B(n8673), .ZN(n8653) );
  AOI21_X1 U6001 ( .B1(n8501), .B2(n6336), .A(n4648), .ZN(n4647) );
  XNOR2_X2 U6002 ( .A(n8608), .B(n8420), .ZN(n6704) );
  AOI21_X1 U6003 ( .B1(n6366), .B2(n8895), .A(n4423), .ZN(n8776) );
  NAND2_X2 U6004 ( .A1(n6325), .A2(n6324), .ZN(n7452) );
  OAI22_X1 U6005 ( .A1(n7105), .A2(n6304), .B1(n10072), .B2(n6844), .ZN(n7090)
         );
  AOI21_X1 U6006 ( .B1(n6348), .B2(n8806), .A(n6347), .ZN(n8787) );
  NAND2_X1 U6007 ( .A1(n4427), .A2(n4426), .ZN(P1_U3262) );
  NAND2_X1 U6008 ( .A1(n7347), .A2(n7348), .ZN(n7580) );
  NAND2_X1 U6009 ( .A1(n6887), .A2(n6888), .ZN(n7017) );
  INV_X1 U6010 ( .A(n9550), .ZN(n4429) );
  NAND2_X1 U6011 ( .A1(n9524), .A2(n9523), .ZN(n9539) );
  AOI21_X1 U6012 ( .B1(n9910), .B2(P1_REG2_REG_4__SCAN_IN), .A(n9911), .ZN(
        n6653) );
  AOI21_X1 U6013 ( .B1(P1_REG2_REG_6__SCAN_IN), .B2(n6669), .A(n6664), .ZN(
        n6667) );
  AOI21_X1 U6014 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(n7682), .A(n7675), .ZN(
        n7678) );
  AOI21_X2 U6015 ( .B1(n7929), .B2(n7928), .A(n4431), .ZN(n7932) );
  AOI21_X2 U6016 ( .B1(n8264), .B2(n8265), .A(n4432), .ZN(n8324) );
  AOI22_X2 U6017 ( .A1(n6758), .A2(n6759), .B1(n6754), .B2(n6729), .ZN(n6736)
         );
  NAND2_X2 U6018 ( .A1(n4435), .A2(n6726), .ZN(n6728) );
  OAI21_X1 U6019 ( .B1(n6725), .B2(n8426), .A(n8568), .ZN(n4435) );
  NAND2_X1 U6020 ( .A1(n7465), .A2(n7464), .ZN(n7573) );
  INV_X1 U6021 ( .A(n6845), .ZN(n4889) );
  NOR2_X2 U6022 ( .A1(n5991), .A2(n5919), .ZN(n6060) );
  NOR2_X1 U6023 ( .A1(n8651), .A2(n4420), .ZN(n8672) );
  NOR2_X1 U6024 ( .A1(n8700), .A2(n4783), .ZN(n8709) );
  NOR2_X1 U6025 ( .A1(n8754), .A2(n8753), .ZN(n4788) );
  INV_X1 U6026 ( .A(n6859), .ZN(n4439) );
  NAND2_X1 U6027 ( .A1(n6290), .A2(n4401), .ZN(n4610) );
  NAND2_X1 U6028 ( .A1(n4643), .A2(n4642), .ZN(n8894) );
  OAI211_X2 U6029 ( .C1(n8368), .C2(P1_DATAO_REG_1__SCAN_IN), .A(n5955), .B(
        n4354), .ZN(n6859) );
  NOR2_X1 U6030 ( .A1(n6681), .A2(n6680), .ZN(n6679) );
  NAND2_X1 U6031 ( .A1(n6871), .A2(n6872), .ZN(n6870) );
  NAND3_X1 U6032 ( .A1(n4731), .A2(n5746), .A3(n4726), .ZN(n7487) );
  NAND2_X1 U6033 ( .A1(n6691), .A2(n5693), .ZN(n4441) );
  INV_X1 U6034 ( .A(n6691), .ZN(n4444) );
  NAND2_X1 U6035 ( .A1(n4442), .A2(n4441), .ZN(n6833) );
  AND2_X1 U6036 ( .A1(n6835), .A2(n4443), .ZN(n4442) );
  NAND2_X1 U6037 ( .A1(n6694), .A2(n5693), .ZN(n4443) );
  NAND2_X1 U6038 ( .A1(n6692), .A2(n5693), .ZN(n6834) );
  NAND2_X1 U6039 ( .A1(n4444), .A2(n5692), .ZN(n6692) );
  NAND4_X2 U6040 ( .A1(n4940), .A2(n4939), .A3(n4937), .A4(n4938), .ZN(n9469)
         );
  NAND2_X1 U6041 ( .A1(n9970), .A2(n9469), .ZN(n9333) );
  OAI21_X1 U6042 ( .B1(n7536), .B2(n4448), .A(n4447), .ZN(n5756) );
  NAND2_X1 U6043 ( .A1(n4454), .A2(n9079), .ZN(n4453) );
  INV_X1 U6044 ( .A(n5838), .ZN(n4454) );
  NAND2_X1 U6045 ( .A1(n7804), .A2(n4458), .ZN(n4455) );
  OAI21_X1 U6046 ( .B1(n7804), .B2(n4746), .A(n4744), .ZN(n4457) );
  NAND2_X1 U6047 ( .A1(n4455), .A2(n4456), .ZN(n5787) );
  AND3_X1 U6048 ( .A1(n4920), .A2(n4926), .A3(n4919), .ZN(n4724) );
  AND4_X1 U6049 ( .A1(n4920), .A2(n4926), .A3(n4466), .A4(n4919), .ZN(n4931)
         );
  MUX2_X1 U6050 ( .A(n10050), .B(P1_REG1_REG_1__SCAN_IN), .S(n6637), .Z(n9476)
         );
  AND2_X2 U6051 ( .A1(n4918), .A2(n5053), .ZN(n4920) );
  NAND2_X1 U6052 ( .A1(n7370), .A2(n10013), .ZN(n7422) );
  NAND2_X1 U6053 ( .A1(n7699), .A2(n4345), .ZN(n9711) );
  NAND2_X1 U6054 ( .A1(n9610), .A2(n4489), .ZN(n8194) );
  NAND2_X1 U6055 ( .A1(n9610), .A2(n9596), .ZN(n9595) );
  OR2_X1 U6056 ( .A1(n4500), .A2(n5088), .ZN(n4506) );
  NAND3_X1 U6057 ( .A1(n4506), .A2(n4504), .A3(n4501), .ZN(n6484) );
  NAND3_X1 U6058 ( .A1(n5088), .A2(n4507), .A3(n4505), .ZN(n4504) );
  NAND2_X1 U6059 ( .A1(n4514), .A2(n4515), .ZN(n8514) );
  NAND2_X1 U6060 ( .A1(n8494), .A2(n4516), .ZN(n4514) );
  NAND3_X1 U6061 ( .A1(n8417), .A2(n8416), .A3(n8567), .ZN(n4522) );
  OAI21_X1 U6062 ( .B1(n8534), .B2(n4529), .A(n4524), .ZN(n8538) );
  NAND2_X1 U6063 ( .A1(n4534), .A2(n8568), .ZN(n4796) );
  NAND2_X1 U6064 ( .A1(n4537), .A2(n4535), .ZN(n4534) );
  NAND2_X1 U6065 ( .A1(n4536), .A2(n8567), .ZN(n4535) );
  NAND2_X1 U6066 ( .A1(n8566), .A2(n8565), .ZN(n4536) );
  AOI21_X1 U6067 ( .B1(n8566), .B2(n4340), .A(n8569), .ZN(n4537) );
  INV_X2 U6068 ( .A(n4332), .ZN(n8358) );
  NAND2_X1 U6069 ( .A1(n5319), .A2(n5340), .ZN(n5538) );
  NAND2_X1 U6070 ( .A1(n4545), .A2(n4544), .ZN(n9243) );
  OAI21_X1 U6071 ( .B1(n4549), .B2(n4402), .A(n4346), .ZN(n4544) );
  NAND2_X1 U6072 ( .A1(n4546), .A2(n4552), .ZN(n4545) );
  OAI21_X1 U6073 ( .B1(n4549), .B2(n9360), .A(n4548), .ZN(n4547) );
  INV_X1 U6074 ( .A(n9364), .ZN(n4548) );
  OAI21_X1 U6075 ( .B1(n9217), .B2(n9209), .A(n9342), .ZN(n9210) );
  AND2_X1 U6076 ( .A1(n4551), .A2(n4550), .ZN(n9217) );
  AOI21_X1 U6077 ( .B1(n9207), .B2(n9278), .A(n9209), .ZN(n4550) );
  NAND3_X1 U6078 ( .A1(n4563), .A2(n4559), .A3(n4555), .ZN(n4554) );
  NAND2_X1 U6079 ( .A1(n4565), .A2(n4566), .ZN(n9213) );
  NAND2_X1 U6080 ( .A1(n9211), .A2(n4567), .ZN(n4565) );
  NAND2_X1 U6081 ( .A1(n4573), .A2(n4574), .ZN(n9267) );
  NAND2_X1 U6082 ( .A1(n9255), .A2(n4338), .ZN(n4573) );
  OAI21_X1 U6083 ( .B1(n9255), .B2(n4577), .A(n4576), .ZN(n9266) );
  NAND3_X1 U6084 ( .A1(n4920), .A2(n4584), .A3(n4926), .ZN(n4941) );
  INV_X1 U6085 ( .A(n4724), .ZN(n5596) );
  NAND2_X1 U6086 ( .A1(n4586), .A2(n6589), .ZN(n4589) );
  XNOR2_X1 U6087 ( .A(n8658), .B(n8673), .ZN(n8639) );
  INV_X1 U6088 ( .A(n6770), .ZN(n4603) );
  INV_X1 U6089 ( .A(n6822), .ZN(n4601) );
  OAI21_X1 U6090 ( .B1(n6770), .B2(n4599), .A(n4598), .ZN(n8621) );
  NAND2_X2 U6091 ( .A1(n6369), .A2(n5943), .ZN(n6374) );
  NAND2_X2 U6092 ( .A1(n4610), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6369) );
  OR2_X1 U6093 ( .A1(n8368), .A2(n6446), .ZN(n5971) );
  NAND2_X1 U6094 ( .A1(n6238), .A2(n4614), .ZN(n4613) );
  NAND2_X1 U6095 ( .A1(n8903), .A2(n4394), .ZN(n4622) );
  NAND2_X1 U6096 ( .A1(n4622), .A2(n4624), .ZN(n8862) );
  NAND3_X1 U6097 ( .A1(n4626), .A2(n8532), .A3(n4628), .ZN(n4625) );
  NAND2_X1 U6098 ( .A1(n4632), .A2(n4631), .ZN(n7124) );
  INV_X1 U6099 ( .A(n10072), .ZN(n7108) );
  INV_X1 U6100 ( .A(n4640), .ZN(n4639) );
  NAND2_X1 U6101 ( .A1(n7913), .A2(n4644), .ZN(n4643) );
  NAND2_X1 U6102 ( .A1(n7836), .A2(n6336), .ZN(n4649) );
  NAND2_X1 U6103 ( .A1(n4651), .A2(n4650), .ZN(n6345) );
  NAND2_X1 U6104 ( .A1(n6343), .A2(n4655), .ZN(n4651) );
  NAND2_X1 U6105 ( .A1(n7452), .A2(n4664), .ZN(n4662) );
  XNOR2_X1 U6106 ( .A(n8787), .B(n8786), .ZN(n4673) );
  NAND4_X1 U6107 ( .A1(n6060), .A2(n5925), .A3(n4675), .A4(n5949), .ZN(n5934)
         );
  CLKBUF_X1 U6108 ( .A(n6290), .Z(n4674) );
  NAND2_X1 U6109 ( .A1(n7420), .A2(n4687), .ZN(n4686) );
  NAND2_X1 U6110 ( .A1(n4686), .A2(n4690), .ZN(n7429) );
  NAND2_X1 U6111 ( .A1(n7199), .A2(n4694), .ZN(n4693) );
  NAND2_X1 U6112 ( .A1(n4693), .A2(n4695), .ZN(n9943) );
  OR2_X1 U6113 ( .A1(n7632), .A2(n4704), .ZN(n4699) );
  NAND2_X1 U6114 ( .A1(n4698), .A2(n4700), .ZN(n5273) );
  NAND2_X1 U6115 ( .A1(n7632), .A2(n4702), .ZN(n4698) );
  NAND2_X1 U6116 ( .A1(n4707), .A2(n4705), .ZN(n5359) );
  NAND2_X1 U6117 ( .A1(n5500), .A2(n4713), .ZN(n4712) );
  NAND2_X1 U6118 ( .A1(n5500), .A2(n5499), .ZN(n9581) );
  NAND2_X1 U6119 ( .A1(n9681), .A2(n5373), .ZN(n4719) );
  NAND2_X1 U6120 ( .A1(n4720), .A2(n4721), .ZN(n5315) );
  NAND2_X1 U6121 ( .A1(n7885), .A2(n5295), .ZN(n4720) );
  NAND2_X1 U6122 ( .A1(n5183), .A2(n5182), .ZN(n4722) );
  NAND2_X1 U6123 ( .A1(n4722), .A2(n4396), .ZN(n5207) );
  NAND2_X1 U6124 ( .A1(n5785), .A2(n5784), .ZN(n5788) );
  NAND2_X1 U6125 ( .A1(n5787), .A2(n5786), .ZN(n4725) );
  NAND3_X1 U6126 ( .A1(n4361), .A2(n5734), .A3(n4729), .ZN(n4728) );
  INV_X1 U6127 ( .A(n9166), .ZN(n4737) );
  NAND2_X1 U6128 ( .A1(n5859), .A2(n4740), .ZN(n4739) );
  NAND2_X1 U6129 ( .A1(n5859), .A2(n9144), .ZN(n9147) );
  NAND2_X1 U6130 ( .A1(n9123), .A2(n4751), .ZN(n4750) );
  NAND3_X1 U6131 ( .A1(n4753), .A2(n4756), .A3(n4752), .ZN(n4749) );
  NAND2_X1 U6132 ( .A1(n4920), .A2(n4763), .ZN(n5537) );
  INV_X1 U6133 ( .A(n5537), .ZN(n5540) );
  CLKBUF_X1 U6134 ( .A(n4920), .Z(n4761) );
  NOR2_X1 U6135 ( .A1(n6986), .A2(n6987), .ZN(n7077) );
  XNOR2_X1 U6136 ( .A(n7075), .B(n7076), .ZN(n6986) );
  OAI21_X1 U6137 ( .B1(n6776), .B2(n4388), .A(n4771), .ZN(n6907) );
  OR2_X2 U6138 ( .A1(n8703), .A2(n8704), .ZN(n4782) );
  NAND2_X1 U6139 ( .A1(n5440), .A2(n5439), .ZN(n5458) );
  NAND2_X1 U6140 ( .A1(n5377), .A2(n4801), .ZN(n4800) );
  NAND2_X1 U6141 ( .A1(n5512), .A2(n4813), .ZN(n4812) );
  NAND3_X1 U6142 ( .A1(n5301), .A2(n4818), .A3(n5302), .ZN(n4816) );
  NAND3_X1 U6143 ( .A1(n5301), .A2(n5302), .A3(n4820), .ZN(n4821) );
  NAND2_X1 U6144 ( .A1(n4821), .A2(n5316), .ZN(n5335) );
  NAND2_X1 U6145 ( .A1(n5259), .A2(n4831), .ZN(n4826) );
  OAI21_X1 U6146 ( .B1(n5259), .B2(n4830), .A(n4827), .ZN(n5300) );
  AOI21_X1 U6147 ( .B1(n4839), .B2(n4838), .A(n4837), .ZN(n4836) );
  OAI21_X1 U6148 ( .B1(n7311), .B2(n5559), .A(n9337), .ZN(n7200) );
  NAND2_X1 U6149 ( .A1(n7328), .A2(n9346), .ZN(n4850) );
  NAND2_X1 U6150 ( .A1(n9620), .A2(n4862), .ZN(n5580) );
  NAND2_X2 U6151 ( .A1(n7714), .A2(n4865), .ZN(n7853) );
  NAND2_X1 U6152 ( .A1(n4869), .A2(n7816), .ZN(n4867) );
  INV_X1 U6153 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n4868) );
  XNOR2_X1 U6154 ( .A(n7764), .B(P2_B_REG_SCAN_IN), .ZN(n4869) );
  NAND2_X1 U6155 ( .A1(n8303), .A2(n4873), .ZN(n4871) );
  NAND2_X1 U6156 ( .A1(n7725), .A2(n4880), .ZN(n4876) );
  NOR2_X1 U6157 ( .A1(n7819), .A2(n4883), .ZN(n7822) );
  INV_X1 U6158 ( .A(n8597), .ZN(n4882) );
  NAND2_X1 U6159 ( .A1(n7820), .A2(n8598), .ZN(n4884) );
  NAND2_X1 U6160 ( .A1(n8241), .A2(n4400), .ZN(n8310) );
  NAND2_X1 U6161 ( .A1(n8201), .A2(n4885), .ZN(n8279) );
  NAND2_X1 U6162 ( .A1(n8279), .A2(n8290), .ZN(n8207) );
  OR2_X1 U6163 ( .A1(n8202), .A2(n8203), .ZN(n4887) );
  OAI22_X1 U6164 ( .A1(n7150), .A2(n4894), .B1(n8605), .B2(n7149), .ZN(n4893)
         );
  AND2_X2 U6165 ( .A1(n4892), .A2(n4890), .ZN(n7249) );
  INV_X1 U6166 ( .A(n4895), .ZN(n6949) );
  NAND2_X1 U6167 ( .A1(n6951), .A2(n6950), .ZN(n4894) );
  NAND3_X1 U6168 ( .A1(n6513), .A2(n4896), .A3(n5914), .ZN(n5978) );
  NOR2_X1 U6169 ( .A1(n6429), .A2(n6428), .ZN(n6438) );
  OAI21_X1 U6170 ( .B1(n6423), .B2(n10150), .A(n6422), .ZN(n6425) );
  INV_X2 U6171 ( .A(n6865), .ZN(n8420) );
  NAND2_X1 U6172 ( .A1(n5931), .A2(n5930), .ZN(n9054) );
  NAND2_X1 U6173 ( .A1(n5300), .A2(n5299), .ZN(n5301) );
  NAND2_X1 U6174 ( .A1(n5255), .A2(n5254), .ZN(n5259) );
  NAND2_X1 U6175 ( .A1(n5504), .A2(n5503), .ZN(n5512) );
  INV_X1 U6176 ( .A(n6298), .ZN(n6752) );
  NOR2_X1 U6177 ( .A1(n8556), .A2(n8555), .ZN(n8564) );
  OAI21_X1 U6178 ( .B1(n8357), .B2(n8356), .A(n8355), .ZN(n8361) );
  NAND2_X1 U6179 ( .A1(n4979), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n4937) );
  INV_X1 U6180 ( .A(n5252), .ZN(n5255) );
  XNOR2_X1 U6181 ( .A(n8175), .B(SI_29_), .ZN(n8185) );
  INV_X1 U6182 ( .A(n6093), .ZN(n6094) );
  NAND2_X1 U6183 ( .A1(n6094), .A2(n5920), .ZN(n6137) );
  NAND2_X1 U6184 ( .A1(n6975), .A2(n9380), .ZN(n6974) );
  OR2_X1 U6185 ( .A1(n4931), .A2(n9844), .ZN(n4932) );
  CLKBUF_X1 U6186 ( .A(n6725), .Z(n8760) );
  AOI22_X2 U6187 ( .A1(n7853), .A2(n7723), .B1(n7722), .B2(n7721), .ZN(n7725)
         );
  NOR2_X1 U6188 ( .A1(n5190), .A2(n5189), .ZN(n4897) );
  AND3_X1 U6189 ( .A1(n8144), .A2(n5945), .A3(n6394), .ZN(n4898) );
  AND2_X1 U6190 ( .A1(n7226), .A2(n5733), .ZN(n4899) );
  AND2_X1 U6191 ( .A1(n5894), .A2(n4912), .ZN(n4900) );
  AND2_X1 U6192 ( .A1(n8249), .A2(n8788), .ZN(n4901) );
  INV_X1 U6193 ( .A(n9348), .ZN(n5569) );
  INV_X1 U6194 ( .A(n5590), .ZN(n9623) );
  AND2_X1 U6195 ( .A1(n5703), .A2(n7182), .ZN(n4902) );
  OR2_X1 U6196 ( .A1(n7796), .A2(n7717), .ZN(n4904) );
  OR2_X1 U6197 ( .A1(n6439), .A2(n5686), .ZN(n4905) );
  NAND2_X1 U6198 ( .A1(n8164), .A2(n9777), .ZN(n4906) );
  NAND2_X1 U6199 ( .A1(n8164), .A2(n9832), .ZN(n4907) );
  AND2_X1 U6200 ( .A1(n5669), .A2(n5668), .ZN(n4908) );
  AND2_X1 U6201 ( .A1(n9061), .A2(n9062), .ZN(n4909) );
  OR2_X1 U6202 ( .A1(n9812), .A2(n9445), .ZN(n4910) );
  AND3_X1 U6203 ( .A1(n5897), .A2(n5896), .A3(n9865), .ZN(n4911) );
  NOR2_X1 U6204 ( .A1(n5896), .A2(n9188), .ZN(n4912) );
  NAND2_X1 U6205 ( .A1(n9363), .A2(n9241), .ZN(n9242) );
  INV_X1 U6206 ( .A(n8562), .ZN(n8563) );
  NAND2_X1 U6207 ( .A1(n8564), .A2(n8563), .ZN(n8566) );
  INV_X1 U6208 ( .A(n5942), .ZN(n5929) );
  NAND2_X1 U6209 ( .A1(n6564), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6551) );
  INV_X1 U6210 ( .A(n7517), .ZN(n7518) );
  INV_X1 U6211 ( .A(n8603), .ZN(n7463) );
  OAI21_X1 U6212 ( .B1(n6564), .B2(P2_REG2_REG_2__SCAN_IN), .A(n6551), .ZN(
        n6555) );
  INV_X1 U6213 ( .A(n7519), .ZN(n7398) );
  INV_X1 U6214 ( .A(n8501), .ZN(n6335) );
  NOR2_X1 U6215 ( .A1(n9010), .A2(n8816), .ZN(n6342) );
  AND2_X1 U6216 ( .A1(n5924), .A2(n6059), .ZN(n5925) );
  AND2_X1 U6217 ( .A1(n7973), .A2(n7974), .ZN(n5768) );
  INV_X1 U6218 ( .A(n5431), .ZN(n5429) );
  INV_X1 U6219 ( .A(n5394), .ZN(n5393) );
  INV_X1 U6220 ( .A(n5266), .ZN(n5264) );
  OR2_X1 U6221 ( .A1(n9343), .A2(n5566), .ZN(n9341) );
  AND2_X1 U6222 ( .A1(n8170), .A2(n8166), .ZN(n5664) );
  INV_X1 U6223 ( .A(n8227), .ZN(n8200) );
  INV_X1 U6224 ( .A(n6243), .ZN(n6242) );
  INV_X1 U6225 ( .A(n8808), .ZN(n8802) );
  INV_X1 U6226 ( .A(n5934), .ZN(n5931) );
  INV_X1 U6227 ( .A(n5801), .ZN(n5802) );
  INV_X1 U6228 ( .A(n5784), .ZN(n5786) );
  INV_X1 U6229 ( .A(n5490), .ZN(n5489) );
  OR2_X1 U6230 ( .A1(n5468), .A2(n9118), .ZN(n5490) );
  OR2_X1 U6231 ( .A1(n5383), .A2(n5382), .ZN(n5394) );
  NAND2_X1 U6232 ( .A1(n5173), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5199) );
  NAND2_X1 U6233 ( .A1(n5393), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n5431) );
  NAND2_X1 U6234 ( .A1(n5264), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5286) );
  OR2_X1 U6235 ( .A1(n5199), .A2(n5198), .ZN(n5223) );
  AND2_X1 U6236 ( .A1(n5948), .A2(n5947), .ZN(n5951) );
  NAND2_X1 U6237 ( .A1(n8570), .A2(n8371), .ZN(n8558) );
  INV_X1 U6238 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n6421) );
  INV_X1 U6239 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n6404) );
  NAND2_X1 U6240 ( .A1(n6107), .A2(n6106), .ZN(n7654) );
  INV_X1 U6241 ( .A(n8601), .ZN(n7716) );
  OR2_X1 U6242 ( .A1(n6743), .A2(n8552), .ZN(n8858) );
  NAND2_X1 U6243 ( .A1(n6181), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6183) );
  INV_X1 U6244 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n6059) );
  INV_X1 U6245 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n6003) );
  NOR2_X1 U6246 ( .A1(n5599), .A2(n7799), .ZN(n5606) );
  AND2_X1 U6247 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5026) );
  NAND2_X1 U6248 ( .A1(n5348), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n5383) );
  AND2_X1 U6249 ( .A1(n6504), .A2(n9899), .ZN(n9291) );
  AND2_X1 U6250 ( .A1(n9362), .A2(n9238), .ZN(n9402) );
  INV_X1 U6251 ( .A(n9296), .ZN(n5677) );
  INV_X1 U6252 ( .A(n9400), .ZN(n5294) );
  NAND2_X1 U6253 ( .A1(n5013), .A2(n6447), .ZN(n5052) );
  OR2_X1 U6254 ( .A1(n8771), .A2(n6285), .ZN(n7410) );
  AND2_X1 U6255 ( .A1(n6190), .A2(n6189), .ZN(n8334) );
  INV_X1 U6256 ( .A(n6568), .ZN(n8584) );
  INV_X1 U6257 ( .A(n8860), .ZN(n8899) );
  INV_X1 U6258 ( .A(n9044), .ZN(n9033) );
  OAI21_X1 U6259 ( .B1(n9596), .B2(n9863), .A(n6434), .ZN(n6435) );
  OR3_X1 U6260 ( .A1(n5528), .A2(n5527), .A3(n5906), .ZN(n8162) );
  INV_X1 U6261 ( .A(n9376), .ZN(n9549) );
  INV_X1 U6262 ( .A(n9671), .ZN(n9960) );
  INV_X1 U6263 ( .A(n9716), .ZN(n9953) );
  AND2_X1 U6264 ( .A1(n10068), .A2(n9993), .ZN(n9777) );
  OR2_X1 U6265 ( .A1(n5607), .A2(P1_U3086), .ZN(n9292) );
  XNOR2_X1 U6266 ( .A(n5048), .B(SI_5_), .ZN(n5046) );
  AND2_X1 U6267 ( .A1(n6723), .A2(n6722), .ZN(n8258) );
  AND2_X1 U6268 ( .A1(n6734), .A2(n6733), .ZN(n8353) );
  INV_X1 U6269 ( .A(n7717), .ZN(n8600) );
  INV_X1 U6270 ( .A(n10152), .ZN(n10150) );
  INV_X1 U6271 ( .A(n6406), .ZN(n6407) );
  INV_X1 U6272 ( .A(n8238), .ZN(n9017) );
  INV_X1 U6273 ( .A(n6564), .ZN(n6583) );
  NOR2_X1 U6274 ( .A1(n4911), .A2(n5910), .ZN(n5911) );
  INV_X1 U6275 ( .A(n6435), .ZN(n6436) );
  OR2_X1 U6276 ( .A1(n4334), .A2(n7044), .ZN(n9716) );
  INV_X1 U6277 ( .A(n10068), .ZN(n10066) );
  INV_X1 U6278 ( .A(n9611), .ZN(n9817) );
  INV_X1 U6279 ( .A(n10049), .ZN(n10047) );
  INV_X1 U6280 ( .A(n5670), .ZN(n9295) );
  INV_X1 U6281 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6455) );
  NOR2_X1 U6282 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n4917) );
  NOR2_X1 U6283 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n4916) );
  NOR2_X1 U6284 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n4915) );
  NOR2_X1 U6285 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n4914) );
  INV_X1 U6286 ( .A(n5538), .ZN(n4922) );
  NOR2_X1 U6287 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n4921) );
  NAND4_X1 U6288 ( .A1(n4922), .A2(n4921), .A3(n5602), .A4(n5546), .ZN(n4925)
         );
  INV_X1 U6289 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n4923) );
  NAND4_X1 U6290 ( .A1(n4765), .A2(n5343), .A3(n5600), .A4(n4923), .ZN(n4924)
         );
  INV_X1 U6291 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n4929) );
  XNOR2_X2 U6292 ( .A(n4932), .B(n4928), .ZN(n4934) );
  NAND2_X2 U6293 ( .A1(n9848), .A2(n4934), .ZN(n4980) );
  INV_X1 U6294 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n4933) );
  OR2_X1 U6295 ( .A1(n4980), .A2(n4933), .ZN(n4940) );
  INV_X1 U6296 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n9470) );
  NAND2_X2 U6297 ( .A1(n4934), .A2(n4936), .ZN(n4982) );
  NAND2_X1 U6298 ( .A1(n4935), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n4938) );
  NAND2_X1 U6299 ( .A1(n4941), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5595) );
  NAND2_X1 U6300 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_26__SCAN_IN), 
        .ZN(n4942) );
  NAND2_X1 U6301 ( .A1(n5595), .A2(n4942), .ZN(n4943) );
  NAND2_X1 U6302 ( .A1(n4944), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4946) );
  INV_X1 U6303 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n4945) );
  BUF_X4 U6304 ( .A(n4331), .Z(n6447) );
  INV_X1 U6305 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6445) );
  INV_X1 U6306 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6451) );
  AND2_X1 U6307 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n4948) );
  NAND2_X1 U6308 ( .A1(n4332), .A2(n4948), .ZN(n4955) );
  NAND3_X1 U6309 ( .A1(n8358), .A2(SI_0_), .A3(P1_DATAO_REG_0__SCAN_IN), .ZN(
        n4949) );
  NAND2_X1 U6310 ( .A1(n4955), .A2(n4949), .ZN(n4966) );
  XNOR2_X1 U6311 ( .A(n4967), .B(n4966), .ZN(n6452) );
  AND2_X2 U6312 ( .A1(n5013), .A2(n8358), .ZN(n4997) );
  NAND2_X1 U6313 ( .A1(n4997), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4951) );
  NAND2_X1 U6314 ( .A1(n4957), .A2(n5672), .ZN(n5552) );
  INV_X1 U6315 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n4952) );
  INV_X1 U6316 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n7190) );
  INV_X1 U6317 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n5686) );
  INV_X1 U6318 ( .A(SI_0_), .ZN(n4954) );
  INV_X1 U6319 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n4953) );
  OAI21_X1 U6320 ( .B1(n8358), .B2(n4954), .A(n4953), .ZN(n4956) );
  AND2_X1 U6321 ( .A1(n4956), .A2(n4955), .ZN(n9854) );
  MUX2_X1 U6322 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9854), .S(n5013), .Z(n7182) );
  NAND2_X1 U6323 ( .A1(n6695), .A2(n7182), .ZN(n7036) );
  NAND2_X1 U6324 ( .A1(n7038), .A2(n7036), .ZN(n4959) );
  NAND2_X1 U6325 ( .A1(n4957), .A2(n9970), .ZN(n4958) );
  NAND2_X1 U6326 ( .A1(n4959), .A2(n4958), .ZN(n6972) );
  INV_X1 U6327 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n4960) );
  OR2_X1 U6328 ( .A1(n4984), .A2(n4960), .ZN(n4965) );
  INV_X1 U6329 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n7193) );
  OR2_X1 U6330 ( .A1(n4980), .A2(n7193), .ZN(n4964) );
  INV_X1 U6331 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n4961) );
  OR2_X1 U6332 ( .A1(n4982), .A2(n4961), .ZN(n4963) );
  NAND2_X1 U6333 ( .A1(n4979), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n4962) );
  NAND2_X1 U6334 ( .A1(n4967), .A2(n4966), .ZN(n4971) );
  INV_X1 U6335 ( .A(n4968), .ZN(n4969) );
  NAND2_X1 U6336 ( .A1(n4969), .A2(SI_1_), .ZN(n4970) );
  NAND2_X1 U6337 ( .A1(n4971), .A2(n4970), .ZN(n4990) );
  INV_X1 U6338 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6446) );
  INV_X1 U6339 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n4972) );
  MUX2_X1 U6340 ( .A(n6446), .B(n4972), .S(n4332), .Z(n4991) );
  XNOR2_X1 U6341 ( .A(n4991), .B(SI_2_), .ZN(n4989) );
  XNOR2_X1 U6342 ( .A(n4990), .B(n4989), .ZN(n6450) );
  NAND2_X1 U6343 ( .A1(n4997), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n4976) );
  NAND2_X1 U6344 ( .A1(n5345), .A2(n9891), .ZN(n4975) );
  XNOR2_X1 U6345 ( .A(n9468), .B(n9336), .ZN(n5553) );
  NAND2_X1 U6346 ( .A1(n6972), .A2(n5553), .ZN(n4978) );
  INV_X1 U6347 ( .A(n9468), .ZN(n6874) );
  NAND2_X1 U6348 ( .A1(n6874), .A2(n9336), .ZN(n4977) );
  NAND2_X1 U6349 ( .A1(n4978), .A2(n4977), .ZN(n7301) );
  NAND2_X1 U6350 ( .A1(n4979), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n4988) );
  INV_X1 U6351 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n4981) );
  OR2_X1 U6352 ( .A1(n4980), .A2(n4981), .ZN(n4987) );
  INV_X1 U6353 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n4983) );
  OR2_X1 U6354 ( .A1(n4984), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n4985) );
  NAND2_X1 U6355 ( .A1(n4990), .A2(n4989), .ZN(n4994) );
  INV_X1 U6356 ( .A(n4991), .ZN(n4992) );
  NAND2_X1 U6357 ( .A1(n4992), .A2(SI_2_), .ZN(n4993) );
  INV_X1 U6358 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6453) );
  INV_X1 U6359 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n4996) );
  MUX2_X1 U6360 ( .A(n6453), .B(n4996), .S(n4331), .Z(n5017) );
  XNOR2_X1 U6361 ( .A(n5017), .B(SI_3_), .ZN(n5015) );
  XNOR2_X1 U6362 ( .A(n5016), .B(n5015), .ZN(n8184) );
  NAND2_X1 U6363 ( .A1(n5465), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n5001) );
  NAND2_X1 U6364 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n4364), .ZN(n4999) );
  XNOR2_X1 U6365 ( .A(n4999), .B(P1_IR_REG_3__SCAN_IN), .ZN(n8182) );
  NAND2_X1 U6366 ( .A1(n5345), .A2(n8182), .ZN(n5000) );
  OAI211_X1 U6367 ( .C1(n5052), .C2(n8184), .A(n5001), .B(n5000), .ZN(n7302)
         );
  XNOR2_X1 U6368 ( .A(n9467), .B(n9976), .ZN(n9384) );
  NAND2_X1 U6369 ( .A1(n7301), .A2(n9384), .ZN(n5003) );
  INV_X1 U6370 ( .A(n9467), .ZN(n5555) );
  NAND2_X1 U6371 ( .A1(n5555), .A2(n9976), .ZN(n5002) );
  NAND2_X1 U6372 ( .A1(n5003), .A2(n5002), .ZN(n7315) );
  NAND2_X1 U6373 ( .A1(n4935), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5012) );
  INV_X1 U6374 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n5004) );
  OR2_X1 U6375 ( .A1(n5290), .A2(n5004), .ZN(n5011) );
  INV_X1 U6376 ( .A(n5026), .ZN(n5007) );
  INV_X1 U6377 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n7306) );
  INV_X1 U6378 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n5005) );
  NAND2_X1 U6379 ( .A1(n7306), .A2(n5005), .ZN(n5006) );
  NAND2_X1 U6380 ( .A1(n5007), .A2(n5006), .ZN(n7322) );
  INV_X1 U6381 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n5008) );
  OR2_X1 U6382 ( .A1(n4980), .A2(n5008), .ZN(n5009) );
  INV_X1 U6383 ( .A(n9466), .ZN(n6873) );
  OR2_X1 U6384 ( .A1(n5014), .A2(n9844), .ZN(n5039) );
  XNOR2_X1 U6385 ( .A(n5039), .B(P1_IR_REG_4__SCAN_IN), .ZN(n9910) );
  INV_X1 U6386 ( .A(n9910), .ZN(n6457) );
  NAND2_X1 U6387 ( .A1(n5016), .A2(n5015), .ZN(n5020) );
  INV_X1 U6388 ( .A(n5017), .ZN(n5018) );
  NAND2_X1 U6389 ( .A1(n5018), .A2(SI_3_), .ZN(n5019) );
  MUX2_X1 U6390 ( .A(n6454), .B(n6455), .S(n6447), .Z(n5033) );
  XNOR2_X1 U6391 ( .A(n5032), .B(n5031), .ZN(n6456) );
  OR2_X1 U6392 ( .A1(n6456), .A2(n5052), .ZN(n5022) );
  NAND2_X1 U6393 ( .A1(n5465), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n5021) );
  OAI211_X1 U6394 ( .C1(n5013), .C2(n6457), .A(n5022), .B(n5021), .ZN(n7317)
         );
  NAND2_X1 U6395 ( .A1(n6873), .A2(n7317), .ZN(n5558) );
  NAND2_X1 U6396 ( .A1(n9466), .A2(n9985), .ZN(n9337) );
  NAND2_X1 U6397 ( .A1(n5558), .A2(n9337), .ZN(n7316) );
  NAND2_X1 U6398 ( .A1(n7315), .A2(n7316), .ZN(n5024) );
  NAND2_X1 U6399 ( .A1(n6873), .A2(n9985), .ZN(n5023) );
  NAND2_X1 U6400 ( .A1(n5024), .A2(n5023), .ZN(n7199) );
  NAND2_X1 U6401 ( .A1(n6530), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5030) );
  INV_X1 U6402 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n5025) );
  OR2_X1 U6403 ( .A1(n4982), .A2(n5025), .ZN(n5029) );
  OAI21_X1 U6404 ( .B1(n5026), .B2(P1_REG3_REG_5__SCAN_IN), .A(n5059), .ZN(
        n7206) );
  OR2_X1 U6405 ( .A1(n4984), .A2(n7206), .ZN(n5028) );
  INV_X1 U6406 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n7207) );
  OR2_X1 U6407 ( .A1(n4980), .A2(n7207), .ZN(n5027) );
  INV_X1 U6408 ( .A(n9465), .ZN(n5044) );
  NAND2_X1 U6409 ( .A1(n5032), .A2(n5031), .ZN(n5036) );
  INV_X1 U6410 ( .A(n5033), .ZN(n5034) );
  NAND2_X1 U6411 ( .A1(n5034), .A2(SI_4_), .ZN(n5035) );
  NAND2_X1 U6412 ( .A1(n5036), .A2(n5035), .ZN(n5047) );
  INV_X1 U6413 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6460) );
  INV_X1 U6414 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n5037) );
  MUX2_X1 U6415 ( .A(n6460), .B(n5037), .S(n6447), .Z(n5048) );
  XNOR2_X1 U6416 ( .A(n5047), .B(n5046), .ZN(n6459) );
  OR2_X1 U6417 ( .A1(n6459), .A2(n5052), .ZN(n5043) );
  INV_X1 U6418 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5038) );
  NAND2_X1 U6419 ( .A1(n5039), .A2(n5038), .ZN(n5040) );
  NAND2_X1 U6420 ( .A1(n5040), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5041) );
  AOI22_X1 U6421 ( .A1(n5465), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n5345), .B2(
        n6658), .ZN(n5042) );
  NAND2_X1 U6422 ( .A1(n5043), .A2(n5042), .ZN(n9992) );
  NAND2_X1 U6423 ( .A1(n5044), .A2(n9992), .ZN(n5560) );
  INV_X1 U6424 ( .A(n9992), .ZN(n7205) );
  NAND2_X1 U6425 ( .A1(n7205), .A2(n9465), .ZN(n9338) );
  NAND2_X1 U6426 ( .A1(n5560), .A2(n9338), .ZN(n9383) );
  NAND2_X1 U6427 ( .A1(n5044), .A2(n7205), .ZN(n5045) );
  NAND2_X1 U6428 ( .A1(n5047), .A2(n5046), .ZN(n5051) );
  INV_X1 U6429 ( .A(n5048), .ZN(n5049) );
  NAND2_X1 U6430 ( .A1(n5049), .A2(SI_5_), .ZN(n5050) );
  NAND2_X1 U6431 ( .A1(n5051), .A2(n5050), .ZN(n5068) );
  MUX2_X1 U6432 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n6447), .Z(n5069) );
  XNOR2_X1 U6433 ( .A(n5068), .B(n5066), .ZN(n6463) );
  NAND2_X1 U6434 ( .A1(n6463), .A2(n5114), .ZN(n5056) );
  OR2_X1 U6435 ( .A1(n5053), .A2(n9844), .ZN(n5054) );
  XNOR2_X1 U6436 ( .A(n5054), .B(P1_IR_REG_6__SCAN_IN), .ZN(n6669) );
  AOI22_X1 U6437 ( .A1(n5465), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n5345), .B2(
        n6669), .ZN(n5055) );
  NAND2_X1 U6438 ( .A1(n5056), .A2(n5055), .ZN(n7179) );
  NAND2_X1 U6439 ( .A1(n4979), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5065) );
  INV_X1 U6440 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n5057) );
  OR2_X1 U6441 ( .A1(n4980), .A2(n5057), .ZN(n5064) );
  AND2_X1 U6442 ( .A1(n5059), .A2(n5058), .ZN(n5060) );
  OR2_X1 U6443 ( .A1(n5060), .A2(n5077), .ZN(n7231) );
  OR2_X1 U6444 ( .A1(n4984), .A2(n7231), .ZN(n5063) );
  INV_X1 U6445 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n5061) );
  OR2_X1 U6446 ( .A1(n4982), .A2(n5061), .ZN(n5062) );
  NAND4_X1 U6447 ( .A1(n5065), .A2(n5064), .A3(n5063), .A4(n5062), .ZN(n9464)
         );
  INV_X1 U6448 ( .A(n9464), .ZN(n5565) );
  XNOR2_X1 U6449 ( .A(n7179), .B(n5565), .ZN(n7174) );
  NAND2_X1 U6450 ( .A1(n5068), .A2(n5067), .ZN(n5071) );
  NAND2_X1 U6451 ( .A1(n5069), .A2(SI_6_), .ZN(n5070) );
  MUX2_X1 U6452 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n6447), .Z(n5089) );
  XNOR2_X1 U6453 ( .A(n5088), .B(n5086), .ZN(n6468) );
  NAND2_X1 U6454 ( .A1(n6468), .A2(n5114), .ZN(n5075) );
  INV_X1 U6455 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5072) );
  NAND2_X1 U6456 ( .A1(n5053), .A2(n5072), .ZN(n5096) );
  NAND2_X1 U6457 ( .A1(n5096), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5073) );
  XNOR2_X1 U6458 ( .A(n5073), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6798) );
  AOI22_X1 U6459 ( .A1(n5465), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n5345), .B2(
        n6798), .ZN(n5074) );
  NAND2_X1 U6460 ( .A1(n4979), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5083) );
  INV_X1 U6461 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n5076) );
  OR2_X1 U6462 ( .A1(n4980), .A2(n5076), .ZN(n5082) );
  NOR2_X1 U6463 ( .A1(n5077), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5078) );
  OR2_X1 U6464 ( .A1(n5100), .A2(n5078), .ZN(n9950) );
  OR2_X1 U6465 ( .A1(n4984), .A2(n9950), .ZN(n5081) );
  INV_X1 U6466 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n5079) );
  OR2_X1 U6467 ( .A1(n4982), .A2(n5079), .ZN(n5080) );
  NAND4_X1 U6468 ( .A1(n5083), .A2(n5082), .A3(n5081), .A4(n5080), .ZN(n9463)
         );
  INV_X1 U6469 ( .A(n9463), .ZN(n5563) );
  XNOR2_X1 U6470 ( .A(n9954), .B(n5563), .ZN(n9946) );
  NAND2_X1 U6471 ( .A1(n9943), .A2(n9946), .ZN(n5085) );
  OR2_X1 U6472 ( .A1(n9954), .A2(n9463), .ZN(n5084) );
  NAND2_X1 U6473 ( .A1(n5085), .A2(n5084), .ZN(n7376) );
  NAND2_X1 U6474 ( .A1(n5089), .A2(SI_7_), .ZN(n5090) );
  INV_X1 U6475 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6479) );
  INV_X1 U6476 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n5091) );
  MUX2_X1 U6477 ( .A(n6479), .B(n5091), .S(n6447), .Z(n5093) );
  INV_X1 U6478 ( .A(SI_8_), .ZN(n5092) );
  INV_X1 U6479 ( .A(n5093), .ZN(n5094) );
  NAND2_X1 U6480 ( .A1(n5094), .A2(SI_8_), .ZN(n5095) );
  NAND2_X1 U6481 ( .A1(n6472), .A2(n5114), .ZN(n5098) );
  NAND2_X1 U6482 ( .A1(n5142), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5115) );
  XNOR2_X1 U6483 ( .A(n5115), .B(P1_IR_REG_8__SCAN_IN), .ZN(n6886) );
  AOI22_X1 U6484 ( .A1(n5465), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n5345), .B2(
        n6886), .ZN(n5097) );
  NAND2_X2 U6485 ( .A1(n5098), .A2(n5097), .ZN(n7495) );
  NAND2_X1 U6486 ( .A1(n4979), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5106) );
  INV_X1 U6487 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n5099) );
  OR2_X1 U6488 ( .A1(n4980), .A2(n5099), .ZN(n5105) );
  NOR2_X1 U6489 ( .A1(n5100), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5101) );
  OR2_X1 U6490 ( .A1(n5121), .A2(n5101), .ZN(n7493) );
  OR2_X1 U6491 ( .A1(n4984), .A2(n7493), .ZN(n5104) );
  INV_X1 U6492 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n5102) );
  OR2_X1 U6493 ( .A1(n4982), .A2(n5102), .ZN(n5103) );
  NAND4_X1 U6494 ( .A1(n5106), .A2(n5105), .A3(n5104), .A4(n5103), .ZN(n9462)
         );
  INV_X1 U6495 ( .A(n9462), .ZN(n7418) );
  NAND2_X1 U6496 ( .A1(n7495), .A2(n7418), .ZN(n9205) );
  NAND2_X1 U6497 ( .A1(n7415), .A2(n9205), .ZN(n7377) );
  NAND2_X1 U6498 ( .A1(n7376), .A2(n7377), .ZN(n5108) );
  OR2_X1 U6499 ( .A1(n7495), .A2(n9462), .ZN(n5107) );
  NAND2_X1 U6500 ( .A1(n5108), .A2(n5107), .ZN(n7420) );
  INV_X1 U6501 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6498) );
  INV_X1 U6502 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n5109) );
  MUX2_X1 U6503 ( .A(n6498), .B(n5109), .S(n6447), .Z(n5111) );
  INV_X1 U6504 ( .A(SI_9_), .ZN(n5110) );
  NAND2_X1 U6505 ( .A1(n5111), .A2(n5110), .ZN(n5132) );
  INV_X1 U6506 ( .A(n5111), .ZN(n5112) );
  AND2_X1 U6507 ( .A1(n5132), .A2(n5156), .ZN(n5113) );
  NAND2_X1 U6508 ( .A1(n6484), .A2(n5114), .ZN(n5119) );
  INV_X1 U6509 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5139) );
  NAND2_X1 U6510 ( .A1(n5115), .A2(n5139), .ZN(n5116) );
  NAND2_X1 U6511 ( .A1(n5116), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5117) );
  XNOR2_X1 U6512 ( .A(n5117), .B(P1_IR_REG_9__SCAN_IN), .ZN(n7022) );
  AOI22_X1 U6513 ( .A1(n4997), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n5345), .B2(
        n7022), .ZN(n5118) );
  NAND2_X1 U6514 ( .A1(n6530), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5126) );
  INV_X1 U6515 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n5120) );
  OR2_X1 U6516 ( .A1(n4982), .A2(n5120), .ZN(n5125) );
  OR2_X1 U6517 ( .A1(n5121), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n5122) );
  NAND2_X1 U6518 ( .A1(n5148), .A2(n5122), .ZN(n7542) );
  OR2_X1 U6519 ( .A1(n4984), .A2(n7542), .ZN(n5124) );
  INV_X1 U6520 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n7424) );
  OR2_X1 U6521 ( .A1(n4980), .A2(n7424), .ZN(n5123) );
  NAND4_X1 U6522 ( .A1(n5126), .A2(n5125), .A3(n5124), .A4(n5123), .ZN(n9461)
         );
  INV_X1 U6523 ( .A(n9461), .ZN(n5127) );
  NAND2_X1 U6524 ( .A1(n10017), .A2(n5127), .ZN(n9208) );
  NAND2_X1 U6525 ( .A1(n9214), .A2(n9208), .ZN(n9391) );
  OR2_X1 U6526 ( .A1(n10017), .A2(n9461), .ZN(n5128) );
  INV_X1 U6527 ( .A(n5156), .ZN(n5134) );
  OR2_X1 U6528 ( .A1(n5129), .A2(n5134), .ZN(n5130) );
  OR2_X1 U6529 ( .A1(n5131), .A2(n5130), .ZN(n5136) );
  OR2_X1 U6530 ( .A1(n5134), .A2(n5155), .ZN(n5135) );
  NAND2_X1 U6531 ( .A1(n5136), .A2(n5135), .ZN(n5138) );
  MUX2_X1 U6532 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .S(n6447), .Z(n5158) );
  INV_X1 U6533 ( .A(n5157), .ZN(n5137) );
  NAND2_X1 U6534 ( .A1(n6480), .A2(n5114), .ZN(n5145) );
  INV_X1 U6535 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n5140) );
  NAND2_X1 U6536 ( .A1(n5140), .A2(n5139), .ZN(n5141) );
  NOR2_X1 U6537 ( .A1(n5142), .A2(n5141), .ZN(n5169) );
  OR2_X1 U6538 ( .A1(n5169), .A2(n9844), .ZN(n5143) );
  XNOR2_X1 U6539 ( .A(n5143), .B(P1_IR_REG_10__SCAN_IN), .ZN(n7266) );
  AOI22_X1 U6540 ( .A1(n4997), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5345), .B2(
        n7266), .ZN(n5144) );
  NAND2_X1 U6541 ( .A1(n5145), .A2(n5144), .ZN(n7338) );
  NAND2_X1 U6542 ( .A1(n6530), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5153) );
  INV_X1 U6543 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n5146) );
  OR2_X1 U6544 ( .A1(n4982), .A2(n5146), .ZN(n5152) );
  INV_X1 U6545 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7335) );
  OR2_X1 U6546 ( .A1(n4980), .A2(n7335), .ZN(n5151) );
  INV_X1 U6547 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n5147) );
  NAND2_X1 U6548 ( .A1(n5148), .A2(n5147), .ZN(n5149) );
  NAND2_X1 U6549 ( .A1(n5175), .A2(n5149), .ZN(n9869) );
  OR2_X1 U6550 ( .A1(n4984), .A2(n9869), .ZN(n5150) );
  NAND4_X1 U6551 ( .A1(n5153), .A2(n5152), .A3(n5151), .A4(n5150), .ZN(n9460)
         );
  INV_X1 U6552 ( .A(n9460), .ZN(n5154) );
  NAND2_X1 U6553 ( .A1(n7338), .A2(n5154), .ZN(n9215) );
  NAND2_X1 U6554 ( .A1(n9342), .A2(n9215), .ZN(n7334) );
  INV_X1 U6555 ( .A(n7429), .ZN(n5183) );
  NAND2_X1 U6556 ( .A1(n5192), .A2(n5184), .ZN(n5161) );
  NAND2_X1 U6557 ( .A1(n5158), .A2(SI_10_), .ZN(n5159) );
  NAND2_X1 U6558 ( .A1(n5161), .A2(n5187), .ZN(n5167) );
  INV_X1 U6559 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6524) );
  INV_X1 U6560 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n5162) );
  MUX2_X1 U6561 ( .A(n6524), .B(n5162), .S(n6447), .Z(n5164) );
  INV_X1 U6562 ( .A(SI_11_), .ZN(n5163) );
  INV_X1 U6563 ( .A(n5164), .ZN(n5165) );
  NAND2_X1 U6564 ( .A1(n5165), .A2(SI_11_), .ZN(n5166) );
  NAND2_X1 U6565 ( .A1(n5185), .A2(n5166), .ZN(n5186) );
  XNOR2_X1 U6566 ( .A(n5167), .B(n5186), .ZN(n6500) );
  NAND2_X1 U6567 ( .A1(n6500), .A2(n5114), .ZN(n5172) );
  INV_X1 U6568 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5168) );
  NAND2_X1 U6569 ( .A1(n5169), .A2(n5168), .ZN(n5193) );
  NAND2_X1 U6570 ( .A1(n5193), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5170) );
  XNOR2_X1 U6571 ( .A(n5170), .B(P1_IR_REG_11__SCAN_IN), .ZN(n7346) );
  AOI22_X1 U6572 ( .A1(n4997), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5345), .B2(
        n7346), .ZN(n5171) );
  NAND2_X1 U6573 ( .A1(n6530), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5181) );
  INV_X1 U6574 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5174) );
  NAND2_X1 U6575 ( .A1(n5175), .A2(n5174), .ZN(n5176) );
  NAND2_X1 U6576 ( .A1(n5199), .A2(n5176), .ZN(n7809) );
  OR2_X1 U6577 ( .A1(n4984), .A2(n7809), .ZN(n5180) );
  INV_X1 U6578 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7446) );
  OR2_X1 U6579 ( .A1(n4980), .A2(n7446), .ZN(n5179) );
  INV_X1 U6580 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n5177) );
  OR2_X1 U6581 ( .A1(n4982), .A2(n5177), .ZN(n5178) );
  NAND4_X1 U6582 ( .A1(n5181), .A2(n5180), .A3(n5179), .A4(n5178), .ZN(n9459)
         );
  NOR2_X1 U6583 ( .A1(n7802), .A2(n9459), .ZN(n7432) );
  INV_X1 U6584 ( .A(n7432), .ZN(n5182) );
  NAND2_X1 U6585 ( .A1(n7802), .A2(n9459), .ZN(n7430) );
  INV_X1 U6586 ( .A(n5185), .ZN(n5190) );
  INV_X1 U6587 ( .A(n5186), .ZN(n5188) );
  INV_X1 U6588 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6527) );
  INV_X1 U6589 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6528) );
  MUX2_X1 U6590 ( .A(n6527), .B(n6528), .S(n6447), .Z(n5209) );
  XNOR2_X1 U6591 ( .A(n5213), .B(n5208), .ZN(n6526) );
  NAND2_X1 U6592 ( .A1(n6526), .A2(n5114), .ZN(n5196) );
  OR2_X1 U6593 ( .A1(n5193), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n5194) );
  NAND2_X1 U6594 ( .A1(n5194), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5216) );
  XNOR2_X1 U6595 ( .A(n5216), .B(P1_IR_REG_12__SCAN_IN), .ZN(n7585) );
  AOI22_X1 U6596 ( .A1(n4997), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n5345), .B2(
        n7585), .ZN(n5195) );
  NAND2_X1 U6597 ( .A1(n4935), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5204) );
  INV_X1 U6598 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n5197) );
  OR2_X1 U6599 ( .A1(n5290), .A2(n5197), .ZN(n5203) );
  INV_X1 U6600 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5198) );
  NAND2_X1 U6601 ( .A1(n5199), .A2(n5198), .ZN(n5200) );
  NAND2_X1 U6602 ( .A1(n5223), .A2(n5200), .ZN(n7972) );
  OR2_X1 U6603 ( .A1(n4984), .A2(n7972), .ZN(n5202) );
  INV_X1 U6604 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7555) );
  OR2_X1 U6605 ( .A1(n4980), .A2(n7555), .ZN(n5201) );
  NAND4_X1 U6606 ( .A1(n5204), .A2(n5203), .A3(n5202), .A4(n5201), .ZN(n9458)
         );
  INV_X1 U6607 ( .A(n9458), .ZN(n7636) );
  OR2_X1 U6608 ( .A1(n7979), .A2(n7636), .ZN(n9223) );
  NAND2_X1 U6609 ( .A1(n7979), .A2(n7636), .ZN(n9221) );
  INV_X1 U6610 ( .A(n9394), .ZN(n5205) );
  OR2_X1 U6611 ( .A1(n7979), .A2(n9458), .ZN(n5206) );
  NAND2_X1 U6612 ( .A1(n5207), .A2(n5206), .ZN(n7632) );
  INV_X1 U6613 ( .A(n5209), .ZN(n5210) );
  MUX2_X1 U6614 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n6447), .Z(n5232) );
  XNOR2_X1 U6615 ( .A(n5232), .B(SI_13_), .ZN(n5214) );
  XNOR2_X1 U6616 ( .A(n5236), .B(n5214), .ZN(n6538) );
  NAND2_X1 U6617 ( .A1(n6538), .A2(n5114), .ZN(n5220) );
  INV_X1 U6618 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5215) );
  NAND2_X1 U6619 ( .A1(n5216), .A2(n5215), .ZN(n5217) );
  NAND2_X1 U6620 ( .A1(n5217), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5218) );
  XNOR2_X1 U6621 ( .A(n5218), .B(P1_IR_REG_13__SCAN_IN), .ZN(n7682) );
  AOI22_X1 U6622 ( .A1(n4997), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n7682), .B2(
        n5345), .ZN(n5219) );
  NAND2_X1 U6623 ( .A1(n6530), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5229) );
  INV_X1 U6624 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n5221) );
  OR2_X1 U6625 ( .A1(n4980), .A2(n5221), .ZN(n5228) );
  INV_X1 U6626 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5222) );
  NAND2_X1 U6627 ( .A1(n5223), .A2(n5222), .ZN(n5224) );
  NAND2_X1 U6628 ( .A1(n5245), .A2(n5224), .ZN(n9726) );
  OR2_X1 U6629 ( .A1(n4984), .A2(n9726), .ZN(n5227) );
  INV_X1 U6630 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n5225) );
  OR2_X1 U6631 ( .A1(n4982), .A2(n5225), .ZN(n5226) );
  NAND4_X1 U6632 ( .A1(n5229), .A2(n5228), .A3(n5227), .A4(n5226), .ZN(n9457)
         );
  INV_X1 U6633 ( .A(n9457), .ZN(n5230) );
  OR2_X1 U6634 ( .A1(n9729), .A2(n5230), .ZN(n9228) );
  NAND2_X1 U6635 ( .A1(n9729), .A2(n5230), .ZN(n9348) );
  NAND2_X1 U6636 ( .A1(n9228), .A2(n9348), .ZN(n9396) );
  OR2_X1 U6637 ( .A1(n9729), .A2(n9457), .ZN(n5231) );
  INV_X1 U6638 ( .A(SI_13_), .ZN(n8067) );
  NAND2_X1 U6639 ( .A1(n5233), .A2(n8067), .ZN(n5234) );
  INV_X1 U6640 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6712) );
  INV_X1 U6641 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n6756) );
  MUX2_X1 U6642 ( .A(n6712), .B(n6756), .S(n6447), .Z(n5256) );
  XNOR2_X1 U6643 ( .A(n5256), .B(SI_14_), .ZN(n5237) );
  XNOR2_X1 U6644 ( .A(n5252), .B(n5237), .ZN(n6711) );
  NAND2_X1 U6645 ( .A1(n6711), .A2(n5114), .ZN(n5242) );
  NAND2_X1 U6646 ( .A1(n5238), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5239) );
  MUX2_X1 U6647 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5239), .S(
        P1_IR_REG_14__SCAN_IN), .Z(n5240) );
  AND2_X1 U6648 ( .A1(n5240), .A2(n5281), .ZN(n9487) );
  AOI22_X1 U6649 ( .A1(n4997), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n5345), .B2(
        n9487), .ZN(n5241) );
  NAND2_X1 U6650 ( .A1(n4935), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5250) );
  INV_X1 U6651 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n7679) );
  OR2_X1 U6652 ( .A1(n5290), .A2(n7679), .ZN(n5249) );
  INV_X1 U6653 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n5244) );
  NAND2_X1 U6654 ( .A1(n5245), .A2(n5244), .ZN(n5246) );
  NAND2_X1 U6655 ( .A1(n5266), .A2(n5246), .ZN(n9074) );
  OR2_X1 U6656 ( .A1(n4984), .A2(n9074), .ZN(n5248) );
  INV_X1 U6657 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7698) );
  OR2_X1 U6658 ( .A1(n4980), .A2(n7698), .ZN(n5247) );
  NAND4_X1 U6659 ( .A1(n5250), .A2(n5249), .A3(n5248), .A4(n5247), .ZN(n9456)
         );
  NAND2_X1 U6660 ( .A1(n9076), .A2(n9456), .ZN(n5251) );
  INV_X1 U6661 ( .A(SI_14_), .ZN(n5253) );
  NAND2_X1 U6662 ( .A1(n5256), .A2(n5253), .ZN(n5254) );
  INV_X1 U6663 ( .A(n5256), .ZN(n5257) );
  NAND2_X1 U6664 ( .A1(n5257), .A2(SI_14_), .ZN(n5258) );
  MUX2_X1 U6665 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n6447), .Z(n5278) );
  XNOR2_X1 U6666 ( .A(n5278), .B(SI_15_), .ZN(n5260) );
  XNOR2_X1 U6667 ( .A(n5277), .B(n5260), .ZN(n6852) );
  NAND2_X1 U6668 ( .A1(n6852), .A2(n5114), .ZN(n5263) );
  NAND2_X1 U6669 ( .A1(n5281), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5261) );
  XNOR2_X1 U6670 ( .A(n5261), .B(P1_IR_REG_15__SCAN_IN), .ZN(n9490) );
  AOI22_X1 U6671 ( .A1(n4997), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n5345), .B2(
        n9490), .ZN(n5262) );
  NAND2_X1 U6672 ( .A1(n4979), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5272) );
  INV_X1 U6673 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n7774) );
  OR2_X1 U6674 ( .A1(n4980), .A2(n7774), .ZN(n5271) );
  INV_X1 U6675 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n5265) );
  NAND2_X1 U6676 ( .A1(n5266), .A2(n5265), .ZN(n5267) );
  NAND2_X1 U6677 ( .A1(n5286), .A2(n5267), .ZN(n9194) );
  OR2_X1 U6678 ( .A1(n4984), .A2(n9194), .ZN(n5270) );
  INV_X1 U6679 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n5268) );
  OR2_X1 U6680 ( .A1(n4982), .A2(n5268), .ZN(n5269) );
  NAND4_X1 U6681 ( .A1(n5272), .A2(n5271), .A3(n5270), .A4(n5269), .ZN(n9455)
         );
  INV_X1 U6682 ( .A(n9455), .ZN(n5572) );
  NAND2_X1 U6683 ( .A1(n5273), .A2(n5572), .ZN(n5276) );
  INV_X1 U6684 ( .A(n7777), .ZN(n5274) );
  NAND2_X1 U6685 ( .A1(n5274), .A2(n4701), .ZN(n5275) );
  NAND2_X1 U6686 ( .A1(n5276), .A2(n5275), .ZN(n7885) );
  INV_X1 U6687 ( .A(n5278), .ZN(n5279) );
  INV_X1 U6688 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n8140) );
  INV_X1 U6689 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n6930) );
  MUX2_X1 U6690 ( .A(n8140), .B(n6930), .S(n6447), .Z(n5298) );
  XNOR2_X1 U6691 ( .A(n5298), .B(SI_16_), .ZN(n5280) );
  XNOR2_X1 U6692 ( .A(n5297), .B(n5280), .ZN(n6921) );
  NAND2_X1 U6693 ( .A1(n6921), .A2(n5114), .ZN(n5284) );
  NAND2_X1 U6694 ( .A1(n4411), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5282) );
  XNOR2_X1 U6695 ( .A(n5282), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9938) );
  AOI22_X1 U6696 ( .A1(n4997), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n5345), .B2(
        n9938), .ZN(n5283) );
  INV_X1 U6697 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n5285) );
  NAND2_X1 U6698 ( .A1(n5286), .A2(n5285), .ZN(n5287) );
  NAND2_X1 U6699 ( .A1(n5310), .A2(n5287), .ZN(n9126) );
  INV_X1 U6700 ( .A(n4980), .ZN(n5492) );
  NAND2_X1 U6701 ( .A1(n5492), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n5288) );
  OAI21_X1 U6702 ( .B1(n9126), .B2(n4984), .A(n5288), .ZN(n5292) );
  INV_X1 U6703 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9501) );
  NAND2_X1 U6704 ( .A1(n4935), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5289) );
  OAI21_X1 U6705 ( .B1(n9501), .B2(n5290), .A(n5289), .ZN(n5291) );
  OR2_X1 U6706 ( .A1(n5292), .A2(n5291), .ZN(n9454) );
  INV_X1 U6707 ( .A(n9454), .ZN(n5293) );
  NAND2_X1 U6708 ( .A1(n7890), .A2(n5293), .ZN(n9357) );
  NAND2_X1 U6709 ( .A1(n7890), .A2(n9454), .ZN(n5295) );
  INV_X1 U6710 ( .A(SI_16_), .ZN(n5296) );
  INV_X1 U6711 ( .A(n5298), .ZN(n5299) );
  INV_X1 U6712 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7014) );
  INV_X1 U6713 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n7016) );
  MUX2_X1 U6714 ( .A(n7014), .B(n7016), .S(n6447), .Z(n5303) );
  INV_X1 U6715 ( .A(SI_17_), .ZN(n8064) );
  NAND2_X1 U6716 ( .A1(n5303), .A2(n8064), .ZN(n5316) );
  INV_X1 U6717 ( .A(n5303), .ZN(n5304) );
  NAND2_X1 U6718 ( .A1(n5304), .A2(SI_17_), .ZN(n5305) );
  NAND2_X1 U6719 ( .A1(n5316), .A2(n5305), .ZN(n5317) );
  XNOR2_X1 U6720 ( .A(n5318), .B(n5317), .ZN(n7013) );
  NAND2_X1 U6721 ( .A1(n7013), .A2(n5114), .ZN(n5307) );
  NAND2_X1 U6722 ( .A1(n5537), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5320) );
  XNOR2_X1 U6723 ( .A(n5320), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9519) );
  AOI22_X1 U6724 ( .A1(n4997), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n5345), .B2(
        n9519), .ZN(n5306) );
  INV_X1 U6725 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n9504) );
  INV_X1 U6726 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n5309) );
  NAND2_X1 U6727 ( .A1(n5310), .A2(n5309), .ZN(n5311) );
  NAND2_X1 U6728 ( .A1(n5324), .A2(n5311), .ZN(n7947) );
  OR2_X1 U6729 ( .A1(n7947), .A2(n4984), .ZN(n5313) );
  AOI22_X1 U6730 ( .A1(n4935), .A2(P1_REG0_REG_17__SCAN_IN), .B1(n4979), .B2(
        P1_REG1_REG_17__SCAN_IN), .ZN(n5312) );
  OAI211_X1 U6731 ( .C1(n4980), .C2(n9504), .A(n5313), .B(n5312), .ZN(n9453)
         );
  NAND2_X1 U6732 ( .A1(n7946), .A2(n9453), .ZN(n5314) );
  NAND2_X1 U6733 ( .A1(n5315), .A2(n5314), .ZN(n9704) );
  INV_X1 U6734 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7146) );
  INV_X1 U6735 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n7103) );
  MUX2_X1 U6736 ( .A(n7146), .B(n7103), .S(n6447), .Z(n5331) );
  XNOR2_X1 U6737 ( .A(n5331), .B(SI_18_), .ZN(n5330) );
  XNOR2_X1 U6738 ( .A(n5335), .B(n5330), .ZN(n7102) );
  NAND2_X1 U6739 ( .A1(n7102), .A2(n5114), .ZN(n5323) );
  NAND2_X1 U6740 ( .A1(n5320), .A2(n5319), .ZN(n5321) );
  XNOR2_X1 U6741 ( .A(n5341), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9530) );
  AOI22_X1 U6742 ( .A1(n4997), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n5345), .B2(
        n9530), .ZN(n5322) );
  INV_X1 U6743 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n9182) );
  NAND2_X1 U6744 ( .A1(n5324), .A2(n9182), .ZN(n5325) );
  NAND2_X1 U6745 ( .A1(n5350), .A2(n5325), .ZN(n9712) );
  AOI22_X1 U6746 ( .A1(n4935), .A2(P1_REG0_REG_18__SCAN_IN), .B1(n6530), .B2(
        P1_REG1_REG_18__SCAN_IN), .ZN(n5327) );
  NAND2_X1 U6747 ( .A1(n5492), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n5326) );
  OAI211_X1 U6748 ( .C1(n9712), .C2(n4984), .A(n5327), .B(n5326), .ZN(n9452)
         );
  OR2_X1 U6749 ( .A1(n9793), .A2(n9452), .ZN(n5328) );
  NAND2_X1 U6750 ( .A1(n9793), .A2(n9452), .ZN(n5329) );
  INV_X1 U6751 ( .A(n5330), .ZN(n5334) );
  INV_X1 U6752 ( .A(n5331), .ZN(n5332) );
  NAND2_X1 U6753 ( .A1(n5332), .A2(SI_18_), .ZN(n5333) );
  INV_X1 U6754 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n8160) );
  INV_X1 U6755 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7276) );
  MUX2_X1 U6756 ( .A(n8160), .B(n7276), .S(n6447), .Z(n5337) );
  INV_X1 U6757 ( .A(SI_19_), .ZN(n5336) );
  NAND2_X1 U6758 ( .A1(n5337), .A2(n5336), .ZN(n5364) );
  INV_X1 U6759 ( .A(n5337), .ZN(n5338) );
  NAND2_X1 U6760 ( .A1(n5338), .A2(SI_19_), .ZN(n5339) );
  NAND2_X1 U6761 ( .A1(n5364), .A2(n5339), .ZN(n5361) );
  XNOR2_X1 U6762 ( .A(n5360), .B(n5361), .ZN(n7275) );
  NAND2_X1 U6763 ( .A1(n7275), .A2(n5114), .ZN(n5347) );
  NAND2_X1 U6764 ( .A1(n5341), .A2(n5340), .ZN(n5342) );
  NAND2_X1 U6765 ( .A1(n5342), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5344) );
  XNOR2_X1 U6766 ( .A(n5344), .B(n5343), .ZN(n9376) );
  AOI22_X1 U6767 ( .A1(n5465), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9549), .B2(
        n5345), .ZN(n5346) );
  INV_X1 U6768 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n5349) );
  NAND2_X1 U6769 ( .A1(n5350), .A2(n5349), .ZN(n5351) );
  NAND2_X1 U6770 ( .A1(n5383), .A2(n5351), .ZN(n9691) );
  OR2_X1 U6771 ( .A1(n9691), .A2(n4984), .ZN(n5357) );
  INV_X1 U6772 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n5354) );
  NAND2_X1 U6773 ( .A1(n6530), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n5353) );
  NAND2_X1 U6774 ( .A1(n4935), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n5352) );
  OAI211_X1 U6775 ( .C1(n5354), .C2(n4980), .A(n5353), .B(n5352), .ZN(n5355)
         );
  INV_X1 U6776 ( .A(n5355), .ZN(n5356) );
  NAND2_X1 U6777 ( .A1(n5357), .A2(n5356), .ZN(n9451) );
  OR2_X1 U6778 ( .A1(n9787), .A2(n9451), .ZN(n5358) );
  NAND2_X1 U6779 ( .A1(n5359), .A2(n5358), .ZN(n9681) );
  INV_X1 U6780 ( .A(n5361), .ZN(n5362) );
  NAND2_X1 U6781 ( .A1(n5363), .A2(n5362), .ZN(n5365) );
  MUX2_X1 U6782 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(P2_DATAO_REG_20__SCAN_IN), 
        .S(n6447), .Z(n5374) );
  INV_X1 U6783 ( .A(SI_20_), .ZN(n5376) );
  XNOR2_X1 U6784 ( .A(n5374), .B(n5376), .ZN(n5366) );
  XNOR2_X1 U6785 ( .A(n5377), .B(n5366), .ZN(n7356) );
  NAND2_X1 U6786 ( .A1(n7356), .A2(n5114), .ZN(n5368) );
  NAND2_X1 U6787 ( .A1(n5465), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n5367) );
  XNOR2_X1 U6788 ( .A(n5383), .B(P1_REG3_REG_20__SCAN_IN), .ZN(n9683) );
  INV_X1 U6789 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n7993) );
  NAND2_X1 U6790 ( .A1(n5492), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n5370) );
  NAND2_X1 U6791 ( .A1(n4979), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n5369) );
  OAI211_X1 U6792 ( .C1(n4982), .C2(n7993), .A(n5370), .B(n5369), .ZN(n5371)
         );
  AOI21_X1 U6793 ( .B1(n9683), .B2(n5516), .A(n5371), .ZN(n9107) );
  INV_X1 U6794 ( .A(n9107), .ZN(n6536) );
  OR2_X1 U6795 ( .A1(n9781), .A2(n6536), .ZN(n9246) );
  NAND2_X1 U6796 ( .A1(n9781), .A2(n6536), .ZN(n9245) );
  OR2_X1 U6797 ( .A1(n9781), .A2(n9107), .ZN(n5373) );
  INV_X1 U6798 ( .A(n5374), .ZN(n5375) );
  INV_X1 U6799 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7533) );
  INV_X1 U6800 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n8190) );
  MUX2_X1 U6801 ( .A(n7533), .B(n8190), .S(n6447), .Z(n5401) );
  XNOR2_X1 U6802 ( .A(n5401), .B(SI_21_), .ZN(n5378) );
  XNOR2_X1 U6803 ( .A(n5404), .B(n5378), .ZN(n7532) );
  NAND2_X1 U6804 ( .A1(n7532), .A2(n5114), .ZN(n5380) );
  NAND2_X1 U6805 ( .A1(n5465), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n5379) );
  INV_X1 U6806 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n9160) );
  INV_X1 U6807 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n5381) );
  OAI21_X1 U6808 ( .B1(n5383), .B2(n9160), .A(n5381), .ZN(n5384) );
  NAND2_X1 U6809 ( .A1(P1_REG3_REG_20__SCAN_IN), .A2(P1_REG3_REG_21__SCAN_IN), 
        .ZN(n5382) );
  NAND2_X1 U6810 ( .A1(n5384), .A2(n5394), .ZN(n9668) );
  OR2_X1 U6811 ( .A1(n9668), .A2(n4984), .ZN(n5390) );
  INV_X1 U6812 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n5387) );
  NAND2_X1 U6813 ( .A1(n4979), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n5386) );
  NAND2_X1 U6814 ( .A1(n4935), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5385) );
  OAI211_X1 U6815 ( .C1(n5387), .C2(n4980), .A(n5386), .B(n5385), .ZN(n5388)
         );
  INV_X1 U6816 ( .A(n5388), .ZN(n5389) );
  NAND2_X1 U6817 ( .A1(n5390), .A2(n5389), .ZN(n9450) );
  INV_X1 U6818 ( .A(n9450), .ZN(n5391) );
  OR2_X1 U6819 ( .A1(n9831), .A2(n5391), .ZN(n9304) );
  NAND2_X1 U6820 ( .A1(n9831), .A2(n5391), .ZN(n9247) );
  NAND2_X1 U6821 ( .A1(n9304), .A2(n9247), .ZN(n9662) );
  NAND2_X1 U6822 ( .A1(n9831), .A2(n9450), .ZN(n5392) );
  NAND2_X1 U6823 ( .A1(n9665), .A2(n5392), .ZN(n9646) );
  INV_X1 U6824 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9170) );
  NAND2_X1 U6825 ( .A1(n5394), .A2(n9170), .ZN(n5395) );
  NAND2_X1 U6826 ( .A1(n5431), .A2(n5395), .ZN(n9648) );
  OR2_X1 U6827 ( .A1(n9648), .A2(n4984), .ZN(n5400) );
  INV_X1 U6828 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n9649) );
  NAND2_X1 U6829 ( .A1(n6530), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n5397) );
  NAND2_X1 U6830 ( .A1(n4935), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5396) );
  OAI211_X1 U6831 ( .C1(n4980), .C2(n9649), .A(n5397), .B(n5396), .ZN(n5398)
         );
  INV_X1 U6832 ( .A(n5398), .ZN(n5399) );
  NAND2_X1 U6833 ( .A1(n5400), .A2(n5399), .ZN(n9449) );
  INV_X1 U6834 ( .A(n5401), .ZN(n5402) );
  NOR2_X1 U6835 ( .A1(n5402), .A2(SI_21_), .ZN(n5403) );
  INV_X1 U6836 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n8076) );
  INV_X1 U6837 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n5405) );
  MUX2_X1 U6838 ( .A(n8076), .B(n5405), .S(n6447), .Z(n5407) );
  INV_X1 U6839 ( .A(SI_22_), .ZN(n5406) );
  NAND2_X1 U6840 ( .A1(n5407), .A2(n5406), .ZN(n5415) );
  INV_X1 U6841 ( .A(n5407), .ZN(n5408) );
  NAND2_X1 U6842 ( .A1(n5408), .A2(SI_22_), .ZN(n5409) );
  NAND2_X1 U6843 ( .A1(n5415), .A2(n5409), .ZN(n5416) );
  XNOR2_X1 U6844 ( .A(n5417), .B(n5416), .ZN(n7595) );
  NAND2_X1 U6845 ( .A1(n7595), .A2(n5114), .ZN(n5411) );
  NAND2_X1 U6846 ( .A1(n5465), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n5410) );
  OR2_X1 U6847 ( .A1(n9449), .A2(n9647), .ZN(n5412) );
  NAND2_X1 U6848 ( .A1(n9646), .A2(n5412), .ZN(n5414) );
  NAND2_X1 U6849 ( .A1(n9647), .A2(n9449), .ZN(n5413) );
  NAND2_X1 U6850 ( .A1(n5414), .A2(n5413), .ZN(n9632) );
  INV_X1 U6851 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n5419) );
  INV_X1 U6852 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n5418) );
  MUX2_X1 U6853 ( .A(n5419), .B(n5418), .S(n6447), .Z(n5421) );
  INV_X1 U6854 ( .A(SI_23_), .ZN(n5420) );
  NAND2_X1 U6855 ( .A1(n5421), .A2(n5420), .ZN(n5439) );
  INV_X1 U6856 ( .A(n5421), .ZN(n5422) );
  NAND2_X1 U6857 ( .A1(n5422), .A2(SI_23_), .ZN(n5423) );
  AND2_X1 U6858 ( .A1(n5439), .A2(n5423), .ZN(n5424) );
  OR2_X1 U6859 ( .A1(n5425), .A2(n5424), .ZN(n5426) );
  NAND2_X1 U6860 ( .A1(n5440), .A2(n5426), .ZN(n7644) );
  NAND2_X1 U6861 ( .A1(n7644), .A2(n5114), .ZN(n5428) );
  NAND2_X1 U6862 ( .A1(n5465), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n5427) );
  INV_X1 U6863 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n5430) );
  NAND2_X1 U6864 ( .A1(n5431), .A2(n5430), .ZN(n5432) );
  NAND2_X1 U6865 ( .A1(n5448), .A2(n5432), .ZN(n9639) );
  OR2_X1 U6866 ( .A1(n9639), .A2(n4984), .ZN(n5438) );
  INV_X1 U6867 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n5435) );
  NAND2_X1 U6868 ( .A1(n4935), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5434) );
  NAND2_X1 U6869 ( .A1(n4979), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n5433) );
  OAI211_X1 U6870 ( .C1(n5435), .C2(n4980), .A(n5434), .B(n5433), .ZN(n5436)
         );
  INV_X1 U6871 ( .A(n5436), .ZN(n5437) );
  NAND2_X1 U6872 ( .A1(n5438), .A2(n5437), .ZN(n9448) );
  INV_X1 U6873 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7763) );
  INV_X1 U6874 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n5441) );
  MUX2_X1 U6875 ( .A(n7763), .B(n5441), .S(n6447), .Z(n5443) );
  INV_X1 U6876 ( .A(SI_24_), .ZN(n5442) );
  NAND2_X1 U6877 ( .A1(n5443), .A2(n5442), .ZN(n5477) );
  INV_X1 U6878 ( .A(n5443), .ZN(n5444) );
  NAND2_X1 U6879 ( .A1(n5444), .A2(SI_24_), .ZN(n5445) );
  AND2_X1 U6880 ( .A1(n5477), .A2(n5445), .ZN(n5457) );
  NAND2_X1 U6881 ( .A1(n7761), .A2(n5114), .ZN(n5447) );
  NAND2_X1 U6882 ( .A1(n5465), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n5446) );
  INV_X1 U6883 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9152) );
  NAND2_X1 U6884 ( .A1(n5448), .A2(n9152), .ZN(n5449) );
  NAND2_X1 U6885 ( .A1(n5468), .A2(n5449), .ZN(n9150) );
  OR2_X1 U6886 ( .A1(n9150), .A2(n4984), .ZN(n5455) );
  INV_X1 U6887 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n5452) );
  NAND2_X1 U6888 ( .A1(n4979), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n5451) );
  NAND2_X1 U6889 ( .A1(n4935), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5450) );
  OAI211_X1 U6890 ( .C1(n5452), .C2(n4980), .A(n5451), .B(n5450), .ZN(n5453)
         );
  INV_X1 U6891 ( .A(n5453), .ZN(n5454) );
  NAND2_X1 U6892 ( .A1(n5455), .A2(n5454), .ZN(n9447) );
  NOR2_X1 U6893 ( .A1(n9624), .A2(n9447), .ZN(n5456) );
  NAND2_X1 U6894 ( .A1(n9624), .A2(n9447), .ZN(n9261) );
  NAND2_X1 U6895 ( .A1(n5481), .A2(n5477), .ZN(n5464) );
  INV_X1 U6896 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7815) );
  INV_X1 U6897 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n5459) );
  MUX2_X1 U6898 ( .A(n7815), .B(n5459), .S(n6447), .Z(n5461) );
  INV_X1 U6899 ( .A(SI_25_), .ZN(n5460) );
  NAND2_X1 U6900 ( .A1(n5461), .A2(n5460), .ZN(n5476) );
  INV_X1 U6901 ( .A(n5461), .ZN(n5462) );
  NAND2_X1 U6902 ( .A1(n5462), .A2(SI_25_), .ZN(n5478) );
  AND2_X1 U6903 ( .A1(n5476), .A2(n5478), .ZN(n5463) );
  NAND2_X1 U6904 ( .A1(n7798), .A2(n5114), .ZN(n5467) );
  NAND2_X1 U6905 ( .A1(n4997), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n5466) );
  INV_X1 U6906 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n9118) );
  NAND2_X1 U6907 ( .A1(n5468), .A2(n9118), .ZN(n5469) );
  AND2_X1 U6908 ( .A1(n5490), .A2(n5469), .ZN(n9612) );
  NAND2_X1 U6909 ( .A1(n9612), .A2(n5516), .ZN(n5475) );
  INV_X1 U6910 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n5472) );
  NAND2_X1 U6911 ( .A1(n6530), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n5471) );
  NAND2_X1 U6912 ( .A1(n4935), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n5470) );
  OAI211_X1 U6913 ( .C1(n5472), .C2(n4980), .A(n5471), .B(n5470), .ZN(n5473)
         );
  INV_X1 U6914 ( .A(n5473), .ZN(n5474) );
  NAND2_X1 U6915 ( .A1(n5475), .A2(n5474), .ZN(n9446) );
  AND2_X1 U6916 ( .A1(n5477), .A2(n5476), .ZN(n5480) );
  INV_X1 U6917 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7872) );
  INV_X1 U6918 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n5482) );
  MUX2_X1 U6919 ( .A(n7872), .B(n5482), .S(n6447), .Z(n5484) );
  INV_X1 U6920 ( .A(SI_26_), .ZN(n5483) );
  NAND2_X1 U6921 ( .A1(n5484), .A2(n5483), .ZN(n5503) );
  INV_X1 U6922 ( .A(n5484), .ZN(n5485) );
  NAND2_X1 U6923 ( .A1(n5485), .A2(SI_26_), .ZN(n5486) );
  AND2_X1 U6924 ( .A1(n5503), .A2(n5486), .ZN(n5501) );
  NAND2_X1 U6925 ( .A1(n7830), .A2(n5114), .ZN(n5488) );
  NAND2_X1 U6926 ( .A1(n4997), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n5487) );
  INV_X1 U6927 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n6432) );
  NAND2_X1 U6928 ( .A1(n5490), .A2(n6432), .ZN(n5491) );
  NAND2_X1 U6929 ( .A1(n5528), .A2(n5491), .ZN(n9598) );
  OR2_X1 U6930 ( .A1(n9598), .A2(n4984), .ZN(n5497) );
  INV_X1 U6931 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n8085) );
  NAND2_X1 U6932 ( .A1(n5492), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n5494) );
  NAND2_X1 U6933 ( .A1(n6530), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n5493) );
  OAI211_X1 U6934 ( .C1(n4982), .C2(n8085), .A(n5494), .B(n5493), .ZN(n5495)
         );
  INV_X1 U6935 ( .A(n5495), .ZN(n5496) );
  NAND2_X1 U6936 ( .A1(n5497), .A2(n5496), .ZN(n9445) );
  NAND2_X1 U6937 ( .A1(n5498), .A2(n4910), .ZN(n5500) );
  NAND2_X1 U6938 ( .A1(n9812), .A2(n9445), .ZN(n5499) );
  INV_X1 U6939 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n5506) );
  INV_X1 U6940 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n5505) );
  MUX2_X1 U6941 ( .A(n5506), .B(n5505), .S(n6447), .Z(n5508) );
  INV_X1 U6942 ( .A(SI_27_), .ZN(n5507) );
  NAND2_X1 U6943 ( .A1(n5508), .A2(n5507), .ZN(n5523) );
  INV_X1 U6944 ( .A(n5508), .ZN(n5509) );
  NAND2_X1 U6945 ( .A1(n5509), .A2(SI_27_), .ZN(n5510) );
  AND2_X1 U6946 ( .A1(n5523), .A2(n5510), .ZN(n5511) );
  OR2_X1 U6947 ( .A1(n5512), .A2(n5511), .ZN(n5513) );
  NAND2_X1 U6948 ( .A1(n5524), .A2(n5513), .ZN(n7921) );
  NAND2_X1 U6949 ( .A1(n7921), .A2(n5114), .ZN(n5515) );
  NAND2_X1 U6950 ( .A1(n5465), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n5514) );
  XNOR2_X1 U6951 ( .A(n5528), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n9584) );
  NAND2_X1 U6952 ( .A1(n9584), .A2(n5516), .ZN(n5522) );
  INV_X1 U6953 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n5519) );
  NAND2_X1 U6954 ( .A1(n6530), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n5518) );
  NAND2_X1 U6955 ( .A1(n4935), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n5517) );
  OAI211_X1 U6956 ( .C1(n5519), .C2(n4980), .A(n5518), .B(n5517), .ZN(n5520)
         );
  INV_X1 U6957 ( .A(n5520), .ZN(n5521) );
  NAND2_X1 U6958 ( .A1(n5522), .A2(n5521), .ZN(n9444) );
  INV_X1 U6959 ( .A(n9444), .ZN(n6431) );
  NAND2_X1 U6960 ( .A1(n9583), .A2(n6431), .ZN(n9315) );
  MUX2_X1 U6961 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n6447), .Z(n5642) );
  INV_X1 U6962 ( .A(SI_28_), .ZN(n5643) );
  XNOR2_X1 U6963 ( .A(n5642), .B(n5643), .ZN(n5640) );
  NAND2_X1 U6964 ( .A1(n5465), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n5525) );
  INV_X1 U6965 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n5527) );
  INV_X1 U6966 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n5906) );
  OAI21_X1 U6967 ( .B1(n5528), .B2(n5527), .A(n5906), .ZN(n5529) );
  NAND2_X1 U6968 ( .A1(n5529), .A2(n8162), .ZN(n9566) );
  OR2_X1 U6969 ( .A1(n9566), .A2(n4984), .ZN(n5534) );
  INV_X1 U6970 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n9565) );
  NAND2_X1 U6971 ( .A1(n6530), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n5531) );
  NAND2_X1 U6972 ( .A1(n4935), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5530) );
  OAI211_X1 U6973 ( .C1(n9565), .C2(n4980), .A(n5531), .B(n5530), .ZN(n5532)
         );
  INV_X1 U6974 ( .A(n5532), .ZN(n5533) );
  NAND2_X1 U6975 ( .A1(n5534), .A2(n5533), .ZN(n9443) );
  INV_X1 U6976 ( .A(n9443), .ZN(n9272) );
  NAND2_X1 U6977 ( .A1(n9568), .A2(n9272), .ZN(n9316) );
  NAND2_X1 U6978 ( .A1(n5535), .A2(n9407), .ZN(n5536) );
  NOR2_X1 U6979 ( .A1(n5538), .A2(P1_IR_REG_19__SCAN_IN), .ZN(n5539) );
  NAND2_X1 U6980 ( .A1(n5540), .A2(n5539), .ZN(n5545) );
  INV_X1 U6981 ( .A(n5545), .ZN(n5541) );
  NAND2_X1 U6982 ( .A1(n5541), .A2(n5546), .ZN(n5604) );
  INV_X1 U6983 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5601) );
  NAND2_X1 U6984 ( .A1(n5548), .A2(n5601), .ZN(n5542) );
  NAND2_X1 U6985 ( .A1(n5542), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5543) );
  OR2_X1 U6986 ( .A1(n5543), .A2(n5602), .ZN(n5544) );
  NAND2_X1 U6987 ( .A1(n5543), .A2(n5602), .ZN(n5593) );
  NAND2_X1 U6988 ( .A1(n5545), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5547) );
  NAND2_X1 U6989 ( .A1(n9376), .A2(n9298), .ZN(n9373) );
  AND2_X1 U6990 ( .A1(n5675), .A2(n9373), .ZN(n5549) );
  NAND2_X1 U6991 ( .A1(n9296), .A2(n5670), .ZN(n9432) );
  AND2_X1 U6992 ( .A1(n5677), .A2(n9295), .ZN(n5630) );
  INV_X1 U6993 ( .A(n5630), .ZN(n6625) );
  OAI21_X1 U6994 ( .B1(n9432), .B2(n9373), .A(n6625), .ZN(n7185) );
  OR2_X1 U6995 ( .A1(n5549), .A2(n7185), .ZN(n7434) );
  AND2_X1 U6996 ( .A1(n5677), .A2(n9549), .ZN(n9278) );
  NAND2_X1 U6997 ( .A1(n9278), .A2(n9298), .ZN(n10041) );
  NAND2_X1 U6998 ( .A1(n7434), .A2(n10041), .ZN(n10029) );
  INV_X1 U6999 ( .A(n10029), .ZN(n9995) );
  INV_X1 U7000 ( .A(n6695), .ZN(n5550) );
  INV_X1 U7001 ( .A(n7037), .ZN(n5551) );
  NAND2_X1 U7002 ( .A1(n7040), .A2(n5552), .ZN(n6975) );
  INV_X1 U7003 ( .A(n5553), .ZN(n9380) );
  NAND2_X1 U7004 ( .A1(n6874), .A2(n6982), .ZN(n5554) );
  NAND2_X1 U7005 ( .A1(n9467), .A2(n9976), .ZN(n9331) );
  NAND2_X1 U7006 ( .A1(n7298), .A2(n9331), .ZN(n5557) );
  NAND2_X1 U7007 ( .A1(n5555), .A2(n7302), .ZN(n5556) );
  INV_X1 U7008 ( .A(n5558), .ZN(n5559) );
  NAND2_X1 U7009 ( .A1(n7179), .A2(n5565), .ZN(n5561) );
  NAND2_X1 U7010 ( .A1(n9954), .A2(n5563), .ZN(n7364) );
  AND2_X1 U7011 ( .A1(n9205), .A2(n7364), .ZN(n9388) );
  NAND3_X1 U7012 ( .A1(n7358), .A2(n9388), .A3(n9208), .ZN(n5567) );
  INV_X1 U7013 ( .A(n9388), .ZN(n7361) );
  NAND3_X1 U7014 ( .A1(n9214), .A2(n7415), .A3(n7361), .ZN(n5562) );
  NAND2_X1 U7015 ( .A1(n5562), .A2(n9208), .ZN(n9343) );
  OR2_X1 U7016 ( .A1(n9954), .A2(n5563), .ZN(n5564) );
  AND2_X1 U7017 ( .A1(n7415), .A2(n5564), .ZN(n9389) );
  OR2_X1 U7018 ( .A1(n5565), .A2(n7179), .ZN(n7359) );
  AND3_X1 U7019 ( .A1(n9214), .A2(n9389), .A3(n7359), .ZN(n5566) );
  NAND2_X1 U7020 ( .A1(n5567), .A2(n9341), .ZN(n7328) );
  INV_X1 U7021 ( .A(n9459), .ZN(n5568) );
  NAND2_X1 U7022 ( .A1(n7802), .A2(n5568), .ZN(n9220) );
  AND2_X1 U7023 ( .A1(n9220), .A2(n9215), .ZN(n9346) );
  OR2_X1 U7024 ( .A1(n7802), .A2(n5568), .ZN(n9218) );
  NAND2_X1 U7025 ( .A1(n7547), .A2(n9394), .ZN(n7546) );
  NAND2_X1 U7026 ( .A1(n7546), .A2(n9223), .ZN(n7635) );
  INV_X1 U7027 ( .A(n7635), .ZN(n5571) );
  INV_X1 U7028 ( .A(n9396), .ZN(n5570) );
  AOI21_X2 U7029 ( .B1(n5571), .B2(n5570), .A(n5569), .ZN(n7691) );
  INV_X1 U7030 ( .A(n9456), .ZN(n7637) );
  OR2_X1 U7031 ( .A1(n9076), .A2(n7637), .ZN(n9351) );
  NAND2_X1 U7032 ( .A1(n9076), .A2(n7637), .ZN(n9226) );
  OR2_X1 U7033 ( .A1(n7773), .A2(n5572), .ZN(n9229) );
  NAND2_X1 U7034 ( .A1(n7773), .A2(n5572), .ZN(n9227) );
  NAND2_X1 U7035 ( .A1(n9229), .A2(n9227), .ZN(n7766) );
  INV_X1 U7036 ( .A(n9453), .ZN(n5573) );
  OR2_X1 U7037 ( .A1(n7946), .A2(n5573), .ZN(n9362) );
  NAND2_X1 U7038 ( .A1(n7946), .A2(n5573), .ZN(n9238) );
  NAND2_X1 U7039 ( .A1(n7941), .A2(n9402), .ZN(n7940) );
  NAND2_X1 U7040 ( .A1(n7940), .A2(n9362), .ZN(n9706) );
  INV_X1 U7041 ( .A(n9452), .ZN(n5574) );
  OR2_X1 U7042 ( .A1(n9793), .A2(n5574), .ZN(n9240) );
  NAND2_X1 U7043 ( .A1(n9793), .A2(n5574), .ZN(n9241) );
  NAND2_X1 U7044 ( .A1(n9240), .A2(n9241), .ZN(n9703) );
  INV_X1 U7045 ( .A(n9451), .ZN(n5576) );
  OR2_X1 U7046 ( .A1(n9787), .A2(n5576), .ZN(n9239) );
  NAND2_X1 U7047 ( .A1(n9787), .A2(n5576), .ZN(n9363) );
  INV_X1 U7048 ( .A(n9449), .ZN(n9085) );
  OR2_X1 U7049 ( .A1(n9647), .A2(n9085), .ZN(n9253) );
  NAND2_X1 U7050 ( .A1(n9647), .A2(n9085), .ZN(n9251) );
  NAND2_X1 U7051 ( .A1(n9652), .A2(n9653), .ZN(n5578) );
  XNOR2_X1 U7052 ( .A(n9824), .B(n9448), .ZN(n9633) );
  NAND2_X1 U7053 ( .A1(n9634), .A2(n9633), .ZN(n5579) );
  INV_X1 U7054 ( .A(n9448), .ZN(n9252) );
  NAND2_X1 U7055 ( .A1(n9824), .A2(n9252), .ZN(n9300) );
  INV_X1 U7056 ( .A(n9447), .ZN(n9086) );
  NAND2_X1 U7057 ( .A1(n9624), .A2(n9086), .ZN(n9309) );
  NAND2_X1 U7058 ( .A1(n9301), .A2(n9309), .ZN(n9619) );
  INV_X1 U7059 ( .A(n9446), .ZN(n6430) );
  NOR2_X1 U7060 ( .A1(n9611), .A2(n6430), .ZN(n9378) );
  NAND2_X1 U7061 ( .A1(n9611), .A2(n6430), .ZN(n9310) );
  XNOR2_X1 U7062 ( .A(n9812), .B(n9445), .ZN(n9594) );
  NAND2_X1 U7063 ( .A1(n9590), .A2(n9594), .ZN(n5581) );
  INV_X1 U7064 ( .A(n9445), .ZN(n9262) );
  NAND2_X1 U7065 ( .A1(n9812), .A2(n9262), .ZN(n9317) );
  NAND2_X1 U7066 ( .A1(n5581), .A2(n9317), .ZN(n9576) );
  NAND2_X1 U7067 ( .A1(n9576), .A2(n9580), .ZN(n9575) );
  XNOR2_X1 U7068 ( .A(n5639), .B(n9407), .ZN(n5588) );
  OR2_X1 U7069 ( .A1(n9295), .A2(n9298), .ZN(n9286) );
  OAI21_X2 U7070 ( .B1(n5677), .B2(n9376), .A(n9286), .ZN(n9698) );
  INV_X1 U7071 ( .A(n9432), .ZN(n6504) );
  INV_X1 U7072 ( .A(n9878), .ZN(n9899) );
  INV_X1 U7073 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n8161) );
  NAND2_X1 U7074 ( .A1(n6530), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n5584) );
  INV_X1 U7075 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n5582) );
  OR2_X1 U7076 ( .A1(n4982), .A2(n5582), .ZN(n5583) );
  OAI211_X1 U7077 ( .C1(n8161), .C2(n4980), .A(n5584), .B(n5583), .ZN(n5585)
         );
  INV_X1 U7078 ( .A(n5585), .ZN(n5586) );
  OAI21_X1 U7079 ( .B1(n8162), .B2(n4984), .A(n5586), .ZN(n9442) );
  AND2_X1 U7080 ( .A1(n6504), .A2(n9878), .ZN(n9169) );
  INV_X1 U7081 ( .A(n9169), .ZN(n9096) );
  INV_X1 U7082 ( .A(n9096), .ZN(n9181) );
  AOI22_X1 U7083 ( .A1(n9444), .A2(n9291), .B1(n9442), .B2(n9181), .ZN(n5900)
         );
  INV_X1 U7084 ( .A(n5900), .ZN(n5587) );
  AOI21_X2 U7085 ( .B1(n5588), .B2(n9698), .A(n5587), .ZN(n9574) );
  INV_X1 U7086 ( .A(n9812), .ZN(n9596) );
  INV_X1 U7087 ( .A(n9824), .ZN(n9638) );
  NAND2_X1 U7088 ( .A1(n7045), .A2(n9336), .ZN(n7303) );
  OR2_X1 U7089 ( .A1(n7303), .A2(n7302), .ZN(n7318) );
  INV_X1 U7090 ( .A(n7179), .ZN(n10001) );
  NOR2_X1 U7091 ( .A1(n7422), .A2(n10017), .ZN(n7421) );
  INV_X1 U7092 ( .A(n7338), .ZN(n10026) );
  NAND2_X1 U7093 ( .A1(n7421), .A2(n10026), .ZN(n7444) );
  INV_X1 U7094 ( .A(n9729), .ZN(n7902) );
  INV_X1 U7095 ( .A(n9076), .ZN(n10040) );
  INV_X1 U7096 ( .A(n9957), .ZN(n9977) );
  AOI21_X1 U7097 ( .B1(n9568), .B2(n9582), .A(n9977), .ZN(n5591) );
  NAND2_X1 U7098 ( .A1(n5591), .A2(n4366), .ZN(n9570) );
  OAI21_X1 U7099 ( .B1(n9564), .B2(n9995), .A(n5592), .ZN(n5634) );
  NAND2_X1 U7100 ( .A1(n5593), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5594) );
  XNOR2_X1 U7101 ( .A(n5594), .B(n5600), .ZN(n7645) );
  XNOR2_X1 U7102 ( .A(n5595), .B(P1_IR_REG_26__SCAN_IN), .ZN(n7831) );
  INV_X1 U7103 ( .A(n7831), .ZN(n5599) );
  NAND2_X1 U7104 ( .A1(n5596), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5598) );
  INV_X1 U7105 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5597) );
  XNOR2_X1 U7106 ( .A(n5598), .B(n5597), .ZN(n7799) );
  NAND3_X1 U7107 ( .A1(n5602), .A2(n5601), .A3(n5600), .ZN(n5603) );
  INV_X1 U7108 ( .A(n5904), .ZN(n5607) );
  NAND2_X1 U7109 ( .A1(n7799), .A2(P1_B_REG_SCAN_IN), .ZN(n5609) );
  MUX2_X1 U7110 ( .A(n5609), .B(P1_B_REG_SCAN_IN), .S(n5608), .Z(n5610) );
  NAND2_X1 U7111 ( .A1(n5610), .A2(n7831), .ZN(n5891) );
  INV_X1 U7112 ( .A(n5891), .ZN(n5611) );
  OR2_X2 U7113 ( .A1(n9292), .A2(n5611), .ZN(n9966) );
  NOR2_X1 U7114 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_2__SCAN_IN), .ZN(
        n5615) );
  NOR4_X1 U7115 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_3__SCAN_IN), .A4(P1_D_REG_4__SCAN_IN), .ZN(n5614) );
  NOR4_X1 U7116 ( .A1(P1_D_REG_9__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_11__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n5613) );
  NOR4_X1 U7117 ( .A1(P1_D_REG_5__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_7__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n5612) );
  NAND4_X1 U7118 ( .A1(n5615), .A2(n5614), .A3(n5613), .A4(n5612), .ZN(n5621)
         );
  NOR4_X1 U7119 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .A3(
        P1_D_REG_19__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n5619) );
  NOR4_X1 U7120 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_13__SCAN_IN), .A3(
        P1_D_REG_14__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n5618) );
  NOR4_X1 U7121 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5617) );
  NOR4_X1 U7122 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_23__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n5616) );
  NAND4_X1 U7123 ( .A1(n5619), .A2(n5618), .A3(n5617), .A4(n5616), .ZN(n5620)
         );
  NOR2_X1 U7124 ( .A1(n5621), .A2(n5620), .ZN(n5892) );
  INV_X1 U7125 ( .A(n5892), .ZN(n5622) );
  OR2_X1 U7126 ( .A1(n9292), .A2(n5622), .ZN(n5623) );
  INV_X1 U7127 ( .A(n9373), .ZN(n9290) );
  NOR2_X1 U7128 ( .A1(n9432), .A2(n9290), .ZN(n5901) );
  AOI21_X1 U7129 ( .B1(n9966), .B2(n5623), .A(n5901), .ZN(n7033) );
  OR2_X1 U7130 ( .A1(n5891), .A2(P1_D_REG_1__SCAN_IN), .ZN(n5624) );
  NAND2_X1 U7131 ( .A1(n5599), .A2(n7799), .ZN(n9841) );
  NAND2_X1 U7132 ( .A1(n9957), .A2(n9549), .ZN(n5902) );
  INV_X1 U7133 ( .A(n5902), .ZN(n5625) );
  NOR2_X1 U7134 ( .A1(n7032), .A2(n5625), .ZN(n5626) );
  AND2_X1 U7135 ( .A1(n7033), .A2(n5626), .ZN(n5633) );
  OR2_X1 U7136 ( .A1(n5891), .A2(P1_D_REG_0__SCAN_IN), .ZN(n5628) );
  INV_X1 U7137 ( .A(n5608), .ZN(n5627) );
  NAND2_X1 U7138 ( .A1(n5627), .A2(n5599), .ZN(n9842) );
  AND2_X2 U7139 ( .A1(n5633), .A2(n5890), .ZN(n10068) );
  MUX2_X1 U7140 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n5634), .S(n10068), .Z(n5629) );
  INV_X1 U7141 ( .A(n5629), .ZN(n5632) );
  AND2_X1 U7142 ( .A1(n5630), .A2(n9373), .ZN(n9993) );
  NAND2_X1 U7143 ( .A1(n5632), .A2(n5631), .ZN(P1_U3550) );
  INV_X1 U7144 ( .A(n5890), .ZN(n7031) );
  AND2_X2 U7145 ( .A1(n5633), .A2(n7031), .ZN(n10049) );
  MUX2_X1 U7146 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n5634), .S(n10049), .Z(n5635) );
  INV_X1 U7147 ( .A(n5635), .ZN(n5637) );
  NAND2_X1 U7148 ( .A1(n5637), .A2(n5636), .ZN(P1_U3518) );
  INV_X1 U7149 ( .A(n9316), .ZN(n5638) );
  AOI21_X1 U7150 ( .B1(n5639), .B2(n9407), .A(n5638), .ZN(n5649) );
  INV_X1 U7151 ( .A(n5642), .ZN(n5644) );
  INV_X1 U7152 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n5645) );
  INV_X1 U7153 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8187) );
  MUX2_X1 U7154 ( .A(n5645), .B(n8187), .S(n8358), .Z(n8171) );
  NAND2_X1 U7155 ( .A1(n8185), .A2(n5114), .ZN(n5647) );
  NAND2_X1 U7156 ( .A1(n4997), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n5646) );
  INV_X1 U7157 ( .A(n9442), .ZN(n5648) );
  NAND2_X1 U7158 ( .A1(n8164), .A2(n5648), .ZN(n9366) );
  XNOR2_X1 U7159 ( .A(n5649), .B(n9277), .ZN(n5659) );
  NAND2_X1 U7160 ( .A1(n4979), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n5653) );
  INV_X1 U7161 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n9559) );
  OR2_X1 U7162 ( .A1(n4980), .A2(n9559), .ZN(n5652) );
  INV_X1 U7163 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n5650) );
  OR2_X1 U7164 ( .A1(n4982), .A2(n5650), .ZN(n5651) );
  AND3_X1 U7165 ( .A1(n5653), .A2(n5652), .A3(n5651), .ZN(n9368) );
  INV_X1 U7166 ( .A(P1_B_REG_SCAN_IN), .ZN(n5655) );
  OR2_X1 U7167 ( .A1(n5654), .A2(n5655), .ZN(n5656) );
  NAND2_X1 U7168 ( .A1(n9181), .A2(n5656), .ZN(n8197) );
  NAND2_X1 U7169 ( .A1(n9443), .A2(n9291), .ZN(n5657) );
  OAI21_X1 U7170 ( .B1(n9368), .B2(n8197), .A(n5657), .ZN(n5658) );
  AOI21_X1 U7171 ( .B1(n8164), .B2(n4366), .A(n9977), .ZN(n5660) );
  NAND2_X1 U7172 ( .A1(n5660), .A2(n8194), .ZN(n8166) );
  NAND2_X1 U7173 ( .A1(n8168), .A2(n10029), .ZN(n5663) );
  NAND2_X1 U7174 ( .A1(n5664), .A2(n5663), .ZN(n5667) );
  NAND2_X1 U7175 ( .A1(n5667), .A2(n10049), .ZN(n5666) );
  NAND2_X1 U7176 ( .A1(n10047), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n5665) );
  NAND2_X1 U7177 ( .A1(n5667), .A2(n10068), .ZN(n5669) );
  NAND2_X1 U7178 ( .A1(n10066), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n5668) );
  NAND2_X1 U7179 ( .A1(n4908), .A2(n4906), .ZN(P1_U3551) );
  AND2_X2 U7180 ( .A1(n6439), .A2(n5671), .ZN(n5703) );
  NAND2_X1 U7181 ( .A1(n5674), .A2(n5673), .ZN(n5676) );
  INV_X1 U7182 ( .A(n5684), .ZN(n5681) );
  NAND2_X1 U7183 ( .A1(n9290), .A2(n5677), .ZN(n5678) );
  OR2_X1 U7184 ( .A1(n5671), .A2(n9376), .ZN(n7191) );
  AND3_X2 U7185 ( .A1(n5678), .A2(n7191), .A3(n6439), .ZN(n5707) );
  NAND2_X1 U7186 ( .A1(n5780), .A2(n5672), .ZN(n5679) );
  NAND2_X1 U7187 ( .A1(n5680), .A2(n5679), .ZN(n5682) );
  NAND2_X1 U7188 ( .A1(n5681), .A2(n5682), .ZN(n5685) );
  INV_X1 U7189 ( .A(n5682), .ZN(n5683) );
  NAND2_X1 U7190 ( .A1(n5684), .A2(n5683), .ZN(n5693) );
  NAND2_X1 U7191 ( .A1(n5685), .A2(n5693), .ZN(n6691) );
  NAND2_X1 U7192 ( .A1(n5689), .A2(n4905), .ZN(n6615) );
  NAND2_X1 U7193 ( .A1(n6695), .A2(n5707), .ZN(n5688) );
  INV_X1 U7194 ( .A(n6439), .ZN(n6502) );
  AOI22_X1 U7195 ( .A1(n5780), .A2(n7182), .B1(P1_IR_REG_0__SCAN_IN), .B2(
        n6502), .ZN(n5687) );
  NAND2_X1 U7196 ( .A1(n5688), .A2(n5687), .ZN(n6616) );
  NAND2_X1 U7197 ( .A1(n6615), .A2(n6616), .ZN(n5691) );
  NAND2_X1 U7198 ( .A1(n5689), .A2(n5874), .ZN(n5690) );
  NAND2_X1 U7199 ( .A1(n5691), .A2(n5690), .ZN(n6694) );
  INV_X1 U7200 ( .A(n6694), .ZN(n5692) );
  NAND2_X1 U7201 ( .A1(n5703), .A2(n6982), .ZN(n5695) );
  NAND2_X1 U7202 ( .A1(n9468), .A2(n5780), .ZN(n5694) );
  NAND2_X1 U7203 ( .A1(n5695), .A2(n5694), .ZN(n5696) );
  XNOR2_X1 U7204 ( .A(n5696), .B(n5874), .ZN(n5697) );
  AOI22_X1 U7205 ( .A1(n9468), .A2(n5707), .B1(n5780), .B2(n6982), .ZN(n5698)
         );
  NAND2_X1 U7206 ( .A1(n5697), .A2(n5698), .ZN(n5702) );
  INV_X1 U7207 ( .A(n5697), .ZN(n5700) );
  INV_X1 U7208 ( .A(n5698), .ZN(n5699) );
  NAND2_X1 U7209 ( .A1(n5700), .A2(n5699), .ZN(n5701) );
  AND2_X1 U7210 ( .A1(n5702), .A2(n5701), .ZN(n6835) );
  NAND2_X1 U7211 ( .A1(n6833), .A2(n5702), .ZN(n6871) );
  NAND2_X1 U7212 ( .A1(n9467), .A2(n5780), .ZN(n5705) );
  NAND2_X1 U7213 ( .A1(n5703), .A2(n7302), .ZN(n5704) );
  NAND2_X1 U7214 ( .A1(n5705), .A2(n5704), .ZN(n5706) );
  XNOR2_X1 U7215 ( .A(n5706), .B(n5886), .ZN(n5708) );
  AOI22_X1 U7216 ( .A1(n9467), .A2(n5707), .B1(n5780), .B2(n7302), .ZN(n5709)
         );
  XNOR2_X1 U7217 ( .A(n5708), .B(n5709), .ZN(n6872) );
  INV_X1 U7218 ( .A(n5708), .ZN(n5710) );
  NAND2_X1 U7219 ( .A1(n5710), .A2(n5709), .ZN(n5711) );
  NAND2_X1 U7220 ( .A1(n9466), .A2(n5780), .ZN(n5713) );
  NAND2_X1 U7221 ( .A1(n5703), .A2(n7317), .ZN(n5712) );
  NAND2_X1 U7222 ( .A1(n5713), .A2(n5712), .ZN(n5714) );
  AOI22_X1 U7223 ( .A1(n9466), .A2(n5707), .B1(n5780), .B2(n7317), .ZN(n5717)
         );
  XNOR2_X1 U7224 ( .A(n5716), .B(n5717), .ZN(n6922) );
  INV_X1 U7225 ( .A(n6922), .ZN(n5715) );
  INV_X1 U7226 ( .A(n5716), .ZN(n5719) );
  INV_X1 U7227 ( .A(n5717), .ZN(n5718) );
  NAND2_X1 U7228 ( .A1(n5719), .A2(n5718), .ZN(n5720) );
  NAND2_X1 U7229 ( .A1(n6924), .A2(n5720), .ZN(n7161) );
  NAND2_X1 U7230 ( .A1(n9465), .A2(n5780), .ZN(n5722) );
  NAND2_X1 U7231 ( .A1(n9992), .A2(n5703), .ZN(n5721) );
  NAND2_X1 U7232 ( .A1(n5722), .A2(n5721), .ZN(n5723) );
  XNOR2_X1 U7233 ( .A(n5723), .B(n5886), .ZN(n7162) );
  NAND2_X1 U7234 ( .A1(n9465), .A2(n5707), .ZN(n5726) );
  NAND2_X1 U7235 ( .A1(n9992), .A2(n5853), .ZN(n5725) );
  NAND2_X1 U7236 ( .A1(n5726), .A2(n5725), .ZN(n7167) );
  NAND2_X1 U7237 ( .A1(n7179), .A2(n5703), .ZN(n5728) );
  NAND2_X1 U7238 ( .A1(n9464), .A2(n5780), .ZN(n5727) );
  NAND2_X1 U7239 ( .A1(n5728), .A2(n5727), .ZN(n5729) );
  XNOR2_X1 U7240 ( .A(n5729), .B(n5874), .ZN(n5731) );
  AOI22_X1 U7241 ( .A1(n7179), .A2(n5853), .B1(n5707), .B2(n9464), .ZN(n5730)
         );
  NAND2_X1 U7242 ( .A1(n5731), .A2(n5730), .ZN(n7239) );
  OAI21_X1 U7243 ( .B1(n5731), .B2(n5730), .A(n7239), .ZN(n5732) );
  INV_X1 U7244 ( .A(n5732), .ZN(n7226) );
  NAND2_X1 U7245 ( .A1(n9954), .A2(n5703), .ZN(n5736) );
  NAND2_X1 U7246 ( .A1(n9463), .A2(n5780), .ZN(n5735) );
  NAND2_X1 U7247 ( .A1(n5736), .A2(n5735), .ZN(n5737) );
  XNOR2_X1 U7248 ( .A(n5737), .B(n5874), .ZN(n5739) );
  AND2_X1 U7249 ( .A1(n9463), .A2(n5707), .ZN(n5738) );
  AOI21_X1 U7250 ( .B1(n9954), .B2(n5853), .A(n5738), .ZN(n5740) );
  NAND2_X1 U7251 ( .A1(n5739), .A2(n5740), .ZN(n5744) );
  INV_X1 U7252 ( .A(n5739), .ZN(n5742) );
  INV_X1 U7253 ( .A(n5740), .ZN(n5741) );
  NAND2_X1 U7254 ( .A1(n5742), .A2(n5741), .ZN(n5743) );
  NAND2_X1 U7255 ( .A1(n5744), .A2(n5743), .ZN(n7238) );
  AOI22_X1 U7256 ( .A1(n7495), .A2(n5703), .B1(n5780), .B2(n9462), .ZN(n5745)
         );
  XOR2_X1 U7257 ( .A(n5886), .B(n5745), .Z(n5746) );
  AOI22_X1 U7258 ( .A1(n7495), .A2(n5853), .B1(n5707), .B2(n9462), .ZN(n7489)
         );
  OAI21_X1 U7259 ( .B1(n7486), .B2(n7489), .A(n7487), .ZN(n7536) );
  NAND2_X1 U7260 ( .A1(n10017), .A2(n5703), .ZN(n5748) );
  NAND2_X1 U7261 ( .A1(n9461), .A2(n5780), .ZN(n5747) );
  NAND2_X1 U7262 ( .A1(n5748), .A2(n5747), .ZN(n5749) );
  XNOR2_X1 U7263 ( .A(n5749), .B(n5874), .ZN(n5752) );
  AND2_X1 U7264 ( .A1(n9461), .A2(n5707), .ZN(n5750) );
  AOI21_X1 U7265 ( .B1(n10017), .B2(n5853), .A(n5750), .ZN(n5751) );
  NAND2_X1 U7266 ( .A1(n5752), .A2(n5751), .ZN(n5753) );
  OAI21_X1 U7267 ( .B1(n5752), .B2(n5751), .A(n5753), .ZN(n7537) );
  INV_X1 U7268 ( .A(n5753), .ZN(n5754) );
  AOI22_X1 U7269 ( .A1(n7338), .A2(n5703), .B1(n5780), .B2(n9460), .ZN(n5755)
         );
  AOI22_X1 U7270 ( .A1(n7338), .A2(n5853), .B1(n5707), .B2(n9460), .ZN(n9857)
         );
  NAND2_X1 U7271 ( .A1(n9856), .A2(n9857), .ZN(n9855) );
  INV_X1 U7272 ( .A(n5756), .ZN(n5757) );
  NAND2_X1 U7273 ( .A1(n9855), .A2(n5757), .ZN(n7803) );
  NAND2_X1 U7274 ( .A1(n7802), .A2(n5703), .ZN(n5759) );
  NAND2_X1 U7275 ( .A1(n9459), .A2(n5853), .ZN(n5758) );
  NAND2_X1 U7276 ( .A1(n5759), .A2(n5758), .ZN(n5760) );
  XNOR2_X1 U7277 ( .A(n5760), .B(n5886), .ZN(n5765) );
  AOI22_X1 U7278 ( .A1(n7802), .A2(n5853), .B1(n5707), .B2(n9459), .ZN(n5766)
         );
  XNOR2_X1 U7279 ( .A(n5765), .B(n5766), .ZN(n7806) );
  NAND2_X1 U7280 ( .A1(n7803), .A2(n7806), .ZN(n7804) );
  NAND2_X1 U7281 ( .A1(n7979), .A2(n5703), .ZN(n5762) );
  NAND2_X1 U7282 ( .A1(n9458), .A2(n5853), .ZN(n5761) );
  NAND2_X1 U7283 ( .A1(n5762), .A2(n5761), .ZN(n5763) );
  XNOR2_X1 U7284 ( .A(n5763), .B(n5886), .ZN(n5775) );
  AND2_X1 U7285 ( .A1(n9458), .A2(n5707), .ZN(n5764) );
  AOI21_X1 U7286 ( .B1(n7979), .B2(n5853), .A(n5764), .ZN(n5773) );
  XNOR2_X1 U7287 ( .A(n5775), .B(n5773), .ZN(n7973) );
  INV_X1 U7288 ( .A(n5765), .ZN(n5767) );
  NAND2_X1 U7289 ( .A1(n5767), .A2(n5766), .ZN(n7974) );
  NAND2_X1 U7290 ( .A1(n9729), .A2(n5703), .ZN(n5770) );
  NAND2_X1 U7291 ( .A1(n9457), .A2(n5853), .ZN(n5769) );
  NAND2_X1 U7292 ( .A1(n5770), .A2(n5769), .ZN(n5771) );
  XNOR2_X1 U7293 ( .A(n5771), .B(n5886), .ZN(n5779) );
  AND2_X1 U7294 ( .A1(n9457), .A2(n5707), .ZN(n5772) );
  AOI21_X1 U7295 ( .B1(n9729), .B2(n5853), .A(n5772), .ZN(n5777) );
  XNOR2_X1 U7296 ( .A(n5779), .B(n5777), .ZN(n7894) );
  INV_X1 U7297 ( .A(n5773), .ZN(n5774) );
  NAND2_X1 U7298 ( .A1(n5775), .A2(n5774), .ZN(n7895) );
  INV_X1 U7299 ( .A(n5777), .ZN(n5778) );
  AOI22_X1 U7300 ( .A1(n9076), .A2(n5703), .B1(n5780), .B2(n9456), .ZN(n5781)
         );
  OAI22_X1 U7301 ( .A1(n10040), .A2(n5724), .B1(n7637), .B2(n5782), .ZN(n9070)
         );
  AOI22_X1 U7302 ( .A1(n7773), .A2(n5703), .B1(n5780), .B2(n9455), .ZN(n5783)
         );
  XNOR2_X1 U7303 ( .A(n5783), .B(n5886), .ZN(n5784) );
  AOI22_X1 U7304 ( .A1(n7773), .A2(n5853), .B1(n5707), .B2(n9455), .ZN(n9191)
         );
  NAND2_X1 U7305 ( .A1(n7890), .A2(n5703), .ZN(n5790) );
  NAND2_X1 U7306 ( .A1(n9454), .A2(n5780), .ZN(n5789) );
  NAND2_X1 U7307 ( .A1(n5790), .A2(n5789), .ZN(n5791) );
  XNOR2_X1 U7308 ( .A(n5791), .B(n5886), .ZN(n5795) );
  NAND2_X1 U7309 ( .A1(n7890), .A2(n5853), .ZN(n5793) );
  NAND2_X1 U7310 ( .A1(n9454), .A2(n5707), .ZN(n5792) );
  NAND2_X1 U7311 ( .A1(n5793), .A2(n5792), .ZN(n5794) );
  NOR2_X1 U7312 ( .A1(n5795), .A2(n5794), .ZN(n5799) );
  AOI21_X1 U7313 ( .B1(n5795), .B2(n5794), .A(n5799), .ZN(n9124) );
  NAND2_X1 U7314 ( .A1(n7946), .A2(n5703), .ZN(n5797) );
  NAND2_X1 U7315 ( .A1(n9453), .A2(n5780), .ZN(n5796) );
  NAND2_X1 U7316 ( .A1(n5797), .A2(n5796), .ZN(n5798) );
  XNOR2_X1 U7317 ( .A(n5798), .B(n5886), .ZN(n5806) );
  AOI22_X1 U7318 ( .A1(n7946), .A2(n5853), .B1(n5707), .B2(n9453), .ZN(n5804)
         );
  XNOR2_X1 U7319 ( .A(n5806), .B(n5804), .ZN(n9136) );
  AND2_X1 U7320 ( .A1(n9124), .A2(n9136), .ZN(n5803) );
  INV_X1 U7321 ( .A(n9136), .ZN(n5800) );
  INV_X1 U7322 ( .A(n5799), .ZN(n9132) );
  INV_X1 U7323 ( .A(n5804), .ZN(n5805) );
  NAND2_X1 U7324 ( .A1(n9793), .A2(n5703), .ZN(n5808) );
  NAND2_X1 U7325 ( .A1(n9452), .A2(n5853), .ZN(n5807) );
  NAND2_X1 U7326 ( .A1(n5808), .A2(n5807), .ZN(n5809) );
  XNOR2_X1 U7327 ( .A(n5809), .B(n5886), .ZN(n5813) );
  NAND2_X1 U7328 ( .A1(n9793), .A2(n5853), .ZN(n5811) );
  NAND2_X1 U7329 ( .A1(n9452), .A2(n5707), .ZN(n5810) );
  NAND2_X1 U7330 ( .A1(n5811), .A2(n5810), .ZN(n5812) );
  NOR2_X1 U7331 ( .A1(n5813), .A2(n5812), .ZN(n9175) );
  NAND2_X1 U7332 ( .A1(n5813), .A2(n5812), .ZN(n9176) );
  NAND2_X1 U7333 ( .A1(n9787), .A2(n5703), .ZN(n5815) );
  NAND2_X1 U7334 ( .A1(n9451), .A2(n5853), .ZN(n5814) );
  NAND2_X1 U7335 ( .A1(n5815), .A2(n5814), .ZN(n5816) );
  XNOR2_X1 U7336 ( .A(n5816), .B(n5874), .ZN(n5819) );
  AND2_X1 U7337 ( .A1(n9451), .A2(n5707), .ZN(n5817) );
  AOI21_X1 U7338 ( .B1(n9787), .B2(n5853), .A(n5817), .ZN(n5818) );
  NOR2_X1 U7339 ( .A1(n5819), .A2(n5818), .ZN(n9093) );
  NAND2_X1 U7340 ( .A1(n5819), .A2(n5818), .ZN(n9091) );
  OAI22_X1 U7341 ( .A1(n9781), .A2(n5820), .B1(n9107), .B2(n5724), .ZN(n5821)
         );
  XNOR2_X1 U7342 ( .A(n5821), .B(n5886), .ZN(n5823) );
  OAI22_X1 U7343 ( .A1(n9781), .A2(n5724), .B1(n9107), .B2(n5782), .ZN(n5822)
         );
  NOR2_X1 U7344 ( .A1(n5823), .A2(n5822), .ZN(n5824) );
  AOI21_X1 U7345 ( .B1(n5823), .B2(n5822), .A(n5824), .ZN(n9158) );
  NAND2_X1 U7346 ( .A1(n9157), .A2(n9158), .ZN(n9156) );
  INV_X1 U7347 ( .A(n5824), .ZN(n5825) );
  NAND2_X1 U7348 ( .A1(n9156), .A2(n5825), .ZN(n9104) );
  NAND2_X1 U7349 ( .A1(n9831), .A2(n5703), .ZN(n5827) );
  NAND2_X1 U7350 ( .A1(n9450), .A2(n5853), .ZN(n5826) );
  NAND2_X1 U7351 ( .A1(n5827), .A2(n5826), .ZN(n5828) );
  XNOR2_X1 U7352 ( .A(n5828), .B(n5886), .ZN(n5831) );
  AOI22_X1 U7353 ( .A1(n9831), .A2(n5853), .B1(n5707), .B2(n9450), .ZN(n5829)
         );
  XNOR2_X1 U7354 ( .A(n5831), .B(n5829), .ZN(n9105) );
  NAND2_X1 U7355 ( .A1(n9104), .A2(n9105), .ZN(n9103) );
  INV_X1 U7356 ( .A(n5829), .ZN(n5830) );
  NAND2_X1 U7357 ( .A1(n9103), .A2(n5832), .ZN(n5837) );
  INV_X1 U7358 ( .A(n5837), .ZN(n5835) );
  AOI22_X1 U7359 ( .A1(n9647), .A2(n5703), .B1(n5853), .B2(n9449), .ZN(n5833)
         );
  XNOR2_X1 U7360 ( .A(n5833), .B(n5886), .ZN(n5836) );
  INV_X1 U7361 ( .A(n5836), .ZN(n5834) );
  NAND2_X1 U7362 ( .A1(n5835), .A2(n5834), .ZN(n5838) );
  NAND2_X1 U7363 ( .A1(n5837), .A2(n5836), .ZN(n9079) );
  OAI22_X1 U7364 ( .A1(n4482), .A2(n5724), .B1(n9085), .B2(n5782), .ZN(n9167)
         );
  NAND2_X1 U7365 ( .A1(n9824), .A2(n5703), .ZN(n5841) );
  NAND2_X1 U7366 ( .A1(n9448), .A2(n5780), .ZN(n5840) );
  NAND2_X1 U7367 ( .A1(n5841), .A2(n5840), .ZN(n5842) );
  XNOR2_X1 U7368 ( .A(n5842), .B(n5874), .ZN(n5844) );
  AND2_X1 U7369 ( .A1(n9448), .A2(n5707), .ZN(n5843) );
  AOI21_X1 U7370 ( .B1(n9824), .B2(n5853), .A(n5843), .ZN(n5845) );
  INV_X1 U7371 ( .A(n5844), .ZN(n5847) );
  INV_X1 U7372 ( .A(n5845), .ZN(n5846) );
  NAND2_X1 U7373 ( .A1(n5847), .A2(n5846), .ZN(n5848) );
  NAND2_X1 U7374 ( .A1(n9624), .A2(n5703), .ZN(n5850) );
  NAND2_X1 U7375 ( .A1(n9447), .A2(n5780), .ZN(n5849) );
  NAND2_X1 U7376 ( .A1(n5850), .A2(n5849), .ZN(n5851) );
  XNOR2_X1 U7377 ( .A(n5851), .B(n5874), .ZN(n5854) );
  AND2_X1 U7378 ( .A1(n9447), .A2(n5707), .ZN(n5852) );
  AOI21_X1 U7379 ( .B1(n9624), .B2(n5853), .A(n5852), .ZN(n5855) );
  NAND2_X1 U7380 ( .A1(n5854), .A2(n5855), .ZN(n5860) );
  INV_X1 U7381 ( .A(n5854), .ZN(n5857) );
  INV_X1 U7382 ( .A(n5855), .ZN(n5856) );
  NAND2_X1 U7383 ( .A1(n5857), .A2(n5856), .ZN(n5858) );
  OAI22_X1 U7384 ( .A1(n9817), .A2(n5724), .B1(n6430), .B2(n5782), .ZN(n5869)
         );
  NAND2_X1 U7385 ( .A1(n9611), .A2(n5703), .ZN(n5862) );
  NAND2_X1 U7386 ( .A1(n9446), .A2(n5780), .ZN(n5861) );
  NAND2_X1 U7387 ( .A1(n5862), .A2(n5861), .ZN(n5863) );
  XNOR2_X1 U7388 ( .A(n5863), .B(n5886), .ZN(n5868) );
  NAND2_X1 U7389 ( .A1(n9812), .A2(n5703), .ZN(n5865) );
  NAND2_X1 U7390 ( .A1(n9445), .A2(n5780), .ZN(n5864) );
  NAND2_X1 U7391 ( .A1(n5865), .A2(n5864), .ZN(n5866) );
  XNOR2_X1 U7392 ( .A(n5866), .B(n5886), .ZN(n5883) );
  AND2_X1 U7393 ( .A1(n9445), .A2(n5707), .ZN(n5867) );
  AOI21_X1 U7394 ( .B1(n9812), .B2(n5853), .A(n5867), .ZN(n5881) );
  XNOR2_X1 U7395 ( .A(n5883), .B(n5881), .ZN(n6428) );
  INV_X1 U7396 ( .A(n5868), .ZN(n5871) );
  INV_X1 U7397 ( .A(n5869), .ZN(n5870) );
  NAND2_X1 U7398 ( .A1(n5871), .A2(n5870), .ZN(n6427) );
  NAND2_X1 U7399 ( .A1(n9583), .A2(n5703), .ZN(n5873) );
  NAND2_X1 U7400 ( .A1(n9444), .A2(n5780), .ZN(n5872) );
  NAND2_X1 U7401 ( .A1(n5873), .A2(n5872), .ZN(n5875) );
  XNOR2_X1 U7402 ( .A(n5875), .B(n5874), .ZN(n5878) );
  INV_X1 U7403 ( .A(n5878), .ZN(n5880) );
  AND2_X1 U7404 ( .A1(n9444), .A2(n5707), .ZN(n5876) );
  AOI21_X1 U7405 ( .B1(n9583), .B2(n5853), .A(n5876), .ZN(n5877) );
  INV_X1 U7406 ( .A(n5877), .ZN(n5879) );
  AOI21_X1 U7407 ( .B1(n5880), .B2(n5879), .A(n5896), .ZN(n9061) );
  INV_X1 U7408 ( .A(n5881), .ZN(n5882) );
  NAND2_X1 U7409 ( .A1(n5883), .A2(n5882), .ZN(n9062) );
  AND2_X2 U7410 ( .A1(n9063), .A2(n4909), .ZN(n9065) );
  INV_X1 U7411 ( .A(n9065), .ZN(n5895) );
  NAND2_X1 U7412 ( .A1(n9568), .A2(n5703), .ZN(n5885) );
  NAND2_X1 U7413 ( .A1(n9443), .A2(n5780), .ZN(n5884) );
  NAND2_X1 U7414 ( .A1(n5885), .A2(n5884), .ZN(n5887) );
  XNOR2_X1 U7415 ( .A(n5887), .B(n5886), .ZN(n5889) );
  AOI22_X1 U7416 ( .A1(n9568), .A2(n5853), .B1(n5707), .B2(n9443), .ZN(n5888)
         );
  XNOR2_X1 U7417 ( .A(n5889), .B(n5888), .ZN(n5897) );
  INV_X1 U7418 ( .A(n5897), .ZN(n5894) );
  OAI211_X1 U7419 ( .C1(n5892), .C2(n5891), .A(n5890), .B(n7032), .ZN(n5903)
         );
  NOR2_X1 U7420 ( .A1(n5903), .A2(n9292), .ZN(n5899) );
  INV_X1 U7421 ( .A(n9993), .ZN(n10039) );
  AND2_X1 U7422 ( .A1(n10039), .A2(n9432), .ZN(n5893) );
  NAND2_X1 U7423 ( .A1(n5895), .A2(n4900), .ZN(n5913) );
  NAND3_X1 U7424 ( .A1(n9065), .A2(n9865), .A3(n5897), .ZN(n5912) );
  NOR2_X1 U7425 ( .A1(n6625), .A2(n9298), .ZN(n7043) );
  NAND2_X1 U7426 ( .A1(n5899), .A2(n7043), .ZN(n5898) );
  NAND2_X1 U7427 ( .A1(n5898), .A2(n9727), .ZN(n9186) );
  NAND2_X1 U7428 ( .A1(n5899), .A2(n9290), .ZN(n9183) );
  NOR2_X1 U7429 ( .A1(n5900), .A2(n9183), .ZN(n5908) );
  AOI21_X1 U7430 ( .B1(n5903), .B2(n5902), .A(n5901), .ZN(n6618) );
  NAND2_X1 U7431 ( .A1(n6618), .A2(n5904), .ZN(n5905) );
  NAND2_X1 U7432 ( .A1(n5905), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9868) );
  OAI22_X1 U7433 ( .A1(n9566), .A2(n9868), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n5906), .ZN(n5907) );
  AOI211_X1 U7434 ( .C1(n9568), .C2(n9186), .A(n5908), .B(n5907), .ZN(n5909)
         );
  INV_X1 U7435 ( .A(n5909), .ZN(n5910) );
  NAND3_X1 U7436 ( .A1(n5913), .A2(n5912), .A3(n5911), .ZN(P1_U3220) );
  NOR2_X1 U7437 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n5918) );
  NAND4_X1 U7438 ( .A1(n5918), .A2(n5917), .A3(n6003), .A4(n5916), .ZN(n5919)
         );
  INV_X1 U7439 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5920) );
  NAND4_X1 U7440 ( .A1(n5921), .A2(n5920), .A3(n6135), .A4(n6134), .ZN(n5923)
         );
  NAND4_X1 U7441 ( .A1(n6150), .A2(n6133), .A3(n6082), .A4(n6163), .ZN(n5922)
         );
  NOR2_X1 U7442 ( .A1(n5923), .A2(n5922), .ZN(n5924) );
  INV_X1 U7443 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5926) );
  AND2_X1 U7444 ( .A1(n5926), .A2(n6294), .ZN(n5927) );
  INV_X1 U7445 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n6293) );
  INV_X1 U7446 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5945) );
  INV_X1 U7447 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6394) );
  INV_X1 U7448 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6368) );
  INV_X1 U7449 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n6372) );
  NAND2_X1 U7450 ( .A1(n6368), .A2(n6372), .ZN(n5942) );
  INV_X1 U7451 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5949) );
  INV_X1 U7452 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n5932) );
  NAND2_X1 U7453 ( .A1(n5934), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5935) );
  XNOR2_X1 U7454 ( .A(n5935), .B(P2_IR_REG_29__SCAN_IN), .ZN(n5936) );
  NAND2_X1 U7455 ( .A1(n5983), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5941) );
  NAND2_X1 U7456 ( .A1(n6197), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5940) );
  INV_X1 U7457 ( .A(n8181), .ZN(n5937) );
  NAND2_X1 U7458 ( .A1(n5973), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5938) );
  NAND2_X1 U7459 ( .A1(n5942), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5943) );
  NAND2_X1 U7460 ( .A1(n8144), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n5944) );
  NAND2_X1 U7461 ( .A1(n6374), .A2(n5945), .ZN(n5948) );
  OAI21_X1 U7462 ( .B1(n8144), .B2(P2_IR_REG_27__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5946) );
  OAI21_X1 U7463 ( .B1(P2_IR_REG_31__SCAN_IN), .B2(P2_IR_REG_27__SCAN_IN), .A(
        n5946), .ZN(n5947) );
  NAND2_X1 U7464 ( .A1(n6443), .A2(n6447), .ZN(n8368) );
  NAND2_X1 U7465 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5953) );
  XNOR2_X1 U7466 ( .A(n4896), .B(n5953), .ZN(n6509) );
  INV_X1 U7467 ( .A(n6540), .ZN(n5954) );
  NAND2_X1 U7468 ( .A1(n6299), .A2(n6859), .ZN(n8431) );
  NAND2_X1 U7469 ( .A1(n5983), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5960) );
  NAND2_X1 U7470 ( .A1(n6197), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5959) );
  INV_X1 U7471 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n5956) );
  NAND2_X1 U7472 ( .A1(n5973), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5957) );
  NAND2_X1 U7473 ( .A1(n8358), .A2(SI_0_), .ZN(n5962) );
  INV_X1 U7474 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5961) );
  XNOR2_X1 U7475 ( .A(n5962), .B(n5961), .ZN(n9059) );
  MUX2_X1 U7476 ( .A(n6513), .B(n9059), .S(n6443), .Z(n8972) );
  NAND2_X1 U7477 ( .A1(n6752), .A2(n8425), .ZN(n6750) );
  NAND2_X1 U7478 ( .A1(n6750), .A2(n8428), .ZN(n6702) );
  NAND2_X1 U7479 ( .A1(n5983), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5966) );
  NAND2_X1 U7480 ( .A1(n6197), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5965) );
  NAND2_X1 U7481 ( .A1(n5972), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n5964) );
  NAND2_X1 U7482 ( .A1(n5973), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5963) );
  XNOR2_X2 U7483 ( .A(n5969), .B(P2_IR_REG_2__SCAN_IN), .ZN(n6564) );
  NAND2_X1 U7484 ( .A1(n6184), .A2(n6564), .ZN(n5970) );
  OAI211_X2 U7485 ( .C1(n6022), .C2(n6450), .A(n5971), .B(n5970), .ZN(n6865)
         );
  INV_X1 U7486 ( .A(n6704), .ZN(n8434) );
  NAND2_X1 U7487 ( .A1(n6702), .A2(n8434), .ZN(n6701) );
  OR2_X1 U7488 ( .A1(n8608), .A2(n8420), .ZN(n8419) );
  NAND2_X1 U7489 ( .A1(n6701), .A2(n8419), .ZN(n7107) );
  NAND2_X1 U7490 ( .A1(n5983), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5977) );
  NAND2_X1 U7491 ( .A1(n6197), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5976) );
  NAND2_X1 U7492 ( .A1(n5972), .A2(n5985), .ZN(n5975) );
  NAND2_X1 U7493 ( .A1(n5973), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5974) );
  NAND4_X1 U7494 ( .A1(n5977), .A2(n5976), .A3(n5975), .A4(n5974), .ZN(n8607)
         );
  NAND2_X1 U7495 ( .A1(n6282), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n5981) );
  NAND2_X1 U7496 ( .A1(n5978), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5979) );
  XNOR2_X1 U7497 ( .A(n5979), .B(P2_IR_REG_3__SCAN_IN), .ZN(n6611) );
  NAND2_X1 U7498 ( .A1(n6184), .A2(n6611), .ZN(n5980) );
  INV_X1 U7499 ( .A(n7104), .ZN(n8381) );
  NAND2_X1 U7500 ( .A1(n7107), .A2(n8381), .ZN(n5982) );
  NAND2_X1 U7501 ( .A1(n5982), .A2(n8441), .ZN(n7094) );
  NAND2_X1 U7502 ( .A1(n5983), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5990) );
  NAND2_X1 U7503 ( .A1(n6197), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5989) );
  NAND2_X1 U7504 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5986) );
  NAND2_X1 U7505 ( .A1(n6009), .A2(n5986), .ZN(n7097) );
  NAND2_X1 U7506 ( .A1(n6216), .A2(n7097), .ZN(n5988) );
  NAND2_X1 U7507 ( .A1(n5973), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5987) );
  NAND4_X1 U7508 ( .A1(n5990), .A2(n5989), .A3(n5988), .A4(n5987), .ZN(n8606)
         );
  NAND2_X1 U7509 ( .A1(n6282), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n5994) );
  NAND2_X1 U7510 ( .A1(n5991), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5992) );
  XNOR2_X1 U7511 ( .A(n5992), .B(P2_IR_REG_4__SCAN_IN), .ZN(n6774) );
  NAND2_X1 U7512 ( .A1(n6184), .A2(n6774), .ZN(n5993) );
  OAI211_X1 U7513 ( .C1(n6022), .C2(n6456), .A(n5994), .B(n5993), .ZN(n10076)
         );
  XNOR2_X1 U7514 ( .A(n8606), .B(n10076), .ZN(n8439) );
  NAND2_X1 U7515 ( .A1(n7094), .A2(n8439), .ZN(n7096) );
  INV_X1 U7516 ( .A(n10076), .ZN(n8442) );
  OR2_X1 U7517 ( .A1(n8606), .A2(n8442), .ZN(n8459) );
  NAND2_X1 U7518 ( .A1(n5983), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6000) );
  INV_X2 U7519 ( .A(n6256), .ZN(n6359) );
  NAND2_X1 U7520 ( .A1(n6359), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5999) );
  OR2_X2 U7521 ( .A1(n6011), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6038) );
  NAND2_X1 U7522 ( .A1(n6011), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5996) );
  NAND2_X1 U7523 ( .A1(n6038), .A2(n5996), .ZN(n7158) );
  NAND2_X1 U7524 ( .A1(n5972), .A2(n7158), .ZN(n5998) );
  NAND2_X1 U7525 ( .A1(n5973), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5997) );
  NAND4_X1 U7526 ( .A1(n6000), .A2(n5999), .A3(n5998), .A4(n5997), .ZN(n8604)
         );
  OR2_X2 U7527 ( .A1(n5991), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n6016) );
  NOR2_X2 U7528 ( .A1(n6016), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n6004) );
  INV_X1 U7529 ( .A(n6004), .ZN(n6001) );
  NAND2_X1 U7530 ( .A1(n6001), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6002) );
  MUX2_X1 U7531 ( .A(n6002), .B(P2_IR_REG_31__SCAN_IN), .S(n6003), .Z(n6006)
         );
  AND2_X2 U7532 ( .A1(n6004), .A2(n6003), .ZN(n6032) );
  INV_X1 U7533 ( .A(n6032), .ZN(n6005) );
  INV_X2 U7534 ( .A(n6022), .ZN(n8365) );
  NAND2_X1 U7535 ( .A1(n6463), .A2(n8365), .ZN(n6008) );
  NAND2_X1 U7536 ( .A1(n6282), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n6007) );
  OAI211_X1 U7537 ( .C1(n6443), .C2(n6908), .A(n6008), .B(n6007), .ZN(n7147)
         );
  INV_X1 U7538 ( .A(n7147), .ZN(n10089) );
  NAND2_X1 U7539 ( .A1(n8604), .A2(n10089), .ZN(n6020) );
  NAND2_X1 U7540 ( .A1(n5983), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6015) );
  NAND2_X1 U7541 ( .A1(n6359), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n6014) );
  NAND2_X1 U7542 ( .A1(n6009), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n6010) );
  NAND2_X1 U7543 ( .A1(n6011), .A2(n6010), .ZN(n7214) );
  NAND2_X1 U7544 ( .A1(n5972), .A2(n7214), .ZN(n6013) );
  NAND2_X1 U7545 ( .A1(n6049), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6012) );
  NAND4_X1 U7546 ( .A1(n6015), .A2(n6014), .A3(n6013), .A4(n6012), .ZN(n8605)
         );
  NAND2_X1 U7547 ( .A1(n6282), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n6019) );
  NAND2_X1 U7548 ( .A1(n6016), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6017) );
  XNOR2_X1 U7549 ( .A(n6017), .B(P2_IR_REG_5__SCAN_IN), .ZN(n6810) );
  NAND2_X1 U7550 ( .A1(n6184), .A2(n6810), .ZN(n6018) );
  OAI211_X1 U7551 ( .C1(n6022), .C2(n6459), .A(n6019), .B(n6018), .ZN(n7212)
         );
  INV_X1 U7552 ( .A(n7212), .ZN(n10083) );
  NAND2_X1 U7553 ( .A1(n8605), .A2(n10083), .ZN(n7116) );
  AND2_X1 U7554 ( .A1(n6020), .A2(n7116), .ZN(n8462) );
  NOR2_X1 U7555 ( .A1(n8605), .A2(n10083), .ZN(n8457) );
  NAND2_X1 U7556 ( .A1(n8457), .A2(n6020), .ZN(n6021) );
  OR2_X1 U7557 ( .A1(n8604), .A2(n10089), .ZN(n8464) );
  AND2_X1 U7558 ( .A1(n6021), .A2(n8464), .ZN(n8445) );
  NAND2_X1 U7559 ( .A1(n6468), .A2(n8365), .ZN(n6025) );
  NOR2_X1 U7560 ( .A1(n6032), .A2(n6138), .ZN(n6023) );
  INV_X1 U7561 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n6031) );
  XNOR2_X1 U7562 ( .A(n6023), .B(n6031), .ZN(n6909) );
  AOI22_X1 U7563 ( .A1(n8362), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n6184), .B2(
        n6909), .ZN(n6024) );
  NAND2_X1 U7564 ( .A1(n6025), .A2(n6024), .ZN(n10094) );
  INV_X1 U7565 ( .A(n10094), .ZN(n6030) );
  NAND2_X1 U7566 ( .A1(n5983), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6029) );
  NAND2_X1 U7567 ( .A1(n6359), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n6028) );
  XNOR2_X1 U7568 ( .A(n6038), .B(P2_REG3_REG_7__SCAN_IN), .ZN(n7253) );
  NAND2_X1 U7569 ( .A1(n6216), .A2(n7253), .ZN(n6027) );
  NAND2_X1 U7570 ( .A1(n6049), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6026) );
  NAND4_X1 U7571 ( .A1(n6029), .A2(n6028), .A3(n6027), .A4(n6026), .ZN(n8603)
         );
  NAND2_X1 U7572 ( .A1(n6030), .A2(n8603), .ZN(n7051) );
  NAND2_X1 U7573 ( .A1(n7463), .A2(n10094), .ZN(n8449) );
  NAND2_X1 U7574 ( .A1(n7051), .A2(n8449), .ZN(n8466) );
  NAND2_X1 U7575 ( .A1(n6472), .A2(n8365), .ZN(n6035) );
  NAND2_X1 U7576 ( .A1(n6032), .A2(n6031), .ZN(n6045) );
  NAND2_X1 U7577 ( .A1(n6045), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6033) );
  XNOR2_X1 U7578 ( .A(n6033), .B(P2_IR_REG_8__SCAN_IN), .ZN(n8619) );
  AOI22_X1 U7579 ( .A1(n8362), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6184), .B2(
        n8619), .ZN(n6034) );
  NAND2_X1 U7580 ( .A1(n6035), .A2(n6034), .ZN(n7578) );
  NAND2_X1 U7581 ( .A1(n5983), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n6043) );
  NAND2_X1 U7582 ( .A1(n6359), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n6042) );
  NOR2_X1 U7583 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_REG3_REG_7__SCAN_IN), 
        .ZN(n6036) );
  OAI21_X1 U7584 ( .B1(n6038), .B2(P2_REG3_REG_7__SCAN_IN), .A(
        P2_REG3_REG_8__SCAN_IN), .ZN(n6039) );
  NAND2_X1 U7585 ( .A1(n6050), .A2(n6039), .ZN(n7055) );
  NAND2_X1 U7586 ( .A1(n5972), .A2(n7055), .ZN(n6041) );
  NAND2_X1 U7587 ( .A1(n6049), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n6040) );
  NAND4_X1 U7588 ( .A1(n6043), .A2(n6042), .A3(n6041), .A4(n6040), .ZN(n8602)
         );
  OR2_X1 U7589 ( .A1(n7578), .A2(n7474), .ZN(n8416) );
  AND2_X1 U7590 ( .A1(n8416), .A2(n7051), .ZN(n8418) );
  NAND2_X1 U7591 ( .A1(n7124), .A2(n8418), .ZN(n6044) );
  NAND2_X1 U7592 ( .A1(n7578), .A2(n7474), .ZN(n8450) );
  NAND2_X1 U7593 ( .A1(n6044), .A2(n8450), .ZN(n7134) );
  INV_X1 U7594 ( .A(n7134), .ZN(n6057) );
  NAND2_X1 U7595 ( .A1(n6484), .A2(n8365), .ZN(n6048) );
  OAI21_X1 U7596 ( .B1(n6045), .B2(P2_IR_REG_8__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6046) );
  XNOR2_X1 U7597 ( .A(n6046), .B(P2_IR_REG_9__SCAN_IN), .ZN(n7076) );
  AOI22_X1 U7598 ( .A1(n8362), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6184), .B2(
        n7076), .ZN(n6047) );
  NAND2_X1 U7599 ( .A1(n6048), .A2(n6047), .ZN(n7468) );
  NAND2_X1 U7600 ( .A1(n6359), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n6055) );
  NAND2_X1 U7601 ( .A1(n6049), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6054) );
  NAND2_X1 U7602 ( .A1(n6050), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n6051) );
  NAND2_X1 U7603 ( .A1(n6065), .A2(n6051), .ZN(n7141) );
  NAND2_X1 U7604 ( .A1(n5972), .A2(n7141), .ZN(n6053) );
  NAND2_X1 U7605 ( .A1(n5983), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n6052) );
  NAND4_X1 U7606 ( .A1(n6055), .A2(n6054), .A3(n6053), .A4(n6052), .ZN(n8601)
         );
  NAND2_X1 U7607 ( .A1(n7468), .A2(n7716), .ZN(n8452) );
  NAND2_X1 U7608 ( .A1(n8417), .A2(n8452), .ZN(n8387) );
  INV_X1 U7609 ( .A(n8387), .ZN(n6056) );
  NAND2_X1 U7610 ( .A1(n6480), .A2(n8365), .ZN(n6063) );
  NOR2_X1 U7611 ( .A1(n6060), .A2(n6138), .ZN(n6058) );
  MUX2_X1 U7612 ( .A(n6138), .B(n6058), .S(P2_IR_REG_10__SCAN_IN), .Z(n6061)
         );
  OR2_X1 U7613 ( .A1(n6061), .A2(n6083), .ZN(n7395) );
  INV_X1 U7614 ( .A(n7395), .ZN(n7067) );
  AOI22_X1 U7615 ( .A1(n8362), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6184), .B2(
        n7067), .ZN(n6062) );
  NAND2_X1 U7616 ( .A1(n5983), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n6071) );
  NAND2_X1 U7617 ( .A1(n6359), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n6070) );
  INV_X1 U7618 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n7083) );
  NAND2_X1 U7619 ( .A1(n6065), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6066) );
  NAND2_X1 U7620 ( .A1(n6075), .A2(n6066), .ZN(n7456) );
  NAND2_X1 U7621 ( .A1(n6216), .A2(n7456), .ZN(n6069) );
  NAND2_X1 U7622 ( .A1(n6049), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6068) );
  NAND2_X1 U7623 ( .A1(n7796), .A2(n7717), .ZN(n8473) );
  NAND2_X1 U7624 ( .A1(n6500), .A2(n8365), .ZN(n6074) );
  OR2_X1 U7625 ( .A1(n6083), .A2(n6138), .ZN(n6072) );
  XNOR2_X1 U7626 ( .A(n6072), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7519) );
  AOI22_X1 U7627 ( .A1(n8362), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6184), .B2(
        n7519), .ZN(n6073) );
  NAND2_X1 U7628 ( .A1(n5983), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n6080) );
  NAND2_X1 U7629 ( .A1(n6359), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n6079) );
  NAND2_X1 U7630 ( .A1(n6075), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6076) );
  NAND2_X1 U7631 ( .A1(n6087), .A2(n6076), .ZN(n7482) );
  NAND2_X1 U7632 ( .A1(n6216), .A2(n7482), .ZN(n6078) );
  NAND2_X1 U7633 ( .A1(n6049), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n6077) );
  NAND4_X1 U7634 ( .A1(n6080), .A2(n6079), .A3(n6078), .A4(n6077), .ZN(n8599)
         );
  INV_X1 U7635 ( .A(n8599), .ZN(n7792) );
  NAND2_X1 U7636 ( .A1(n10124), .A2(n7792), .ZN(n8478) );
  NAND2_X1 U7637 ( .A1(n7479), .A2(n8478), .ZN(n6081) );
  OR2_X1 U7638 ( .A1(n10124), .A2(n7792), .ZN(n8476) );
  NAND2_X1 U7639 ( .A1(n6081), .A2(n8476), .ZN(n7625) );
  NAND2_X1 U7640 ( .A1(n6526), .A2(n8365), .ZN(n6086) );
  NAND2_X1 U7641 ( .A1(n6083), .A2(n6082), .ZN(n6093) );
  NAND2_X1 U7642 ( .A1(n6093), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6084) );
  XNOR2_X1 U7643 ( .A(n6084), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7528) );
  AOI22_X1 U7644 ( .A1(n8362), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6184), .B2(
        n7528), .ZN(n6085) );
  NAND2_X1 U7645 ( .A1(n6359), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n6092) );
  NAND2_X1 U7646 ( .A1(n5983), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n6091) );
  NAND2_X1 U7647 ( .A1(n6087), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6088) );
  NAND2_X1 U7648 ( .A1(n6099), .A2(n6088), .ZN(n7623) );
  NAND2_X1 U7649 ( .A1(n6216), .A2(n7623), .ZN(n6090) );
  NAND2_X1 U7650 ( .A1(n6049), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n6089) );
  NAND4_X1 U7651 ( .A1(n6092), .A2(n6091), .A3(n6090), .A4(n6089), .ZN(n8598)
         );
  XNOR2_X1 U7652 ( .A(n10131), .B(n8598), .ZN(n8377) );
  NAND2_X1 U7653 ( .A1(n7625), .A2(n8377), .ZN(n7626) );
  INV_X1 U7654 ( .A(n8598), .ZN(n8482) );
  OR2_X1 U7655 ( .A1(n10131), .A2(n8482), .ZN(n8484) );
  NAND2_X1 U7656 ( .A1(n7626), .A2(n8484), .ZN(n7669) );
  NAND2_X1 U7657 ( .A1(n6538), .A2(n8365), .ZN(n6096) );
  NAND2_X1 U7658 ( .A1(n6137), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6108) );
  XNOR2_X1 U7659 ( .A(n6108), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7751) );
  AOI22_X1 U7660 ( .A1(n8362), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6184), .B2(
        n7751), .ZN(n6095) );
  NAND2_X1 U7661 ( .A1(n5983), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n6104) );
  NAND2_X1 U7662 ( .A1(n6359), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n6103) );
  INV_X1 U7663 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n6097) );
  NAND2_X1 U7664 ( .A1(n6099), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n6100) );
  NAND2_X1 U7665 ( .A1(n6116), .A2(n6100), .ZN(n7826) );
  NAND2_X1 U7666 ( .A1(n6216), .A2(n7826), .ZN(n6102) );
  NAND2_X1 U7667 ( .A1(n6049), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n6101) );
  NAND4_X1 U7668 ( .A1(n6104), .A2(n6103), .A3(n6102), .A4(n6101), .ZN(n8597)
         );
  NAND2_X1 U7669 ( .A1(n8488), .A2(n4882), .ZN(n6105) );
  NAND2_X1 U7670 ( .A1(n7669), .A2(n6105), .ZN(n6107) );
  OR2_X1 U7671 ( .A1(n8488), .A2(n4882), .ZN(n6106) );
  NAND2_X1 U7672 ( .A1(n6711), .A2(n8365), .ZN(n6113) );
  NAND2_X1 U7673 ( .A1(n6108), .A2(n6134), .ZN(n6109) );
  NAND2_X1 U7674 ( .A1(n6109), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6110) );
  NAND2_X1 U7675 ( .A1(n6110), .A2(n6135), .ZN(n6122) );
  OR2_X1 U7676 ( .A1(n6110), .A2(n6135), .ZN(n6111) );
  NAND2_X1 U7677 ( .A1(n6122), .A2(n6111), .ZN(n8652) );
  INV_X1 U7678 ( .A(n8652), .ZN(n7748) );
  AOI22_X1 U7679 ( .A1(n8362), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6184), .B2(
        n7748), .ZN(n6112) );
  NAND2_X1 U7680 ( .A1(n6359), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n6121) );
  NAND2_X1 U7681 ( .A1(n6049), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n6120) );
  INV_X1 U7682 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n6114) );
  NAND2_X1 U7683 ( .A1(n6116), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6117) );
  NAND2_X1 U7684 ( .A1(n6126), .A2(n6117), .ZN(n7905) );
  NAND2_X1 U7685 ( .A1(n6216), .A2(n7905), .ZN(n6119) );
  NAND2_X1 U7686 ( .A1(n5983), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n6118) );
  NAND4_X1 U7687 ( .A1(n6121), .A2(n6120), .A3(n6119), .A4(n6118), .ZN(n8596)
         );
  INV_X1 U7688 ( .A(n8596), .ZN(n7927) );
  NOR2_X1 U7689 ( .A1(n7909), .A2(n7927), .ZN(n8498) );
  NAND2_X1 U7690 ( .A1(n7909), .A2(n7927), .ZN(n7650) );
  NAND2_X1 U7691 ( .A1(n6852), .A2(n8365), .ZN(n6125) );
  NAND2_X1 U7692 ( .A1(n6122), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6123) );
  XNOR2_X1 U7693 ( .A(n6123), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8673) );
  AOI22_X1 U7694 ( .A1(n6282), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n6184), .B2(
        n8673), .ZN(n6124) );
  NAND2_X1 U7695 ( .A1(n5983), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n6131) );
  NAND2_X1 U7696 ( .A1(n6359), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n6130) );
  OR2_X2 U7697 ( .A1(n6126), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6144) );
  NAND2_X1 U7698 ( .A1(n6126), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6127) );
  NAND2_X1 U7699 ( .A1(n6144), .A2(n6127), .ZN(n7935) );
  NAND2_X1 U7700 ( .A1(n6216), .A2(n7935), .ZN(n6129) );
  NAND2_X1 U7701 ( .A1(n6049), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n6128) );
  NAND4_X1 U7702 ( .A1(n6131), .A2(n6130), .A3(n6129), .A4(n6128), .ZN(n8595)
         );
  INV_X1 U7703 ( .A(n8595), .ZN(n8203) );
  NAND2_X1 U7704 ( .A1(n7930), .A2(n8203), .ZN(n8502) );
  INV_X1 U7705 ( .A(n8502), .ZN(n6132) );
  OR2_X1 U7706 ( .A1(n7930), .A2(n8203), .ZN(n8513) );
  NAND2_X1 U7707 ( .A1(n6921), .A2(n8365), .ZN(n6141) );
  NAND3_X1 U7708 ( .A1(n6135), .A2(n6134), .A3(n6133), .ZN(n6136) );
  OR2_X1 U7709 ( .A1(n6151), .A2(n6138), .ZN(n6139) );
  XNOR2_X1 U7710 ( .A(n6139), .B(P2_IR_REG_16__SCAN_IN), .ZN(n8675) );
  AOI22_X1 U7711 ( .A1(n8362), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6184), .B2(
        n8675), .ZN(n6140) );
  NAND2_X1 U7712 ( .A1(n5983), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n6149) );
  NAND2_X1 U7713 ( .A1(n6359), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n6148) );
  INV_X1 U7714 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n6142) );
  NAND2_X1 U7715 ( .A1(n6144), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6145) );
  NAND2_X1 U7716 ( .A1(n6155), .A2(n6145), .ZN(n8285) );
  NAND2_X1 U7717 ( .A1(n6216), .A2(n8285), .ZN(n6147) );
  NAND2_X1 U7718 ( .A1(n6049), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n6146) );
  NAND4_X1 U7719 ( .A1(n6149), .A2(n6148), .A3(n6147), .A4(n6146), .ZN(n8594)
         );
  INV_X1 U7720 ( .A(n8594), .ZN(n8204) );
  OR2_X1 U7721 ( .A1(n8966), .A2(n8204), .ZN(n8512) );
  NAND2_X1 U7722 ( .A1(n8966), .A2(n8204), .ZN(n8515) );
  NAND2_X1 U7723 ( .A1(n8512), .A2(n8515), .ZN(n7866) );
  NAND2_X1 U7724 ( .A1(n7013), .A2(n8365), .ZN(n6154) );
  NAND2_X1 U7725 ( .A1(n6151), .A2(n6150), .ZN(n6162) );
  NAND2_X1 U7726 ( .A1(n6162), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6152) );
  XNOR2_X1 U7727 ( .A(n6152), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8728) );
  AOI22_X1 U7728 ( .A1(n8362), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6184), .B2(
        n8728), .ZN(n6153) );
  NAND2_X1 U7729 ( .A1(n6359), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n6160) );
  NAND2_X1 U7730 ( .A1(n5983), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n6159) );
  OR2_X2 U7731 ( .A1(n6155), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n6173) );
  NAND2_X1 U7732 ( .A1(n6155), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n6156) );
  NAND2_X1 U7733 ( .A1(n6173), .A2(n6156), .ZN(n8300) );
  NAND2_X1 U7734 ( .A1(n6216), .A2(n8300), .ZN(n6158) );
  NAND2_X1 U7735 ( .A1(n6049), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n6157) );
  NAND4_X1 U7736 ( .A1(n6160), .A2(n6159), .A3(n6158), .A4(n6157), .ZN(n8593)
         );
  INV_X1 U7737 ( .A(n8593), .ZN(n8283) );
  NAND2_X1 U7738 ( .A1(n8289), .A2(n8283), .ZN(n8505) );
  NAND2_X1 U7739 ( .A1(n6161), .A2(n8505), .ZN(n7953) );
  INV_X1 U7740 ( .A(n7953), .ZN(n6180) );
  NAND2_X1 U7741 ( .A1(n7102), .A2(n8365), .ZN(n6170) );
  INV_X1 U7742 ( .A(n6162), .ZN(n6164) );
  NAND2_X1 U7743 ( .A1(n6164), .A2(n6163), .ZN(n6165) );
  INV_X1 U7744 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n6166) );
  NAND2_X1 U7745 ( .A1(n6167), .A2(n6166), .ZN(n6181) );
  OR2_X1 U7746 ( .A1(n6167), .A2(n6166), .ZN(n6168) );
  AND2_X1 U7747 ( .A1(n6181), .A2(n6168), .ZN(n8747) );
  AOI22_X1 U7748 ( .A1(n8362), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6184), .B2(
        n8747), .ZN(n6169) );
  NAND2_X1 U7749 ( .A1(n6359), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n6178) );
  NAND2_X1 U7750 ( .A1(n6049), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n6177) );
  INV_X1 U7751 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n6171) );
  NAND2_X1 U7752 ( .A1(n6173), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6174) );
  NAND2_X1 U7753 ( .A1(n6187), .A2(n6174), .ZN(n8336) );
  NAND2_X1 U7754 ( .A1(n6216), .A2(n8336), .ZN(n6176) );
  NAND2_X1 U7755 ( .A1(n5983), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n6175) );
  NAND4_X1 U7756 ( .A1(n6178), .A2(n6177), .A3(n6176), .A4(n6175), .ZN(n8897)
         );
  INV_X1 U7757 ( .A(n8897), .ZN(n8298) );
  NAND2_X1 U7758 ( .A1(n8959), .A2(n8298), .ZN(n8506) );
  NAND2_X1 U7759 ( .A1(n8521), .A2(n8506), .ZN(n8397) );
  INV_X1 U7760 ( .A(n8397), .ZN(n6179) );
  NAND2_X1 U7761 ( .A1(n6180), .A2(n6179), .ZN(n7955) );
  NAND2_X1 U7762 ( .A1(n7955), .A2(n8521), .ZN(n8903) );
  NAND2_X1 U7763 ( .A1(n7275), .A2(n8365), .ZN(n6186) );
  INV_X1 U7764 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n6182) );
  XNOR2_X1 U7765 ( .A(n6183), .B(n6182), .ZN(n6725) );
  AOI22_X1 U7766 ( .A1(n8362), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n6184), .B2(
        n6399), .ZN(n6185) );
  OR2_X2 U7767 ( .A1(n6187), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6195) );
  NAND2_X1 U7768 ( .A1(n6187), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6188) );
  NAND2_X1 U7769 ( .A1(n6195), .A2(n6188), .ZN(n8907) );
  AOI22_X1 U7770 ( .A1(n8907), .A2(n6216), .B1(n5983), .B2(
        P2_REG1_REG_19__SCAN_IN), .ZN(n6190) );
  AOI22_X1 U7771 ( .A1(n6359), .A2(P2_REG0_REG_19__SCAN_IN), .B1(n6049), .B2(
        P2_REG2_REG_19__SCAN_IN), .ZN(n6189) );
  NAND2_X1 U7772 ( .A1(n8954), .A2(n8334), .ZN(n8507) );
  NAND2_X1 U7773 ( .A1(n8411), .A2(n8507), .ZN(n8904) );
  INV_X1 U7774 ( .A(n8904), .ZN(n8893) );
  NAND2_X1 U7775 ( .A1(n7356), .A2(n8365), .ZN(n6192) );
  NAND2_X1 U7776 ( .A1(n6282), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n6191) );
  INV_X1 U7777 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8886) );
  INV_X1 U7778 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n6193) );
  NAND2_X1 U7779 ( .A1(n6195), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6196) );
  NAND2_X1 U7780 ( .A1(n6203), .A2(n6196), .ZN(n8887) );
  NAND2_X1 U7781 ( .A1(n8887), .A2(n6216), .ZN(n6199) );
  AOI22_X1 U7782 ( .A1(n5983), .A2(P2_REG1_REG_20__SCAN_IN), .B1(n6197), .B2(
        P2_REG0_REG_20__SCAN_IN), .ZN(n6198) );
  OAI211_X1 U7783 ( .C1(n6067), .C2(n8886), .A(n6199), .B(n6198), .ZN(n8900)
         );
  INV_X1 U7784 ( .A(n8900), .ZN(n8268) );
  INV_X1 U7785 ( .A(n8408), .ZN(n6200) );
  NAND2_X1 U7786 ( .A1(n9032), .A2(n8268), .ZN(n8508) );
  NAND2_X1 U7787 ( .A1(n7532), .A2(n8365), .ZN(n6202) );
  NAND2_X1 U7788 ( .A1(n6282), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n6201) );
  INV_X1 U7789 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n8875) );
  NAND2_X1 U7790 ( .A1(n6203), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n6204) );
  NAND2_X1 U7791 ( .A1(n6211), .A2(n6204), .ZN(n8876) );
  NAND2_X1 U7792 ( .A1(n8876), .A2(n6216), .ZN(n6206) );
  AOI22_X1 U7793 ( .A1(n5983), .A2(P2_REG1_REG_21__SCAN_IN), .B1(n6359), .B2(
        P2_REG0_REG_21__SCAN_IN), .ZN(n6205) );
  OAI211_X1 U7794 ( .C1(n6067), .C2(n8875), .A(n6206), .B(n6205), .ZN(n8884)
         );
  INV_X1 U7795 ( .A(n8884), .ZN(n8857) );
  NAND2_X1 U7796 ( .A1(n9026), .A2(n8857), .ZN(n8532) );
  NAND2_X1 U7797 ( .A1(n7595), .A2(n8365), .ZN(n6208) );
  NAND2_X1 U7798 ( .A1(n6282), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n6207) );
  INV_X1 U7799 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n6209) );
  NAND2_X1 U7800 ( .A1(n6211), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6212) );
  NAND2_X1 U7801 ( .A1(n6228), .A2(n6212), .ZN(n8861) );
  INV_X1 U7802 ( .A(n5983), .ZN(n6277) );
  INV_X1 U7803 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8941) );
  NAND2_X1 U7804 ( .A1(n6049), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n6214) );
  NAND2_X1 U7805 ( .A1(n6359), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n6213) );
  OAI211_X1 U7806 ( .C1(n6277), .C2(n8941), .A(n6214), .B(n6213), .ZN(n6215)
         );
  AOI21_X1 U7807 ( .B1(n8861), .B2(n6216), .A(n6215), .ZN(n8843) );
  NAND2_X1 U7808 ( .A1(n9020), .A2(n8843), .ZN(n8531) );
  NAND2_X1 U7809 ( .A1(n8862), .A2(n8531), .ZN(n6217) );
  NAND2_X1 U7810 ( .A1(n6217), .A2(n8535), .ZN(n8845) );
  NAND2_X1 U7811 ( .A1(n7761), .A2(n8365), .ZN(n6219) );
  NAND2_X1 U7812 ( .A1(n6282), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n6218) );
  OR2_X2 U7813 ( .A1(n6228), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6230) );
  OR2_X2 U7814 ( .A1(n6230), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6243) );
  NAND2_X1 U7815 ( .A1(n6230), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6220) );
  NAND2_X1 U7816 ( .A1(n6243), .A2(n6220), .ZN(n8838) );
  NAND2_X1 U7817 ( .A1(n8838), .A2(n6216), .ZN(n6225) );
  INV_X1 U7818 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n9009) );
  NAND2_X1 U7819 ( .A1(n6049), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n6222) );
  NAND2_X1 U7820 ( .A1(n5983), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n6221) );
  OAI211_X1 U7821 ( .C1(n6256), .C2(n9009), .A(n6222), .B(n6221), .ZN(n6223)
         );
  INV_X1 U7822 ( .A(n6223), .ZN(n6224) );
  NAND2_X1 U7823 ( .A1(n6225), .A2(n6224), .ZN(n8816) );
  NAND2_X1 U7824 ( .A1(n9010), .A2(n8844), .ZN(n8404) );
  NAND2_X1 U7825 ( .A1(n7644), .A2(n8365), .ZN(n6227) );
  NAND2_X1 U7826 ( .A1(n6282), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n6226) );
  NAND2_X1 U7827 ( .A1(n6228), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6229) );
  NAND2_X1 U7828 ( .A1(n6230), .A2(n6229), .ZN(n8847) );
  NAND2_X1 U7829 ( .A1(n8847), .A2(n6216), .ZN(n6235) );
  INV_X1 U7830 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n8938) );
  NAND2_X1 U7831 ( .A1(n6049), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n6232) );
  NAND2_X1 U7832 ( .A1(n6359), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n6231) );
  OAI211_X1 U7833 ( .C1(n6277), .C2(n8938), .A(n6232), .B(n6231), .ZN(n6233)
         );
  INV_X1 U7834 ( .A(n6233), .ZN(n6234) );
  NAND2_X1 U7835 ( .A1(n8238), .A2(n8859), .ZN(n8827) );
  NAND2_X1 U7836 ( .A1(n8845), .A2(n8406), .ZN(n6238) );
  INV_X1 U7837 ( .A(n8406), .ZN(n6236) );
  NAND2_X1 U7838 ( .A1(n7798), .A2(n8365), .ZN(n6240) );
  NAND2_X1 U7839 ( .A1(n8362), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n6239) );
  INV_X1 U7840 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n6241) );
  NAND2_X1 U7841 ( .A1(n6243), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6244) );
  NAND2_X1 U7842 ( .A1(n6252), .A2(n6244), .ZN(n8820) );
  NAND2_X1 U7843 ( .A1(n8820), .A2(n6216), .ZN(n6249) );
  INV_X1 U7844 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n8930) );
  NAND2_X1 U7845 ( .A1(n6359), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n6246) );
  NAND2_X1 U7846 ( .A1(n6049), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n6245) );
  OAI211_X1 U7847 ( .C1(n8930), .C2(n6277), .A(n6246), .B(n6245), .ZN(n6247)
         );
  INV_X1 U7848 ( .A(n6247), .ZN(n6248) );
  NAND2_X1 U7849 ( .A1(n6249), .A2(n6248), .ZN(n8832) );
  NOR2_X1 U7850 ( .A1(n9004), .A2(n8805), .ZN(n8541) );
  NAND2_X1 U7851 ( .A1(n9004), .A2(n8805), .ZN(n8540) );
  NAND2_X1 U7852 ( .A1(n7830), .A2(n8365), .ZN(n6251) );
  NAND2_X1 U7853 ( .A1(n8362), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n6250) );
  NAND2_X1 U7854 ( .A1(n6252), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6253) );
  NAND2_X1 U7855 ( .A1(n6262), .A2(n6253), .ZN(n8807) );
  NAND2_X1 U7856 ( .A1(n8807), .A2(n6216), .ZN(n6259) );
  INV_X1 U7857 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8997) );
  NAND2_X1 U7858 ( .A1(n5983), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n6255) );
  NAND2_X1 U7859 ( .A1(n6049), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n6254) );
  OAI211_X1 U7860 ( .C1(n6256), .C2(n8997), .A(n6255), .B(n6254), .ZN(n6257)
         );
  INV_X1 U7861 ( .A(n6257), .ZN(n6258) );
  NAND2_X1 U7862 ( .A1(n7921), .A2(n8365), .ZN(n6261) );
  NAND2_X1 U7863 ( .A1(n8362), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n6260) );
  NAND2_X1 U7864 ( .A1(n6262), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6263) );
  NAND2_X1 U7865 ( .A1(n6273), .A2(n6263), .ZN(n8799) );
  NAND2_X1 U7866 ( .A1(n8799), .A2(n6216), .ZN(n6268) );
  INV_X1 U7867 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n8924) );
  NAND2_X1 U7868 ( .A1(n6359), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n6265) );
  NAND2_X1 U7869 ( .A1(n5973), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n6264) );
  OAI211_X1 U7870 ( .C1(n6277), .C2(n8924), .A(n6265), .B(n6264), .ZN(n6266)
         );
  INV_X1 U7871 ( .A(n6266), .ZN(n6267) );
  NAND2_X1 U7872 ( .A1(n8991), .A2(n8806), .ZN(n8547) );
  NAND2_X1 U7873 ( .A1(n7963), .A2(n8365), .ZN(n6271) );
  NAND2_X1 U7874 ( .A1(n8362), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n6270) );
  INV_X1 U7875 ( .A(n6273), .ZN(n6272) );
  INV_X1 U7876 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n8257) );
  NAND2_X1 U7877 ( .A1(n6272), .A2(n8257), .ZN(n8771) );
  NAND2_X1 U7878 ( .A1(n6273), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n6274) );
  NAND2_X1 U7879 ( .A1(n8771), .A2(n6274), .ZN(n8791) );
  NAND2_X1 U7880 ( .A1(n8791), .A2(n6216), .ZN(n6280) );
  INV_X1 U7881 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n8921) );
  NAND2_X1 U7882 ( .A1(n6359), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6276) );
  NAND2_X1 U7883 ( .A1(n5973), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n6275) );
  OAI211_X1 U7884 ( .C1(n8921), .C2(n6277), .A(n6276), .B(n6275), .ZN(n6278)
         );
  INV_X1 U7885 ( .A(n6278), .ZN(n6279) );
  NAND2_X1 U7886 ( .A1(n8985), .A2(n8551), .ZN(n8252) );
  NAND2_X1 U7887 ( .A1(n8785), .A2(n8252), .ZN(n6281) );
  NAND2_X1 U7888 ( .A1(n6281), .A2(n8253), .ZN(n8573) );
  NAND2_X1 U7889 ( .A1(n8185), .A2(n8365), .ZN(n6284) );
  NAND2_X1 U7890 ( .A1(n6282), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n6283) );
  INV_X1 U7891 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n8777) );
  NAND2_X1 U7892 ( .A1(n6359), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6287) );
  NAND2_X1 U7893 ( .A1(n5983), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6286) );
  OAI211_X1 U7894 ( .C1(n6067), .C2(n8777), .A(n6287), .B(n6286), .ZN(n6288)
         );
  INV_X1 U7895 ( .A(n6288), .ZN(n6289) );
  NAND2_X1 U7896 ( .A1(n8780), .A2(n8592), .ZN(n8371) );
  INV_X1 U7897 ( .A(n8782), .ZN(n6367) );
  INV_X1 U7898 ( .A(n4674), .ZN(n6291) );
  NAND2_X1 U7899 ( .A1(n6291), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6292) );
  XNOR2_X1 U7900 ( .A(n6292), .B(P2_IR_REG_20__SCAN_IN), .ZN(n6410) );
  INV_X1 U7901 ( .A(n6410), .ZN(n8568) );
  NAND2_X1 U7902 ( .A1(n6399), .A2(n8568), .ZN(n6940) );
  AND2_X1 U7903 ( .A1(n4674), .A2(n6293), .ZN(n6351) );
  NAND2_X1 U7904 ( .A1(n6351), .A2(n6294), .ZN(n6354) );
  NAND2_X1 U7905 ( .A1(n6354), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6295) );
  MUX2_X1 U7906 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6295), .S(
        P2_IR_REG_22__SCAN_IN), .Z(n6297) );
  NAND2_X1 U7907 ( .A1(n6297), .A2(n6296), .ZN(n7597) );
  INV_X1 U7908 ( .A(n7597), .ZN(n8588) );
  INV_X1 U7909 ( .A(n8991), .ZN(n6348) );
  INV_X1 U7910 ( .A(n8843), .ZN(n8873) );
  INV_X1 U7911 ( .A(n8972), .ZN(n6969) );
  NAND2_X1 U7912 ( .A1(n8610), .A2(n6969), .ZN(n6751) );
  NAND2_X1 U7913 ( .A1(n6298), .A2(n6751), .ZN(n6301) );
  NAND2_X1 U7914 ( .A1(n4438), .A2(n6859), .ZN(n6300) );
  NAND2_X1 U7915 ( .A1(n6301), .A2(n6300), .ZN(n6703) );
  NAND2_X1 U7916 ( .A1(n6703), .A2(n6704), .ZN(n6303) );
  INV_X1 U7917 ( .A(n8608), .ZN(n6754) );
  NAND2_X1 U7918 ( .A1(n6754), .A2(n8420), .ZN(n6302) );
  NOR2_X1 U7919 ( .A1(n8607), .A2(n7108), .ZN(n6304) );
  INV_X1 U7920 ( .A(n8607), .ZN(n6844) );
  OR2_X1 U7921 ( .A1(n8606), .A2(n10076), .ZN(n6305) );
  NAND2_X1 U7922 ( .A1(n7090), .A2(n6305), .ZN(n6307) );
  NAND2_X1 U7923 ( .A1(n8606), .A2(n10076), .ZN(n6306) );
  NAND2_X1 U7924 ( .A1(n6307), .A2(n6306), .ZN(n7216) );
  INV_X1 U7925 ( .A(n8605), .ZN(n7155) );
  NAND2_X1 U7926 ( .A1(n7155), .A2(n10083), .ZN(n6308) );
  NAND2_X1 U7927 ( .A1(n7216), .A2(n6308), .ZN(n6310) );
  NAND2_X1 U7928 ( .A1(n8605), .A2(n7212), .ZN(n6309) );
  NAND2_X1 U7929 ( .A1(n6310), .A2(n6309), .ZN(n7114) );
  OR2_X1 U7930 ( .A1(n8604), .A2(n7147), .ZN(n7113) );
  OR2_X1 U7931 ( .A1(n8603), .A2(n10094), .ZN(n6319) );
  AND2_X1 U7932 ( .A1(n7113), .A2(n6319), .ZN(n6311) );
  NAND2_X1 U7933 ( .A1(n7114), .A2(n6311), .ZN(n6315) );
  INV_X1 U7934 ( .A(n6319), .ZN(n6313) );
  NAND2_X1 U7935 ( .A1(n8604), .A2(n7147), .ZN(n7125) );
  NAND2_X1 U7936 ( .A1(n10094), .A2(n8603), .ZN(n6312) );
  AND2_X1 U7937 ( .A1(n7125), .A2(n6312), .ZN(n6317) );
  OR2_X1 U7938 ( .A1(n6313), .A2(n6317), .ZN(n6314) );
  NAND2_X1 U7939 ( .A1(n6315), .A2(n6314), .ZN(n7053) );
  NAND2_X1 U7940 ( .A1(n7053), .A2(n8602), .ZN(n6316) );
  INV_X1 U7941 ( .A(n7578), .ZN(n10102) );
  NAND2_X1 U7942 ( .A1(n6316), .A2(n10102), .ZN(n6323) );
  NAND2_X1 U7943 ( .A1(n7114), .A2(n7113), .ZN(n7126) );
  AND2_X1 U7944 ( .A1(n6317), .A2(n7474), .ZN(n6318) );
  NAND2_X1 U7945 ( .A1(n7126), .A2(n6318), .ZN(n6321) );
  OR2_X1 U7946 ( .A1(n8602), .A2(n6319), .ZN(n6320) );
  AND2_X1 U7947 ( .A1(n6321), .A2(n6320), .ZN(n6322) );
  NAND2_X1 U7948 ( .A1(n6323), .A2(n6322), .ZN(n7137) );
  NAND2_X1 U7949 ( .A1(n7137), .A2(n8387), .ZN(n6325) );
  OR2_X1 U7950 ( .A1(n7468), .A2(n8601), .ZN(n6324) );
  NOR2_X1 U7951 ( .A1(n7796), .A2(n8600), .ZN(n6326) );
  NAND2_X1 U7952 ( .A1(n7796), .A2(n8600), .ZN(n6327) );
  AND2_X1 U7953 ( .A1(n10124), .A2(n8599), .ZN(n6328) );
  NOR2_X1 U7954 ( .A1(n10131), .A2(n8598), .ZN(n7659) );
  INV_X1 U7955 ( .A(n6330), .ZN(n8492) );
  OR2_X1 U7956 ( .A1(n7659), .A2(n8492), .ZN(n6329) );
  NAND2_X1 U7957 ( .A1(n10131), .A2(n8598), .ZN(n7661) );
  NAND2_X1 U7958 ( .A1(n8488), .A2(n8597), .ZN(n8489) );
  NAND2_X1 U7959 ( .A1(n6330), .A2(n8489), .ZN(n8392) );
  INV_X1 U7960 ( .A(n8392), .ZN(n7665) );
  AND2_X1 U7961 ( .A1(n7661), .A2(n7665), .ZN(n7662) );
  NAND2_X1 U7962 ( .A1(n7909), .A2(n8596), .ZN(n6332) );
  NAND2_X1 U7963 ( .A1(n7651), .A2(n6332), .ZN(n6334) );
  OR2_X1 U7964 ( .A1(n7909), .A2(n8596), .ZN(n6333) );
  NAND2_X1 U7965 ( .A1(n7930), .A2(n8595), .ZN(n6336) );
  NAND2_X1 U7966 ( .A1(n8966), .A2(n8594), .ZN(n6337) );
  NAND2_X1 U7967 ( .A1(n8520), .A2(n8505), .ZN(n8516) );
  NAND2_X1 U7968 ( .A1(n8289), .A2(n8593), .ZN(n6338) );
  OR2_X1 U7969 ( .A1(n8959), .A2(n8897), .ZN(n6339) );
  INV_X1 U7970 ( .A(n8334), .ZN(n8883) );
  NAND2_X1 U7971 ( .A1(n8408), .A2(n8508), .ZN(n8881) );
  INV_X1 U7972 ( .A(n9032), .ZN(n6340) );
  NAND2_X1 U7973 ( .A1(n6340), .A2(n8268), .ZN(n8869) );
  NOR2_X1 U7974 ( .A1(n9026), .A2(n8884), .ZN(n8853) );
  NAND2_X1 U7975 ( .A1(n8535), .A2(n8531), .ZN(n8863) );
  OAI21_X1 U7976 ( .B1(n8868), .B2(n8853), .A(n8863), .ZN(n8852) );
  INV_X1 U7977 ( .A(n8859), .ZN(n8833) );
  NAND2_X1 U7978 ( .A1(n8238), .A2(n8833), .ZN(n6341) );
  INV_X1 U7979 ( .A(n9010), .ZN(n8836) );
  INV_X1 U7980 ( .A(n9004), .ZN(n8813) );
  OAI21_X1 U7981 ( .B1(n6346), .B2(n4658), .A(n6345), .ZN(n8795) );
  AOI21_X1 U7982 ( .B1(n8788), .B2(n8991), .A(n8795), .ZN(n6347) );
  INV_X1 U7983 ( .A(n8985), .ZN(n8550) );
  NAND2_X1 U7984 ( .A1(n8550), .A2(n8551), .ZN(n6349) );
  INV_X1 U7985 ( .A(n8551), .ZN(n8796) );
  AOI22_X1 U7986 ( .A1(n8787), .A2(n6349), .B1(n8985), .B2(n8796), .ZN(n6350)
         );
  XNOR2_X1 U7987 ( .A(n6350), .B(n8558), .ZN(n6366) );
  AND2_X1 U7988 ( .A1(n6399), .A2(n8588), .ZN(n6397) );
  INV_X1 U7989 ( .A(n6351), .ZN(n6352) );
  NAND2_X1 U7990 ( .A1(n6352), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6353) );
  MUX2_X1 U7991 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6353), .S(
        P2_IR_REG_21__SCAN_IN), .Z(n6355) );
  NAND2_X1 U7992 ( .A1(n6355), .A2(n6354), .ZN(n7534) );
  NOR2_X1 U7993 ( .A1(n7534), .A2(n8568), .ZN(n8578) );
  AND2_X1 U7994 ( .A1(n8760), .A2(n8568), .ZN(n6412) );
  NOR2_X1 U7995 ( .A1(n7597), .A2(n7534), .ZN(n8430) );
  AND2_X1 U7996 ( .A1(n6412), .A2(n8567), .ZN(n6741) );
  NAND2_X1 U7997 ( .A1(n7597), .A2(n7534), .ZN(n10114) );
  OAI21_X1 U7998 ( .B1(n8588), .B2(n8568), .A(n10114), .ZN(n6356) );
  OR3_X1 U7999 ( .A1(n6741), .A2(n6399), .A3(n6356), .ZN(n10107) );
  INV_X1 U8000 ( .A(n10107), .ZN(n7217) );
  OR2_X2 U8001 ( .A1(n6374), .A2(P2_IR_REG_26__SCAN_IN), .ZN(n6376) );
  NAND2_X1 U8002 ( .A1(n6376), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6357) );
  INV_X1 U8003 ( .A(n6489), .ZN(n8585) );
  NAND2_X1 U8004 ( .A1(n6568), .A2(n8585), .ZN(n6358) );
  NAND2_X1 U8005 ( .A1(n6358), .A2(n6443), .ZN(n6743) );
  NAND2_X1 U8006 ( .A1(n5973), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n6362) );
  NAND2_X1 U8007 ( .A1(n5983), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n6361) );
  NAND2_X1 U8008 ( .A1(n6359), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n6360) );
  AND3_X1 U8009 ( .A1(n6362), .A2(n6361), .A3(n6360), .ZN(n6363) );
  AND2_X1 U8010 ( .A1(n7410), .A2(n6363), .ZN(n8374) );
  NAND2_X1 U8011 ( .A1(n6743), .A2(n8567), .ZN(n8860) );
  AND2_X1 U8012 ( .A1(n6443), .A2(P2_B_REG_SCAN_IN), .ZN(n6364) );
  OR2_X1 U8013 ( .A1(n8860), .A2(n6364), .ZN(n8768) );
  OAI22_X1 U8014 ( .A1(n8551), .A2(n8858), .B1(n8374), .B2(n8768), .ZN(n6365)
         );
  OAI21_X1 U8015 ( .B1(n6367), .B2(n10116), .A(n8776), .ZN(n6423) );
  OR2_X1 U8016 ( .A1(n6369), .A2(n6368), .ZN(n6370) );
  NAND2_X1 U8017 ( .A1(n6371), .A2(n6370), .ZN(n7764) );
  NAND2_X1 U8018 ( .A1(n6371), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6373) );
  NAND2_X1 U8019 ( .A1(n6374), .A2(P2_IR_REG_26__SCAN_IN), .ZN(n6375) );
  AND2_X2 U8020 ( .A1(n6376), .A2(n6375), .ZN(n6391) );
  OR2_X1 U8021 ( .A1(n6461), .A2(P2_D_REG_1__SCAN_IN), .ZN(n6378) );
  INV_X1 U8022 ( .A(n6391), .ZN(n7873) );
  NAND2_X1 U8023 ( .A1(n7816), .A2(n7873), .ZN(n6377) );
  NAND2_X1 U8024 ( .A1(n6378), .A2(n6377), .ZN(n6931) );
  INV_X1 U8025 ( .A(n6931), .ZN(n9052) );
  NAND2_X1 U8026 ( .A1(n7873), .A2(n7764), .ZN(n6475) );
  AND2_X1 U8027 ( .A1(n9052), .A2(n6724), .ZN(n6409) );
  NOR2_X1 U8028 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .ZN(
        n6383) );
  NOR4_X1 U8029 ( .A1(P2_D_REG_5__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_23__SCAN_IN), .A4(P2_D_REG_4__SCAN_IN), .ZN(n6382) );
  NOR4_X1 U8030 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_16__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_27__SCAN_IN), .ZN(n6381) );
  NOR4_X1 U8031 ( .A1(P2_D_REG_20__SCAN_IN), .A2(P2_D_REG_29__SCAN_IN), .A3(
        P2_D_REG_30__SCAN_IN), .A4(P2_D_REG_22__SCAN_IN), .ZN(n6380) );
  NAND4_X1 U8032 ( .A1(n6383), .A2(n6382), .A3(n6381), .A4(n6380), .ZN(n6389)
         );
  NOR4_X1 U8033 ( .A1(P2_D_REG_9__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_14__SCAN_IN), .ZN(n6387) );
  NOR4_X1 U8034 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_24__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n6386) );
  NOR4_X1 U8035 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_6__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6385) );
  NOR4_X1 U8036 ( .A1(P2_D_REG_13__SCAN_IN), .A2(P2_D_REG_21__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_11__SCAN_IN), .ZN(n6384) );
  NAND4_X1 U8037 ( .A1(n6387), .A2(n6386), .A3(n6385), .A4(n6384), .ZN(n6388)
         );
  NOR2_X1 U8038 ( .A1(n6389), .A2(n6388), .ZN(n6390) );
  OR2_X1 U8039 ( .A1(n6461), .A2(n6390), .ZN(n6414) );
  NAND2_X1 U8040 ( .A1(n6409), .A2(n6414), .ZN(n6714) );
  INV_X1 U8041 ( .A(n6714), .ZN(n6396) );
  INV_X1 U8042 ( .A(n7816), .ZN(n6393) );
  INV_X1 U8043 ( .A(n7764), .ZN(n6392) );
  NAND3_X1 U8044 ( .A1(n6393), .A2(n6392), .A3(n6391), .ZN(n6715) );
  NAND2_X1 U8045 ( .A1(n6296), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6395) );
  XNOR2_X1 U8046 ( .A(n6395), .B(n6394), .ZN(n7647) );
  AND2_X1 U8047 ( .A1(n7647), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6477) );
  NAND2_X1 U8048 ( .A1(n6715), .A2(n6477), .ZN(n9051) );
  INV_X1 U8049 ( .A(n9051), .ZN(n6738) );
  AND2_X1 U8050 ( .A1(n6396), .A2(n6738), .ZN(n6737) );
  AND2_X1 U8051 ( .A1(n7534), .A2(n6410), .ZN(n8378) );
  AND2_X1 U8052 ( .A1(n6397), .A2(n8378), .ZN(n6732) );
  OR2_X1 U8053 ( .A1(n6741), .A2(n6732), .ZN(n6398) );
  NAND2_X1 U8054 ( .A1(n6737), .A2(n6398), .ZN(n6403) );
  INV_X1 U8055 ( .A(n6724), .ZN(n6932) );
  NAND3_X1 U8056 ( .A1(n6931), .A2(n6932), .A3(n6414), .ZN(n6721) );
  NOR2_X1 U8057 ( .A1(n6721), .A2(n9051), .ZN(n6742) );
  INV_X1 U8058 ( .A(n10114), .ZN(n10132) );
  NAND2_X1 U8059 ( .A1(n6940), .A2(n10132), .ZN(n8835) );
  NAND2_X1 U8060 ( .A1(n6399), .A2(n8378), .ZN(n6401) );
  NOR2_X1 U8061 ( .A1(n8567), .A2(n10132), .ZN(n6400) );
  NAND2_X1 U8062 ( .A1(n6401), .A2(n6400), .ZN(n6730) );
  NAND2_X1 U8063 ( .A1(n8835), .A2(n6730), .ZN(n6713) );
  NAND2_X1 U8064 ( .A1(n6742), .A2(n6713), .ZN(n6402) );
  INV_X2 U8065 ( .A(n10135), .ZN(n10133) );
  NAND2_X1 U8066 ( .A1(n6423), .A2(n10133), .ZN(n6408) );
  INV_X1 U8067 ( .A(n8780), .ZN(n6405) );
  OR2_X1 U8068 ( .A1(n10135), .A2(n10114), .ZN(n9044) );
  OAI22_X1 U8069 ( .A1(n6405), .A2(n9044), .B1(n10133), .B2(n6404), .ZN(n6406)
         );
  NAND2_X1 U8070 ( .A1(n6408), .A2(n6407), .ZN(P2_U3456) );
  INV_X1 U8071 ( .A(n6409), .ZN(n6420) );
  NAND3_X1 U8072 ( .A1(n8760), .A2(n8588), .A3(n6410), .ZN(n6411) );
  NAND2_X1 U8073 ( .A1(n6411), .A2(n8552), .ZN(n6935) );
  AND2_X1 U8074 ( .A1(n6931), .A2(n6935), .ZN(n6415) );
  INV_X1 U8075 ( .A(n6412), .ZN(n6413) );
  NAND2_X1 U8076 ( .A1(n6413), .A2(n8567), .ZN(n6716) );
  NAND3_X1 U8077 ( .A1(n6738), .A2(n6414), .A3(n6716), .ZN(n6933) );
  NOR2_X1 U8078 ( .A1(n6415), .A2(n6933), .ZN(n6419) );
  INV_X1 U8079 ( .A(n7534), .ZN(n8426) );
  NOR2_X1 U8080 ( .A1(n10116), .A2(n8426), .ZN(n6739) );
  INV_X1 U8081 ( .A(n6739), .ZN(n6416) );
  NAND2_X1 U8082 ( .A1(n6416), .A2(n6724), .ZN(n6417) );
  INV_X1 U8083 ( .A(n6935), .ZN(n6934) );
  NAND2_X1 U8084 ( .A1(n6417), .A2(n6934), .ZN(n6418) );
  AND3_X2 U8085 ( .A1(n6420), .A2(n6419), .A3(n6418), .ZN(n10152) );
  NAND2_X1 U8086 ( .A1(n10150), .A2(n6421), .ZN(n6422) );
  NAND2_X1 U8087 ( .A1(n8780), .A2(n8948), .ZN(n6424) );
  NAND2_X1 U8088 ( .A1(n6425), .A2(n6424), .ZN(P2_U3488) );
  NAND2_X1 U8089 ( .A1(n9063), .A2(n9865), .ZN(n6437) );
  INV_X1 U8090 ( .A(n9291), .ZN(n9106) );
  OAI22_X1 U8091 ( .A1(n6431), .A2(n9096), .B1(n6430), .B2(n9106), .ZN(n9591)
         );
  OAI22_X1 U8092 ( .A1(n9598), .A2(n9868), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6432), .ZN(n6433) );
  AOI21_X1 U8093 ( .B1(n9591), .B2(n9861), .A(n6433), .ZN(n6434) );
  OAI21_X1 U8094 ( .B1(n6438), .B2(n6437), .A(n6436), .ZN(P1_U3240) );
  NOR2_X1 U8095 ( .A1(n6439), .A2(P1_U3086), .ZN(n6440) );
  INV_X1 U8096 ( .A(n6477), .ZN(n6441) );
  OR2_X2 U8097 ( .A1(n6715), .A2(n6441), .ZN(n8719) );
  INV_X1 U8098 ( .A(n8719), .ZN(P2_U3893) );
  NAND2_X1 U8099 ( .A1(n6715), .A2(n8552), .ZN(n6442) );
  NAND2_X1 U8100 ( .A1(n6442), .A2(n7647), .ZN(n6490) );
  NAND2_X1 U8101 ( .A1(n6490), .A2(n6443), .ZN(n6444) );
  NAND2_X1 U8102 ( .A1(n6444), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  NOR2_X1 U8103 ( .A1(n8358), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9056) );
  NAND2_X1 U8104 ( .A1(n8358), .A2(P2_U3151), .ZN(n9058) );
  CLKBUF_X1 U8105 ( .A(n9058), .Z(n8159) );
  OAI222_X1 U8106 ( .A1(n8186), .A2(n6445), .B1(n8159), .B2(n6452), .C1(
        P2_U3151), .C2(n6540), .ZN(P2_U3294) );
  OAI222_X1 U8107 ( .A1(n8186), .A2(n6446), .B1(n8159), .B2(n6450), .C1(
        P2_U3151), .C2(n6583), .ZN(P2_U3293) );
  AOI22_X1 U8108 ( .A1(n6448), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(
        P1_STATE_REG_SCAN_IN), .B2(n9891), .ZN(n6449) );
  OAI21_X1 U8109 ( .B1(n6450), .B2(n7965), .A(n6449), .ZN(P1_U3353) );
  INV_X1 U8110 ( .A(n6448), .ZN(n8191) );
  OAI222_X1 U8111 ( .A1(n6637), .A2(P1_U3086), .B1(n7965), .B2(n6452), .C1(
        n6451), .C2(n8191), .ZN(P1_U3354) );
  OAI222_X1 U8112 ( .A1(n8186), .A2(n6453), .B1(n9058), .B2(n8184), .C1(
        P2_U3151), .C2(n6586), .ZN(P2_U3292) );
  INV_X1 U8113 ( .A(n6774), .ZN(n6765) );
  OAI222_X1 U8114 ( .A1(n8186), .A2(n6454), .B1(n9058), .B2(n6456), .C1(
        P2_U3151), .C2(n6765), .ZN(P2_U3291) );
  OAI222_X1 U8115 ( .A1(n6457), .A2(P1_U3086), .B1(n7965), .B2(n6456), .C1(
        n6455), .C2(n8191), .ZN(P1_U3351) );
  AOI22_X1 U8116 ( .A1(n6658), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n6448), .ZN(n6458) );
  OAI21_X1 U8117 ( .B1(n6459), .B2(n7965), .A(n6458), .ZN(P1_U3350) );
  OAI222_X1 U8118 ( .A1(n8186), .A2(n6460), .B1(n8159), .B2(n6459), .C1(
        P2_U3151), .C2(n6777), .ZN(P2_U3290) );
  AND2_X1 U8119 ( .A1(n6461), .A2(n6738), .ZN(n6474) );
  INV_X1 U8120 ( .A(P2_D_REG_4__SCAN_IN), .ZN(n7982) );
  NOR2_X1 U8121 ( .A1(n6474), .A2(n7982), .ZN(P2_U3261) );
  INV_X1 U8122 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n6462) );
  NOR2_X1 U8123 ( .A1(n6474), .A2(n6462), .ZN(P2_U3248) );
  INV_X1 U8124 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n7983) );
  NOR2_X1 U8125 ( .A1(n6474), .A2(n7983), .ZN(P2_U3242) );
  INV_X1 U8126 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n7995) );
  NOR2_X1 U8127 ( .A1(n6474), .A2(n7995), .ZN(P2_U3258) );
  INV_X1 U8128 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n8096) );
  NOR2_X1 U8129 ( .A1(n6474), .A2(n8096), .ZN(P2_U3245) );
  INV_X1 U8130 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6464) );
  INV_X1 U8131 ( .A(n6463), .ZN(n6466) );
  OAI222_X1 U8132 ( .A1(n8186), .A2(n6464), .B1(n8159), .B2(n6466), .C1(
        P2_U3151), .C2(n6908), .ZN(P2_U3289) );
  INV_X1 U8133 ( .A(n6669), .ZN(n6627) );
  INV_X1 U8134 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6465) );
  OAI222_X1 U8135 ( .A1(n6627), .A2(P1_U3086), .B1(n7965), .B2(n6466), .C1(
        n6465), .C2(n8191), .ZN(P1_U3349) );
  INV_X1 U8136 ( .A(n6474), .ZN(n6467) );
  AND2_X1 U8137 ( .A1(n6467), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U8138 ( .A1(n6467), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U8139 ( .A1(n6467), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U8140 ( .A1(n6467), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  AND2_X1 U8141 ( .A1(n6467), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U8142 ( .A1(n6467), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U8143 ( .A1(n6467), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U8144 ( .A1(n6467), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  INV_X1 U8145 ( .A(n6798), .ZN(n6469) );
  INV_X1 U8146 ( .A(n6468), .ZN(n6470) );
  INV_X1 U8147 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n8142) );
  OAI222_X1 U8148 ( .A1(n6469), .A2(P1_U3086), .B1(n7965), .B2(n6470), .C1(
        n8142), .C2(n8191), .ZN(P1_U3348) );
  INV_X1 U8149 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6471) );
  OAI222_X1 U8150 ( .A1(n8186), .A2(n6471), .B1(n8159), .B2(n6470), .C1(
        P2_U3151), .C2(n4604), .ZN(P2_U3288) );
  INV_X1 U8151 ( .A(n6472), .ZN(n6478) );
  AOI22_X1 U8152 ( .A1(n6886), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n6448), .ZN(n6473) );
  OAI21_X1 U8153 ( .B1(n6478), .B2(n7965), .A(n6473), .ZN(P1_U3347) );
  AND2_X1 U8154 ( .A1(n6467), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3255) );
  AND2_X1 U8155 ( .A1(n6467), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  AND2_X1 U8156 ( .A1(n6467), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U8157 ( .A1(n6467), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  AND2_X1 U8158 ( .A1(n6467), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U8159 ( .A1(n6467), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U8160 ( .A1(n6467), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U8161 ( .A1(n6467), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3262) );
  AND2_X1 U8162 ( .A1(n6467), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  AND2_X1 U8163 ( .A1(n6467), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U8164 ( .A1(n6467), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U8165 ( .A1(n6467), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U8166 ( .A1(n6467), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  AND2_X1 U8167 ( .A1(n6467), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U8168 ( .A1(n6467), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  AND2_X1 U8169 ( .A1(n6467), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U8170 ( .A1(n6467), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  INV_X1 U8171 ( .A(n6475), .ZN(n6476) );
  AOI22_X1 U8172 ( .A1(n6467), .A2(n4868), .B1(n6477), .B2(n6476), .ZN(
        P2_U3376) );
  INV_X1 U8173 ( .A(n8619), .ZN(n7004) );
  OAI222_X1 U8174 ( .A1(n8186), .A2(n6479), .B1(n8159), .B2(n6478), .C1(
        P2_U3151), .C2(n7004), .ZN(P2_U3287) );
  INV_X1 U8175 ( .A(n6480), .ZN(n6483) );
  AOI22_X1 U8176 ( .A1(n7266), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n6448), .ZN(n6481) );
  OAI21_X1 U8177 ( .B1(n6483), .B2(n7965), .A(n6481), .ZN(P1_U3345) );
  INV_X1 U8178 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6482) );
  OAI222_X1 U8179 ( .A1(n8159), .A2(n6483), .B1(n7395), .B2(P2_U3151), .C1(
        n6482), .C2(n8186), .ZN(P2_U3285) );
  INV_X1 U8180 ( .A(n6484), .ZN(n6499) );
  AOI22_X1 U8181 ( .A1(n7022), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n6448), .ZN(n6485) );
  OAI21_X1 U8182 ( .B1(n6499), .B2(n7965), .A(n6485), .ZN(P1_U3346) );
  AND2_X1 U8183 ( .A1(n6568), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7923) );
  NAND2_X1 U8184 ( .A1(n6490), .A2(n7923), .ZN(n6486) );
  MUX2_X1 U8185 ( .A(n6486), .B(n8719), .S(n8585), .Z(n8761) );
  INV_X1 U8186 ( .A(n7647), .ZN(n6487) );
  NOR2_X1 U8187 ( .A1(n6715), .A2(n6487), .ZN(n6488) );
  OR2_X1 U8188 ( .A1(P2_U3150), .A2(n6488), .ZN(n8724) );
  INV_X1 U8189 ( .A(n8724), .ZN(n8757) );
  AOI22_X1 U8190 ( .A1(n8757), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3151), .ZN(n6497) );
  NOR2_X1 U8191 ( .A1(n6489), .A2(P2_U3151), .ZN(n7966) );
  NAND2_X1 U8192 ( .A1(n6490), .A2(n7966), .ZN(n6517) );
  INV_X1 U8193 ( .A(n6517), .ZN(n6495) );
  NOR2_X2 U8194 ( .A1(n8719), .A2(n8585), .ZN(n8763) );
  INV_X1 U8195 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n6492) );
  INV_X1 U8196 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6491) );
  MUX2_X1 U8197 ( .A(n6492), .B(n6491), .S(n6568), .Z(n6493) );
  NAND2_X1 U8198 ( .A1(n6493), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6542) );
  OAI21_X1 U8199 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n6493), .A(n6542), .ZN(n6494) );
  OAI21_X1 U8200 ( .B1(n6495), .B2(n8763), .A(n6494), .ZN(n6496) );
  OAI211_X1 U8201 ( .C1(n8761), .C2(n6513), .A(n6497), .B(n6496), .ZN(P2_U3182) );
  INV_X1 U8202 ( .A(n7076), .ZN(n7005) );
  OAI222_X1 U8203 ( .A1(n8159), .A2(n6499), .B1(n7005), .B2(P2_U3151), .C1(
        n6498), .C2(n8186), .ZN(P2_U3286) );
  INV_X1 U8204 ( .A(n6500), .ZN(n6523) );
  AOI22_X1 U8205 ( .A1(n7346), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n6448), .ZN(n6501) );
  OAI21_X1 U8206 ( .B1(n6523), .B2(n7965), .A(n6501), .ZN(P1_U3344) );
  NAND2_X1 U8207 ( .A1(n7645), .A2(n6502), .ZN(n6503) );
  NAND2_X1 U8208 ( .A1(n6503), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6632) );
  INV_X1 U8209 ( .A(n6632), .ZN(n6506) );
  NAND2_X1 U8210 ( .A1(n6504), .A2(n7645), .ZN(n6505) );
  NAND2_X1 U8211 ( .A1(n6505), .A2(n5013), .ZN(n6633) );
  NAND2_X1 U8212 ( .A1(n6506), .A2(n6633), .ZN(n9553) );
  INV_X1 U8213 ( .A(n9553), .ZN(n9933) );
  NOR2_X1 U8214 ( .A1(n9933), .A2(P1_U3973), .ZN(P1_U3085) );
  MUX2_X1 U8215 ( .A(P2_REG1_REG_1__SCAN_IN), .B(P2_REG2_REG_1__SCAN_IN), .S(
        n4333), .Z(n6541) );
  XOR2_X1 U8216 ( .A(n6540), .B(n6541), .Z(n6543) );
  XOR2_X1 U8217 ( .A(n6542), .B(n6543), .Z(n6507) );
  NAND2_X1 U8218 ( .A1(n6507), .A2(n8763), .ZN(n6522) );
  OR2_X1 U8219 ( .A1(n6517), .A2(n8584), .ZN(n8756) );
  AND2_X1 U8220 ( .A1(n6513), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6508) );
  NAND2_X1 U8221 ( .A1(n5968), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6552) );
  OAI21_X1 U8222 ( .B1(n6509), .B2(n6508), .A(n6552), .ZN(n6510) );
  INV_X1 U8223 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n8013) );
  OR2_X1 U8224 ( .A1(n6510), .A2(n8013), .ZN(n6553) );
  NAND2_X1 U8225 ( .A1(n6510), .A2(n8013), .ZN(n6511) );
  AND2_X1 U8226 ( .A1(n6553), .A2(n6511), .ZN(n6512) );
  OAI22_X1 U8227 ( .A1(n8756), .A2(n6512), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n4641), .ZN(n6520) );
  AND2_X1 U8228 ( .A1(n6513), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6514) );
  NAND2_X1 U8229 ( .A1(n5968), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6545) );
  OAI21_X1 U8230 ( .B1(n6540), .B2(n6514), .A(n6545), .ZN(n6516) );
  INV_X1 U8231 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6515) );
  OR2_X1 U8232 ( .A1(n6516), .A2(n6515), .ZN(n6546) );
  NAND2_X1 U8233 ( .A1(n6516), .A2(n6515), .ZN(n6518) );
  OR2_X1 U8234 ( .A1(n6517), .A2(n6568), .ZN(n8766) );
  AOI21_X1 U8235 ( .B1(n6546), .B2(n6518), .A(n8766), .ZN(n6519) );
  AOI211_X1 U8236 ( .C1(n8757), .C2(P2_ADDR_REG_1__SCAN_IN), .A(n6520), .B(
        n6519), .ZN(n6521) );
  OAI211_X1 U8237 ( .C1(n8761), .C2(n6540), .A(n6522), .B(n6521), .ZN(P2_U3183) );
  OAI222_X1 U8238 ( .A1(n8186), .A2(n6524), .B1(n8159), .B2(n6523), .C1(
        P2_U3151), .C2(n7398), .ZN(P2_U3284) );
  NAND2_X1 U8239 ( .A1(n6695), .A2(P1_U3973), .ZN(n6525) );
  OAI21_X1 U8240 ( .B1(P1_U3973), .B2(n5961), .A(n6525), .ZN(P1_U3554) );
  INV_X1 U8241 ( .A(n6526), .ZN(n6529) );
  INV_X1 U8242 ( .A(n7528), .ZN(n7507) );
  OAI222_X1 U8243 ( .A1(n8159), .A2(n6529), .B1(n7507), .B2(P2_U3151), .C1(
        n6527), .C2(n8186), .ZN(P2_U3283) );
  INV_X1 U8244 ( .A(n7585), .ZN(n7355) );
  OAI222_X1 U8245 ( .A1(P1_U3086), .A2(n7355), .B1(n7965), .B2(n6529), .C1(
        n6528), .C2(n8191), .ZN(P1_U3343) );
  INV_X1 U8246 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6535) );
  INV_X1 U8247 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n6533) );
  NAND2_X1 U8248 ( .A1(n6530), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n6532) );
  INV_X1 U8249 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n9804) );
  OR2_X1 U8250 ( .A1(n4982), .A2(n9804), .ZN(n6531) );
  OAI211_X1 U8251 ( .C1(n4980), .C2(n6533), .A(n6532), .B(n6531), .ZN(n9425)
         );
  NAND2_X1 U8252 ( .A1(P1_U3973), .A2(n9425), .ZN(n6534) );
  OAI21_X1 U8253 ( .B1(P1_U3973), .B2(n6535), .A(n6534), .ZN(P1_U3585) );
  INV_X1 U8254 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7357) );
  NAND2_X1 U8255 ( .A1(n6536), .A2(P1_U3973), .ZN(n6537) );
  OAI21_X1 U8256 ( .B1(n7357), .B2(P1_U3973), .A(n6537), .ZN(P1_U3574) );
  INV_X1 U8257 ( .A(n6538), .ZN(n6622) );
  AOI22_X1 U8258 ( .A1(n7682), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n6448), .ZN(n6539) );
  OAI21_X1 U8259 ( .B1(n6622), .B2(n7965), .A(n6539), .ZN(P1_U3342) );
  MUX2_X1 U8260 ( .A(P2_REG1_REG_2__SCAN_IN), .B(P2_REG2_REG_2__SCAN_IN), .S(
        n6568), .Z(n6562) );
  XNOR2_X1 U8261 ( .A(n6562), .B(n6583), .ZN(n6565) );
  AOI22_X1 U8262 ( .A1(n6543), .A2(n6542), .B1(n6541), .B2(n6540), .ZN(n6566)
         );
  XOR2_X1 U8263 ( .A(n6565), .B(n6566), .Z(n6560) );
  INV_X1 U8264 ( .A(n8766), .ZN(n8735) );
  INV_X1 U8265 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6544) );
  MUX2_X1 U8266 ( .A(n6544), .B(P2_REG1_REG_2__SCAN_IN), .S(n6564), .Z(n6548)
         );
  NAND2_X1 U8267 ( .A1(n6546), .A2(n6545), .ZN(n6547) );
  NAND2_X1 U8268 ( .A1(n6548), .A2(n6547), .ZN(n6585) );
  OAI21_X1 U8269 ( .B1(n6548), .B2(n6547), .A(n6585), .ZN(n6549) );
  AOI22_X1 U8270 ( .A1(n8757), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(n8735), .B2(
        n6549), .ZN(n6558) );
  INV_X1 U8271 ( .A(n8756), .ZN(n8631) );
  INV_X1 U8272 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6550) );
  NAND2_X1 U8273 ( .A1(n6553), .A2(n6552), .ZN(n6554) );
  NAND2_X1 U8274 ( .A1(n6555), .A2(n6554), .ZN(n6574) );
  OAI21_X1 U8275 ( .B1(n6555), .B2(n6554), .A(n6574), .ZN(n6556) );
  INV_X1 U8276 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n8139) );
  AOI22_X1 U8277 ( .A1(n8631), .A2(n6556), .B1(P2_U3151), .B2(
        P2_REG3_REG_2__SCAN_IN), .ZN(n6557) );
  OAI211_X1 U8278 ( .C1(n6583), .C2(n8761), .A(n6558), .B(n6557), .ZN(n6559)
         );
  AOI21_X1 U8279 ( .B1(n6560), .B2(n8763), .A(n6559), .ZN(n6561) );
  INV_X1 U8280 ( .A(n6561), .ZN(P2_U3184) );
  INV_X1 U8281 ( .A(n6562), .ZN(n6563) );
  OAI22_X1 U8282 ( .A1(n6566), .A2(n6565), .B1(n6564), .B2(n6563), .ZN(n6597)
         );
  MUX2_X1 U8283 ( .A(P2_REG1_REG_3__SCAN_IN), .B(P2_REG2_REG_3__SCAN_IN), .S(
        n6568), .Z(n6567) );
  XOR2_X1 U8284 ( .A(n6611), .B(n6567), .Z(n6598) );
  NOR2_X1 U8285 ( .A1(n6597), .A2(n6598), .ZN(n6596) );
  NOR2_X1 U8286 ( .A1(n6567), .A2(n6586), .ZN(n6570) );
  MUX2_X1 U8287 ( .A(P2_REG1_REG_4__SCAN_IN), .B(P2_REG2_REG_4__SCAN_IN), .S(
        n8748), .Z(n6766) );
  XNOR2_X1 U8288 ( .A(n6766), .B(n6765), .ZN(n6569) );
  NOR3_X1 U8289 ( .A1(n6596), .A2(n6570), .A3(n6569), .ZN(n6764) );
  INV_X1 U8290 ( .A(n6764), .ZN(n6572) );
  OAI21_X1 U8291 ( .B1(n6596), .B2(n6570), .A(n6569), .ZN(n6571) );
  NAND3_X1 U8292 ( .A1(n6572), .A2(n8763), .A3(n6571), .ZN(n6595) );
  NAND2_X1 U8293 ( .A1(n6583), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6573) );
  NAND2_X1 U8294 ( .A1(n6574), .A2(n6573), .ZN(n6576) );
  INV_X1 U8295 ( .A(n6577), .ZN(n6575) );
  INV_X1 U8296 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n7099) );
  MUX2_X1 U8297 ( .A(n7099), .B(P2_REG2_REG_4__SCAN_IN), .S(n6774), .Z(n6578)
         );
  NOR2_X1 U8298 ( .A1(n6575), .A2(n6578), .ZN(n6581) );
  INV_X1 U8299 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n7110) );
  OR2_X2 U8300 ( .A1(n6601), .A2(n7110), .ZN(n6599) );
  NAND2_X1 U8301 ( .A1(n6599), .A2(n6577), .ZN(n6579) );
  INV_X1 U8302 ( .A(n6776), .ZN(n6580) );
  AOI21_X1 U8303 ( .B1(n6581), .B2(n6599), .A(n6580), .ZN(n6582) );
  NAND2_X1 U8304 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3151), .ZN(n6847) );
  OAI21_X1 U8305 ( .B1(n8756), .B2(n6582), .A(n6847), .ZN(n6593) );
  NAND2_X1 U8306 ( .A1(n6583), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6584) );
  NAND2_X1 U8307 ( .A1(n6585), .A2(n6584), .ZN(n6587) );
  NAND2_X1 U8308 ( .A1(n6587), .A2(n6586), .ZN(n6589) );
  INV_X1 U8309 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10136) );
  INV_X1 U8310 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10138) );
  MUX2_X1 U8311 ( .A(n10138), .B(P2_REG1_REG_4__SCAN_IN), .S(n6774), .Z(n6588)
         );
  INV_X1 U8312 ( .A(n6588), .ZN(n6590) );
  NAND3_X1 U8313 ( .A1(n6604), .A2(n6590), .A3(n6589), .ZN(n6591) );
  AOI21_X1 U8314 ( .B1(n6768), .B2(n6591), .A(n8766), .ZN(n6592) );
  AOI211_X1 U8315 ( .C1(n8757), .C2(P2_ADDR_REG_4__SCAN_IN), .A(n6593), .B(
        n6592), .ZN(n6594) );
  OAI211_X1 U8316 ( .C1(n8761), .C2(n6765), .A(n6595), .B(n6594), .ZN(P2_U3186) );
  AOI21_X1 U8317 ( .B1(n6598), .B2(n6597), .A(n6596), .ZN(n6613) );
  INV_X1 U8318 ( .A(n8763), .ZN(n8695) );
  INV_X1 U8319 ( .A(n8761), .ZN(n8699) );
  INV_X1 U8320 ( .A(n6599), .ZN(n6600) );
  AOI21_X1 U8321 ( .B1(n7110), .B2(n6601), .A(n6600), .ZN(n6603) );
  NOR2_X1 U8322 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5985), .ZN(n6747) );
  INV_X1 U8323 ( .A(n6747), .ZN(n6602) );
  OAI21_X1 U8324 ( .B1(n8756), .B2(n6603), .A(n6602), .ZN(n6610) );
  INV_X1 U8325 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n6608) );
  INV_X1 U8326 ( .A(n6604), .ZN(n6605) );
  AOI21_X1 U8327 ( .B1(n10136), .B2(n6606), .A(n6605), .ZN(n6607) );
  OAI22_X1 U8328 ( .A1(n8724), .A2(n6608), .B1(n8766), .B2(n6607), .ZN(n6609)
         );
  AOI211_X1 U8329 ( .C1(n6611), .C2(n8699), .A(n6610), .B(n6609), .ZN(n6612)
         );
  OAI21_X1 U8330 ( .B1(n6613), .B2(n8695), .A(n6612), .ZN(P2_U3185) );
  INV_X1 U8331 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7414) );
  NAND2_X1 U8332 ( .A1(n8900), .A2(P2_U3893), .ZN(n6614) );
  OAI21_X1 U8333 ( .B1(P2_U3893), .B2(n7414), .A(n6614), .ZN(P2_U3511) );
  XNOR2_X1 U8334 ( .A(n6615), .B(n6616), .ZN(n9898) );
  INV_X1 U8335 ( .A(n9292), .ZN(n6617) );
  NAND2_X1 U8336 ( .A1(n6618), .A2(n6617), .ZN(n6839) );
  AOI22_X1 U8337 ( .A1(n9186), .A2(n7182), .B1(n6839), .B2(
        P1_REG3_REG_0__SCAN_IN), .ZN(n6621) );
  NAND2_X1 U8338 ( .A1(n9469), .A2(n9169), .ZN(n7184) );
  INV_X1 U8339 ( .A(n7184), .ZN(n6619) );
  NAND2_X1 U8340 ( .A1(n9861), .A2(n6619), .ZN(n6620) );
  OAI211_X1 U8341 ( .C1(n9898), .C2(n9188), .A(n6621), .B(n6620), .ZN(P1_U3232) );
  INV_X1 U8342 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6623) );
  INV_X1 U8343 ( .A(n7751), .ZN(n7616) );
  OAI222_X1 U8344 ( .A1(n8186), .A2(n6623), .B1(n8159), .B2(n6622), .C1(
        P2_U3151), .C2(n7616), .ZN(P2_U3282) );
  INV_X1 U8345 ( .A(n7182), .ZN(n7047) );
  NAND2_X1 U8346 ( .A1(n6695), .A2(n7047), .ZN(n9332) );
  NAND2_X1 U8347 ( .A1(n7037), .A2(n9332), .ZN(n9379) );
  OAI21_X1 U8348 ( .B1(n10029), .B2(n9698), .A(n9379), .ZN(n6624) );
  OAI211_X1 U8349 ( .C1(n6625), .C2(n7047), .A(n6624), .B(n7184), .ZN(n9802)
         );
  NAND2_X1 U8350 ( .A1(n10049), .A2(n9802), .ZN(n6626) );
  OAI21_X1 U8351 ( .B1(n10049), .B2(n4852), .A(n6626), .ZN(P1_U3453) );
  AOI22_X1 U8352 ( .A1(n6669), .A2(n5057), .B1(P1_REG2_REG_6__SCAN_IN), .B2(
        n6627), .ZN(n6636) );
  MUX2_X1 U8353 ( .A(n4933), .B(P1_REG2_REG_1__SCAN_IN), .S(n6637), .Z(n9478)
         );
  AND2_X1 U8354 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n9897) );
  NAND2_X1 U8355 ( .A1(n9478), .A2(n9897), .ZN(n9477) );
  INV_X1 U8356 ( .A(n6637), .ZN(n9473) );
  NAND2_X1 U8357 ( .A1(n9473), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6628) );
  NAND2_X1 U8358 ( .A1(n9477), .A2(n6628), .ZN(n9889) );
  NAND2_X1 U8359 ( .A1(n8182), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6629) );
  OAI21_X1 U8360 ( .B1(n8182), .B2(P1_REG2_REG_3__SCAN_IN), .A(n6629), .ZN(
        n6681) );
  NAND2_X1 U8361 ( .A1(P1_REG2_REG_4__SCAN_IN), .A2(n9910), .ZN(n6630) );
  OAI21_X1 U8362 ( .B1(P1_REG2_REG_4__SCAN_IN), .B2(n9910), .A(n6630), .ZN(
        n9913) );
  NOR2_X1 U8363 ( .A1(n9912), .A2(n9913), .ZN(n9911) );
  NAND2_X1 U8364 ( .A1(n6658), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6631) );
  OAI21_X1 U8365 ( .B1(n6658), .B2(P1_REG2_REG_5__SCAN_IN), .A(n6631), .ZN(
        n6654) );
  NOR2_X1 U8366 ( .A1(n6653), .A2(n6654), .ZN(n6652) );
  NOR2_X1 U8367 ( .A1(n6635), .A2(n6636), .ZN(n6664) );
  OR2_X1 U8368 ( .A1(n6633), .A2(n6632), .ZN(n9881) );
  INV_X1 U8369 ( .A(n5654), .ZN(n9896) );
  NAND2_X1 U8370 ( .A1(n9899), .A2(n9896), .ZN(n6634) );
  NOR2_X1 U8371 ( .A1(n9881), .A2(n6634), .ZN(n9915) );
  INV_X1 U8372 ( .A(n9915), .ZN(n9928) );
  AOI211_X1 U8373 ( .C1(n6636), .C2(n6635), .A(n6664), .B(n9928), .ZN(n6651)
         );
  INV_X1 U8374 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10050) );
  AND2_X1 U8375 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n9475) );
  NAND2_X1 U8376 ( .A1(n9473), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6638) );
  NAND2_X1 U8377 ( .A1(n9474), .A2(n6638), .ZN(n9885) );
  INV_X1 U8378 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6639) );
  MUX2_X1 U8379 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n6639), .S(n9891), .Z(n9886)
         );
  NAND2_X1 U8380 ( .A1(n9885), .A2(n9886), .ZN(n9884) );
  NAND2_X1 U8381 ( .A1(n8182), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6640) );
  OAI21_X1 U8382 ( .B1(n8182), .B2(P1_REG1_REG_3__SCAN_IN), .A(n6640), .ZN(
        n6683) );
  NAND2_X1 U8383 ( .A1(P1_REG1_REG_4__SCAN_IN), .A2(n9910), .ZN(n6641) );
  OAI21_X1 U8384 ( .B1(n9910), .B2(P1_REG1_REG_4__SCAN_IN), .A(n6641), .ZN(
        n9906) );
  NOR2_X1 U8385 ( .A1(n9905), .A2(n9906), .ZN(n9907) );
  NAND2_X1 U8386 ( .A1(n6658), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6642) );
  OAI21_X1 U8387 ( .B1(n6658), .B2(P1_REG1_REG_5__SCAN_IN), .A(n6642), .ZN(
        n6656) );
  NAND2_X1 U8388 ( .A1(n6669), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6643) );
  OAI21_X1 U8389 ( .B1(n6669), .B2(P1_REG1_REG_6__SCAN_IN), .A(n6643), .ZN(
        n6645) );
  INV_X1 U8390 ( .A(n9881), .ZN(n6644) );
  NAND2_X1 U8391 ( .A1(n6644), .A2(n5654), .ZN(n9919) );
  AOI211_X1 U8392 ( .C1(n6646), .C2(n6645), .A(n6668), .B(n9919), .ZN(n6650)
         );
  INV_X1 U8393 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n6648) );
  NOR2_X2 U8394 ( .A1(n9881), .A2(n9899), .ZN(n9937) );
  NAND2_X1 U8395 ( .A1(n9937), .A2(n6669), .ZN(n6647) );
  NAND2_X1 U8396 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n7232) );
  OAI211_X1 U8397 ( .C1(n6648), .C2(n9553), .A(n6647), .B(n7232), .ZN(n6649)
         );
  OR3_X1 U8398 ( .A1(n6651), .A2(n6650), .A3(n6649), .ZN(P1_U3249) );
  AOI211_X1 U8399 ( .C1(n6654), .C2(n6653), .A(n6652), .B(n9928), .ZN(n6663)
         );
  AOI211_X1 U8400 ( .C1(n6657), .C2(n6656), .A(n6655), .B(n9919), .ZN(n6662)
         );
  INV_X1 U8401 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n6660) );
  NAND2_X1 U8402 ( .A1(n9937), .A2(n6658), .ZN(n6659) );
  NAND2_X1 U8403 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n7168) );
  OAI211_X1 U8404 ( .C1(n6660), .C2(n9553), .A(n6659), .B(n7168), .ZN(n6661)
         );
  OR3_X1 U8405 ( .A1(n6663), .A2(n6662), .A3(n6661), .ZN(P1_U3248) );
  NAND2_X1 U8406 ( .A1(n6798), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6665) );
  OAI21_X1 U8407 ( .B1(n6798), .B2(P1_REG2_REG_7__SCAN_IN), .A(n6665), .ZN(
        n6666) );
  NOR2_X1 U8408 ( .A1(n6667), .A2(n6666), .ZN(n6793) );
  AOI211_X1 U8409 ( .C1(n6667), .C2(n6666), .A(n6793), .B(n9928), .ZN(n6678)
         );
  AOI21_X1 U8410 ( .B1(n6669), .B2(P1_REG1_REG_6__SCAN_IN), .A(n6668), .ZN(
        n6672) );
  NAND2_X1 U8411 ( .A1(n6798), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6670) );
  OAI21_X1 U8412 ( .B1(n6798), .B2(P1_REG1_REG_7__SCAN_IN), .A(n6670), .ZN(
        n6671) );
  NOR2_X1 U8413 ( .A1(n6672), .A2(n6671), .ZN(n6797) );
  AOI211_X1 U8414 ( .C1(n6672), .C2(n6671), .A(n6797), .B(n9919), .ZN(n6677)
         );
  INV_X1 U8415 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n6675) );
  NAND2_X1 U8416 ( .A1(n9937), .A2(n6798), .ZN(n6674) );
  INV_X1 U8417 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n8005) );
  NOR2_X1 U8418 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8005), .ZN(n7245) );
  INV_X1 U8419 ( .A(n7245), .ZN(n6673) );
  OAI211_X1 U8420 ( .C1(n6675), .C2(n9553), .A(n6674), .B(n6673), .ZN(n6676)
         );
  OR3_X1 U8421 ( .A1(n6678), .A2(n6677), .A3(n6676), .ZN(P1_U3250) );
  AOI211_X1 U8422 ( .C1(n6681), .C2(n6680), .A(n6679), .B(n9928), .ZN(n6690)
         );
  AOI211_X1 U8423 ( .C1(n6684), .C2(n6683), .A(n6682), .B(n9919), .ZN(n6689)
         );
  INV_X1 U8424 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n6687) );
  NAND2_X1 U8425 ( .A1(n9937), .A2(n8182), .ZN(n6686) );
  NAND2_X1 U8426 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_U3086), .ZN(n6685) );
  OAI211_X1 U8427 ( .C1(n6687), .C2(n9553), .A(n6686), .B(n6685), .ZN(n6688)
         );
  OR3_X1 U8428 ( .A1(n6690), .A2(n6689), .A3(n6688), .ZN(P1_U3246) );
  INV_X1 U8429 ( .A(n6692), .ZN(n6693) );
  AOI21_X1 U8430 ( .B1(n6694), .B2(n6691), .A(n6693), .ZN(n6700) );
  NAND2_X1 U8431 ( .A1(n6695), .A2(n9291), .ZN(n6697) );
  NAND2_X1 U8432 ( .A1(n9468), .A2(n9169), .ZN(n6696) );
  NAND2_X1 U8433 ( .A1(n6697), .A2(n6696), .ZN(n7041) );
  AOI22_X1 U8434 ( .A1(n9861), .A2(n7041), .B1(n6839), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n6699) );
  NAND2_X1 U8435 ( .A1(n9186), .A2(n5672), .ZN(n6698) );
  OAI211_X1 U8436 ( .C1(n6700), .C2(n9188), .A(n6699), .B(n6698), .ZN(P1_U3222) );
  NAND2_X1 U8437 ( .A1(n10107), .A2(n10116), .ZN(n10091) );
  OAI21_X1 U8438 ( .B1(n6702), .B2(n8434), .A(n6701), .ZN(n6943) );
  XNOR2_X1 U8439 ( .A(n6704), .B(n6703), .ZN(n6705) );
  NAND2_X1 U8440 ( .A1(n6705), .A2(n8895), .ZN(n6707) );
  AOI22_X1 U8441 ( .A1(n8898), .A2(n8609), .B1(n8607), .B2(n8899), .ZN(n6706)
         );
  NAND2_X1 U8442 ( .A1(n6707), .A2(n6706), .ZN(n6945) );
  AOI21_X1 U8443 ( .B1(n10091), .B2(n6943), .A(n6945), .ZN(n6867) );
  INV_X1 U8444 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n6708) );
  OAI22_X1 U8445 ( .A1(n8420), .A2(n9044), .B1(n10133), .B2(n6708), .ZN(n6709)
         );
  INV_X1 U8446 ( .A(n6709), .ZN(n6710) );
  OAI21_X1 U8447 ( .B1(n6867), .B2(n10135), .A(n6710), .ZN(P2_U3396) );
  INV_X1 U8448 ( .A(n6711), .ZN(n6757) );
  OAI222_X1 U8449 ( .A1(n8159), .A2(n6757), .B1(n8652), .B2(P2_U3151), .C1(
        n6712), .C2(n8186), .ZN(P2_U3281) );
  NAND2_X1 U8450 ( .A1(n6714), .A2(n6713), .ZN(n6719) );
  NAND3_X1 U8451 ( .A1(n6716), .A2(n6715), .A3(n7647), .ZN(n6717) );
  AOI21_X1 U8452 ( .B1(n6721), .B2(n6732), .A(n6717), .ZN(n6718) );
  NAND2_X1 U8453 ( .A1(n6719), .A2(n6718), .ZN(n6720) );
  NAND2_X1 U8454 ( .A1(n6720), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6723) );
  INV_X1 U8455 ( .A(n6741), .ZN(n6966) );
  NOR2_X1 U8456 ( .A1(n9051), .A2(n6966), .ZN(n8586) );
  NAND2_X1 U8457 ( .A1(n6721), .A2(n8586), .ZN(n6722) );
  NAND2_X1 U8458 ( .A1(n6724), .A2(n8378), .ZN(n6726) );
  XNOR2_X1 U8459 ( .A(n6728), .B(n6859), .ZN(n6727) );
  XNOR2_X1 U8460 ( .A(n6727), .B(n8609), .ZN(n6856) );
  AOI21_X1 U8461 ( .B1(n8227), .B2(n8972), .A(n8425), .ZN(n6857) );
  OAI22_X1 U8462 ( .A1(n6856), .A2(n6857), .B1(n8609), .B2(n6727), .ZN(n6758)
         );
  XNOR2_X1 U8463 ( .A(n6865), .B(n6728), .ZN(n6729) );
  XNOR2_X1 U8464 ( .A(n6729), .B(n8608), .ZN(n6759) );
  XNOR2_X1 U8465 ( .A(n6728), .B(n7108), .ZN(n6843) );
  XNOR2_X1 U8466 ( .A(n6843), .B(n8607), .ZN(n6735) );
  NAND2_X1 U8467 ( .A1(n6736), .A2(n6735), .ZN(n6842) );
  INV_X1 U8468 ( .A(n6730), .ZN(n6731) );
  NAND2_X1 U8469 ( .A1(n6737), .A2(n6731), .ZN(n6734) );
  NAND2_X1 U8470 ( .A1(n6742), .A2(n6732), .ZN(n6733) );
  INV_X1 U8471 ( .A(n8353), .ZN(n8321) );
  OAI211_X1 U8472 ( .C1(n6736), .C2(n6735), .A(n6842), .B(n8321), .ZN(n6749)
         );
  NAND2_X1 U8473 ( .A1(n6737), .A2(n10132), .ZN(n6740) );
  NAND2_X1 U8474 ( .A1(n6739), .A2(n6738), .ZN(n8770) );
  NAND2_X1 U8475 ( .A1(n6740), .A2(n8770), .ZN(n8351) );
  INV_X1 U8476 ( .A(n8606), .ZN(n6951) );
  AND2_X1 U8477 ( .A1(n6742), .A2(n6741), .ZN(n6745) );
  NAND2_X1 U8478 ( .A1(n6745), .A2(n6743), .ZN(n8349) );
  INV_X1 U8479 ( .A(n6743), .ZN(n6744) );
  NAND2_X1 U8480 ( .A1(n6745), .A2(n6744), .ZN(n8317) );
  OAI22_X1 U8481 ( .A1(n6951), .A2(n8349), .B1(n8317), .B2(n6754), .ZN(n6746)
         );
  AOI211_X1 U8482 ( .C1(n7108), .C2(n8351), .A(n6747), .B(n6746), .ZN(n6748)
         );
  OAI211_X1 U8483 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n8258), .A(n6749), .B(
        n6748), .ZN(P2_U3158) );
  OAI21_X1 U8484 ( .B1(n6752), .B2(n8425), .A(n6750), .ZN(n6958) );
  INV_X1 U8485 ( .A(n8610), .ZN(n6858) );
  INV_X1 U8486 ( .A(n8895), .ZN(n8970) );
  XNOR2_X1 U8487 ( .A(n6752), .B(n6751), .ZN(n6753) );
  OAI222_X1 U8488 ( .A1(n8860), .A2(n6754), .B1(n8858), .B2(n6858), .C1(n8970), 
        .C2(n6753), .ZN(n6959) );
  AOI21_X1 U8489 ( .B1(n10091), .B2(n6958), .A(n6959), .ZN(n6869) );
  INV_X1 U8490 ( .A(n6859), .ZN(n6962) );
  INV_X1 U8491 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n8084) );
  AOI22_X1 U8492 ( .A1(n9033), .A2(n6962), .B1(n10135), .B2(
        P2_REG0_REG_1__SCAN_IN), .ZN(n6755) );
  OAI21_X1 U8493 ( .B1(n6869), .B2(n10135), .A(n6755), .ZN(P2_U3393) );
  INV_X1 U8494 ( .A(n9487), .ZN(n7676) );
  OAI222_X1 U8495 ( .A1(P1_U3086), .A2(n7676), .B1(n7965), .B2(n6757), .C1(
        n6756), .C2(n8191), .ZN(P1_U3341) );
  XOR2_X1 U8496 ( .A(n6759), .B(n6758), .Z(n6763) );
  NAND2_X1 U8497 ( .A1(n8258), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6789) );
  INV_X1 U8498 ( .A(n8317), .ZN(n8345) );
  AOI22_X1 U8499 ( .A1(n8345), .A2(n8609), .B1(n8351), .B2(n6865), .ZN(n6760)
         );
  OAI21_X1 U8500 ( .B1(n6844), .B2(n8349), .A(n6760), .ZN(n6761) );
  AOI21_X1 U8501 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(n6789), .A(n6761), .ZN(
        n6762) );
  OAI21_X1 U8502 ( .B1(n6763), .B2(n8353), .A(n6762), .ZN(P2_U3177) );
  MUX2_X1 U8503 ( .A(P2_REG1_REG_5__SCAN_IN), .B(P2_REG2_REG_5__SCAN_IN), .S(
        n8748), .Z(n6808) );
  XOR2_X1 U8504 ( .A(n6810), .B(n6808), .Z(n6811) );
  AOI21_X1 U8505 ( .B1(n6766), .B2(n6765), .A(n6764), .ZN(n6812) );
  XOR2_X1 U8506 ( .A(n6811), .B(n6812), .Z(n6787) );
  OR2_X1 U8507 ( .A1(n6774), .A2(n10138), .ZN(n6767) );
  NAND2_X1 U8508 ( .A1(n6768), .A2(n6767), .ZN(n6769) );
  NAND2_X1 U8509 ( .A1(n6769), .A2(n6777), .ZN(n6822) );
  OAI21_X1 U8510 ( .B1(n6769), .B2(n6777), .A(n6822), .ZN(n6770) );
  INV_X1 U8511 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n10140) );
  NAND2_X1 U8512 ( .A1(n6770), .A2(n10140), .ZN(n6771) );
  NAND2_X1 U8513 ( .A1(n6824), .A2(n6771), .ZN(n6772) );
  AOI22_X1 U8514 ( .A1(n8757), .A2(P2_ADDR_REG_5__SCAN_IN), .B1(n8735), .B2(
        n6772), .ZN(n6785) );
  NOR2_X1 U8515 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6773), .ZN(n6954) );
  INV_X1 U8516 ( .A(n6954), .ZN(n6784) );
  NAND2_X1 U8517 ( .A1(n8699), .A2(n6810), .ZN(n6783) );
  OR2_X1 U8518 ( .A1(n6774), .A2(n7099), .ZN(n6775) );
  INV_X1 U8519 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n6778) );
  NAND2_X1 U8520 ( .A1(n6779), .A2(n6778), .ZN(n6780) );
  NAND2_X1 U8521 ( .A1(n6819), .A2(n6780), .ZN(n6781) );
  NAND2_X1 U8522 ( .A1(n8631), .A2(n6781), .ZN(n6782) );
  NAND4_X1 U8523 ( .A1(n6785), .A2(n6784), .A3(n6783), .A4(n6782), .ZN(n6786)
         );
  AOI21_X1 U8524 ( .B1(n6787), .B2(n8763), .A(n6786), .ZN(n6788) );
  INV_X1 U8525 ( .A(n6788), .ZN(P2_U3187) );
  INV_X1 U8526 ( .A(n6789), .ZN(n6860) );
  INV_X1 U8527 ( .A(n8349), .ZN(n8314) );
  INV_X1 U8528 ( .A(n8351), .ZN(n8329) );
  NAND2_X1 U8529 ( .A1(n8610), .A2(n8972), .ZN(n8433) );
  INV_X1 U8530 ( .A(n8433), .ZN(n6790) );
  OR2_X1 U8531 ( .A1(n6790), .A2(n8425), .ZN(n8975) );
  INV_X1 U8532 ( .A(n8975), .ZN(n8382) );
  OAI22_X1 U8533 ( .A1(n8329), .A2(n8972), .B1(n8353), .B2(n8382), .ZN(n6791)
         );
  AOI21_X1 U8534 ( .B1(n8314), .B2(n8609), .A(n6791), .ZN(n6792) );
  OAI21_X1 U8535 ( .B1(n6860), .B2(n5956), .A(n6792), .ZN(P2_U3172) );
  NAND2_X1 U8536 ( .A1(n6886), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6794) );
  OAI21_X1 U8537 ( .B1(n6886), .B2(P1_REG2_REG_8__SCAN_IN), .A(n6794), .ZN(
        n6795) );
  NOR2_X1 U8538 ( .A1(n6796), .A2(n6795), .ZN(n6885) );
  AOI211_X1 U8539 ( .C1(n6796), .C2(n6795), .A(n6885), .B(n9928), .ZN(n6807)
         );
  NAND2_X1 U8540 ( .A1(n6886), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6799) );
  OAI21_X1 U8541 ( .B1(n6886), .B2(P1_REG1_REG_8__SCAN_IN), .A(n6799), .ZN(
        n6800) );
  AOI211_X1 U8542 ( .C1(n6801), .C2(n6800), .A(n6881), .B(n9919), .ZN(n6806)
         );
  INV_X1 U8543 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n6804) );
  NAND2_X1 U8544 ( .A1(n9937), .A2(n6886), .ZN(n6803) );
  NAND2_X1 U8545 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n6802) );
  OAI211_X1 U8546 ( .C1(n6804), .C2(n9553), .A(n6803), .B(n6802), .ZN(n6805)
         );
  OR3_X1 U8547 ( .A1(n6807), .A2(n6806), .A3(n6805), .ZN(P1_U3251) );
  INV_X1 U8548 ( .A(n6808), .ZN(n6809) );
  OAI22_X1 U8549 ( .A1(n6812), .A2(n6811), .B1(n6810), .B2(n6809), .ZN(n6815)
         );
  INV_X1 U8550 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6821) );
  INV_X1 U8551 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6816) );
  MUX2_X1 U8552 ( .A(n6821), .B(n6816), .S(n8748), .Z(n6813) );
  INV_X1 U8553 ( .A(n6908), .ZN(n6830) );
  NAND2_X1 U8554 ( .A1(n6813), .A2(n6830), .ZN(n6898) );
  OAI21_X1 U8555 ( .B1(n6813), .B2(n6830), .A(n6898), .ZN(n6814) );
  NOR2_X1 U8556 ( .A1(n6815), .A2(n6814), .ZN(n6904) );
  AOI21_X1 U8557 ( .B1(n6815), .B2(n6814), .A(n6904), .ZN(n6832) );
  NAND2_X1 U8558 ( .A1(n8757), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n6828) );
  MUX2_X1 U8559 ( .A(n6816), .B(P2_REG2_REG_6__SCAN_IN), .S(n6908), .Z(n6818)
         );
  AND3_X1 U8560 ( .A1(n6819), .A2(n6818), .A3(n6817), .ZN(n6820) );
  OAI21_X1 U8561 ( .B1(n6907), .B2(n6820), .A(n8631), .ZN(n6827) );
  MUX2_X1 U8562 ( .A(n6821), .B(P2_REG1_REG_6__SCAN_IN), .S(n6908), .Z(n6823)
         );
  AND3_X1 U8563 ( .A1(n6824), .A2(n6823), .A3(n6822), .ZN(n6825) );
  OAI21_X1 U8564 ( .B1(n6895), .B2(n6825), .A(n8735), .ZN(n6826) );
  NAND2_X1 U8565 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3151), .ZN(n7154) );
  NAND4_X1 U8566 ( .A1(n6828), .A2(n6827), .A3(n6826), .A4(n7154), .ZN(n6829)
         );
  AOI21_X1 U8567 ( .B1(n6830), .B2(n8699), .A(n6829), .ZN(n6831) );
  OAI21_X1 U8568 ( .B1(n6832), .B2(n8695), .A(n6831), .ZN(P2_U3188) );
  OAI21_X1 U8569 ( .B1(n6835), .B2(n6834), .A(n6833), .ZN(n6836) );
  NAND2_X1 U8570 ( .A1(n6836), .A2(n9865), .ZN(n6841) );
  NAND2_X1 U8571 ( .A1(n9469), .A2(n9291), .ZN(n6838) );
  NAND2_X1 U8572 ( .A1(n9467), .A2(n9181), .ZN(n6837) );
  NAND2_X1 U8573 ( .A1(n6838), .A2(n6837), .ZN(n6977) );
  AOI22_X1 U8574 ( .A1(n9861), .A2(n6977), .B1(n6839), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n6840) );
  OAI211_X1 U8575 ( .C1(n9336), .C2(n9863), .A(n6841), .B(n6840), .ZN(P1_U3237) );
  XNOR2_X1 U8576 ( .A(n6728), .B(n10076), .ZN(n6950) );
  XOR2_X1 U8577 ( .A(n8606), .B(n6950), .Z(n6846) );
  AOI21_X1 U8578 ( .B1(n6846), .B2(n6845), .A(n6949), .ZN(n6851) );
  AOI22_X1 U8579 ( .A1(n8314), .A2(n8605), .B1(n8345), .B2(n8607), .ZN(n6848)
         );
  OAI211_X1 U8580 ( .C1(n8442), .C2(n8329), .A(n6848), .B(n6847), .ZN(n6849)
         );
  AOI21_X1 U8581 ( .B1(n7097), .B2(n8346), .A(n6849), .ZN(n6850) );
  OAI21_X1 U8582 ( .B1(n6851), .B2(n8353), .A(n6850), .ZN(P2_U3170) );
  INV_X1 U8583 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n8145) );
  INV_X1 U8584 ( .A(n6852), .ZN(n6855) );
  INV_X1 U8585 ( .A(n8673), .ZN(n6853) );
  OAI222_X1 U8586 ( .A1(n8186), .A2(n8145), .B1(n8159), .B2(n6855), .C1(
        P2_U3151), .C2(n6853), .ZN(P2_U3280) );
  INV_X1 U8587 ( .A(n9490), .ZN(n9505) );
  INV_X1 U8588 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6854) );
  OAI222_X1 U8589 ( .A1(n9505), .A2(P1_U3086), .B1(n7965), .B2(n6855), .C1(
        n6854), .C2(n8191), .ZN(P1_U3340) );
  XOR2_X1 U8590 ( .A(n6857), .B(n6856), .Z(n6864) );
  OAI22_X1 U8591 ( .A1(n8329), .A2(n6859), .B1(n6858), .B2(n8317), .ZN(n6862)
         );
  NOR2_X1 U8592 ( .A1(n6860), .A2(n4641), .ZN(n6861) );
  AOI211_X1 U8593 ( .C1(n8314), .C2(n8608), .A(n6862), .B(n6861), .ZN(n6863)
         );
  OAI21_X1 U8594 ( .B1(n8353), .B2(n6864), .A(n6863), .ZN(P2_U3162) );
  AOI22_X1 U8595 ( .A1(n8948), .A2(n6865), .B1(n10150), .B2(
        P2_REG1_REG_2__SCAN_IN), .ZN(n6866) );
  OAI21_X1 U8596 ( .B1(n6867), .B2(n10150), .A(n6866), .ZN(P2_U3461) );
  AOI22_X1 U8597 ( .A1(n8948), .A2(n6962), .B1(n10150), .B2(
        P2_REG1_REG_1__SCAN_IN), .ZN(n6868) );
  OAI21_X1 U8598 ( .B1(n6869), .B2(n10150), .A(n6868), .ZN(P2_U3460) );
  OAI21_X1 U8599 ( .B1(n6872), .B2(n6871), .A(n6870), .ZN(n6878) );
  OAI22_X1 U8600 ( .A1(n6874), .A2(n9106), .B1(n6873), .B2(n9096), .ZN(n7299)
         );
  AOI22_X1 U8601 ( .A1(n9861), .A2(n7299), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        P1_U3086), .ZN(n6876) );
  INV_X1 U8602 ( .A(n9868), .ZN(n9162) );
  NAND2_X1 U8603 ( .A1(n9162), .A2(n7306), .ZN(n6875) );
  OAI211_X1 U8604 ( .C1(n9976), .C2(n9863), .A(n6876), .B(n6875), .ZN(n6877)
         );
  AOI21_X1 U8605 ( .B1(n6878), .B2(n9865), .A(n6877), .ZN(n6879) );
  INV_X1 U8606 ( .A(n6879), .ZN(P1_U3218) );
  INV_X1 U8607 ( .A(n9919), .ZN(n9939) );
  NOR2_X1 U8608 ( .A1(n7022), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6880) );
  AOI21_X1 U8609 ( .B1(n7022), .B2(P1_REG1_REG_9__SCAN_IN), .A(n6880), .ZN(
        n6883) );
  OAI21_X1 U8610 ( .B1(n6883), .B2(n6882), .A(n7021), .ZN(n6890) );
  NOR2_X1 U8611 ( .A1(n7022), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6884) );
  AOI21_X1 U8612 ( .B1(P1_REG2_REG_9__SCAN_IN), .B2(n7022), .A(n6884), .ZN(
        n6888) );
  AOI21_X1 U8613 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n6886), .A(n6885), .ZN(
        n6887) );
  OAI21_X1 U8614 ( .B1(n6888), .B2(n6887), .A(n7017), .ZN(n6889) );
  AOI22_X1 U8615 ( .A1(n9939), .A2(n6890), .B1(n9915), .B2(n6889), .ZN(n6894)
         );
  INV_X1 U8616 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n6891) );
  NAND2_X1 U8617 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3086), .ZN(n7540) );
  OAI21_X1 U8618 ( .B1(n9553), .B2(n6891), .A(n7540), .ZN(n6892) );
  AOI21_X1 U8619 ( .B1(n7022), .B2(n9937), .A(n6892), .ZN(n6893) );
  NAND2_X1 U8620 ( .A1(n6894), .A2(n6893), .ZN(P1_U3252) );
  INV_X1 U8621 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n10143) );
  AOI21_X1 U8622 ( .B1(n4342), .B2(n6909), .A(n8621), .ZN(n6896) );
  INV_X1 U8623 ( .A(n6896), .ZN(n6897) );
  NAND2_X1 U8624 ( .A1(n6896), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n7003) );
  INV_X1 U8625 ( .A(n7003), .ZN(n8623) );
  AOI21_X1 U8626 ( .B1(n10143), .B2(n6897), .A(n8623), .ZN(n6920) );
  INV_X1 U8627 ( .A(n6898), .ZN(n6903) );
  INV_X1 U8628 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n7131) );
  MUX2_X1 U8629 ( .A(n10143), .B(n7131), .S(n8748), .Z(n6899) );
  NAND2_X1 U8630 ( .A1(n6899), .A2(n6909), .ZN(n8612) );
  INV_X1 U8631 ( .A(n6899), .ZN(n6900) );
  NAND2_X1 U8632 ( .A1(n6900), .A2(n4604), .ZN(n6901) );
  AND2_X1 U8633 ( .A1(n8612), .A2(n6901), .ZN(n6902) );
  OAI21_X1 U8634 ( .B1(n6904), .B2(n6903), .A(n6902), .ZN(n8613) );
  INV_X1 U8635 ( .A(n8613), .ZN(n6906) );
  NOR3_X1 U8636 ( .A1(n6904), .A2(n6903), .A3(n6902), .ZN(n6905) );
  OAI21_X1 U8637 ( .B1(n6906), .B2(n6905), .A(n8763), .ZN(n6919) );
  AOI21_X1 U8638 ( .B1(P2_REG2_REG_6__SCAN_IN), .B2(n6908), .A(n6907), .ZN(
        n6910) );
  NOR2_X1 U8639 ( .A1(n6910), .A2(n6909), .ZN(n8628) );
  OAI21_X1 U8640 ( .B1(n6912), .B2(P2_REG2_REG_7__SCAN_IN), .A(n8626), .ZN(
        n6917) );
  NAND2_X1 U8641 ( .A1(n8757), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n6915) );
  INV_X1 U8642 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n6913) );
  NOR2_X1 U8643 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6913), .ZN(n7254) );
  INV_X1 U8644 ( .A(n7254), .ZN(n6914) );
  OAI211_X1 U8645 ( .C1(n8761), .C2(n4604), .A(n6915), .B(n6914), .ZN(n6916)
         );
  AOI21_X1 U8646 ( .B1(n6917), .B2(n8631), .A(n6916), .ZN(n6918) );
  OAI211_X1 U8647 ( .C1(n6920), .C2(n8766), .A(n6919), .B(n6918), .ZN(P2_U3189) );
  INV_X1 U8648 ( .A(n6921), .ZN(n6929) );
  INV_X1 U8649 ( .A(n8675), .ZN(n8701) );
  OAI222_X1 U8650 ( .A1(n8159), .A2(n6929), .B1(n8701), .B2(P2_U3151), .C1(
        n8140), .C2(n8186), .ZN(P2_U3279) );
  AOI21_X1 U8651 ( .B1(n6923), .B2(n6922), .A(n9188), .ZN(n6925) );
  NAND2_X1 U8652 ( .A1(n6925), .A2(n6924), .ZN(n6928) );
  AOI22_X1 U8653 ( .A1(n9291), .A2(n9467), .B1(n9465), .B2(n9181), .ZN(n7312)
         );
  NAND2_X1 U8654 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3086), .ZN(n9923) );
  OAI21_X1 U8655 ( .B1(n9183), .B2(n7312), .A(n9923), .ZN(n6926) );
  AOI21_X1 U8656 ( .B1(n7317), .B2(n9186), .A(n6926), .ZN(n6927) );
  OAI211_X1 U8657 ( .C1(n9868), .C2(n7322), .A(n6928), .B(n6927), .ZN(P1_U3230) );
  INV_X1 U8658 ( .A(n9938), .ZN(n9503) );
  OAI222_X1 U8659 ( .A1(n8191), .A2(n6930), .B1(n7965), .B2(n6929), .C1(
        P1_U3086), .C2(n9503), .ZN(P1_U3339) );
  NAND2_X1 U8660 ( .A1(n6932), .A2(n6931), .ZN(n6939) );
  INV_X1 U8661 ( .A(n6933), .ZN(n6938) );
  NAND2_X1 U8662 ( .A1(n6724), .A2(n6934), .ZN(n6937) );
  NAND2_X1 U8663 ( .A1(n9052), .A2(n6935), .ZN(n6936) );
  NAND4_X1 U8664 ( .A1(n6939), .A2(n6938), .A3(n6937), .A4(n6936), .ZN(n6961)
         );
  OR2_X1 U8665 ( .A1(n6940), .A2(n7534), .ZN(n6941) );
  OR2_X1 U8666 ( .A1(n6961), .A2(n6941), .ZN(n7461) );
  NAND2_X1 U8667 ( .A1(n7461), .A2(n10107), .ZN(n6942) );
  NAND2_X1 U8668 ( .A1(n6942), .A2(n8915), .ZN(n8891) );
  INV_X1 U8669 ( .A(n6943), .ZN(n6948) );
  OAI22_X1 U8670 ( .A1(n8770), .A2(n8139), .B1(n8420), .B2(n8835), .ZN(n6944)
         );
  NOR2_X1 U8671 ( .A1(n6945), .A2(n6944), .ZN(n6946) );
  INV_X2 U8672 ( .A(n8915), .ZN(n8909) );
  MUX2_X1 U8673 ( .A(n6946), .B(n6550), .S(n8909), .Z(n6947) );
  OAI21_X1 U8674 ( .B1(n8891), .B2(n6948), .A(n6947), .ZN(P2_U3231) );
  XNOR2_X1 U8675 ( .A(n6728), .B(n7212), .ZN(n7148) );
  XOR2_X1 U8676 ( .A(n8605), .B(n7148), .Z(n7150) );
  XOR2_X1 U8677 ( .A(n7150), .B(n4421), .Z(n6957) );
  INV_X1 U8678 ( .A(n8604), .ZN(n6952) );
  OAI22_X1 U8679 ( .A1(n6952), .A2(n8349), .B1(n8317), .B2(n6951), .ZN(n6953)
         );
  AOI211_X1 U8680 ( .C1(n7212), .C2(n8351), .A(n6954), .B(n6953), .ZN(n6956)
         );
  NAND2_X1 U8681 ( .A1(n8346), .A2(n7214), .ZN(n6955) );
  OAI211_X1 U8682 ( .C1(n6957), .C2(n8353), .A(n6956), .B(n6955), .ZN(P2_U3167) );
  INV_X1 U8683 ( .A(n6958), .ZN(n6965) );
  INV_X1 U8684 ( .A(n6959), .ZN(n6960) );
  MUX2_X1 U8685 ( .A(n8013), .B(n6960), .S(n8915), .Z(n6964) );
  OR2_X1 U8686 ( .A1(n6961), .A2(n8835), .ZN(n8912) );
  INV_X1 U8687 ( .A(n8770), .ZN(n8908) );
  AOI22_X1 U8688 ( .A1(n8888), .A2(n6962), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n8908), .ZN(n6963) );
  OAI211_X1 U8689 ( .C1(n8891), .C2(n6965), .A(n6964), .B(n6963), .ZN(P2_U3232) );
  NAND2_X1 U8690 ( .A1(n8609), .A2(n8899), .ZN(n8971) );
  NAND3_X1 U8691 ( .A1(n8975), .A2(n6966), .A3(n10114), .ZN(n6967) );
  AOI21_X1 U8692 ( .B1(n8971), .B2(n6967), .A(n8909), .ZN(n6968) );
  AOI21_X1 U8693 ( .B1(n8888), .B2(n6969), .A(n6968), .ZN(n6971) );
  NAND2_X1 U8694 ( .A1(n8908), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n6970) );
  OAI211_X1 U8695 ( .C1(n6491), .C2(n8915), .A(n6971), .B(n6970), .ZN(P2_U3233) );
  XNOR2_X1 U8696 ( .A(n6972), .B(n9380), .ZN(n7198) );
  INV_X1 U8697 ( .A(n7198), .ZN(n6980) );
  INV_X1 U8698 ( .A(n10041), .ZN(n10033) );
  OR2_X1 U8699 ( .A1(n7045), .A2(n9336), .ZN(n6973) );
  AND3_X1 U8700 ( .A1(n7303), .A2(n9957), .A3(n6973), .ZN(n7195) );
  OAI21_X1 U8701 ( .B1(n9380), .B2(n6975), .A(n6974), .ZN(n6978) );
  NOR2_X1 U8702 ( .A1(n7198), .A2(n7434), .ZN(n6976) );
  AOI211_X1 U8703 ( .C1(n9698), .C2(n6978), .A(n6977), .B(n6976), .ZN(n7192)
         );
  INV_X1 U8704 ( .A(n7192), .ZN(n6979) );
  AOI211_X1 U8705 ( .C1(n6980), .C2(n10033), .A(n7195), .B(n6979), .ZN(n6984)
         );
  AOI22_X1 U8706 ( .A1(n9777), .A2(n6982), .B1(n10066), .B2(
        P1_REG1_REG_2__SCAN_IN), .ZN(n6981) );
  OAI21_X1 U8707 ( .B1(n6984), .B2(n10066), .A(n6981), .ZN(P1_U3524) );
  AOI22_X1 U8708 ( .A1(n9832), .A2(n6982), .B1(n10047), .B2(
        P1_REG0_REG_2__SCAN_IN), .ZN(n6983) );
  OAI21_X1 U8709 ( .B1(n6984), .B2(n10047), .A(n6983), .ZN(P1_U3459) );
  INV_X1 U8710 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n6987) );
  INV_X1 U8711 ( .A(n8628), .ZN(n6985) );
  INV_X1 U8712 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7056) );
  MUX2_X1 U8713 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n7056), .S(n8619), .Z(n8627)
         );
  AOI21_X1 U8714 ( .B1(n6987), .B2(n6986), .A(n7077), .ZN(n7012) );
  INV_X1 U8715 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n7001) );
  MUX2_X1 U8716 ( .A(n7001), .B(n7056), .S(n8748), .Z(n6988) );
  NAND2_X1 U8717 ( .A1(n6988), .A2(n8619), .ZN(n6991) );
  INV_X1 U8718 ( .A(n6988), .ZN(n6989) );
  NAND2_X1 U8719 ( .A1(n6989), .A2(n7004), .ZN(n6990) );
  NAND2_X1 U8720 ( .A1(n6991), .A2(n6990), .ZN(n8611) );
  AOI21_X1 U8721 ( .B1(n8613), .B2(n8612), .A(n8611), .ZN(n8615) );
  INV_X1 U8722 ( .A(n6991), .ZN(n6997) );
  INV_X1 U8723 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n6992) );
  MUX2_X1 U8724 ( .A(n6992), .B(n6987), .S(n8748), .Z(n6993) );
  NAND2_X1 U8725 ( .A1(n6993), .A2(n7076), .ZN(n7072) );
  INV_X1 U8726 ( .A(n6993), .ZN(n6994) );
  NAND2_X1 U8727 ( .A1(n6994), .A2(n7005), .ZN(n6995) );
  AND2_X1 U8728 ( .A1(n7072), .A2(n6995), .ZN(n6996) );
  OAI21_X1 U8729 ( .B1(n8615), .B2(n6997), .A(n6996), .ZN(n7073) );
  INV_X1 U8730 ( .A(n7073), .ZN(n6999) );
  NOR3_X1 U8731 ( .A1(n8615), .A2(n6997), .A3(n6996), .ZN(n6998) );
  OAI21_X1 U8732 ( .B1(n6999), .B2(n6998), .A(n8763), .ZN(n7011) );
  INV_X1 U8733 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n7000) );
  NAND2_X1 U8734 ( .A1(P2_U3151), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n7472) );
  OAI21_X1 U8735 ( .B1(n8724), .B2(n7000), .A(n7472), .ZN(n7009) );
  INV_X1 U8736 ( .A(n8621), .ZN(n7002) );
  MUX2_X1 U8737 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n7001), .S(n8619), .Z(n8620)
         );
  AOI21_X1 U8738 ( .B1(n7003), .B2(n7002), .A(n8620), .ZN(n8625) );
  AOI21_X1 U8739 ( .B1(P2_REG1_REG_8__SCAN_IN), .B2(n7004), .A(n8625), .ZN(
        n7060) );
  XOR2_X1 U8740 ( .A(n7060), .B(n7005), .Z(n7006) );
  NOR2_X1 U8741 ( .A1(n6992), .A2(n7006), .ZN(n7061) );
  AOI21_X1 U8742 ( .B1(n6992), .B2(n7006), .A(n7061), .ZN(n7007) );
  NOR2_X1 U8743 ( .A1(n7007), .A2(n8766), .ZN(n7008) );
  AOI211_X1 U8744 ( .C1(n8699), .C2(n7076), .A(n7009), .B(n7008), .ZN(n7010)
         );
  OAI211_X1 U8745 ( .C1(n7012), .C2(n8756), .A(n7011), .B(n7010), .ZN(P2_U3191) );
  INV_X1 U8746 ( .A(n7013), .ZN(n7015) );
  INV_X1 U8747 ( .A(n8728), .ZN(n8702) );
  OAI222_X1 U8748 ( .A1(n8186), .A2(n7014), .B1(n8159), .B2(n7015), .C1(
        P2_U3151), .C2(n8702), .ZN(P2_U3278) );
  INV_X1 U8749 ( .A(n9519), .ZN(n9527) );
  OAI222_X1 U8750 ( .A1(n8191), .A2(n7016), .B1(n7965), .B2(n7015), .C1(n9527), 
        .C2(P1_U3086), .ZN(P1_U3338) );
  OAI21_X1 U8751 ( .B1(n7022), .B2(P1_REG2_REG_9__SCAN_IN), .A(n7017), .ZN(
        n7020) );
  NAND2_X1 U8752 ( .A1(n7266), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n7018) );
  OAI21_X1 U8753 ( .B1(n7266), .B2(P1_REG2_REG_10__SCAN_IN), .A(n7018), .ZN(
        n7019) );
  NOR2_X1 U8754 ( .A1(n7019), .A2(n7020), .ZN(n7262) );
  AOI211_X1 U8755 ( .C1(n7020), .C2(n7019), .A(n7262), .B(n9928), .ZN(n7030)
         );
  OAI21_X1 U8756 ( .B1(n7022), .B2(P1_REG1_REG_9__SCAN_IN), .A(n7021), .ZN(
        n7025) );
  INV_X1 U8757 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n7023) );
  MUX2_X1 U8758 ( .A(n7023), .B(P1_REG1_REG_10__SCAN_IN), .S(n7266), .Z(n7024)
         );
  NOR2_X1 U8759 ( .A1(n7024), .A2(n7025), .ZN(n7265) );
  AOI211_X1 U8760 ( .C1(n7025), .C2(n7024), .A(n7265), .B(n9919), .ZN(n7029)
         );
  INV_X1 U8761 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n7027) );
  NAND2_X1 U8762 ( .A1(n9937), .A2(n7266), .ZN(n7026) );
  NAND2_X1 U8763 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n9858) );
  OAI211_X1 U8764 ( .C1(n7027), .C2(n9553), .A(n7026), .B(n9858), .ZN(n7028)
         );
  OR3_X1 U8765 ( .A1(n7030), .A2(n7029), .A3(n7028), .ZN(P1_U3253) );
  NAND3_X1 U8766 ( .A1(n7033), .A2(n7032), .A3(n7031), .ZN(n7034) );
  AND2_X1 U8767 ( .A1(n7434), .A2(n7191), .ZN(n7035) );
  XNOR2_X1 U8768 ( .A(n7036), .B(n4543), .ZN(n9967) );
  NAND2_X1 U8769 ( .A1(n7038), .A2(n7037), .ZN(n7039) );
  NAND2_X1 U8770 ( .A1(n7040), .A2(n7039), .ZN(n7042) );
  AOI21_X1 U8771 ( .B1(n7042), .B2(n9698), .A(n7041), .ZN(n9969) );
  OAI22_X1 U8772 ( .A1(n9969), .A2(n4334), .B1(n9470), .B2(n9727), .ZN(n7049)
         );
  INV_X1 U8773 ( .A(n7043), .ZN(n7044) );
  INV_X1 U8774 ( .A(n7045), .ZN(n7046) );
  OAI211_X1 U8775 ( .C1(n9970), .C2(n7047), .A(n7046), .B(n9957), .ZN(n9968)
         );
  OAI22_X1 U8776 ( .A1(n9970), .A2(n9716), .B1(n9671), .B2(n9968), .ZN(n7048)
         );
  AOI211_X1 U8777 ( .C1(n4334), .C2(P1_REG2_REG_1__SCAN_IN), .A(n7049), .B(
        n7048), .ZN(n7050) );
  OAI21_X1 U8778 ( .B1(n9720), .B2(n9967), .A(n7050), .ZN(P1_U3292) );
  NAND2_X1 U8779 ( .A1(n8416), .A2(n8450), .ZN(n8386) );
  NAND2_X1 U8780 ( .A1(n7124), .A2(n7051), .ZN(n7052) );
  XOR2_X1 U8781 ( .A(n8386), .B(n7052), .Z(n10103) );
  XNOR2_X1 U8782 ( .A(n7053), .B(n8386), .ZN(n7054) );
  OAI222_X1 U8783 ( .A1(n8858), .A2(n7463), .B1(n8860), .B2(n7716), .C1(n7054), 
        .C2(n8970), .ZN(n10105) );
  NAND2_X1 U8784 ( .A1(n10105), .A2(n8915), .ZN(n7059) );
  INV_X1 U8785 ( .A(n7055), .ZN(n7572) );
  OAI22_X1 U8786 ( .A1(n8915), .A2(n7056), .B1(n7572), .B2(n8770), .ZN(n7057)
         );
  AOI21_X1 U8787 ( .B1(n8888), .B2(n7578), .A(n7057), .ZN(n7058) );
  OAI211_X1 U8788 ( .C1(n10103), .C2(n8891), .A(n7059), .B(n7058), .ZN(
        P2_U3225) );
  NOR2_X1 U8789 ( .A1(n7076), .A2(n7060), .ZN(n7062) );
  INV_X1 U8790 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n7066) );
  MUX2_X1 U8791 ( .A(n7066), .B(P2_REG1_REG_10__SCAN_IN), .S(n7395), .Z(n7064)
         );
  INV_X1 U8792 ( .A(n7381), .ZN(n7063) );
  AOI21_X1 U8793 ( .B1(n7065), .B2(n7064), .A(n7063), .ZN(n7089) );
  INV_X1 U8794 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7457) );
  MUX2_X1 U8795 ( .A(n7066), .B(n7457), .S(n8748), .Z(n7068) );
  NAND2_X1 U8796 ( .A1(n7068), .A2(n7067), .ZN(n7383) );
  INV_X1 U8797 ( .A(n7068), .ZN(n7069) );
  NAND2_X1 U8798 ( .A1(n7069), .A2(n7395), .ZN(n7070) );
  NAND2_X1 U8799 ( .A1(n7383), .A2(n7070), .ZN(n7071) );
  AOI21_X1 U8800 ( .B1(n7073), .B2(n7072), .A(n7071), .ZN(n7390) );
  AND3_X1 U8801 ( .A1(n7073), .A2(n7072), .A3(n7071), .ZN(n7074) );
  OAI21_X1 U8802 ( .B1(n7390), .B2(n7074), .A(n8763), .ZN(n7088) );
  NOR2_X1 U8803 ( .A1(n7076), .A2(n7075), .ZN(n7078) );
  INV_X1 U8804 ( .A(n7080), .ZN(n7082) );
  MUX2_X1 U8805 ( .A(n7457), .B(P2_REG2_REG_10__SCAN_IN), .S(n7395), .Z(n7079)
         );
  INV_X1 U8806 ( .A(n7079), .ZN(n7081) );
  OAI21_X1 U8807 ( .B1(n7082), .B2(n7081), .A(n7397), .ZN(n7086) );
  NOR2_X1 U8808 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7083), .ZN(n7788) );
  AOI21_X1 U8809 ( .B1(n8757), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n7788), .ZN(
        n7084) );
  OAI21_X1 U8810 ( .B1(n7395), .B2(n8761), .A(n7084), .ZN(n7085) );
  AOI21_X1 U8811 ( .B1(n7086), .B2(n8631), .A(n7085), .ZN(n7087) );
  OAI211_X1 U8812 ( .C1(n7089), .C2(n8766), .A(n7088), .B(n7087), .ZN(P2_U3192) );
  XNOR2_X1 U8813 ( .A(n7090), .B(n8439), .ZN(n7091) );
  NAND2_X1 U8814 ( .A1(n7091), .A2(n8895), .ZN(n7093) );
  AOI22_X1 U8815 ( .A1(n8898), .A2(n8607), .B1(n8605), .B2(n8899), .ZN(n7092)
         );
  AND2_X1 U8816 ( .A1(n7093), .A2(n7092), .ZN(n10079) );
  OR2_X1 U8817 ( .A1(n7094), .A2(n8439), .ZN(n7095) );
  NAND2_X1 U8818 ( .A1(n7096), .A2(n7095), .ZN(n10078) );
  INV_X1 U8819 ( .A(n8891), .ZN(n8906) );
  AOI22_X1 U8820 ( .A1(n8888), .A2(n10076), .B1(n8908), .B2(n7097), .ZN(n7098)
         );
  OAI21_X1 U8821 ( .B1(n7099), .B2(n8915), .A(n7098), .ZN(n7100) );
  AOI21_X1 U8822 ( .B1(n10078), .B2(n8906), .A(n7100), .ZN(n7101) );
  OAI21_X1 U8823 ( .B1(n10079), .B2(n8909), .A(n7101), .ZN(P2_U3229) );
  INV_X1 U8824 ( .A(n7102), .ZN(n7145) );
  INV_X1 U8825 ( .A(n9530), .ZN(n9531) );
  OAI222_X1 U8826 ( .A1(n8191), .A2(n7103), .B1(n7965), .B2(n7145), .C1(
        P1_U3086), .C2(n9531), .ZN(P1_U3337) );
  XNOR2_X1 U8827 ( .A(n7105), .B(n7104), .ZN(n7106) );
  AOI222_X1 U8828 ( .A1(n8895), .A2(n7106), .B1(n8608), .B2(n8898), .C1(n8606), 
        .C2(n8899), .ZN(n10071) );
  XNOR2_X1 U8829 ( .A(n8381), .B(n7107), .ZN(n10074) );
  AOI22_X1 U8830 ( .A1(n8888), .A2(n7108), .B1(n5985), .B2(n8908), .ZN(n7109)
         );
  OAI21_X1 U8831 ( .B1(n7110), .B2(n8915), .A(n7109), .ZN(n7111) );
  AOI21_X1 U8832 ( .B1(n10074), .B2(n8906), .A(n7111), .ZN(n7112) );
  OAI21_X1 U8833 ( .B1(n10071), .B2(n8909), .A(n7112), .ZN(P2_U3230) );
  NAND2_X1 U8834 ( .A1(n7113), .A2(n7125), .ZN(n8383) );
  XNOR2_X1 U8835 ( .A(n7114), .B(n8383), .ZN(n7115) );
  AOI222_X1 U8836 ( .A1(n8895), .A2(n7115), .B1(n8603), .B2(n8899), .C1(n8605), 
        .C2(n8898), .ZN(n10088) );
  OAI21_X1 U8837 ( .B1(n7213), .B2(n8457), .A(n7116), .ZN(n7117) );
  XOR2_X1 U8838 ( .A(n8383), .B(n7117), .Z(n10092) );
  NOR2_X1 U8839 ( .A1(n8912), .A2(n10089), .ZN(n7120) );
  INV_X1 U8840 ( .A(n7158), .ZN(n7118) );
  OAI22_X1 U8841 ( .A1(n8915), .A2(n6816), .B1(n7118), .B2(n8770), .ZN(n7119)
         );
  AOI211_X1 U8842 ( .C1(n10092), .C2(n8906), .A(n7120), .B(n7119), .ZN(n7121)
         );
  OAI21_X1 U8843 ( .B1(n10088), .B2(n8909), .A(n7121), .ZN(P2_U3227) );
  NAND2_X1 U8844 ( .A1(n7122), .A2(n8466), .ZN(n7123) );
  NAND2_X1 U8845 ( .A1(n7124), .A2(n7123), .ZN(n10097) );
  NAND2_X1 U8846 ( .A1(n7126), .A2(n7125), .ZN(n7127) );
  INV_X1 U8847 ( .A(n8466), .ZN(n8448) );
  XNOR2_X1 U8848 ( .A(n7127), .B(n8448), .ZN(n7128) );
  NAND2_X1 U8849 ( .A1(n7128), .A2(n8895), .ZN(n7130) );
  AOI22_X1 U8850 ( .A1(n8898), .A2(n8604), .B1(n8602), .B2(n8899), .ZN(n7129)
         );
  AND2_X1 U8851 ( .A1(n7130), .A2(n7129), .ZN(n10099) );
  MUX2_X1 U8852 ( .A(n10099), .B(n7131), .S(n8909), .Z(n7133) );
  AOI22_X1 U8853 ( .A1(n8888), .A2(n10094), .B1(n8908), .B2(n7253), .ZN(n7132)
         );
  OAI211_X1 U8854 ( .C1(n8891), .C2(n10097), .A(n7133), .B(n7132), .ZN(
        P2_U3226) );
  NAND2_X1 U8855 ( .A1(n7134), .A2(n8387), .ZN(n7135) );
  NAND2_X1 U8856 ( .A1(n7136), .A2(n7135), .ZN(n10109) );
  XNOR2_X1 U8857 ( .A(n7137), .B(n8387), .ZN(n7138) );
  NAND2_X1 U8858 ( .A1(n7138), .A2(n8895), .ZN(n7140) );
  AOI22_X1 U8859 ( .A1(n8600), .A2(n8899), .B1(n8898), .B2(n8602), .ZN(n7139)
         );
  NAND2_X1 U8860 ( .A1(n7140), .A2(n7139), .ZN(n10112) );
  NAND2_X1 U8861 ( .A1(n10112), .A2(n8915), .ZN(n7144) );
  INV_X1 U8862 ( .A(n7141), .ZN(n7471) );
  OAI22_X1 U8863 ( .A1(n8915), .A2(n6987), .B1(n7471), .B2(n8770), .ZN(n7142)
         );
  AOI21_X1 U8864 ( .B1(n8888), .B2(n7468), .A(n7142), .ZN(n7143) );
  OAI211_X1 U8865 ( .C1(n8891), .C2(n10109), .A(n7144), .B(n7143), .ZN(
        P2_U3224) );
  INV_X1 U8866 ( .A(n8747), .ZN(n8730) );
  OAI222_X1 U8867 ( .A1(n8186), .A2(n7146), .B1(n8730), .B2(P2_U3151), .C1(
        n8159), .C2(n7145), .ZN(P2_U3277) );
  XNOR2_X1 U8868 ( .A(n8200), .B(n7147), .ZN(n7248) );
  XOR2_X1 U8869 ( .A(n8604), .B(n7248), .Z(n7152) );
  INV_X1 U8870 ( .A(n7148), .ZN(n7149) );
  AOI211_X1 U8871 ( .C1(n7152), .C2(n7151), .A(n8353), .B(n7249), .ZN(n7153)
         );
  INV_X1 U8872 ( .A(n7153), .ZN(n7160) );
  NOR2_X1 U8873 ( .A1(n8349), .A2(n7463), .ZN(n7157) );
  OAI21_X1 U8874 ( .B1(n8317), .B2(n7155), .A(n7154), .ZN(n7156) );
  AOI211_X1 U8875 ( .C1(n7158), .C2(n8346), .A(n7157), .B(n7156), .ZN(n7159)
         );
  OAI211_X1 U8876 ( .C1(n10089), .C2(n8329), .A(n7160), .B(n7159), .ZN(
        P2_U3179) );
  INV_X1 U8877 ( .A(n7161), .ZN(n7163) );
  INV_X1 U8878 ( .A(n7162), .ZN(n7164) );
  NAND2_X1 U8879 ( .A1(n7163), .A2(n7164), .ZN(n7224) );
  NAND2_X1 U8880 ( .A1(n7161), .A2(n7162), .ZN(n7165) );
  NAND2_X1 U8881 ( .A1(n7224), .A2(n7165), .ZN(n7166) );
  NOR2_X1 U8882 ( .A1(n7166), .A2(n7167), .ZN(n7227) );
  AOI21_X1 U8883 ( .B1(n7167), .B2(n7166), .A(n7227), .ZN(n7172) );
  AOI22_X1 U8884 ( .A1(n9169), .A2(n9464), .B1(n9466), .B2(n9291), .ZN(n7201)
         );
  OAI21_X1 U8885 ( .B1(n9183), .B2(n7201), .A(n7168), .ZN(n7170) );
  NOR2_X1 U8886 ( .A1(n9868), .A2(n7206), .ZN(n7169) );
  AOI211_X1 U8887 ( .C1(n9992), .C2(n9186), .A(n7170), .B(n7169), .ZN(n7171)
         );
  OAI21_X1 U8888 ( .B1(n7172), .B2(n9188), .A(n7171), .ZN(P1_U3227) );
  INV_X1 U8889 ( .A(n7174), .ZN(n9386) );
  XNOR2_X1 U8890 ( .A(n7173), .B(n9386), .ZN(n9999) );
  XNOR2_X1 U8891 ( .A(n7175), .B(n9386), .ZN(n7176) );
  INV_X1 U8892 ( .A(n9698), .ZN(n9945) );
  AOI22_X1 U8893 ( .A1(n9291), .A2(n9465), .B1(n9463), .B2(n9181), .ZN(n7233)
         );
  OAI21_X1 U8894 ( .B1(n7176), .B2(n9945), .A(n7233), .ZN(n10002) );
  NAND2_X1 U8895 ( .A1(n10002), .A2(n9723), .ZN(n7181) );
  OAI22_X1 U8896 ( .A1(n9723), .A2(n5057), .B1(n7231), .B2(n9727), .ZN(n7178)
         );
  OAI211_X1 U8897 ( .C1(n7203), .C2(n10001), .A(n9957), .B(n9955), .ZN(n10000)
         );
  NOR2_X1 U8898 ( .A1(n10000), .A2(n9671), .ZN(n7177) );
  AOI211_X1 U8899 ( .C1(n9953), .C2(n7179), .A(n7178), .B(n7177), .ZN(n7180)
         );
  OAI211_X1 U8900 ( .C1(n9999), .C2(n9720), .A(n7181), .B(n7180), .ZN(P1_U3287) );
  NOR2_X1 U8901 ( .A1(n9671), .A2(n9977), .ZN(n7305) );
  OAI21_X1 U8902 ( .B1(n7305), .B2(n9953), .A(n7182), .ZN(n7189) );
  INV_X1 U8903 ( .A(n9379), .ZN(n7186) );
  INV_X1 U8904 ( .A(n9727), .ZN(n9951) );
  NAND2_X1 U8905 ( .A1(n9951), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n7183) );
  OAI211_X1 U8906 ( .C1(n7186), .C2(n7185), .A(n7184), .B(n7183), .ZN(n7187)
         );
  NAND2_X1 U8907 ( .A1(n9723), .A2(n7187), .ZN(n7188) );
  OAI211_X1 U8908 ( .C1(n9723), .C2(n7190), .A(n7189), .B(n7188), .ZN(P1_U3293) );
  OR2_X1 U8909 ( .A1(n4334), .A2(n7191), .ZN(n7443) );
  MUX2_X1 U8910 ( .A(n7193), .B(n7192), .S(n9723), .Z(n7197) );
  OAI22_X1 U8911 ( .A1(n9716), .A2(n9336), .B1(n4960), .B2(n9727), .ZN(n7194)
         );
  AOI21_X1 U8912 ( .B1(n9960), .B2(n7195), .A(n7194), .ZN(n7196) );
  OAI211_X1 U8913 ( .C1(n7198), .C2(n7443), .A(n7197), .B(n7196), .ZN(P1_U3291) );
  XOR2_X1 U8914 ( .A(n7199), .B(n9383), .Z(n9996) );
  XOR2_X1 U8915 ( .A(n7200), .B(n9383), .Z(n7202) );
  OAI21_X1 U8916 ( .B1(n7202), .B2(n9945), .A(n7201), .ZN(n9998) );
  NAND2_X1 U8917 ( .A1(n9998), .A2(n9723), .ZN(n7211) );
  INV_X1 U8918 ( .A(n7321), .ZN(n7204) );
  AOI211_X1 U8919 ( .C1(n9992), .C2(n7204), .A(n9977), .B(n7203), .ZN(n9991)
         );
  NOR2_X1 U8920 ( .A1(n9716), .A2(n7205), .ZN(n7209) );
  OAI22_X1 U8921 ( .A1(n9723), .A2(n7207), .B1(n7206), .B2(n9727), .ZN(n7208)
         );
  AOI211_X1 U8922 ( .C1(n9991), .C2(n9960), .A(n7209), .B(n7208), .ZN(n7210)
         );
  OAI211_X1 U8923 ( .C1(n9996), .C2(n9720), .A(n7211), .B(n7210), .ZN(P1_U3288) );
  INV_X1 U8924 ( .A(n7461), .ZN(n8781) );
  XNOR2_X1 U8925 ( .A(n8605), .B(n7212), .ZN(n8384) );
  XNOR2_X1 U8926 ( .A(n7213), .B(n8384), .ZN(n10082) );
  INV_X1 U8927 ( .A(n7214), .ZN(n7215) );
  OAI22_X1 U8928 ( .A1(n8912), .A2(n10083), .B1(n7215), .B2(n8770), .ZN(n7222)
         );
  XOR2_X1 U8929 ( .A(n7216), .B(n8384), .Z(n7220) );
  NAND2_X1 U8930 ( .A1(n10082), .A2(n7217), .ZN(n7219) );
  AOI22_X1 U8931 ( .A1(n8898), .A2(n8606), .B1(n8604), .B2(n8899), .ZN(n7218)
         );
  OAI211_X1 U8932 ( .C1(n7220), .C2(n8970), .A(n7219), .B(n7218), .ZN(n10086)
         );
  MUX2_X1 U8933 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n10086), .S(n8915), .Z(n7221)
         );
  AOI211_X1 U8934 ( .C1(n8781), .C2(n10082), .A(n7222), .B(n7221), .ZN(n7223)
         );
  INV_X1 U8935 ( .A(n7223), .ZN(P2_U3228) );
  INV_X1 U8936 ( .A(n7224), .ZN(n7225) );
  NOR3_X1 U8937 ( .A1(n7227), .A2(n7226), .A3(n7225), .ZN(n7230) );
  INV_X1 U8938 ( .A(n7228), .ZN(n7229) );
  OAI21_X1 U8939 ( .B1(n7230), .B2(n7229), .A(n9865), .ZN(n7237) );
  INV_X1 U8940 ( .A(n7231), .ZN(n7235) );
  OAI21_X1 U8941 ( .B1(n9183), .B2(n7233), .A(n7232), .ZN(n7234) );
  AOI21_X1 U8942 ( .B1(n7235), .B2(n9162), .A(n7234), .ZN(n7236) );
  OAI211_X1 U8943 ( .C1(n10001), .C2(n9863), .A(n7237), .B(n7236), .ZN(
        P1_U3239) );
  AND3_X1 U8944 ( .A1(n7228), .A2(n7239), .A3(n7238), .ZN(n7240) );
  OAI21_X1 U8945 ( .B1(n7241), .B2(n7240), .A(n9865), .ZN(n7247) );
  NAND2_X1 U8946 ( .A1(n9462), .A2(n9181), .ZN(n7243) );
  NAND2_X1 U8947 ( .A1(n9464), .A2(n9291), .ZN(n7242) );
  NAND2_X1 U8948 ( .A1(n7243), .A2(n7242), .ZN(n9949) );
  NOR2_X1 U8949 ( .A1(n9868), .A2(n9950), .ZN(n7244) );
  AOI211_X1 U8950 ( .C1(n9861), .C2(n9949), .A(n7245), .B(n7244), .ZN(n7246)
         );
  OAI211_X1 U8951 ( .C1(n4479), .C2(n9863), .A(n7247), .B(n7246), .ZN(P1_U3213) );
  INV_X1 U8952 ( .A(n7248), .ZN(n7250) );
  XNOR2_X1 U8953 ( .A(n8200), .B(n10094), .ZN(n7462) );
  XNOR2_X1 U8954 ( .A(n7462), .B(n8603), .ZN(n7251) );
  OAI21_X1 U8955 ( .B1(n7252), .B2(n7251), .A(n7465), .ZN(n7260) );
  AND2_X1 U8956 ( .A1(n8351), .A2(n10094), .ZN(n7259) );
  INV_X1 U8957 ( .A(n7253), .ZN(n7257) );
  AOI21_X1 U8958 ( .B1(n8345), .B2(n8604), .A(n7254), .ZN(n7256) );
  OR2_X1 U8959 ( .A1(n8349), .A2(n7474), .ZN(n7255) );
  OAI211_X1 U8960 ( .C1(n8258), .C2(n7257), .A(n7256), .B(n7255), .ZN(n7258)
         );
  AOI211_X1 U8961 ( .C1(n7260), .C2(n8321), .A(n7259), .B(n7258), .ZN(n7261)
         );
  INV_X1 U8962 ( .A(n7261), .ZN(P2_U3153) );
  XNOR2_X1 U8963 ( .A(n7346), .B(P1_REG2_REG_11__SCAN_IN), .ZN(n7263) );
  NOR2_X1 U8964 ( .A1(n7263), .A2(n7264), .ZN(n7345) );
  AOI211_X1 U8965 ( .C1(n7264), .C2(n7263), .A(n7345), .B(n9928), .ZN(n7274)
         );
  INV_X1 U8966 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n7267) );
  MUX2_X1 U8967 ( .A(n7267), .B(P1_REG1_REG_11__SCAN_IN), .S(n7346), .Z(n7268)
         );
  AOI211_X1 U8968 ( .C1(n7269), .C2(n7268), .A(n7341), .B(n9919), .ZN(n7273)
         );
  INV_X1 U8969 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n7271) );
  NAND2_X1 U8970 ( .A1(n9937), .A2(n7346), .ZN(n7270) );
  NAND2_X1 U8971 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n7808) );
  OAI211_X1 U8972 ( .C1(n7271), .C2(n9553), .A(n7270), .B(n7808), .ZN(n7272)
         );
  OR3_X1 U8973 ( .A1(n7274), .A2(n7273), .A3(n7272), .ZN(P1_U3254) );
  INV_X1 U8974 ( .A(n7275), .ZN(n8158) );
  OAI222_X1 U8975 ( .A1(n9376), .A2(P1_U3086), .B1(n7965), .B2(n8158), .C1(
        n7276), .C2(n8191), .ZN(P1_U3336) );
  INV_X1 U8976 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10159) );
  NOR2_X1 U8977 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7277) );
  AOI21_X1 U8978 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n7277), .ZN(n10164) );
  NOR2_X1 U8979 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7278) );
  AOI21_X1 U8980 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n7278), .ZN(n10167) );
  NOR2_X1 U8981 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7279) );
  AOI21_X1 U8982 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n7279), .ZN(n10170) );
  NOR2_X1 U8983 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7280) );
  AOI21_X1 U8984 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n7280), .ZN(n10173) );
  NOR2_X1 U8985 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7281) );
  AOI21_X1 U8986 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n7281), .ZN(n10176) );
  NOR2_X1 U8987 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7282) );
  AOI21_X1 U8988 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n7282), .ZN(n10179) );
  NOR2_X1 U8989 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n7283) );
  AOI21_X1 U8990 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n7283), .ZN(n10182) );
  NOR2_X1 U8991 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n7284) );
  AOI21_X1 U8992 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n7284), .ZN(n10185) );
  NOR2_X1 U8993 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n7285) );
  AOI21_X1 U8994 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(P2_ADDR_REG_9__SCAN_IN), 
        .A(n7285), .ZN(n10194) );
  NOR2_X1 U8995 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n7286) );
  AOI21_X1 U8996 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(P2_ADDR_REG_8__SCAN_IN), 
        .A(n7286), .ZN(n10200) );
  NOR2_X1 U8997 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n7287) );
  AOI21_X1 U8998 ( .B1(P1_ADDR_REG_7__SCAN_IN), .B2(P2_ADDR_REG_7__SCAN_IN), 
        .A(n7287), .ZN(n10197) );
  NOR2_X1 U8999 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n7288) );
  AOI21_X1 U9000 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(P2_ADDR_REG_6__SCAN_IN), 
        .A(n7288), .ZN(n10191) );
  NOR2_X1 U9001 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n7289) );
  AOI21_X1 U9002 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(P2_ADDR_REG_5__SCAN_IN), 
        .A(n7289), .ZN(n10188) );
  AND2_X1 U9003 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n7290) );
  NOR2_X1 U9004 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n7290), .ZN(n10154) );
  INV_X1 U9005 ( .A(n10154), .ZN(n10155) );
  INV_X1 U9006 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10157) );
  NAND3_X1 U9007 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .A3(P2_ADDR_REG_0__SCAN_IN), .ZN(n10156) );
  NAND2_X1 U9008 ( .A1(n10157), .A2(n10156), .ZN(n10153) );
  NAND2_X1 U9009 ( .A1(n10155), .A2(n10153), .ZN(n10203) );
  NAND2_X1 U9010 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n7291) );
  OAI21_X1 U9011 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(P1_ADDR_REG_2__SCAN_IN), 
        .A(n7291), .ZN(n10202) );
  NOR2_X1 U9012 ( .A1(n10203), .A2(n10202), .ZN(n10201) );
  AOI21_X1 U9013 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(P2_ADDR_REG_2__SCAN_IN), 
        .A(n10201), .ZN(n10206) );
  NAND2_X1 U9014 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7292) );
  OAI21_X1 U9015 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(P2_ADDR_REG_3__SCAN_IN), 
        .A(n7292), .ZN(n10205) );
  NOR2_X1 U9016 ( .A1(n10206), .A2(n10205), .ZN(n10204) );
  AOI21_X1 U9017 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(P1_ADDR_REG_3__SCAN_IN), 
        .A(n10204), .ZN(n10209) );
  NOR2_X1 U9018 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7293) );
  AOI21_X1 U9019 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(P1_ADDR_REG_4__SCAN_IN), 
        .A(n7293), .ZN(n10208) );
  NAND2_X1 U9020 ( .A1(n10209), .A2(n10208), .ZN(n10207) );
  OAI21_X1 U9021 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(P2_ADDR_REG_4__SCAN_IN), 
        .A(n10207), .ZN(n10187) );
  NAND2_X1 U9022 ( .A1(n10188), .A2(n10187), .ZN(n10186) );
  OAI21_X1 U9023 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(P1_ADDR_REG_5__SCAN_IN), 
        .A(n10186), .ZN(n10190) );
  NAND2_X1 U9024 ( .A1(n10191), .A2(n10190), .ZN(n10189) );
  OAI21_X1 U9025 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(P1_ADDR_REG_6__SCAN_IN), 
        .A(n10189), .ZN(n10196) );
  NAND2_X1 U9026 ( .A1(n10197), .A2(n10196), .ZN(n10195) );
  OAI21_X1 U9027 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(P1_ADDR_REG_7__SCAN_IN), 
        .A(n10195), .ZN(n10199) );
  NAND2_X1 U9028 ( .A1(n10200), .A2(n10199), .ZN(n10198) );
  OAI21_X1 U9029 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(P1_ADDR_REG_8__SCAN_IN), 
        .A(n10198), .ZN(n10193) );
  NAND2_X1 U9030 ( .A1(n10194), .A2(n10193), .ZN(n10192) );
  OAI21_X1 U9031 ( .B1(P2_ADDR_REG_9__SCAN_IN), .B2(P1_ADDR_REG_9__SCAN_IN), 
        .A(n10192), .ZN(n10184) );
  NAND2_X1 U9032 ( .A1(n10185), .A2(n10184), .ZN(n10183) );
  OAI21_X1 U9033 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10183), .ZN(n10181) );
  NAND2_X1 U9034 ( .A1(n10182), .A2(n10181), .ZN(n10180) );
  OAI21_X1 U9035 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10180), .ZN(n10178) );
  NAND2_X1 U9036 ( .A1(n10179), .A2(n10178), .ZN(n10177) );
  OAI21_X1 U9037 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10177), .ZN(n10175) );
  NAND2_X1 U9038 ( .A1(n10176), .A2(n10175), .ZN(n10174) );
  OAI21_X1 U9039 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10174), .ZN(n10172) );
  NAND2_X1 U9040 ( .A1(n10173), .A2(n10172), .ZN(n10171) );
  OAI21_X1 U9041 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10171), .ZN(n10169) );
  NAND2_X1 U9042 ( .A1(n10170), .A2(n10169), .ZN(n10168) );
  OAI21_X1 U9043 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10168), .ZN(n10166) );
  NAND2_X1 U9044 ( .A1(n10167), .A2(n10166), .ZN(n10165) );
  OAI21_X1 U9045 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10165), .ZN(n10163) );
  NAND2_X1 U9046 ( .A1(n10164), .A2(n10163), .ZN(n10162) );
  OAI21_X1 U9047 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10162), .ZN(n10160) );
  NOR2_X1 U9048 ( .A1(n10159), .A2(n10160), .ZN(n7294) );
  NAND2_X1 U9049 ( .A1(n10159), .A2(n10160), .ZN(n10158) );
  OAI21_X1 U9050 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n7294), .A(n10158), .ZN(
        n7296) );
  XNOR2_X1 U9051 ( .A(n4541), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n7295) );
  XNOR2_X1 U9052 ( .A(n7296), .B(n7295), .ZN(ADD_1068_U4) );
  NAND2_X1 U9053 ( .A1(n8719), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n7297) );
  OAI21_X1 U9054 ( .B1(n8374), .B2(n8719), .A(n7297), .ZN(P2_U3521) );
  XOR2_X1 U9055 ( .A(n7298), .B(n9384), .Z(n7300) );
  AOI21_X1 U9056 ( .B1(n7300), .B2(n9698), .A(n7299), .ZN(n9979) );
  XNOR2_X1 U9057 ( .A(n7301), .B(n9384), .ZN(n9982) );
  NAND2_X1 U9058 ( .A1(n7303), .A2(n7302), .ZN(n7304) );
  AND2_X1 U9059 ( .A1(n7318), .A2(n7304), .ZN(n9975) );
  NAND2_X1 U9060 ( .A1(n7305), .A2(n9975), .ZN(n7308) );
  AOI22_X1 U9061 ( .A1(n4334), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n9951), .B2(
        n7306), .ZN(n7307) );
  OAI211_X1 U9062 ( .C1(n9976), .C2(n9716), .A(n7308), .B(n7307), .ZN(n7309)
         );
  AOI21_X1 U9063 ( .B1(n9721), .B2(n9982), .A(n7309), .ZN(n7310) );
  OAI21_X1 U9064 ( .B1(n4334), .B2(n9979), .A(n7310), .ZN(P1_U3290) );
  INV_X1 U9065 ( .A(n7316), .ZN(n9381) );
  XNOR2_X1 U9066 ( .A(n7311), .B(n9381), .ZN(n7314) );
  INV_X1 U9067 ( .A(n7312), .ZN(n7313) );
  AOI21_X1 U9068 ( .B1(n7314), .B2(n9698), .A(n7313), .ZN(n9986) );
  XNOR2_X1 U9069 ( .A(n7315), .B(n7316), .ZN(n9989) );
  NAND2_X1 U9070 ( .A1(n7318), .A2(n7317), .ZN(n7319) );
  NAND2_X1 U9071 ( .A1(n7319), .A2(n9957), .ZN(n7320) );
  NOR2_X1 U9072 ( .A1(n7321), .A2(n7320), .ZN(n9983) );
  NAND2_X1 U9073 ( .A1(n9960), .A2(n9983), .ZN(n7325) );
  NOR2_X1 U9074 ( .A1(n9727), .A2(n7322), .ZN(n7323) );
  AOI21_X1 U9075 ( .B1(n4334), .B2(P1_REG2_REG_4__SCAN_IN), .A(n7323), .ZN(
        n7324) );
  OAI211_X1 U9076 ( .C1(n9985), .C2(n9716), .A(n7325), .B(n7324), .ZN(n7326)
         );
  AOI21_X1 U9077 ( .B1(n9721), .B2(n9989), .A(n7326), .ZN(n7327) );
  OAI21_X1 U9078 ( .B1(n9986), .B2(n4334), .A(n7327), .ZN(P1_U3289) );
  INV_X1 U9079 ( .A(n7328), .ZN(n7329) );
  OAI21_X1 U9080 ( .B1(n7329), .B2(n4688), .A(n7435), .ZN(n7332) );
  NAND2_X1 U9081 ( .A1(n9461), .A2(n9291), .ZN(n7331) );
  NAND2_X1 U9082 ( .A1(n9459), .A2(n9169), .ZN(n7330) );
  NAND2_X1 U9083 ( .A1(n7331), .A2(n7330), .ZN(n9860) );
  AOI21_X1 U9084 ( .B1(n7332), .B2(n9698), .A(n9860), .ZN(n10025) );
  XNOR2_X1 U9085 ( .A(n7333), .B(n7334), .ZN(n10028) );
  NAND2_X1 U9086 ( .A1(n10028), .A2(n9721), .ZN(n7340) );
  OAI22_X1 U9087 ( .A1(n9723), .A2(n7335), .B1(n9869), .B2(n9727), .ZN(n7337)
         );
  OAI211_X1 U9088 ( .C1(n7421), .C2(n10026), .A(n7444), .B(n9957), .ZN(n10024)
         );
  NOR2_X1 U9089 ( .A1(n10024), .A2(n9671), .ZN(n7336) );
  AOI211_X1 U9090 ( .C1(n9953), .C2(n7338), .A(n7337), .B(n7336), .ZN(n7339)
         );
  OAI211_X1 U9091 ( .C1(n10025), .C2(n4334), .A(n7340), .B(n7339), .ZN(
        P1_U3283) );
  INV_X1 U9092 ( .A(n9937), .ZN(n7354) );
  AOI22_X1 U9093 ( .A1(n7585), .A2(P1_REG1_REG_12__SCAN_IN), .B1(n5197), .B2(
        n7355), .ZN(n7342) );
  OAI21_X1 U9094 ( .B1(n7343), .B2(n7342), .A(n7584), .ZN(n7350) );
  NOR2_X1 U9095 ( .A1(n7585), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n7344) );
  AOI21_X1 U9096 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n7585), .A(n7344), .ZN(
        n7348) );
  OAI21_X1 U9097 ( .B1(n7348), .B2(n7347), .A(n7580), .ZN(n7349) );
  AOI22_X1 U9098 ( .A1(n9939), .A2(n7350), .B1(n9915), .B2(n7349), .ZN(n7353)
         );
  NAND2_X1 U9099 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n7970) );
  INV_X1 U9100 ( .A(n7970), .ZN(n7351) );
  AOI21_X1 U9101 ( .B1(n9933), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n7351), .ZN(
        n7352) );
  OAI211_X1 U9102 ( .C1(n7355), .C2(n7354), .A(n7353), .B(n7352), .ZN(P1_U3255) );
  INV_X1 U9103 ( .A(n7356), .ZN(n7413) );
  OAI222_X1 U9104 ( .A1(n8159), .A2(n7413), .B1(n8186), .B2(n7357), .C1(n8568), 
        .C2(P2_U3151), .ZN(P2_U3275) );
  NAND2_X1 U9105 ( .A1(n7360), .A2(n7359), .ZN(n9204) );
  NOR2_X1 U9106 ( .A1(n7362), .A2(n7361), .ZN(n7417) );
  INV_X1 U9107 ( .A(n7362), .ZN(n7365) );
  INV_X1 U9108 ( .A(n7377), .ZN(n7363) );
  AOI21_X1 U9109 ( .B1(n7365), .B2(n7364), .A(n7363), .ZN(n7366) );
  AOI211_X1 U9110 ( .C1(n7417), .C2(n7415), .A(n9945), .B(n7366), .ZN(n7369)
         );
  NAND2_X1 U9111 ( .A1(n9463), .A2(n9291), .ZN(n7368) );
  NAND2_X1 U9112 ( .A1(n9461), .A2(n9181), .ZN(n7367) );
  NAND2_X1 U9113 ( .A1(n7368), .A2(n7367), .ZN(n7491) );
  NOR2_X1 U9114 ( .A1(n7369), .A2(n7491), .ZN(n10012) );
  INV_X1 U9115 ( .A(n7370), .ZN(n9956) );
  AOI21_X1 U9116 ( .B1(n9956), .B2(n7495), .A(n9977), .ZN(n7371) );
  NAND2_X1 U9117 ( .A1(n7371), .A2(n7422), .ZN(n10011) );
  INV_X1 U9118 ( .A(n10011), .ZN(n7375) );
  INV_X1 U9119 ( .A(n7495), .ZN(n10013) );
  NOR2_X1 U9120 ( .A1(n9727), .A2(n7493), .ZN(n7372) );
  AOI21_X1 U9121 ( .B1(n4334), .B2(P1_REG2_REG_8__SCAN_IN), .A(n7372), .ZN(
        n7373) );
  OAI21_X1 U9122 ( .B1(n9716), .B2(n10013), .A(n7373), .ZN(n7374) );
  AOI21_X1 U9123 ( .B1(n7375), .B2(n9960), .A(n7374), .ZN(n7379) );
  XOR2_X1 U9124 ( .A(n7376), .B(n7377), .Z(n10010) );
  INV_X1 U9125 ( .A(n10010), .ZN(n10016) );
  NAND2_X1 U9126 ( .A1(n10016), .A2(n9721), .ZN(n7378) );
  OAI211_X1 U9127 ( .C1(n10012), .C2(n4334), .A(n7379), .B(n7378), .ZN(
        P1_U3285) );
  INV_X1 U9128 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n10148) );
  NAND2_X1 U9129 ( .A1(n7395), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n7380) );
  NOR2_X1 U9130 ( .A1(n10148), .A2(n7382), .ZN(n7499) );
  AOI21_X1 U9131 ( .B1(n10148), .B2(n7382), .A(n7499), .ZN(n7405) );
  INV_X1 U9132 ( .A(n7383), .ZN(n7389) );
  INV_X1 U9133 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7384) );
  MUX2_X1 U9134 ( .A(n10148), .B(n7384), .S(n8748), .Z(n7385) );
  NAND2_X1 U9135 ( .A1(n7385), .A2(n7519), .ZN(n7511) );
  INV_X1 U9136 ( .A(n7385), .ZN(n7386) );
  NAND2_X1 U9137 ( .A1(n7386), .A2(n7398), .ZN(n7387) );
  AND2_X1 U9138 ( .A1(n7511), .A2(n7387), .ZN(n7388) );
  OAI21_X1 U9139 ( .B1(n7390), .B2(n7389), .A(n7388), .ZN(n7512) );
  INV_X1 U9140 ( .A(n7512), .ZN(n7392) );
  NOR3_X1 U9141 ( .A1(n7390), .A2(n7389), .A3(n7388), .ZN(n7391) );
  OAI21_X1 U9142 ( .B1(n7392), .B2(n7391), .A(n8763), .ZN(n7404) );
  INV_X1 U9143 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n7394) );
  AND2_X1 U9144 ( .A1(P2_U3151), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n7848) );
  INV_X1 U9145 ( .A(n7848), .ZN(n7393) );
  OAI21_X1 U9146 ( .B1(n8724), .B2(n7394), .A(n7393), .ZN(n7402) );
  NAND2_X1 U9147 ( .A1(n7395), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n7396) );
  AOI21_X1 U9148 ( .B1(n7384), .B2(n7399), .A(n7521), .ZN(n7400) );
  NOR2_X1 U9149 ( .A1(n7400), .A2(n8756), .ZN(n7401) );
  AOI211_X1 U9150 ( .C1(n8699), .C2(n7519), .A(n7402), .B(n7401), .ZN(n7403)
         );
  OAI211_X1 U9151 ( .C1(n7405), .C2(n8766), .A(n7404), .B(n7403), .ZN(P2_U3193) );
  INV_X1 U9152 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n7412) );
  NAND2_X1 U9153 ( .A1(n5983), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n7408) );
  NAND2_X1 U9154 ( .A1(n6359), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n7407) );
  NAND2_X1 U9155 ( .A1(n5973), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n7406) );
  AND3_X1 U9156 ( .A1(n7408), .A2(n7407), .A3(n7406), .ZN(n7409) );
  INV_X1 U9157 ( .A(n8769), .ZN(n8582) );
  NAND2_X1 U9158 ( .A1(n8582), .A2(P2_U3893), .ZN(n7411) );
  OAI21_X1 U9159 ( .B1(P2_U3893), .B2(n7412), .A(n7411), .ZN(P2_U3522) );
  OAI222_X1 U9160 ( .A1(n9298), .A2(P1_U3086), .B1(n8191), .B2(n7414), .C1(
        n7413), .C2(n7965), .ZN(P1_U3335) );
  INV_X1 U9161 ( .A(n7415), .ZN(n7416) );
  XOR2_X1 U9162 ( .A(n9391), .B(n9203), .Z(n7419) );
  NOR2_X1 U9163 ( .A1(n7418), .A2(n9106), .ZN(n7538) );
  AOI21_X1 U9164 ( .B1(n7419), .B2(n9698), .A(n7538), .ZN(n10020) );
  XNOR2_X1 U9165 ( .A(n7420), .B(n9391), .ZN(n10023) );
  AOI211_X1 U9166 ( .C1(n10017), .C2(n7422), .A(n9977), .B(n7421), .ZN(n7423)
         );
  AND2_X1 U9167 ( .A1(n9169), .A2(n9460), .ZN(n7539) );
  NOR2_X1 U9168 ( .A1(n7423), .A2(n7539), .ZN(n10018) );
  OAI22_X1 U9169 ( .A1(n9723), .A2(n7424), .B1(n7542), .B2(n9727), .ZN(n7425)
         );
  AOI21_X1 U9170 ( .B1(n9953), .B2(n10017), .A(n7425), .ZN(n7426) );
  OAI21_X1 U9171 ( .B1(n10018), .B2(n9671), .A(n7426), .ZN(n7427) );
  AOI21_X1 U9172 ( .B1(n9721), .B2(n10023), .A(n7427), .ZN(n7428) );
  OAI21_X1 U9173 ( .B1(n10020), .B2(n4334), .A(n7428), .ZN(P1_U3284) );
  INV_X1 U9174 ( .A(n7430), .ZN(n7431) );
  OR2_X1 U9175 ( .A1(n7432), .A2(n7431), .ZN(n9392) );
  INV_X1 U9176 ( .A(n9392), .ZN(n7433) );
  XNOR2_X1 U9177 ( .A(n7429), .B(n7433), .ZN(n10034) );
  INV_X1 U9178 ( .A(n7434), .ZN(n10046) );
  NAND2_X1 U9179 ( .A1(n7435), .A2(n9215), .ZN(n7436) );
  XNOR2_X1 U9180 ( .A(n7436), .B(n9392), .ZN(n7437) );
  NAND2_X1 U9181 ( .A1(n7437), .A2(n9698), .ZN(n7441) );
  NAND2_X1 U9182 ( .A1(n9458), .A2(n9181), .ZN(n7439) );
  NAND2_X1 U9183 ( .A1(n9460), .A2(n9291), .ZN(n7438) );
  NAND2_X1 U9184 ( .A1(n7439), .A2(n7438), .ZN(n7812) );
  INV_X1 U9185 ( .A(n7812), .ZN(n7440) );
  NAND2_X1 U9186 ( .A1(n7441), .A2(n7440), .ZN(n7442) );
  AOI21_X1 U9187 ( .B1(n10034), .B2(n10046), .A(n7442), .ZN(n10036) );
  INV_X1 U9188 ( .A(n7443), .ZN(n9961) );
  AOI21_X1 U9189 ( .B1(n7444), .B2(n7802), .A(n9977), .ZN(n7445) );
  NAND2_X1 U9190 ( .A1(n7445), .A2(n7553), .ZN(n10030) );
  OAI22_X1 U9191 ( .A1(n9723), .A2(n7446), .B1(n7809), .B2(n9727), .ZN(n7447)
         );
  AOI21_X1 U9192 ( .B1(n7802), .B2(n9953), .A(n7447), .ZN(n7448) );
  OAI21_X1 U9193 ( .B1(n10030), .B2(n9671), .A(n7448), .ZN(n7449) );
  AOI21_X1 U9194 ( .B1(n10034), .B2(n9961), .A(n7449), .ZN(n7450) );
  OAI21_X1 U9195 ( .B1(n10036), .B2(n4334), .A(n7450), .ZN(P1_U3282) );
  XNOR2_X1 U9196 ( .A(n7796), .B(n8600), .ZN(n8389) );
  XNOR2_X1 U9197 ( .A(n7451), .B(n8389), .ZN(n10117) );
  XOR2_X1 U9198 ( .A(n7452), .B(n8389), .Z(n7453) );
  NAND2_X1 U9199 ( .A1(n7453), .A2(n8895), .ZN(n7455) );
  AOI22_X1 U9200 ( .A1(n8898), .A2(n8601), .B1(n8599), .B2(n8899), .ZN(n7454)
         );
  OAI211_X1 U9201 ( .C1(n10107), .C2(n10117), .A(n7455), .B(n7454), .ZN(n10119) );
  NAND2_X1 U9202 ( .A1(n10119), .A2(n8915), .ZN(n7460) );
  INV_X1 U9203 ( .A(n7456), .ZN(n7789) );
  OAI22_X1 U9204 ( .A1(n8915), .A2(n7457), .B1(n7789), .B2(n8770), .ZN(n7458)
         );
  AOI21_X1 U9205 ( .B1(n8888), .B2(n7796), .A(n7458), .ZN(n7459) );
  OAI211_X1 U9206 ( .C1(n10117), .C2(n7461), .A(n7460), .B(n7459), .ZN(
        P2_U3223) );
  INV_X1 U9207 ( .A(n7468), .ZN(n10108) );
  NAND2_X1 U9208 ( .A1(n7462), .A2(n7463), .ZN(n7464) );
  XNOR2_X1 U9209 ( .A(n7578), .B(n8254), .ZN(n7466) );
  XNOR2_X1 U9210 ( .A(n7466), .B(n8602), .ZN(n7574) );
  AND2_X1 U9211 ( .A1(n7466), .A2(n7474), .ZN(n7467) );
  XNOR2_X1 U9212 ( .A(n7468), .B(n8200), .ZN(n7715) );
  XNOR2_X1 U9213 ( .A(n7715), .B(n8601), .ZN(n7469) );
  OAI211_X1 U9214 ( .C1(n7470), .C2(n7469), .A(n7714), .B(n8321), .ZN(n7478)
         );
  NOR2_X1 U9215 ( .A1(n8258), .A2(n7471), .ZN(n7476) );
  OR2_X1 U9216 ( .A1(n8349), .A2(n7717), .ZN(n7473) );
  OAI211_X1 U9217 ( .C1(n8317), .C2(n7474), .A(n7473), .B(n7472), .ZN(n7475)
         );
  NOR2_X1 U9218 ( .A1(n7476), .A2(n7475), .ZN(n7477) );
  OAI211_X1 U9219 ( .C1(n10108), .C2(n8329), .A(n7478), .B(n7477), .ZN(
        P2_U3171) );
  XNOR2_X1 U9220 ( .A(n10124), .B(n8599), .ZN(n8390) );
  XNOR2_X1 U9221 ( .A(n7479), .B(n8390), .ZN(n10121) );
  INV_X1 U9222 ( .A(n8390), .ZN(n7719) );
  XNOR2_X1 U9223 ( .A(n7480), .B(n7719), .ZN(n7481) );
  OAI222_X1 U9224 ( .A1(n8860), .A2(n8482), .B1(n8858), .B2(n7717), .C1(n8970), 
        .C2(n7481), .ZN(n10122) );
  NAND2_X1 U9225 ( .A1(n10122), .A2(n8915), .ZN(n7485) );
  INV_X1 U9226 ( .A(n7482), .ZN(n7849) );
  OAI22_X1 U9227 ( .A1(n8915), .A2(n7384), .B1(n7849), .B2(n8770), .ZN(n7483)
         );
  AOI21_X1 U9228 ( .B1(n10124), .B2(n8888), .A(n7483), .ZN(n7484) );
  OAI211_X1 U9229 ( .C1(n10121), .C2(n8891), .A(n7485), .B(n7484), .ZN(
        P2_U3222) );
  INV_X1 U9230 ( .A(n7486), .ZN(n7488) );
  NAND2_X1 U9231 ( .A1(n7488), .A2(n7487), .ZN(n7490) );
  XNOR2_X1 U9232 ( .A(n7490), .B(n7489), .ZN(n7497) );
  AOI22_X1 U9233 ( .A1(n9861), .A2(n7491), .B1(P1_REG3_REG_8__SCAN_IN), .B2(
        P1_U3086), .ZN(n7492) );
  OAI21_X1 U9234 ( .B1(n7493), .B2(n9868), .A(n7492), .ZN(n7494) );
  AOI21_X1 U9235 ( .B1(n7495), .B2(n9186), .A(n7494), .ZN(n7496) );
  OAI21_X1 U9236 ( .B1(n7497), .B2(n9188), .A(n7496), .ZN(P1_U3221) );
  NOR2_X1 U9237 ( .A1(n7519), .A2(n7498), .ZN(n7500) );
  NOR2_X1 U9238 ( .A1(n7500), .A2(n7499), .ZN(n7504) );
  INV_X1 U9239 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7505) );
  OR2_X1 U9240 ( .A1(n7528), .A2(n7505), .ZN(n7599) );
  NAND2_X1 U9241 ( .A1(n7528), .A2(n7505), .ZN(n7501) );
  NAND2_X1 U9242 ( .A1(n7599), .A2(n7501), .ZN(n7503) );
  INV_X1 U9243 ( .A(n7600), .ZN(n7502) );
  AOI21_X1 U9244 ( .B1(n7504), .B2(n7503), .A(n7502), .ZN(n7531) );
  INV_X1 U9245 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7624) );
  MUX2_X1 U9246 ( .A(n7505), .B(n7624), .S(n8748), .Z(n7506) );
  NAND2_X1 U9247 ( .A1(n7506), .A2(n7528), .ZN(n7603) );
  INV_X1 U9248 ( .A(n7506), .ZN(n7508) );
  NAND2_X1 U9249 ( .A1(n7508), .A2(n7507), .ZN(n7509) );
  NAND2_X1 U9250 ( .A1(n7603), .A2(n7509), .ZN(n7510) );
  AOI21_X1 U9251 ( .B1(n7512), .B2(n7511), .A(n7510), .ZN(n7610) );
  AND3_X1 U9252 ( .A1(n7512), .A2(n7511), .A3(n7510), .ZN(n7513) );
  OAI21_X1 U9253 ( .B1(n7610), .B2(n7513), .A(n8763), .ZN(n7530) );
  INV_X1 U9254 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7516) );
  INV_X1 U9255 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n7514) );
  NOR2_X1 U9256 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7514), .ZN(n7710) );
  INV_X1 U9257 ( .A(n7710), .ZN(n7515) );
  OAI21_X1 U9258 ( .B1(n8724), .B2(n7516), .A(n7515), .ZN(n7527) );
  NOR2_X1 U9259 ( .A1(n7519), .A2(n7518), .ZN(n7520) );
  OR2_X1 U9260 ( .A1(n7528), .A2(n7624), .ZN(n7614) );
  NAND2_X1 U9261 ( .A1(n7528), .A2(n7624), .ZN(n7522) );
  NAND2_X1 U9262 ( .A1(n7614), .A2(n7522), .ZN(n7523) );
  NAND2_X1 U9263 ( .A1(n7524), .A2(n7523), .ZN(n7525) );
  AOI21_X1 U9264 ( .B1(n7615), .B2(n7525), .A(n8756), .ZN(n7526) );
  AOI211_X1 U9265 ( .C1(n8699), .C2(n7528), .A(n7527), .B(n7526), .ZN(n7529)
         );
  OAI211_X1 U9266 ( .C1(n7531), .C2(n8766), .A(n7530), .B(n7529), .ZN(P2_U3194) );
  INV_X1 U9267 ( .A(n7532), .ZN(n8189) );
  OAI222_X1 U9268 ( .A1(n9058), .A2(n8189), .B1(P2_U3151), .B2(n7534), .C1(
        n7533), .C2(n8186), .ZN(P2_U3274) );
  AOI21_X1 U9269 ( .B1(n7537), .B2(n7536), .A(n7535), .ZN(n7545) );
  OAI21_X1 U9270 ( .B1(n7539), .B2(n7538), .A(n9861), .ZN(n7541) );
  OAI211_X1 U9271 ( .C1(n9868), .C2(n7542), .A(n7541), .B(n7540), .ZN(n7543)
         );
  AOI21_X1 U9272 ( .B1(n10017), .B2(n9186), .A(n7543), .ZN(n7544) );
  OAI21_X1 U9273 ( .B1(n7545), .B2(n9188), .A(n7544), .ZN(P1_U3231) );
  OAI211_X1 U9274 ( .C1(n7547), .C2(n9394), .A(n7546), .B(n9698), .ZN(n7551)
         );
  NAND2_X1 U9275 ( .A1(n9457), .A2(n9169), .ZN(n7549) );
  NAND2_X1 U9276 ( .A1(n9459), .A2(n9291), .ZN(n7548) );
  NAND2_X1 U9277 ( .A1(n7549), .A2(n7548), .ZN(n7969) );
  INV_X1 U9278 ( .A(n7969), .ZN(n7550) );
  NAND2_X1 U9279 ( .A1(n7551), .A2(n7550), .ZN(n7561) );
  INV_X1 U9280 ( .A(n7561), .ZN(n7560) );
  XNOR2_X1 U9281 ( .A(n7552), .B(n9394), .ZN(n7563) );
  NAND2_X1 U9282 ( .A1(n7563), .A2(n9721), .ZN(n7559) );
  AOI211_X1 U9283 ( .C1(n7979), .C2(n7553), .A(n9977), .B(n7633), .ZN(n7562)
         );
  INV_X1 U9284 ( .A(n7979), .ZN(n7554) );
  NOR2_X1 U9285 ( .A1(n7554), .A2(n9716), .ZN(n7557) );
  OAI22_X1 U9286 ( .A1(n9723), .A2(n7555), .B1(n7972), .B2(n9727), .ZN(n7556)
         );
  AOI211_X1 U9287 ( .C1(n7562), .C2(n9960), .A(n7557), .B(n7556), .ZN(n7558)
         );
  OAI211_X1 U9288 ( .C1(n4334), .C2(n7560), .A(n7559), .B(n7558), .ZN(P1_U3281) );
  AOI211_X1 U9289 ( .C1(n7563), .C2(n10029), .A(n7562), .B(n7561), .ZN(n7568)
         );
  INV_X1 U9290 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n7564) );
  NOR2_X1 U9291 ( .A1(n10049), .A2(n7564), .ZN(n7565) );
  AOI21_X1 U9292 ( .B1(n7979), .B2(n9832), .A(n7565), .ZN(n7566) );
  OAI21_X1 U9293 ( .B1(n7568), .B2(n10047), .A(n7566), .ZN(P1_U3489) );
  AOI22_X1 U9294 ( .A1(n7979), .A2(n9777), .B1(n10066), .B2(
        P1_REG1_REG_12__SCAN_IN), .ZN(n7567) );
  OAI21_X1 U9295 ( .B1(n7568), .B2(n10066), .A(n7567), .ZN(P1_U3534) );
  INV_X1 U9296 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n7569) );
  NOR2_X1 U9297 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7569), .ZN(n8618) );
  AOI21_X1 U9298 ( .B1(n8345), .B2(n8603), .A(n8618), .ZN(n7571) );
  OR2_X1 U9299 ( .A1(n8349), .A2(n7716), .ZN(n7570) );
  OAI211_X1 U9300 ( .C1(n7572), .C2(n8258), .A(n7571), .B(n7570), .ZN(n7577)
         );
  XOR2_X1 U9301 ( .A(n7574), .B(n7573), .Z(n7575) );
  NOR2_X1 U9302 ( .A1(n7575), .A2(n8353), .ZN(n7576) );
  AOI211_X1 U9303 ( .C1(n7578), .C2(n8351), .A(n7577), .B(n7576), .ZN(n7579)
         );
  INV_X1 U9304 ( .A(n7579), .ZN(P2_U3161) );
  NAND2_X1 U9305 ( .A1(n7682), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n7581) );
  OAI21_X1 U9306 ( .B1(n7682), .B2(P1_REG2_REG_13__SCAN_IN), .A(n7581), .ZN(
        n7582) );
  NOR2_X1 U9307 ( .A1(n7582), .A2(n7583), .ZN(n7675) );
  AOI211_X1 U9308 ( .C1(n7583), .C2(n7582), .A(n7675), .B(n9928), .ZN(n7594)
         );
  OAI21_X1 U9309 ( .B1(n7585), .B2(P1_REG1_REG_12__SCAN_IN), .A(n7584), .ZN(
        n7588) );
  INV_X1 U9310 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n7586) );
  MUX2_X1 U9311 ( .A(n7586), .B(P1_REG1_REG_13__SCAN_IN), .S(n7682), .Z(n7587)
         );
  NOR2_X1 U9312 ( .A1(n7587), .A2(n7588), .ZN(n7681) );
  AOI211_X1 U9313 ( .C1(n7588), .C2(n7587), .A(n7681), .B(n9919), .ZN(n7593)
         );
  INV_X1 U9314 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n7591) );
  NAND2_X1 U9315 ( .A1(n9937), .A2(n7682), .ZN(n7590) );
  AND2_X1 U9316 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n7898) );
  INV_X1 U9317 ( .A(n7898), .ZN(n7589) );
  OAI211_X1 U9318 ( .C1(n7591), .C2(n9553), .A(n7590), .B(n7589), .ZN(n7592)
         );
  OR3_X1 U9319 ( .A1(n7594), .A2(n7593), .A3(n7592), .ZN(P1_U3256) );
  INV_X1 U9320 ( .A(n7595), .ZN(n7598) );
  AOI22_X1 U9321 ( .A1(n9296), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n6448), .ZN(n7596) );
  OAI21_X1 U9322 ( .B1(n7598), .B2(n7965), .A(n7596), .ZN(P1_U3333) );
  OAI222_X1 U9323 ( .A1(n8186), .A2(n8076), .B1(n8159), .B2(n7598), .C1(n7597), 
        .C2(P2_U3151), .ZN(P2_U3273) );
  INV_X1 U9324 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n7668) );
  AOI21_X1 U9325 ( .B1(n7668), .B2(n7601), .A(n7729), .ZN(n7621) );
  INV_X1 U9326 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n7602) );
  OAI22_X1 U9327 ( .A1(n8724), .A2(n7602), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6097), .ZN(n7613) );
  INV_X1 U9328 ( .A(n7603), .ZN(n7609) );
  INV_X1 U9329 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n7604) );
  MUX2_X1 U9330 ( .A(n7668), .B(n7604), .S(n8748), .Z(n7605) );
  NAND2_X1 U9331 ( .A1(n7605), .A2(n7751), .ZN(n7742) );
  INV_X1 U9332 ( .A(n7605), .ZN(n7606) );
  NAND2_X1 U9333 ( .A1(n7606), .A2(n7616), .ZN(n7607) );
  AND2_X1 U9334 ( .A1(n7742), .A2(n7607), .ZN(n7608) );
  OAI21_X1 U9335 ( .B1(n7610), .B2(n7609), .A(n7608), .ZN(n7743) );
  OR3_X1 U9336 ( .A1(n7610), .A2(n7609), .A3(n7608), .ZN(n7611) );
  AOI21_X1 U9337 ( .B1(n7743), .B2(n7611), .A(n8695), .ZN(n7612) );
  AOI211_X1 U9338 ( .C1(n8699), .C2(n7751), .A(n7613), .B(n7612), .ZN(n7620)
         );
  AOI21_X1 U9339 ( .B1(n7604), .B2(n7617), .A(n7752), .ZN(n7618) );
  OR2_X1 U9340 ( .A1(n7618), .A2(n8756), .ZN(n7619) );
  OAI211_X1 U9341 ( .C1(n7621), .C2(n8766), .A(n7620), .B(n7619), .ZN(P2_U3195) );
  XNOR2_X1 U9342 ( .A(n7660), .B(n8377), .ZN(n7622) );
  OAI222_X1 U9343 ( .A1(n8858), .A2(n7792), .B1(n8860), .B2(n4882), .C1(n7622), 
        .C2(n8970), .ZN(n10129) );
  INV_X1 U9344 ( .A(n10129), .ZN(n7630) );
  INV_X1 U9345 ( .A(n7623), .ZN(n7713) );
  OAI22_X1 U9346 ( .A1(n8915), .A2(n7624), .B1(n7713), .B2(n8770), .ZN(n7628)
         );
  NOR2_X1 U9347 ( .A1(n7625), .A2(n8377), .ZN(n10128) );
  INV_X1 U9348 ( .A(n7626), .ZN(n10127) );
  NOR3_X1 U9349 ( .A1(n10128), .A2(n10127), .A3(n8891), .ZN(n7627) );
  AOI211_X1 U9350 ( .C1(n8888), .C2(n10131), .A(n7628), .B(n7627), .ZN(n7629)
         );
  OAI21_X1 U9351 ( .B1(n8909), .B2(n7630), .A(n7629), .ZN(P2_U3221) );
  OAI21_X1 U9352 ( .B1(n7632), .B2(n9396), .A(n7631), .ZN(n9722) );
  OAI21_X1 U9353 ( .B1(n7633), .B2(n7902), .A(n9957), .ZN(n7634) );
  NOR2_X1 U9354 ( .A1(n7634), .A2(n7699), .ZN(n9730) );
  XOR2_X1 U9355 ( .A(n7635), .B(n9396), .Z(n7639) );
  OAI22_X1 U9356 ( .A1(n7637), .A2(n9096), .B1(n7636), .B2(n9106), .ZN(n7899)
         );
  INV_X1 U9357 ( .A(n7899), .ZN(n7638) );
  OAI21_X1 U9358 ( .B1(n7639), .B2(n9945), .A(n7638), .ZN(n9724) );
  AOI211_X1 U9359 ( .C1(n10029), .C2(n9722), .A(n9730), .B(n9724), .ZN(n7643)
         );
  AOI22_X1 U9360 ( .A1(n9729), .A2(n9777), .B1(n10066), .B2(
        P1_REG1_REG_13__SCAN_IN), .ZN(n7640) );
  OAI21_X1 U9361 ( .B1(n7643), .B2(n10066), .A(n7640), .ZN(P1_U3535) );
  INV_X1 U9362 ( .A(n9832), .ZN(n9840) );
  OAI22_X1 U9363 ( .A1(n7902), .A2(n9840), .B1(n10049), .B2(n5225), .ZN(n7641)
         );
  INV_X1 U9364 ( .A(n7641), .ZN(n7642) );
  OAI21_X1 U9365 ( .B1(n7643), .B2(n10047), .A(n7642), .ZN(P1_U3492) );
  INV_X1 U9366 ( .A(n7644), .ZN(n7649) );
  NAND2_X1 U9367 ( .A1(n6448), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n7646) );
  OR2_X1 U9368 ( .A1(n7645), .A2(P1_U3086), .ZN(n9416) );
  OAI211_X1 U9369 ( .C1(n7649), .C2(n7965), .A(n7646), .B(n9416), .ZN(P1_U3332) );
  OR2_X1 U9370 ( .A1(n7647), .A2(P2_U3151), .ZN(n8590) );
  NAND2_X1 U9371 ( .A1(n9056), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n7648) );
  OAI211_X1 U9372 ( .C1(n7649), .C2(n9058), .A(n8590), .B(n7648), .ZN(P2_U3272) );
  INV_X1 U9373 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n7653) );
  INV_X1 U9374 ( .A(n7650), .ZN(n8497) );
  OR2_X1 U9375 ( .A1(n8498), .A2(n8497), .ZN(n8495) );
  XNOR2_X1 U9376 ( .A(n7651), .B(n8495), .ZN(n7652) );
  AOI222_X1 U9377 ( .A1(n8895), .A2(n7652), .B1(n8595), .B2(n8899), .C1(n8597), 
        .C2(n8898), .ZN(n7782) );
  MUX2_X1 U9378 ( .A(n7653), .B(n7782), .S(n10133), .Z(n7656) );
  XNOR2_X1 U9379 ( .A(n7654), .B(n8495), .ZN(n7785) );
  INV_X1 U9380 ( .A(n10091), .ZN(n10126) );
  OR2_X1 U9381 ( .A1(n10135), .A2(n10126), .ZN(n9046) );
  INV_X1 U9382 ( .A(n9046), .ZN(n9034) );
  AOI22_X1 U9383 ( .A1(n7785), .A2(n9034), .B1(n9033), .B2(n7909), .ZN(n7655)
         );
  NAND2_X1 U9384 ( .A1(n7656), .A2(n7655), .ZN(P2_U3432) );
  INV_X1 U9385 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n7737) );
  MUX2_X1 U9386 ( .A(n7737), .B(n7782), .S(n10152), .Z(n7658) );
  NAND2_X1 U9387 ( .A1(n10152), .A2(n10091), .ZN(n8963) );
  INV_X1 U9388 ( .A(n8963), .ZN(n8949) );
  AOI22_X1 U9389 ( .A1(n7785), .A2(n8949), .B1(n8948), .B2(n7909), .ZN(n7657)
         );
  NAND2_X1 U9390 ( .A1(n7658), .A2(n7657), .ZN(P2_U3473) );
  OR2_X1 U9391 ( .A1(n7660), .A2(n7659), .ZN(n7663) );
  AND2_X1 U9392 ( .A1(n7663), .A2(n7661), .ZN(n7666) );
  NAND2_X1 U9393 ( .A1(n7663), .A2(n7662), .ZN(n7664) );
  OAI21_X1 U9394 ( .B1(n7666), .B2(n7665), .A(n7664), .ZN(n7667) );
  AOI222_X1 U9395 ( .A1(n8895), .A2(n7667), .B1(n8598), .B2(n8898), .C1(n8596), 
        .C2(n8899), .ZN(n7704) );
  MUX2_X1 U9396 ( .A(n7668), .B(n7704), .S(n10152), .Z(n7671) );
  XOR2_X1 U9397 ( .A(n7669), .B(n8392), .Z(n7707) );
  AOI22_X1 U9398 ( .A1(n7707), .A2(n8949), .B1(n8948), .B2(n8488), .ZN(n7670)
         );
  NAND2_X1 U9399 ( .A1(n7671), .A2(n7670), .ZN(P2_U3472) );
  INV_X1 U9400 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n7672) );
  MUX2_X1 U9401 ( .A(n7672), .B(n7704), .S(n10133), .Z(n7674) );
  AOI22_X1 U9402 ( .A1(n7707), .A2(n9034), .B1(n9033), .B2(n8488), .ZN(n7673)
         );
  NAND2_X1 U9403 ( .A1(n7674), .A2(n7673), .ZN(P2_U3429) );
  AOI22_X1 U9404 ( .A1(n9487), .A2(n7698), .B1(P1_REG2_REG_14__SCAN_IN), .B2(
        n7676), .ZN(n7677) );
  NOR2_X1 U9405 ( .A1(n7678), .A2(n7677), .ZN(n9482) );
  AOI211_X1 U9406 ( .C1(n7678), .C2(n7677), .A(n9482), .B(n9928), .ZN(n7690)
         );
  NOR2_X1 U9407 ( .A1(n9487), .A2(n7679), .ZN(n7680) );
  AOI21_X1 U9408 ( .B1(n9487), .B2(n7679), .A(n7680), .ZN(n7684) );
  AOI211_X1 U9409 ( .C1(n7684), .C2(n7683), .A(n9486), .B(n9919), .ZN(n7689)
         );
  INV_X1 U9410 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n7687) );
  NAND2_X1 U9411 ( .A1(n9937), .A2(n9487), .ZN(n7686) );
  NAND2_X1 U9412 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n7685) );
  OAI211_X1 U9413 ( .C1(n7687), .C2(n9553), .A(n7686), .B(n7685), .ZN(n7688)
         );
  OR3_X1 U9414 ( .A1(n7690), .A2(n7689), .A3(n7688), .ZN(P1_U3257) );
  INV_X1 U9415 ( .A(n7691), .ZN(n7692) );
  AOI21_X1 U9416 ( .B1(n7692), .B2(n4845), .A(n9945), .ZN(n7696) );
  NAND2_X1 U9417 ( .A1(n9455), .A2(n9169), .ZN(n7694) );
  NAND2_X1 U9418 ( .A1(n9457), .A2(n9291), .ZN(n7693) );
  NAND2_X1 U9419 ( .A1(n7694), .A2(n7693), .ZN(n9072) );
  AOI21_X1 U9420 ( .B1(n7696), .B2(n7695), .A(n9072), .ZN(n10038) );
  XNOR2_X1 U9421 ( .A(n7697), .B(n9399), .ZN(n10042) );
  INV_X1 U9422 ( .A(n10042), .ZN(n10045) );
  NAND2_X1 U9423 ( .A1(n10045), .A2(n9721), .ZN(n7703) );
  OAI22_X1 U9424 ( .A1(n9723), .A2(n7698), .B1(n9074), .B2(n9727), .ZN(n7701)
         );
  OAI211_X1 U9425 ( .C1(n7699), .C2(n10040), .A(n9957), .B(n7772), .ZN(n10037)
         );
  NOR2_X1 U9426 ( .A1(n10037), .A2(n9671), .ZN(n7700) );
  AOI211_X1 U9427 ( .C1(n9953), .C2(n9076), .A(n7701), .B(n7700), .ZN(n7702)
         );
  OAI211_X1 U9428 ( .C1(n4334), .C2(n10038), .A(n7703), .B(n7702), .ZN(
        P1_U3279) );
  INV_X1 U9429 ( .A(n8488), .ZN(n7829) );
  NOR2_X1 U9430 ( .A1(n7829), .A2(n8835), .ZN(n7706) );
  INV_X1 U9431 ( .A(n7704), .ZN(n7705) );
  AOI211_X1 U9432 ( .C1(n8908), .C2(n7826), .A(n7706), .B(n7705), .ZN(n7709)
         );
  AOI22_X1 U9433 ( .A1(n7707), .A2(n8906), .B1(P2_REG2_REG_13__SCAN_IN), .B2(
        n8909), .ZN(n7708) );
  OAI21_X1 U9434 ( .B1(n7709), .B2(n8909), .A(n7708), .ZN(P2_U3220) );
  AOI21_X1 U9435 ( .B1(n8345), .B2(n8599), .A(n7710), .ZN(n7712) );
  OR2_X1 U9436 ( .A1(n8349), .A2(n4882), .ZN(n7711) );
  OAI211_X1 U9437 ( .C1(n7713), .C2(n8258), .A(n7712), .B(n7711), .ZN(n7727)
         );
  XNOR2_X1 U9438 ( .A(n7796), .B(n8254), .ZN(n7852) );
  XOR2_X1 U9439 ( .A(n8254), .B(n8390), .Z(n7856) );
  AOI21_X1 U9440 ( .B1(n7717), .B2(n7852), .A(n7856), .ZN(n7723) );
  NAND3_X1 U9441 ( .A1(n7796), .A2(n8227), .A3(n8600), .ZN(n7718) );
  OAI211_X1 U9442 ( .C1(n7792), .C2(n8227), .A(n7719), .B(n7718), .ZN(n7722)
         );
  INV_X1 U9443 ( .A(n7796), .ZN(n10115) );
  NAND3_X1 U9444 ( .A1(n10115), .A2(n8600), .A3(n8254), .ZN(n7720) );
  OAI211_X1 U9445 ( .C1(n7792), .C2(n8200), .A(n8390), .B(n7720), .ZN(n7721)
         );
  XNOR2_X1 U9446 ( .A(n10131), .B(n8200), .ZN(n7818) );
  XOR2_X1 U9447 ( .A(n8598), .B(n7818), .Z(n7724) );
  AOI211_X1 U9448 ( .C1(n10131), .C2(n8351), .A(n7727), .B(n7726), .ZN(n7728)
         );
  INV_X1 U9449 ( .A(n7728), .ZN(P2_U3164) );
  NOR2_X1 U9450 ( .A1(n7751), .A2(n4369), .ZN(n7730) );
  NAND2_X1 U9451 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n8652), .ZN(n7731) );
  OAI21_X1 U9452 ( .B1(P2_REG1_REG_14__SCAN_IN), .B2(n8652), .A(n7731), .ZN(
        n7732) );
  NOR2_X1 U9453 ( .A1(n7733), .A2(n7732), .ZN(n8638) );
  AOI21_X1 U9454 ( .B1(n7733), .B2(n7732), .A(n8638), .ZN(n7760) );
  INV_X1 U9455 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7735) );
  NAND2_X1 U9456 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3151), .ZN(n7734) );
  OAI21_X1 U9457 ( .B1(n8724), .B2(n7735), .A(n7734), .ZN(n7747) );
  INV_X1 U9458 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n7736) );
  MUX2_X1 U9459 ( .A(n7737), .B(n7736), .S(n8748), .Z(n7738) );
  NAND2_X1 U9460 ( .A1(n7738), .A2(n7748), .ZN(n8643) );
  INV_X1 U9461 ( .A(n7738), .ZN(n7739) );
  NAND2_X1 U9462 ( .A1(n7739), .A2(n8652), .ZN(n7740) );
  NAND2_X1 U9463 ( .A1(n8643), .A2(n7740), .ZN(n7741) );
  AOI21_X1 U9464 ( .B1(n7743), .B2(n7742), .A(n7741), .ZN(n8645) );
  INV_X1 U9465 ( .A(n8645), .ZN(n7745) );
  NAND3_X1 U9466 ( .A1(n7743), .A2(n7742), .A3(n7741), .ZN(n7744) );
  AOI21_X1 U9467 ( .B1(n7745), .B2(n7744), .A(n8695), .ZN(n7746) );
  AOI211_X1 U9468 ( .C1(n8699), .C2(n7748), .A(n7747), .B(n7746), .ZN(n7759)
         );
  NOR2_X1 U9469 ( .A1(n7751), .A2(n7750), .ZN(n7753) );
  NAND2_X1 U9470 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n8652), .ZN(n7754) );
  OAI21_X1 U9471 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n8652), .A(n7754), .ZN(
        n7755) );
  NOR2_X1 U9472 ( .A1(n7756), .A2(n7755), .ZN(n8651) );
  AOI21_X1 U9473 ( .B1(n7756), .B2(n7755), .A(n8651), .ZN(n7757) );
  OR2_X1 U9474 ( .A1(n7757), .A2(n8756), .ZN(n7758) );
  OAI211_X1 U9475 ( .C1(n7760), .C2(n8766), .A(n7759), .B(n7758), .ZN(P2_U3196) );
  INV_X1 U9476 ( .A(n7761), .ZN(n7765) );
  AOI22_X1 U9477 ( .A1(n5608), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n6448), .ZN(n7762) );
  OAI21_X1 U9478 ( .B1(n7765), .B2(n7965), .A(n7762), .ZN(P1_U3331) );
  OAI222_X1 U9479 ( .A1(n9058), .A2(n7765), .B1(P2_U3151), .B2(n7764), .C1(
        n7763), .C2(n8186), .ZN(P2_U3271) );
  INV_X1 U9480 ( .A(n7766), .ZN(n9398) );
  XNOR2_X1 U9481 ( .A(n7767), .B(n9398), .ZN(n7771) );
  NAND2_X1 U9482 ( .A1(n9454), .A2(n9169), .ZN(n7769) );
  NAND2_X1 U9483 ( .A1(n9456), .A2(n9291), .ZN(n7768) );
  NAND2_X1 U9484 ( .A1(n7769), .A2(n7768), .ZN(n9196) );
  INV_X1 U9485 ( .A(n9196), .ZN(n7770) );
  OAI21_X1 U9486 ( .B1(n7771), .B2(n9945), .A(n7770), .ZN(n7875) );
  INV_X1 U9487 ( .A(n7875), .ZN(n7780) );
  AOI211_X1 U9488 ( .C1(n7773), .C2(n7772), .A(n9977), .B(n4405), .ZN(n7876)
         );
  NOR2_X1 U9489 ( .A1(n4701), .A2(n9716), .ZN(n7776) );
  OAI22_X1 U9490 ( .A1(n9723), .A2(n7774), .B1(n9194), .B2(n9727), .ZN(n7775)
         );
  AOI211_X1 U9491 ( .C1(n7876), .C2(n9960), .A(n7776), .B(n7775), .ZN(n7779)
         );
  XNOR2_X1 U9492 ( .A(n7777), .B(n9398), .ZN(n7877) );
  NAND2_X1 U9493 ( .A1(n7877), .A2(n9721), .ZN(n7778) );
  OAI211_X1 U9494 ( .C1(n7780), .C2(n4334), .A(n7779), .B(n7778), .ZN(P1_U3278) );
  INV_X1 U9495 ( .A(n7909), .ZN(n7781) );
  NOR2_X1 U9496 ( .A1(n7781), .A2(n8835), .ZN(n7784) );
  INV_X1 U9497 ( .A(n7782), .ZN(n7783) );
  AOI211_X1 U9498 ( .C1(n8908), .C2(n7905), .A(n7784), .B(n7783), .ZN(n7787)
         );
  AOI22_X1 U9499 ( .A1(n7785), .A2(n8906), .B1(P2_REG2_REG_14__SCAN_IN), .B2(
        n8909), .ZN(n7786) );
  OAI21_X1 U9500 ( .B1(n7787), .B2(n8909), .A(n7786), .ZN(P2_U3219) );
  AOI21_X1 U9501 ( .B1(n8345), .B2(n8601), .A(n7788), .ZN(n7791) );
  OR2_X1 U9502 ( .A1(n8258), .A2(n7789), .ZN(n7790) );
  OAI211_X1 U9503 ( .C1(n7792), .C2(n8349), .A(n7791), .B(n7790), .ZN(n7795)
         );
  XNOR2_X1 U9504 ( .A(n7853), .B(n8600), .ZN(n7855) );
  XNOR2_X1 U9505 ( .A(n7855), .B(n7852), .ZN(n7793) );
  NOR2_X1 U9506 ( .A1(n7793), .A2(n8353), .ZN(n7794) );
  AOI211_X1 U9507 ( .C1(n7796), .C2(n8351), .A(n7795), .B(n7794), .ZN(n7797)
         );
  INV_X1 U9508 ( .A(n7797), .ZN(P2_U3157) );
  INV_X1 U9509 ( .A(n7798), .ZN(n7817) );
  INV_X1 U9510 ( .A(n7799), .ZN(n7800) );
  AOI22_X1 U9511 ( .A1(n7800), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n6448), .ZN(n7801) );
  OAI21_X1 U9512 ( .B1(n7817), .B2(n7965), .A(n7801), .ZN(P1_U3330) );
  INV_X1 U9513 ( .A(n7802), .ZN(n10031) );
  OAI21_X1 U9514 ( .B1(n7806), .B2(n7803), .A(n7805), .ZN(n7807) );
  NAND2_X1 U9515 ( .A1(n7807), .A2(n9865), .ZN(n7814) );
  INV_X1 U9516 ( .A(n7808), .ZN(n7811) );
  NOR2_X1 U9517 ( .A1(n9868), .A2(n7809), .ZN(n7810) );
  AOI211_X1 U9518 ( .C1(n9861), .C2(n7812), .A(n7811), .B(n7810), .ZN(n7813)
         );
  OAI211_X1 U9519 ( .C1(n10031), .C2(n9863), .A(n7814), .B(n7813), .ZN(
        P1_U3236) );
  OAI222_X1 U9520 ( .A1(n9058), .A2(n7817), .B1(P2_U3151), .B2(n7816), .C1(
        n7815), .C2(n8186), .ZN(P2_U3270) );
  INV_X1 U9521 ( .A(n7818), .ZN(n7820) );
  XNOR2_X1 U9522 ( .A(n8488), .B(n8200), .ZN(n7903) );
  XNOR2_X1 U9523 ( .A(n7903), .B(n8597), .ZN(n7821) );
  OAI21_X1 U9524 ( .B1(n7822), .B2(n7821), .A(n7904), .ZN(n7823) );
  NAND2_X1 U9525 ( .A1(n7823), .A2(n8321), .ZN(n7828) );
  AOI22_X1 U9526 ( .A1(n8345), .A2(n8598), .B1(P2_REG3_REG_13__SCAN_IN), .B2(
        P2_U3151), .ZN(n7824) );
  OAI21_X1 U9527 ( .B1(n7927), .B2(n8349), .A(n7824), .ZN(n7825) );
  AOI21_X1 U9528 ( .B1(n7826), .B2(n8346), .A(n7825), .ZN(n7827) );
  OAI211_X1 U9529 ( .C1(n7829), .C2(n8329), .A(n7828), .B(n7827), .ZN(P2_U3174) );
  INV_X1 U9530 ( .A(n7830), .ZN(n7874) );
  AOI22_X1 U9531 ( .A1(n7831), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n6448), .ZN(n7832) );
  OAI21_X1 U9532 ( .B1(n7874), .B2(n7965), .A(n7832), .ZN(P1_U3329) );
  XOR2_X1 U9533 ( .A(n7833), .B(n8501), .Z(n7847) );
  INV_X1 U9534 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n8074) );
  AND2_X1 U9535 ( .A1(n8898), .A2(n8596), .ZN(n7838) );
  INV_X1 U9536 ( .A(n7834), .ZN(n7835) );
  AOI211_X1 U9537 ( .C1(n8501), .C2(n7836), .A(n8970), .B(n7835), .ZN(n7837)
         );
  AOI211_X1 U9538 ( .C1(n8899), .C2(n8594), .A(n7838), .B(n7837), .ZN(n7843)
         );
  MUX2_X1 U9539 ( .A(n8074), .B(n7843), .S(n10133), .Z(n7840) );
  NAND2_X1 U9540 ( .A1(n7930), .A2(n9033), .ZN(n7839) );
  OAI211_X1 U9541 ( .C1(n7847), .C2(n9046), .A(n7840), .B(n7839), .ZN(P2_U3435) );
  INV_X1 U9542 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8640) );
  MUX2_X1 U9543 ( .A(n8640), .B(n7843), .S(n10152), .Z(n7842) );
  NAND2_X1 U9544 ( .A1(n7930), .A2(n8948), .ZN(n7841) );
  OAI211_X1 U9545 ( .C1(n8963), .C2(n7847), .A(n7842), .B(n7841), .ZN(P2_U3474) );
  INV_X1 U9546 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n7844) );
  MUX2_X1 U9547 ( .A(n7844), .B(n7843), .S(n8915), .Z(n7846) );
  AOI22_X1 U9548 ( .A1(n7930), .A2(n8888), .B1(n8908), .B2(n7935), .ZN(n7845)
         );
  OAI211_X1 U9549 ( .C1(n7847), .C2(n8891), .A(n7846), .B(n7845), .ZN(P2_U3218) );
  AOI21_X1 U9550 ( .B1(n8345), .B2(n8600), .A(n7848), .ZN(n7851) );
  OR2_X1 U9551 ( .A1(n8258), .A2(n7849), .ZN(n7850) );
  OAI211_X1 U9552 ( .C1(n8482), .C2(n8349), .A(n7851), .B(n7850), .ZN(n7860)
         );
  INV_X1 U9553 ( .A(n7852), .ZN(n7854) );
  OAI22_X1 U9554 ( .A1(n7855), .A2(n7854), .B1(n8600), .B2(n7853), .ZN(n7857)
         );
  XNOR2_X1 U9555 ( .A(n7857), .B(n7856), .ZN(n7858) );
  NOR2_X1 U9556 ( .A1(n7858), .A2(n8353), .ZN(n7859) );
  AOI211_X1 U9557 ( .C1(n10124), .C2(n8351), .A(n7860), .B(n7859), .ZN(n7861)
         );
  INV_X1 U9558 ( .A(n7861), .ZN(P2_U3176) );
  OAI211_X1 U9559 ( .C1(n7863), .C2(n7866), .A(n7862), .B(n8895), .ZN(n7865)
         );
  AOI22_X1 U9560 ( .A1(n8898), .A2(n8595), .B1(n8593), .B2(n8899), .ZN(n7864)
         );
  AND2_X1 U9561 ( .A1(n7865), .A2(n7864), .ZN(n8968) );
  OAI21_X1 U9562 ( .B1(n4409), .B2(n4648), .A(n7867), .ZN(n8967) );
  INV_X1 U9563 ( .A(n8966), .ZN(n7869) );
  AOI22_X1 U9564 ( .A1(n8909), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n8908), .B2(
        n8285), .ZN(n7868) );
  OAI21_X1 U9565 ( .B1(n7869), .B2(n8912), .A(n7868), .ZN(n7870) );
  AOI21_X1 U9566 ( .B1(n8967), .B2(n8906), .A(n7870), .ZN(n7871) );
  OAI21_X1 U9567 ( .B1(n8968), .B2(n8909), .A(n7871), .ZN(P2_U3217) );
  OAI222_X1 U9568 ( .A1(n9058), .A2(n7874), .B1(P2_U3151), .B2(n7873), .C1(
        n7872), .C2(n8186), .ZN(P2_U3269) );
  INV_X1 U9569 ( .A(n9777), .ZN(n9801) );
  INV_X1 U9570 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9489) );
  AOI211_X1 U9571 ( .C1(n7877), .C2(n10029), .A(n7876), .B(n7875), .ZN(n7879)
         );
  MUX2_X1 U9572 ( .A(n9489), .B(n7879), .S(n10068), .Z(n7878) );
  OAI21_X1 U9573 ( .B1(n4701), .B2(n9801), .A(n7878), .ZN(P1_U3537) );
  MUX2_X1 U9574 ( .A(n5268), .B(n7879), .S(n10049), .Z(n7880) );
  OAI21_X1 U9575 ( .B1(n4701), .B2(n9840), .A(n7880), .ZN(P1_U3498) );
  AOI21_X1 U9576 ( .B1(n7881), .B2(n5294), .A(n9945), .ZN(n7884) );
  AOI22_X1 U9577 ( .A1(n9453), .A2(n9169), .B1(n9291), .B2(n9455), .ZN(n9127)
         );
  INV_X1 U9578 ( .A(n9127), .ZN(n7882) );
  AOI21_X1 U9579 ( .B1(n7884), .B2(n7883), .A(n7882), .ZN(n9872) );
  AND2_X1 U9580 ( .A1(n7885), .A2(n9400), .ZN(n9870) );
  INV_X1 U9581 ( .A(n9870), .ZN(n7886) );
  NAND3_X1 U9582 ( .A1(n7886), .A2(n9721), .A3(n9874), .ZN(n7892) );
  INV_X1 U9583 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n7887) );
  OAI22_X1 U9584 ( .A1(n9723), .A2(n7887), .B1(n9126), .B2(n9727), .ZN(n7889)
         );
  OAI211_X1 U9585 ( .C1(n5589), .C2(n4405), .A(n9957), .B(n7945), .ZN(n9871)
         );
  NOR2_X1 U9586 ( .A1(n9871), .A2(n9671), .ZN(n7888) );
  AOI211_X1 U9587 ( .C1(n9953), .C2(n7890), .A(n7889), .B(n7888), .ZN(n7891)
         );
  OAI211_X1 U9588 ( .C1(n4334), .C2(n9872), .A(n7892), .B(n7891), .ZN(P1_U3277) );
  AOI21_X1 U9589 ( .B1(n7893), .B2(n7895), .A(n7894), .ZN(n7896) );
  OAI21_X1 U9590 ( .B1(n4410), .B2(n7896), .A(n9865), .ZN(n7901) );
  NOR2_X1 U9591 ( .A1(n9868), .A2(n9726), .ZN(n7897) );
  AOI211_X1 U9592 ( .C1(n9861), .C2(n7899), .A(n7898), .B(n7897), .ZN(n7900)
         );
  OAI211_X1 U9593 ( .C1(n7902), .C2(n9863), .A(n7901), .B(n7900), .ZN(P1_U3234) );
  XNOR2_X1 U9594 ( .A(n7909), .B(n8254), .ZN(n7926) );
  XNOR2_X1 U9595 ( .A(n7926), .B(n8596), .ZN(n7928) );
  XOR2_X1 U9596 ( .A(n7928), .B(n7929), .Z(n7911) );
  AOI22_X1 U9597 ( .A1(n8314), .A2(n8595), .B1(P2_REG3_REG_14__SCAN_IN), .B2(
        P2_U3151), .ZN(n7907) );
  NAND2_X1 U9598 ( .A1(n8346), .A2(n7905), .ZN(n7906) );
  OAI211_X1 U9599 ( .C1(n4882), .C2(n8317), .A(n7907), .B(n7906), .ZN(n7908)
         );
  AOI21_X1 U9600 ( .B1(n7909), .B2(n8351), .A(n7908), .ZN(n7910) );
  OAI21_X1 U9601 ( .B1(n7911), .B2(n8353), .A(n7910), .ZN(P2_U3155) );
  XNOR2_X1 U9602 ( .A(n7912), .B(n8516), .ZN(n9047) );
  OR2_X1 U9603 ( .A1(n7913), .A2(n8516), .ZN(n7914) );
  NAND3_X1 U9604 ( .A1(n7915), .A2(n7914), .A3(n8895), .ZN(n7917) );
  AOI22_X1 U9605 ( .A1(n8898), .A2(n8594), .B1(n8897), .B2(n8899), .ZN(n7916)
         );
  NAND2_X1 U9606 ( .A1(n7917), .A2(n7916), .ZN(n9043) );
  MUX2_X1 U9607 ( .A(n9043), .B(P2_REG2_REG_17__SCAN_IN), .S(n8909), .Z(n7918)
         );
  INV_X1 U9608 ( .A(n7918), .ZN(n7920) );
  AOI22_X1 U9609 ( .A1(n8289), .A2(n8888), .B1(n8908), .B2(n8300), .ZN(n7919)
         );
  OAI211_X1 U9610 ( .C1(n9047), .C2(n8891), .A(n7920), .B(n7919), .ZN(P2_U3216) );
  INV_X1 U9611 ( .A(n7921), .ZN(n7925) );
  AOI22_X1 U9612 ( .A1(n9896), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n6448), .ZN(n7922) );
  OAI21_X1 U9613 ( .B1(n7925), .B2(n7965), .A(n7922), .ZN(P1_U3328) );
  AOI21_X1 U9614 ( .B1(n9056), .B2(P1_DATAO_REG_27__SCAN_IN), .A(n7923), .ZN(
        n7924) );
  OAI21_X1 U9615 ( .B1(n7925), .B2(n9058), .A(n7924), .ZN(P2_U3268) );
  INV_X1 U9616 ( .A(n7930), .ZN(n7938) );
  XNOR2_X1 U9617 ( .A(n7930), .B(n8200), .ZN(n8202) );
  XNOR2_X1 U9618 ( .A(n8202), .B(n8595), .ZN(n7931) );
  NAND2_X1 U9619 ( .A1(n7932), .A2(n7931), .ZN(n8201) );
  OAI211_X1 U9620 ( .C1(n7932), .C2(n7931), .A(n8201), .B(n8321), .ZN(n7937)
         );
  NAND2_X1 U9621 ( .A1(n8345), .A2(n8596), .ZN(n7933) );
  NAND2_X1 U9622 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8641) );
  OAI211_X1 U9623 ( .C1(n8204), .C2(n8349), .A(n7933), .B(n8641), .ZN(n7934)
         );
  AOI21_X1 U9624 ( .B1(n7935), .B2(n8346), .A(n7934), .ZN(n7936) );
  OAI211_X1 U9625 ( .C1(n7938), .C2(n8329), .A(n7937), .B(n7936), .ZN(P2_U3181) );
  XNOR2_X1 U9626 ( .A(n7939), .B(n9402), .ZN(n9798) );
  INV_X1 U9627 ( .A(n9798), .ZN(n7952) );
  OAI211_X1 U9628 ( .C1(n7941), .C2(n9402), .A(n7940), .B(n9698), .ZN(n7943)
         );
  AND2_X1 U9629 ( .A1(n9454), .A2(n9291), .ZN(n7942) );
  AOI21_X1 U9630 ( .B1(n9452), .B2(n9169), .A(n7942), .ZN(n9138) );
  NAND2_X1 U9631 ( .A1(n7943), .A2(n9138), .ZN(n9796) );
  INV_X1 U9632 ( .A(n9711), .ZN(n7944) );
  AOI211_X1 U9633 ( .C1(n7946), .C2(n7945), .A(n9977), .B(n7944), .ZN(n9797)
         );
  NAND2_X1 U9634 ( .A1(n9797), .A2(n9960), .ZN(n7949) );
  INV_X1 U9635 ( .A(n7947), .ZN(n9140) );
  AOI22_X1 U9636 ( .A1(n4334), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9140), .B2(
        n9951), .ZN(n7948) );
  OAI211_X1 U9637 ( .C1(n4485), .C2(n9716), .A(n7949), .B(n7948), .ZN(n7950)
         );
  AOI21_X1 U9638 ( .B1(n9723), .B2(n9796), .A(n7950), .ZN(n7951) );
  OAI21_X1 U9639 ( .B1(n7952), .B2(n9720), .A(n7951), .ZN(P1_U3276) );
  NAND2_X1 U9640 ( .A1(n7953), .A2(n8397), .ZN(n7954) );
  NAND2_X1 U9641 ( .A1(n7955), .A2(n7954), .ZN(n9042) );
  XNOR2_X1 U9642 ( .A(n7956), .B(n8397), .ZN(n7957) );
  OAI222_X1 U9643 ( .A1(n8860), .A2(n8334), .B1(n8858), .B2(n8283), .C1(n7957), 
        .C2(n8970), .ZN(n8958) );
  NAND2_X1 U9644 ( .A1(n8958), .A2(n8915), .ZN(n7962) );
  INV_X1 U9645 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n7959) );
  INV_X1 U9646 ( .A(n8336), .ZN(n7958) );
  OAI22_X1 U9647 ( .A1(n8915), .A2(n7959), .B1(n7958), .B2(n8770), .ZN(n7960)
         );
  AOI21_X1 U9648 ( .B1(n8959), .B2(n8888), .A(n7960), .ZN(n7961) );
  OAI211_X1 U9649 ( .C1(n9042), .C2(n8891), .A(n7962), .B(n7961), .ZN(P2_U3215) );
  INV_X1 U9650 ( .A(n7963), .ZN(n7968) );
  AOI22_X1 U9651 ( .A1(n9899), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n6448), .ZN(n7964) );
  OAI21_X1 U9652 ( .B1(n7968), .B2(n7965), .A(n7964), .ZN(P1_U3327) );
  AOI21_X1 U9653 ( .B1(n9056), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n7966), .ZN(
        n7967) );
  OAI21_X1 U9654 ( .B1(n7968), .B2(n9058), .A(n7967), .ZN(P2_U3267) );
  NAND2_X1 U9655 ( .A1(n9861), .A2(n7969), .ZN(n7971) );
  OAI211_X1 U9656 ( .C1(n9868), .C2(n7972), .A(n7971), .B(n7970), .ZN(n7978)
         );
  INV_X1 U9657 ( .A(n7893), .ZN(n7976) );
  AOI21_X1 U9658 ( .B1(n7805), .B2(n7974), .A(n7973), .ZN(n7975) );
  NOR3_X1 U9659 ( .A1(n7976), .A2(n7975), .A3(n9188), .ZN(n7977) );
  AOI211_X1 U9660 ( .C1(n7979), .C2(n9186), .A(n7978), .B(n7977), .ZN(n8157)
         );
  AOI22_X1 U9661 ( .A1(n8139), .A2(keyinput122), .B1(n8190), .B2(keyinput117), 
        .ZN(n7980) );
  OAI221_X1 U9662 ( .B1(n8139), .B2(keyinput122), .C1(n8190), .C2(keyinput117), 
        .A(n7980), .ZN(n7989) );
  AOI22_X1 U9663 ( .A1(n7983), .A2(keyinput103), .B1(keyinput73), .B2(n7982), 
        .ZN(n7981) );
  OAI221_X1 U9664 ( .B1(n7983), .B2(keyinput103), .C1(n7982), .C2(keyinput73), 
        .A(n7981), .ZN(n7988) );
  INV_X1 U9665 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n8723) );
  AOI22_X1 U9666 ( .A1(n5120), .A2(keyinput64), .B1(keyinput72), .B2(n8723), 
        .ZN(n7984) );
  OAI221_X1 U9667 ( .B1(n5120), .B2(keyinput64), .C1(n8723), .C2(keyinput72), 
        .A(n7984), .ZN(n7987) );
  AOI22_X1 U9668 ( .A1(n5079), .A2(keyinput90), .B1(keyinput86), .B2(n5057), 
        .ZN(n7985) );
  OAI221_X1 U9669 ( .B1(n5079), .B2(keyinput90), .C1(n5057), .C2(keyinput86), 
        .A(n7985), .ZN(n7986) );
  NOR4_X1 U9670 ( .A1(n7989), .A2(n7988), .A3(n7987), .A4(n7986), .ZN(n8023)
         );
  INV_X1 U9671 ( .A(SI_4_), .ZN(n7991) );
  INV_X1 U9672 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8367) );
  AOI22_X1 U9673 ( .A1(n7991), .A2(keyinput127), .B1(keyinput71), .B2(n8367), 
        .ZN(n7990) );
  OAI221_X1 U9674 ( .B1(n7991), .B2(keyinput127), .C1(n8367), .C2(keyinput71), 
        .A(n7990), .ZN(n8001) );
  INV_X1 U9675 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10134) );
  AOI22_X1 U9676 ( .A1(n7993), .A2(keyinput66), .B1(keyinput84), .B2(n10134), 
        .ZN(n7992) );
  OAI221_X1 U9677 ( .B1(n7993), .B2(keyinput66), .C1(n10134), .C2(keyinput84), 
        .A(n7992), .ZN(n8000) );
  INV_X1 U9678 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n7996) );
  AOI22_X1 U9679 ( .A1(n7996), .A2(keyinput97), .B1(keyinput77), .B2(n7995), 
        .ZN(n7994) );
  OAI221_X1 U9680 ( .B1(n7996), .B2(keyinput97), .C1(n7995), .C2(keyinput77), 
        .A(n7994), .ZN(n7999) );
  AOI22_X1 U9681 ( .A1(n8085), .A2(keyinput105), .B1(keyinput70), .B2(n8074), 
        .ZN(n7997) );
  OAI221_X1 U9682 ( .B1(n8085), .B2(keyinput105), .C1(n8074), .C2(keyinput70), 
        .A(n7997), .ZN(n7998) );
  NOR4_X1 U9683 ( .A1(n8001), .A2(n8000), .A3(n7999), .A4(n7998), .ZN(n8022)
         );
  INV_X1 U9684 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n8920) );
  INV_X1 U9685 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8960) );
  AOI22_X1 U9686 ( .A1(n8920), .A2(keyinput120), .B1(keyinput126), .B2(n8960), 
        .ZN(n8002) );
  OAI221_X1 U9687 ( .B1(n8920), .B2(keyinput120), .C1(n8960), .C2(keyinput126), 
        .A(n8002), .ZN(n8010) );
  AOI22_X1 U9688 ( .A1(n10140), .A2(keyinput69), .B1(n8064), .B2(keyinput76), 
        .ZN(n8003) );
  OAI221_X1 U9689 ( .B1(n10140), .B2(keyinput69), .C1(n8064), .C2(keyinput76), 
        .A(n8003), .ZN(n8009) );
  AOI22_X1 U9690 ( .A1(n6533), .A2(keyinput108), .B1(n8005), .B2(keyinput106), 
        .ZN(n8004) );
  OAI221_X1 U9691 ( .B1(n6533), .B2(keyinput108), .C1(n8005), .C2(keyinput106), 
        .A(n8004), .ZN(n8008) );
  AOI22_X1 U9692 ( .A1(n9170), .A2(keyinput89), .B1(n8142), .B2(keyinput114), 
        .ZN(n8006) );
  OAI221_X1 U9693 ( .B1(n9170), .B2(keyinput89), .C1(n8142), .C2(keyinput114), 
        .A(n8006), .ZN(n8007) );
  NOR4_X1 U9694 ( .A1(n8010), .A2(n8009), .A3(n8008), .A4(n8007), .ZN(n8021)
         );
  INV_X1 U9695 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n8087) );
  INV_X1 U9696 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10120) );
  AOI22_X1 U9697 ( .A1(n8087), .A2(keyinput74), .B1(keyinput68), .B2(n10120), 
        .ZN(n8011) );
  OAI221_X1 U9698 ( .B1(n8087), .B2(keyinput74), .C1(n10120), .C2(keyinput68), 
        .A(n8011), .ZN(n8019) );
  AOI22_X1 U9699 ( .A1(n4960), .A2(keyinput121), .B1(keyinput83), .B2(n8013), 
        .ZN(n8012) );
  OAI221_X1 U9700 ( .B1(n4960), .B2(keyinput121), .C1(n8013), .C2(keyinput83), 
        .A(n8012), .ZN(n8018) );
  AOI22_X1 U9701 ( .A1(n5102), .A2(keyinput93), .B1(keyinput94), .B2(n4641), 
        .ZN(n8014) );
  OAI221_X1 U9702 ( .B1(n5102), .B2(keyinput93), .C1(n4641), .C2(keyinput94), 
        .A(n8014), .ZN(n8017) );
  AOI22_X1 U9703 ( .A1(P2_U3151), .A2(keyinput107), .B1(n8067), .B2(
        keyinput113), .ZN(n8015) );
  OAI221_X1 U9704 ( .B1(P2_U3151), .B2(keyinput107), .C1(n8067), .C2(
        keyinput113), .A(n8015), .ZN(n8016) );
  NOR4_X1 U9705 ( .A1(n8019), .A2(n8018), .A3(n8017), .A4(n8016), .ZN(n8020)
         );
  NAND4_X1 U9706 ( .A1(n8023), .A2(n8022), .A3(n8021), .A4(n8020), .ZN(n8033)
         );
  AOI22_X1 U9707 ( .A1(P2_IR_REG_29__SCAN_IN), .A2(keyinput109), .B1(n8875), 
        .B2(keyinput119), .ZN(n8024) );
  OAI221_X1 U9708 ( .B1(P2_IR_REG_29__SCAN_IN), .B2(keyinput109), .C1(n8875), 
        .C2(keyinput119), .A(n8024), .ZN(n8032) );
  AOI22_X1 U9709 ( .A1(P2_REG0_REG_3__SCAN_IN), .A2(keyinput87), .B1(
        P2_REG2_REG_7__SCAN_IN), .B2(keyinput102), .ZN(n8025) );
  OAI221_X1 U9710 ( .B1(P2_REG0_REG_3__SCAN_IN), .B2(keyinput87), .C1(
        P2_REG2_REG_7__SCAN_IN), .C2(keyinput102), .A(n8025), .ZN(n8030) );
  AOI22_X1 U9711 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(keyinput104), .B1(
        P1_DATAO_REG_4__SCAN_IN), .B2(keyinput67), .ZN(n8026) );
  OAI221_X1 U9712 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(keyinput104), .C1(
        P1_DATAO_REG_4__SCAN_IN), .C2(keyinput67), .A(n8026), .ZN(n8029) );
  XNOR2_X1 U9713 ( .A(n9009), .B(keyinput99), .ZN(n8028) );
  XOR2_X1 U9714 ( .A(SI_2_), .B(keyinput123), .Z(n8027) );
  OR4_X1 U9715 ( .A1(n8030), .A2(n8029), .A3(n8028), .A4(n8027), .ZN(n8031) );
  NOR3_X1 U9716 ( .A1(n8033), .A2(n8032), .A3(n8031), .ZN(n8061) );
  AOI22_X1 U9717 ( .A1(P2_REG1_REG_10__SCAN_IN), .A2(keyinput96), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(keyinput88), .ZN(n8034) );
  OAI221_X1 U9718 ( .B1(P2_REG1_REG_10__SCAN_IN), .B2(keyinput96), .C1(
        P1_DATAO_REG_16__SCAN_IN), .C2(keyinput88), .A(n8034), .ZN(n8041) );
  AOI22_X1 U9719 ( .A1(P2_REG0_REG_1__SCAN_IN), .A2(keyinput78), .B1(
        P2_IR_REG_26__SCAN_IN), .B2(keyinput80), .ZN(n8035) );
  OAI221_X1 U9720 ( .B1(P2_REG0_REG_1__SCAN_IN), .B2(keyinput78), .C1(
        P2_IR_REG_26__SCAN_IN), .C2(keyinput80), .A(n8035), .ZN(n8040) );
  AOI22_X1 U9721 ( .A1(P2_REG2_REG_20__SCAN_IN), .A2(keyinput111), .B1(
        P1_REG3_REG_23__SCAN_IN), .B2(keyinput115), .ZN(n8036) );
  OAI221_X1 U9722 ( .B1(P2_REG2_REG_20__SCAN_IN), .B2(keyinput111), .C1(
        P1_REG3_REG_23__SCAN_IN), .C2(keyinput115), .A(n8036), .ZN(n8039) );
  AOI22_X1 U9723 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(keyinput124), .B1(
        P1_D_REG_0__SCAN_IN), .B2(keyinput118), .ZN(n8037) );
  OAI221_X1 U9724 ( .B1(P1_DATAO_REG_15__SCAN_IN), .B2(keyinput124), .C1(
        P1_D_REG_0__SCAN_IN), .C2(keyinput118), .A(n8037), .ZN(n8038) );
  NOR4_X1 U9725 ( .A1(n8041), .A2(n8040), .A3(n8039), .A4(n8038), .ZN(n8060)
         );
  AOI22_X1 U9726 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(keyinput110), .B1(SI_7_), 
        .B2(keyinput92), .ZN(n8042) );
  OAI221_X1 U9727 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(keyinput110), .C1(SI_7_), 
        .C2(keyinput92), .A(n8042), .ZN(n8049) );
  AOI22_X1 U9728 ( .A1(P2_REG2_REG_29__SCAN_IN), .A2(keyinput101), .B1(
        P1_D_REG_25__SCAN_IN), .B2(keyinput95), .ZN(n8043) );
  OAI221_X1 U9729 ( .B1(P2_REG2_REG_29__SCAN_IN), .B2(keyinput101), .C1(
        P1_D_REG_25__SCAN_IN), .C2(keyinput95), .A(n8043), .ZN(n8048) );
  AOI22_X1 U9730 ( .A1(P1_REG0_REG_11__SCAN_IN), .A2(keyinput125), .B1(
        P1_IR_REG_10__SCAN_IN), .B2(keyinput82), .ZN(n8044) );
  OAI221_X1 U9731 ( .B1(P1_REG0_REG_11__SCAN_IN), .B2(keyinput125), .C1(
        P1_IR_REG_10__SCAN_IN), .C2(keyinput82), .A(n8044), .ZN(n8047) );
  AOI22_X1 U9732 ( .A1(P2_REG1_REG_25__SCAN_IN), .A2(keyinput81), .B1(
        P1_DATAO_REG_22__SCAN_IN), .B2(keyinput79), .ZN(n8045) );
  OAI221_X1 U9733 ( .B1(P2_REG1_REG_25__SCAN_IN), .B2(keyinput81), .C1(
        P1_DATAO_REG_22__SCAN_IN), .C2(keyinput79), .A(n8045), .ZN(n8046) );
  NOR4_X1 U9734 ( .A1(n8049), .A2(n8048), .A3(n8047), .A4(n8046), .ZN(n8059)
         );
  AOI22_X1 U9735 ( .A1(P2_D_REG_17__SCAN_IN), .A2(keyinput116), .B1(
        P1_IR_REG_9__SCAN_IN), .B2(keyinput75), .ZN(n8050) );
  OAI221_X1 U9736 ( .B1(P2_D_REG_17__SCAN_IN), .B2(keyinput116), .C1(
        P1_IR_REG_9__SCAN_IN), .C2(keyinput75), .A(n8050), .ZN(n8057) );
  AOI22_X1 U9737 ( .A1(P2_REG0_REG_26__SCAN_IN), .A2(keyinput98), .B1(
        P2_D_REG_20__SCAN_IN), .B2(keyinput112), .ZN(n8051) );
  OAI221_X1 U9738 ( .B1(P2_REG0_REG_26__SCAN_IN), .B2(keyinput98), .C1(
        P2_D_REG_20__SCAN_IN), .C2(keyinput112), .A(n8051), .ZN(n8056) );
  AOI22_X1 U9739 ( .A1(P2_REG2_REG_19__SCAN_IN), .A2(keyinput100), .B1(
        P1_REG2_REG_17__SCAN_IN), .B2(keyinput85), .ZN(n8052) );
  OAI221_X1 U9740 ( .B1(P2_REG2_REG_19__SCAN_IN), .B2(keyinput100), .C1(
        P1_REG2_REG_17__SCAN_IN), .C2(keyinput85), .A(n8052), .ZN(n8055) );
  AOI22_X1 U9741 ( .A1(SI_28_), .A2(keyinput91), .B1(P2_DATAO_REG_2__SCAN_IN), 
        .B2(keyinput65), .ZN(n8053) );
  OAI221_X1 U9742 ( .B1(SI_28_), .B2(keyinput91), .C1(P2_DATAO_REG_2__SCAN_IN), 
        .C2(keyinput65), .A(n8053), .ZN(n8054) );
  NOR4_X1 U9743 ( .A1(n8057), .A2(n8056), .A3(n8055), .A4(n8054), .ZN(n8058)
         );
  AND4_X1 U9744 ( .A1(n8061), .A2(n8060), .A3(n8059), .A4(n8058), .ZN(n8155)
         );
  AOI22_X1 U9745 ( .A1(n8875), .A2(keyinput55), .B1(keyinput62), .B2(n8960), 
        .ZN(n8062) );
  OAI221_X1 U9746 ( .B1(n8875), .B2(keyinput55), .C1(n8960), .C2(keyinput62), 
        .A(n8062), .ZN(n8071) );
  AOI22_X1 U9747 ( .A1(n7066), .A2(keyinput32), .B1(n8064), .B2(keyinput12), 
        .ZN(n8063) );
  OAI221_X1 U9748 ( .B1(n7066), .B2(keyinput32), .C1(n8064), .C2(keyinput12), 
        .A(n8063), .ZN(n8070) );
  AOI22_X1 U9749 ( .A1(n8367), .A2(keyinput7), .B1(P2_U3151), .B2(keyinput43), 
        .ZN(n8065) );
  OAI221_X1 U9750 ( .B1(n8367), .B2(keyinput7), .C1(P2_U3151), .C2(keyinput43), 
        .A(n8065), .ZN(n8069) );
  AOI22_X1 U9751 ( .A1(n7131), .A2(keyinput38), .B1(n8067), .B2(keyinput49), 
        .ZN(n8066) );
  OAI221_X1 U9752 ( .B1(n7131), .B2(keyinput38), .C1(n8067), .C2(keyinput49), 
        .A(n8066), .ZN(n8068) );
  NOR4_X1 U9753 ( .A1(n8071), .A2(n8070), .A3(n8069), .A4(n8068), .ZN(n8102)
         );
  OAI22_X1 U9754 ( .A1(n10140), .A2(keyinput5), .B1(n6533), .B2(keyinput44), 
        .ZN(n8072) );
  AOI221_X1 U9755 ( .B1(n10140), .B2(keyinput5), .C1(keyinput44), .C2(n6533), 
        .A(n8072), .ZN(n8094) );
  OAI22_X1 U9756 ( .A1(n9504), .A2(keyinput21), .B1(n8074), .B2(keyinput6), 
        .ZN(n8073) );
  AOI221_X1 U9757 ( .B1(n9504), .B2(keyinput21), .C1(keyinput6), .C2(n8074), 
        .A(n8073), .ZN(n8093) );
  AOI22_X1 U9758 ( .A1(n8723), .A2(keyinput8), .B1(n8076), .B2(keyinput15), 
        .ZN(n8075) );
  OAI221_X1 U9759 ( .B1(n8723), .B2(keyinput8), .C1(n8076), .C2(keyinput15), 
        .A(n8075), .ZN(n8082) );
  XNOR2_X1 U9760 ( .A(P1_REG3_REG_7__SCAN_IN), .B(keyinput42), .ZN(n8080) );
  XNOR2_X1 U9761 ( .A(P1_IR_REG_10__SCAN_IN), .B(keyinput18), .ZN(n8079) );
  XNOR2_X1 U9762 ( .A(SI_2_), .B(keyinput59), .ZN(n8078) );
  XNOR2_X1 U9763 ( .A(keyinput26), .B(P1_REG0_REG_7__SCAN_IN), .ZN(n8077) );
  NAND4_X1 U9764 ( .A1(n8080), .A2(n8079), .A3(n8078), .A4(n8077), .ZN(n8081)
         );
  NOR2_X1 U9765 ( .A1(n8082), .A2(n8081), .ZN(n8092) );
  AOI22_X1 U9766 ( .A1(n8085), .A2(keyinput41), .B1(keyinput14), .B2(n8084), 
        .ZN(n8083) );
  OAI221_X1 U9767 ( .B1(n8085), .B2(keyinput41), .C1(n8084), .C2(keyinput14), 
        .A(n8083), .ZN(n8090) );
  INV_X1 U9768 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n8088) );
  AOI22_X1 U9769 ( .A1(n8088), .A2(keyinput46), .B1(n8087), .B2(keyinput10), 
        .ZN(n8086) );
  OAI221_X1 U9770 ( .B1(n8088), .B2(keyinput46), .C1(n8087), .C2(keyinput10), 
        .A(n8086), .ZN(n8089) );
  NOR2_X1 U9771 ( .A1(n8090), .A2(n8089), .ZN(n8091) );
  AND4_X1 U9772 ( .A1(n8094), .A2(n8093), .A3(n8092), .A4(n8091), .ZN(n8101)
         );
  INV_X1 U9773 ( .A(SI_7_), .ZN(n8097) );
  OAI22_X1 U9774 ( .A1(n8097), .A2(keyinput28), .B1(n8096), .B2(keyinput48), 
        .ZN(n8095) );
  AOI221_X1 U9775 ( .B1(n8097), .B2(keyinput28), .C1(keyinput48), .C2(n8096), 
        .A(n8095), .ZN(n8100) );
  OAI22_X1 U9776 ( .A1(n5102), .A2(keyinput29), .B1(n9009), .B2(keyinput35), 
        .ZN(n8098) );
  AOI221_X1 U9777 ( .B1(n5102), .B2(keyinput29), .C1(keyinput35), .C2(n9009), 
        .A(n8098), .ZN(n8099) );
  NAND4_X1 U9778 ( .A1(n8102), .A2(n8101), .A3(n8100), .A4(n8099), .ZN(n8154)
         );
  AOI22_X1 U9779 ( .A1(P2_DATAO_REG_2__SCAN_IN), .A2(keyinput1), .B1(
        P1_D_REG_0__SCAN_IN), .B2(keyinput54), .ZN(n8103) );
  OAI221_X1 U9780 ( .B1(P2_DATAO_REG_2__SCAN_IN), .B2(keyinput1), .C1(
        P1_D_REG_0__SCAN_IN), .C2(keyinput54), .A(n8103), .ZN(n8110) );
  AOI22_X1 U9781 ( .A1(P2_REG3_REG_1__SCAN_IN), .A2(keyinput30), .B1(
        P2_REG1_REG_30__SCAN_IN), .B2(keyinput56), .ZN(n8104) );
  OAI221_X1 U9782 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(keyinput30), .C1(
        P2_REG1_REG_30__SCAN_IN), .C2(keyinput56), .A(n8104), .ZN(n8109) );
  AOI22_X1 U9783 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(keyinput33), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(keyinput53), .ZN(n8105) );
  OAI221_X1 U9784 ( .B1(P1_DATAO_REG_28__SCAN_IN), .B2(keyinput33), .C1(
        P2_DATAO_REG_21__SCAN_IN), .C2(keyinput53), .A(n8105), .ZN(n8108) );
  AOI22_X1 U9785 ( .A1(P2_D_REG_17__SCAN_IN), .A2(keyinput52), .B1(SI_4_), 
        .B2(keyinput63), .ZN(n8106) );
  OAI221_X1 U9786 ( .B1(P2_D_REG_17__SCAN_IN), .B2(keyinput52), .C1(SI_4_), 
        .C2(keyinput63), .A(n8106), .ZN(n8107) );
  NOR4_X1 U9787 ( .A1(n8110), .A2(n8109), .A3(n8108), .A4(n8107), .ZN(n8120)
         );
  AOI22_X1 U9788 ( .A1(P2_D_REG_23__SCAN_IN), .A2(keyinput39), .B1(
        P1_REG0_REG_20__SCAN_IN), .B2(keyinput2), .ZN(n8111) );
  OAI221_X1 U9789 ( .B1(P2_D_REG_23__SCAN_IN), .B2(keyinput39), .C1(
        P1_REG0_REG_20__SCAN_IN), .C2(keyinput2), .A(n8111), .ZN(n8118) );
  AOI22_X1 U9790 ( .A1(P1_REG0_REG_9__SCAN_IN), .A2(keyinput0), .B1(
        P1_REG3_REG_22__SCAN_IN), .B2(keyinput25), .ZN(n8112) );
  OAI221_X1 U9791 ( .B1(P1_REG0_REG_9__SCAN_IN), .B2(keyinput0), .C1(
        P1_REG3_REG_22__SCAN_IN), .C2(keyinput25), .A(n8112), .ZN(n8117) );
  AOI22_X1 U9792 ( .A1(P2_REG0_REG_12__SCAN_IN), .A2(keyinput20), .B1(SI_28_), 
        .B2(keyinput27), .ZN(n8113) );
  OAI221_X1 U9793 ( .B1(P2_REG0_REG_12__SCAN_IN), .B2(keyinput20), .C1(SI_28_), 
        .C2(keyinput27), .A(n8113), .ZN(n8116) );
  AOI22_X1 U9794 ( .A1(P2_D_REG_4__SCAN_IN), .A2(keyinput9), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(keyinput57), .ZN(n8114) );
  OAI221_X1 U9795 ( .B1(P2_D_REG_4__SCAN_IN), .B2(keyinput9), .C1(
        P1_REG3_REG_2__SCAN_IN), .C2(keyinput57), .A(n8114), .ZN(n8115) );
  NOR4_X1 U9796 ( .A1(n8118), .A2(n8117), .A3(n8116), .A4(n8115), .ZN(n8119)
         );
  NAND2_X1 U9797 ( .A1(n8120), .A2(n8119), .ZN(n8153) );
  AOI22_X1 U9798 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(keyinput40), .B1(
        P2_REG2_REG_20__SCAN_IN), .B2(keyinput47), .ZN(n8121) );
  OAI221_X1 U9799 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(keyinput40), .C1(
        P2_REG2_REG_20__SCAN_IN), .C2(keyinput47), .A(n8121), .ZN(n8129) );
  AOI22_X1 U9800 ( .A1(P1_REG0_REG_11__SCAN_IN), .A2(keyinput61), .B1(
        P1_DATAO_REG_4__SCAN_IN), .B2(keyinput3), .ZN(n8122) );
  OAI221_X1 U9801 ( .B1(P1_REG0_REG_11__SCAN_IN), .B2(keyinput61), .C1(
        P1_DATAO_REG_4__SCAN_IN), .C2(keyinput3), .A(n8122), .ZN(n8128) );
  AOI22_X1 U9802 ( .A1(P1_REG2_REG_6__SCAN_IN), .A2(keyinput22), .B1(
        P1_REG3_REG_23__SCAN_IN), .B2(keyinput51), .ZN(n8123) );
  OAI221_X1 U9803 ( .B1(P1_REG2_REG_6__SCAN_IN), .B2(keyinput22), .C1(
        P1_REG3_REG_23__SCAN_IN), .C2(keyinput51), .A(n8123), .ZN(n8127) );
  INV_X1 U9804 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8125) );
  AOI22_X1 U9805 ( .A1(n10120), .A2(keyinput4), .B1(n8125), .B2(keyinput36), 
        .ZN(n8124) );
  OAI221_X1 U9806 ( .B1(n10120), .B2(keyinput4), .C1(n8125), .C2(keyinput36), 
        .A(n8124), .ZN(n8126) );
  NOR4_X1 U9807 ( .A1(n8129), .A2(n8128), .A3(n8127), .A4(n8126), .ZN(n8151)
         );
  AOI22_X1 U9808 ( .A1(P2_REG1_REG_25__SCAN_IN), .A2(keyinput17), .B1(
        P2_IR_REG_29__SCAN_IN), .B2(keyinput45), .ZN(n8130) );
  OAI221_X1 U9809 ( .B1(P2_REG1_REG_25__SCAN_IN), .B2(keyinput17), .C1(
        P2_IR_REG_29__SCAN_IN), .C2(keyinput45), .A(n8130), .ZN(n8137) );
  AOI22_X1 U9810 ( .A1(P2_REG0_REG_3__SCAN_IN), .A2(keyinput23), .B1(
        P2_REG2_REG_29__SCAN_IN), .B2(keyinput37), .ZN(n8131) );
  OAI221_X1 U9811 ( .B1(P2_REG0_REG_3__SCAN_IN), .B2(keyinput23), .C1(
        P2_REG2_REG_29__SCAN_IN), .C2(keyinput37), .A(n8131), .ZN(n8136) );
  AOI22_X1 U9812 ( .A1(P2_REG2_REG_1__SCAN_IN), .A2(keyinput19), .B1(
        P1_IR_REG_9__SCAN_IN), .B2(keyinput11), .ZN(n8132) );
  OAI221_X1 U9813 ( .B1(P2_REG2_REG_1__SCAN_IN), .B2(keyinput19), .C1(
        P1_IR_REG_9__SCAN_IN), .C2(keyinput11), .A(n8132), .ZN(n8135) );
  AOI22_X1 U9814 ( .A1(P2_REG0_REG_26__SCAN_IN), .A2(keyinput34), .B1(
        P2_D_REG_7__SCAN_IN), .B2(keyinput13), .ZN(n8133) );
  OAI221_X1 U9815 ( .B1(P2_REG0_REG_26__SCAN_IN), .B2(keyinput34), .C1(
        P2_D_REG_7__SCAN_IN), .C2(keyinput13), .A(n8133), .ZN(n8134) );
  NOR4_X1 U9816 ( .A1(n8137), .A2(n8136), .A3(n8135), .A4(n8134), .ZN(n8150)
         );
  OAI22_X1 U9817 ( .A1(n8140), .A2(keyinput24), .B1(n8139), .B2(keyinput58), 
        .ZN(n8138) );
  AOI221_X1 U9818 ( .B1(n8140), .B2(keyinput24), .C1(keyinput58), .C2(n8139), 
        .A(n8138), .ZN(n8149) );
  INV_X1 U9819 ( .A(P1_D_REG_25__SCAN_IN), .ZN(n9964) );
  OAI22_X1 U9820 ( .A1(n9964), .A2(keyinput31), .B1(n8142), .B2(keyinput50), 
        .ZN(n8141) );
  AOI221_X1 U9821 ( .B1(n9964), .B2(keyinput31), .C1(keyinput50), .C2(n8142), 
        .A(n8141), .ZN(n8147) );
  OAI22_X1 U9822 ( .A1(n8145), .A2(keyinput60), .B1(n8144), .B2(keyinput16), 
        .ZN(n8143) );
  AOI221_X1 U9823 ( .B1(n8145), .B2(keyinput60), .C1(keyinput16), .C2(n8144), 
        .A(n8143), .ZN(n8146) );
  AND2_X1 U9824 ( .A1(n8147), .A2(n8146), .ZN(n8148) );
  NAND4_X1 U9825 ( .A1(n8151), .A2(n8150), .A3(n8149), .A4(n8148), .ZN(n8152)
         );
  NOR4_X1 U9826 ( .A1(n8155), .A2(n8154), .A3(n8153), .A4(n8152), .ZN(n8156)
         );
  XNOR2_X1 U9827 ( .A(n8157), .B(n8156), .ZN(P1_U3224) );
  OAI222_X1 U9828 ( .A1(n8186), .A2(n8160), .B1(n8159), .B2(n8158), .C1(n8760), 
        .C2(P2_U3151), .ZN(P2_U3276) );
  OAI22_X1 U9829 ( .A1(n8162), .A2(n9727), .B1(n8161), .B2(n9723), .ZN(n8163)
         );
  AOI21_X1 U9830 ( .B1(n8164), .B2(n9953), .A(n8163), .ZN(n8165) );
  OAI21_X1 U9831 ( .B1(n8166), .B2(n9671), .A(n8165), .ZN(n8167) );
  AOI21_X1 U9832 ( .B1(n8168), .B2(n9721), .A(n8167), .ZN(n8169) );
  OAI21_X1 U9833 ( .B1(n8170), .B2(n4334), .A(n8169), .ZN(P1_U3356) );
  INV_X1 U9834 ( .A(SI_29_), .ZN(n8174) );
  INV_X1 U9835 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8176) );
  MUX2_X1 U9836 ( .A(n8176), .B(n8367), .S(n8358), .Z(n8178) );
  INV_X1 U9837 ( .A(SI_30_), .ZN(n8177) );
  NAND2_X1 U9838 ( .A1(n8178), .A2(n8177), .ZN(n8355) );
  INV_X1 U9839 ( .A(n8178), .ZN(n8179) );
  NAND2_X1 U9840 ( .A1(n8179), .A2(SI_30_), .ZN(n8180) );
  NAND2_X1 U9841 ( .A1(n8355), .A2(n8180), .ZN(n8356) );
  INV_X1 U9842 ( .A(n8366), .ZN(n9850) );
  OAI222_X1 U9843 ( .A1(n8186), .A2(n8367), .B1(n9058), .B2(n9850), .C1(
        P2_U3151), .C2(n8181), .ZN(P2_U3265) );
  AOI22_X1 U9844 ( .A1(n6448), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(
        P1_STATE_REG_SCAN_IN), .B2(n8182), .ZN(n8183) );
  OAI21_X1 U9845 ( .B1(n8184), .B2(n7965), .A(n8183), .ZN(P1_U3352) );
  INV_X1 U9846 ( .A(n8185), .ZN(n9853) );
  OAI222_X1 U9847 ( .A1(n9058), .A2(n9853), .B1(n8188), .B2(P2_U3151), .C1(
        n8187), .C2(n8186), .ZN(P2_U3266) );
  OAI222_X1 U9848 ( .A1(n8191), .A2(n8190), .B1(n7965), .B2(n8189), .C1(
        P1_U3086), .C2(n9295), .ZN(P1_U3334) );
  NAND2_X1 U9849 ( .A1(n8366), .A2(n5114), .ZN(n8193) );
  NAND2_X1 U9850 ( .A1(n5465), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n8192) );
  NAND2_X1 U9851 ( .A1(n9741), .A2(n8194), .ZN(n8195) );
  NAND2_X1 U9852 ( .A1(n8195), .A2(n9957), .ZN(n8196) );
  INV_X1 U9853 ( .A(n9425), .ZN(n9202) );
  NOR2_X1 U9854 ( .A1(n8197), .A2(n9202), .ZN(n9735) );
  INV_X1 U9855 ( .A(n9735), .ZN(n9556) );
  NAND2_X1 U9856 ( .A1(n9563), .A2(n9556), .ZN(n9739) );
  MUX2_X1 U9857 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n9739), .S(n10049), .Z(n8198) );
  AOI21_X1 U9858 ( .B1(n9832), .B2(n9741), .A(n8198), .ZN(n8199) );
  INV_X1 U9859 ( .A(n8199), .ZN(P1_U3520) );
  XNOR2_X1 U9860 ( .A(n8289), .B(n8200), .ZN(n8206) );
  XNOR2_X1 U9861 ( .A(n8966), .B(n8254), .ZN(n8205) );
  XOR2_X1 U9862 ( .A(n8594), .B(n8205), .Z(n8281) );
  NAND2_X1 U9863 ( .A1(n8205), .A2(n8204), .ZN(n8290) );
  XNOR2_X1 U9864 ( .A(n8206), .B(n8593), .ZN(n8291) );
  NAND2_X1 U9865 ( .A1(n8207), .A2(n8291), .ZN(n8294) );
  XNOR2_X1 U9866 ( .A(n8959), .B(n8254), .ZN(n8208) );
  XNOR2_X1 U9867 ( .A(n8208), .B(n8897), .ZN(n8332) );
  XNOR2_X1 U9868 ( .A(n8954), .B(n8254), .ZN(n8209) );
  XOR2_X1 U9869 ( .A(n8334), .B(n8209), .Z(n8242) );
  INV_X1 U9870 ( .A(n8209), .ZN(n8210) );
  NAND2_X1 U9871 ( .A1(n8210), .A2(n8883), .ZN(n8211) );
  XNOR2_X1 U9872 ( .A(n9032), .B(n8254), .ZN(n8213) );
  XOR2_X1 U9873 ( .A(n8900), .B(n8213), .Z(n8313) );
  INV_X1 U9874 ( .A(n8313), .ZN(n8212) );
  NAND2_X1 U9875 ( .A1(n8213), .A2(n8268), .ZN(n8214) );
  XNOR2_X1 U9876 ( .A(n9026), .B(n8254), .ZN(n8215) );
  XNOR2_X1 U9877 ( .A(n8215), .B(n8884), .ZN(n8265) );
  XNOR2_X1 U9878 ( .A(n9020), .B(n8254), .ZN(n8216) );
  XOR2_X1 U9879 ( .A(n8843), .B(n8216), .Z(n8323) );
  NAND2_X1 U9880 ( .A1(n8324), .A2(n8323), .ZN(n8322) );
  INV_X1 U9881 ( .A(n8216), .ZN(n8217) );
  NAND2_X1 U9882 ( .A1(n8217), .A2(n8873), .ZN(n8218) );
  XNOR2_X1 U9883 ( .A(n8238), .B(n8254), .ZN(n8220) );
  NAND2_X1 U9884 ( .A1(n8234), .A2(n8859), .ZN(n8223) );
  INV_X1 U9885 ( .A(n8219), .ZN(n8221) );
  NAND2_X1 U9886 ( .A1(n8221), .A2(n8220), .ZN(n8222) );
  XNOR2_X1 U9887 ( .A(n9010), .B(n8254), .ZN(n8224) );
  XNOR2_X1 U9888 ( .A(n8224), .B(n8816), .ZN(n8304) );
  NAND2_X1 U9889 ( .A1(n8224), .A2(n8844), .ZN(n8225) );
  XNOR2_X1 U9890 ( .A(n9004), .B(n8254), .ZN(n8226) );
  XNOR2_X1 U9891 ( .A(n8226), .B(n8832), .ZN(n8273) );
  XNOR2_X1 U9892 ( .A(n8998), .B(n8227), .ZN(n8228) );
  NAND2_X1 U9893 ( .A1(n8228), .A2(n8815), .ZN(n8342) );
  NOR2_X1 U9894 ( .A1(n8228), .A2(n8815), .ZN(n8341) );
  AOI21_X2 U9895 ( .B1(n8340), .B2(n8342), .A(n8341), .ZN(n8251) );
  XNOR2_X1 U9896 ( .A(n8991), .B(n8254), .ZN(n8248) );
  XNOR2_X1 U9897 ( .A(n8248), .B(n8788), .ZN(n8250) );
  XNOR2_X1 U9898 ( .A(n8251), .B(n8250), .ZN(n8233) );
  AOI22_X1 U9899 ( .A1(n8815), .A2(n8345), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n8230) );
  NAND2_X1 U9900 ( .A1(n8799), .A2(n8346), .ZN(n8229) );
  OAI211_X1 U9901 ( .C1(n8551), .C2(n8349), .A(n8230), .B(n8229), .ZN(n8231)
         );
  AOI21_X1 U9902 ( .B1(n8991), .B2(n8351), .A(n8231), .ZN(n8232) );
  OAI21_X1 U9903 ( .B1(n8233), .B2(n8353), .A(n8232), .ZN(P2_U3154) );
  XNOR2_X1 U9904 ( .A(n8234), .B(n8833), .ZN(n8240) );
  AOI22_X1 U9905 ( .A1(n8873), .A2(n8345), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n8236) );
  NAND2_X1 U9906 ( .A1(n8346), .A2(n8847), .ZN(n8235) );
  OAI211_X1 U9907 ( .C1(n8844), .C2(n8349), .A(n8236), .B(n8235), .ZN(n8237)
         );
  AOI21_X1 U9908 ( .B1(n8238), .B2(n8351), .A(n8237), .ZN(n8239) );
  OAI21_X1 U9909 ( .B1(n8240), .B2(n8353), .A(n8239), .ZN(P2_U3156) );
  INV_X1 U9910 ( .A(n8954), .ZN(n8913) );
  OAI211_X1 U9911 ( .C1(n8243), .C2(n8242), .A(n8241), .B(n8321), .ZN(n8247)
         );
  NAND2_X1 U9912 ( .A1(n8345), .A2(n8897), .ZN(n8244) );
  NAND2_X1 U9913 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8758) );
  OAI211_X1 U9914 ( .C1(n8268), .C2(n8349), .A(n8244), .B(n8758), .ZN(n8245)
         );
  AOI21_X1 U9915 ( .B1(n8907), .B2(n8346), .A(n8245), .ZN(n8246) );
  OAI211_X1 U9916 ( .C1(n8913), .C2(n8329), .A(n8247), .B(n8246), .ZN(P2_U3159) );
  INV_X1 U9917 ( .A(n8248), .ZN(n8249) );
  AOI21_X2 U9918 ( .B1(n8251), .B2(n8250), .A(n4901), .ZN(n8256) );
  XNOR2_X1 U9919 ( .A(n8375), .B(n8254), .ZN(n8255) );
  XNOR2_X1 U9920 ( .A(n8256), .B(n8255), .ZN(n8263) );
  INV_X1 U9921 ( .A(n8791), .ZN(n8259) );
  OAI22_X1 U9922 ( .A1(n8259), .A2(n8258), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8257), .ZN(n8261) );
  OAI22_X1 U9923 ( .A1(n8592), .A2(n8349), .B1(n8806), .B2(n8317), .ZN(n8260)
         );
  AOI211_X1 U9924 ( .C1(n8985), .C2(n8351), .A(n8261), .B(n8260), .ZN(n8262)
         );
  OAI21_X1 U9925 ( .B1(n8263), .B2(n8353), .A(n8262), .ZN(P2_U3160) );
  XOR2_X1 U9926 ( .A(n8265), .B(n8264), .Z(n8271) );
  AOI22_X1 U9927 ( .A1(n8873), .A2(n8314), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n8267) );
  NAND2_X1 U9928 ( .A1(n8346), .A2(n8876), .ZN(n8266) );
  OAI211_X1 U9929 ( .C1(n8268), .C2(n8317), .A(n8267), .B(n8266), .ZN(n8269)
         );
  AOI21_X1 U9930 ( .B1(n9026), .B2(n8351), .A(n8269), .ZN(n8270) );
  OAI21_X1 U9931 ( .B1(n8271), .B2(n8353), .A(n8270), .ZN(P2_U3163) );
  XOR2_X1 U9932 ( .A(n8273), .B(n8272), .Z(n8278) );
  AOI22_X1 U9933 ( .A1(n8815), .A2(n8314), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n8275) );
  NAND2_X1 U9934 ( .A1(n8820), .A2(n8346), .ZN(n8274) );
  OAI211_X1 U9935 ( .C1(n8844), .C2(n8317), .A(n8275), .B(n8274), .ZN(n8276)
         );
  AOI21_X1 U9936 ( .B1(n9004), .B2(n8351), .A(n8276), .ZN(n8277) );
  OAI21_X1 U9937 ( .B1(n8278), .B2(n8353), .A(n8277), .ZN(P2_U3165) );
  INV_X1 U9938 ( .A(n8279), .ZN(n8293) );
  AOI21_X1 U9939 ( .B1(n8281), .B2(n8280), .A(n8293), .ZN(n8288) );
  NAND2_X1 U9940 ( .A1(n8345), .A2(n8595), .ZN(n8282) );
  NAND2_X1 U9941 ( .A1(P2_U3151), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8679) );
  OAI211_X1 U9942 ( .C1(n8283), .C2(n8349), .A(n8282), .B(n8679), .ZN(n8284)
         );
  AOI21_X1 U9943 ( .B1(n8285), .B2(n8346), .A(n8284), .ZN(n8287) );
  NAND2_X1 U9944 ( .A1(n8966), .A2(n8351), .ZN(n8286) );
  OAI211_X1 U9945 ( .C1(n8288), .C2(n8353), .A(n8287), .B(n8286), .ZN(P2_U3166) );
  INV_X1 U9946 ( .A(n8289), .ZN(n9045) );
  INV_X1 U9947 ( .A(n8290), .ZN(n8292) );
  NOR3_X1 U9948 ( .A1(n8293), .A2(n8292), .A3(n8291), .ZN(n8296) );
  INV_X1 U9949 ( .A(n8294), .ZN(n8295) );
  OAI21_X1 U9950 ( .B1(n8296), .B2(n8295), .A(n8321), .ZN(n8302) );
  NAND2_X1 U9951 ( .A1(n8345), .A2(n8594), .ZN(n8297) );
  NAND2_X1 U9952 ( .A1(P2_U3151), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8689) );
  OAI211_X1 U9953 ( .C1(n8298), .C2(n8349), .A(n8297), .B(n8689), .ZN(n8299)
         );
  AOI21_X1 U9954 ( .B1(n8300), .B2(n8346), .A(n8299), .ZN(n8301) );
  OAI211_X1 U9955 ( .C1(n9045), .C2(n8329), .A(n8302), .B(n8301), .ZN(P2_U3168) );
  XOR2_X1 U9956 ( .A(n8304), .B(n8303), .Z(n8309) );
  AOI22_X1 U9957 ( .A1(n8832), .A2(n8314), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n8306) );
  NAND2_X1 U9958 ( .A1(n8346), .A2(n8838), .ZN(n8305) );
  OAI211_X1 U9959 ( .C1(n8859), .C2(n8317), .A(n8306), .B(n8305), .ZN(n8307)
         );
  AOI21_X1 U9960 ( .B1(n9010), .B2(n8351), .A(n8307), .ZN(n8308) );
  OAI21_X1 U9961 ( .B1(n8309), .B2(n8353), .A(n8308), .ZN(P2_U3169) );
  INV_X1 U9962 ( .A(n8310), .ZN(n8311) );
  AOI21_X1 U9963 ( .B1(n8313), .B2(n8312), .A(n8311), .ZN(n8320) );
  AOI22_X1 U9964 ( .A1(n8314), .A2(n8884), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n8316) );
  NAND2_X1 U9965 ( .A1(n8346), .A2(n8887), .ZN(n8315) );
  OAI211_X1 U9966 ( .C1(n8334), .C2(n8317), .A(n8316), .B(n8315), .ZN(n8318)
         );
  AOI21_X1 U9967 ( .B1(n9032), .B2(n8351), .A(n8318), .ZN(n8319) );
  OAI21_X1 U9968 ( .B1(n8320), .B2(n8353), .A(n8319), .ZN(P2_U3173) );
  INV_X1 U9969 ( .A(n9020), .ZN(n8330) );
  OAI211_X1 U9970 ( .C1(n8324), .C2(n8323), .A(n8322), .B(n8321), .ZN(n8328)
         );
  AOI22_X1 U9971 ( .A1(n8345), .A2(n8884), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n8325) );
  OAI21_X1 U9972 ( .B1(n8859), .B2(n8349), .A(n8325), .ZN(n8326) );
  AOI21_X1 U9973 ( .B1(n8861), .B2(n8346), .A(n8326), .ZN(n8327) );
  OAI211_X1 U9974 ( .C1(n8330), .C2(n8329), .A(n8328), .B(n8327), .ZN(P2_U3175) );
  XOR2_X1 U9975 ( .A(n8332), .B(n8331), .Z(n8339) );
  NAND2_X1 U9976 ( .A1(n8345), .A2(n8593), .ZN(n8333) );
  NAND2_X1 U9977 ( .A1(P2_U3151), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8721) );
  OAI211_X1 U9978 ( .C1(n8334), .C2(n8349), .A(n8333), .B(n8721), .ZN(n8335)
         );
  AOI21_X1 U9979 ( .B1(n8336), .B2(n8346), .A(n8335), .ZN(n8338) );
  NAND2_X1 U9980 ( .A1(n8959), .A2(n8351), .ZN(n8337) );
  OAI211_X1 U9981 ( .C1(n8339), .C2(n8353), .A(n8338), .B(n8337), .ZN(P2_U3178) );
  INV_X1 U9982 ( .A(n8341), .ZN(n8343) );
  NAND2_X1 U9983 ( .A1(n8343), .A2(n8342), .ZN(n8344) );
  XNOR2_X1 U9984 ( .A(n8340), .B(n8344), .ZN(n8354) );
  AOI22_X1 U9985 ( .A1(n8832), .A2(n8345), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n8348) );
  NAND2_X1 U9986 ( .A1(n8807), .A2(n8346), .ZN(n8347) );
  OAI211_X1 U9987 ( .C1(n8806), .C2(n8349), .A(n8348), .B(n8347), .ZN(n8350)
         );
  AOI21_X1 U9988 ( .B1(n8998), .B2(n8351), .A(n8350), .ZN(n8352) );
  OAI21_X1 U9989 ( .B1(n8354), .B2(n8353), .A(n8352), .ZN(P2_U3180) );
  MUX2_X1 U9990 ( .A(n7412), .B(n6535), .S(n8358), .Z(n8359) );
  XNOR2_X1 U9991 ( .A(n8359), .B(SI_31_), .ZN(n8360) );
  NAND2_X1 U9992 ( .A1(n9199), .A2(n8365), .ZN(n8364) );
  NAND2_X1 U9993 ( .A1(n8362), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n8363) );
  NOR2_X1 U9994 ( .A1(n8575), .A2(n8769), .ZN(n8569) );
  INV_X1 U9995 ( .A(n8569), .ZN(n8373) );
  NAND2_X1 U9996 ( .A1(n8366), .A2(n8365), .ZN(n8370) );
  OR2_X1 U9997 ( .A1(n8368), .A2(n8367), .ZN(n8369) );
  NAND2_X1 U9998 ( .A1(n8571), .A2(n8374), .ZN(n8565) );
  NAND2_X1 U9999 ( .A1(n8565), .A2(n8371), .ZN(n8553) );
  INV_X1 U10000 ( .A(n8553), .ZN(n8372) );
  NAND2_X1 U10001 ( .A1(n8373), .A2(n8372), .ZN(n8581) );
  NAND2_X1 U10002 ( .A1(n8574), .A2(n8570), .ZN(n8554) );
  INV_X1 U10003 ( .A(n8554), .ZN(n8402) );
  INV_X1 U10004 ( .A(n8794), .ZN(n8400) );
  INV_X1 U10005 ( .A(n8376), .ZN(n8544) );
  NAND2_X1 U10006 ( .A1(n8405), .A2(n8404), .ZN(n8831) );
  INV_X1 U10007 ( .A(n8863), .ZN(n8533) );
  INV_X1 U10008 ( .A(n8516), .ZN(n8395) );
  INV_X1 U10009 ( .A(n8377), .ZN(n8486) );
  INV_X1 U10010 ( .A(n8378), .ZN(n8379) );
  NOR2_X1 U10011 ( .A1(n6298), .A2(n8379), .ZN(n8380) );
  AND4_X1 U10012 ( .A1(n8382), .A2(n8381), .A3(n8380), .A4(n8434), .ZN(n8385)
         );
  NAND4_X1 U10013 ( .A1(n8385), .A2(n8384), .A3(n8383), .A4(n8439), .ZN(n8388)
         );
  NOR4_X1 U10014 ( .A1(n8388), .A2(n8387), .A3(n8466), .A4(n8386), .ZN(n8391)
         );
  NAND4_X1 U10015 ( .A1(n8392), .A2(n8391), .A3(n8390), .A4(n8389), .ZN(n8393)
         );
  NOR3_X1 U10016 ( .A1(n8495), .A2(n8486), .A3(n8393), .ZN(n8394) );
  NAND4_X1 U10017 ( .A1(n8395), .A2(n8501), .A3(n4648), .A4(n8394), .ZN(n8396)
         );
  NOR4_X1 U10018 ( .A1(n8881), .A2(n8904), .A3(n8397), .A4(n8396), .ZN(n8398)
         );
  NAND4_X1 U10019 ( .A1(n8846), .A2(n8533), .A3(n8870), .A4(n8398), .ZN(n8399)
         );
  NOR4_X1 U10020 ( .A1(n8400), .A2(n8802), .A3(n8831), .A4(n8399), .ZN(n8401)
         );
  XNOR2_X1 U10021 ( .A(n9004), .B(n8805), .ZN(n8537) );
  INV_X1 U10022 ( .A(n8537), .ZN(n8821) );
  MUX2_X1 U10023 ( .A(n8404), .B(n8403), .S(n8567), .Z(n8539) );
  AND2_X1 U10024 ( .A1(n8405), .A2(n8826), .ZN(n8407) );
  MUX2_X1 U10025 ( .A(n8407), .B(n8406), .S(n8567), .Z(n8536) );
  AND2_X1 U10026 ( .A1(n8532), .A2(n8508), .ZN(n8410) );
  AND2_X1 U10027 ( .A1(n8530), .A2(n8408), .ZN(n8409) );
  MUX2_X1 U10028 ( .A(n8410), .B(n8409), .S(n8567), .Z(n8529) );
  NOR2_X1 U10029 ( .A1(n8881), .A2(n4630), .ZN(n8511) );
  NAND2_X1 U10030 ( .A1(n8521), .A2(n8567), .ZN(n8415) );
  AND2_X1 U10031 ( .A1(n8506), .A2(n8552), .ZN(n8412) );
  NAND2_X1 U10032 ( .A1(n8507), .A2(n8412), .ZN(n8519) );
  INV_X1 U10033 ( .A(n8515), .ZN(n8413) );
  OR2_X1 U10034 ( .A1(n8519), .A2(n8413), .ZN(n8414) );
  OAI21_X1 U10035 ( .B1(n8904), .B2(n8415), .A(n8414), .ZN(n8504) );
  NAND2_X1 U10036 ( .A1(n8441), .A2(n8419), .ZN(n8423) );
  NAND2_X1 U10037 ( .A1(n8608), .A2(n8420), .ZN(n8421) );
  NAND2_X1 U10038 ( .A1(n8456), .A2(n8421), .ZN(n8422) );
  MUX2_X1 U10039 ( .A(n8423), .B(n8422), .S(n8430), .Z(n8424) );
  INV_X1 U10040 ( .A(n8424), .ZN(n8438) );
  INV_X1 U10041 ( .A(n8425), .ZN(n8429) );
  NAND2_X1 U10042 ( .A1(n8433), .A2(n8426), .ZN(n8427) );
  NAND4_X1 U10043 ( .A1(n8429), .A2(n8552), .A3(n8428), .A4(n8427), .ZN(n8436)
         );
  XNOR2_X1 U10044 ( .A(n8431), .B(n8430), .ZN(n8432) );
  OAI21_X1 U10045 ( .B1(n6298), .B2(n8433), .A(n8432), .ZN(n8435) );
  NAND3_X1 U10046 ( .A1(n8436), .A2(n8435), .A3(n8434), .ZN(n8437) );
  NAND2_X1 U10047 ( .A1(n8438), .A2(n8437), .ZN(n8440) );
  NAND2_X1 U10048 ( .A1(n8440), .A2(n8439), .ZN(n8461) );
  INV_X1 U10049 ( .A(n8441), .ZN(n8444) );
  NAND2_X1 U10050 ( .A1(n8606), .A2(n8442), .ZN(n8443) );
  OAI211_X1 U10051 ( .C1(n8461), .C2(n8444), .A(n8462), .B(n8443), .ZN(n8447)
         );
  AND2_X1 U10052 ( .A1(n8445), .A2(n8567), .ZN(n8446) );
  NAND2_X1 U10053 ( .A1(n8447), .A2(n8446), .ZN(n8470) );
  NAND2_X1 U10054 ( .A1(n8470), .A2(n8448), .ZN(n8451) );
  NAND3_X1 U10055 ( .A1(n8451), .A2(n8450), .A3(n8449), .ZN(n8454) );
  NAND2_X1 U10056 ( .A1(n8473), .A2(n8452), .ZN(n8453) );
  AOI21_X1 U10057 ( .B1(n8454), .B2(n8469), .A(n8453), .ZN(n8455) );
  MUX2_X1 U10058 ( .A(n4395), .B(n8455), .S(n8567), .Z(n8472) );
  INV_X1 U10059 ( .A(n8456), .ZN(n8460) );
  INV_X1 U10060 ( .A(n8457), .ZN(n8458) );
  OAI211_X1 U10061 ( .C1(n8461), .C2(n8460), .A(n8459), .B(n8458), .ZN(n8463)
         );
  NAND2_X1 U10062 ( .A1(n8463), .A2(n8462), .ZN(n8468) );
  INV_X1 U10063 ( .A(n8464), .ZN(n8465) );
  NOR2_X1 U10064 ( .A1(n8466), .A2(n8465), .ZN(n8467) );
  NAND4_X1 U10065 ( .A1(n8470), .A2(n8469), .A3(n8468), .A4(n8467), .ZN(n8471)
         );
  NAND2_X1 U10066 ( .A1(n8472), .A2(n8471), .ZN(n8475) );
  NAND3_X1 U10067 ( .A1(n8475), .A2(n8473), .A3(n8478), .ZN(n8474) );
  NAND2_X1 U10068 ( .A1(n8474), .A2(n8476), .ZN(n8481) );
  NAND2_X1 U10069 ( .A1(n8475), .A2(n4904), .ZN(n8479) );
  INV_X1 U10070 ( .A(n8476), .ZN(n8477) );
  AOI21_X1 U10071 ( .B1(n8479), .B2(n8478), .A(n8477), .ZN(n8480) );
  MUX2_X1 U10072 ( .A(n8481), .B(n8480), .S(n8567), .Z(n8487) );
  NAND2_X1 U10073 ( .A1(n10131), .A2(n8482), .ZN(n8483) );
  MUX2_X1 U10074 ( .A(n8484), .B(n8483), .S(n8552), .Z(n8485) );
  OAI21_X1 U10075 ( .B1(n8487), .B2(n8486), .A(n8485), .ZN(n8491) );
  MUX2_X1 U10076 ( .A(n8597), .B(n8488), .S(n8567), .Z(n8493) );
  NAND2_X1 U10077 ( .A1(n8493), .A2(n8489), .ZN(n8490) );
  NAND2_X1 U10078 ( .A1(n8491), .A2(n8490), .ZN(n8494) );
  INV_X1 U10079 ( .A(n8495), .ZN(n8496) );
  MUX2_X1 U10080 ( .A(n8498), .B(n8497), .S(n8552), .Z(n8499) );
  INV_X1 U10081 ( .A(n8499), .ZN(n8500) );
  NAND2_X1 U10082 ( .A1(n8514), .A2(n8502), .ZN(n8503) );
  NAND2_X1 U10083 ( .A1(n8506), .A2(n8505), .ZN(n8510) );
  NAND2_X1 U10084 ( .A1(n8508), .A2(n8507), .ZN(n8509) );
  NAND3_X1 U10085 ( .A1(n8514), .A2(n8513), .A3(n8512), .ZN(n8518) );
  AND2_X1 U10086 ( .A1(n8515), .A2(n8567), .ZN(n8517) );
  AOI21_X1 U10087 ( .B1(n8518), .B2(n8517), .A(n8516), .ZN(n8524) );
  INV_X1 U10088 ( .A(n8519), .ZN(n8523) );
  NAND2_X1 U10089 ( .A1(n8521), .A2(n8520), .ZN(n8522) );
  AOI22_X1 U10090 ( .A1(n8525), .A2(n8524), .B1(n8523), .B2(n8522), .ZN(n8526)
         );
  NAND2_X1 U10091 ( .A1(n8527), .A2(n8526), .ZN(n8528) );
  NAND2_X1 U10092 ( .A1(n8529), .A2(n8528), .ZN(n8534) );
  AOI21_X1 U10093 ( .B1(n8539), .B2(n8538), .A(n8537), .ZN(n8543) );
  MUX2_X1 U10094 ( .A(n4616), .B(n8541), .S(n8567), .Z(n8542) );
  MUX2_X1 U10095 ( .A(n8545), .B(n8544), .S(n8552), .Z(n8546) );
  MUX2_X1 U10096 ( .A(n8548), .B(n8547), .S(n8567), .Z(n8549) );
  MUX2_X1 U10097 ( .A(n8551), .B(n8550), .S(n8552), .Z(n8557) );
  NOR2_X1 U10098 ( .A1(n8561), .A2(n8557), .ZN(n8556) );
  MUX2_X1 U10099 ( .A(n8554), .B(n8553), .S(n8552), .Z(n8555) );
  OR2_X1 U10100 ( .A1(n8558), .A2(n8557), .ZN(n8560) );
  MUX2_X1 U10101 ( .A(n8796), .B(n8985), .S(n8567), .Z(n8559) );
  AOI21_X1 U10102 ( .B1(n8561), .B2(n8560), .A(n8559), .ZN(n8562) );
  INV_X1 U10103 ( .A(n8570), .ZN(n8572) );
  INV_X1 U10104 ( .A(n8571), .ZN(n8775) );
  OAI22_X1 U10105 ( .A1(n8573), .A2(n8572), .B1(n8775), .B2(n8575), .ZN(n8579)
         );
  INV_X1 U10106 ( .A(n8574), .ZN(n8576) );
  NAND2_X1 U10107 ( .A1(n8576), .A2(n8575), .ZN(n8577) );
  OAI211_X1 U10108 ( .C1(n8579), .C2(n8581), .A(n8578), .B(n8577), .ZN(n8580)
         );
  XNOR2_X1 U10109 ( .A(n8583), .B(n8760), .ZN(n8591) );
  NAND3_X1 U10110 ( .A1(n8586), .A2(n8585), .A3(n8584), .ZN(n8587) );
  OAI211_X1 U10111 ( .C1(n8588), .C2(n8590), .A(n8587), .B(P2_B_REG_SCAN_IN), 
        .ZN(n8589) );
  OAI21_X1 U10112 ( .B1(n8591), .B2(n8590), .A(n8589), .ZN(P2_U3296) );
  INV_X1 U10113 ( .A(n8592), .ZN(n8789) );
  MUX2_X1 U10114 ( .A(n8789), .B(P2_DATAO_REG_29__SCAN_IN), .S(n8719), .Z(
        P2_U3520) );
  MUX2_X1 U10115 ( .A(n8796), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8719), .Z(
        P2_U3519) );
  MUX2_X1 U10116 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8788), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U10117 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n8815), .S(P2_U3893), .Z(
        P2_U3517) );
  MUX2_X1 U10118 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8832), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U10119 ( .A(n8816), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8719), .Z(
        P2_U3515) );
  MUX2_X1 U10120 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n8833), .S(P2_U3893), .Z(
        P2_U3514) );
  MUX2_X1 U10121 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8873), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U10122 ( .A(n8884), .B(P2_DATAO_REG_21__SCAN_IN), .S(n8719), .Z(
        P2_U3512) );
  MUX2_X1 U10123 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8883), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U10124 ( .A(n8897), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8719), .Z(
        P2_U3509) );
  MUX2_X1 U10125 ( .A(n8593), .B(P2_DATAO_REG_17__SCAN_IN), .S(n8719), .Z(
        P2_U3508) );
  MUX2_X1 U10126 ( .A(n8594), .B(P2_DATAO_REG_16__SCAN_IN), .S(n8719), .Z(
        P2_U3507) );
  MUX2_X1 U10127 ( .A(n8595), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8719), .Z(
        P2_U3506) );
  MUX2_X1 U10128 ( .A(n8596), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8719), .Z(
        P2_U3505) );
  MUX2_X1 U10129 ( .A(n8597), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8719), .Z(
        P2_U3504) );
  MUX2_X1 U10130 ( .A(n8598), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8719), .Z(
        P2_U3503) );
  MUX2_X1 U10131 ( .A(n8599), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8719), .Z(
        P2_U3502) );
  MUX2_X1 U10132 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n8600), .S(P2_U3893), .Z(
        P2_U3501) );
  MUX2_X1 U10133 ( .A(n8601), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8719), .Z(
        P2_U3500) );
  MUX2_X1 U10134 ( .A(n8602), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8719), .Z(
        P2_U3499) );
  MUX2_X1 U10135 ( .A(n8603), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8719), .Z(
        P2_U3498) );
  MUX2_X1 U10136 ( .A(n8604), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8719), .Z(
        P2_U3497) );
  MUX2_X1 U10137 ( .A(n8605), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8719), .Z(
        P2_U3496) );
  MUX2_X1 U10138 ( .A(n8606), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8719), .Z(
        P2_U3495) );
  MUX2_X1 U10139 ( .A(n8607), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8719), .Z(
        P2_U3494) );
  MUX2_X1 U10140 ( .A(n8608), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8719), .Z(
        P2_U3493) );
  MUX2_X1 U10141 ( .A(n8609), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8719), .Z(
        P2_U3492) );
  MUX2_X1 U10142 ( .A(n8610), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8719), .Z(
        P2_U3491) );
  AND3_X1 U10143 ( .A1(n8613), .A2(n8612), .A3(n8611), .ZN(n8614) );
  OAI21_X1 U10144 ( .B1(n8615), .B2(n8614), .A(n8763), .ZN(n8637) );
  INV_X1 U10145 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n8616) );
  NOR2_X1 U10146 ( .A1(n8724), .A2(n8616), .ZN(n8617) );
  AOI211_X1 U10147 ( .C1(n8699), .C2(n8619), .A(n8618), .B(n8617), .ZN(n8636)
         );
  INV_X1 U10148 ( .A(n8620), .ZN(n8622) );
  NOR3_X1 U10149 ( .A1(n8623), .A2(n8622), .A3(n8621), .ZN(n8624) );
  OAI21_X1 U10150 ( .B1(n8625), .B2(n8624), .A(n8735), .ZN(n8635) );
  INV_X1 U10151 ( .A(n8626), .ZN(n8630) );
  INV_X1 U10152 ( .A(n8627), .ZN(n8629) );
  NOR3_X1 U10153 ( .A1(n8630), .A2(n8629), .A3(n8628), .ZN(n8632) );
  OAI21_X1 U10154 ( .B1(n8633), .B2(n8632), .A(n8631), .ZN(n8634) );
  NAND4_X1 U10155 ( .A1(n8637), .A2(n8636), .A3(n8635), .A4(n8634), .ZN(
        P2_U3190) );
  AOI21_X1 U10156 ( .B1(P2_REG1_REG_14__SCAN_IN), .B2(n8652), .A(n8638), .ZN(
        n8658) );
  AOI21_X1 U10157 ( .B1(n8640), .B2(n8639), .A(n8659), .ZN(n8657) );
  INV_X1 U10158 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n8642) );
  OAI21_X1 U10159 ( .B1(n8724), .B2(n8642), .A(n8641), .ZN(n8650) );
  INV_X1 U10160 ( .A(n8643), .ZN(n8644) );
  NOR2_X1 U10161 ( .A1(n8645), .A2(n8644), .ZN(n8647) );
  MUX2_X1 U10162 ( .A(P2_REG1_REG_15__SCAN_IN), .B(P2_REG2_REG_15__SCAN_IN), 
        .S(n8748), .Z(n8662) );
  XOR2_X1 U10163 ( .A(n8673), .B(n8662), .Z(n8646) );
  NOR2_X1 U10164 ( .A1(n8647), .A2(n8646), .ZN(n8663) );
  AOI21_X1 U10165 ( .B1(n8647), .B2(n8646), .A(n8663), .ZN(n8648) );
  NOR2_X1 U10166 ( .A1(n8648), .A2(n8695), .ZN(n8649) );
  AOI211_X1 U10167 ( .C1(n8699), .C2(n8673), .A(n8650), .B(n8649), .ZN(n8656)
         );
  AOI21_X1 U10168 ( .B1(n7844), .B2(n8653), .A(n8674), .ZN(n8654) );
  OR2_X1 U10169 ( .A1(n8654), .A2(n8756), .ZN(n8655) );
  OAI211_X1 U10170 ( .C1(n8657), .C2(n8766), .A(n8656), .B(n8655), .ZN(
        P2_U3197) );
  NOR2_X1 U10171 ( .A1(n8673), .A2(n8658), .ZN(n8660) );
  INV_X1 U10172 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8666) );
  AOI22_X1 U10173 ( .A1(P2_REG1_REG_16__SCAN_IN), .A2(n8675), .B1(n8701), .B2(
        n8666), .ZN(n8661) );
  AOI21_X1 U10174 ( .B1(n4375), .B2(n8661), .A(n8686), .ZN(n8685) );
  INV_X1 U10175 ( .A(n8662), .ZN(n8664) );
  AOI21_X1 U10176 ( .B1(n8673), .B2(n8664), .A(n8663), .ZN(n8668) );
  INV_X1 U10177 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8665) );
  MUX2_X1 U10178 ( .A(n8666), .B(n8665), .S(n6568), .Z(n8667) );
  NOR2_X1 U10179 ( .A1(n8667), .A2(n8675), .ZN(n8669) );
  NOR2_X1 U10180 ( .A1(n8668), .A2(n8669), .ZN(n8692) );
  INV_X1 U10181 ( .A(n8692), .ZN(n8671) );
  AND2_X1 U10182 ( .A1(n8667), .A2(n8675), .ZN(n8691) );
  OAI21_X1 U10183 ( .B1(n8691), .B2(n8669), .A(n8668), .ZN(n8670) );
  OAI21_X1 U10184 ( .B1(n8671), .B2(n8691), .A(n8670), .ZN(n8683) );
  AOI22_X1 U10185 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n8675), .B1(n8701), .B2(
        n8665), .ZN(n8676) );
  NOR2_X1 U10186 ( .A1(n8677), .A2(n8676), .ZN(n8700) );
  AOI21_X1 U10187 ( .B1(n8677), .B2(n8676), .A(n8700), .ZN(n8678) );
  NOR2_X1 U10188 ( .A1(n8678), .A2(n8756), .ZN(n8682) );
  NAND2_X1 U10189 ( .A1(n8757), .A2(P2_ADDR_REG_16__SCAN_IN), .ZN(n8680) );
  OAI211_X1 U10190 ( .C1(n8761), .C2(n8701), .A(n8680), .B(n8679), .ZN(n8681)
         );
  AOI211_X1 U10191 ( .C1(n8683), .C2(n8763), .A(n8682), .B(n8681), .ZN(n8684)
         );
  OAI21_X1 U10192 ( .B1(n8685), .B2(n8766), .A(n8684), .ZN(P2_U3198) );
  INV_X1 U10193 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8688) );
  AOI21_X1 U10194 ( .B1(P2_REG1_REG_16__SCAN_IN), .B2(n8701), .A(n8686), .ZN(
        n8729) );
  AOI21_X1 U10195 ( .B1(n8688), .B2(n8687), .A(n8727), .ZN(n8708) );
  INV_X1 U10196 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n8690) );
  OAI21_X1 U10197 ( .B1(n8724), .B2(n8690), .A(n8689), .ZN(n8698) );
  NOR2_X1 U10198 ( .A1(n8692), .A2(n8691), .ZN(n8694) );
  MUX2_X1 U10199 ( .A(P2_REG1_REG_17__SCAN_IN), .B(P2_REG2_REG_17__SCAN_IN), 
        .S(n6568), .Z(n8713) );
  XNOR2_X1 U10200 ( .A(n8713), .B(n8702), .ZN(n8693) );
  NOR2_X1 U10201 ( .A1(n8694), .A2(n8693), .ZN(n8714) );
  AOI21_X1 U10202 ( .B1(n8694), .B2(n8693), .A(n8714), .ZN(n8696) );
  NOR2_X1 U10203 ( .A1(n8696), .A2(n8695), .ZN(n8697) );
  AOI211_X1 U10204 ( .C1(n8699), .C2(n8728), .A(n8698), .B(n8697), .ZN(n8707)
         );
  INV_X1 U10205 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8704) );
  AOI21_X1 U10206 ( .B1(n8704), .B2(n8703), .A(n8710), .ZN(n8705) );
  OR2_X1 U10207 ( .A1(n8705), .A2(n8756), .ZN(n8706) );
  OAI211_X1 U10208 ( .C1(n8708), .C2(n8766), .A(n8707), .B(n8706), .ZN(
        P2_U3199) );
  NAND2_X1 U10209 ( .A1(n8730), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n8752) );
  OAI21_X1 U10210 ( .B1(n8730), .B2(P2_REG2_REG_18__SCAN_IN), .A(n8752), .ZN(
        n8711) );
  AOI21_X1 U10211 ( .B1(n8712), .B2(n8711), .A(n8754), .ZN(n8739) );
  INV_X1 U10212 ( .A(n8713), .ZN(n8715) );
  AOI21_X1 U10213 ( .B1(n8728), .B2(n8715), .A(n8714), .ZN(n8717) );
  MUX2_X1 U10214 ( .A(P2_REG1_REG_18__SCAN_IN), .B(P2_REG2_REG_18__SCAN_IN), 
        .S(n6568), .Z(n8716) );
  NOR2_X1 U10215 ( .A1(n8717), .A2(n8716), .ZN(n8745) );
  INV_X1 U10216 ( .A(n8745), .ZN(n8718) );
  NAND2_X1 U10217 ( .A1(n8717), .A2(n8716), .ZN(n8746) );
  NAND2_X1 U10218 ( .A1(n8718), .A2(n8746), .ZN(n8720) );
  OAI21_X1 U10219 ( .B1(n8720), .B2(n8719), .A(n8761), .ZN(n8726) );
  NAND3_X1 U10220 ( .A1(n8720), .A2(n8763), .A3(n8730), .ZN(n8722) );
  OAI211_X1 U10221 ( .C1(n8724), .C2(n8723), .A(n8722), .B(n8721), .ZN(n8725)
         );
  AOI21_X1 U10222 ( .B1(n8747), .B2(n8726), .A(n8725), .ZN(n8738) );
  OR2_X1 U10223 ( .A1(n8729), .A2(n8728), .ZN(n8733) );
  NAND2_X1 U10224 ( .A1(n8730), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8740) );
  NAND2_X1 U10225 ( .A1(n8747), .A2(n8960), .ZN(n8731) );
  NAND2_X1 U10226 ( .A1(n8740), .A2(n8731), .ZN(n8732) );
  AND3_X1 U10227 ( .A1(n8734), .A2(n8733), .A3(n8732), .ZN(n8736) );
  OAI21_X1 U10228 ( .B1(n8742), .B2(n8736), .A(n8735), .ZN(n8737) );
  OAI211_X1 U10229 ( .C1(n8739), .C2(n8756), .A(n8738), .B(n8737), .ZN(
        P2_U3200) );
  INV_X1 U10230 ( .A(n8740), .ZN(n8741) );
  NOR2_X1 U10231 ( .A1(n8742), .A2(n8741), .ZN(n8744) );
  XNOR2_X1 U10232 ( .A(n8760), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8749) );
  INV_X1 U10233 ( .A(n8749), .ZN(n8743) );
  XNOR2_X1 U10234 ( .A(n8744), .B(n8743), .ZN(n8767) );
  AOI21_X1 U10235 ( .B1(n8747), .B2(n8746), .A(n8745), .ZN(n8751) );
  XNOR2_X1 U10236 ( .A(n8760), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n8755) );
  MUX2_X1 U10237 ( .A(n8749), .B(n8755), .S(n6568), .Z(n8750) );
  XNOR2_X1 U10238 ( .A(n8751), .B(n8750), .ZN(n8764) );
  INV_X1 U10239 ( .A(n8752), .ZN(n8753) );
  NAND2_X1 U10240 ( .A1(n8757), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n8759) );
  OAI211_X1 U10241 ( .C1(n8761), .C2(n8760), .A(n8759), .B(n8758), .ZN(n8762)
         );
  OAI21_X1 U10242 ( .B1(n8767), .B2(n8766), .A(n8765), .ZN(P2_U3201) );
  NOR2_X1 U10243 ( .A1(n8769), .A2(n8768), .ZN(n8977) );
  NOR2_X1 U10244 ( .A1(n8771), .A2(n8770), .ZN(n8778) );
  AOI21_X1 U10245 ( .B1(n8977), .B2(n8915), .A(n8778), .ZN(n8774) );
  NAND2_X1 U10246 ( .A1(n8909), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n8772) );
  OAI211_X1 U10247 ( .C1(n8979), .C2(n8912), .A(n8774), .B(n8772), .ZN(
        P2_U3202) );
  NAND2_X1 U10248 ( .A1(n8909), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8773) );
  OAI211_X1 U10249 ( .C1(n8775), .C2(n8912), .A(n8774), .B(n8773), .ZN(
        P2_U3203) );
  NOR2_X1 U10250 ( .A1(n8915), .A2(n8777), .ZN(n8779) );
  AOI211_X1 U10251 ( .C1(n8780), .C2(n8888), .A(n8779), .B(n8778), .ZN(n8784)
         );
  NAND2_X1 U10252 ( .A1(n8782), .A2(n8781), .ZN(n8783) );
  OAI211_X1 U10253 ( .C1(n8776), .C2(n8909), .A(n8784), .B(n8783), .ZN(
        P2_U3204) );
  INV_X1 U10254 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n8790) );
  AOI22_X1 U10255 ( .A1(n8985), .A2(n8888), .B1(n8908), .B2(n8791), .ZN(n8792)
         );
  XNOR2_X1 U10256 ( .A(n8793), .B(n8794), .ZN(n8994) );
  INV_X1 U10257 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n8798) );
  XNOR2_X1 U10258 ( .A(n8795), .B(n8794), .ZN(n8797) );
  AOI222_X1 U10259 ( .A1(n8895), .A2(n8797), .B1(n8796), .B2(n8899), .C1(n8815), .C2(n8898), .ZN(n8989) );
  MUX2_X1 U10260 ( .A(n8798), .B(n8989), .S(n8915), .Z(n8801) );
  AOI22_X1 U10261 ( .A1(n8991), .A2(n8888), .B1(n8908), .B2(n8799), .ZN(n8800)
         );
  OAI211_X1 U10262 ( .C1(n8994), .C2(n8891), .A(n8801), .B(n8800), .ZN(
        P2_U3206) );
  XNOR2_X1 U10263 ( .A(n8803), .B(n8802), .ZN(n8804) );
  OAI222_X1 U10264 ( .A1(n8860), .A2(n8806), .B1(n8858), .B2(n8805), .C1(n8970), .C2(n8804), .ZN(n8995) );
  AOI21_X1 U10265 ( .B1(n8908), .B2(n8807), .A(n8995), .ZN(n8812) );
  AOI22_X1 U10266 ( .A1(n8998), .A2(n8888), .B1(P2_REG2_REG_26__SCAN_IN), .B2(
        n8909), .ZN(n8811) );
  XNOR2_X1 U10267 ( .A(n8809), .B(n8808), .ZN(n8927) );
  NAND2_X1 U10268 ( .A1(n8927), .A2(n8906), .ZN(n8810) );
  OAI211_X1 U10269 ( .C1(n8812), .C2(n8909), .A(n8811), .B(n8810), .ZN(
        P2_U3207) );
  NOR2_X1 U10270 ( .A1(n8813), .A2(n8835), .ZN(n8819) );
  XNOR2_X1 U10271 ( .A(n8814), .B(n8821), .ZN(n8817) );
  AOI222_X1 U10272 ( .A1(n8895), .A2(n8817), .B1(n8816), .B2(n8898), .C1(n8815), .C2(n8899), .ZN(n9002) );
  INV_X1 U10273 ( .A(n9002), .ZN(n8818) );
  AOI211_X1 U10274 ( .C1(n8908), .C2(n8820), .A(n8819), .B(n8818), .ZN(n8825)
         );
  XNOR2_X1 U10275 ( .A(n8822), .B(n8821), .ZN(n9007) );
  INV_X1 U10276 ( .A(n9007), .ZN(n8823) );
  AOI22_X1 U10277 ( .A1(n8823), .A2(n8906), .B1(P2_REG2_REG_25__SCAN_IN), .B2(
        n8909), .ZN(n8824) );
  OAI21_X1 U10278 ( .B1(n8825), .B2(n8909), .A(n8824), .ZN(P2_U3208) );
  INV_X1 U10279 ( .A(n8826), .ZN(n8828) );
  OAI21_X1 U10280 ( .B1(n8845), .B2(n8828), .A(n8827), .ZN(n8829) );
  XNOR2_X1 U10281 ( .A(n8829), .B(n8831), .ZN(n9013) );
  XOR2_X1 U10282 ( .A(n8831), .B(n8830), .Z(n8834) );
  AOI222_X1 U10283 ( .A1(n8895), .A2(n8834), .B1(n8833), .B2(n8898), .C1(n8832), .C2(n8899), .ZN(n9008) );
  OAI21_X1 U10284 ( .B1(n8836), .B2(n8835), .A(n9008), .ZN(n8837) );
  NAND2_X1 U10285 ( .A1(n8837), .A2(n8915), .ZN(n8840) );
  AOI22_X1 U10286 ( .A1(n8838), .A2(n8908), .B1(n8909), .B2(
        P2_REG2_REG_24__SCAN_IN), .ZN(n8839) );
  OAI211_X1 U10287 ( .C1(n9013), .C2(n8891), .A(n8840), .B(n8839), .ZN(
        P2_U3209) );
  XNOR2_X1 U10288 ( .A(n8841), .B(n8846), .ZN(n8842) );
  OAI222_X1 U10289 ( .A1(n8860), .A2(n8844), .B1(n8858), .B2(n8843), .C1(n8970), .C2(n8842), .ZN(n8936) );
  INV_X1 U10290 ( .A(n8936), .ZN(n8851) );
  XOR2_X1 U10291 ( .A(n8846), .B(n8845), .Z(n8937) );
  AOI22_X1 U10292 ( .A1(n8909), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n8847), .B2(
        n8908), .ZN(n8848) );
  OAI21_X1 U10293 ( .B1(n9017), .B2(n8912), .A(n8848), .ZN(n8849) );
  AOI21_X1 U10294 ( .B1(n8937), .B2(n8906), .A(n8849), .ZN(n8850) );
  OAI21_X1 U10295 ( .B1(n8851), .B2(n8909), .A(n8850), .ZN(P2_U3210) );
  INV_X1 U10296 ( .A(n8852), .ZN(n8855) );
  NOR3_X1 U10297 ( .A1(n8868), .A2(n8853), .A3(n8863), .ZN(n8854) );
  NOR2_X1 U10298 ( .A1(n8855), .A2(n8854), .ZN(n8856) );
  OAI222_X1 U10299 ( .A1(n8860), .A2(n8859), .B1(n8858), .B2(n8857), .C1(n8970), .C2(n8856), .ZN(n8940) );
  AOI21_X1 U10300 ( .B1(n8908), .B2(n8861), .A(n8940), .ZN(n8866) );
  AOI22_X1 U10301 ( .A1(n9020), .A2(n8888), .B1(P2_REG2_REG_22__SCAN_IN), .B2(
        n8909), .ZN(n8865) );
  XNOR2_X1 U10302 ( .A(n8862), .B(n8863), .ZN(n9021) );
  NAND2_X1 U10303 ( .A1(n9021), .A2(n8906), .ZN(n8864) );
  OAI211_X1 U10304 ( .C1(n8866), .C2(n8909), .A(n8865), .B(n8864), .ZN(
        P2_U3211) );
  XOR2_X1 U10305 ( .A(n8870), .B(n8867), .Z(n9029) );
  INV_X1 U10306 ( .A(n8868), .ZN(n8872) );
  NAND3_X1 U10307 ( .A1(n8880), .A2(n8870), .A3(n8869), .ZN(n8871) );
  NAND2_X1 U10308 ( .A1(n8872), .A2(n8871), .ZN(n8874) );
  AOI222_X1 U10309 ( .A1(n8895), .A2(n8874), .B1(n8900), .B2(n8898), .C1(n8873), .C2(n8899), .ZN(n9024) );
  MUX2_X1 U10310 ( .A(n8875), .B(n9024), .S(n8915), .Z(n8878) );
  AOI22_X1 U10311 ( .A1(n9026), .A2(n8888), .B1(n8908), .B2(n8876), .ZN(n8877)
         );
  OAI211_X1 U10312 ( .C1(n9029), .C2(n8891), .A(n8878), .B(n8877), .ZN(
        P2_U3212) );
  XNOR2_X1 U10313 ( .A(n8879), .B(n8881), .ZN(n9035) );
  INV_X1 U10314 ( .A(n9035), .ZN(n8892) );
  OAI21_X1 U10315 ( .B1(n8882), .B2(n8881), .A(n8880), .ZN(n8885) );
  AOI222_X1 U10316 ( .A1(n8895), .A2(n8885), .B1(n8884), .B2(n8899), .C1(n8883), .C2(n8898), .ZN(n9030) );
  MUX2_X1 U10317 ( .A(n8886), .B(n9030), .S(n8915), .Z(n8890) );
  AOI22_X1 U10318 ( .A1(n9032), .A2(n8888), .B1(n8908), .B2(n8887), .ZN(n8889)
         );
  OAI211_X1 U10319 ( .C1(n8892), .C2(n8891), .A(n8890), .B(n8889), .ZN(
        P2_U3213) );
  XNOR2_X1 U10320 ( .A(n8894), .B(n8893), .ZN(n8896) );
  NAND2_X1 U10321 ( .A1(n8896), .A2(n8895), .ZN(n8902) );
  AOI22_X1 U10322 ( .A1(n8900), .A2(n8899), .B1(n8898), .B2(n8897), .ZN(n8901)
         );
  NAND2_X1 U10323 ( .A1(n8902), .A2(n8901), .ZN(n8955) );
  INV_X1 U10324 ( .A(n8903), .ZN(n8905) );
  NAND2_X1 U10325 ( .A1(n8905), .A2(n8904), .ZN(n8953) );
  NAND3_X1 U10326 ( .A1(n8953), .A2(n8906), .A3(n8952), .ZN(n8911) );
  AOI22_X1 U10327 ( .A1(n8909), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n8908), .B2(
        n8907), .ZN(n8910) );
  OAI211_X1 U10328 ( .C1(n8913), .C2(n8912), .A(n8911), .B(n8910), .ZN(n8914)
         );
  AOI21_X1 U10329 ( .B1(n8955), .B2(n8915), .A(n8914), .ZN(n8916) );
  INV_X1 U10330 ( .A(n8916), .ZN(P2_U3214) );
  INV_X1 U10331 ( .A(n8948), .ZN(n8962) );
  NAND2_X1 U10332 ( .A1(n8977), .A2(n10152), .ZN(n8918) );
  NAND2_X1 U10333 ( .A1(n10150), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n8917) );
  OAI211_X1 U10334 ( .C1(n8979), .C2(n8962), .A(n8918), .B(n8917), .ZN(
        P2_U3490) );
  NAND2_X1 U10335 ( .A1(n8571), .A2(n8948), .ZN(n8919) );
  OAI211_X1 U10336 ( .C1(n10152), .C2(n8920), .A(n8919), .B(n8918), .ZN(
        P2_U3489) );
  MUX2_X1 U10337 ( .A(n8921), .B(n8983), .S(n10152), .Z(n8923) );
  NAND2_X1 U10338 ( .A1(n8985), .A2(n8948), .ZN(n8922) );
  OAI211_X1 U10339 ( .C1(n8988), .C2(n8963), .A(n8923), .B(n8922), .ZN(
        P2_U3487) );
  MUX2_X1 U10340 ( .A(n8924), .B(n8989), .S(n10152), .Z(n8926) );
  NAND2_X1 U10341 ( .A1(n8991), .A2(n8948), .ZN(n8925) );
  OAI211_X1 U10342 ( .C1(n8994), .C2(n8963), .A(n8926), .B(n8925), .ZN(
        P2_U3486) );
  MUX2_X1 U10343 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n8995), .S(n10152), .Z(
        n8929) );
  INV_X1 U10344 ( .A(n8927), .ZN(n9001) );
  OAI22_X1 U10345 ( .A1(n9001), .A2(n8963), .B1(n4658), .B2(n8962), .ZN(n8928)
         );
  OR2_X1 U10346 ( .A1(n8929), .A2(n8928), .ZN(P2_U3485) );
  MUX2_X1 U10347 ( .A(n8930), .B(n9002), .S(n10152), .Z(n8932) );
  NAND2_X1 U10348 ( .A1(n9004), .A2(n8948), .ZN(n8931) );
  OAI211_X1 U10349 ( .C1(n8963), .C2(n9007), .A(n8932), .B(n8931), .ZN(
        P2_U3484) );
  INV_X1 U10350 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n8933) );
  MUX2_X1 U10351 ( .A(n8933), .B(n9008), .S(n10152), .Z(n8935) );
  NAND2_X1 U10352 ( .A1(n9010), .A2(n8948), .ZN(n8934) );
  OAI211_X1 U10353 ( .C1(n8963), .C2(n9013), .A(n8935), .B(n8934), .ZN(
        P2_U3483) );
  AOI21_X1 U10354 ( .B1(n10091), .B2(n8937), .A(n8936), .ZN(n9014) );
  MUX2_X1 U10355 ( .A(n8938), .B(n9014), .S(n10152), .Z(n8939) );
  OAI21_X1 U10356 ( .B1(n9017), .B2(n8962), .A(n8939), .ZN(P2_U3482) );
  INV_X1 U10357 ( .A(n8940), .ZN(n9018) );
  MUX2_X1 U10358 ( .A(n8941), .B(n9018), .S(n10152), .Z(n8943) );
  AOI22_X1 U10359 ( .A1(n9021), .A2(n8949), .B1(n8948), .B2(n9020), .ZN(n8942)
         );
  NAND2_X1 U10360 ( .A1(n8943), .A2(n8942), .ZN(P2_U3481) );
  INV_X1 U10361 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8944) );
  MUX2_X1 U10362 ( .A(n8944), .B(n9024), .S(n10152), .Z(n8946) );
  NAND2_X1 U10363 ( .A1(n9026), .A2(n8948), .ZN(n8945) );
  OAI211_X1 U10364 ( .C1(n8963), .C2(n9029), .A(n8946), .B(n8945), .ZN(
        P2_U3480) );
  INV_X1 U10365 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n8947) );
  MUX2_X1 U10366 ( .A(n8947), .B(n9030), .S(n10152), .Z(n8951) );
  AOI22_X1 U10367 ( .A1(n9035), .A2(n8949), .B1(n8948), .B2(n9032), .ZN(n8950)
         );
  NAND2_X1 U10368 ( .A1(n8951), .A2(n8950), .ZN(P2_U3479) );
  AND3_X1 U10369 ( .A1(n8953), .A2(n8952), .A3(n10091), .ZN(n8957) );
  AND2_X1 U10370 ( .A1(n8954), .A2(n10132), .ZN(n8956) );
  MUX2_X1 U10371 ( .A(n9038), .B(P2_REG1_REG_19__SCAN_IN), .S(n10150), .Z(
        P2_U3478) );
  AOI21_X1 U10372 ( .B1(n10132), .B2(n8959), .A(n8958), .ZN(n9039) );
  MUX2_X1 U10373 ( .A(n8960), .B(n9039), .S(n10152), .Z(n8961) );
  OAI21_X1 U10374 ( .B1(n8963), .B2(n9042), .A(n8961), .ZN(P2_U3477) );
  MUX2_X1 U10375 ( .A(n9043), .B(P2_REG1_REG_17__SCAN_IN), .S(n10150), .Z(
        n8965) );
  OAI22_X1 U10376 ( .A1(n9047), .A2(n8963), .B1(n9045), .B2(n8962), .ZN(n8964)
         );
  OR2_X1 U10377 ( .A1(n8965), .A2(n8964), .ZN(P2_U3476) );
  AOI22_X1 U10378 ( .A1(n8967), .A2(n10091), .B1(n10132), .B2(n8966), .ZN(
        n8969) );
  NAND2_X1 U10379 ( .A1(n8969), .A2(n8968), .ZN(n9050) );
  MUX2_X1 U10380 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n9050), .S(n10152), .Z(
        P2_U3475) );
  NAND2_X1 U10381 ( .A1(n10126), .A2(n8970), .ZN(n8974) );
  OAI21_X1 U10382 ( .B1(n10114), .B2(n8972), .A(n8971), .ZN(n8973) );
  AOI21_X1 U10383 ( .B1(n8975), .B2(n8974), .A(n8973), .ZN(n10069) );
  INV_X1 U10384 ( .A(n10069), .ZN(n8976) );
  MUX2_X1 U10385 ( .A(P2_REG1_REG_0__SCAN_IN), .B(n8976), .S(n10152), .Z(
        P2_U3459) );
  NAND2_X1 U10386 ( .A1(n8977), .A2(n10133), .ZN(n8980) );
  NAND2_X1 U10387 ( .A1(n10135), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n8978) );
  OAI211_X1 U10388 ( .C1(n8979), .C2(n9044), .A(n8980), .B(n8978), .ZN(
        P2_U3458) );
  INV_X1 U10389 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n8982) );
  NAND2_X1 U10390 ( .A1(n8571), .A2(n9033), .ZN(n8981) );
  OAI211_X1 U10391 ( .C1(n8982), .C2(n10133), .A(n8981), .B(n8980), .ZN(
        P2_U3457) );
  INV_X1 U10392 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n8984) );
  MUX2_X1 U10393 ( .A(n8984), .B(n8983), .S(n10133), .Z(n8987) );
  NAND2_X1 U10394 ( .A1(n8985), .A2(n9033), .ZN(n8986) );
  OAI211_X1 U10395 ( .C1(n8988), .C2(n9046), .A(n8987), .B(n8986), .ZN(
        P2_U3455) );
  INV_X1 U10396 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n8990) );
  MUX2_X1 U10397 ( .A(n8990), .B(n8989), .S(n10133), .Z(n8993) );
  NAND2_X1 U10398 ( .A1(n8991), .A2(n9033), .ZN(n8992) );
  OAI211_X1 U10399 ( .C1(n8994), .C2(n9046), .A(n8993), .B(n8992), .ZN(
        P2_U3454) );
  INV_X1 U10400 ( .A(n8995), .ZN(n8996) );
  MUX2_X1 U10401 ( .A(n8997), .B(n8996), .S(n10133), .Z(n9000) );
  NAND2_X1 U10402 ( .A1(n8998), .A2(n9033), .ZN(n8999) );
  OAI211_X1 U10403 ( .C1(n9001), .C2(n9046), .A(n9000), .B(n8999), .ZN(
        P2_U3453) );
  INV_X1 U10404 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n9003) );
  MUX2_X1 U10405 ( .A(n9003), .B(n9002), .S(n10133), .Z(n9006) );
  NAND2_X1 U10406 ( .A1(n9004), .A2(n9033), .ZN(n9005) );
  OAI211_X1 U10407 ( .C1(n9007), .C2(n9046), .A(n9006), .B(n9005), .ZN(
        P2_U3452) );
  MUX2_X1 U10408 ( .A(n9009), .B(n9008), .S(n10133), .Z(n9012) );
  NAND2_X1 U10409 ( .A1(n9010), .A2(n9033), .ZN(n9011) );
  OAI211_X1 U10410 ( .C1(n9013), .C2(n9046), .A(n9012), .B(n9011), .ZN(
        P2_U3451) );
  INV_X1 U10411 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n9015) );
  MUX2_X1 U10412 ( .A(n9015), .B(n9014), .S(n10133), .Z(n9016) );
  OAI21_X1 U10413 ( .B1(n9017), .B2(n9044), .A(n9016), .ZN(P2_U3450) );
  INV_X1 U10414 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n9019) );
  MUX2_X1 U10415 ( .A(n9019), .B(n9018), .S(n10133), .Z(n9023) );
  AOI22_X1 U10416 ( .A1(n9021), .A2(n9034), .B1(n9033), .B2(n9020), .ZN(n9022)
         );
  NAND2_X1 U10417 ( .A1(n9023), .A2(n9022), .ZN(P2_U3449) );
  INV_X1 U10418 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n9025) );
  MUX2_X1 U10419 ( .A(n9025), .B(n9024), .S(n10133), .Z(n9028) );
  NAND2_X1 U10420 ( .A1(n9026), .A2(n9033), .ZN(n9027) );
  OAI211_X1 U10421 ( .C1(n9029), .C2(n9046), .A(n9028), .B(n9027), .ZN(
        P2_U3448) );
  INV_X1 U10422 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n9031) );
  MUX2_X1 U10423 ( .A(n9031), .B(n9030), .S(n10133), .Z(n9037) );
  AOI22_X1 U10424 ( .A1(n9035), .A2(n9034), .B1(n9033), .B2(n9032), .ZN(n9036)
         );
  NAND2_X1 U10425 ( .A1(n9037), .A2(n9036), .ZN(P2_U3447) );
  MUX2_X1 U10426 ( .A(n9038), .B(P2_REG0_REG_19__SCAN_IN), .S(n10135), .Z(
        P2_U3446) );
  INV_X1 U10427 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n9040) );
  MUX2_X1 U10428 ( .A(n9040), .B(n9039), .S(n10133), .Z(n9041) );
  OAI21_X1 U10429 ( .B1(n9042), .B2(n9046), .A(n9041), .ZN(P2_U3444) );
  MUX2_X1 U10430 ( .A(n9043), .B(P2_REG0_REG_17__SCAN_IN), .S(n10135), .Z(
        n9049) );
  OAI22_X1 U10431 ( .A1(n9047), .A2(n9046), .B1(n9045), .B2(n9044), .ZN(n9048)
         );
  OR2_X1 U10432 ( .A1(n9049), .A2(n9048), .ZN(P2_U3441) );
  MUX2_X1 U10433 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n9050), .S(n10133), .Z(
        P2_U3438) );
  MUX2_X1 U10434 ( .A(n9052), .B(P2_D_REG_1__SCAN_IN), .S(n9051), .Z(P2_U3377)
         );
  INV_X1 U10435 ( .A(n9199), .ZN(n9847) );
  NOR4_X1 U10436 ( .A1(n9054), .A2(P2_IR_REG_30__SCAN_IN), .A3(P2_U3151), .A4(
        n6138), .ZN(n9055) );
  AOI21_X1 U10437 ( .B1(n9056), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n9055), .ZN(
        n9057) );
  OAI21_X1 U10438 ( .B1(n9847), .B2(n9058), .A(n9057), .ZN(P2_U3264) );
  INV_X1 U10439 ( .A(n9059), .ZN(n9060) );
  MUX2_X1 U10440 ( .A(n9060), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  AOI21_X1 U10441 ( .B1(n9063), .B2(n9062), .A(n9061), .ZN(n9064) );
  OAI21_X1 U10442 ( .B1(n9065), .B2(n9064), .A(n9865), .ZN(n9069) );
  AOI22_X1 U10443 ( .A1(n9443), .A2(n9169), .B1(n9291), .B2(n9445), .ZN(n9578)
         );
  AOI22_X1 U10444 ( .A1(n9584), .A2(n9162), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3086), .ZN(n9066) );
  OAI21_X1 U10445 ( .B1(n9578), .B2(n9183), .A(n9066), .ZN(n9067) );
  AOI21_X1 U10446 ( .B1(n9583), .B2(n9186), .A(n9067), .ZN(n9068) );
  NAND2_X1 U10447 ( .A1(n9069), .A2(n9068), .ZN(P1_U3214) );
  NOR2_X1 U10448 ( .A1(n4414), .A2(n4347), .ZN(n9071) );
  XNOR2_X1 U10449 ( .A(n9071), .B(n9070), .ZN(n9078) );
  AOI22_X1 U10450 ( .A1(n9861), .A2(n9072), .B1(P1_REG3_REG_14__SCAN_IN), .B2(
        P1_U3086), .ZN(n9073) );
  OAI21_X1 U10451 ( .B1(n9074), .B2(n9868), .A(n9073), .ZN(n9075) );
  AOI21_X1 U10452 ( .B1(n9076), .B2(n9186), .A(n9075), .ZN(n9077) );
  OAI21_X1 U10453 ( .B1(n9078), .B2(n9188), .A(n9077), .ZN(P1_U3215) );
  INV_X1 U10454 ( .A(n9079), .ZN(n9081) );
  NOR2_X1 U10455 ( .A1(n9081), .A2(n9080), .ZN(n9084) );
  INV_X1 U10456 ( .A(n9083), .ZN(n9146) );
  AOI21_X1 U10457 ( .B1(n9084), .B2(n9082), .A(n9146), .ZN(n9090) );
  OAI22_X1 U10458 ( .A1(n9086), .A2(n9096), .B1(n9085), .B2(n9106), .ZN(n9635)
         );
  AOI22_X1 U10459 ( .A1(n9635), .A2(n9861), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3086), .ZN(n9087) );
  OAI21_X1 U10460 ( .B1(n9639), .B2(n9868), .A(n9087), .ZN(n9088) );
  AOI21_X1 U10461 ( .B1(n9824), .B2(n9186), .A(n9088), .ZN(n9089) );
  OAI21_X1 U10462 ( .B1(n9090), .B2(n9188), .A(n9089), .ZN(P1_U3216) );
  INV_X1 U10463 ( .A(n9091), .ZN(n9092) );
  NOR2_X1 U10464 ( .A1(n9093), .A2(n9092), .ZN(n9094) );
  XNOR2_X1 U10465 ( .A(n9095), .B(n9094), .ZN(n9102) );
  OR2_X1 U10466 ( .A1(n9107), .A2(n9096), .ZN(n9098) );
  NAND2_X1 U10467 ( .A1(n9452), .A2(n9291), .ZN(n9097) );
  NAND2_X1 U10468 ( .A1(n9098), .A2(n9097), .ZN(n9697) );
  AOI22_X1 U10469 ( .A1(n9697), .A2(n9861), .B1(P1_REG3_REG_19__SCAN_IN), .B2(
        P1_U3086), .ZN(n9099) );
  OAI21_X1 U10470 ( .B1(n9691), .B2(n9868), .A(n9099), .ZN(n9100) );
  AOI21_X1 U10471 ( .B1(n9787), .B2(n9186), .A(n9100), .ZN(n9101) );
  OAI21_X1 U10472 ( .B1(n9102), .B2(n9188), .A(n9101), .ZN(P1_U3219) );
  OAI21_X1 U10473 ( .B1(n9105), .B2(n9104), .A(n9103), .ZN(n9113) );
  NAND2_X1 U10474 ( .A1(n9831), .A2(n9186), .ZN(n9111) );
  NAND2_X1 U10475 ( .A1(n9449), .A2(n9181), .ZN(n9109) );
  OR2_X1 U10476 ( .A1(n9107), .A2(n9106), .ZN(n9108) );
  NAND2_X1 U10477 ( .A1(n9109), .A2(n9108), .ZN(n9660) );
  AOI22_X1 U10478 ( .A1(n9660), .A2(n9861), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3086), .ZN(n9110) );
  OAI211_X1 U10479 ( .C1(n9868), .C2(n9668), .A(n9111), .B(n9110), .ZN(n9112)
         );
  AOI21_X1 U10480 ( .B1(n9113), .B2(n9865), .A(n9112), .ZN(n9114) );
  INV_X1 U10481 ( .A(n9114), .ZN(P1_U3223) );
  NAND2_X1 U10482 ( .A1(n9445), .A2(n9181), .ZN(n9117) );
  NAND2_X1 U10483 ( .A1(n9447), .A2(n9291), .ZN(n9116) );
  NAND2_X1 U10484 ( .A1(n9117), .A2(n9116), .ZN(n9607) );
  INV_X1 U10485 ( .A(n9612), .ZN(n9119) );
  OAI22_X1 U10486 ( .A1(n9119), .A2(n9868), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9118), .ZN(n9120) );
  AOI21_X1 U10487 ( .B1(n9607), .B2(n9861), .A(n9120), .ZN(n9121) );
  OAI211_X1 U10488 ( .C1(n9817), .C2(n9863), .A(n9122), .B(n9121), .ZN(
        P1_U3225) );
  NAND2_X1 U10489 ( .A1(n9123), .A2(n9124), .ZN(n9133) );
  OAI21_X1 U10490 ( .B1(n9124), .B2(n9123), .A(n9133), .ZN(n9125) );
  NAND2_X1 U10491 ( .A1(n9125), .A2(n9865), .ZN(n9131) );
  INV_X1 U10492 ( .A(n9126), .ZN(n9129) );
  NAND2_X1 U10493 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9925) );
  OAI21_X1 U10494 ( .B1(n9183), .B2(n9127), .A(n9925), .ZN(n9128) );
  AOI21_X1 U10495 ( .B1(n9129), .B2(n9162), .A(n9128), .ZN(n9130) );
  OAI211_X1 U10496 ( .C1(n5589), .C2(n9863), .A(n9131), .B(n9130), .ZN(
        P1_U3226) );
  NAND2_X1 U10497 ( .A1(n9133), .A2(n9132), .ZN(n9135) );
  OAI21_X1 U10498 ( .B1(n9136), .B2(n9135), .A(n9134), .ZN(n9137) );
  NAND2_X1 U10499 ( .A1(n9137), .A2(n9865), .ZN(n9142) );
  NAND2_X1 U10500 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9513) );
  OAI21_X1 U10501 ( .B1(n9183), .B2(n9138), .A(n9513), .ZN(n9139) );
  AOI21_X1 U10502 ( .B1(n9140), .B2(n9162), .A(n9139), .ZN(n9141) );
  OAI211_X1 U10503 ( .C1(n4485), .C2(n9863), .A(n9142), .B(n9141), .ZN(
        P1_U3228) );
  INV_X1 U10504 ( .A(n9624), .ZN(n9821) );
  INV_X1 U10505 ( .A(n9143), .ZN(n9145) );
  NOR3_X1 U10506 ( .A1(n9146), .A2(n9145), .A3(n9144), .ZN(n9149) );
  INV_X1 U10507 ( .A(n9147), .ZN(n9148) );
  OAI21_X1 U10508 ( .B1(n9149), .B2(n9148), .A(n9865), .ZN(n9155) );
  INV_X1 U10509 ( .A(n9150), .ZN(n9625) );
  AND2_X1 U10510 ( .A1(n9448), .A2(n9291), .ZN(n9151) );
  AOI21_X1 U10511 ( .B1(n9446), .B2(n9169), .A(n9151), .ZN(n9621) );
  OAI22_X1 U10512 ( .A1(n9621), .A2(n9183), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9152), .ZN(n9153) );
  AOI21_X1 U10513 ( .B1(n9625), .B2(n9162), .A(n9153), .ZN(n9154) );
  OAI211_X1 U10514 ( .C1(n9821), .C2(n9863), .A(n9155), .B(n9154), .ZN(
        P1_U3229) );
  OAI21_X1 U10515 ( .B1(n9158), .B2(n9157), .A(n9156), .ZN(n9159) );
  NAND2_X1 U10516 ( .A1(n9159), .A2(n9865), .ZN(n9164) );
  AOI22_X1 U10517 ( .A1(n9450), .A2(n9169), .B1(n9291), .B2(n9451), .ZN(n9676)
         );
  OAI22_X1 U10518 ( .A1(n9676), .A2(n9183), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9160), .ZN(n9161) );
  AOI21_X1 U10519 ( .B1(n9683), .B2(n9162), .A(n9161), .ZN(n9163) );
  OAI211_X1 U10520 ( .C1(n9781), .C2(n9863), .A(n9164), .B(n9163), .ZN(
        P1_U3233) );
  INV_X1 U10521 ( .A(n9082), .ZN(n9165) );
  AOI21_X1 U10522 ( .B1(n9167), .B2(n9166), .A(n9165), .ZN(n9174) );
  NOR2_X1 U10523 ( .A1(n9868), .A2(n9648), .ZN(n9172) );
  AND2_X1 U10524 ( .A1(n9450), .A2(n9291), .ZN(n9168) );
  AOI21_X1 U10525 ( .B1(n9448), .B2(n9169), .A(n9168), .ZN(n9654) );
  OAI22_X1 U10526 ( .A1(n9654), .A2(n9183), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9170), .ZN(n9171) );
  AOI211_X1 U10527 ( .C1(n9647), .C2(n9186), .A(n9172), .B(n9171), .ZN(n9173)
         );
  OAI21_X1 U10528 ( .B1(n9174), .B2(n9188), .A(n9173), .ZN(P1_U3235) );
  INV_X1 U10529 ( .A(n9175), .ZN(n9177) );
  NAND2_X1 U10530 ( .A1(n9177), .A2(n9176), .ZN(n9178) );
  XNOR2_X1 U10531 ( .A(n9179), .B(n9178), .ZN(n9189) );
  NOR2_X1 U10532 ( .A1(n9868), .A2(n9712), .ZN(n9185) );
  AND2_X1 U10533 ( .A1(n9453), .A2(n9291), .ZN(n9180) );
  AOI21_X1 U10534 ( .B1(n9451), .B2(n9181), .A(n9180), .ZN(n9707) );
  OAI22_X1 U10535 ( .A1(n9183), .A2(n9707), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9182), .ZN(n9184) );
  AOI211_X1 U10536 ( .C1(n9793), .C2(n9186), .A(n9185), .B(n9184), .ZN(n9187)
         );
  OAI21_X1 U10537 ( .B1(n9189), .B2(n9188), .A(n9187), .ZN(P1_U3238) );
  OAI21_X1 U10538 ( .B1(n9192), .B2(n9191), .A(n9190), .ZN(n9193) );
  NAND2_X1 U10539 ( .A1(n9193), .A2(n9865), .ZN(n9198) );
  AND2_X1 U10540 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9491) );
  NOR2_X1 U10541 ( .A1(n9868), .A2(n9194), .ZN(n9195) );
  AOI211_X1 U10542 ( .C1(n9861), .C2(n9196), .A(n9491), .B(n9195), .ZN(n9197)
         );
  OAI211_X1 U10543 ( .C1(n4701), .C2(n9863), .A(n9198), .B(n9197), .ZN(
        P1_U3241) );
  NAND2_X1 U10544 ( .A1(n9199), .A2(n5114), .ZN(n9201) );
  NAND2_X1 U10545 ( .A1(n4997), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n9200) );
  INV_X1 U10546 ( .A(n9806), .ZN(n9282) );
  INV_X1 U10547 ( .A(n9417), .ZN(n9370) );
  MUX2_X1 U10548 ( .A(n9624), .B(n9447), .S(n9278), .Z(n9260) );
  NAND2_X1 U10549 ( .A1(n9245), .A2(n9239), .ZN(n9244) );
  INV_X1 U10550 ( .A(n9204), .ZN(n9947) );
  NOR2_X1 U10551 ( .A1(n9947), .A2(n9946), .ZN(n9944) );
  INV_X1 U10552 ( .A(n9389), .ZN(n9206) );
  OAI21_X1 U10553 ( .B1(n9944), .B2(n9206), .A(n9205), .ZN(n9207) );
  INV_X1 U10554 ( .A(n9208), .ZN(n9209) );
  NAND2_X1 U10555 ( .A1(n9223), .A2(n9218), .ZN(n9345) );
  AOI21_X1 U10556 ( .B1(n9210), .B2(n9346), .A(n9345), .ZN(n9211) );
  INV_X1 U10557 ( .A(n9221), .ZN(n9349) );
  INV_X1 U10558 ( .A(n9357), .ZN(n9212) );
  AOI21_X1 U10559 ( .B1(n9213), .B2(n9353), .A(n9212), .ZN(n9235) );
  INV_X1 U10560 ( .A(n9214), .ZN(n9216) );
  NAND3_X1 U10561 ( .A1(n9219), .A2(n9342), .A3(n9218), .ZN(n9222) );
  NAND3_X1 U10562 ( .A1(n9222), .A2(n9221), .A3(n9220), .ZN(n9224) );
  NAND2_X1 U10563 ( .A1(n9224), .A2(n9223), .ZN(n9225) );
  AOI21_X1 U10564 ( .B1(n9225), .B2(n9348), .A(n4845), .ZN(n9231) );
  NAND2_X1 U10565 ( .A1(n9227), .A2(n9226), .ZN(n9354) );
  OR2_X1 U10566 ( .A1(n9354), .A2(n9228), .ZN(n9230) );
  AND2_X1 U10567 ( .A1(n9230), .A2(n9229), .ZN(n9356) );
  OAI21_X1 U10568 ( .B1(n9231), .B2(n9354), .A(n9356), .ZN(n9233) );
  INV_X1 U10569 ( .A(n9353), .ZN(n9232) );
  AOI21_X1 U10570 ( .B1(n9233), .B2(n9357), .A(n9232), .ZN(n9234) );
  MUX2_X1 U10571 ( .A(n9235), .B(n9234), .S(n9278), .Z(n9237) );
  INV_X1 U10572 ( .A(n9402), .ZN(n9236) );
  NAND2_X1 U10573 ( .A1(n9241), .A2(n9238), .ZN(n9360) );
  NAND2_X1 U10574 ( .A1(n9239), .A2(n9240), .ZN(n9364) );
  NAND2_X1 U10575 ( .A1(n9304), .A2(n9245), .ZN(n9320) );
  NAND2_X1 U10576 ( .A1(n9247), .A2(n9246), .ZN(n9305) );
  MUX2_X1 U10577 ( .A(n9320), .B(n9305), .S(n9278), .Z(n9249) );
  MUX2_X1 U10578 ( .A(n9247), .B(n9304), .S(n9278), .Z(n9248) );
  OAI21_X1 U10579 ( .B1(n9250), .B2(n9249), .A(n9248), .ZN(n9255) );
  NAND2_X1 U10580 ( .A1(n9300), .A2(n9251), .ZN(n9307) );
  OR2_X1 U10581 ( .A1(n9824), .A2(n9252), .ZN(n9256) );
  NAND2_X1 U10582 ( .A1(n9256), .A2(n9253), .ZN(n9299) );
  MUX2_X1 U10583 ( .A(n9307), .B(n9299), .S(n9278), .Z(n9254) );
  INV_X1 U10584 ( .A(n9256), .ZN(n9258) );
  INV_X1 U10585 ( .A(n9300), .ZN(n9257) );
  MUX2_X1 U10586 ( .A(n9258), .B(n9257), .S(n9278), .Z(n9259) );
  INV_X1 U10587 ( .A(n9266), .ZN(n9263) );
  INV_X1 U10588 ( .A(n9310), .ZN(n9377) );
  NOR2_X1 U10589 ( .A1(n9812), .A2(n9262), .ZN(n9312) );
  NOR2_X1 U10590 ( .A1(n9312), .A2(n9378), .ZN(n9265) );
  OAI21_X1 U10591 ( .B1(n9263), .B2(n9377), .A(n9265), .ZN(n9264) );
  NAND2_X1 U10592 ( .A1(n9267), .A2(n9317), .ZN(n9269) );
  INV_X1 U10593 ( .A(n9315), .ZN(n9268) );
  NOR2_X1 U10594 ( .A1(n9444), .A2(n9278), .ZN(n9270) );
  NAND2_X1 U10595 ( .A1(n9583), .A2(n9270), .ZN(n9271) );
  OAI21_X1 U10596 ( .B1(n9278), .B2(n9443), .A(n9271), .ZN(n9274) );
  INV_X1 U10597 ( .A(n9271), .ZN(n9273) );
  AOI22_X1 U10598 ( .A1(n9568), .A2(n9274), .B1(n9273), .B2(n9272), .ZN(n9275)
         );
  MUX2_X1 U10599 ( .A(n9327), .B(n9366), .S(n9278), .Z(n9276) );
  INV_X1 U10600 ( .A(n9368), .ZN(n9441) );
  AOI21_X1 U10601 ( .B1(n9441), .B2(n9425), .A(n9427), .ZN(n9279) );
  MUX2_X1 U10602 ( .A(n4552), .B(n9281), .S(n9741), .Z(n9283) );
  NAND3_X1 U10603 ( .A1(n9283), .A2(n9441), .A3(n9282), .ZN(n9284) );
  NAND2_X1 U10604 ( .A1(n9285), .A2(n9284), .ZN(n9297) );
  OAI21_X1 U10605 ( .B1(n9370), .B2(n4552), .A(n9297), .ZN(n9288) );
  AOI21_X1 U10606 ( .B1(n9427), .B2(n9549), .A(n9286), .ZN(n9287) );
  OR2_X1 U10607 ( .A1(n9416), .A2(n9296), .ZN(n9289) );
  AOI21_X1 U10608 ( .B1(n9288), .B2(n9287), .A(n9289), .ZN(n9440) );
  INV_X1 U10609 ( .A(n9289), .ZN(n9294) );
  NAND3_X1 U10610 ( .A1(n9291), .A2(n9290), .A3(n9896), .ZN(n9293) );
  OAI22_X1 U10611 ( .A1(n9294), .A2(P1_B_REG_SCAN_IN), .B1(n9293), .B2(n9292), 
        .ZN(n9439) );
  INV_X1 U10612 ( .A(n9298), .ZN(n9375) );
  NAND2_X1 U10613 ( .A1(n9549), .A2(n9375), .ZN(n9414) );
  NAND2_X1 U10614 ( .A1(n9549), .A2(n9298), .ZN(n9374) );
  NAND3_X1 U10615 ( .A1(n9309), .A2(n9300), .A3(n9299), .ZN(n9302) );
  NAND2_X1 U10616 ( .A1(n9302), .A2(n9301), .ZN(n9303) );
  OR2_X1 U10617 ( .A1(n9378), .A2(n9303), .ZN(n9319) );
  AND2_X1 U10618 ( .A1(n9305), .A2(n9304), .ZN(n9306) );
  NOR2_X1 U10619 ( .A1(n9307), .A2(n9306), .ZN(n9308) );
  AND2_X1 U10620 ( .A1(n9309), .A2(n9308), .ZN(n9311) );
  OAI21_X1 U10621 ( .B1(n9319), .B2(n9311), .A(n9310), .ZN(n9313) );
  INV_X1 U10622 ( .A(n9312), .ZN(n9321) );
  NAND3_X1 U10623 ( .A1(n9313), .A2(n9321), .A3(n9325), .ZN(n9314) );
  NAND3_X1 U10624 ( .A1(n9316), .A2(n9315), .A3(n9314), .ZN(n9326) );
  INV_X1 U10625 ( .A(n9317), .ZN(n9318) );
  NOR2_X1 U10626 ( .A1(n9326), .A2(n9318), .ZN(n9418) );
  INV_X1 U10627 ( .A(n9319), .ZN(n9323) );
  INV_X1 U10628 ( .A(n9320), .ZN(n9322) );
  NAND3_X1 U10629 ( .A1(n9323), .A2(n9322), .A3(n9321), .ZN(n9330) );
  OAI21_X1 U10630 ( .B1(n9326), .B2(n9325), .A(n9324), .ZN(n9329) );
  INV_X1 U10631 ( .A(n9327), .ZN(n9328) );
  AOI211_X1 U10632 ( .C1(n9418), .C2(n9330), .A(n9329), .B(n9328), .ZN(n9419)
         );
  INV_X1 U10633 ( .A(n9331), .ZN(n9335) );
  NAND3_X1 U10634 ( .A1(n9333), .A2(n9332), .A3(n5670), .ZN(n9334) );
  AOI211_X1 U10635 ( .C1(n9336), .C2(n9468), .A(n9335), .B(n9334), .ZN(n9339)
         );
  NAND3_X1 U10636 ( .A1(n9339), .A2(n9338), .A3(n9337), .ZN(n9340) );
  NAND2_X1 U10637 ( .A1(n7358), .A2(n9340), .ZN(n9344) );
  OAI211_X1 U10638 ( .C1(n9344), .C2(n9343), .A(n9342), .B(n9341), .ZN(n9347)
         );
  AOI21_X1 U10639 ( .B1(n9347), .B2(n9346), .A(n9345), .ZN(n9350) );
  NOR3_X1 U10640 ( .A1(n9350), .A2(n9349), .A3(n5569), .ZN(n9352) );
  NOR2_X1 U10641 ( .A1(n9352), .A2(n4848), .ZN(n9355) );
  OAI21_X1 U10642 ( .B1(n9355), .B2(n9354), .A(n9353), .ZN(n9359) );
  INV_X1 U10643 ( .A(n9356), .ZN(n9358) );
  OAI21_X1 U10644 ( .B1(n9359), .B2(n9358), .A(n9357), .ZN(n9361) );
  AOI21_X1 U10645 ( .B1(n9362), .B2(n9361), .A(n9360), .ZN(n9365) );
  OAI211_X1 U10646 ( .C1(n9365), .C2(n9364), .A(n9418), .B(n9363), .ZN(n9367)
         );
  NAND2_X1 U10647 ( .A1(n9741), .A2(n9368), .ZN(n9408) );
  NAND2_X1 U10648 ( .A1(n9408), .A2(n9366), .ZN(n9421) );
  AOI21_X1 U10649 ( .B1(n9419), .B2(n9367), .A(n9421), .ZN(n9369) );
  NOR2_X1 U10650 ( .A1(n9741), .A2(n9368), .ZN(n9426) );
  NOR2_X1 U10651 ( .A1(n9369), .A2(n9426), .ZN(n9371) );
  OAI21_X1 U10652 ( .B1(n9371), .B2(n9427), .A(n9370), .ZN(n9372) );
  MUX2_X1 U10653 ( .A(n9374), .B(n9373), .S(n9372), .Z(n9436) );
  AND2_X1 U10654 ( .A1(n9376), .A2(n9375), .ZN(n9431) );
  INV_X1 U10655 ( .A(n9427), .ZN(n9413) );
  INV_X1 U10656 ( .A(n9426), .ZN(n9410) );
  OR2_X1 U10657 ( .A1(n9378), .A2(n9377), .ZN(n9605) );
  INV_X1 U10658 ( .A(n9633), .ZN(n9631) );
  INV_X1 U10659 ( .A(n9703), .ZN(n9705) );
  NOR2_X1 U10660 ( .A1(n9379), .A2(n5670), .ZN(n9382) );
  NAND4_X1 U10661 ( .A1(n9382), .A2(n4543), .A3(n9381), .A4(n9380), .ZN(n9385)
         );
  NOR3_X1 U10662 ( .A1(n9385), .A2(n9384), .A3(n9383), .ZN(n9387) );
  NAND4_X1 U10663 ( .A1(n9389), .A2(n9388), .A3(n9387), .A4(n9386), .ZN(n9390)
         );
  NOR2_X1 U10664 ( .A1(n9391), .A2(n9390), .ZN(n9393) );
  NAND4_X1 U10665 ( .A1(n9394), .A2(n4688), .A3(n9393), .A4(n9392), .ZN(n9395)
         );
  NOR2_X1 U10666 ( .A1(n9396), .A2(n9395), .ZN(n9397) );
  AND4_X1 U10667 ( .A1(n9400), .A2(n9399), .A3(n9398), .A4(n9397), .ZN(n9401)
         );
  AND4_X1 U10668 ( .A1(n9695), .A2(n9402), .A3(n9705), .A4(n9401), .ZN(n9403)
         );
  NAND4_X1 U10669 ( .A1(n9653), .A2(n4718), .A3(n9680), .A4(n9403), .ZN(n9404)
         );
  OR3_X1 U10670 ( .A1(n9619), .A2(n9631), .A3(n9404), .ZN(n9405) );
  NOR2_X1 U10671 ( .A1(n9605), .A2(n9405), .ZN(n9406) );
  AND4_X1 U10672 ( .A1(n9407), .A2(n9580), .A3(n9406), .A4(n9594), .ZN(n9409)
         );
  AND4_X1 U10673 ( .A1(n9411), .A2(n9410), .A3(n9409), .A4(n9408), .ZN(n9412)
         );
  NAND2_X1 U10674 ( .A1(n9413), .A2(n9412), .ZN(n9430) );
  NOR3_X1 U10675 ( .A1(n9430), .A2(n9417), .A3(n9414), .ZN(n9415) );
  AOI211_X1 U10676 ( .C1(n9417), .C2(n9431), .A(n9416), .B(n9415), .ZN(n9435)
         );
  INV_X1 U10677 ( .A(n9741), .ZN(n9424) );
  INV_X1 U10678 ( .A(n9418), .ZN(n9420) );
  OAI21_X1 U10679 ( .B1(n9420), .B2(n9675), .A(n9419), .ZN(n9423) );
  INV_X1 U10680 ( .A(n9421), .ZN(n9422) );
  OAI211_X1 U10681 ( .C1(n9424), .C2(n9425), .A(n9423), .B(n9422), .ZN(n9429)
         );
  NAND2_X1 U10682 ( .A1(n9426), .A2(n9425), .ZN(n9428) );
  AOI21_X1 U10683 ( .B1(n9429), .B2(n9428), .A(n9427), .ZN(n9433) );
  OAI211_X1 U10684 ( .C1(n9433), .C2(n9432), .A(n9431), .B(n9430), .ZN(n9434)
         );
  NAND3_X1 U10685 ( .A1(n9436), .A2(n9435), .A3(n9434), .ZN(n9437) );
  OAI22_X1 U10686 ( .A1(n9440), .A2(n9439), .B1(n9438), .B2(n9437), .ZN(
        P1_U3242) );
  MUX2_X1 U10687 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9441), .S(P1_U3973), .Z(
        P1_U3584) );
  MUX2_X1 U10688 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9442), .S(P1_U3973), .Z(
        P1_U3583) );
  MUX2_X1 U10689 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9443), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U10690 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9444), .S(P1_U3973), .Z(
        P1_U3581) );
  MUX2_X1 U10691 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9445), .S(P1_U3973), .Z(
        P1_U3580) );
  MUX2_X1 U10692 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9446), .S(P1_U3973), .Z(
        P1_U3579) );
  MUX2_X1 U10693 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9447), .S(P1_U3973), .Z(
        P1_U3578) );
  MUX2_X1 U10694 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9448), .S(P1_U3973), .Z(
        P1_U3577) );
  MUX2_X1 U10695 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9449), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U10696 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9450), .S(P1_U3973), .Z(
        P1_U3575) );
  MUX2_X1 U10697 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9451), .S(P1_U3973), .Z(
        P1_U3573) );
  MUX2_X1 U10698 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9452), .S(P1_U3973), .Z(
        P1_U3572) );
  MUX2_X1 U10699 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9453), .S(P1_U3973), .Z(
        P1_U3571) );
  MUX2_X1 U10700 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9454), .S(P1_U3973), .Z(
        P1_U3570) );
  MUX2_X1 U10701 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9455), .S(P1_U3973), .Z(
        P1_U3569) );
  MUX2_X1 U10702 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9456), .S(P1_U3973), .Z(
        P1_U3568) );
  MUX2_X1 U10703 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9457), .S(P1_U3973), .Z(
        P1_U3567) );
  MUX2_X1 U10704 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9458), .S(P1_U3973), .Z(
        P1_U3566) );
  MUX2_X1 U10705 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9459), .S(P1_U3973), .Z(
        P1_U3565) );
  MUX2_X1 U10706 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9460), .S(P1_U3973), .Z(
        P1_U3564) );
  MUX2_X1 U10707 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9461), .S(P1_U3973), .Z(
        P1_U3563) );
  MUX2_X1 U10708 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9462), .S(P1_U3973), .Z(
        P1_U3562) );
  MUX2_X1 U10709 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9463), .S(P1_U3973), .Z(
        P1_U3561) );
  MUX2_X1 U10710 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9464), .S(P1_U3973), .Z(
        P1_U3560) );
  MUX2_X1 U10711 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9465), .S(P1_U3973), .Z(
        P1_U3559) );
  MUX2_X1 U10712 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9466), .S(P1_U3973), .Z(
        P1_U3558) );
  MUX2_X1 U10713 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9467), .S(P1_U3973), .Z(
        P1_U3557) );
  MUX2_X1 U10714 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n9468), .S(P1_U3973), .Z(
        P1_U3556) );
  MUX2_X1 U10715 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n9469), .S(P1_U3973), .Z(
        P1_U3555) );
  INV_X1 U10716 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9471) );
  OAI22_X1 U10717 ( .A1(n9553), .A2(n9471), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9470), .ZN(n9472) );
  AOI21_X1 U10718 ( .B1(n9473), .B2(n9937), .A(n9472), .ZN(n9481) );
  OAI211_X1 U10719 ( .C1(n9476), .C2(n9475), .A(n9939), .B(n9474), .ZN(n9480)
         );
  OAI211_X1 U10720 ( .C1(n9478), .C2(n9897), .A(n9915), .B(n9477), .ZN(n9479)
         );
  NAND3_X1 U10721 ( .A1(n9481), .A2(n9480), .A3(n9479), .ZN(P1_U3244) );
  NOR2_X1 U10722 ( .A1(n7774), .A2(n9485), .ZN(n9507) );
  INV_X1 U10723 ( .A(n9507), .ZN(n9483) );
  NAND2_X1 U10724 ( .A1(n9915), .A2(n9483), .ZN(n9484) );
  AOI21_X1 U10725 ( .B1(n9485), .B2(n7774), .A(n9484), .ZN(n9497) );
  NOR2_X1 U10726 ( .A1(n9489), .A2(n9488), .ZN(n9499) );
  AOI211_X1 U10727 ( .C1(n9489), .C2(n9488), .A(n9499), .B(n9919), .ZN(n9496)
         );
  INV_X1 U10728 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n9494) );
  NAND2_X1 U10729 ( .A1(n9937), .A2(n9490), .ZN(n9493) );
  INV_X1 U10730 ( .A(n9491), .ZN(n9492) );
  OAI211_X1 U10731 ( .C1(n9494), .C2(n9553), .A(n9493), .B(n9492), .ZN(n9495)
         );
  OR3_X1 U10732 ( .A1(n9497), .A2(n9496), .A3(n9495), .ZN(P1_U3258) );
  XOR2_X1 U10733 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9519), .Z(n9528) );
  NOR2_X1 U10734 ( .A1(n9498), .A2(n9505), .ZN(n9500) );
  NOR2_X1 U10735 ( .A1(n9500), .A2(n9499), .ZN(n9936) );
  NOR2_X1 U10736 ( .A1(n9503), .A2(n9501), .ZN(n9502) );
  AOI21_X1 U10737 ( .B1(n9501), .B2(n9503), .A(n9502), .ZN(n9935) );
  NAND2_X1 U10738 ( .A1(n9936), .A2(n9935), .ZN(n9934) );
  OAI21_X1 U10739 ( .B1(n9938), .B2(P1_REG1_REG_16__SCAN_IN), .A(n9934), .ZN(
        n9529) );
  XOR2_X1 U10740 ( .A(n9528), .B(n9529), .Z(n9518) );
  XNOR2_X1 U10741 ( .A(n9519), .B(n9504), .ZN(n9511) );
  NOR2_X1 U10742 ( .A1(n9506), .A2(n9505), .ZN(n9508) );
  XNOR2_X1 U10743 ( .A(n9938), .B(P1_REG2_REG_16__SCAN_IN), .ZN(n9929) );
  NAND2_X1 U10744 ( .A1(n9938), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n9509) );
  NAND2_X1 U10745 ( .A1(n9510), .A2(n9511), .ZN(n9521) );
  OAI21_X1 U10746 ( .B1(n9511), .B2(n9510), .A(n9521), .ZN(n9512) );
  NAND2_X1 U10747 ( .A1(n9512), .A2(n9915), .ZN(n9517) );
  INV_X1 U10748 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9514) );
  OAI21_X1 U10749 ( .B1(n9553), .B2(n9514), .A(n9513), .ZN(n9515) );
  AOI21_X1 U10750 ( .B1(n9519), .B2(n9937), .A(n9515), .ZN(n9516) );
  OAI211_X1 U10751 ( .C1(n9919), .C2(n9518), .A(n9517), .B(n9516), .ZN(
        P1_U3260) );
  OR2_X1 U10752 ( .A1(n9519), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9520) );
  NAND2_X1 U10753 ( .A1(n9530), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9538) );
  OR2_X1 U10754 ( .A1(n9530), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9522) );
  AND2_X1 U10755 ( .A1(n9538), .A2(n9522), .ZN(n9523) );
  OAI211_X1 U10756 ( .C1(n9524), .C2(n9523), .A(n9539), .B(n9915), .ZN(n9537)
         );
  NAND2_X1 U10757 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_U3086), .ZN(n9525) );
  OAI21_X1 U10758 ( .B1(n9553), .B2(n10159), .A(n9525), .ZN(n9526) );
  AOI21_X1 U10759 ( .B1(n9530), .B2(n9937), .A(n9526), .ZN(n9536) );
  INV_X1 U10760 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9799) );
  AOI22_X1 U10761 ( .A1(n9529), .A2(n9528), .B1(n9527), .B2(n9799), .ZN(n9534)
         );
  INV_X1 U10762 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9532) );
  AND2_X1 U10763 ( .A1(n9530), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9541) );
  AOI21_X1 U10764 ( .B1(n9532), .B2(n9531), .A(n9541), .ZN(n9533) );
  NAND2_X1 U10765 ( .A1(n9534), .A2(n9533), .ZN(n9543) );
  OAI211_X1 U10766 ( .C1(n9534), .C2(n9533), .A(n9543), .B(n9939), .ZN(n9535)
         );
  NAND3_X1 U10767 ( .A1(n9537), .A2(n9536), .A3(n9535), .ZN(P1_U3261) );
  NAND2_X1 U10768 ( .A1(n9539), .A2(n9538), .ZN(n9540) );
  INV_X1 U10769 ( .A(n9548), .ZN(n9545) );
  INV_X1 U10770 ( .A(n9541), .ZN(n9542) );
  NAND2_X1 U10771 ( .A1(n9543), .A2(n9542), .ZN(n9544) );
  XOR2_X1 U10772 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9544), .Z(n9546) );
  AOI22_X1 U10773 ( .A1(n9545), .A2(n9915), .B1(n9939), .B2(n9546), .ZN(n9551)
         );
  NOR2_X1 U10774 ( .A1(n9546), .A2(n9919), .ZN(n9547) );
  NAND2_X1 U10775 ( .A1(P1_REG3_REG_19__SCAN_IN), .A2(P1_U3086), .ZN(n9552) );
  XNOR2_X1 U10776 ( .A(n9806), .B(n9554), .ZN(n9555) );
  NAND2_X1 U10777 ( .A1(n9736), .A2(n9960), .ZN(n9558) );
  NOR2_X1 U10778 ( .A1(n4334), .A2(n9556), .ZN(n9560) );
  AOI21_X1 U10779 ( .B1(n4334), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9560), .ZN(
        n9557) );
  OAI211_X1 U10780 ( .C1(n9806), .C2(n9716), .A(n9558), .B(n9557), .ZN(
        P1_U3263) );
  NOR2_X1 U10781 ( .A1(n9723), .A2(n9559), .ZN(n9561) );
  AOI211_X1 U10782 ( .C1(n9741), .C2(n9953), .A(n9561), .B(n9560), .ZN(n9562)
         );
  OAI21_X1 U10783 ( .B1(n9563), .B2(n9671), .A(n9562), .ZN(P1_U3264) );
  INV_X1 U10784 ( .A(n9564), .ZN(n9572) );
  OAI22_X1 U10785 ( .A1(n9566), .A2(n9727), .B1(n9565), .B2(n9723), .ZN(n9567)
         );
  AOI21_X1 U10786 ( .B1(n9568), .B2(n9953), .A(n9567), .ZN(n9569) );
  OAI21_X1 U10787 ( .B1(n9570), .B2(n9671), .A(n9569), .ZN(n9571) );
  AOI21_X1 U10788 ( .B1(n9572), .B2(n9721), .A(n9571), .ZN(n9573) );
  OAI21_X1 U10789 ( .B1(n4334), .B2(n9574), .A(n9573), .ZN(P1_U3265) );
  OAI21_X1 U10790 ( .B1(n9580), .B2(n9576), .A(n9575), .ZN(n9577) );
  NAND2_X1 U10791 ( .A1(n9577), .A2(n9698), .ZN(n9579) );
  NAND2_X1 U10792 ( .A1(n9579), .A2(n9578), .ZN(n9743) );
  INV_X1 U10793 ( .A(n9743), .ZN(n9589) );
  XNOR2_X1 U10794 ( .A(n9581), .B(n9580), .ZN(n9745) );
  AOI211_X1 U10795 ( .C1(n9583), .C2(n9595), .A(n9977), .B(n4491), .ZN(n9744)
         );
  NAND2_X1 U10796 ( .A1(n9744), .A2(n9960), .ZN(n9586) );
  AOI22_X1 U10797 ( .A1(n9584), .A2(n9951), .B1(P1_REG2_REG_27__SCAN_IN), .B2(
        n4334), .ZN(n9585) );
  OAI211_X1 U10798 ( .C1(n4493), .C2(n9716), .A(n9586), .B(n9585), .ZN(n9587)
         );
  AOI21_X1 U10799 ( .B1(n9745), .B2(n9721), .A(n9587), .ZN(n9588) );
  OAI21_X1 U10800 ( .B1(n4334), .B2(n9589), .A(n9588), .ZN(P1_U3266) );
  XNOR2_X1 U10801 ( .A(n9590), .B(n9594), .ZN(n9592) );
  AOI21_X1 U10802 ( .B1(n9592), .B2(n9698), .A(n9591), .ZN(n9749) );
  XNOR2_X1 U10803 ( .A(n9593), .B(n9594), .ZN(n9750) );
  INV_X1 U10804 ( .A(n9750), .ZN(n9602) );
  OAI211_X1 U10805 ( .C1(n9596), .C2(n9610), .A(n9957), .B(n9595), .ZN(n9748)
         );
  INV_X1 U10806 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n9597) );
  OAI22_X1 U10807 ( .A1(n9598), .A2(n9727), .B1(n9597), .B2(n9723), .ZN(n9599)
         );
  AOI21_X1 U10808 ( .B1(n9812), .B2(n9953), .A(n9599), .ZN(n9600) );
  OAI21_X1 U10809 ( .B1(n9748), .B2(n9671), .A(n9600), .ZN(n9601) );
  AOI21_X1 U10810 ( .B1(n9602), .B2(n9721), .A(n9601), .ZN(n9603) );
  OAI21_X1 U10811 ( .B1(n4334), .B2(n9749), .A(n9603), .ZN(P1_U3267) );
  XOR2_X1 U10812 ( .A(n9605), .B(n9604), .Z(n9755) );
  INV_X1 U10813 ( .A(n9755), .ZN(n9617) );
  XOR2_X1 U10814 ( .A(n9606), .B(n9605), .Z(n9609) );
  INV_X1 U10815 ( .A(n9607), .ZN(n9608) );
  OAI21_X1 U10816 ( .B1(n9609), .B2(n9945), .A(n9608), .ZN(n9753) );
  AOI211_X1 U10817 ( .C1(n9611), .C2(n9623), .A(n9977), .B(n9610), .ZN(n9754)
         );
  NAND2_X1 U10818 ( .A1(n9754), .A2(n9960), .ZN(n9614) );
  AOI22_X1 U10819 ( .A1(n9612), .A2(n9951), .B1(P1_REG2_REG_25__SCAN_IN), .B2(
        n4334), .ZN(n9613) );
  OAI211_X1 U10820 ( .C1(n9817), .C2(n9716), .A(n9614), .B(n9613), .ZN(n9615)
         );
  AOI21_X1 U10821 ( .B1(n9753), .B2(n9723), .A(n9615), .ZN(n9616) );
  OAI21_X1 U10822 ( .B1(n9617), .B2(n9720), .A(n9616), .ZN(P1_U3268) );
  XNOR2_X1 U10823 ( .A(n9618), .B(n9619), .ZN(n9760) );
  INV_X1 U10824 ( .A(n9760), .ZN(n9630) );
  OAI211_X1 U10825 ( .C1(n4376), .C2(n4864), .A(n9620), .B(n9698), .ZN(n9622)
         );
  NAND2_X1 U10826 ( .A1(n9622), .A2(n9621), .ZN(n9758) );
  AOI211_X1 U10827 ( .C1(n9624), .C2(n9637), .A(n9977), .B(n5590), .ZN(n9759)
         );
  NAND2_X1 U10828 ( .A1(n9759), .A2(n9960), .ZN(n9627) );
  AOI22_X1 U10829 ( .A1(n9625), .A2(n9951), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n4334), .ZN(n9626) );
  OAI211_X1 U10830 ( .C1(n9821), .C2(n9716), .A(n9627), .B(n9626), .ZN(n9628)
         );
  AOI21_X1 U10831 ( .B1(n9723), .B2(n9758), .A(n9628), .ZN(n9629) );
  OAI21_X1 U10832 ( .B1(n9630), .B2(n9720), .A(n9629), .ZN(P1_U3269) );
  XNOR2_X1 U10833 ( .A(n9632), .B(n9631), .ZN(n9765) );
  XNOR2_X1 U10834 ( .A(n9634), .B(n9633), .ZN(n9636) );
  AOI21_X1 U10835 ( .B1(n9636), .B2(n9698), .A(n9635), .ZN(n9764) );
  INV_X1 U10836 ( .A(n9764), .ZN(n9644) );
  OAI211_X1 U10837 ( .C1(n9638), .C2(n4404), .A(n9957), .B(n9637), .ZN(n9763)
         );
  INV_X1 U10838 ( .A(n9639), .ZN(n9640) );
  AOI22_X1 U10839 ( .A1(n9640), .A2(n9951), .B1(P1_REG2_REG_23__SCAN_IN), .B2(
        n4334), .ZN(n9642) );
  NAND2_X1 U10840 ( .A1(n9824), .A2(n9953), .ZN(n9641) );
  OAI211_X1 U10841 ( .C1(n9763), .C2(n9671), .A(n9642), .B(n9641), .ZN(n9643)
         );
  AOI21_X1 U10842 ( .B1(n9644), .B2(n9723), .A(n9643), .ZN(n9645) );
  OAI21_X1 U10843 ( .B1(n9765), .B2(n9720), .A(n9645), .ZN(P1_U3270) );
  XNOR2_X1 U10844 ( .A(n9646), .B(n9653), .ZN(n9770) );
  INV_X1 U10845 ( .A(n9770), .ZN(n9658) );
  AOI211_X1 U10846 ( .C1(n9647), .C2(n4903), .A(n9977), .B(n4404), .ZN(n9769)
         );
  NOR2_X1 U10847 ( .A1(n4482), .A2(n9716), .ZN(n9651) );
  OAI22_X1 U10848 ( .A1(n9723), .A2(n9649), .B1(n9648), .B2(n9727), .ZN(n9650)
         );
  AOI211_X1 U10849 ( .C1(n9769), .C2(n9960), .A(n9651), .B(n9650), .ZN(n9657)
         );
  XOR2_X1 U10850 ( .A(n9653), .B(n9652), .Z(n9655) );
  OAI21_X1 U10851 ( .B1(n9655), .B2(n9945), .A(n9654), .ZN(n9768) );
  NAND2_X1 U10852 ( .A1(n9768), .A2(n9723), .ZN(n9656) );
  OAI211_X1 U10853 ( .C1(n9658), .C2(n9720), .A(n9657), .B(n9656), .ZN(
        P1_U3271) );
  XNOR2_X1 U10854 ( .A(n9659), .B(n9662), .ZN(n9661) );
  AOI21_X1 U10855 ( .B1(n9661), .B2(n9698), .A(n9660), .ZN(n9774) );
  OR2_X1 U10856 ( .A1(n9663), .A2(n9662), .ZN(n9664) );
  NAND2_X1 U10857 ( .A1(n9665), .A2(n9664), .ZN(n9775) );
  INV_X1 U10858 ( .A(n9775), .ZN(n9673) );
  AOI21_X1 U10859 ( .B1(n9831), .B2(n9682), .A(n9977), .ZN(n9666) );
  NAND2_X1 U10860 ( .A1(n9666), .A2(n4903), .ZN(n9773) );
  NAND2_X1 U10861 ( .A1(n4334), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n9667) );
  OAI21_X1 U10862 ( .B1(n9727), .B2(n9668), .A(n9667), .ZN(n9669) );
  AOI21_X1 U10863 ( .B1(n9831), .B2(n9953), .A(n9669), .ZN(n9670) );
  OAI21_X1 U10864 ( .B1(n9773), .B2(n9671), .A(n9670), .ZN(n9672) );
  AOI21_X1 U10865 ( .B1(n9673), .B2(n9721), .A(n9672), .ZN(n9674) );
  OAI21_X1 U10866 ( .B1(n4334), .B2(n9774), .A(n9674), .ZN(P1_U3272) );
  AOI21_X1 U10867 ( .B1(n9675), .B2(n5372), .A(n9945), .ZN(n9679) );
  INV_X1 U10868 ( .A(n9676), .ZN(n9677) );
  AOI21_X1 U10869 ( .B1(n9679), .B2(n9678), .A(n9677), .ZN(n9784) );
  NAND2_X1 U10870 ( .A1(n9681), .A2(n9680), .ZN(n9779) );
  NAND3_X1 U10871 ( .A1(n9780), .A2(n9779), .A3(n9721), .ZN(n9688) );
  OAI211_X1 U10872 ( .C1(n9781), .C2(n9690), .A(n9957), .B(n9682), .ZN(n9783)
         );
  INV_X1 U10873 ( .A(n9783), .ZN(n9686) );
  AOI22_X1 U10874 ( .A1(n4334), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9683), .B2(
        n9951), .ZN(n9684) );
  OAI21_X1 U10875 ( .B1(n9781), .B2(n9716), .A(n9684), .ZN(n9685) );
  AOI21_X1 U10876 ( .B1(n9686), .B2(n9960), .A(n9685), .ZN(n9687) );
  OAI211_X1 U10877 ( .C1(n9784), .C2(n4334), .A(n9688), .B(n9687), .ZN(
        P1_U3273) );
  XOR2_X1 U10878 ( .A(n9689), .B(n9695), .Z(n9790) );
  AOI211_X1 U10879 ( .C1(n9787), .C2(n9709), .A(n9977), .B(n9690), .ZN(n9786)
         );
  INV_X1 U10880 ( .A(n9787), .ZN(n9694) );
  INV_X1 U10881 ( .A(n9691), .ZN(n9692) );
  AOI22_X1 U10882 ( .A1(n4334), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9692), .B2(
        n9951), .ZN(n9693) );
  OAI21_X1 U10883 ( .B1(n9694), .B2(n9716), .A(n9693), .ZN(n9701) );
  XNOR2_X1 U10884 ( .A(n9696), .B(n9695), .ZN(n9699) );
  AOI21_X1 U10885 ( .B1(n9699), .B2(n9698), .A(n9697), .ZN(n9789) );
  NOR2_X1 U10886 ( .A1(n9789), .A2(n4334), .ZN(n9700) );
  AOI211_X1 U10887 ( .C1(n9786), .C2(n9960), .A(n9701), .B(n9700), .ZN(n9702)
         );
  OAI21_X1 U10888 ( .B1(n9720), .B2(n9790), .A(n9702), .ZN(P1_U3274) );
  XNOR2_X1 U10889 ( .A(n9704), .B(n9703), .ZN(n9795) );
  XNOR2_X1 U10890 ( .A(n9706), .B(n9705), .ZN(n9708) );
  OAI21_X1 U10891 ( .B1(n9708), .B2(n9945), .A(n9707), .ZN(n9791) );
  INV_X1 U10892 ( .A(n9793), .ZN(n9717) );
  INV_X1 U10893 ( .A(n9709), .ZN(n9710) );
  AOI211_X1 U10894 ( .C1(n9793), .C2(n9711), .A(n9977), .B(n9710), .ZN(n9792)
         );
  NAND2_X1 U10895 ( .A1(n9792), .A2(n9960), .ZN(n9715) );
  INV_X1 U10896 ( .A(n9712), .ZN(n9713) );
  AOI22_X1 U10897 ( .A1(n4334), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9713), .B2(
        n9951), .ZN(n9714) );
  OAI211_X1 U10898 ( .C1(n9717), .C2(n9716), .A(n9715), .B(n9714), .ZN(n9718)
         );
  AOI21_X1 U10899 ( .B1(n9723), .B2(n9791), .A(n9718), .ZN(n9719) );
  OAI21_X1 U10900 ( .B1(n9720), .B2(n9795), .A(n9719), .ZN(P1_U3275) );
  NAND2_X1 U10901 ( .A1(n9722), .A2(n9721), .ZN(n9734) );
  NAND2_X1 U10902 ( .A1(n9724), .A2(n9723), .ZN(n9733) );
  NAND2_X1 U10903 ( .A1(n4334), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n9725) );
  OAI21_X1 U10904 ( .B1(n9727), .B2(n9726), .A(n9725), .ZN(n9728) );
  AOI21_X1 U10905 ( .B1(n9729), .B2(n9953), .A(n9728), .ZN(n9732) );
  NAND2_X1 U10906 ( .A1(n9730), .A2(n9960), .ZN(n9731) );
  NAND4_X1 U10907 ( .A1(n9734), .A2(n9733), .A3(n9732), .A4(n9731), .ZN(
        P1_U3280) );
  INV_X1 U10908 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9737) );
  NOR2_X1 U10909 ( .A1(n9736), .A2(n9735), .ZN(n9803) );
  MUX2_X1 U10910 ( .A(n9737), .B(n9803), .S(n10068), .Z(n9738) );
  OAI21_X1 U10911 ( .B1(n9806), .B2(n9801), .A(n9738), .ZN(P1_U3553) );
  MUX2_X1 U10912 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n9739), .S(n10068), .Z(
        n9740) );
  AOI21_X1 U10913 ( .B1(n9777), .B2(n9741), .A(n9740), .ZN(n9742) );
  INV_X1 U10914 ( .A(n9742), .ZN(P1_U3552) );
  INV_X1 U10915 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n9746) );
  AOI211_X1 U10916 ( .C1(n9745), .C2(n10029), .A(n9744), .B(n9743), .ZN(n9807)
         );
  MUX2_X1 U10917 ( .A(n9746), .B(n9807), .S(n10068), .Z(n9747) );
  OAI21_X1 U10918 ( .B1(n4493), .B2(n9801), .A(n9747), .ZN(P1_U3549) );
  OAI211_X1 U10919 ( .C1(n9750), .C2(n9995), .A(n9749), .B(n9748), .ZN(n9810)
         );
  MUX2_X1 U10920 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9810), .S(n10068), .Z(
        n9751) );
  AOI21_X1 U10921 ( .B1(n9777), .B2(n9812), .A(n9751), .ZN(n9752) );
  INV_X1 U10922 ( .A(n9752), .ZN(P1_U3548) );
  INV_X1 U10923 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n9756) );
  AOI211_X1 U10924 ( .C1(n9755), .C2(n10029), .A(n9754), .B(n9753), .ZN(n9814)
         );
  MUX2_X1 U10925 ( .A(n9756), .B(n9814), .S(n10068), .Z(n9757) );
  OAI21_X1 U10926 ( .B1(n9817), .B2(n9801), .A(n9757), .ZN(P1_U3547) );
  INV_X1 U10927 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n9761) );
  AOI211_X1 U10928 ( .C1(n9760), .C2(n10029), .A(n9759), .B(n9758), .ZN(n9818)
         );
  MUX2_X1 U10929 ( .A(n9761), .B(n9818), .S(n10068), .Z(n9762) );
  OAI21_X1 U10930 ( .B1(n9821), .B2(n9801), .A(n9762), .ZN(P1_U3546) );
  OAI211_X1 U10931 ( .C1(n9765), .C2(n9995), .A(n9764), .B(n9763), .ZN(n9822)
         );
  MUX2_X1 U10932 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9822), .S(n10068), .Z(
        n9766) );
  AOI21_X1 U10933 ( .B1(n9777), .B2(n9824), .A(n9766), .ZN(n9767) );
  INV_X1 U10934 ( .A(n9767), .ZN(P1_U3545) );
  INV_X1 U10935 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n9771) );
  AOI211_X1 U10936 ( .C1(n9770), .C2(n10029), .A(n9769), .B(n9768), .ZN(n9826)
         );
  MUX2_X1 U10937 ( .A(n9771), .B(n9826), .S(n10068), .Z(n9772) );
  OAI21_X1 U10938 ( .B1(n4482), .B2(n9801), .A(n9772), .ZN(P1_U3544) );
  OAI211_X1 U10939 ( .C1(n9775), .C2(n9995), .A(n9774), .B(n9773), .ZN(n9829)
         );
  MUX2_X1 U10940 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9829), .S(n10068), .Z(
        n9776) );
  AOI21_X1 U10941 ( .B1(n9777), .B2(n9831), .A(n9776), .ZN(n9778) );
  INV_X1 U10942 ( .A(n9778), .ZN(P1_U3543) );
  NAND3_X1 U10943 ( .A1(n9780), .A2(n10029), .A3(n9779), .ZN(n9785) );
  NAND2_X1 U10944 ( .A1(n4484), .A2(n9993), .ZN(n9782) );
  NAND4_X1 U10945 ( .A1(n9785), .A2(n9784), .A3(n9783), .A4(n9782), .ZN(n9834)
         );
  MUX2_X1 U10946 ( .A(n9834), .B(P1_REG1_REG_20__SCAN_IN), .S(n10066), .Z(
        P1_U3542) );
  AOI21_X1 U10947 ( .B1(n9993), .B2(n9787), .A(n9786), .ZN(n9788) );
  OAI211_X1 U10948 ( .C1(n9790), .C2(n9995), .A(n9789), .B(n9788), .ZN(n9835)
         );
  MUX2_X1 U10949 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9835), .S(n10068), .Z(
        P1_U3541) );
  AOI211_X1 U10950 ( .C1(n9993), .C2(n9793), .A(n9792), .B(n9791), .ZN(n9794)
         );
  OAI21_X1 U10951 ( .B1(n9995), .B2(n9795), .A(n9794), .ZN(n9836) );
  MUX2_X1 U10952 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9836), .S(n10068), .Z(
        P1_U3540) );
  AOI211_X1 U10953 ( .C1(n9798), .C2(n10029), .A(n9797), .B(n9796), .ZN(n9837)
         );
  MUX2_X1 U10954 ( .A(n9799), .B(n9837), .S(n10068), .Z(n9800) );
  OAI21_X1 U10955 ( .B1(n4485), .B2(n9801), .A(n9800), .ZN(P1_U3539) );
  MUX2_X1 U10956 ( .A(P1_REG1_REG_0__SCAN_IN), .B(n9802), .S(n10068), .Z(
        P1_U3522) );
  MUX2_X1 U10957 ( .A(n9804), .B(n9803), .S(n10049), .Z(n9805) );
  OAI21_X1 U10958 ( .B1(n9806), .B2(n9840), .A(n9805), .ZN(P1_U3521) );
  INV_X1 U10959 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n9808) );
  MUX2_X1 U10960 ( .A(n9808), .B(n9807), .S(n10049), .Z(n9809) );
  OAI21_X1 U10961 ( .B1(n4493), .B2(n9840), .A(n9809), .ZN(P1_U3517) );
  MUX2_X1 U10962 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9810), .S(n10049), .Z(
        n9811) );
  AOI21_X1 U10963 ( .B1(n9832), .B2(n9812), .A(n9811), .ZN(n9813) );
  INV_X1 U10964 ( .A(n9813), .ZN(P1_U3516) );
  INV_X1 U10965 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n9815) );
  MUX2_X1 U10966 ( .A(n9815), .B(n9814), .S(n10049), .Z(n9816) );
  OAI21_X1 U10967 ( .B1(n9817), .B2(n9840), .A(n9816), .ZN(P1_U3515) );
  INV_X1 U10968 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n9819) );
  MUX2_X1 U10969 ( .A(n9819), .B(n9818), .S(n10049), .Z(n9820) );
  OAI21_X1 U10970 ( .B1(n9821), .B2(n9840), .A(n9820), .ZN(P1_U3514) );
  MUX2_X1 U10971 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9822), .S(n10049), .Z(
        n9823) );
  AOI21_X1 U10972 ( .B1(n9832), .B2(n9824), .A(n9823), .ZN(n9825) );
  INV_X1 U10973 ( .A(n9825), .ZN(P1_U3513) );
  INV_X1 U10974 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n9827) );
  MUX2_X1 U10975 ( .A(n9827), .B(n9826), .S(n10049), .Z(n9828) );
  OAI21_X1 U10976 ( .B1(n4482), .B2(n9840), .A(n9828), .ZN(P1_U3512) );
  MUX2_X1 U10977 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9829), .S(n10049), .Z(
        n9830) );
  AOI21_X1 U10978 ( .B1(n9832), .B2(n9831), .A(n9830), .ZN(n9833) );
  INV_X1 U10979 ( .A(n9833), .ZN(P1_U3511) );
  MUX2_X1 U10980 ( .A(n9834), .B(P1_REG0_REG_20__SCAN_IN), .S(n10047), .Z(
        P1_U3510) );
  MUX2_X1 U10981 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9835), .S(n10049), .Z(
        P1_U3509) );
  MUX2_X1 U10982 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9836), .S(n10049), .Z(
        P1_U3507) );
  INV_X1 U10983 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n9838) );
  MUX2_X1 U10984 ( .A(n9838), .B(n9837), .S(n10049), .Z(n9839) );
  OAI21_X1 U10985 ( .B1(n4485), .B2(n9840), .A(n9839), .ZN(P1_U3504) );
  MUX2_X1 U10986 ( .A(n9841), .B(P1_D_REG_1__SCAN_IN), .S(n9966), .Z(P1_U3440)
         );
  MUX2_X1 U10987 ( .A(n9842), .B(P1_D_REG_0__SCAN_IN), .S(n9966), .Z(P1_U3439)
         );
  NOR4_X1 U10988 ( .A1(n9843), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3086), .A4(
        n9844), .ZN(n9845) );
  AOI21_X1 U10989 ( .B1(n6448), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9845), .ZN(
        n9846) );
  OAI21_X1 U10990 ( .B1(n9847), .B2(n7965), .A(n9846), .ZN(P1_U3324) );
  AOI22_X1 U10991 ( .A1(n9848), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n6448), .ZN(n9849) );
  OAI21_X1 U10992 ( .B1(n9850), .B2(n7965), .A(n9849), .ZN(P1_U3325) );
  AOI22_X1 U10993 ( .A1(n9851), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n6448), .ZN(n9852) );
  OAI21_X1 U10994 ( .B1(n9853), .B2(n7965), .A(n9852), .ZN(P1_U3326) );
  MUX2_X1 U10995 ( .A(n9854), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  OAI21_X1 U10996 ( .B1(n9857), .B2(n9856), .A(n9855), .ZN(n9866) );
  INV_X1 U10997 ( .A(n9858), .ZN(n9859) );
  AOI21_X1 U10998 ( .B1(n9861), .B2(n9860), .A(n9859), .ZN(n9862) );
  OAI21_X1 U10999 ( .B1(n10026), .B2(n9863), .A(n9862), .ZN(n9864) );
  AOI21_X1 U11000 ( .B1(n9866), .B2(n9865), .A(n9864), .ZN(n9867) );
  OAI21_X1 U11001 ( .B1(n9869), .B2(n9868), .A(n9867), .ZN(P1_U3217) );
  NOR2_X1 U11002 ( .A1(n9870), .A2(n9995), .ZN(n9875) );
  OAI211_X1 U11003 ( .C1(n5589), .C2(n10039), .A(n9872), .B(n9871), .ZN(n9873)
         );
  AOI21_X1 U11004 ( .B1(n9875), .B2(n9874), .A(n9873), .ZN(n9877) );
  AOI22_X1 U11005 ( .A1(n10068), .A2(n9877), .B1(n9501), .B2(n10066), .ZN(
        P1_U3538) );
  INV_X1 U11006 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n9876) );
  AOI22_X1 U11007 ( .A1(n10049), .A2(n9877), .B1(n9876), .B2(n10047), .ZN(
        P1_U3501) );
  XNOR2_X1 U11008 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U11009 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  AOI21_X1 U11010 ( .B1(n9896), .B2(n7190), .A(n9878), .ZN(n9902) );
  OAI21_X1 U11011 ( .B1(P1_REG1_REG_0__SCAN_IN), .B2(n9896), .A(n9902), .ZN(
        n9879) );
  XOR2_X1 U11012 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9879), .Z(n9882) );
  AOI22_X1 U11013 ( .A1(n9933), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n9880) );
  OAI21_X1 U11014 ( .B1(n9882), .B2(n9881), .A(n9880), .ZN(P1_U3243) );
  AOI22_X1 U11015 ( .A1(n9933), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n9904) );
  OAI21_X1 U11016 ( .B1(n9886), .B2(n9885), .A(n9884), .ZN(n9894) );
  INV_X1 U11017 ( .A(n9887), .ZN(n9888) );
  OAI211_X1 U11018 ( .C1(n9890), .C2(n9889), .A(n9915), .B(n9888), .ZN(n9893)
         );
  NAND2_X1 U11019 ( .A1(n9937), .A2(n9891), .ZN(n9892) );
  OAI211_X1 U11020 ( .C1(n9919), .C2(n9894), .A(n9893), .B(n9892), .ZN(n9895)
         );
  INV_X1 U11021 ( .A(n9895), .ZN(n9903) );
  MUX2_X1 U11022 ( .A(n9898), .B(n9897), .S(n9896), .Z(n9900) );
  NAND2_X1 U11023 ( .A1(n9900), .A2(n9899), .ZN(n9901) );
  OAI211_X1 U11024 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n9902), .A(n9901), .B(
        P1_U3973), .ZN(n9922) );
  NAND3_X1 U11025 ( .A1(n9904), .A2(n9903), .A3(n9922), .ZN(P1_U3245) );
  NAND2_X1 U11026 ( .A1(n9906), .A2(n9905), .ZN(n9909) );
  INV_X1 U11027 ( .A(n9907), .ZN(n9908) );
  NAND2_X1 U11028 ( .A1(n9909), .A2(n9908), .ZN(n9918) );
  NAND2_X1 U11029 ( .A1(n9937), .A2(n9910), .ZN(n9917) );
  AOI21_X1 U11030 ( .B1(n9913), .B2(n9912), .A(n9911), .ZN(n9914) );
  NAND2_X1 U11031 ( .A1(n9915), .A2(n9914), .ZN(n9916) );
  OAI211_X1 U11032 ( .C1(n9919), .C2(n9918), .A(n9917), .B(n9916), .ZN(n9920)
         );
  INV_X1 U11033 ( .A(n9920), .ZN(n9924) );
  NAND2_X1 U11034 ( .A1(n9933), .A2(P1_ADDR_REG_4__SCAN_IN), .ZN(n9921) );
  NAND4_X1 U11035 ( .A1(n9924), .A2(n9923), .A3(n9922), .A4(n9921), .ZN(
        P1_U3247) );
  INV_X1 U11036 ( .A(n9925), .ZN(n9932) );
  INV_X1 U11037 ( .A(n9926), .ZN(n9927) );
  AOI211_X1 U11038 ( .C1(n9930), .C2(n9929), .A(n9928), .B(n9927), .ZN(n9931)
         );
  AOI211_X1 U11039 ( .C1(n9933), .C2(P1_ADDR_REG_16__SCAN_IN), .A(n9932), .B(
        n9931), .ZN(n9942) );
  OAI21_X1 U11040 ( .B1(n9936), .B2(n9935), .A(n9934), .ZN(n9940) );
  AOI22_X1 U11041 ( .A1(n9940), .A2(n9939), .B1(n9938), .B2(n9937), .ZN(n9941)
         );
  NAND2_X1 U11042 ( .A1(n9942), .A2(n9941), .ZN(P1_U3259) );
  XNOR2_X1 U11043 ( .A(n9943), .B(n9946), .ZN(n10009) );
  AOI211_X1 U11044 ( .C1(n9947), .C2(n9946), .A(n9945), .B(n9944), .ZN(n9948)
         );
  AOI211_X1 U11045 ( .C1(n10046), .C2(n10009), .A(n9949), .B(n9948), .ZN(
        n10006) );
  INV_X1 U11046 ( .A(n9950), .ZN(n9952) );
  AOI222_X1 U11047 ( .A1(n9954), .A2(n9953), .B1(n9952), .B2(n9951), .C1(
        P1_REG2_REG_7__SCAN_IN), .C2(n4334), .ZN(n9963) );
  INV_X1 U11048 ( .A(n9955), .ZN(n9958) );
  OAI211_X1 U11049 ( .C1(n9958), .C2(n4479), .A(n9957), .B(n9956), .ZN(n10005)
         );
  INV_X1 U11050 ( .A(n10005), .ZN(n9959) );
  AOI22_X1 U11051 ( .A1(n10009), .A2(n9961), .B1(n9960), .B2(n9959), .ZN(n9962) );
  OAI211_X1 U11052 ( .C1(n4334), .C2(n10006), .A(n9963), .B(n9962), .ZN(
        P1_U3286) );
  AND2_X1 U11053 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9966), .ZN(P1_U3294) );
  AND2_X1 U11054 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9966), .ZN(P1_U3295) );
  AND2_X1 U11055 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9966), .ZN(P1_U3296) );
  AND2_X1 U11056 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9966), .ZN(P1_U3297) );
  AND2_X1 U11057 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9966), .ZN(P1_U3298) );
  AND2_X1 U11058 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9966), .ZN(P1_U3299) );
  INV_X1 U11059 ( .A(n9966), .ZN(n9965) );
  NOR2_X1 U11060 ( .A1(n9965), .A2(n9964), .ZN(P1_U3300) );
  AND2_X1 U11061 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9966), .ZN(P1_U3301) );
  AND2_X1 U11062 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9966), .ZN(P1_U3302) );
  AND2_X1 U11063 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9966), .ZN(P1_U3303) );
  AND2_X1 U11064 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9966), .ZN(P1_U3304) );
  AND2_X1 U11065 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9966), .ZN(P1_U3305) );
  AND2_X1 U11066 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9966), .ZN(P1_U3306) );
  AND2_X1 U11067 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9966), .ZN(P1_U3307) );
  AND2_X1 U11068 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9966), .ZN(P1_U3308) );
  AND2_X1 U11069 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9966), .ZN(P1_U3309) );
  AND2_X1 U11070 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9966), .ZN(P1_U3310) );
  AND2_X1 U11071 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9966), .ZN(P1_U3311) );
  AND2_X1 U11072 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9966), .ZN(P1_U3312) );
  AND2_X1 U11073 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9966), .ZN(P1_U3313) );
  AND2_X1 U11074 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9966), .ZN(P1_U3314) );
  AND2_X1 U11075 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9966), .ZN(P1_U3315) );
  AND2_X1 U11076 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9966), .ZN(P1_U3316) );
  AND2_X1 U11077 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9966), .ZN(P1_U3317) );
  AND2_X1 U11078 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9966), .ZN(P1_U3318) );
  AND2_X1 U11079 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9966), .ZN(P1_U3319) );
  AND2_X1 U11080 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9966), .ZN(P1_U3320) );
  AND2_X1 U11081 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n9966), .ZN(P1_U3321) );
  AND2_X1 U11082 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9966), .ZN(P1_U3322) );
  AND2_X1 U11083 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9966), .ZN(P1_U3323) );
  INV_X1 U11084 ( .A(n9967), .ZN(n9973) );
  NOR2_X1 U11085 ( .A1(n9967), .A2(n10041), .ZN(n9972) );
  OAI211_X1 U11086 ( .C1(n9970), .C2(n10039), .A(n9969), .B(n9968), .ZN(n9971)
         );
  AOI211_X1 U11087 ( .C1(n10046), .C2(n9973), .A(n9972), .B(n9971), .ZN(n10051) );
  INV_X1 U11088 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9974) );
  AOI22_X1 U11089 ( .A1(n10049), .A2(n10051), .B1(n9974), .B2(n10047), .ZN(
        P1_U3456) );
  INV_X1 U11090 ( .A(n9975), .ZN(n9978) );
  OAI22_X1 U11091 ( .A1(n9978), .A2(n9977), .B1(n9976), .B2(n10039), .ZN(n9981) );
  INV_X1 U11092 ( .A(n9979), .ZN(n9980) );
  AOI211_X1 U11093 ( .C1(n9982), .C2(n10029), .A(n9981), .B(n9980), .ZN(n10053) );
  AOI22_X1 U11094 ( .A1(n10049), .A2(n10053), .B1(n4983), .B2(n10047), .ZN(
        P1_U3462) );
  INV_X1 U11095 ( .A(n9983), .ZN(n9984) );
  OAI21_X1 U11096 ( .B1(n9985), .B2(n10039), .A(n9984), .ZN(n9988) );
  INV_X1 U11097 ( .A(n9986), .ZN(n9987) );
  AOI211_X1 U11098 ( .C1(n10029), .C2(n9989), .A(n9988), .B(n9987), .ZN(n10054) );
  INV_X1 U11099 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n9990) );
  AOI22_X1 U11100 ( .A1(n10049), .A2(n10054), .B1(n9990), .B2(n10047), .ZN(
        P1_U3465) );
  AOI21_X1 U11101 ( .B1(n9993), .B2(n9992), .A(n9991), .ZN(n9994) );
  OAI21_X1 U11102 ( .B1(n9996), .B2(n9995), .A(n9994), .ZN(n9997) );
  NOR2_X1 U11103 ( .A1(n9998), .A2(n9997), .ZN(n10056) );
  AOI22_X1 U11104 ( .A1(n10049), .A2(n10056), .B1(n5025), .B2(n10047), .ZN(
        P1_U3468) );
  INV_X1 U11105 ( .A(n9999), .ZN(n10004) );
  OAI21_X1 U11106 ( .B1(n10001), .B2(n10039), .A(n10000), .ZN(n10003) );
  AOI211_X1 U11107 ( .C1(n10004), .C2(n10029), .A(n10003), .B(n10002), .ZN(
        n10058) );
  AOI22_X1 U11108 ( .A1(n10049), .A2(n10058), .B1(n5061), .B2(n10047), .ZN(
        P1_U3471) );
  OAI21_X1 U11109 ( .B1(n4479), .B2(n10039), .A(n10005), .ZN(n10008) );
  INV_X1 U11110 ( .A(n10006), .ZN(n10007) );
  AOI211_X1 U11111 ( .C1(n10033), .C2(n10009), .A(n10008), .B(n10007), .ZN(
        n10060) );
  AOI22_X1 U11112 ( .A1(n10049), .A2(n10060), .B1(n5079), .B2(n10047), .ZN(
        P1_U3474) );
  NOR2_X1 U11113 ( .A1(n10010), .A2(n10041), .ZN(n10015) );
  OAI211_X1 U11114 ( .C1(n10013), .C2(n10039), .A(n10012), .B(n10011), .ZN(
        n10014) );
  AOI211_X1 U11115 ( .C1(n10046), .C2(n10016), .A(n10015), .B(n10014), .ZN(
        n10061) );
  AOI22_X1 U11116 ( .A1(n10049), .A2(n10061), .B1(n5102), .B2(n10047), .ZN(
        P1_U3477) );
  INV_X1 U11117 ( .A(n10017), .ZN(n10019) );
  OAI21_X1 U11118 ( .B1(n10019), .B2(n10039), .A(n10018), .ZN(n10022) );
  INV_X1 U11119 ( .A(n10020), .ZN(n10021) );
  AOI211_X1 U11120 ( .C1(n10029), .C2(n10023), .A(n10022), .B(n10021), .ZN(
        n10063) );
  AOI22_X1 U11121 ( .A1(n10049), .A2(n10063), .B1(n5120), .B2(n10047), .ZN(
        P1_U3480) );
  OAI211_X1 U11122 ( .C1(n10026), .C2(n10039), .A(n10025), .B(n10024), .ZN(
        n10027) );
  AOI21_X1 U11123 ( .B1(n10029), .B2(n10028), .A(n10027), .ZN(n10064) );
  AOI22_X1 U11124 ( .A1(n10049), .A2(n10064), .B1(n5146), .B2(n10047), .ZN(
        P1_U3483) );
  OAI21_X1 U11125 ( .B1(n10031), .B2(n10039), .A(n10030), .ZN(n10032) );
  AOI21_X1 U11126 ( .B1(n10034), .B2(n10033), .A(n10032), .ZN(n10035) );
  AND2_X1 U11127 ( .A1(n10036), .A2(n10035), .ZN(n10065) );
  AOI22_X1 U11128 ( .A1(n10049), .A2(n10065), .B1(n5177), .B2(n10047), .ZN(
        P1_U3486) );
  OAI211_X1 U11129 ( .C1(n10040), .C2(n10039), .A(n10038), .B(n10037), .ZN(
        n10044) );
  NOR2_X1 U11130 ( .A1(n10042), .A2(n10041), .ZN(n10043) );
  AOI211_X1 U11131 ( .C1(n10046), .C2(n10045), .A(n10044), .B(n10043), .ZN(
        n10067) );
  INV_X1 U11132 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n10048) );
  AOI22_X1 U11133 ( .A1(n10049), .A2(n10067), .B1(n10048), .B2(n10047), .ZN(
        P1_U3495) );
  AOI22_X1 U11134 ( .A1(n10068), .A2(n10051), .B1(n10050), .B2(n10066), .ZN(
        P1_U3523) );
  INV_X1 U11135 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n10052) );
  AOI22_X1 U11136 ( .A1(n10068), .A2(n10053), .B1(n10052), .B2(n10066), .ZN(
        P1_U3525) );
  AOI22_X1 U11137 ( .A1(n10068), .A2(n10054), .B1(n5004), .B2(n10066), .ZN(
        P1_U3526) );
  INV_X1 U11138 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n10055) );
  AOI22_X1 U11139 ( .A1(n10068), .A2(n10056), .B1(n10055), .B2(n10066), .ZN(
        P1_U3527) );
  INV_X1 U11140 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n10057) );
  AOI22_X1 U11141 ( .A1(n10068), .A2(n10058), .B1(n10057), .B2(n10066), .ZN(
        P1_U3528) );
  INV_X1 U11142 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n10059) );
  AOI22_X1 U11143 ( .A1(n10068), .A2(n10060), .B1(n10059), .B2(n10066), .ZN(
        P1_U3529) );
  AOI22_X1 U11144 ( .A1(n10068), .A2(n10061), .B1(n4471), .B2(n10066), .ZN(
        P1_U3530) );
  INV_X1 U11145 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10062) );
  AOI22_X1 U11146 ( .A1(n10068), .A2(n10063), .B1(n10062), .B2(n10066), .ZN(
        P1_U3531) );
  AOI22_X1 U11147 ( .A1(n10068), .A2(n10064), .B1(n7023), .B2(n10066), .ZN(
        P1_U3532) );
  AOI22_X1 U11148 ( .A1(n10068), .A2(n10065), .B1(n7267), .B2(n10066), .ZN(
        P1_U3533) );
  AOI22_X1 U11149 ( .A1(n10068), .A2(n10067), .B1(n7679), .B2(n10066), .ZN(
        P1_U3536) );
  INV_X1 U11150 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n10070) );
  AOI22_X1 U11151 ( .A1(n10135), .A2(n10070), .B1(n10069), .B2(n10133), .ZN(
        P2_U3390) );
  INV_X1 U11152 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10075) );
  OAI21_X1 U11153 ( .B1(n10072), .B2(n10114), .A(n10071), .ZN(n10073) );
  AOI21_X1 U11154 ( .B1(n10074), .B2(n10091), .A(n10073), .ZN(n10137) );
  AOI22_X1 U11155 ( .A1(n10135), .A2(n10075), .B1(n10137), .B2(n10133), .ZN(
        P2_U3399) );
  INV_X1 U11156 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10081) );
  AND2_X1 U11157 ( .A1(n10076), .A2(n10132), .ZN(n10077) );
  AOI21_X1 U11158 ( .B1(n10078), .B2(n10091), .A(n10077), .ZN(n10080) );
  AND2_X1 U11159 ( .A1(n10080), .A2(n10079), .ZN(n10139) );
  AOI22_X1 U11160 ( .A1(n10135), .A2(n10081), .B1(n10139), .B2(n10133), .ZN(
        P2_U3402) );
  INV_X1 U11161 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10087) );
  INV_X1 U11162 ( .A(n10082), .ZN(n10084) );
  OAI22_X1 U11163 ( .A1(n10084), .A2(n10116), .B1(n10083), .B2(n10114), .ZN(
        n10085) );
  NOR2_X1 U11164 ( .A1(n10086), .A2(n10085), .ZN(n10141) );
  AOI22_X1 U11165 ( .A1(n10135), .A2(n10087), .B1(n10141), .B2(n10133), .ZN(
        P2_U3405) );
  INV_X1 U11166 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10093) );
  OAI21_X1 U11167 ( .B1(n10089), .B2(n10114), .A(n10088), .ZN(n10090) );
  AOI21_X1 U11168 ( .B1(n10092), .B2(n10091), .A(n10090), .ZN(n10142) );
  AOI22_X1 U11169 ( .A1(n10135), .A2(n10093), .B1(n10142), .B2(n10133), .ZN(
        P2_U3408) );
  INV_X1 U11170 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10101) );
  OR2_X1 U11171 ( .A1(n10097), .A2(n10107), .ZN(n10096) );
  NAND2_X1 U11172 ( .A1(n10094), .A2(n10132), .ZN(n10095) );
  OAI211_X1 U11173 ( .C1(n10097), .C2(n10116), .A(n10096), .B(n10095), .ZN(
        n10098) );
  INV_X1 U11174 ( .A(n10098), .ZN(n10100) );
  AND2_X1 U11175 ( .A1(n10100), .A2(n10099), .ZN(n10144) );
  AOI22_X1 U11176 ( .A1(n10135), .A2(n10101), .B1(n10144), .B2(n10133), .ZN(
        P2_U3411) );
  INV_X1 U11177 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10106) );
  OAI22_X1 U11178 ( .A1(n10103), .A2(n10126), .B1(n10102), .B2(n10114), .ZN(
        n10104) );
  NOR2_X1 U11179 ( .A1(n10105), .A2(n10104), .ZN(n10145) );
  AOI22_X1 U11180 ( .A1(n10135), .A2(n10106), .B1(n10145), .B2(n10133), .ZN(
        P2_U3414) );
  INV_X1 U11181 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10113) );
  NOR2_X1 U11182 ( .A1(n10109), .A2(n10107), .ZN(n10111) );
  OAI22_X1 U11183 ( .A1(n10109), .A2(n10116), .B1(n10108), .B2(n10114), .ZN(
        n10110) );
  NOR3_X1 U11184 ( .A1(n10112), .A2(n10111), .A3(n10110), .ZN(n10146) );
  AOI22_X1 U11185 ( .A1(n10135), .A2(n10113), .B1(n10146), .B2(n10133), .ZN(
        P2_U3417) );
  OAI22_X1 U11186 ( .A1(n10117), .A2(n10116), .B1(n10115), .B2(n10114), .ZN(
        n10118) );
  NOR2_X1 U11187 ( .A1(n10119), .A2(n10118), .ZN(n10147) );
  AOI22_X1 U11188 ( .A1(n10135), .A2(n10120), .B1(n10147), .B2(n10133), .ZN(
        P2_U3420) );
  INV_X1 U11189 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10125) );
  NOR2_X1 U11190 ( .A1(n10121), .A2(n10126), .ZN(n10123) );
  AOI211_X1 U11191 ( .C1(n10132), .C2(n10124), .A(n10123), .B(n10122), .ZN(
        n10149) );
  AOI22_X1 U11192 ( .A1(n10135), .A2(n10125), .B1(n10149), .B2(n10133), .ZN(
        P2_U3423) );
  NOR3_X1 U11193 ( .A1(n10128), .A2(n10127), .A3(n10126), .ZN(n10130) );
  AOI211_X1 U11194 ( .C1(n10132), .C2(n10131), .A(n10130), .B(n10129), .ZN(
        n10151) );
  AOI22_X1 U11195 ( .A1(n10135), .A2(n10134), .B1(n10151), .B2(n10133), .ZN(
        P2_U3426) );
  AOI22_X1 U11196 ( .A1(n10152), .A2(n10137), .B1(n10136), .B2(n10150), .ZN(
        P2_U3462) );
  AOI22_X1 U11197 ( .A1(n10152), .A2(n10139), .B1(n10138), .B2(n10150), .ZN(
        P2_U3463) );
  AOI22_X1 U11198 ( .A1(n10152), .A2(n10141), .B1(n10140), .B2(n10150), .ZN(
        P2_U3464) );
  AOI22_X1 U11199 ( .A1(n10152), .A2(n10142), .B1(n6821), .B2(n10150), .ZN(
        P2_U3465) );
  AOI22_X1 U11200 ( .A1(n10152), .A2(n10144), .B1(n10143), .B2(n10150), .ZN(
        P2_U3466) );
  AOI22_X1 U11201 ( .A1(n10152), .A2(n10145), .B1(n7001), .B2(n10150), .ZN(
        P2_U3467) );
  AOI22_X1 U11202 ( .A1(n10152), .A2(n10146), .B1(n6992), .B2(n10150), .ZN(
        P2_U3468) );
  AOI22_X1 U11203 ( .A1(n10152), .A2(n10147), .B1(n7066), .B2(n10150), .ZN(
        P2_U3469) );
  AOI22_X1 U11204 ( .A1(n10152), .A2(n10149), .B1(n10148), .B2(n10150), .ZN(
        P2_U3470) );
  AOI22_X1 U11205 ( .A1(n10152), .A2(n10151), .B1(n7505), .B2(n10150), .ZN(
        P2_U3471) );
  OAI222_X1 U11206 ( .A1(n10157), .A2(n10156), .B1(n10157), .B2(n10155), .C1(
        n10154), .C2(n10153), .ZN(ADD_1068_U5) );
  XOR2_X1 U11207 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  OAI21_X1 U11208 ( .B1(n10160), .B2(n10159), .A(n10158), .ZN(n10161) );
  XNOR2_X1 U11209 ( .A(n10161), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(ADD_1068_U55)
         );
  OAI21_X1 U11210 ( .B1(n10164), .B2(n10163), .A(n10162), .ZN(ADD_1068_U56) );
  OAI21_X1 U11211 ( .B1(n10167), .B2(n10166), .A(n10165), .ZN(ADD_1068_U57) );
  OAI21_X1 U11212 ( .B1(n10170), .B2(n10169), .A(n10168), .ZN(ADD_1068_U58) );
  OAI21_X1 U11213 ( .B1(n10173), .B2(n10172), .A(n10171), .ZN(ADD_1068_U59) );
  OAI21_X1 U11214 ( .B1(n10176), .B2(n10175), .A(n10174), .ZN(ADD_1068_U60) );
  OAI21_X1 U11215 ( .B1(n10179), .B2(n10178), .A(n10177), .ZN(ADD_1068_U61) );
  OAI21_X1 U11216 ( .B1(n10182), .B2(n10181), .A(n10180), .ZN(ADD_1068_U62) );
  OAI21_X1 U11217 ( .B1(n10185), .B2(n10184), .A(n10183), .ZN(ADD_1068_U63) );
  OAI21_X1 U11218 ( .B1(n10188), .B2(n10187), .A(n10186), .ZN(ADD_1068_U51) );
  OAI21_X1 U11219 ( .B1(n10191), .B2(n10190), .A(n10189), .ZN(ADD_1068_U50) );
  OAI21_X1 U11220 ( .B1(n10194), .B2(n10193), .A(n10192), .ZN(ADD_1068_U47) );
  OAI21_X1 U11221 ( .B1(n10197), .B2(n10196), .A(n10195), .ZN(ADD_1068_U49) );
  OAI21_X1 U11222 ( .B1(n10200), .B2(n10199), .A(n10198), .ZN(ADD_1068_U48) );
  AOI21_X1 U11223 ( .B1(n10203), .B2(n10202), .A(n10201), .ZN(ADD_1068_U54) );
  AOI21_X1 U11224 ( .B1(n10206), .B2(n10205), .A(n10204), .ZN(ADD_1068_U53) );
  OAI21_X1 U11225 ( .B1(n10209), .B2(n10208), .A(n10207), .ZN(ADD_1068_U52) );
  INV_X1 U4845 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9844) );
  CLKBUF_X1 U4850 ( .A(n8430), .Z(n8567) );
  CLKBUF_X1 U4855 ( .A(n4979), .Z(n6530) );
endmodule

