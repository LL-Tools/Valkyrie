

module b21_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, P2_WR_REG_SCAN_IN, SI_31_, 
        SI_30_, SI_29_, SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, 
        SI_21_, SI_20_, SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, 
        SI_12_, SI_11_, SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, 
        SI_3_, SI_2_, SI_1_, SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, 
        ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, 
        ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, 
        ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, 
        ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, P1_U3352, P1_U3351, 
        P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, 
        P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, 
        P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, 
        P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, 
        P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, 
        P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, 
        P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, 
        P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, 
        P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, 
        P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, 
        P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, 
        P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, 
        P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, 
        P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, 
        P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, 
        P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, 
        P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, 
        P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, 
        P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, 
        P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, 
        P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, 
        P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, 
        P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, 
        P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, 
        P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, 
        P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, 
        P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, 
        P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, 
        P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, 
        P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, 
        P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, 
        P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, 
        P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, 
        P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, 
        P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, 
        P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, 
        P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, 
        P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, 
        P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, 
        P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, 
        P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, 
        P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, 
        P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, 
        P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, 
        P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, 
        P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, 
        P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, 
        P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3152, P2_U3151, P2_U3966 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_,
         SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_,
         SI_20_, SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_,
         SI_12_, SI_11_, SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_,
         SI_3_, SI_2_, SI_1_, SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_REG3_REG_7__SCAN_IN, P2_REG3_REG_27__SCAN_IN,
         P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_23__SCAN_IN,
         P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_3__SCAN_IN,
         P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_28__SCAN_IN,
         P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_1__SCAN_IN,
         P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_12__SCAN_IN,
         P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_16__SCAN_IN,
         P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_17__SCAN_IN,
         P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_4__SCAN_IN,
         P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN,
         P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN,
         P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN,
         P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN,
         P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN,
         P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855,
         n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865,
         n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875,
         n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885,
         n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895,
         n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905,
         n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915,
         n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925,
         n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935,
         n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945,
         n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955,
         n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965,
         n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975,
         n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985,
         n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995,
         n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005,
         n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015,
         n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025,
         n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035,
         n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045,
         n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055,
         n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065,
         n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075,
         n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085,
         n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095,
         n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105,
         n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115,
         n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125,
         n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135,
         n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145,
         n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155,
         n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165,
         n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175,
         n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185,
         n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195,
         n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205,
         n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215,
         n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225,
         n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235,
         n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245,
         n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255,
         n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265,
         n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275,
         n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285,
         n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295,
         n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305,
         n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315,
         n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325,
         n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335,
         n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345,
         n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355,
         n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365,
         n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375,
         n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385,
         n5386, n5387, n5388, n5389, n5390, n5392, n5393, n5394, n5395, n5396,
         n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406,
         n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416,
         n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426,
         n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436,
         n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446,
         n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456,
         n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466,
         n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476,
         n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486,
         n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496,
         n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506,
         n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516,
         n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526,
         n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536,
         n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546,
         n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556,
         n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566,
         n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576,
         n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586,
         n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596,
         n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606,
         n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616,
         n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626,
         n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636,
         n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646,
         n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656,
         n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666,
         n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676,
         n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686,
         n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696,
         n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706,
         n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716,
         n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726,
         n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736,
         n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746,
         n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756,
         n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766,
         n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776,
         n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786,
         n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796,
         n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806,
         n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816,
         n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826,
         n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836,
         n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846,
         n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856,
         n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866,
         n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876,
         n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886,
         n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896,
         n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906,
         n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916,
         n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926,
         n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936,
         n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946,
         n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956,
         n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966,
         n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976,
         n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986,
         n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996,
         n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006,
         n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016,
         n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026,
         n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036,
         n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046,
         n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056,
         n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066,
         n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076,
         n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086,
         n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096,
         n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106,
         n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116,
         n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126,
         n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136,
         n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146,
         n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156,
         n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166,
         n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176,
         n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186,
         n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196,
         n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206,
         n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216,
         n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226,
         n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236,
         n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246,
         n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256,
         n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266,
         n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276,
         n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286,
         n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296,
         n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306,
         n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316,
         n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326,
         n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336,
         n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346,
         n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356,
         n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366,
         n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376,
         n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386,
         n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396,
         n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406,
         n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416,
         n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426,
         n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436,
         n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446,
         n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456,
         n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466,
         n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476,
         n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486,
         n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496,
         n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506,
         n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516,
         n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526,
         n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536,
         n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546,
         n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556,
         n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566,
         n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576,
         n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586,
         n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596,
         n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606,
         n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616,
         n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626,
         n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636,
         n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646,
         n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656,
         n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666,
         n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676,
         n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686,
         n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696,
         n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706,
         n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716,
         n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726,
         n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736,
         n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746,
         n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756,
         n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766,
         n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776,
         n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786,
         n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796,
         n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806,
         n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816,
         n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826,
         n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836,
         n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846,
         n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856,
         n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866,
         n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876,
         n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886,
         n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896,
         n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906,
         n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916,
         n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926,
         n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936,
         n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946,
         n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956,
         n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966,
         n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976,
         n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986,
         n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996,
         n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006,
         n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016,
         n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026,
         n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036,
         n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046,
         n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056,
         n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066,
         n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076,
         n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086,
         n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096,
         n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106,
         n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116,
         n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126,
         n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136,
         n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146,
         n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156,
         n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166,
         n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176,
         n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186,
         n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196,
         n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206,
         n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216,
         n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226,
         n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236,
         n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246,
         n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256,
         n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266,
         n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276,
         n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286,
         n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296,
         n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306,
         n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316,
         n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326,
         n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336,
         n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346,
         n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356,
         n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366,
         n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376,
         n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386,
         n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396,
         n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406,
         n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416,
         n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426,
         n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436,
         n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446,
         n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456,
         n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466,
         n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476,
         n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486,
         n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496,
         n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506,
         n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516,
         n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526,
         n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536,
         n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546,
         n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556,
         n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566,
         n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576,
         n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586,
         n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596,
         n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606,
         n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616,
         n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626,
         n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636,
         n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646,
         n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656,
         n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666,
         n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676,
         n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686,
         n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696,
         n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706,
         n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716,
         n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726,
         n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736,
         n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746,
         n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756,
         n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766,
         n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776,
         n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786,
         n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796,
         n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806,
         n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816,
         n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826,
         n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836,
         n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846,
         n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856,
         n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866,
         n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876,
         n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886,
         n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896,
         n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906,
         n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916,
         n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926,
         n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936,
         n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946,
         n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956,
         n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966,
         n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976,
         n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986,
         n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996,
         n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006,
         n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016,
         n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026,
         n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036,
         n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046,
         n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056,
         n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066,
         n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076,
         n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086,
         n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096,
         n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106,
         n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116,
         n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126,
         n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136,
         n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146,
         n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156,
         n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166,
         n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176,
         n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186,
         n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196,
         n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206,
         n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216,
         n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226,
         n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236,
         n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246,
         n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256,
         n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266,
         n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276,
         n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286,
         n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296,
         n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306,
         n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316,
         n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326,
         n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336,
         n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346,
         n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356,
         n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366,
         n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376,
         n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386,
         n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396,
         n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406,
         n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416,
         n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426,
         n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436,
         n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446,
         n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456,
         n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466,
         n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476,
         n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486,
         n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496,
         n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506,
         n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516,
         n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526,
         n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536,
         n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546,
         n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556,
         n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566,
         n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576,
         n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586,
         n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596,
         n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606,
         n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616,
         n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626,
         n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636,
         n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646,
         n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656,
         n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666,
         n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676,
         n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686,
         n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696,
         n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706,
         n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716,
         n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726,
         n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736,
         n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746,
         n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756,
         n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766,
         n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776,
         n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786,
         n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796,
         n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806,
         n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816,
         n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826,
         n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836,
         n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846,
         n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856,
         n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866,
         n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876,
         n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886,
         n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896,
         n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906,
         n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916,
         n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926,
         n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936,
         n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946,
         n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956,
         n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966,
         n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976,
         n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986,
         n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996,
         n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006,
         n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016,
         n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026,
         n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036,
         n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046,
         n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056,
         n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066,
         n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076,
         n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086,
         n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096,
         n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106,
         n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116,
         n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126,
         n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136,
         n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146,
         n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156,
         n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166,
         n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176,
         n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186,
         n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196,
         n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206,
         n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216,
         n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226,
         n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236,
         n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246,
         n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256,
         n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266,
         n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276,
         n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286,
         n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296,
         n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306,
         n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316,
         n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326,
         n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336,
         n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346,
         n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356,
         n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366,
         n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376,
         n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386,
         n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396,
         n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406,
         n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416,
         n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426,
         n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436,
         n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446,
         n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456,
         n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466,
         n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476,
         n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486,
         n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496,
         n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506,
         n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516,
         n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526,
         n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536,
         n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546,
         n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556,
         n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566,
         n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576,
         n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586,
         n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596,
         n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606,
         n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616,
         n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626,
         n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636,
         n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646,
         n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656,
         n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666,
         n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676,
         n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686,
         n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696,
         n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706,
         n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716,
         n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726,
         n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736,
         n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746,
         n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756,
         n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766,
         n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776,
         n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786,
         n9787, n9788, n9789, n9790, n9791, n9794, n9795, n9796, n9797, n9798,
         n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808,
         n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818,
         n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828,
         n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838,
         n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848,
         n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858,
         n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868,
         n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878,
         n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888,
         n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898,
         n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908,
         n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918,
         n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928,
         n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938,
         n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948,
         n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958,
         n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968,
         n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978,
         n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988,
         n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998,
         n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
         n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
         n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
         n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
         n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
         n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,
         n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
         n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
         n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656,
         n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664,
         n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672,
         n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680,
         n10681, n10682, n10683, n10684;

  INV_X1 U4909 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  AND2_X1 U4910 ( .A1(n7667), .A2(n7375), .ZN(n8711) );
  AND2_X1 U4911 ( .A1(n7989), .A2(n7096), .ZN(n7098) );
  INV_X2 U4912 ( .A(n8702), .ZN(n8718) );
  XNOR2_X1 U4913 ( .A(n7491), .B(n7766), .ZN(n6077) );
  NAND4_X2 U4914 ( .A1(n5719), .A2(n5718), .A3(n5717), .A4(n5716), .ZN(n7491)
         );
  NAND2_X1 U4915 ( .A1(n7377), .A2(n7663), .ZN(n8701) );
  INV_X1 U4916 ( .A(n10491), .ZN(n9791) );
  NAND2_X1 U4917 ( .A1(n9385), .A2(n6841), .ZN(n7172) );
  NAND2_X1 U4918 ( .A1(n5551), .A2(n5550), .ZN(n10260) );
  INV_X1 U4921 ( .A(P2_STATE_REG_SCAN_IN), .ZN(n4846) );
  CLKBUF_X3 U4923 ( .A(n6259), .Z(n4852) );
  AND2_X1 U4924 ( .A1(n7948), .A2(n6676), .ZN(n8138) );
  INV_X4 U4925 ( .A(n6960), .ZN(n6976) );
  INV_X1 U4926 ( .A(n6498), .ZN(n6482) );
  OR2_X1 U4927 ( .A1(n6841), .A2(n7180), .ZN(n10611) );
  INV_X1 U4928 ( .A(n8720), .ZN(n8713) );
  INV_X1 U4929 ( .A(n8711), .ZN(n7496) );
  AND2_X1 U4930 ( .A1(n7597), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n7595) );
  INV_X1 U4931 ( .A(n7914), .ZN(n10518) );
  INV_X1 U4932 ( .A(n7929), .ZN(n10502) );
  INV_X1 U4934 ( .A(n6228), .ZN(n9379) );
  OAI22_X1 U4935 ( .A1(n7595), .A2(n7711), .B1(P1_REG2_REG_11__SCAN_IN), .B2(
        n7597), .ZN(n7718) );
  INV_X2 U4936 ( .A(n5774), .ZN(n6041) );
  AOI211_X1 U4937 ( .C1(n10071), .C2(n10026), .A(n8822), .B(n8821), .ZN(n8823)
         );
  AND4_X1 U4938 ( .A1(n6431), .A2(n6415), .A3(n6401), .A4(n6386), .ZN(n4847)
         );
  OAI211_X1 U4939 ( .C1(n5745), .C2(n7307), .A(n5795), .B(n5794), .ZN(n7997)
         );
  NOR2_X2 U4940 ( .A1(n8513), .A2(n6430), .ZN(n8512) );
  INV_X1 U4941 ( .A(n7753), .ZN(n7633) );
  OAI21_X2 U4942 ( .B1(n8279), .B2(n8284), .A(n6697), .ZN(n8367) );
  INV_X1 U4943 ( .A(n5774), .ZN(n4848) );
  NAND2_X1 U4944 ( .A1(n4853), .A2(n6238), .ZN(n5774) );
  XNOR2_X1 U4945 ( .A(n6626), .B(P2_IR_REG_19__SCAN_IN), .ZN(n6624) );
  NAND2_X1 U4946 ( .A1(n9135), .A2(n9056), .ZN(n9121) );
  NAND2_X1 U4947 ( .A1(n7051), .A2(n7050), .ZN(n9953) );
  AND2_X1 U4948 ( .A1(n4990), .A2(n4989), .ZN(n9163) );
  NOR2_X1 U4949 ( .A1(n5081), .A2(n9141), .ZN(n5080) );
  NAND2_X1 U4950 ( .A1(n6752), .A2(n6755), .ZN(n9162) );
  NAND2_X1 U4951 ( .A1(n10051), .A2(n10050), .ZN(n5175) );
  OAI21_X1 U4952 ( .B1(n8551), .B2(n7042), .A(n7041), .ZN(n10051) );
  NAND2_X1 U4953 ( .A1(n8524), .A2(n7039), .ZN(n8551) );
  NAND2_X1 U4954 ( .A1(n5917), .A2(n5916), .ZN(n10152) );
  AOI21_X1 U4955 ( .B1(n7255), .B2(n5250), .A(n5095), .ZN(n10595) );
  AND2_X1 U4956 ( .A1(n10483), .A2(n10485), .ZN(n7993) );
  INV_X1 U4957 ( .A(n9496), .ZN(n10423) );
  INV_X1 U4958 ( .A(n7997), .ZN(n10463) );
  NAND2_X1 U4959 ( .A1(n7687), .A2(n7885), .ZN(n6797) );
  INV_X2 U4960 ( .A(n6975), .ZN(n7701) );
  INV_X1 U4963 ( .A(n7064), .ZN(n4850) );
  NAND2_X1 U4965 ( .A1(n8311), .A2(n9991), .ZN(n7064) );
  INV_X4 U4966 ( .A(n5745), .ZN(n6007) );
  NAND2_X1 U4967 ( .A1(n9371), .A2(n6223), .ZN(n6228) );
  AND2_X1 U4968 ( .A1(n7172), .A2(n6238), .ZN(n6259) );
  NAND2_X1 U4969 ( .A1(n6631), .A2(n4855), .ZN(n6236) );
  INV_X4 U4970 ( .A(n5552), .ZN(n5418) );
  NAND2_X2 U4971 ( .A1(n5292), .A2(n5293), .ZN(n5552) );
  AOI21_X1 U4972 ( .B1(n8592), .B2(n10522), .A(n8591), .ZN(n10089) );
  XNOR2_X1 U4973 ( .A(n8584), .B(n8586), .ZN(n10090) );
  OAI22_X1 U4974 ( .A1(n6617), .A2(n6634), .B1(n8203), .B2(n8929), .ZN(n6619)
         );
  NAND2_X1 U4975 ( .A1(n9084), .A2(n6595), .ZN(n9065) );
  CLKBUF_X1 U4976 ( .A(n9112), .Z(n9122) );
  OAI21_X1 U4977 ( .B1(n9953), .B2(n7053), .A(n7052), .ZN(n9929) );
  AOI21_X1 U4978 ( .B1(n5365), .B2(n5369), .A(n4889), .ZN(n5364) );
  NAND2_X1 U4979 ( .A1(n9205), .A2(n9212), .ZN(n9204) );
  AND2_X1 U4980 ( .A1(n7054), .A2(n6131), .ZN(n9928) );
  NAND2_X1 U4981 ( .A1(n9221), .A2(n9224), .ZN(n9222) );
  OR2_X1 U4982 ( .A1(n10092), .A2(n9543), .ZN(n6133) );
  OR2_X1 U4983 ( .A1(n9159), .A2(n9143), .ZN(n6752) );
  NAND2_X1 U4984 ( .A1(n6043), .A2(n6042), .ZN(n10092) );
  XNOR2_X1 U4985 ( .A(n5623), .B(n5622), .ZN(n10205) );
  NAND2_X1 U4986 ( .A1(n5336), .A2(n5337), .ZN(n9238) );
  NAND2_X1 U4987 ( .A1(n6541), .A2(n6540), .ZN(n9304) );
  NAND2_X1 U4988 ( .A1(n6530), .A2(n6529), .ZN(n9159) );
  NAND2_X1 U4989 ( .A1(n6917), .A2(n8782), .ZN(n8789) );
  NOR2_X1 U4990 ( .A1(n8322), .A2(n5242), .ZN(n5023) );
  NAND2_X1 U4991 ( .A1(n5658), .A2(n5509), .ZN(n5661) );
  NAND2_X1 U4992 ( .A1(n6493), .A2(n6492), .ZN(n9333) );
  NAND2_X1 U4993 ( .A1(n6523), .A2(n6522), .ZN(n9316) );
  NAND2_X1 U4994 ( .A1(n6481), .A2(n6480), .ZN(n9336) );
  NAND2_X1 U4995 ( .A1(n10532), .A2(n7102), .ZN(n8075) );
  NAND2_X1 U4996 ( .A1(n5978), .A2(n5977), .ZN(n10135) );
  NAND2_X1 U4997 ( .A1(n6462), .A2(n6461), .ZN(n9343) );
  AND2_X1 U4998 ( .A1(n5321), .A2(n8316), .ZN(n5320) );
  NAND2_X1 U4999 ( .A1(n5687), .A2(n5686), .ZN(n10117) );
  NAND2_X1 U5000 ( .A1(n5180), .A2(n5181), .ZN(n8293) );
  NAND2_X1 U5001 ( .A1(n5955), .A2(n5954), .ZN(n10141) );
  NAND2_X1 U5002 ( .A1(n6391), .A2(n6390), .ZN(n8411) );
  AND2_X1 U5003 ( .A1(n6100), .A2(n7030), .ZN(n8192) );
  NOR2_X1 U5004 ( .A1(n5343), .A2(n5342), .ZN(n5341) );
  NAND2_X1 U5005 ( .A1(n6374), .A2(n6373), .ZN(n10640) );
  NAND2_X1 U5006 ( .A1(n10542), .A2(n6163), .ZN(n8013) );
  AND2_X1 U5007 ( .A1(n5145), .A2(n5294), .ZN(n7782) );
  NAND2_X1 U5008 ( .A1(n5454), .A2(n9614), .ZN(n5290) );
  INV_X1 U5009 ( .A(n10595), .ZN(n8179) );
  OR2_X1 U5010 ( .A1(n5453), .A2(n5452), .ZN(n5455) );
  OAI21_X1 U5011 ( .B1(n7247), .B2(n6328), .A(n4991), .ZN(n10525) );
  XNOR2_X1 U5012 ( .A(n5823), .B(n5822), .ZN(n7247) );
  NAND2_X1 U5013 ( .A1(n9791), .A2(n10463), .ZN(n10485) );
  AND3_X1 U5014 ( .A1(n6313), .A2(n6312), .A3(n6311), .ZN(n10509) );
  NAND2_X1 U5015 ( .A1(n4966), .A2(n5434), .ZN(n5835) );
  INV_X2 U5016 ( .A(n6242), .ZN(n6860) );
  AND2_X2 U5017 ( .A1(n5253), .A2(n8718), .ZN(n8720) );
  NAND2_X2 U5019 ( .A1(n5322), .A2(n5323), .ZN(n6960) );
  NAND2_X1 U5020 ( .A1(n5768), .A2(n5767), .ZN(n5777) );
  NAND2_X1 U5021 ( .A1(n6265), .A2(n5247), .ZN(n7738) );
  AND2_X2 U5022 ( .A1(n7262), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U4006) );
  AND4_X1 U5023 ( .A1(n5738), .A2(n5737), .A3(n5736), .A4(n5735), .ZN(n7763)
         );
  AND2_X1 U5024 ( .A1(n5128), .A2(n4860), .ZN(n5127) );
  BUF_X2 U5025 ( .A(n5762), .Z(n6047) );
  OAI211_X1 U5026 ( .C1(n6328), .C2(n7237), .A(n5139), .B(n5138), .ZN(n7885)
         );
  NAND2_X1 U5027 ( .A1(n7377), .A2(n7375), .ZN(n8702) );
  NAND2_X2 U5028 ( .A1(n9375), .A2(n6228), .ZN(n6498) );
  NAND2_X1 U5029 ( .A1(n6203), .A2(n5025), .ZN(n7377) );
  AND2_X1 U5030 ( .A1(n5603), .A2(n5602), .ZN(n5762) );
  AND2_X1 U5031 ( .A1(n8825), .A2(n5603), .ZN(n5763) );
  NAND2_X1 U5032 ( .A1(n5395), .A2(n5022), .ZN(n7766) );
  NAND2_X1 U5033 ( .A1(n5559), .A2(n5560), .ZN(n8825) );
  NAND2_X1 U5034 ( .A1(n4959), .A2(n5417), .ZN(n5773) );
  OR2_X1 U5035 ( .A1(n6221), .A2(n9370), .ZN(n6220) );
  NAND2_X1 U5036 ( .A1(n6491), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6626) );
  NAND2_X1 U5037 ( .A1(n6237), .A2(n6236), .ZN(n9385) );
  MUX2_X1 U5038 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6232), .S(
        P2_IR_REG_28__SCAN_IN), .Z(n6234) );
  NAND2_X1 U5039 ( .A1(n5543), .A2(n5542), .ZN(n5544) );
  NAND2_X1 U5040 ( .A1(n5436), .A2(n9586), .ZN(n5439) );
  NAND2_X2 U5041 ( .A1(n5021), .A2(P2_U3152), .ZN(n8243) );
  XNOR2_X1 U5042 ( .A(n5259), .B(P1_IR_REG_19__SCAN_IN), .ZN(n9991) );
  AND2_X1 U5043 ( .A1(n5381), .A2(n5379), .ZN(n4998) );
  AND2_X1 U5044 ( .A1(n4897), .A2(n4847), .ZN(n5219) );
  AND2_X1 U5045 ( .A1(n5380), .A2(n5185), .ZN(n4999) );
  AND2_X1 U5046 ( .A1(n5188), .A2(n4875), .ZN(n5185) );
  AND2_X1 U5047 ( .A1(n5375), .A2(n5540), .ZN(n5374) );
  AND2_X1 U5048 ( .A1(n5404), .A2(n5189), .ZN(n5188) );
  AND2_X1 U5049 ( .A1(n6323), .A2(n6385), .ZN(n5222) );
  AND4_X1 U5050 ( .A1(n5398), .A2(n5399), .A3(n5403), .A4(n5402), .ZN(n5381)
         );
  INV_X1 U5051 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n6198) );
  INV_X1 U5052 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n6201) );
  NOR2_X1 U5053 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n5397) );
  NOR2_X1 U5054 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n5403) );
  NOR2_X1 U5055 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n5402) );
  NOR2_X1 U5056 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n5401) );
  NOR2_X1 U5057 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n5396) );
  INV_X1 U5058 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5404) );
  INV_X1 U5059 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n6211) );
  INV_X1 U5060 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n6625) );
  INV_X1 U5061 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n6323) );
  INV_X1 U5062 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n6489) );
  NOR2_X1 U5063 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n5400) );
  INV_X1 U5064 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n6385) );
  INV_X1 U5065 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n6386) );
  INV_X1 U5066 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n6401) );
  INV_X1 U5067 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n6415) );
  INV_X1 U5068 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n6431) );
  INV_X1 U5069 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6834) );
  INV_X1 U5070 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n6216) );
  NOR2_X2 U5071 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n5326) );
  OAI21_X1 U5072 ( .B1(n8296), .B2(n5372), .A(n5370), .ZN(n7111) );
  OR3_X2 U5073 ( .A1(n6703), .A2(n6702), .A3(n8377), .ZN(n6710) );
  OAI22_X2 U5074 ( .A1(n7858), .A2(n6314), .B1(n10509), .B2(n8941), .ZN(n7978)
         );
  NAND2_X1 U5075 ( .A1(n6205), .A2(n10260), .ZN(n4853) );
  NAND2_X1 U5076 ( .A1(n6205), .A2(n10260), .ZN(n4854) );
  NAND2_X4 U5077 ( .A1(n6205), .A2(n10260), .ZN(n5745) );
  OR2_X1 U5078 ( .A1(n8919), .A2(n4913), .ZN(n5310) );
  OR2_X1 U5079 ( .A1(n9304), .A2(n8868), .ZN(n6763) );
  NAND2_X1 U5080 ( .A1(n4976), .A2(n4973), .ZN(n10604) );
  NAND2_X1 U5081 ( .A1(n7970), .A2(n5341), .ZN(n4976) );
  AND2_X1 U5082 ( .A1(n4903), .A2(n4974), .ZN(n4973) );
  AND2_X1 U5083 ( .A1(n6213), .A2(n6458), .ZN(n6214) );
  NAND2_X1 U5084 ( .A1(n7640), .A2(n5028), .ZN(n7641) );
  NAND2_X1 U5085 ( .A1(n8720), .A2(n5029), .ZN(n5028) );
  INV_X1 U5086 ( .A(n8825), .ZN(n5602) );
  NAND2_X1 U5087 ( .A1(n8464), .A2(n8463), .ZN(n5027) );
  INV_X1 U5088 ( .A(n5771), .ZN(n6008) );
  NAND2_X1 U5089 ( .A1(n5137), .A2(n5134), .ZN(n5133) );
  NOR2_X1 U5090 ( .A1(n5136), .A2(n5135), .ZN(n5134) );
  NAND2_X1 U5091 ( .A1(n6780), .A2(n6779), .ZN(n5135) );
  NOR2_X1 U5092 ( .A1(n9162), .A2(n5228), .ZN(n5227) );
  INV_X1 U5093 ( .A(n6751), .ZN(n5228) );
  AOI21_X1 U5094 ( .B1(n4860), .B2(n5271), .A(n4886), .ZN(n5267) );
  NAND2_X1 U5095 ( .A1(n5127), .A2(n5130), .ZN(n5125) );
  AND2_X1 U5096 ( .A1(n5132), .A2(n5389), .ZN(n5131) );
  NAND2_X1 U5097 ( .A1(n5834), .A2(n5439), .ZN(n5132) );
  NAND2_X1 U5098 ( .A1(n6854), .A2(n6842), .ZN(n5323) );
  NAND3_X1 U5099 ( .A1(n6853), .A2(n6852), .A3(n6854), .ZN(n5322) );
  INV_X1 U5100 ( .A(n7431), .ZN(n6854) );
  XNOR2_X1 U5101 ( .A(n7707), .B(n6960), .ZN(n6862) );
  INV_X1 U5102 ( .A(n9115), .ZN(n5335) );
  OR2_X1 U5103 ( .A1(n9295), .A2(n8829), .ZN(n6792) );
  NAND2_X1 U5104 ( .A1(n9123), .A2(n9124), .ZN(n9112) );
  AOI21_X1 U5105 ( .B1(n5227), .B2(n5225), .A(n5224), .ZN(n5223) );
  OR2_X1 U5106 ( .A1(n9326), .A2(n9196), .ZN(n6743) );
  OR2_X1 U5107 ( .A1(n9321), .A2(n9214), .ZN(n6645) );
  INV_X1 U5108 ( .A(n8132), .ZN(n5342) );
  NAND2_X1 U5109 ( .A1(n10595), .A2(n8939), .ZN(n6680) );
  NOR2_X1 U5110 ( .A1(n5170), .A2(n10525), .ZN(n5168) );
  NAND2_X1 U5111 ( .A1(n6658), .A2(n6657), .ZN(n7860) );
  INV_X1 U5112 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5348) );
  INV_X1 U5113 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6215) );
  AND2_X1 U5114 ( .A1(n10072), .A2(n9899), .ZN(n6072) );
  OR2_X1 U5115 ( .A1(n6044), .A2(n9447), .ZN(n6046) );
  OR2_X1 U5116 ( .A1(n10146), .A2(n9465), .ZN(n6109) );
  NAND2_X1 U5117 ( .A1(n9897), .A2(n8810), .ZN(n8812) );
  OR2_X1 U5118 ( .A1(n7388), .A2(n7650), .ZN(n7409) );
  AND2_X1 U5119 ( .A1(n5522), .A2(n5521), .ZN(n5634) );
  INV_X1 U5120 ( .A(n4998), .ZN(n5190) );
  NAND2_X1 U5121 ( .A1(n6006), .A2(n5489), .ZN(n5685) );
  NAND2_X1 U5122 ( .A1(n4894), .A2(n4863), .ZN(n5265) );
  NAND2_X1 U5123 ( .A1(n5481), .A2(n5480), .ZN(n5266) );
  INV_X1 U5124 ( .A(n5990), .ZN(n5484) );
  AND2_X1 U5125 ( .A1(n5910), .A2(n5909), .ZN(n5914) );
  INV_X1 U5126 ( .A(SI_14_), .ZN(n5463) );
  OAI21_X1 U5127 ( .B1(n5552), .B2(n4986), .A(n4985), .ZN(n5425) );
  NAND2_X1 U5128 ( .A1(n5552), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n4985) );
  OR2_X1 U5129 ( .A1(n5702), .A2(P1_IR_REG_3__SCAN_IN), .ZN(n5752) );
  AND2_X1 U5130 ( .A1(n5308), .A2(n7000), .ZN(n5307) );
  NAND2_X1 U5131 ( .A1(n7829), .A2(n5150), .ZN(n7142) );
  NOR2_X1 U5132 ( .A1(n6860), .A2(n7701), .ZN(n6861) );
  INV_X1 U5133 ( .A(n6273), .ZN(n6612) );
  AND3_X1 U5134 ( .A1(n6839), .A2(n10308), .A3(n10307), .ZN(n7157) );
  AOI21_X1 U5135 ( .B1(n5330), .B2(n5332), .A(n4880), .ZN(n5328) );
  NAND2_X1 U5136 ( .A1(n9164), .A2(n4878), .ZN(n9135) );
  OR2_X1 U5137 ( .A1(n9316), .A2(n9197), .ZN(n6751) );
  NAND2_X1 U5138 ( .A1(n9175), .A2(n9174), .ZN(n9173) );
  OR2_X1 U5139 ( .A1(n9321), .A2(n9176), .ZN(n9052) );
  OR2_X1 U5140 ( .A1(n10661), .A2(n8783), .ZN(n6712) );
  OR2_X1 U5141 ( .A1(n6301), .A2(n6300), .ZN(n5246) );
  NAND2_X1 U5142 ( .A1(n7861), .A2(n7860), .ZN(n5345) );
  NOR2_X1 U5143 ( .A1(n7431), .A2(n7430), .ZN(n10436) );
  AND2_X1 U5144 ( .A1(n10307), .A2(n6987), .ZN(n10212) );
  AND2_X1 U5145 ( .A1(n6211), .A2(n6610), .ZN(n5218) );
  OR2_X1 U5146 ( .A1(n9538), .A2(n5048), .ZN(n5047) );
  NAND2_X1 U5147 ( .A1(n7376), .A2(n8311), .ZN(n5253) );
  NAND2_X1 U5148 ( .A1(n5027), .A2(n4911), .ZN(n8610) );
  NOR2_X1 U5149 ( .A1(n8452), .A2(n5026), .ZN(n5025) );
  OR2_X1 U5150 ( .A1(n7390), .A2(n7388), .ZN(n7514) );
  AND2_X1 U5151 ( .A1(n5579), .A2(n9884), .ZN(n6184) );
  NAND2_X1 U5152 ( .A1(n4937), .A2(n4873), .ZN(n6148) );
  OR2_X1 U5153 ( .A1(n6063), .A2(n4938), .ZN(n4937) );
  AND3_X1 U5154 ( .A1(n5683), .A2(n5682), .A3(n5681), .ZN(n10000) );
  NAND2_X1 U5155 ( .A1(n10538), .A2(n10580), .ZN(n5377) );
  NAND2_X1 U5156 ( .A1(n8075), .A2(n5378), .ZN(n5376) );
  OR2_X1 U5157 ( .A1(n10538), .A2(n10580), .ZN(n5378) );
  NAND2_X1 U5158 ( .A1(n6010), .A2(n6009), .ZN(n10123) );
  OR2_X1 U5159 ( .A1(n7064), .A2(n7063), .ZN(n10370) );
  INV_X1 U5160 ( .A(n5551), .ZN(n5545) );
  AND2_X1 U5161 ( .A1(n6070), .A2(n6071), .ZN(n7130) );
  NOR2_X1 U5162 ( .A1(n6849), .A2(n8203), .ZN(n7431) );
  NAND2_X1 U5163 ( .A1(n5625), .A2(n5624), .ZN(n10082) );
  AND2_X1 U5164 ( .A1(n5841), .A2(n7028), .ZN(n4931) );
  NOR2_X1 U5165 ( .A1(n4928), .A2(n8207), .ZN(n4927) );
  INV_X1 U5166 ( .A(n5871), .ZN(n4928) );
  NAND2_X1 U5167 ( .A1(n6055), .A2(n9921), .ZN(n4923) );
  INV_X1 U5168 ( .A(n6056), .ZN(n4924) );
  NAND2_X1 U5169 ( .A1(n6636), .A2(n6775), .ZN(n5272) );
  NAND2_X1 U5170 ( .A1(n6789), .A2(n6782), .ZN(n5274) );
  INV_X1 U5171 ( .A(n5462), .ZN(n5115) );
  INV_X1 U5172 ( .A(SI_13_), .ZN(n9675) );
  INV_X1 U5173 ( .A(n4969), .ZN(n4968) );
  OAI21_X1 U5174 ( .B1(n5429), .B2(n4970), .A(n5822), .ZN(n4969) );
  INV_X1 U5175 ( .A(n5431), .ZN(n4970) );
  NOR2_X1 U5176 ( .A1(n9280), .A2(n5154), .ZN(n5153) );
  NAND2_X1 U5177 ( .A1(n5155), .A2(n9097), .ZN(n5154) );
  OR2_X1 U5178 ( .A1(n9316), .A2(n9321), .ZN(n5160) );
  AND2_X1 U5179 ( .A1(n6731), .A2(n6732), .ZN(n6738) );
  AND2_X1 U5180 ( .A1(n5165), .A2(n5164), .ZN(n5163) );
  OR2_X1 U5181 ( .A1(n8781), .A2(n8505), .ZN(n6716) );
  AND2_X1 U5182 ( .A1(n6705), .A2(n6704), .ZN(n6805) );
  INV_X1 U5183 ( .A(n7967), .ZN(n4994) );
  NAND2_X1 U5184 ( .A1(n8059), .A2(n10509), .ZN(n5170) );
  NAND2_X1 U5185 ( .A1(n8057), .A2(n7864), .ZN(n5349) );
  INV_X1 U5186 ( .A(n6849), .ZN(n5144) );
  NAND2_X1 U5187 ( .A1(n6849), .A2(n7180), .ZN(n6850) );
  OR2_X1 U5188 ( .A1(n6849), .A2(n8307), .ZN(n6851) );
  INV_X1 U5189 ( .A(n8708), .ZN(n5048) );
  NAND2_X1 U5190 ( .A1(n8097), .A2(n8096), .ZN(n5036) );
  NOR2_X1 U5191 ( .A1(n5032), .A2(n5035), .ZN(n5031) );
  INV_X1 U5192 ( .A(n8096), .ZN(n5032) );
  NOR2_X1 U5193 ( .A1(n8152), .A2(n8101), .ZN(n5035) );
  INV_X1 U5194 ( .A(n8157), .ZN(n5251) );
  INV_X1 U5195 ( .A(n8693), .ZN(n5237) );
  OR2_X1 U5196 ( .A1(n10067), .A2(n6087), .ZN(n6089) );
  OR2_X1 U5197 ( .A1(n10076), .A2(n9396), .ZN(n8810) );
  NAND2_X1 U5198 ( .A1(n5599), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n6044) );
  OR2_X1 U5199 ( .A1(n10097), .A2(n9448), .ZN(n7054) );
  NAND2_X1 U5200 ( .A1(n4869), .A2(n7119), .ZN(n5360) );
  NOR2_X1 U5201 ( .A1(n9997), .A2(n5362), .ZN(n5361) );
  INV_X1 U5202 ( .A(n7119), .ZN(n5362) );
  OR2_X1 U5203 ( .A1(n10135), .A2(n10035), .ZN(n7043) );
  INV_X1 U5204 ( .A(n7108), .ZN(n5372) );
  OR2_X1 U5205 ( .A1(n10152), .A2(n8525), .ZN(n7037) );
  NOR2_X1 U5206 ( .A1(n10544), .A2(n5355), .ZN(n5354) );
  INV_X1 U5207 ( .A(n7100), .ZN(n5355) );
  NAND2_X1 U5208 ( .A1(n6075), .A2(n10407), .ZN(n7743) );
  NOR2_X1 U5209 ( .A1(n5514), .A2(n5289), .ZN(n5288) );
  INV_X1 U5210 ( .A(n5510), .ZN(n5289) );
  INV_X1 U5211 ( .A(n5121), .ZN(n5120) );
  AND2_X1 U5212 ( .A1(n5118), .A2(n5262), .ZN(n5117) );
  AOI21_X1 U5213 ( .B1(n5265), .B2(n5263), .A(n6004), .ZN(n5262) );
  NAND2_X1 U5214 ( .A1(n5123), .A2(n5478), .ZN(n5969) );
  NAND2_X1 U5215 ( .A1(n5290), .A2(n5455), .ZN(n5891) );
  NAND2_X1 U5216 ( .A1(n5891), .A2(n5461), .ZN(n5894) );
  AND2_X1 U5217 ( .A1(n5876), .A2(n5875), .ZN(n5910) );
  AOI21_X1 U5218 ( .B1(n5390), .B2(n5270), .A(n5269), .ZN(n5268) );
  INV_X1 U5219 ( .A(n5444), .ZN(n5270) );
  INV_X1 U5220 ( .A(n5449), .ZN(n5269) );
  INV_X1 U5221 ( .A(SI_11_), .ZN(n5450) );
  NAND2_X1 U5222 ( .A1(n5126), .A2(n5131), .ZN(n5445) );
  XNOR2_X1 U5223 ( .A(n5430), .B(SI_6_), .ZN(n5806) );
  INV_X1 U5224 ( .A(n5423), .ZN(n5099) );
  INV_X1 U5225 ( .A(SI_4_), .ZN(n4984) );
  OAI21_X1 U5226 ( .B1(n5418), .B2(n5420), .A(n5419), .ZN(n5422) );
  NAND2_X1 U5227 ( .A1(n5418), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n5419) );
  OAI21_X1 U5228 ( .B1(n5418), .B2(n5415), .A(n5414), .ZN(n5416) );
  NAND2_X1 U5229 ( .A1(n5730), .A2(n6250), .ZN(n5412) );
  NAND2_X1 U5230 ( .A1(n8864), .A2(n5143), .ZN(n5142) );
  OR2_X1 U5231 ( .A1(n6524), .A2(n8895), .ZN(n6532) );
  AND2_X1 U5232 ( .A1(n5305), .A2(n5311), .ZN(n5304) );
  NAND2_X1 U5233 ( .A1(n5308), .A2(n5306), .ZN(n5305) );
  INV_X1 U5234 ( .A(n7005), .ZN(n5311) );
  INV_X1 U5235 ( .A(n5304), .ZN(n5302) );
  INV_X1 U5236 ( .A(n6316), .ZN(n6315) );
  OR2_X1 U5237 ( .A1(n6331), .A2(n8068), .ZN(n6346) );
  NAND2_X1 U5238 ( .A1(n8574), .A2(n5250), .ZN(n5112) );
  INV_X1 U5239 ( .A(n6376), .ZN(n6375) );
  XNOR2_X1 U5240 ( .A(n7885), .B(n6960), .ZN(n6856) );
  OAI21_X1 U5241 ( .B1(n6874), .B2(n5317), .A(n6877), .ZN(n5316) );
  AND2_X1 U5242 ( .A1(n7445), .A2(n7690), .ZN(n7007) );
  OR2_X1 U5243 ( .A1(n6908), .A2(n4857), .ZN(n5321) );
  INV_X1 U5244 ( .A(n5320), .ZN(n5148) );
  AND4_X1 U5245 ( .A1(n6364), .A2(n6363), .A3(n6362), .A4(n6361), .ZN(n8246)
         );
  NAND2_X1 U5246 ( .A1(n6848), .A2(n6842), .ZN(n7180) );
  OAI21_X1 U5247 ( .B1(n9058), .B2(n5085), .A(n6768), .ZN(n5084) );
  INV_X1 U5248 ( .A(n6791), .ZN(n5085) );
  AND2_X1 U5249 ( .A1(n5335), .A2(n9057), .ZN(n5334) );
  AOI21_X1 U5250 ( .B1(n5335), .B2(n4858), .A(n4888), .ZN(n5333) );
  NOR2_X1 U5251 ( .A1(n9127), .A2(n9295), .ZN(n9107) );
  INV_X1 U5252 ( .A(n9124), .ZN(n9057) );
  AND2_X1 U5253 ( .A1(n6792), .A2(n6791), .ZN(n9115) );
  AND2_X1 U5254 ( .A1(n6762), .A2(n9113), .ZN(n9124) );
  NAND2_X1 U5255 ( .A1(n9055), .A2(n8868), .ZN(n9056) );
  NAND2_X1 U5256 ( .A1(n5082), .A2(n5223), .ZN(n9142) );
  INV_X1 U5257 ( .A(n5223), .ZN(n5081) );
  OR2_X1 U5258 ( .A1(n9175), .A2(n5226), .ZN(n5082) );
  NAND2_X1 U5259 ( .A1(n9172), .A2(n9197), .ZN(n4989) );
  NAND2_X1 U5260 ( .A1(n9168), .A2(n5225), .ZN(n4990) );
  AND3_X1 U5261 ( .A1(n9311), .A2(n5159), .A3(n5158), .ZN(n9155) );
  INV_X1 U5262 ( .A(n5160), .ZN(n5158) );
  NAND2_X1 U5263 ( .A1(n9222), .A2(n9050), .ZN(n9205) );
  INV_X1 U5264 ( .A(n5215), .ZN(n5214) );
  OAI21_X1 U5265 ( .B1(n9237), .B2(n5216), .A(n6738), .ZN(n5215) );
  INV_X1 U5266 ( .A(n9225), .ZN(n5216) );
  AOI21_X1 U5267 ( .B1(n9238), .B2(n9246), .A(n9048), .ZN(n9221) );
  NOR2_X1 U5268 ( .A1(n9336), .A2(n8932), .ZN(n9048) );
  INV_X1 U5269 ( .A(n6738), .ZN(n9224) );
  AND2_X1 U5270 ( .A1(n9263), .A2(n4896), .ZN(n5339) );
  OR2_X1 U5271 ( .A1(n8540), .A2(n8541), .ZN(n5340) );
  AND2_X1 U5272 ( .A1(n9257), .A2(n9256), .ZN(n8541) );
  AND2_X1 U5273 ( .A1(n6716), .A2(n6715), .ZN(n8538) );
  INV_X1 U5274 ( .A(n6805), .ZN(n8377) );
  AND2_X1 U5275 ( .A1(n8284), .A2(n8281), .ZN(n5351) );
  AND2_X1 U5276 ( .A1(n6688), .A2(n6685), .ZN(n10610) );
  AND4_X1 U5277 ( .A1(n6353), .A2(n6352), .A3(n6351), .A4(n6350), .ZN(n10612)
         );
  INV_X1 U5278 ( .A(n10611), .ZN(n9177) );
  AND2_X1 U5279 ( .A1(n10437), .A2(n7862), .ZN(n5344) );
  NOR2_X1 U5280 ( .A1(n7885), .A2(n7565), .ZN(n7703) );
  AND4_X1 U5281 ( .A1(n6271), .A2(n6270), .A3(n6269), .A4(n6268), .ZN(n10438)
         );
  INV_X1 U5282 ( .A(n9178), .ZN(n10613) );
  NAND2_X1 U5283 ( .A1(n7567), .A2(n5144), .ZN(n7699) );
  AND2_X1 U5284 ( .A1(n6841), .A2(n7159), .ZN(n9178) );
  NAND2_X1 U5285 ( .A1(n6853), .A2(n6852), .ZN(n10619) );
  NAND2_X1 U5286 ( .A1(n9280), .A2(n10662), .ZN(n5093) );
  NAND2_X1 U5287 ( .A1(n6582), .A2(n5250), .ZN(n6584) );
  AND2_X1 U5288 ( .A1(n6327), .A2(n6326), .ZN(n4991) );
  AND3_X1 U5289 ( .A1(n6284), .A2(n6283), .A3(n6282), .ZN(n10434) );
  INV_X1 U5290 ( .A(n7442), .ZN(n10213) );
  AND2_X1 U5291 ( .A1(n5388), .A2(n4865), .ZN(n5346) );
  INV_X1 U5292 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5347) );
  INV_X2 U5293 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n6628) );
  AND2_X1 U5294 ( .A1(n6459), .A2(n6458), .ZN(n6479) );
  XNOR2_X1 U5295 ( .A(n4996), .B(P2_IR_REG_1__SCAN_IN), .ZN(n10319) );
  NAND2_X1 U5296 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n4996) );
  NAND2_X1 U5297 ( .A1(n8610), .A2(n8609), .ZN(n5209) );
  INV_X1 U5298 ( .A(n7641), .ZN(n7643) );
  INV_X1 U5299 ( .A(n9528), .ZN(n5069) );
  INV_X1 U5300 ( .A(n5063), .ZN(n5062) );
  OAI21_X1 U5301 ( .B1(n5071), .B2(n5064), .A(n9528), .ZN(n5063) );
  INV_X1 U5302 ( .A(n5066), .ZN(n5065) );
  OAI21_X1 U5303 ( .B1(n5064), .B2(n5067), .A(n9527), .ZN(n5066) );
  NAND2_X1 U5304 ( .A1(n5072), .A2(n5069), .ZN(n5067) );
  XNOR2_X1 U5305 ( .A(n7494), .B(n8711), .ZN(n7506) );
  NAND2_X1 U5306 ( .A1(n5238), .A2(n9482), .ZN(n9479) );
  AND2_X1 U5307 ( .A1(n9481), .A2(n9480), .ZN(n5238) );
  NAND2_X1 U5308 ( .A1(n5036), .A2(n8102), .ZN(n8153) );
  NAND2_X1 U5309 ( .A1(n5033), .A2(n8101), .ZN(n8154) );
  INV_X1 U5310 ( .A(n5036), .ZN(n5033) );
  NOR2_X1 U5311 ( .A1(n7379), .A2(n5254), .ZN(n7384) );
  AND2_X1 U5312 ( .A1(n7380), .A2(n8720), .ZN(n5254) );
  NAND2_X1 U5313 ( .A1(n7383), .A2(n7382), .ZN(n7495) );
  NAND2_X1 U5314 ( .A1(n5596), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n6014) );
  NAND2_X1 U5315 ( .A1(n6007), .A2(n5172), .ZN(n5171) );
  INV_X1 U5316 ( .A(n7234), .ZN(n5174) );
  AOI21_X1 U5317 ( .B1(n5071), .B2(n8630), .A(n4887), .ZN(n5070) );
  NAND2_X1 U5318 ( .A1(n5205), .A2(n5208), .ZN(n5199) );
  NAND2_X1 U5319 ( .A1(n5202), .A2(n5204), .ZN(n5201) );
  NOR2_X1 U5320 ( .A1(n4856), .A2(n8683), .ZN(n5233) );
  NOR2_X1 U5321 ( .A1(n4856), .A2(n5236), .ZN(n5235) );
  INV_X1 U5322 ( .A(n9415), .ZN(n5236) );
  NOR2_X1 U5323 ( .A1(n4856), .A2(n9480), .ZN(n5232) );
  INV_X1 U5324 ( .A(n9443), .ZN(n5234) );
  NAND2_X1 U5325 ( .A1(n8682), .A2(n8683), .ZN(n9413) );
  AND2_X1 U5326 ( .A1(n10076), .A2(n9570), .ZN(n8794) );
  NAND2_X1 U5327 ( .A1(n8801), .A2(n8800), .ZN(n9907) );
  INV_X1 U5328 ( .A(n10076), .ZN(n8800) );
  AND2_X1 U5329 ( .A1(n5633), .A2(n5632), .ZN(n9898) );
  NOR2_X1 U5330 ( .A1(n8595), .A2(n10082), .ZN(n8801) );
  INV_X1 U5331 ( .A(n5368), .ZN(n5367) );
  OAI22_X1 U5332 ( .A1(n7055), .A2(n5369), .B1(n9549), .B2(n9451), .ZN(n5368)
         );
  NAND2_X1 U5333 ( .A1(n8587), .A2(n10546), .ZN(n8590) );
  INV_X1 U5334 ( .A(n5195), .ZN(n5194) );
  AOI21_X1 U5335 ( .B1(n5195), .B2(n5193), .A(n5192), .ZN(n5191) );
  NOR2_X1 U5336 ( .A1(n5197), .A2(n5196), .ZN(n5195) );
  NAND2_X1 U5337 ( .A1(n10020), .A2(n10021), .ZN(n10019) );
  AND2_X1 U5338 ( .A1(n6114), .A2(n7045), .ZN(n10021) );
  NOR2_X1 U5339 ( .A1(n10057), .A2(n10043), .ZN(n10039) );
  NAND2_X1 U5340 ( .A1(n6111), .A2(n7044), .ZN(n10032) );
  NAND2_X1 U5341 ( .A1(n5353), .A2(n4877), .ZN(n8555) );
  NAND2_X1 U5342 ( .A1(n8518), .A2(n7112), .ZN(n5352) );
  AND4_X1 U5343 ( .A1(n5906), .A2(n5905), .A3(n5904), .A4(n5903), .ZN(n8472)
         );
  AOI21_X1 U5344 ( .B1(n7031), .B2(n5183), .A(n5182), .ZN(n5181) );
  NAND2_X1 U5345 ( .A1(n8187), .A2(n4972), .ZN(n5180) );
  INV_X1 U5346 ( .A(n7032), .ZN(n5182) );
  INV_X1 U5347 ( .A(n5865), .ZN(n5591) );
  INV_X1 U5348 ( .A(n8192), .ZN(n7103) );
  OAI21_X1 U5349 ( .B1(n10486), .B2(n7021), .A(n7022), .ZN(n8009) );
  NAND2_X1 U5350 ( .A1(n7664), .A2(n6154), .ZN(n4943) );
  NOR2_X1 U5351 ( .A1(n7758), .A2(n10364), .ZN(n7749) );
  OR2_X1 U5352 ( .A1(n10370), .A2(n7130), .ZN(n7406) );
  NAND2_X1 U5353 ( .A1(n5021), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n5020) );
  NAND2_X1 U5354 ( .A1(n5587), .A2(n5586), .ZN(n10072) );
  NAND2_X1 U5355 ( .A1(n8818), .A2(n8817), .ZN(n8819) );
  AND2_X1 U5356 ( .A1(n7412), .A2(n7668), .ZN(n10365) );
  INV_X1 U5357 ( .A(n7766), .ZN(n10357) );
  NAND2_X1 U5358 ( .A1(n7377), .A2(n6204), .ZN(n7388) );
  OR2_X1 U5359 ( .A1(n7067), .A2(n7066), .ZN(n7403) );
  AOI21_X1 U5360 ( .B1(n5278), .B2(n5280), .A(n4919), .ZN(n5275) );
  XNOR2_X1 U5361 ( .A(n5570), .B(n5569), .ZN(n8790) );
  NAND2_X1 U5362 ( .A1(n5277), .A2(n5537), .ZN(n5570) );
  NAND2_X1 U5363 ( .A1(n5555), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5198) );
  NAND2_X1 U5364 ( .A1(n5547), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5548) );
  AOI21_X1 U5365 ( .B1(n5284), .B2(n4909), .A(n5283), .ZN(n5282) );
  NAND2_X1 U5366 ( .A1(n5539), .A2(n5374), .ZN(n6195) );
  XNOR2_X1 U5367 ( .A(n6149), .B(P1_IR_REG_20__SCAN_IN), .ZN(n7063) );
  OAI21_X1 U5368 ( .B1(n5186), .B2(n5190), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n6149) );
  INV_X1 U5369 ( .A(n5806), .ZN(n5429) );
  NAND2_X1 U5370 ( .A1(n5086), .A2(n5428), .ZN(n5807) );
  NOR2_X1 U5371 ( .A1(n5752), .A2(n5703), .ZN(n5803) );
  XNOR2_X1 U5372 ( .A(n5412), .B(n9728), .ZN(n5721) );
  NAND2_X1 U5373 ( .A1(n7829), .A2(n6881), .ZN(n7144) );
  NAND2_X1 U5374 ( .A1(n6419), .A2(n6418), .ZN(n10661) );
  INV_X1 U5375 ( .A(n7738), .ZN(n10392) );
  INV_X1 U5376 ( .A(n5307), .ZN(n5303) );
  AND3_X1 U5377 ( .A1(n6513), .A2(n6512), .A3(n6511), .ZN(n9196) );
  NAND2_X1 U5378 ( .A1(n7602), .A2(n5295), .ZN(n5294) );
  INV_X1 U5379 ( .A(n6865), .ZN(n5295) );
  OAI21_X1 U5380 ( .B1(n7829), .B2(n4956), .A(n4954), .ZN(n8167) );
  AND2_X1 U5381 ( .A1(n4955), .A2(n8062), .ZN(n4954) );
  OR2_X1 U5382 ( .A1(n5150), .A2(n4956), .ZN(n4955) );
  INV_X1 U5383 ( .A(n6887), .ZN(n4956) );
  AND3_X1 U5384 ( .A1(n6521), .A2(n6520), .A3(n6519), .ZN(n9214) );
  OR2_X1 U5385 ( .A1(n7616), .A2(n7615), .ZN(n4980) );
  OR2_X1 U5386 ( .A1(n8987), .A2(n8986), .ZN(n4993) );
  AND2_X1 U5387 ( .A1(n6561), .A2(n6553), .ZN(n9129) );
  NAND2_X1 U5388 ( .A1(n9173), .A2(n6751), .ZN(n9151) );
  AND2_X1 U5389 ( .A1(n8133), .A2(n8132), .ZN(n8134) );
  XNOR2_X1 U5390 ( .A(n6838), .B(P2_IR_REG_26__SCAN_IN), .ZN(n10307) );
  NAND2_X1 U5391 ( .A1(n9537), .A2(n8708), .ZN(n9392) );
  NAND2_X1 U5392 ( .A1(n5664), .A2(n5663), .ZN(n10102) );
  AND2_X1 U5393 ( .A1(n5045), .A2(n4868), .ZN(n5038) );
  NAND2_X1 U5394 ( .A1(n5882), .A2(n5881), .ZN(n10163) );
  NAND2_X1 U5395 ( .A1(n6027), .A2(n6026), .ZN(n10106) );
  AND2_X1 U5396 ( .A1(n6054), .A2(n6053), .ZN(n9543) );
  INV_X1 U5397 ( .A(n9561), .ZN(n9545) );
  OAI21_X1 U5398 ( .B1(n6148), .B2(n7138), .A(n6092), .ZN(n6146) );
  OR2_X1 U5399 ( .A1(n5017), .A2(n9888), .ZN(n5016) );
  INV_X1 U5400 ( .A(n5018), .ZN(n5017) );
  AOI21_X1 U5401 ( .B1(n9907), .B2(n10072), .A(n10582), .ZN(n5018) );
  AOI21_X1 U5402 ( .B1(n10082), .B2(n10042), .A(n7134), .ZN(n7135) );
  AOI21_X1 U5403 ( .B1(n4965), .B2(n10546), .A(n4964), .ZN(n10084) );
  OAI22_X1 U5404 ( .A1(n9396), .A2(n10489), .B1(n9451), .B2(n7059), .ZN(n4964)
         );
  XNOR2_X1 U5405 ( .A(n7058), .B(n8792), .ZN(n4965) );
  NAND2_X1 U5406 ( .A1(n9913), .A2(n7128), .ZN(n8584) );
  NAND2_X1 U5407 ( .A1(n5408), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5259) );
  OR2_X1 U5408 ( .A1(n7388), .A2(n7406), .ZN(n10005) );
  NAND2_X1 U5409 ( .A1(n10568), .A2(n7132), .ZN(n10565) );
  AND2_X1 U5410 ( .A1(n5541), .A2(n5556), .ZN(n5382) );
  INV_X1 U5411 ( .A(n9991), .ZN(n8116) );
  NOR2_X1 U5412 ( .A1(n8761), .A2(n8760), .ZN(n10244) );
  NOR2_X1 U5413 ( .A1(n10242), .A2(n10241), .ZN(n8760) );
  OAI211_X1 U5414 ( .C1(n4933), .C2(n5840), .A(n10544), .B(n5839), .ZN(n4932)
         );
  NAND2_X1 U5415 ( .A1(n4930), .A2(n5890), .ZN(n5925) );
  NAND2_X1 U5416 ( .A1(n5872), .A2(n4927), .ZN(n4930) );
  NAND2_X1 U5417 ( .A1(n5103), .A2(n4883), .ZN(n5102) );
  NAND2_X1 U5418 ( .A1(n9057), .A2(n4861), .ZN(n5100) );
  OR2_X1 U5419 ( .A1(n5988), .A2(n4850), .ZN(n4942) );
  INV_X1 U5420 ( .A(n6778), .ZN(n5136) );
  INV_X1 U5421 ( .A(SI_16_), .ZN(n9703) );
  INV_X1 U5422 ( .A(SI_15_), .ZN(n9705) );
  INV_X1 U5423 ( .A(n5131), .ZN(n5130) );
  NAND2_X1 U5424 ( .A1(n5131), .A2(n5129), .ZN(n5128) );
  INV_X1 U5425 ( .A(n5439), .ZN(n5129) );
  NAND2_X1 U5426 ( .A1(n5273), .A2(n6779), .ZN(n6636) );
  OR2_X1 U5427 ( .A1(n6781), .A2(n6622), .ZN(n5273) );
  NAND2_X1 U5428 ( .A1(n5341), .A2(n4975), .ZN(n4974) );
  NOR2_X1 U5429 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n5220) );
  NOR2_X1 U5430 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n5221) );
  INV_X1 U5431 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n6210) );
  AOI21_X1 U5432 ( .B1(n5053), .B2(n5055), .A(n5051), .ZN(n5050) );
  INV_X1 U5433 ( .A(n9512), .ZN(n5051) );
  OR2_X1 U5434 ( .A1(n4922), .A2(n4921), .ZN(n6058) );
  NAND2_X1 U5435 ( .A1(n6057), .A2(n8586), .ZN(n4921) );
  AOI21_X1 U5436 ( .B1(n4925), .B2(n4924), .A(n4923), .ZN(n4922) );
  NAND2_X1 U5437 ( .A1(n8532), .A2(n5012), .ZN(n5011) );
  NOR2_X1 U5438 ( .A1(n5264), .A2(n5122), .ZN(n5121) );
  INV_X1 U5439 ( .A(n5478), .ZN(n5122) );
  INV_X1 U5440 ( .A(n5265), .ZN(n5264) );
  INV_X1 U5441 ( .A(n4910), .ZN(n5263) );
  NAND2_X1 U5442 ( .A1(n5121), .A2(n5119), .ZN(n5118) );
  INV_X1 U5443 ( .A(n5950), .ZN(n5119) );
  INV_X1 U5444 ( .A(SI_17_), .ZN(n9700) );
  INV_X1 U5445 ( .A(SI_9_), .ZN(n9712) );
  INV_X1 U5446 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n5440) );
  INV_X1 U5447 ( .A(SI_8_), .ZN(n9586) );
  NAND2_X1 U5448 ( .A1(n6786), .A2(n6785), .ZN(n6788) );
  NAND2_X1 U5449 ( .A1(n5133), .A2(n4881), .ZN(n6786) );
  OAI21_X1 U5450 ( .B1(n9065), .B2(n6637), .A(n6776), .ZN(n6617) );
  INV_X1 U5451 ( .A(n6636), .ZN(n6816) );
  OR2_X1 U5452 ( .A1(n6498), .A2(n6243), .ZN(n6245) );
  OR2_X1 U5453 ( .A1(n6354), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n6388) );
  AND2_X1 U5454 ( .A1(n6776), .A2(n6777), .ZN(n6790) );
  AOI21_X1 U5455 ( .B1(n5331), .B2(n5333), .A(n9099), .ZN(n5330) );
  INV_X1 U5456 ( .A(n5334), .ZN(n5331) );
  INV_X1 U5457 ( .A(n5333), .ZN(n5332) );
  AND2_X1 U5458 ( .A1(n6743), .A2(n6742), .ZN(n6811) );
  NAND2_X1 U5459 ( .A1(n5089), .A2(n5091), .ZN(n5088) );
  OR2_X1 U5460 ( .A1(n6483), .A2(n9773), .ZN(n6496) );
  NAND2_X1 U5461 ( .A1(n5092), .A2(n6715), .ZN(n5091) );
  NAND2_X1 U5462 ( .A1(n8493), .A2(n6712), .ZN(n5092) );
  NAND2_X1 U5463 ( .A1(n6420), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6438) );
  INV_X1 U5464 ( .A(n6422), .ZN(n6420) );
  OR2_X1 U5465 ( .A1(n6406), .A2(n9667), .ZN(n6422) );
  OR2_X1 U5466 ( .A1(n6393), .A2(n6392), .ZN(n6406) );
  NOR2_X1 U5467 ( .A1(n7963), .A2(n7964), .ZN(n7967) );
  INV_X1 U5468 ( .A(n10432), .ZN(n5169) );
  NAND2_X1 U5469 ( .A1(n9155), .A2(n9055), .ZN(n9128) );
  NOR2_X1 U5470 ( .A1(n9128), .A2(n9301), .ZN(n8602) );
  AND2_X1 U5471 ( .A1(n8369), .A2(n4867), .ZN(n9264) );
  NOR2_X2 U5472 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n6239) );
  INV_X1 U5473 ( .A(n8629), .ZN(n5073) );
  INV_X1 U5474 ( .A(n5205), .ZN(n5202) );
  OR2_X1 U5475 ( .A1(n4850), .A2(n6139), .ZN(n5578) );
  INV_X1 U5476 ( .A(n7056), .ZN(n5179) );
  OR2_X1 U5477 ( .A1(n10102), .A2(n8681), .ZN(n7052) );
  NOR2_X1 U5478 ( .A1(n10102), .A2(n5006), .ZN(n5005) );
  INV_X1 U5479 ( .A(n5007), .ZN(n5006) );
  INV_X1 U5480 ( .A(n7046), .ZN(n5192) );
  INV_X1 U5481 ( .A(n10021), .ZN(n5193) );
  NOR2_X1 U5482 ( .A1(n10106), .A2(n10113), .ZN(n5007) );
  NOR2_X1 U5483 ( .A1(n8344), .A2(n5009), .ZN(n8557) );
  NAND2_X1 U5484 ( .A1(n9407), .A2(n5010), .ZN(n5009) );
  NOR2_X1 U5485 ( .A1(n5011), .A2(n10141), .ZN(n5010) );
  OR2_X1 U5486 ( .A1(n10141), .A2(n9562), .ZN(n7041) );
  OAI21_X1 U5487 ( .B1(n5373), .B2(n5372), .A(n7109), .ZN(n5371) );
  NAND2_X1 U5488 ( .A1(n8166), .A2(n7130), .ZN(n7375) );
  AND2_X1 U5489 ( .A1(n8343), .A2(n7107), .ZN(n5373) );
  AND2_X1 U5490 ( .A1(n7031), .A2(n8192), .ZN(n4972) );
  INV_X1 U5491 ( .A(n7030), .ZN(n5183) );
  INV_X1 U5492 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n5851) );
  NAND2_X1 U5493 ( .A1(n10480), .A2(n4866), .ZN(n5002) );
  AND2_X1 U5494 ( .A1(n10518), .A2(n10566), .ZN(n5001) );
  NAND2_X1 U5495 ( .A1(n8012), .A2(n8013), .ZN(n5356) );
  OR2_X1 U5496 ( .A1(n10401), .A2(n7997), .ZN(n7996) );
  INV_X1 U5497 ( .A(n7375), .ZN(n7663) );
  NAND2_X1 U5498 ( .A1(n9570), .A2(n10540), .ZN(n8818) );
  OR2_X1 U5499 ( .A1(n8298), .A2(n10163), .ZN(n8344) );
  NOR2_X1 U5500 ( .A1(n5002), .A2(n8276), .ZN(n8212) );
  INV_X1 U5501 ( .A(n5537), .ZN(n5280) );
  INV_X1 U5502 ( .A(n5279), .ZN(n5278) );
  OAI21_X1 U5503 ( .B1(n5583), .B2(n5280), .A(n5569), .ZN(n5279) );
  AND3_X1 U5504 ( .A1(n4998), .A2(n4999), .A3(n5374), .ZN(n5546) );
  INV_X1 U5505 ( .A(n5634), .ZN(n5283) );
  INV_X1 U5506 ( .A(n5513), .ZN(n5286) );
  INV_X1 U5507 ( .A(n5285), .ZN(n5284) );
  OAI21_X1 U5508 ( .B1(n5288), .B2(n4909), .A(n5518), .ZN(n5285) );
  INV_X1 U5509 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n6188) );
  OAI21_X1 U5510 ( .B1(n5677), .B2(n5499), .A(n5498), .ZN(n6025) );
  NAND2_X1 U5511 ( .A1(n5114), .A2(n5113), .ZN(n5933) );
  NAND2_X1 U5512 ( .A1(n4895), .A2(n5465), .ZN(n5113) );
  OAI21_X1 U5513 ( .B1(n5807), .B2(n4970), .A(n4968), .ZN(n4966) );
  INV_X1 U5514 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5754) );
  NAND2_X1 U5515 ( .A1(n4961), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n4960) );
  INV_X1 U5516 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4961) );
  INV_X1 U5517 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n5409) );
  XNOR2_X1 U5518 ( .A(n6958), .B(n6956), .ZN(n8836) );
  NAND2_X1 U5519 ( .A1(n6345), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n6357) );
  INV_X1 U5520 ( .A(n6346), .ZN(n6345) );
  OR2_X1 U5521 ( .A1(n6509), .A2(n9661), .ZN(n6517) );
  NAND2_X1 U5522 ( .A1(n6516), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n6524) );
  INV_X1 U5523 ( .A(n6517), .ZN(n6516) );
  XNOR2_X1 U5524 ( .A(n10434), .B(n6976), .ZN(n6872) );
  AND2_X1 U5525 ( .A1(n6869), .A2(n6870), .ZN(n7602) );
  AND2_X1 U5526 ( .A1(n6886), .A2(n6881), .ZN(n5150) );
  NAND2_X1 U5527 ( .A1(n8167), .A2(n6893), .ZN(n8176) );
  AND2_X1 U5528 ( .A1(n6953), .A2(n6947), .ZN(n5324) );
  AND2_X1 U5529 ( .A1(n7396), .A2(n6855), .ZN(n7482) );
  INV_X1 U5530 ( .A(n6925), .ZN(n4949) );
  INV_X1 U5531 ( .A(n8566), .ZN(n4945) );
  NAND2_X1 U5532 ( .A1(n6302), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6316) );
  INV_X1 U5533 ( .A(n6631), .ZN(n6632) );
  OR2_X1 U5534 ( .A1(n7435), .A2(n7009), .ZN(n6975) );
  AND2_X1 U5535 ( .A1(n6568), .A2(n6567), .ZN(n8829) );
  OR2_X1 U5536 ( .A1(n9108), .A2(n6574), .ZN(n6568) );
  NOR2_X1 U5537 ( .A1(n6273), .A2(n6224), .ZN(n6226) );
  NAND2_X1 U5538 ( .A1(n7152), .A2(n4995), .ZN(n10322) );
  NAND2_X1 U5539 ( .A1(n10319), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n4995) );
  OR2_X1 U5540 ( .A1(n7189), .A2(n7188), .ZN(n4982) );
  AND2_X1 U5541 ( .A1(n4980), .A2(n4979), .ZN(n8959) );
  NAND2_X1 U5542 ( .A1(n7940), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n4979) );
  NAND2_X1 U5543 ( .A1(n8959), .A2(n8960), .ZN(n8958) );
  NOR2_X1 U5544 ( .A1(n8025), .A2(n4988), .ZN(n8028) );
  AND2_X1 U5545 ( .A1(n8026), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n4988) );
  NAND2_X1 U5546 ( .A1(n8028), .A2(n8027), .ZN(n8121) );
  NAND2_X1 U5547 ( .A1(n8121), .A2(n4987), .ZN(n8123) );
  OR2_X1 U5548 ( .A1(n8122), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n4987) );
  NAND2_X1 U5549 ( .A1(n8123), .A2(n8124), .ZN(n8435) );
  AND2_X1 U5550 ( .A1(n9107), .A2(n4899), .ZN(n9038) );
  XNOR2_X1 U5551 ( .A(n9284), .B(n9069), .ZN(n9060) );
  AND2_X1 U5552 ( .A1(n9107), .A2(n5152), .ZN(n9073) );
  INV_X1 U5553 ( .A(n5154), .ZN(n5152) );
  INV_X1 U5554 ( .A(n9060), .ZN(n6594) );
  NAND2_X1 U5555 ( .A1(n9107), .A2(n9097), .ZN(n9092) );
  NAND2_X1 U5556 ( .A1(n5112), .A2(n5109), .ZN(n9113) );
  NOR2_X1 U5557 ( .A1(n9144), .A2(n5110), .ZN(n5109) );
  INV_X1 U5558 ( .A(n6551), .ZN(n5110) );
  OR2_X1 U5559 ( .A1(n6552), .A2(n9672), .ZN(n6561) );
  NAND2_X1 U5560 ( .A1(n5079), .A2(n5077), .ZN(n9123) );
  AOI21_X1 U5561 ( .B1(n5080), .B2(n5226), .A(n5078), .ZN(n5077) );
  INV_X1 U5562 ( .A(n6763), .ZN(n5078) );
  NOR2_X1 U5563 ( .A1(n9206), .A2(n5160), .ZN(n9169) );
  AND3_X1 U5564 ( .A1(n6528), .A2(n6527), .A3(n6526), .ZN(n9197) );
  AOI21_X1 U5565 ( .B1(n5214), .B2(n5216), .A(n5213), .ZN(n5212) );
  NOR2_X1 U5566 ( .A1(n9239), .A2(n9333), .ZN(n9230) );
  OR2_X1 U5567 ( .A1(n9241), .A2(n9336), .ZN(n9239) );
  AOI21_X1 U5568 ( .B1(n5339), .B2(n8541), .A(n5338), .ZN(n5337) );
  NAND2_X1 U5569 ( .A1(n6463), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n6483) );
  INV_X1 U5570 ( .A(n6464), .ZN(n6463) );
  OR2_X1 U5571 ( .A1(n9349), .A2(n8775), .ZN(n9257) );
  NAND2_X1 U5572 ( .A1(n6437), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6450) );
  INV_X1 U5573 ( .A(n6438), .ZN(n6437) );
  NOR2_X1 U5574 ( .A1(n10661), .A2(n8371), .ZN(n5165) );
  NAND2_X1 U5575 ( .A1(n8369), .A2(n5163), .ZN(n8542) );
  AND4_X1 U5576 ( .A1(n6445), .A2(n6444), .A3(n6443), .A4(n6442), .ZN(n8505)
         );
  NAND2_X1 U5577 ( .A1(n8369), .A2(n10654), .ZN(n8508) );
  NOR2_X1 U5578 ( .A1(n10607), .A2(n10640), .ZN(n8286) );
  AND2_X1 U5579 ( .A1(n8286), .A2(n10647), .ZN(n8369) );
  AOI21_X1 U5580 ( .B1(n5240), .B2(n8136), .A(n5239), .ZN(n5096) );
  INV_X1 U5581 ( .A(n6685), .ZN(n5239) );
  OR2_X1 U5582 ( .A1(n10605), .A2(n10606), .ZN(n10607) );
  NAND2_X1 U5583 ( .A1(n8137), .A2(n5240), .ZN(n10609) );
  AND2_X1 U5584 ( .A1(n8234), .A2(n8233), .ZN(n10602) );
  NAND2_X1 U5585 ( .A1(n8138), .A2(n5343), .ZN(n8137) );
  NOR2_X1 U5586 ( .A1(n5166), .A2(n10432), .ZN(n8142) );
  NAND2_X1 U5587 ( .A1(n5169), .A2(n5168), .ZN(n7981) );
  INV_X1 U5588 ( .A(n7963), .ZN(n6329) );
  NAND2_X1 U5589 ( .A1(n5169), .A2(n5167), .ZN(n7983) );
  INV_X1 U5590 ( .A(n5170), .ZN(n5167) );
  NOR2_X1 U5591 ( .A1(n10432), .A2(n10473), .ZN(n8053) );
  AND4_X1 U5592 ( .A1(n6322), .A2(n6321), .A3(n6320), .A4(n6319), .ZN(n8065)
         );
  AND2_X1 U5593 ( .A1(n6666), .A2(n6665), .ZN(n8058) );
  AND4_X1 U5594 ( .A1(n6295), .A2(n6294), .A3(n6293), .A4(n6292), .ZN(n10439)
         );
  NAND2_X1 U5595 ( .A1(n7729), .A2(n4859), .ZN(n10441) );
  NAND2_X1 U5596 ( .A1(n10438), .A2(n7738), .ZN(n6658) );
  OR2_X1 U5597 ( .A1(n10431), .A2(n10450), .ZN(n10432) );
  OR2_X1 U5598 ( .A1(n7734), .A2(n7738), .ZN(n10431) );
  NAND2_X1 U5599 ( .A1(n5250), .A2(n5249), .ZN(n5248) );
  INV_X1 U5600 ( .A(n7235), .ZN(n5249) );
  NAND2_X1 U5601 ( .A1(n6847), .A2(n7565), .ZN(n7685) );
  NAND2_X1 U5602 ( .A1(n6559), .A2(n6558), .ZN(n9295) );
  AND2_X1 U5603 ( .A1(n8377), .A2(n8375), .ZN(n5350) );
  INV_X1 U5604 ( .A(n6355), .ZN(n5095) );
  INV_X1 U5605 ( .A(n10673), .ZN(n10663) );
  NAND2_X1 U5606 ( .A1(n6459), .A2(n6214), .ZN(n6609) );
  NAND2_X1 U5607 ( .A1(n5157), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6490) );
  AND2_X1 U5608 ( .A1(n6458), .A2(n6478), .ZN(n5156) );
  AND2_X1 U5609 ( .A1(n5219), .A2(n4957), .ZN(n6459) );
  NOR2_X1 U5610 ( .A1(n5217), .A2(n6296), .ZN(n4957) );
  INV_X1 U5611 ( .A(n5222), .ZN(n5217) );
  OR2_X1 U5612 ( .A1(n6339), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n6354) );
  INV_X1 U5613 ( .A(n4868), .ZN(n5043) );
  AOI21_X1 U5614 ( .B1(n5045), .B2(n5048), .A(n4893), .ZN(n5044) );
  NAND2_X1 U5615 ( .A1(n7499), .A2(n7498), .ZN(n7505) );
  NAND2_X1 U5616 ( .A1(n7497), .A2(n7496), .ZN(n7498) );
  NOR2_X1 U5617 ( .A1(n9502), .A2(n5058), .ZN(n5057) );
  INV_X1 U5618 ( .A(n8650), .ZN(n5058) );
  OR2_X1 U5619 ( .A1(n8692), .A2(n8691), .ZN(n8693) );
  NAND2_X1 U5620 ( .A1(n8685), .A2(n8684), .ZN(n9481) );
  NAND2_X1 U5621 ( .A1(n9413), .A2(n9415), .ZN(n9482) );
  NAND2_X1 U5622 ( .A1(n8152), .A2(n8101), .ZN(n5034) );
  NAND2_X1 U5623 ( .A1(n5597), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n5690) );
  OR2_X1 U5624 ( .A1(n5690), .A2(n9435), .ZN(n6028) );
  OR2_X1 U5625 ( .A1(n6028), .A2(n9513), .ZN(n6030) );
  OR2_X1 U5626 ( .A1(n9431), .A2(n5056), .ZN(n5055) );
  INV_X1 U5627 ( .A(n9503), .ZN(n5056) );
  INV_X1 U5628 ( .A(n5054), .ZN(n5053) );
  OAI21_X1 U5629 ( .B1(n5057), .B2(n5055), .A(n9430), .ZN(n5054) );
  NAND2_X1 U5630 ( .A1(n8324), .A2(n8323), .ZN(n5243) );
  AND2_X1 U5631 ( .A1(n7645), .A2(n7646), .ZN(n9521) );
  NAND2_X1 U5632 ( .A1(n5582), .A2(n9882), .ZN(n6142) );
  AOI21_X1 U5633 ( .B1(n5392), .B2(n6091), .A(n7130), .ZN(n6144) );
  NOR2_X1 U5634 ( .A1(n6150), .A2(n6184), .ZN(n6091) );
  AND2_X1 U5635 ( .A1(n5657), .A2(n5656), .ZN(n9448) );
  AND4_X1 U5636 ( .A1(n5818), .A2(n5817), .A3(n5816), .A4(n5815), .ZN(n10490)
         );
  AND4_X1 U5637 ( .A1(n5751), .A2(n5750), .A3(n5749), .A4(n5748), .ZN(n7794)
         );
  AND3_X1 U5638 ( .A1(n5766), .A2(n5765), .A3(n5764), .ZN(n5767) );
  NAND4_X1 U5639 ( .A1(n5727), .A2(n5726), .A3(n5725), .A4(n5724), .ZN(n7380)
         );
  NOR2_X1 U5640 ( .A1(n6073), .A2(n6072), .ZN(n8813) );
  OAI22_X1 U5641 ( .A1(n9920), .A2(n5176), .B1(n8807), .B2(n5177), .ZN(n9897)
         );
  NAND2_X1 U5642 ( .A1(n8586), .A2(n6137), .ZN(n5176) );
  AND2_X1 U5643 ( .A1(n8808), .A2(n5178), .ZN(n5177) );
  NAND2_X1 U5644 ( .A1(n8586), .A2(n5179), .ZN(n5178) );
  NAND2_X1 U5645 ( .A1(n8585), .A2(n8586), .ZN(n8809) );
  AOI21_X1 U5646 ( .B1(n9929), .B2(n9928), .A(n4971), .ZN(n9922) );
  INV_X1 U5647 ( .A(n7054), .ZN(n4971) );
  NAND2_X1 U5648 ( .A1(n9922), .A2(n9921), .ZN(n9920) );
  AND2_X1 U5649 ( .A1(n6046), .A2(n6045), .ZN(n9917) );
  NAND2_X1 U5650 ( .A1(n9995), .A2(n5003), .ZN(n9941) );
  NOR2_X1 U5651 ( .A1(n10097), .A2(n5004), .ZN(n5003) );
  INV_X1 U5652 ( .A(n5005), .ZN(n5004) );
  NOR2_X1 U5653 ( .A1(n9941), .A2(n10092), .ZN(n9916) );
  NAND2_X1 U5654 ( .A1(n9933), .A2(n7125), .ZN(n9934) );
  NAND2_X1 U5655 ( .A1(n9995), .A2(n7062), .ZN(n9978) );
  NAND2_X1 U5656 ( .A1(n9995), .A2(n5007), .ZN(n9961) );
  INV_X1 U5657 ( .A(n5359), .ZN(n5358) );
  OAI22_X1 U5658 ( .A1(n9997), .A2(n5360), .B1(n7120), .B2(n9436), .ZN(n5359)
         );
  NOR2_X1 U5659 ( .A1(n10013), .A2(n10117), .ZN(n9995) );
  NAND2_X1 U5660 ( .A1(n8557), .A2(n7061), .ZN(n10057) );
  NAND2_X1 U5661 ( .A1(n5995), .A2(n5994), .ZN(n10043) );
  NAND2_X1 U5662 ( .A1(n5175), .A2(n4876), .ZN(n10034) );
  AND2_X1 U5663 ( .A1(n7043), .A2(n6095), .ZN(n10050) );
  OR2_X1 U5664 ( .A1(n8517), .A2(n8518), .ZN(n8520) );
  INV_X1 U5665 ( .A(n8419), .ZN(n5184) );
  NOR3_X1 U5666 ( .A1(n8344), .A2(n10152), .A3(n10157), .ZN(n8528) );
  NOR2_X1 U5667 ( .A1(n8344), .A2(n10157), .ZN(n8416) );
  NAND2_X1 U5668 ( .A1(n8296), .A2(n5373), .ZN(n8342) );
  INV_X1 U5669 ( .A(n8295), .ZN(n7106) );
  AND2_X1 U5670 ( .A1(n6103), .A2(n7033), .ZN(n8295) );
  NAND2_X1 U5671 ( .A1(n8186), .A2(n7030), .ZN(n8208) );
  NAND2_X1 U5672 ( .A1(n8187), .A2(n8192), .ZN(n8186) );
  OR2_X1 U5673 ( .A1(n5829), .A2(n5710), .ZN(n5852) );
  NAND2_X1 U5674 ( .A1(n10480), .A2(n5001), .ZN(n10536) );
  NOR2_X1 U5675 ( .A1(n7996), .A2(n7929), .ZN(n10480) );
  NAND2_X1 U5676 ( .A1(n10480), .A2(n10518), .ZN(n10535) );
  AND4_X1 U5677 ( .A1(n5802), .A2(n5801), .A3(n5800), .A4(n5799), .ZN(n8011)
         );
  NAND2_X1 U5678 ( .A1(n7024), .A2(n7023), .ZN(n10543) );
  INV_X1 U5679 ( .A(n8013), .ZN(n7023) );
  NAND2_X1 U5680 ( .A1(n6159), .A2(n6076), .ZN(n10406) );
  AND4_X1 U5681 ( .A1(n5788), .A2(n5787), .A3(n5786), .A4(n5785), .ZN(n10491)
         );
  INV_X1 U5682 ( .A(n5777), .ZN(n10403) );
  INV_X1 U5683 ( .A(n10489), .ZN(n10539) );
  NAND2_X1 U5684 ( .A1(n5637), .A2(n5636), .ZN(n10086) );
  AND2_X1 U5685 ( .A1(n10019), .A2(n7045), .ZN(n9999) );
  OR2_X1 U5686 ( .A1(n7627), .A2(n7063), .ZN(n10582) );
  INV_X1 U5687 ( .A(n10365), .ZN(n10581) );
  NOR2_X1 U5688 ( .A1(n7410), .A2(n7409), .ZN(n7418) );
  XNOR2_X1 U5689 ( .A(n5584), .B(n5583), .ZN(n8824) );
  AND2_X1 U5690 ( .A1(n5527), .A2(n5526), .ZN(n5622) );
  XNOR2_X1 U5691 ( .A(n5635), .B(n5634), .ZN(n8579) );
  OAI21_X1 U5692 ( .B1(n5661), .B2(n4909), .A(n5284), .ZN(n5635) );
  NAND2_X1 U5693 ( .A1(n5287), .A2(n5513), .ZN(n6040) );
  NAND2_X1 U5694 ( .A1(n5661), .A2(n5288), .ZN(n5287) );
  NAND2_X1 U5695 ( .A1(n5380), .A2(n5188), .ZN(n5187) );
  AND2_X1 U5696 ( .A1(n5538), .A2(n6188), .ZN(n5375) );
  NAND2_X1 U5697 ( .A1(n5106), .A2(n5503), .ZN(n5658) );
  NAND2_X1 U5698 ( .A1(n5108), .A2(n5107), .ZN(n5106) );
  INV_X1 U5699 ( .A(n6024), .ZN(n5107) );
  INV_X1 U5700 ( .A(n6025), .ZN(n5108) );
  NAND2_X1 U5701 ( .A1(n5969), .A2(n4910), .ZN(n5261) );
  OR2_X1 U5702 ( .A1(n5952), .A2(P1_IR_REG_15__SCAN_IN), .ZN(n5953) );
  AND2_X1 U5703 ( .A1(n5915), .A2(n5952), .ZN(n9798) );
  NAND2_X1 U5704 ( .A1(n5894), .A2(n5462), .ZN(n5908) );
  NAND2_X1 U5705 ( .A1(n5291), .A2(n5455), .ZN(n5874) );
  INV_X1 U5706 ( .A(n5290), .ZN(n5291) );
  OAI21_X1 U5707 ( .B1(n5445), .B2(n5271), .A(n5268), .ZN(n5859) );
  OR3_X1 U5708 ( .A1(n5844), .A2(P1_IR_REG_8__SCAN_IN), .A3(
        P1_IR_REG_9__SCAN_IN), .ZN(n5846) );
  NOR2_X1 U5709 ( .A1(n5846), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n5876) );
  AND2_X1 U5710 ( .A1(n5803), .A2(n5704), .ZN(n5819) );
  AOI21_X1 U5711 ( .B1(n5424), .B2(n5099), .A(n4882), .ZN(n5097) );
  NAND2_X1 U5712 ( .A1(n5773), .A2(n4864), .ZN(n4958) );
  INV_X1 U5713 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5790) );
  NAND2_X1 U5714 ( .A1(n5260), .A2(n5423), .ZN(n5757) );
  NAND2_X1 U5715 ( .A1(n5773), .A2(n5772), .ZN(n5260) );
  NAND2_X1 U5716 ( .A1(n5721), .A2(n5720), .ZN(n5116) );
  NOR2_X2 U5717 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5741) );
  NOR2_X1 U5718 ( .A1(n10228), .A2(n8739), .ZN(n8740) );
  AND4_X1 U5719 ( .A1(n6338), .A2(n6337), .A3(n6336), .A4(n6335), .ZN(n8175)
         );
  NAND2_X1 U5720 ( .A1(n5141), .A2(n5140), .ZN(n8828) );
  AOI21_X1 U5721 ( .B1(n4862), .B2(n4950), .A(n4913), .ZN(n5140) );
  NAND2_X1 U5722 ( .A1(n6570), .A2(n6569), .ZN(n9289) );
  OR2_X1 U5723 ( .A1(n8871), .A2(n10613), .ZN(n8913) );
  INV_X1 U5724 ( .A(n5300), .ZN(n5299) );
  OAI211_X1 U5725 ( .C1(n5302), .C2(n5308), .A(n5301), .B(n7004), .ZN(n5300)
         );
  NAND2_X1 U5726 ( .A1(n5307), .A2(n5306), .ZN(n5301) );
  NAND2_X1 U5727 ( .A1(n6515), .A2(n6514), .ZN(n9321) );
  AND4_X1 U5728 ( .A1(n6383), .A2(n6382), .A3(n6381), .A4(n6380), .ZN(n10614)
         );
  NAND2_X1 U5729 ( .A1(n6921), .A2(n8456), .ZN(n8461) );
  NAND2_X1 U5730 ( .A1(n8461), .A2(n6925), .ZN(n8568) );
  OR2_X1 U5731 ( .A1(n7685), .A2(n7701), .ZN(n7396) );
  NAND2_X1 U5732 ( .A1(n6506), .A2(n6505), .ZN(n9326) );
  AND4_X1 U5733 ( .A1(n6400), .A2(n6399), .A3(n6398), .A4(n6397), .ZN(n8374)
         );
  NAND2_X1 U5734 ( .A1(n5318), .A2(n5320), .ZN(n8312) );
  OR2_X1 U5735 ( .A1(n8400), .A2(n4857), .ZN(n5318) );
  NAND2_X1 U5736 ( .A1(n8400), .A2(n6908), .ZN(n8408) );
  NAND2_X1 U5737 ( .A1(n5325), .A2(n6947), .ZN(n8894) );
  NAND2_X1 U5738 ( .A1(n5149), .A2(n8245), .ZN(n8400) );
  AND2_X1 U5739 ( .A1(n6865), .A2(n6864), .ZN(n7558) );
  NAND2_X1 U5740 ( .A1(n5296), .A2(n7481), .ZN(n7604) );
  AND2_X1 U5741 ( .A1(n7558), .A2(n6859), .ZN(n5296) );
  AND2_X1 U5742 ( .A1(n7007), .A2(n7002), .ZN(n8905) );
  OAI21_X1 U5743 ( .B1(n6921), .B2(n4947), .A(n4944), .ZN(n8907) );
  INV_X1 U5744 ( .A(n4948), .ZN(n4947) );
  AOI21_X1 U5745 ( .B1(n4948), .B2(n4946), .A(n4945), .ZN(n4944) );
  NOR2_X1 U5746 ( .A1(n8565), .A2(n4949), .ZN(n4948) );
  AOI21_X1 U5747 ( .B1(n5315), .B2(n5317), .A(n4918), .ZN(n5313) );
  AND2_X1 U5748 ( .A1(n6996), .A2(n10446), .ZN(n8922) );
  AND2_X1 U5749 ( .A1(n7397), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8910) );
  NAND2_X1 U5750 ( .A1(n7781), .A2(n6874), .ZN(n5314) );
  OAI21_X1 U5751 ( .B1(n4953), .B2(n5143), .A(n4952), .ZN(n8920) );
  AOI21_X1 U5752 ( .B1(n4951), .B2(n8865), .A(n4950), .ZN(n4952) );
  OAI211_X1 U5753 ( .C1(n5149), .C2(n5148), .A(n5319), .B(n5146), .ZN(n6913)
         );
  NAND2_X1 U5754 ( .A1(n5320), .A2(n5147), .ZN(n5146) );
  AOI21_X1 U5755 ( .B1(n5320), .B2(n4857), .A(n4871), .ZN(n5319) );
  XNOR2_X1 U5756 ( .A(n6827), .B(P2_IR_REG_22__SCAN_IN), .ZN(n6848) );
  AND2_X1 U5757 ( .A1(n6580), .A2(n6579), .ZN(n9059) );
  INV_X1 U5758 ( .A(n8829), .ZN(n9101) );
  INV_X1 U5759 ( .A(n10612), .ZN(n8939) );
  INV_X1 U5760 ( .A(n8175), .ZN(n8135) );
  INV_X1 U5761 ( .A(n10439), .ZN(n8942) );
  OR2_X1 U5762 ( .A1(n6273), .A2(n6274), .ZN(n6275) );
  INV_X1 U5763 ( .A(n10438), .ZN(n8944) );
  NAND2_X1 U5764 ( .A1(n7477), .A2(n7478), .ZN(n7476) );
  NOR2_X1 U5765 ( .A1(n7217), .A2(n7216), .ZN(n7215) );
  AND2_X1 U5766 ( .A1(n7476), .A2(n4997), .ZN(n7217) );
  NAND2_X1 U5767 ( .A1(n7475), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n4997) );
  NOR2_X1 U5768 ( .A1(n7186), .A2(n4983), .ZN(n7189) );
  AND2_X1 U5769 ( .A1(n7191), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n4983) );
  INV_X1 U5770 ( .A(n4982), .ZN(n7200) );
  NOR2_X1 U5771 ( .A1(n7203), .A2(n7202), .ZN(n7518) );
  AND2_X1 U5772 ( .A1(n4982), .A2(n4981), .ZN(n7203) );
  NAND2_X1 U5773 ( .A1(n7205), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n4981) );
  NAND2_X1 U5774 ( .A1(n8958), .A2(n4978), .ZN(n7944) );
  OR2_X1 U5775 ( .A1(n8963), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n4978) );
  NAND2_X1 U5776 ( .A1(n4993), .A2(n4992), .ZN(n9005) );
  NAND2_X1 U5777 ( .A1(n9004), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n4992) );
  NOR2_X1 U5778 ( .A1(n9005), .A2(n9006), .ZN(n9020) );
  NAND2_X1 U5779 ( .A1(n5329), .A2(n5333), .ZN(n9091) );
  NAND2_X1 U5780 ( .A1(n9121), .A2(n5334), .ZN(n5329) );
  AOI21_X1 U5781 ( .B1(n9121), .B2(n9057), .A(n4858), .ZN(n9106) );
  NAND2_X1 U5782 ( .A1(n5082), .A2(n5080), .ZN(n9146) );
  NAND2_X1 U5783 ( .A1(n9164), .A2(n9053), .ZN(n9137) );
  AND2_X1 U5784 ( .A1(n9181), .A2(n9180), .ZN(n9319) );
  NAND2_X1 U5785 ( .A1(n9204), .A2(n5384), .ZN(n9187) );
  OAI21_X1 U5786 ( .B1(n9245), .B2(n5216), .A(n5214), .ZN(n9227) );
  NAND2_X1 U5787 ( .A1(n5340), .A2(n5339), .ZN(n9262) );
  OAI21_X1 U5788 ( .B1(n8503), .B2(n8493), .A(n6712), .ZN(n8496) );
  AND2_X1 U5789 ( .A1(n8376), .A2(n8375), .ZN(n8378) );
  AND2_X1 U5790 ( .A1(n8282), .A2(n8281), .ZN(n8285) );
  INV_X1 U5791 ( .A(n7970), .ZN(n4977) );
  INV_X1 U5792 ( .A(n10525), .ZN(n7985) );
  NAND2_X1 U5793 ( .A1(n5345), .A2(n7862), .ZN(n10430) );
  NAND2_X1 U5794 ( .A1(n7177), .A2(n10319), .ZN(n5139) );
  NAND2_X1 U5795 ( .A1(n4852), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5138) );
  OR2_X1 U5796 ( .A1(n9157), .A2(n7851), .ZN(n9255) );
  AND2_X2 U5797 ( .A1(n7445), .A2(n7444), .ZN(n10681) );
  INV_X1 U5798 ( .A(n9282), .ZN(n5094) );
  OR3_X1 U5799 ( .A1(n9315), .A2(n9314), .A3(n9313), .ZN(n9361) );
  AND2_X1 U5800 ( .A1(n7010), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10312) );
  NAND2_X1 U5801 ( .A1(n10214), .A2(n10213), .ZN(n10309) );
  NAND2_X1 U5802 ( .A1(n5258), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6235) );
  NAND2_X1 U5803 ( .A1(n6631), .A2(n5346), .ZN(n5258) );
  INV_X1 U5804 ( .A(n6848), .ZN(n8307) );
  NAND2_X1 U5805 ( .A1(n6627), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6629) );
  INV_X1 U5806 ( .A(n6624), .ZN(n9029) );
  INV_X1 U5807 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n7258) );
  INV_X1 U5808 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n7254) );
  AND4_X1 U5809 ( .A1(n5833), .A2(n5832), .A3(n5831), .A4(n5830), .ZN(n8098)
         );
  OAI21_X1 U5810 ( .B1(n7925), .B2(n7922), .A(n7921), .ZN(n8092) );
  AND2_X1 U5811 ( .A1(n5621), .A2(n5620), .ZN(n9396) );
  NAND2_X1 U5812 ( .A1(n8610), .A2(n5203), .ZN(n9401) );
  AOI22_X1 U5813 ( .A1(n5062), .A2(n5064), .B1(n5065), .B2(n5068), .ZN(n5060)
         );
  NAND2_X1 U5814 ( .A1(n5070), .A2(n5069), .ZN(n5068) );
  AND2_X1 U5815 ( .A1(n5609), .A2(n5608), .ZN(n9899) );
  OAI21_X1 U5816 ( .B1(n5044), .B2(n4868), .A(n5040), .ZN(n5039) );
  NAND2_X1 U5817 ( .A1(n5044), .A2(n5041), .ZN(n5040) );
  NAND2_X1 U5818 ( .A1(n5046), .A2(n5043), .ZN(n5041) );
  NAND2_X1 U5819 ( .A1(n5044), .A2(n5043), .ZN(n5042) );
  NAND2_X1 U5820 ( .A1(n5052), .A2(n9503), .ZN(n9434) );
  NAND2_X1 U5821 ( .A1(n9422), .A2(n5057), .ZN(n5052) );
  AND4_X1 U5822 ( .A1(n5870), .A2(n5869), .A3(n5868), .A4(n5867), .ZN(n8363)
         );
  NAND2_X1 U5823 ( .A1(n9479), .A2(n8693), .ZN(n9446) );
  AND4_X1 U5824 ( .A1(n6003), .A2(n6002), .A3(n6001), .A4(n6000), .ZN(n9474)
         );
  NAND2_X1 U5825 ( .A1(n5075), .A2(n5076), .ZN(n5074) );
  INV_X1 U5826 ( .A(n9455), .ZN(n5075) );
  AND4_X1 U5827 ( .A1(n5857), .A2(n5856), .A3(n5855), .A4(n5854), .ZN(n8267)
         );
  NAND2_X1 U5828 ( .A1(n8153), .A2(n8152), .ZN(n5252) );
  NAND2_X1 U5829 ( .A1(n9422), .A2(n8650), .ZN(n9505) );
  OAI21_X1 U5830 ( .B1(n9422), .B2(n5055), .A(n5053), .ZN(n9511) );
  AND4_X1 U5831 ( .A1(n5888), .A2(n5887), .A3(n5886), .A4(n5885), .ZN(n8486)
         );
  AND2_X1 U5832 ( .A1(n5243), .A2(n5244), .ZN(n8330) );
  INV_X1 U5833 ( .A(n4936), .ZN(n4935) );
  NAND2_X1 U5834 ( .A1(n4848), .A2(n5174), .ZN(n5173) );
  OAI21_X1 U5835 ( .B1(n5771), .B2(n5746), .A(n5171), .ZN(n4936) );
  NAND2_X1 U5836 ( .A1(n5061), .A2(n5070), .ZN(n9530) );
  NAND2_X1 U5837 ( .A1(n9455), .A2(n5071), .ZN(n5061) );
  NOR2_X1 U5838 ( .A1(n5232), .A2(n5234), .ZN(n5229) );
  NAND2_X1 U5839 ( .A1(n8685), .A2(n5233), .ZN(n5231) );
  INV_X1 U5840 ( .A(n9566), .ZN(n9536) );
  OR2_X1 U5841 ( .A1(n7514), .A2(n7386), .ZN(n9566) );
  OR2_X1 U5842 ( .A1(n7514), .A2(n7393), .ZN(n9561) );
  NAND2_X1 U5843 ( .A1(n5940), .A2(n5939), .ZN(n10146) );
  NAND2_X1 U5844 ( .A1(n7374), .A2(n10005), .ZN(n9564) );
  INV_X1 U5845 ( .A(n9396), .ZN(n9570) );
  OR2_X1 U5846 ( .A1(n8596), .A2(n6035), .ZN(n5646) );
  INV_X1 U5847 ( .A(n9543), .ZN(n9930) );
  INV_X1 U5848 ( .A(n9448), .ZN(n9954) );
  INV_X1 U5849 ( .A(n10000), .ZN(n9970) );
  INV_X1 U5850 ( .A(n7794), .ZN(n7364) );
  NAND2_X1 U5851 ( .A1(n5554), .A2(n5553), .ZN(n10067) );
  NAND2_X1 U5852 ( .A1(n5615), .A2(n5614), .ZN(n10076) );
  INV_X1 U5853 ( .A(n10086), .ZN(n9549) );
  NAND2_X1 U5854 ( .A1(n8590), .A2(n8589), .ZN(n8591) );
  INV_X1 U5855 ( .A(n10090), .ZN(n8592) );
  NAND2_X1 U5856 ( .A1(n7124), .A2(n7123), .ZN(n9946) );
  NAND2_X1 U5857 ( .A1(n10019), .A2(n5195), .ZN(n9982) );
  NAND2_X1 U5858 ( .A1(n5376), .A2(n5377), .ZN(n8191) );
  INV_X1 U5859 ( .A(n10364), .ZN(n7676) );
  NAND2_X1 U5860 ( .A1(n5019), .A2(n5745), .ZN(n5022) );
  OAI21_X1 U5861 ( .B1(n7237), .B2(n5021), .A(n5020), .ZN(n5019) );
  INV_X1 U5862 ( .A(n10046), .ZN(n10558) );
  INV_X1 U5863 ( .A(n5014), .ZN(n5013) );
  OAI21_X1 U5864 ( .B1(n10074), .B2(n10460), .A(n5015), .ZN(n5014) );
  NAND2_X1 U5865 ( .A1(n10072), .A2(n10365), .ZN(n5015) );
  NAND2_X1 U5866 ( .A1(n10084), .A2(n4962), .ZN(n10177) );
  INV_X1 U5867 ( .A(n4963), .ZN(n4962) );
  OAI21_X1 U5868 ( .B1(n10085), .B2(n10460), .A(n10083), .ZN(n4963) );
  AND2_X2 U5869 ( .A1(n7418), .A2(n7417), .ZN(n10594) );
  NAND2_X1 U5870 ( .A1(n7249), .A2(n7403), .ZN(n10211) );
  XNOR2_X1 U5871 ( .A(n5576), .B(n5575), .ZN(n9369) );
  NAND2_X1 U5872 ( .A1(n5276), .A2(n5275), .ZN(n5576) );
  NAND2_X1 U5873 ( .A1(n5560), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5561) );
  NAND2_X1 U5874 ( .A1(n5558), .A2(n5557), .ZN(n5559) );
  NAND2_X1 U5875 ( .A1(n5556), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5557) );
  NAND2_X1 U5876 ( .A1(n6200), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6202) );
  XNOR2_X1 U5877 ( .A(n5407), .B(n5406), .ZN(n8311) );
  INV_X1 U5878 ( .A(n7130), .ZN(n8185) );
  INV_X1 U5879 ( .A(n7063), .ZN(n8166) );
  INV_X1 U5880 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n7819) );
  AND2_X1 U5881 ( .A1(n5880), .A2(n5896), .ZN(n7836) );
  NAND2_X1 U5882 ( .A1(n4967), .A2(n5431), .ZN(n5823) );
  NAND2_X1 U5883 ( .A1(n5807), .A2(n5429), .ZN(n4967) );
  NOR2_X1 U5884 ( .A1(n8764), .A2(n8763), .ZN(n10246) );
  NOR2_X1 U5885 ( .A1(n10244), .A2(n10243), .ZN(n8763) );
  INV_X1 U5886 ( .A(n4980), .ZN(n7939) );
  INV_X1 U5887 ( .A(n4993), .ZN(n9003) );
  OAI21_X1 U5888 ( .B1(n6194), .B2(n6193), .A(n6192), .ZN(n6209) );
  INV_X1 U5889 ( .A(n5016), .ZN(n10071) );
  OAI21_X1 U5890 ( .B1(n10085), .B2(n10028), .A(n7135), .ZN(n7136) );
  INV_X1 U5891 ( .A(n5418), .ZN(n5021) );
  INV_X1 U5892 ( .A(n5070), .ZN(n5064) );
  AND3_X1 U5893 ( .A1(n5388), .A2(n4865), .A3(n5347), .ZN(n4855) );
  INV_X1 U5894 ( .A(n8630), .ZN(n5076) );
  INV_X4 U5895 ( .A(n6328), .ZN(n5250) );
  INV_X1 U5896 ( .A(n9997), .ZN(n5197) );
  OR2_X1 U5897 ( .A1(n5237), .A2(n9442), .ZN(n4856) );
  AND2_X1 U5898 ( .A1(n8317), .A2(n6910), .ZN(n4857) );
  OR2_X1 U5899 ( .A1(n10082), .A2(n9898), .ZN(n6137) );
  INV_X1 U5900 ( .A(n7460), .ZN(n5172) );
  NOR2_X1 U5901 ( .A1(n5111), .A2(n9301), .ZN(n4858) );
  AND4_X1 U5902 ( .A1(n6247), .A2(n6246), .A3(n6245), .A4(n6244), .ZN(n7485)
         );
  AND2_X1 U5903 ( .A1(n6285), .A2(n6658), .ZN(n4859) );
  INV_X1 U5904 ( .A(n9144), .ZN(n5111) );
  AND2_X1 U5905 ( .A1(n5268), .A2(n5860), .ZN(n4860) );
  NAND2_X1 U5906 ( .A1(n6762), .A2(n6782), .ZN(n4861) );
  AND2_X1 U5907 ( .A1(n5142), .A2(n8919), .ZN(n4862) );
  OAI21_X1 U5908 ( .B1(n7127), .B2(n5369), .A(n5367), .ZN(n8793) );
  OAI21_X1 U5909 ( .B1(n5083), .B2(n4898), .A(n6791), .ZN(n9098) );
  OR2_X1 U5910 ( .A1(n5483), .A2(n9677), .ZN(n4863) );
  AND2_X1 U5911 ( .A1(n5772), .A2(n5424), .ZN(n4864) );
  INV_X1 U5912 ( .A(n8864), .ZN(n4950) );
  AND2_X1 U5913 ( .A1(n6216), .A2(n5348), .ZN(n4865) );
  AND2_X1 U5914 ( .A1(n6751), .A2(n6750), .ZN(n9174) );
  INV_X1 U5915 ( .A(n9174), .ZN(n5225) );
  AND2_X1 U5916 ( .A1(n6102), .A2(n7032), .ZN(n7031) );
  INV_X1 U5917 ( .A(n7031), .ZN(n8207) );
  AND2_X1 U5918 ( .A1(n5001), .A2(n5000), .ZN(n4866) );
  OR2_X1 U5919 ( .A1(n9421), .A2(n9424), .ZN(n9422) );
  OR2_X1 U5920 ( .A1(n9289), .A2(n9059), .ZN(n6768) );
  INV_X1 U5921 ( .A(n5090), .ZN(n5089) );
  OAI21_X1 U5922 ( .B1(n5091), .B2(n6712), .A(n6716), .ZN(n5090) );
  AND2_X1 U5923 ( .A1(n5163), .A2(n5162), .ZN(n4867) );
  NAND2_X1 U5924 ( .A1(n8154), .A2(n5252), .ZN(n8155) );
  NAND2_X1 U5925 ( .A1(n6597), .A2(n6596), .ZN(n9280) );
  NAND2_X1 U5926 ( .A1(n6436), .A2(n6435), .ZN(n8781) );
  INV_X1 U5927 ( .A(n8781), .ZN(n5164) );
  INV_X1 U5928 ( .A(n7775), .ZN(n5317) );
  NAND2_X2 U5929 ( .A1(n6227), .A2(n6228), .ZN(n6273) );
  XOR2_X1 U5930 ( .A(n8723), .B(n8722), .Z(n4868) );
  AND2_X1 U5931 ( .A1(n6109), .A2(n7039), .ZN(n8518) );
  NAND3_X1 U5932 ( .A1(n6239), .A2(n5326), .A3(n6211), .ZN(n6296) );
  NAND2_X1 U5933 ( .A1(n9245), .A2(n9237), .ZN(n9223) );
  INV_X1 U5934 ( .A(n5760), .ZN(n5692) );
  INV_X1 U5935 ( .A(n5072), .ZN(n5071) );
  OR2_X1 U5936 ( .A1(n8635), .A2(n5073), .ZN(n5072) );
  AND2_X1 U5937 ( .A1(n10123), .A2(n9572), .ZN(n4869) );
  XNOR2_X1 U5938 ( .A(n5561), .B(n10195), .ZN(n5562) );
  INV_X1 U5939 ( .A(n5579), .ZN(n9882) );
  AOI21_X1 U5940 ( .B1(n9369), .B2(n6041), .A(n5577), .ZN(n5579) );
  NAND2_X1 U5941 ( .A1(n10102), .A2(n9969), .ZN(n4870) );
  XNOR2_X1 U5942 ( .A(n5613), .B(n5612), .ZN(n6582) );
  INV_X1 U5943 ( .A(n6802), .ZN(n4975) );
  NAND2_X1 U5944 ( .A1(n5439), .A2(n5438), .ZN(n5834) );
  INV_X1 U5945 ( .A(n8865), .ZN(n5143) );
  INV_X1 U5946 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n6826) );
  INV_X1 U5947 ( .A(n6842), .ZN(n8203) );
  XNOR2_X1 U5948 ( .A(n6611), .B(P2_IR_REG_21__SCAN_IN), .ZN(n6842) );
  AND2_X1 U5949 ( .A1(n8391), .A2(n6912), .ZN(n4871) );
  NAND2_X1 U5950 ( .A1(n7172), .A2(n5021), .ZN(n6328) );
  AND4_X1 U5951 ( .A1(n5222), .A2(n6239), .A3(n5326), .A4(n5218), .ZN(n4872)
         );
  AND3_X1 U5952 ( .A1(n6067), .A2(n5385), .A3(n6066), .ZN(n4873) );
  OR2_X1 U5953 ( .A1(n9054), .A2(n6782), .ZN(n4874) );
  AND2_X1 U5954 ( .A1(n6198), .A2(n6201), .ZN(n4875) );
  NAND2_X1 U5955 ( .A1(n6604), .A2(n6603), .ZN(n9039) );
  INV_X1 U5956 ( .A(n9039), .ZN(n5151) );
  XNOR2_X1 U5957 ( .A(n5425), .B(n4984), .ZN(n5424) );
  NAND2_X1 U5958 ( .A1(n5175), .A2(n7043), .ZN(n10031) );
  NAND2_X1 U5959 ( .A1(n5539), .A2(n5375), .ZN(n6196) );
  NAND2_X1 U5960 ( .A1(n5326), .A2(n6239), .ZN(n6280) );
  NAND2_X1 U5961 ( .A1(n5650), .A2(n5649), .ZN(n10097) );
  INV_X1 U5962 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n9370) );
  AND2_X1 U5963 ( .A1(n6133), .A2(n7056), .ZN(n9921) );
  NAND2_X1 U5964 ( .A1(n6405), .A2(n6404), .ZN(n8371) );
  NAND2_X1 U5965 ( .A1(n5679), .A2(n5678), .ZN(n10113) );
  AND2_X1 U5966 ( .A1(n10030), .A2(n7043), .ZN(n4876) );
  NAND2_X1 U5967 ( .A1(n9159), .A2(n9143), .ZN(n6755) );
  INV_X1 U5968 ( .A(n6755), .ZN(n5224) );
  XNOR2_X1 U5969 ( .A(n5451), .B(n5450), .ZN(n5860) );
  AND2_X1 U5970 ( .A1(n8827), .A2(n5310), .ZN(n5309) );
  INV_X1 U5971 ( .A(n5309), .ZN(n5306) );
  AND2_X1 U5972 ( .A1(n5352), .A2(n8556), .ZN(n4877) );
  NAND2_X1 U5973 ( .A1(n5112), .A2(n6551), .ZN(n9301) );
  AND2_X1 U5974 ( .A1(n9141), .A2(n9053), .ZN(n4878) );
  AND2_X1 U5975 ( .A1(n7103), .A2(n5377), .ZN(n4879) );
  AND2_X1 U5976 ( .A1(n9097), .A2(n9059), .ZN(n4880) );
  AND2_X1 U5977 ( .A1(n7025), .A2(n8076), .ZN(n10544) );
  AND2_X1 U5978 ( .A1(n5274), .A2(n5272), .ZN(n4881) );
  AND2_X1 U5979 ( .A1(n5425), .A2(SI_4_), .ZN(n4882) );
  NAND2_X1 U5980 ( .A1(n6649), .A2(n6258), .ZN(n7725) );
  NAND2_X1 U5981 ( .A1(n6763), .A2(n4874), .ZN(n4883) );
  AND2_X1 U5982 ( .A1(n5251), .A2(n5034), .ZN(n4884) );
  OR2_X1 U5983 ( .A1(n9333), .A2(n9248), .ZN(n6731) );
  INV_X1 U5984 ( .A(n6731), .ZN(n5213) );
  OR2_X1 U5985 ( .A1(n9343), .A2(n8933), .ZN(n9046) );
  INV_X1 U5986 ( .A(n9046), .ZN(n5338) );
  NAND2_X1 U5987 ( .A1(n6584), .A2(n6583), .ZN(n9284) );
  INV_X1 U5988 ( .A(n9284), .ZN(n5155) );
  AND2_X1 U5989 ( .A1(n6974), .A2(n6973), .ZN(n4885) );
  AND2_X1 U5990 ( .A1(n5451), .A2(SI_11_), .ZN(n4886) );
  NOR2_X1 U5991 ( .A1(n9471), .A2(n9470), .ZN(n4887) );
  NOR2_X1 U5992 ( .A1(n9295), .A2(n9101), .ZN(n4888) );
  NOR2_X1 U5993 ( .A1(n10082), .A2(n9571), .ZN(n4889) );
  NOR2_X1 U5994 ( .A1(n5190), .A2(n5187), .ZN(n5539) );
  AND2_X1 U5995 ( .A1(n5261), .A2(n5265), .ZN(n4890) );
  AOI21_X1 U5996 ( .B1(n5309), .B2(n4913), .A(n4885), .ZN(n5308) );
  NAND2_X1 U5997 ( .A1(n5455), .A2(n5454), .ZN(n4891) );
  OR2_X1 U5998 ( .A1(n10086), .A2(n9923), .ZN(n4892) );
  NAND2_X1 U5999 ( .A1(n4892), .A2(n7128), .ZN(n5369) );
  INV_X1 U6000 ( .A(n5241), .ZN(n5240) );
  NAND2_X1 U6001 ( .A1(n10610), .A2(n6680), .ZN(n5241) );
  INV_X1 U6002 ( .A(n9058), .ZN(n9099) );
  NAND2_X1 U6003 ( .A1(n6768), .A2(n6769), .ZN(n9058) );
  AND2_X1 U6004 ( .A1(n6134), .A2(n7057), .ZN(n8586) );
  AND2_X1 U6005 ( .A1(n6645), .A2(n6644), .ZN(n9188) );
  AND2_X1 U6006 ( .A1(n8716), .A2(n9389), .ZN(n4893) );
  INV_X1 U6007 ( .A(n5046), .ZN(n5045) );
  NAND2_X1 U6008 ( .A1(n5047), .A2(n8717), .ZN(n5046) );
  NAND2_X1 U6009 ( .A1(n5484), .A2(n5266), .ZN(n4894) );
  OR2_X1 U6010 ( .A1(n5466), .A2(n5115), .ZN(n4895) );
  NAND2_X1 U6011 ( .A1(n4958), .A2(n5097), .ZN(n5792) );
  NAND2_X1 U6012 ( .A1(n9349), .A2(n9043), .ZN(n4896) );
  NAND2_X1 U6013 ( .A1(n5741), .A2(n5210), .ZN(n5702) );
  AND3_X1 U6014 ( .A1(n5221), .A2(n5220), .A3(n6210), .ZN(n4897) );
  AND2_X1 U6015 ( .A1(n6137), .A2(n6136), .ZN(n8792) );
  INV_X1 U6016 ( .A(n8792), .ZN(n5366) );
  NAND2_X1 U6017 ( .A1(n6792), .A2(n9113), .ZN(n4898) );
  AND2_X1 U6018 ( .A1(n5153), .A2(n5151), .ZN(n4899) );
  AND2_X1 U6019 ( .A1(n5184), .A2(n7035), .ZN(n4900) );
  AND2_X1 U6020 ( .A1(n7865), .A2(n7962), .ZN(n4901) );
  AND2_X1 U6021 ( .A1(n5461), .A2(n5465), .ZN(n4902) );
  AND2_X1 U6022 ( .A1(n10601), .A2(n8233), .ZN(n4903) );
  AND2_X1 U6023 ( .A1(n4870), .A2(n7123), .ZN(n4904) );
  AND2_X1 U6024 ( .A1(n9051), .A2(n5384), .ZN(n4905) );
  INV_X1 U6025 ( .A(n9304), .ZN(n9055) );
  AND2_X1 U6026 ( .A1(n5387), .A2(n5093), .ZN(n4906) );
  OR2_X1 U6027 ( .A1(n4898), .A2(n6581), .ZN(n4907) );
  OR2_X1 U6028 ( .A1(n5062), .A2(n5065), .ZN(n4908) );
  AND2_X1 U6029 ( .A1(n5367), .A2(n5366), .ZN(n5365) );
  INV_X1 U6030 ( .A(n4852), .ZN(n6504) );
  OR2_X1 U6031 ( .A1(n5286), .A2(n6039), .ZN(n4909) );
  OAI21_X1 U6032 ( .B1(n8503), .B2(n5091), .A(n5089), .ZN(n8535) );
  OAI211_X1 U6033 ( .C1(n6328), .C2(n7244), .A(n6299), .B(n6298), .ZN(n10473)
         );
  NAND2_X1 U6034 ( .A1(n6829), .A2(n6216), .ZN(n6832) );
  AND2_X1 U6035 ( .A1(n4863), .A2(n5480), .ZN(n4910) );
  AND2_X1 U6036 ( .A1(n8475), .A2(n8468), .ZN(n4911) );
  INV_X1 U6037 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n4986) );
  XNOR2_X1 U6038 ( .A(n6202), .B(n6201), .ZN(n7066) );
  NAND2_X1 U6039 ( .A1(n8342), .A2(n7108), .ZN(n8415) );
  NAND2_X1 U6040 ( .A1(n6414), .A2(n6704), .ZN(n8503) );
  OAI21_X1 U6041 ( .B1(n10012), .B2(n4869), .A(n7119), .ZN(n9996) );
  NAND2_X1 U6042 ( .A1(n5074), .A2(n8629), .ZN(n9469) );
  INV_X1 U6043 ( .A(n7045), .ZN(n5196) );
  NAND2_X1 U6044 ( .A1(n5027), .A2(n8468), .ZN(n8480) );
  AND2_X1 U6045 ( .A1(n6631), .A2(n5388), .ZN(n6829) );
  NAND2_X1 U6046 ( .A1(n8297), .A2(n7106), .ZN(n8296) );
  NAND2_X1 U6047 ( .A1(n5539), .A2(n5538), .ZN(n4912) );
  NAND2_X1 U6048 ( .A1(n8520), .A2(n7112), .ZN(n8554) );
  AND2_X1 U6049 ( .A1(n8296), .A2(n7107), .ZN(n8341) );
  NAND2_X1 U6050 ( .A1(n9230), .A2(n9210), .ZN(n9206) );
  AND2_X1 U6051 ( .A1(n6971), .A2(n6970), .ZN(n4913) );
  NAND2_X1 U6052 ( .A1(n8422), .A2(n7037), .ZN(n8521) );
  INV_X1 U6053 ( .A(n5204), .ZN(n5203) );
  NAND2_X1 U6054 ( .A1(n5208), .A2(n8609), .ZN(n5204) );
  INV_X1 U6055 ( .A(n5161), .ZN(n9189) );
  NOR2_X1 U6056 ( .A1(n9206), .A2(n9321), .ZN(n5161) );
  NAND2_X1 U6057 ( .A1(n9995), .A2(n5005), .ZN(n5008) );
  AND2_X1 U6058 ( .A1(n8137), .A2(n6680), .ZN(n4914) );
  AND2_X1 U6059 ( .A1(n5340), .A2(n4896), .ZN(n4915) );
  NAND2_X1 U6060 ( .A1(n5899), .A2(n5898), .ZN(n10157) );
  INV_X1 U6061 ( .A(n10157), .ZN(n5012) );
  INV_X1 U6062 ( .A(n7080), .ZN(n5026) );
  INV_X1 U6063 ( .A(n8456), .ZN(n4946) );
  NAND2_X1 U6064 ( .A1(n8376), .A2(n5350), .ZN(n8492) );
  NAND2_X1 U6065 ( .A1(n5349), .A2(n7865), .ZN(n7961) );
  NAND2_X1 U6066 ( .A1(n5314), .A2(n7775), .ZN(n7770) );
  INV_X1 U6067 ( .A(n8136), .ZN(n5343) );
  NAND2_X1 U6068 ( .A1(n4977), .A2(n6802), .ZN(n8133) );
  NAND2_X1 U6069 ( .A1(n6448), .A2(n6447), .ZN(n9349) );
  INV_X1 U6070 ( .A(n9349), .ZN(n5162) );
  NAND2_X1 U6071 ( .A1(n7729), .A2(n6658), .ZN(n10435) );
  NAND2_X1 U6072 ( .A1(n5030), .A2(n4884), .ZN(n8260) );
  NAND2_X1 U6073 ( .A1(n8282), .A2(n5351), .ZN(n8376) );
  NAND2_X1 U6074 ( .A1(n8133), .A2(n5341), .ZN(n8234) );
  NAND2_X1 U6075 ( .A1(n7098), .A2(n7097), .ZN(n10479) );
  INV_X1 U6076 ( .A(n8245), .ZN(n5147) );
  OR3_X1 U6077 ( .A1(n8344), .A2(n10152), .A3(n5011), .ZN(n4916) );
  NAND2_X1 U6078 ( .A1(n5356), .A2(n7100), .ZN(n10533) );
  AND2_X1 U6079 ( .A1(n8369), .A2(n5165), .ZN(n4917) );
  AND2_X1 U6080 ( .A1(n8266), .A2(n8265), .ZN(n8322) );
  NAND2_X2 U6081 ( .A1(n5555), .A2(n5544), .ZN(n6205) );
  INV_X1 U6082 ( .A(n10580), .ZN(n5000) );
  XOR2_X1 U6083 ( .A(n6878), .B(n6879), .Z(n4918) );
  INV_X1 U6084 ( .A(n7763), .ZN(n5029) );
  AND4_X1 U6085 ( .A1(n6256), .A2(n6255), .A3(n6254), .A4(n6253), .ZN(n7687)
         );
  AND2_X1 U6086 ( .A1(n5572), .A2(n9682), .ZN(n4919) );
  AND2_X1 U6087 ( .A1(n7481), .A2(n6859), .ZN(n4920) );
  INV_X1 U6088 ( .A(n6227), .ZN(n9375) );
  INV_X1 U6089 ( .A(n9516), .ZN(n9556) );
  NAND3_X1 U6090 ( .A1(n4926), .A2(n9952), .A3(n6038), .ZN(n4925) );
  NAND3_X1 U6091 ( .A1(n6036), .A2(n6037), .A3(n9967), .ZN(n4926) );
  NAND2_X1 U6092 ( .A1(n4929), .A2(n6106), .ZN(n5926) );
  NAND2_X1 U6093 ( .A1(n5925), .A2(n7033), .ZN(n4929) );
  NAND2_X1 U6094 ( .A1(n4932), .A2(n4931), .ZN(n5842) );
  AOI21_X1 U6095 ( .B1(n4934), .B2(n7993), .A(n5811), .ZN(n4933) );
  XNOR2_X1 U6096 ( .A(n10486), .B(n4850), .ZN(n4934) );
  NAND2_X2 U6097 ( .A1(n4935), .A2(n5173), .ZN(n10364) );
  NAND2_X1 U6098 ( .A1(n6154), .A2(n6155), .ZN(n7087) );
  NAND2_X1 U6099 ( .A1(n7512), .A2(n7676), .ZN(n6155) );
  NAND3_X1 U6100 ( .A1(n6142), .A2(n6065), .A3(n6139), .ZN(n4938) );
  NAND2_X1 U6101 ( .A1(n4939), .A2(n6020), .ZN(n6023) );
  NAND3_X1 U6102 ( .A1(n4940), .A2(n6019), .A3(n10021), .ZN(n4939) );
  NAND3_X1 U6103 ( .A1(n4942), .A2(n4941), .A3(n10030), .ZN(n4940) );
  OR2_X1 U6104 ( .A1(n5989), .A2(n7064), .ZN(n4941) );
  INV_X1 U6105 ( .A(n4943), .ZN(n5781) );
  OAI21_X1 U6106 ( .B1(n7744), .B2(n4943), .A(n10408), .ZN(n7745) );
  NAND2_X1 U6107 ( .A1(n4943), .A2(n7744), .ZN(n10408) );
  AND4_X2 U6108 ( .A1(n5401), .A2(n5396), .A3(n5397), .A4(n5400), .ZN(n5380)
         );
  NAND2_X1 U6109 ( .A1(n8907), .A2(n8908), .ZN(n8906) );
  NAND2_X1 U6110 ( .A1(n8877), .A2(n8876), .ZN(n4953) );
  INV_X1 U6111 ( .A(n6964), .ZN(n4951) );
  NAND2_X1 U6112 ( .A1(n4953), .A2(n6964), .ZN(n8866) );
  NAND2_X1 U6113 ( .A1(n5739), .A2(n5740), .ZN(n4959) );
  NAND2_X2 U6114 ( .A1(n4960), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n5293) );
  OAI21_X2 U6115 ( .B1(P1_ADDR_REG_19__SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        n5409), .ZN(n5292) );
  NAND2_X2 U6116 ( .A1(n9163), .A2(n9162), .ZN(n9164) );
  NAND3_X1 U6117 ( .A1(n4994), .A2(n5349), .A3(n4901), .ZN(n7969) );
  NAND4_X1 U6118 ( .A1(n4998), .A2(n4999), .A3(n5374), .A4(n5547), .ZN(n5551)
         );
  INV_X1 U6119 ( .A(n5002), .ZN(n8193) );
  INV_X1 U6120 ( .A(n5008), .ZN(n9947) );
  NAND3_X1 U6121 ( .A1(n5016), .A2(n10073), .A3(n5013), .ZN(n10175) );
  NAND2_X2 U6122 ( .A1(n4854), .A2(n5021), .ZN(n5771) );
  NAND2_X1 U6123 ( .A1(n5243), .A2(n5023), .ZN(n8353) );
  NAND2_X1 U6124 ( .A1(n5024), .A2(n8264), .ZN(n8324) );
  INV_X1 U6125 ( .A(n8266), .ZN(n5024) );
  NAND2_X1 U6126 ( .A1(n8097), .A2(n5031), .ZN(n5030) );
  NAND2_X1 U6127 ( .A1(n9539), .A2(n5038), .ZN(n5037) );
  OAI211_X1 U6128 ( .C1(n9539), .C2(n5042), .A(n5039), .B(n5037), .ZN(n8729)
         );
  NAND2_X1 U6129 ( .A1(n9539), .A2(n9538), .ZN(n9537) );
  NAND2_X1 U6130 ( .A1(n9422), .A2(n5053), .ZN(n5049) );
  NAND2_X1 U6131 ( .A1(n5049), .A2(n5050), .ZN(n8677) );
  NAND2_X1 U6132 ( .A1(n9455), .A2(n4908), .ZN(n5059) );
  NAND2_X1 U6133 ( .A1(n5059), .A2(n5060), .ZN(n9421) );
  NAND2_X1 U6134 ( .A1(n9175), .A2(n5080), .ZN(n5079) );
  INV_X1 U6135 ( .A(n9112), .ZN(n5083) );
  OAI21_X1 U6136 ( .B1(n5083), .B2(n4907), .A(n5084), .ZN(n9085) );
  NAND2_X1 U6137 ( .A1(n5792), .A2(n5793), .ZN(n5086) );
  INV_X1 U6138 ( .A(n8503), .ZN(n5087) );
  OAI211_X1 U6139 ( .C1(n5090), .C2(n5087), .A(n5088), .B(n6471), .ZN(n6477)
         );
  NAND3_X1 U6140 ( .A1(n5094), .A2(n9283), .A3(n4906), .ZN(n9355) );
  NAND3_X1 U6141 ( .A1(n5292), .A2(n5293), .A3(P2_DATAO_REG_2__SCAN_IN), .ZN(
        n5414) );
  OAI21_X2 U6142 ( .B1(n8138), .B2(n5241), .A(n5096), .ZN(n8227) );
  INV_X1 U6143 ( .A(n5424), .ZN(n5098) );
  NAND2_X1 U6144 ( .A1(n5102), .A2(n6764), .ZN(n5101) );
  NAND2_X1 U6145 ( .A1(n5101), .A2(n5100), .ZN(n5105) );
  NAND2_X1 U6146 ( .A1(n4861), .A2(n9055), .ZN(n5103) );
  NAND2_X1 U6147 ( .A1(n5104), .A2(n6766), .ZN(n6767) );
  NAND2_X1 U6148 ( .A1(n6765), .A2(n5105), .ZN(n5104) );
  NAND2_X1 U6149 ( .A1(n5891), .A2(n4902), .ZN(n5114) );
  NAND2_X1 U6150 ( .A1(n5116), .A2(n5413), .ZN(n5739) );
  MUX2_X1 U6151 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(P1_DATAO_REG_1__SCAN_IN), 
        .S(n5552), .Z(n5720) );
  OAI21_X1 U6152 ( .B1(n5951), .B2(n5120), .A(n5117), .ZN(n6006) );
  NAND2_X1 U6153 ( .A1(n5951), .A2(n5950), .ZN(n5123) );
  NAND3_X1 U6154 ( .A1(n5124), .A2(n5125), .A3(n5267), .ZN(n5453) );
  NAND2_X1 U6155 ( .A1(n5835), .A2(n5127), .ZN(n5124) );
  NAND2_X1 U6156 ( .A1(n5835), .A2(n5439), .ZN(n5126) );
  OAI21_X1 U6157 ( .B1(n5835), .B2(n5834), .A(n5439), .ZN(n5701) );
  NAND4_X1 U6158 ( .A1(n6774), .A2(n6790), .A3(n6772), .A4(n6773), .ZN(n5137)
         );
  INV_X2 U6159 ( .A(n7172), .ZN(n7177) );
  NAND2_X1 U6160 ( .A1(n8866), .A2(n4862), .ZN(n5141) );
  NAND3_X1 U6161 ( .A1(n7561), .A2(n7857), .A3(n5144), .ZN(n6798) );
  NAND4_X1 U6162 ( .A1(n7602), .A2(n7481), .A3(n7558), .A4(n6859), .ZN(n5145)
         );
  NAND2_X1 U6163 ( .A1(n7483), .A2(n7482), .ZN(n7481) );
  NAND2_X1 U6164 ( .A1(n6871), .A2(n7782), .ZN(n7781) );
  NAND2_X1 U6165 ( .A1(n8845), .A2(n6902), .ZN(n5149) );
  NAND2_X1 U6166 ( .A1(n9107), .A2(n5153), .ZN(n9074) );
  AND3_X2 U6167 ( .A1(n6214), .A2(n4872), .A3(n5219), .ZN(n6631) );
  NAND2_X1 U6168 ( .A1(n6459), .A2(n5156), .ZN(n5157) );
  NAND2_X1 U6169 ( .A1(n6490), .A2(n6489), .ZN(n6491) );
  INV_X1 U6170 ( .A(n9206), .ZN(n5159) );
  NAND2_X1 U6171 ( .A1(n5168), .A2(n10575), .ZN(n5166) );
  NAND2_X1 U6172 ( .A1(n5325), .A2(n5324), .ZN(n8891) );
  NAND2_X1 U6173 ( .A1(n6913), .A2(n8390), .ZN(n8386) );
  NAND2_X1 U6174 ( .A1(n8858), .A2(n8859), .ZN(n5325) );
  NAND2_X2 U6175 ( .A1(n6849), .A2(n9029), .ZN(n7009) );
  AOI21_X2 U6176 ( .B1(n6623), .B2(n6816), .A(n6633), .ZN(n6630) );
  INV_X1 U6177 ( .A(n5227), .ZN(n5226) );
  NAND2_X1 U6178 ( .A1(n5549), .A2(n5548), .ZN(n5550) );
  NAND2_X1 U6179 ( .A1(n8176), .A2(n6897), .ZN(n8844) );
  INV_X1 U6180 ( .A(n5316), .ZN(n5315) );
  NAND2_X1 U6181 ( .A1(n7647), .A2(n7648), .ZN(n9491) );
  NAND2_X1 U6182 ( .A1(n5380), .A2(n5404), .ZN(n5186) );
  NAND2_X1 U6183 ( .A1(n8353), .A2(n8352), .ZN(n8464) );
  NAND2_X1 U6184 ( .A1(n5200), .A2(n5199), .ZN(n9455) );
  NAND2_X1 U6185 ( .A1(n9920), .A2(n7056), .ZN(n8585) );
  NAND2_X1 U6186 ( .A1(n7036), .A2(n4900), .ZN(n8422) );
  NAND2_X1 U6187 ( .A1(n7036), .A2(n7035), .ZN(n8420) );
  INV_X1 U6188 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5189) );
  OAI21_X1 U6189 ( .B1(n10020), .B2(n5194), .A(n5191), .ZN(n7048) );
  OAI21_X2 U6190 ( .B1(n5781), .B2(n6157), .A(n5780), .ZN(n10486) );
  NAND2_X1 U6191 ( .A1(n5198), .A2(P1_IR_REG_29__SCAN_IN), .ZN(n5558) );
  NAND2_X1 U6192 ( .A1(n5545), .A2(n5541), .ZN(n5555) );
  NAND2_X1 U6193 ( .A1(n8610), .A2(n5201), .ZN(n5200) );
  AOI21_X1 U6194 ( .B1(n5207), .B2(n8616), .A(n5206), .ZN(n5205) );
  INV_X1 U6195 ( .A(n9403), .ZN(n5206) );
  INV_X1 U6196 ( .A(n8609), .ZN(n5207) );
  INV_X1 U6197 ( .A(n8616), .ZN(n5208) );
  NAND2_X1 U6198 ( .A1(n5209), .A2(n8616), .ZN(n9400) );
  INV_X1 U6199 ( .A(n5702), .ZN(n5379) );
  INV_X1 U6200 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5210) );
  NAND2_X1 U6201 ( .A1(n9245), .A2(n5214), .ZN(n5211) );
  NAND2_X1 U6202 ( .A1(n5211), .A2(n5212), .ZN(n9211) );
  NAND2_X1 U6203 ( .A1(n9413), .A2(n5235), .ZN(n5230) );
  NAND3_X1 U6204 ( .A1(n5231), .A2(n5230), .A3(n5229), .ZN(n9539) );
  INV_X1 U6205 ( .A(n8322), .ZN(n5244) );
  INV_X1 U6206 ( .A(n8329), .ZN(n5242) );
  NAND2_X1 U6207 ( .A1(n5245), .A2(n5246), .ZN(n7858) );
  NAND3_X1 U6208 ( .A1(n7729), .A2(n6666), .A3(n4859), .ZN(n5245) );
  NAND2_X1 U6209 ( .A1(n8944), .A2(n10392), .ZN(n6657) );
  AND2_X1 U6210 ( .A1(n6264), .A2(n5248), .ZN(n5247) );
  NAND3_X1 U6211 ( .A1(n7638), .A2(n7637), .A3(n9521), .ZN(n9520) );
  NAND2_X1 U6212 ( .A1(n7638), .A2(n7637), .ZN(n5257) );
  NAND2_X1 U6213 ( .A1(n9520), .A2(n5255), .ZN(n9522) );
  NAND2_X1 U6214 ( .A1(n5257), .A2(n5256), .ZN(n5255) );
  INV_X1 U6215 ( .A(n9521), .ZN(n5256) );
  OAI21_X1 U6216 ( .B1(n5969), .B2(n5481), .A(n5480), .ZN(n5991) );
  NAND2_X1 U6217 ( .A1(n5445), .A2(n5444), .ZN(n5843) );
  INV_X1 U6218 ( .A(n5390), .ZN(n5271) );
  NAND2_X1 U6219 ( .A1(n5584), .A2(n5278), .ZN(n5276) );
  NAND2_X1 U6220 ( .A1(n5584), .A2(n5583), .ZN(n5277) );
  NAND2_X1 U6221 ( .A1(n5661), .A2(n5284), .ZN(n5281) );
  NAND2_X1 U6222 ( .A1(n5281), .A2(n5282), .ZN(n5523) );
  NAND2_X1 U6223 ( .A1(n5661), .A2(n5510), .ZN(n5648) );
  NAND3_X1 U6224 ( .A1(n5292), .A2(n5293), .A3(n5410), .ZN(n5730) );
  OR2_X2 U6225 ( .A1(n8844), .A2(n8843), .ZN(n8845) );
  OR2_X1 U6226 ( .A1(n8920), .A2(n5303), .ZN(n5298) );
  NAND3_X1 U6227 ( .A1(n5298), .A2(n5297), .A3(n5299), .ZN(n7018) );
  NAND2_X1 U6228 ( .A1(n8920), .A2(n5304), .ZN(n5297) );
  NAND2_X1 U6229 ( .A1(n7781), .A2(n5315), .ZN(n5312) );
  NAND2_X1 U6230 ( .A1(n5313), .A2(n5312), .ZN(n7829) );
  NAND2_X1 U6231 ( .A1(n9121), .A2(n5330), .ZN(n5327) );
  NAND2_X1 U6232 ( .A1(n5327), .A2(n5328), .ZN(n9081) );
  NAND2_X1 U6233 ( .A1(n9204), .A2(n4905), .ZN(n9185) );
  NAND2_X1 U6234 ( .A1(n8540), .A2(n5339), .ZN(n5336) );
  INV_X1 U6235 ( .A(n5340), .ZN(n9044) );
  NAND2_X1 U6236 ( .A1(n5345), .A2(n5344), .ZN(n10428) );
  NAND2_X1 U6237 ( .A1(n7095), .A2(n7094), .ZN(n7989) );
  NAND3_X1 U6238 ( .A1(n5768), .A2(n5767), .A3(n7753), .ZN(n10407) );
  NAND2_X1 U6239 ( .A1(n8517), .A2(n7112), .ZN(n5353) );
  NAND2_X1 U6240 ( .A1(n5356), .A2(n5354), .ZN(n10532) );
  NAND2_X1 U6241 ( .A1(n10012), .A2(n5361), .ZN(n5357) );
  NAND2_X1 U6242 ( .A1(n5357), .A2(n5358), .ZN(n9976) );
  NAND2_X1 U6243 ( .A1(n7127), .A2(n5365), .ZN(n5363) );
  NAND2_X1 U6244 ( .A1(n5363), .A2(n5364), .ZN(n9895) );
  NAND2_X1 U6245 ( .A1(n7127), .A2(n7055), .ZN(n9913) );
  NAND2_X1 U6246 ( .A1(n7124), .A2(n4904), .ZN(n9933) );
  INV_X1 U6247 ( .A(n5371), .ZN(n5370) );
  NAND2_X1 U6248 ( .A1(n5376), .A2(n4879), .ZN(n8189) );
  NAND3_X1 U6249 ( .A1(n5381), .A2(n5380), .A3(n5379), .ZN(n5408) );
  NAND2_X1 U6250 ( .A1(n5545), .A2(n5382), .ZN(n5560) );
  OR2_X1 U6251 ( .A1(n7491), .A2(n7766), .ZN(n7086) );
  OR2_X1 U6252 ( .A1(n7759), .A2(n8701), .ZN(n7378) );
  INV_X1 U6253 ( .A(n7505), .ZN(n7508) );
  AOI21_X1 U6254 ( .B1(n9129), .B2(n6286), .A(n6557), .ZN(n9144) );
  INV_X1 U6255 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5820) );
  AND2_X2 U6256 ( .A1(n5602), .A2(n5562), .ZN(n5760) );
  INV_X1 U6257 ( .A(n6605), .ZN(n6616) );
  NAND2_X1 U6258 ( .A1(n5763), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5725) );
  INV_X1 U6259 ( .A(n5562), .ZN(n5603) );
  OR2_X1 U6260 ( .A1(n7129), .A2(n8397), .ZN(n5383) );
  INV_X1 U6261 ( .A(n9159), .ZN(n9311) );
  INV_X1 U6262 ( .A(n8371), .ZN(n10654) );
  OR2_X1 U6263 ( .A1(n9210), .A2(n9196), .ZN(n5384) );
  NAND2_X1 U6264 ( .A1(n5581), .A2(n6090), .ZN(n5385) );
  NAND4_X1 U6265 ( .A1(n6148), .A2(n7130), .A3(n6147), .A4(n8311), .ZN(n5386)
         );
  XNOR2_X1 U6266 ( .A(n8943), .B(n10434), .ZN(n10437) );
  OR2_X1 U6267 ( .A1(n9281), .A2(n10673), .ZN(n5387) );
  AND3_X1 U6268 ( .A1(n6826), .A2(n6834), .A3(n6215), .ZN(n5388) );
  INV_X1 U6269 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n5415) );
  AND2_X1 U6270 ( .A1(n7567), .A2(n7009), .ZN(n10662) );
  INV_X1 U6271 ( .A(n10662), .ZN(n10672) );
  INV_X1 U6272 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n6356) );
  AND2_X1 U6273 ( .A1(n5444), .A2(n5443), .ZN(n5389) );
  INV_X1 U6274 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n5435) );
  INV_X1 U6275 ( .A(n10436), .ZN(n10616) );
  AND2_X1 U6276 ( .A1(n5449), .A2(n5448), .ZN(n5390) );
  AND2_X1 U6277 ( .A1(n6593), .A2(n6592), .ZN(n9069) );
  AND4_X1 U6278 ( .A1(n6429), .A2(n6428), .A3(n6427), .A4(n6426), .ZN(n8783)
         );
  OR2_X1 U6279 ( .A1(n7137), .A2(n7136), .ZN(P1_U3264) );
  INV_X1 U6280 ( .A(n8801), .ZN(n9905) );
  INV_X1 U6281 ( .A(n6790), .ZN(n9064) );
  AND4_X1 U6282 ( .A1(n9896), .A2(n8813), .A3(n6088), .A4(n6180), .ZN(n5392)
         );
  NAND2_X1 U6283 ( .A1(n6187), .A2(n7376), .ZN(n5393) );
  OR2_X1 U6284 ( .A1(n6187), .A2(n8116), .ZN(n5394) );
  INV_X1 U6285 ( .A(n10487), .ZN(n7097) );
  AND2_X1 U6286 ( .A1(n8014), .A2(n10005), .ZN(n10563) );
  INV_X1 U6287 ( .A(n10563), .ZN(n10568) );
  NAND2_X1 U6288 ( .A1(n5646), .A2(n5645), .ZN(n9923) );
  OR2_X1 U6289 ( .A1(n5745), .A2(n7323), .ZN(n5395) );
  INV_X1 U6290 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5547) );
  AND2_X1 U6291 ( .A1(n6539), .A2(n6538), .ZN(n9143) );
  INV_X1 U6292 ( .A(n9143), .ZN(n9179) );
  INV_X1 U6293 ( .A(n8868), .ZN(n9054) );
  AND2_X1 U6294 ( .A1(n6549), .A2(n6548), .ZN(n8868) );
  INV_X1 U6295 ( .A(n9141), .ZN(n6550) );
  INV_X1 U6296 ( .A(n8602), .ZN(n9127) );
  INV_X1 U6297 ( .A(n10631), .ZN(n10448) );
  INV_X1 U6298 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5556) );
  AND4_X1 U6299 ( .A1(n6413), .A2(n6412), .A3(n6411), .A4(n6410), .ZN(n8504)
         );
  NOR2_X1 U6300 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(n6212), .ZN(n6213) );
  OR2_X1 U6301 ( .A1(n9280), .A2(n7876), .ZN(n6776) );
  INV_X1 U6302 ( .A(n8783), .ZN(n8494) );
  NAND2_X1 U6303 ( .A1(n6089), .A2(n9884), .ZN(n5582) );
  OAI21_X1 U6304 ( .B1(n6142), .B2(n7064), .A(n5610), .ZN(n5611) );
  INV_X1 U6305 ( .A(n10135), .ZN(n7061) );
  NAND2_X1 U6306 ( .A1(n5541), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5542) );
  INV_X1 U6307 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5541) );
  INV_X1 U6308 ( .A(SI_10_), .ZN(n9716) );
  INV_X1 U6309 ( .A(n6532), .ZN(n6531) );
  INV_X1 U6310 ( .A(n7145), .ZN(n6886) );
  INV_X1 U6311 ( .A(n6561), .ZN(n6560) );
  INV_X1 U6312 ( .A(n6496), .ZN(n6494) );
  OR2_X1 U6313 ( .A1(n6586), .A2(n6585), .ZN(n6598) );
  OR2_X1 U6314 ( .A1(n6450), .A2(n6449), .ZN(n6464) );
  NAND2_X1 U6315 ( .A1(n5155), .A2(n9069), .ZN(n9061) );
  INV_X1 U6316 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n6458) );
  INV_X1 U6317 ( .A(n5667), .ZN(n5599) );
  INV_X1 U6318 ( .A(n6184), .ZN(n6147) );
  INV_X1 U6319 ( .A(n6030), .ZN(n5598) );
  INV_X1 U6320 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5710) );
  OR2_X1 U6321 ( .A1(n5640), .A2(n5626), .ZN(n5628) );
  INV_X1 U6322 ( .A(n6014), .ZN(n5597) );
  OR2_X1 U6323 ( .A1(n5941), .A2(n9557), .ZN(n5957) );
  INV_X1 U6324 ( .A(n10544), .ZN(n7101) );
  NAND2_X1 U6325 ( .A1(n10364), .A2(n7763), .ZN(n6154) );
  INV_X1 U6326 ( .A(n5892), .ZN(n5461) );
  NAND2_X1 U6327 ( .A1(n5441), .A2(n9712), .ZN(n5444) );
  NAND2_X1 U6328 ( .A1(n6531), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6542) );
  NAND2_X1 U6329 ( .A1(n6315), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6331) );
  NAND2_X1 U6330 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n6288) );
  INV_X1 U6331 ( .A(n8893), .ZN(n6953) );
  NAND2_X1 U6332 ( .A1(n6560), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6572) );
  OR2_X1 U6333 ( .A1(n6542), .A2(n9761), .ZN(n6552) );
  NAND2_X1 U6334 ( .A1(n6494), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6509) );
  AND2_X1 U6335 ( .A1(n6605), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6225) );
  INV_X1 U6336 ( .A(n9280), .ZN(n8603) );
  AND2_X1 U6337 ( .A1(n6598), .A2(n6587), .ZN(n9082) );
  INV_X1 U6338 ( .A(n9188), .ZN(n9051) );
  INV_X1 U6339 ( .A(n5919), .ZN(n5593) );
  INV_X1 U6340 ( .A(n6012), .ZN(n5596) );
  INV_X1 U6341 ( .A(n7506), .ZN(n7507) );
  INV_X1 U6342 ( .A(n5957), .ZN(n5594) );
  OR2_X1 U6343 ( .A1(n5852), .A2(n5851), .ZN(n5865) );
  NAND2_X1 U6344 ( .A1(n5598), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n5667) );
  INV_X1 U6345 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n9667) );
  AND2_X1 U6346 ( .A1(n5628), .A2(n5627), .ZN(n9393) );
  INV_X1 U6347 ( .A(n8311), .ZN(n7129) );
  INV_X1 U6348 ( .A(n7403), .ZN(n7405) );
  INV_X1 U6349 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n10195) );
  INV_X1 U6350 ( .A(n5658), .ZN(n5660) );
  INV_X1 U6351 ( .A(n5676), .ZN(n5499) );
  INV_X1 U6352 ( .A(n5934), .ZN(n5471) );
  OR2_X1 U6353 ( .A1(n5910), .A2(n5970), .ZN(n5879) );
  CLKBUF_X3 U6354 ( .A(n5418), .Z(n6238) );
  INV_X1 U6355 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n5420) );
  OR2_X1 U6356 ( .A1(n6357), .A2(n6356), .ZN(n6376) );
  INV_X1 U6357 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n8068) );
  NAND2_X1 U6358 ( .A1(n6375), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6393) );
  INV_X1 U6359 ( .A(n8875), .ZN(n8902) );
  INV_X1 U6360 ( .A(n6286), .ZN(n6574) );
  AND2_X1 U6361 ( .A1(n6794), .A2(n6793), .ZN(n8236) );
  INV_X1 U6362 ( .A(n10437), .ZN(n6285) );
  AND2_X1 U6363 ( .A1(n6991), .A2(n6990), .ZN(n7425) );
  NAND2_X1 U6364 ( .A1(n9211), .A2(n6811), .ZN(n9216) );
  OR2_X1 U6365 ( .A1(n10215), .A2(n6992), .ZN(n7441) );
  NAND2_X1 U6366 ( .A1(n8705), .A2(n8707), .ZN(n8708) );
  NAND2_X1 U6367 ( .A1(n5593), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n5941) );
  INV_X1 U6368 ( .A(n9923), .ZN(n9451) );
  NAND2_X1 U6369 ( .A1(n5594), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5998) );
  OR2_X1 U6370 ( .A1(n5901), .A2(n5900), .ZN(n5919) );
  NAND2_X1 U6371 ( .A1(n5591), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5883) );
  OR2_X1 U6372 ( .A1(n5998), .A2(n5595), .ZN(n6012) );
  OR2_X1 U6373 ( .A1(n7514), .A2(n7513), .ZN(n9542) );
  OR2_X1 U6374 ( .A1(n9903), .A2(n6035), .ZN(n5621) );
  NAND2_X1 U6375 ( .A1(n5763), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5719) );
  AND2_X1 U6376 ( .A1(n8041), .A2(n8040), .ZN(n8042) );
  INV_X1 U6377 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n9877) );
  AND2_X1 U6378 ( .A1(n8810), .A2(n8811), .ZN(n9896) );
  AND4_X1 U6379 ( .A1(n5946), .A2(n5945), .A3(n5944), .A4(n5943), .ZN(n9465)
         );
  AND2_X1 U6380 ( .A1(n7129), .A2(n7130), .ZN(n7385) );
  INV_X1 U6381 ( .A(n10582), .ZN(n10366) );
  AND2_X1 U6382 ( .A1(n5494), .A2(n5493), .ZN(n5684) );
  AND2_X1 U6383 ( .A1(n5478), .A2(n5477), .ZN(n5950) );
  XNOR2_X1 U6384 ( .A(n5464), .B(n5463), .ZN(n5907) );
  OR2_X1 U6385 ( .A1(n7157), .A2(n6840), .ZN(n7442) );
  OAI21_X1 U6386 ( .B1(n7015), .B2(n8871), .A(n7014), .ZN(n7016) );
  INV_X1 U6387 ( .A(n8922), .ZN(n8915) );
  OR2_X1 U6388 ( .A1(n8830), .A2(n6574), .ZN(n6580) );
  AND4_X1 U6389 ( .A1(n6457), .A2(n6456), .A3(n6455), .A4(n6454), .ZN(n8775)
         );
  AND2_X1 U6390 ( .A1(n7164), .A2(n6841), .ZN(n10320) );
  INV_X1 U6391 ( .A(n6811), .ZN(n9212) );
  INV_X1 U6392 ( .A(n10454), .ZN(n10626) );
  NAND2_X1 U6393 ( .A1(n10213), .A2(n6995), .ZN(n10446) );
  INV_X1 U6394 ( .A(n7860), .ZN(n7730) );
  AND2_X1 U6395 ( .A1(n7427), .A2(n7425), .ZN(n7445) );
  INV_X1 U6396 ( .A(n10677), .ZN(n10667) );
  AND2_X1 U6397 ( .A1(n6994), .A2(n6849), .ZN(n10622) );
  AND2_X1 U6398 ( .A1(n7427), .A2(n7426), .ZN(n7691) );
  XNOR2_X1 U6399 ( .A(n6837), .B(P2_IR_REG_24__SCAN_IN), .ZN(n10308) );
  AND2_X1 U6400 ( .A1(n6368), .A2(n6371), .ZN(n7940) );
  INV_X1 U6401 ( .A(n9542), .ZN(n9558) );
  INV_X1 U6402 ( .A(n6032), .ZN(n6050) );
  INV_X1 U6403 ( .A(n6047), .ZN(n6035) );
  AND4_X1 U6404 ( .A1(n5962), .A2(n5961), .A3(n5960), .A4(n5959), .ZN(n9562)
         );
  AND2_X1 U6405 ( .A1(n7266), .A2(n10256), .ZN(n10349) );
  INV_X1 U6406 ( .A(n10067), .ZN(n9889) );
  AND2_X1 U6407 ( .A1(n7049), .A2(n7050), .ZN(n9967) );
  AND2_X1 U6408 ( .A1(n8520), .A2(n8519), .ZN(n10145) );
  AND2_X1 U6409 ( .A1(n7465), .A2(n7385), .ZN(n10540) );
  INV_X1 U6410 ( .A(n8598), .ZN(n10559) );
  INV_X1 U6411 ( .A(n10565), .ZN(n10042) );
  AND2_X1 U6412 ( .A1(n7069), .A2(n10194), .ZN(n7411) );
  AND2_X1 U6413 ( .A1(n10550), .A2(n10370), .ZN(n10460) );
  INV_X1 U6414 ( .A(n7411), .ZN(n7417) );
  XNOR2_X1 U6415 ( .A(n6040), .B(n6039), .ZN(n8574) );
  AND2_X1 U6416 ( .A1(n5976), .A2(n5992), .ZN(n9849) );
  XNOR2_X1 U6417 ( .A(n5432), .B(SI_7_), .ZN(n5822) );
  INV_X1 U6418 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n8731) );
  NOR2_X1 U6419 ( .A1(n10240), .A2(n10239), .ZN(n8757) );
  NAND2_X1 U6420 ( .A1(n8836), .A2(n6955), .ZN(n8842) );
  INV_X1 U6421 ( .A(n9069), .ZN(n9100) );
  AND4_X1 U6422 ( .A1(n6503), .A2(n6502), .A3(n6501), .A4(n6500), .ZN(n9248)
         );
  INV_X1 U6423 ( .A(n10451), .ZN(n10634) );
  AND2_X1 U6424 ( .A1(n7700), .A2(n10446), .ZN(n10631) );
  INV_X1 U6425 ( .A(n10681), .ZN(n10679) );
  INV_X1 U6426 ( .A(n10684), .ZN(n10682) );
  AND2_X2 U6427 ( .A1(n7691), .A2(n7428), .ZN(n10684) );
  INV_X1 U6428 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n7293) );
  INV_X1 U6429 ( .A(n9564), .ZN(n9548) );
  INV_X1 U6430 ( .A(n9898), .ZN(n9571) );
  OR2_X1 U6431 ( .A1(n5695), .A2(n5694), .ZN(n10022) );
  OR2_X1 U6432 ( .A1(P1_U3083), .A2(n7262), .ZN(n10342) );
  INV_X1 U6433 ( .A(n10349), .ZN(n10299) );
  OR2_X1 U6434 ( .A1(n9977), .A2(n7628), .ZN(n10046) );
  INV_X1 U6435 ( .A(n10568), .ZN(n9977) );
  AND2_X1 U6436 ( .A1(n8083), .A2(n8082), .ZN(n10588) );
  OR2_X1 U6437 ( .A1(n9977), .A2(n9998), .ZN(n8598) );
  INV_X1 U6438 ( .A(n10590), .ZN(n10589) );
  AND2_X2 U6439 ( .A1(n7418), .A2(n7411), .ZN(n10590) );
  AND2_X1 U6440 ( .A1(n10588), .A2(n10587), .ZN(n10593) );
  INV_X1 U6441 ( .A(n10594), .ZN(n10591) );
  INV_X1 U6442 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n7291) );
  INV_X1 U6443 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n7246) );
  NOR2_X1 U6444 ( .A1(n8758), .A2(n8757), .ZN(n10242) );
  INV_X1 U6445 ( .A(n8945), .ZN(P2_U3966) );
  NAND2_X1 U6446 ( .A1(n6209), .A2(n6208), .ZN(P1_U3240) );
  INV_X2 U6447 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  NOR2_X1 U6448 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n5399) );
  NOR2_X1 U6449 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n5398) );
  INV_X1 U6450 ( .A(n5539), .ZN(n5405) );
  NAND2_X1 U6451 ( .A1(n5405), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6069) );
  INV_X1 U6452 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n6068) );
  NAND2_X1 U6453 ( .A1(n6069), .A2(n6068), .ZN(n6071) );
  NAND2_X1 U6454 ( .A1(n6071), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5407) );
  INV_X1 U6455 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5406) );
  AND2_X1 U6456 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5410) );
  AND2_X1 U6457 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n5411) );
  NAND2_X1 U6458 ( .A1(n5552), .A2(n5411), .ZN(n6250) );
  INV_X1 U6459 ( .A(SI_1_), .ZN(n9728) );
  NAND2_X1 U6460 ( .A1(n5412), .A2(SI_1_), .ZN(n5413) );
  INV_X1 U6461 ( .A(SI_2_), .ZN(n9729) );
  XNOR2_X1 U6462 ( .A(n5416), .B(n9729), .ZN(n5740) );
  NAND2_X1 U6463 ( .A1(n5416), .A2(SI_2_), .ZN(n5417) );
  INV_X1 U6464 ( .A(SI_3_), .ZN(n5421) );
  XNOR2_X1 U6465 ( .A(n5422), .B(n5421), .ZN(n5772) );
  NAND2_X1 U6466 ( .A1(n5422), .A2(SI_3_), .ZN(n5423) );
  MUX2_X1 U6467 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n6238), .Z(n5427) );
  INV_X1 U6468 ( .A(SI_5_), .ZN(n5426) );
  XNOR2_X1 U6469 ( .A(n5427), .B(n5426), .ZN(n5793) );
  NAND2_X1 U6470 ( .A1(n5427), .A2(SI_5_), .ZN(n5428) );
  MUX2_X1 U6471 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n6238), .Z(n5430) );
  NAND2_X1 U6472 ( .A1(n5430), .A2(SI_6_), .ZN(n5431) );
  MUX2_X1 U6473 ( .A(n7372), .B(n7246), .S(n6238), .Z(n5432) );
  INV_X1 U6474 ( .A(n5432), .ZN(n5433) );
  NAND2_X1 U6475 ( .A1(n5433), .A2(SI_7_), .ZN(n5434) );
  MUX2_X1 U6476 ( .A(n7254), .B(n5435), .S(n6238), .Z(n5436) );
  INV_X1 U6477 ( .A(n5436), .ZN(n5437) );
  NAND2_X1 U6478 ( .A1(n5437), .A2(SI_8_), .ZN(n5438) );
  MUX2_X1 U6479 ( .A(n7258), .B(n5440), .S(n6238), .Z(n5441) );
  INV_X1 U6480 ( .A(n5441), .ZN(n5442) );
  NAND2_X1 U6481 ( .A1(n5442), .A2(SI_9_), .ZN(n5443) );
  MUX2_X1 U6482 ( .A(n7293), .B(n7291), .S(n6238), .Z(n5446) );
  NAND2_X1 U6483 ( .A1(n5446), .A2(n9716), .ZN(n5449) );
  INV_X1 U6484 ( .A(n5446), .ZN(n5447) );
  NAND2_X1 U6485 ( .A1(n5447), .A2(SI_10_), .ZN(n5448) );
  MUX2_X1 U6486 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .S(n6238), .Z(n5451) );
  MUX2_X1 U6487 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .S(n6238), .Z(n5452) );
  NAND2_X1 U6488 ( .A1(n5453), .A2(n5452), .ZN(n5454) );
  INV_X1 U6489 ( .A(SI_12_), .ZN(n9614) );
  INV_X1 U6490 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n5457) );
  INV_X1 U6491 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n5456) );
  MUX2_X1 U6492 ( .A(n5457), .B(n5456), .S(n5418), .Z(n5458) );
  NAND2_X1 U6493 ( .A1(n5458), .A2(n9675), .ZN(n5462) );
  INV_X1 U6494 ( .A(n5458), .ZN(n5459) );
  NAND2_X1 U6495 ( .A1(n5459), .A2(SI_13_), .ZN(n5460) );
  NAND2_X1 U6496 ( .A1(n5462), .A2(n5460), .ZN(n5892) );
  MUX2_X1 U6497 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n5418), .Z(n5464) );
  INV_X1 U6498 ( .A(n5907), .ZN(n5466) );
  NAND2_X1 U6499 ( .A1(n5464), .A2(SI_14_), .ZN(n5465) );
  INV_X1 U6500 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n5467) );
  MUX2_X1 U6501 ( .A(n5467), .B(n7819), .S(n5418), .Z(n5468) );
  NAND2_X1 U6502 ( .A1(n5468), .A2(n9705), .ZN(n5472) );
  INV_X1 U6503 ( .A(n5468), .ZN(n5469) );
  NAND2_X1 U6504 ( .A1(n5469), .A2(SI_15_), .ZN(n5470) );
  NAND2_X1 U6505 ( .A1(n5472), .A2(n5470), .ZN(n5934) );
  NAND2_X1 U6506 ( .A1(n5933), .A2(n5471), .ZN(n5937) );
  NAND2_X1 U6507 ( .A1(n5937), .A2(n5472), .ZN(n5951) );
  INV_X1 U6508 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n5474) );
  INV_X1 U6509 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n5473) );
  MUX2_X1 U6510 ( .A(n5474), .B(n5473), .S(n6238), .Z(n5475) );
  NAND2_X1 U6511 ( .A1(n5475), .A2(n9703), .ZN(n5478) );
  INV_X1 U6512 ( .A(n5475), .ZN(n5476) );
  NAND2_X1 U6513 ( .A1(n5476), .A2(SI_16_), .ZN(n5477) );
  MUX2_X1 U6514 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(P2_DATAO_REG_17__SCAN_IN), 
        .S(n5418), .Z(n5479) );
  XNOR2_X1 U6515 ( .A(n5479), .B(n9700), .ZN(n5968) );
  INV_X1 U6516 ( .A(n5968), .ZN(n5481) );
  NAND2_X1 U6517 ( .A1(n5479), .A2(SI_17_), .ZN(n5480) );
  MUX2_X1 U6518 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n6238), .Z(n5482) );
  XNOR2_X1 U6519 ( .A(n5482), .B(SI_18_), .ZN(n5990) );
  INV_X1 U6520 ( .A(n5482), .ZN(n5483) );
  INV_X1 U6521 ( .A(SI_18_), .ZN(n9677) );
  INV_X1 U6522 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n8113) );
  INV_X1 U6523 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n8114) );
  MUX2_X1 U6524 ( .A(n8113), .B(n8114), .S(n5418), .Z(n5486) );
  INV_X1 U6525 ( .A(SI_19_), .ZN(n5485) );
  NAND2_X1 U6526 ( .A1(n5486), .A2(n5485), .ZN(n5489) );
  INV_X1 U6527 ( .A(n5486), .ZN(n5487) );
  NAND2_X1 U6528 ( .A1(n5487), .A2(SI_19_), .ZN(n5488) );
  NAND2_X1 U6529 ( .A1(n5489), .A2(n5488), .ZN(n6004) );
  INV_X1 U6530 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n8244) );
  INV_X1 U6531 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n8165) );
  MUX2_X1 U6532 ( .A(n8244), .B(n8165), .S(n6238), .Z(n5491) );
  INV_X1 U6533 ( .A(SI_20_), .ZN(n5490) );
  NAND2_X1 U6534 ( .A1(n5491), .A2(n5490), .ZN(n5494) );
  INV_X1 U6535 ( .A(n5491), .ZN(n5492) );
  NAND2_X1 U6536 ( .A1(n5492), .A2(SI_20_), .ZN(n5493) );
  NAND2_X1 U6537 ( .A1(n5685), .A2(n5684), .ZN(n5495) );
  NAND2_X1 U6538 ( .A1(n5495), .A2(n5494), .ZN(n5677) );
  INV_X1 U6539 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n8204) );
  INV_X1 U6540 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n8184) );
  MUX2_X1 U6541 ( .A(n8204), .B(n8184), .S(n5418), .Z(n5496) );
  XNOR2_X1 U6542 ( .A(n5496), .B(SI_21_), .ZN(n5676) );
  INV_X1 U6543 ( .A(n5496), .ZN(n5497) );
  NAND2_X1 U6544 ( .A1(n5497), .A2(SI_21_), .ZN(n5498) );
  INV_X1 U6545 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n8308) );
  INV_X1 U6546 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8309) );
  MUX2_X1 U6547 ( .A(n8308), .B(n8309), .S(n6238), .Z(n5500) );
  INV_X1 U6548 ( .A(SI_22_), .ZN(n9595) );
  NAND2_X1 U6549 ( .A1(n5500), .A2(n9595), .ZN(n5503) );
  INV_X1 U6550 ( .A(n5500), .ZN(n5501) );
  NAND2_X1 U6551 ( .A1(n5501), .A2(SI_22_), .ZN(n5502) );
  NAND2_X1 U6552 ( .A1(n5503), .A2(n5502), .ZN(n6024) );
  INV_X1 U6553 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n5504) );
  INV_X1 U6554 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n8399) );
  MUX2_X1 U6555 ( .A(n5504), .B(n8399), .S(n5418), .Z(n5506) );
  INV_X1 U6556 ( .A(SI_23_), .ZN(n5505) );
  NAND2_X1 U6557 ( .A1(n5506), .A2(n5505), .ZN(n5510) );
  INV_X1 U6558 ( .A(n5506), .ZN(n5507) );
  NAND2_X1 U6559 ( .A1(n5507), .A2(SI_23_), .ZN(n5508) );
  NAND2_X1 U6560 ( .A1(n5510), .A2(n5508), .ZN(n5659) );
  INV_X1 U6561 ( .A(n5659), .ZN(n5509) );
  MUX2_X1 U6562 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(P2_DATAO_REG_24__SCAN_IN), 
        .S(n6238), .Z(n5512) );
  INV_X1 U6563 ( .A(SI_24_), .ZN(n5511) );
  XNOR2_X1 U6564 ( .A(n5512), .B(n5511), .ZN(n5647) );
  INV_X1 U6565 ( .A(n5647), .ZN(n5514) );
  NAND2_X1 U6566 ( .A1(n5512), .A2(SI_24_), .ZN(n5513) );
  INV_X1 U6567 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n8578) );
  INV_X1 U6568 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n8575) );
  MUX2_X1 U6569 ( .A(n8578), .B(n8575), .S(n5418), .Z(n5515) );
  INV_X1 U6570 ( .A(SI_25_), .ZN(n9689) );
  NAND2_X1 U6571 ( .A1(n5515), .A2(n9689), .ZN(n5518) );
  INV_X1 U6572 ( .A(n5515), .ZN(n5516) );
  NAND2_X1 U6573 ( .A1(n5516), .A2(SI_25_), .ZN(n5517) );
  NAND2_X1 U6574 ( .A1(n5518), .A2(n5517), .ZN(n6039) );
  INV_X1 U6575 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n8580) );
  INV_X1 U6576 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n8582) );
  MUX2_X1 U6577 ( .A(n8580), .B(n8582), .S(n6238), .Z(n5519) );
  INV_X1 U6578 ( .A(SI_26_), .ZN(n9687) );
  NAND2_X1 U6579 ( .A1(n5519), .A2(n9687), .ZN(n5522) );
  INV_X1 U6580 ( .A(n5519), .ZN(n5520) );
  NAND2_X1 U6581 ( .A1(n5520), .A2(SI_26_), .ZN(n5521) );
  NAND2_X1 U6582 ( .A1(n5523), .A2(n5522), .ZN(n5623) );
  INV_X1 U6583 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n9386) );
  INV_X1 U6584 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n10208) );
  MUX2_X1 U6585 ( .A(n9386), .B(n10208), .S(n5418), .Z(n5524) );
  INV_X1 U6586 ( .A(SI_27_), .ZN(n9593) );
  NAND2_X1 U6587 ( .A1(n5524), .A2(n9593), .ZN(n5527) );
  INV_X1 U6588 ( .A(n5524), .ZN(n5525) );
  NAND2_X1 U6589 ( .A1(n5525), .A2(SI_27_), .ZN(n5526) );
  NAND2_X1 U6590 ( .A1(n5623), .A2(n5622), .ZN(n5528) );
  NAND2_X1 U6591 ( .A1(n5528), .A2(n5527), .ZN(n5613) );
  MUX2_X1 U6592 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n6238), .Z(n5529) );
  INV_X1 U6593 ( .A(SI_28_), .ZN(n5530) );
  XNOR2_X1 U6594 ( .A(n5529), .B(n5530), .ZN(n5612) );
  NAND2_X1 U6595 ( .A1(n5613), .A2(n5612), .ZN(n5533) );
  INV_X1 U6596 ( .A(n5529), .ZN(n5531) );
  NAND2_X1 U6597 ( .A1(n5531), .A2(n5530), .ZN(n5532) );
  NAND2_X1 U6598 ( .A1(n5533), .A2(n5532), .ZN(n5584) );
  MUX2_X1 U6599 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .S(n5418), .Z(n5534) );
  INV_X1 U6600 ( .A(SI_29_), .ZN(n5535) );
  XNOR2_X1 U6601 ( .A(n5534), .B(n5535), .ZN(n5583) );
  INV_X1 U6602 ( .A(n5534), .ZN(n5536) );
  NAND2_X1 U6603 ( .A1(n5536), .A2(n5535), .ZN(n5537) );
  MUX2_X1 U6604 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .S(n6238), .Z(n5571) );
  INV_X1 U6605 ( .A(SI_30_), .ZN(n9682) );
  XNOR2_X1 U6606 ( .A(n5571), .B(n9682), .ZN(n5569) );
  NOR2_X1 U6607 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n5538) );
  INV_X1 U6608 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5540) );
  OAI21_X1 U6609 ( .B1(n5545), .B2(n5970), .A(P1_IR_REG_28__SCAN_IN), .ZN(
        n5543) );
  OAI21_X1 U6610 ( .B1(n5546), .B2(n5970), .A(P1_IR_REG_27__SCAN_IN), .ZN(
        n5549) );
  NAND2_X1 U6611 ( .A1(n8790), .A2(n6041), .ZN(n5554) );
  INV_X1 U6612 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8791) );
  OR2_X1 U6613 ( .A1(n5771), .A2(n8791), .ZN(n5553) );
  NAND2_X1 U6614 ( .A1(n5760), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n5565) );
  NAND2_X1 U6615 ( .A1(n6032), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n5564) );
  AND2_X2 U6616 ( .A1(n5562), .A2(n8825), .ZN(n5734) );
  NAND2_X1 U6617 ( .A1(n5734), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n5563) );
  NAND3_X1 U6618 ( .A1(n5565), .A2(n5564), .A3(n5563), .ZN(n9884) );
  INV_X1 U6619 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n9890) );
  NAND2_X1 U6620 ( .A1(n5956), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n5567) );
  NAND2_X1 U6621 ( .A1(n6031), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n5566) );
  OAI211_X1 U6622 ( .C1(n6050), .C2(n9890), .A(n5567), .B(n5566), .ZN(n9568)
         );
  NAND2_X1 U6623 ( .A1(n9884), .A2(n9568), .ZN(n5568) );
  NAND2_X1 U6624 ( .A1(n10067), .A2(n5568), .ZN(n6139) );
  INV_X1 U6625 ( .A(n5571), .ZN(n5572) );
  MUX2_X1 U6626 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n5418), .Z(n5574) );
  INV_X1 U6627 ( .A(SI_31_), .ZN(n5573) );
  XNOR2_X1 U6628 ( .A(n5574), .B(n5573), .ZN(n5575) );
  INV_X1 U6629 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n10197) );
  NOR2_X1 U6630 ( .A1(n5771), .A2(n10197), .ZN(n5577) );
  NAND2_X1 U6631 ( .A1(n5578), .A2(n6147), .ZN(n5581) );
  INV_X1 U6632 ( .A(n9884), .ZN(n5580) );
  NAND2_X1 U6633 ( .A1(n9882), .A2(n5580), .ZN(n6090) );
  INV_X1 U6634 ( .A(n9568), .ZN(n6087) );
  NAND2_X1 U6635 ( .A1(n8824), .A2(n6041), .ZN(n5587) );
  INV_X1 U6636 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n5585) );
  OR2_X1 U6637 ( .A1(n5771), .A2(n5585), .ZN(n5586) );
  INV_X1 U6638 ( .A(n10072), .ZN(n8805) );
  NAND3_X1 U6639 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n5797) );
  INV_X1 U6640 ( .A(n5797), .ZN(n5588) );
  NAND2_X1 U6641 ( .A1(n5588), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5813) );
  INV_X1 U6642 ( .A(n5813), .ZN(n5589) );
  NAND2_X1 U6643 ( .A1(n5589), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5827) );
  INV_X1 U6644 ( .A(n5827), .ZN(n5590) );
  NAND2_X1 U6645 ( .A1(n5590), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5829) );
  INV_X1 U6646 ( .A(n5883), .ZN(n5592) );
  NAND2_X1 U6647 ( .A1(n5592), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5901) );
  INV_X1 U6648 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5900) );
  INV_X1 U6649 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n9557) );
  NAND2_X1 U6650 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_REG3_REG_17__SCAN_IN), 
        .ZN(n5595) );
  INV_X1 U6651 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n9435) );
  INV_X1 U6652 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9513) );
  INV_X1 U6653 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n9447) );
  INV_X1 U6654 ( .A(n6046), .ZN(n5600) );
  NAND2_X1 U6655 ( .A1(n5600), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n5640) );
  INV_X1 U6656 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n5626) );
  INV_X1 U6657 ( .A(n5628), .ZN(n5601) );
  NAND2_X1 U6658 ( .A1(n5601), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n8802) );
  OR2_X1 U6659 ( .A1(n8802), .A2(n6035), .ZN(n5609) );
  INV_X1 U6660 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n5606) );
  NAND2_X1 U6661 ( .A1(n5760), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n5605) );
  NAND2_X1 U6662 ( .A1(n5734), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n5604) );
  OAI211_X1 U6663 ( .C1(n5606), .C2(n6050), .A(n5605), .B(n5604), .ZN(n5607)
         );
  INV_X1 U6664 ( .A(n5607), .ZN(n5608) );
  INV_X1 U6665 ( .A(n9899), .ZN(n9569) );
  NAND4_X1 U6666 ( .A1(n6139), .A2(n8805), .A3(n4850), .A4(n9569), .ZN(n5610)
         );
  INV_X1 U6667 ( .A(n5611), .ZN(n6067) );
  NAND4_X1 U6668 ( .A1(n6142), .A2(n9899), .A3(n7064), .A4(n10072), .ZN(n6066)
         );
  NAND2_X1 U6669 ( .A1(n6582), .A2(n6041), .ZN(n5615) );
  INV_X1 U6670 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n10203) );
  OR2_X1 U6671 ( .A1(n5771), .A2(n10203), .ZN(n5614) );
  INV_X1 U6672 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n8724) );
  NAND2_X1 U6673 ( .A1(n5628), .A2(n8724), .ZN(n5616) );
  NAND2_X1 U6674 ( .A1(n8802), .A2(n5616), .ZN(n9903) );
  INV_X1 U6675 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n9902) );
  NAND2_X1 U6676 ( .A1(n5760), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n5618) );
  NAND2_X1 U6677 ( .A1(n5734), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5617) );
  OAI211_X1 U6678 ( .C1(n9902), .C2(n6050), .A(n5618), .B(n5617), .ZN(n5619)
         );
  INV_X1 U6679 ( .A(n5619), .ZN(n5620) );
  NAND2_X1 U6680 ( .A1(n10076), .A2(n9396), .ZN(n8811) );
  INV_X1 U6681 ( .A(n6072), .ZN(n6181) );
  NAND2_X1 U6682 ( .A1(n10205), .A2(n6041), .ZN(n5625) );
  OR2_X1 U6683 ( .A1(n5771), .A2(n10208), .ZN(n5624) );
  NAND2_X1 U6684 ( .A1(n5640), .A2(n5626), .ZN(n5627) );
  NAND2_X1 U6685 ( .A1(n9393), .A2(n6047), .ZN(n5633) );
  INV_X1 U6686 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n7133) );
  NAND2_X1 U6687 ( .A1(n5760), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n5630) );
  NAND2_X1 U6688 ( .A1(n5734), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n5629) );
  OAI211_X1 U6689 ( .C1(n7133), .C2(n6050), .A(n5630), .B(n5629), .ZN(n5631)
         );
  INV_X1 U6690 ( .A(n5631), .ZN(n5632) );
  NAND2_X1 U6691 ( .A1(n10082), .A2(n9898), .ZN(n6136) );
  MUX2_X1 U6692 ( .A(n6136), .B(n6137), .S(n4850), .Z(n6061) );
  NAND2_X1 U6693 ( .A1(n8579), .A2(n6041), .ZN(n5637) );
  OR2_X1 U6694 ( .A1(n5771), .A2(n8582), .ZN(n5636) );
  INV_X1 U6695 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n5638) );
  NAND2_X1 U6696 ( .A1(n6046), .A2(n5638), .ZN(n5639) );
  NAND2_X1 U6697 ( .A1(n5640), .A2(n5639), .ZN(n8596) );
  INV_X1 U6698 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n5643) );
  NAND2_X1 U6699 ( .A1(n6031), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5642) );
  NAND2_X1 U6700 ( .A1(n5956), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n5641) );
  OAI211_X1 U6701 ( .C1(n5643), .C2(n6050), .A(n5642), .B(n5641), .ZN(n5644)
         );
  INV_X1 U6702 ( .A(n5644), .ZN(n5645) );
  NAND2_X1 U6703 ( .A1(n10086), .A2(n9451), .ZN(n7057) );
  OR2_X1 U6704 ( .A1(n10086), .A2(n9451), .ZN(n6134) );
  MUX2_X1 U6705 ( .A(n7057), .B(n6134), .S(n7064), .Z(n6059) );
  XNOR2_X1 U6706 ( .A(n5648), .B(n5647), .ZN(n8447) );
  NAND2_X1 U6707 ( .A1(n8447), .A2(n6041), .ZN(n5650) );
  INV_X1 U6708 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n8450) );
  OR2_X1 U6709 ( .A1(n5771), .A2(n8450), .ZN(n5649) );
  INV_X1 U6710 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n5651) );
  NAND2_X1 U6711 ( .A1(n5667), .A2(n5651), .ZN(n5652) );
  NAND2_X1 U6712 ( .A1(n6044), .A2(n5652), .ZN(n9938) );
  OR2_X1 U6713 ( .A1(n9938), .A2(n6035), .ZN(n5657) );
  INV_X1 U6714 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n9937) );
  NAND2_X1 U6715 ( .A1(n5956), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n5654) );
  NAND2_X1 U6716 ( .A1(n6031), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5653) );
  OAI211_X1 U6717 ( .C1(n9937), .C2(n6050), .A(n5654), .B(n5653), .ZN(n5655)
         );
  INV_X1 U6718 ( .A(n5655), .ZN(n5656) );
  NAND2_X1 U6719 ( .A1(n5660), .A2(n5659), .ZN(n5662) );
  NAND2_X1 U6720 ( .A1(n5662), .A2(n5661), .ZN(n8396) );
  NAND2_X1 U6721 ( .A1(n8396), .A2(n6041), .ZN(n5664) );
  OR2_X1 U6722 ( .A1(n5771), .A2(n8399), .ZN(n5663) );
  INV_X1 U6723 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n5665) );
  NAND2_X1 U6724 ( .A1(n6030), .A2(n5665), .ZN(n5666) );
  NAND2_X1 U6725 ( .A1(n5667), .A2(n5666), .ZN(n9948) );
  OR2_X1 U6726 ( .A1(n9948), .A2(n6035), .ZN(n5673) );
  INV_X1 U6727 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n5670) );
  NAND2_X1 U6728 ( .A1(n6031), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5669) );
  NAND2_X1 U6729 ( .A1(n5956), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n5668) );
  OAI211_X1 U6730 ( .C1(n5670), .C2(n6050), .A(n5669), .B(n5668), .ZN(n5671)
         );
  INV_X1 U6731 ( .A(n5671), .ZN(n5672) );
  NAND2_X1 U6732 ( .A1(n5673), .A2(n5672), .ZN(n9969) );
  INV_X1 U6733 ( .A(n9969), .ZN(n8681) );
  NAND2_X1 U6734 ( .A1(n7054), .A2(n7052), .ZN(n6119) );
  NAND2_X1 U6735 ( .A1(n10097), .A2(n9448), .ZN(n6131) );
  AND2_X1 U6736 ( .A1(n10102), .A2(n8681), .ZN(n7053) );
  INV_X1 U6737 ( .A(n7053), .ZN(n5674) );
  NAND2_X1 U6738 ( .A1(n6131), .A2(n5674), .ZN(n5675) );
  MUX2_X1 U6739 ( .A(n6119), .B(n5675), .S(n7064), .Z(n6056) );
  XNOR2_X1 U6740 ( .A(n5677), .B(n5676), .ZN(n8183) );
  NAND2_X1 U6741 ( .A1(n8183), .A2(n6041), .ZN(n5679) );
  OR2_X1 U6742 ( .A1(n5771), .A2(n8184), .ZN(n5678) );
  NAND2_X1 U6743 ( .A1(n5690), .A2(n9435), .ZN(n5680) );
  NAND2_X1 U6744 ( .A1(n6028), .A2(n5680), .ZN(n9986) );
  OR2_X1 U6745 ( .A1(n9986), .A2(n6035), .ZN(n5683) );
  AOI22_X1 U6746 ( .A1(n6032), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n5760), .B2(
        P1_REG1_REG_21__SCAN_IN), .ZN(n5682) );
  NAND2_X1 U6747 ( .A1(n5734), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5681) );
  OR2_X1 U6748 ( .A1(n10113), .A2(n10000), .ZN(n6021) );
  XNOR2_X1 U6749 ( .A(n5685), .B(n5684), .ZN(n8164) );
  NAND2_X1 U6750 ( .A1(n8164), .A2(n6041), .ZN(n5687) );
  OR2_X1 U6751 ( .A1(n5771), .A2(n8165), .ZN(n5686) );
  INV_X1 U6752 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n5688) );
  NAND2_X1 U6753 ( .A1(n6014), .A2(n5688), .ZN(n5689) );
  NAND2_X1 U6754 ( .A1(n5690), .A2(n5689), .ZN(n10006) );
  INV_X1 U6755 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n10007) );
  OAI22_X1 U6756 ( .A1(n10006), .A2(n6035), .B1(n6050), .B2(n10007), .ZN(n5695) );
  INV_X1 U6757 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n5693) );
  NAND2_X1 U6758 ( .A1(n6031), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n5691) );
  OAI21_X1 U6759 ( .B1(n5693), .B2(n5692), .A(n5691), .ZN(n5694) );
  INV_X1 U6760 ( .A(n10022), .ZN(n9436) );
  OR2_X1 U6761 ( .A1(n10117), .A2(n9436), .ZN(n9981) );
  AND2_X1 U6762 ( .A1(n6021), .A2(n9981), .ZN(n7046) );
  NAND2_X1 U6763 ( .A1(n10113), .A2(n10000), .ZN(n7047) );
  INV_X1 U6764 ( .A(n7047), .ZN(n5696) );
  OR2_X1 U6765 ( .A1(n7046), .A2(n5696), .ZN(n5700) );
  NAND2_X1 U6766 ( .A1(n10117), .A2(n9436), .ZN(n5697) );
  NAND2_X1 U6767 ( .A1(n7047), .A2(n5697), .ZN(n5698) );
  AND2_X1 U6768 ( .A1(n5698), .A2(n6021), .ZN(n6093) );
  INV_X1 U6769 ( .A(n6093), .ZN(n5699) );
  MUX2_X1 U6770 ( .A(n5700), .B(n5699), .S(n7064), .Z(n6037) );
  XNOR2_X1 U6771 ( .A(n5701), .B(n5389), .ZN(n7255) );
  NAND2_X1 U6772 ( .A1(n7255), .A2(n6041), .ZN(n5709) );
  NAND2_X1 U6773 ( .A1(n5754), .A2(n5790), .ZN(n5703) );
  INV_X1 U6774 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5704) );
  NAND2_X1 U6775 ( .A1(n5819), .A2(n5820), .ZN(n5844) );
  NAND2_X1 U6776 ( .A1(n5844), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5836) );
  INV_X1 U6777 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5705) );
  NAND2_X1 U6778 ( .A1(n5836), .A2(n5705), .ZN(n5706) );
  NAND2_X1 U6779 ( .A1(n5706), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5707) );
  XNOR2_X1 U6780 ( .A(n5707), .B(P1_IR_REG_9__SCAN_IN), .ZN(n10281) );
  AOI22_X1 U6781 ( .A1(n6008), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n6007), .B2(
        n10281), .ZN(n5708) );
  NAND2_X1 U6782 ( .A1(n5709), .A2(n5708), .ZN(n10580) );
  NAND2_X1 U6783 ( .A1(n6031), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5715) );
  NAND2_X1 U6784 ( .A1(n5956), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5714) );
  NAND2_X1 U6785 ( .A1(n5829), .A2(n5710), .ZN(n5711) );
  AND2_X1 U6786 ( .A1(n5852), .A2(n5711), .ZN(n8158) );
  NAND2_X1 U6787 ( .A1(n6047), .A2(n8158), .ZN(n5713) );
  NAND2_X1 U6788 ( .A1(n6032), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5712) );
  NAND4_X1 U6789 ( .A1(n5715), .A2(n5714), .A3(n5713), .A4(n5712), .ZN(n10538)
         );
  INV_X1 U6790 ( .A(n10538), .ZN(n8107) );
  NAND2_X1 U6791 ( .A1(n10580), .A2(n8107), .ZN(n7028) );
  NAND2_X1 U6792 ( .A1(n5762), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5718) );
  NAND2_X1 U6793 ( .A1(n5760), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5717) );
  NAND2_X1 U6794 ( .A1(n5734), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5716) );
  XNOR2_X1 U6795 ( .A(n5721), .B(n5720), .ZN(n7237) );
  INV_X1 U6796 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n7238) );
  INV_X1 U6797 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n5723) );
  NAND2_X1 U6798 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5722) );
  XNOR2_X1 U6799 ( .A(n5723), .B(n5722), .ZN(n7323) );
  NAND2_X1 U6800 ( .A1(n5762), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5727) );
  NAND2_X1 U6801 ( .A1(n5734), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5726) );
  NAND2_X1 U6802 ( .A1(n5760), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5724) );
  INV_X1 U6803 ( .A(SI_0_), .ZN(n5729) );
  INV_X1 U6804 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5728) );
  OAI21_X1 U6805 ( .B1(n5021), .B2(n5729), .A(n5728), .ZN(n5731) );
  AND2_X1 U6806 ( .A1(n5731), .A2(n5730), .ZN(n10210) );
  MUX2_X1 U6807 ( .A(P1_IR_REG_0__SCAN_IN), .B(n10210), .S(n5745), .Z(n7629)
         );
  INV_X1 U6808 ( .A(n7629), .ZN(n7759) );
  NOR2_X1 U6809 ( .A1(n7380), .A2(n7759), .ZN(n7761) );
  NAND2_X1 U6810 ( .A1(n6077), .A2(n7761), .ZN(n7760) );
  INV_X1 U6811 ( .A(n7491), .ZN(n5732) );
  NAND2_X1 U6812 ( .A1(n5732), .A2(n7766), .ZN(n5733) );
  NAND2_X1 U6813 ( .A1(n7760), .A2(n5733), .ZN(n7665) );
  NAND2_X1 U6814 ( .A1(n5760), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5738) );
  NAND2_X1 U6815 ( .A1(n5734), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5737) );
  NAND2_X1 U6816 ( .A1(n5762), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5736) );
  NAND2_X1 U6817 ( .A1(n5763), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5735) );
  INV_X1 U6818 ( .A(n7763), .ZN(n7512) );
  XNOR2_X1 U6819 ( .A(n5739), .B(n5740), .ZN(n7234) );
  INV_X1 U6820 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n5746) );
  NOR2_X1 U6821 ( .A1(n5741), .A2(n5970), .ZN(n5742) );
  MUX2_X1 U6822 ( .A(n5970), .B(n5742), .S(P1_IR_REG_2__SCAN_IN), .Z(n5743) );
  INV_X1 U6823 ( .A(n5743), .ZN(n5744) );
  NAND2_X1 U6824 ( .A1(n5744), .A2(n5702), .ZN(n7460) );
  INV_X1 U6825 ( .A(n7087), .ZN(n7666) );
  NAND2_X1 U6826 ( .A1(n7665), .A2(n7666), .ZN(n7664) );
  NAND2_X1 U6827 ( .A1(n5760), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5751) );
  NAND2_X1 U6828 ( .A1(n5734), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5750) );
  INV_X1 U6829 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n5747) );
  XNOR2_X1 U6830 ( .A(n5747), .B(P1_REG3_REG_3__SCAN_IN), .ZN(n10421) );
  NAND2_X1 U6831 ( .A1(n5762), .A2(n10421), .ZN(n5749) );
  NAND2_X1 U6832 ( .A1(n5763), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5748) );
  AND2_X1 U6833 ( .A1(n5752), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5753) );
  NAND2_X1 U6834 ( .A1(n5753), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n5756) );
  INV_X1 U6835 ( .A(n5753), .ZN(n5755) );
  NAND2_X1 U6836 ( .A1(n5755), .A2(n5754), .ZN(n5789) );
  NAND2_X1 U6837 ( .A1(n5756), .A2(n5789), .ZN(n7304) );
  XNOR2_X1 U6838 ( .A(n5757), .B(n5098), .ZN(n6279) );
  INV_X1 U6839 ( .A(n6279), .ZN(n7230) );
  OR2_X1 U6840 ( .A1(n5774), .A2(n7230), .ZN(n5759) );
  OR2_X1 U6841 ( .A1(n5771), .A2(n4986), .ZN(n5758) );
  OAI211_X1 U6842 ( .C1(n5745), .C2(n7304), .A(n5759), .B(n5758), .ZN(n9496)
         );
  NAND2_X1 U6843 ( .A1(n7364), .A2(n10423), .ZN(n6076) );
  NAND2_X1 U6844 ( .A1(n5734), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5768) );
  NAND2_X1 U6845 ( .A1(n5760), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5766) );
  INV_X1 U6846 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n5761) );
  NAND2_X1 U6847 ( .A1(n5762), .A2(n5761), .ZN(n5765) );
  NAND2_X1 U6848 ( .A1(n5763), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5764) );
  NAND2_X1 U6849 ( .A1(n5702), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5770) );
  INV_X1 U6850 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5769) );
  XNOR2_X1 U6851 ( .A(n5770), .B(n5769), .ZN(n7300) );
  INV_X1 U6852 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n7236) );
  OR2_X1 U6853 ( .A1(n5771), .A2(n7236), .ZN(n5776) );
  XNOR2_X1 U6854 ( .A(n5773), .B(n5772), .ZN(n7235) );
  OR2_X1 U6855 ( .A1(n5774), .A2(n7235), .ZN(n5775) );
  OAI211_X1 U6856 ( .C1(n5745), .C2(n7300), .A(n5776), .B(n5775), .ZN(n7753)
         );
  NAND2_X1 U6857 ( .A1(n5777), .A2(n7633), .ZN(n6075) );
  NAND2_X1 U6858 ( .A1(n6076), .A2(n6075), .ZN(n6157) );
  INV_X1 U6859 ( .A(n10407), .ZN(n5779) );
  NAND2_X1 U6860 ( .A1(n7794), .A2(n9496), .ZN(n6159) );
  INV_X1 U6861 ( .A(n6159), .ZN(n5778) );
  OAI21_X1 U6862 ( .B1(n5779), .B2(n5778), .A(n6076), .ZN(n5780) );
  NAND2_X1 U6863 ( .A1(n5734), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5788) );
  NAND2_X1 U6864 ( .A1(n5760), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5787) );
  INV_X1 U6865 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5783) );
  NAND2_X1 U6866 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n5782) );
  NAND2_X1 U6867 ( .A1(n5783), .A2(n5782), .ZN(n5784) );
  AND2_X1 U6868 ( .A1(n5797), .A2(n5784), .ZN(n7998) );
  NAND2_X1 U6869 ( .A1(n6047), .A2(n7998), .ZN(n5786) );
  NAND2_X1 U6870 ( .A1(n6032), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5785) );
  NAND2_X1 U6871 ( .A1(n5789), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5791) );
  XNOR2_X1 U6872 ( .A(n5791), .B(n5790), .ZN(n7307) );
  XNOR2_X1 U6873 ( .A(n5792), .B(n5793), .ZN(n7244) );
  OR2_X1 U6874 ( .A1(n5774), .A2(n7244), .ZN(n5795) );
  INV_X1 U6875 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n7243) );
  OR2_X1 U6876 ( .A1(n5771), .A2(n7243), .ZN(n5794) );
  NAND2_X1 U6877 ( .A1(n10491), .A2(n7997), .ZN(n10483) );
  MUX2_X1 U6878 ( .A(n10485), .B(n10483), .S(n4850), .Z(n5810) );
  NAND2_X1 U6879 ( .A1(n5956), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5802) );
  NAND2_X1 U6880 ( .A1(n6031), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5801) );
  INV_X1 U6881 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n5796) );
  NAND2_X1 U6882 ( .A1(n5797), .A2(n5796), .ZN(n5798) );
  AND2_X1 U6883 ( .A1(n5813), .A2(n5798), .ZN(n10506) );
  NAND2_X1 U6884 ( .A1(n6047), .A2(n10506), .ZN(n5800) );
  NAND2_X1 U6885 ( .A1(n6032), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5799) );
  NOR2_X1 U6886 ( .A1(n5803), .A2(n5970), .ZN(n5804) );
  MUX2_X1 U6887 ( .A(n5970), .B(n5804), .S(P1_IR_REG_6__SCAN_IN), .Z(n5805) );
  OR2_X1 U6888 ( .A1(n5805), .A2(n5819), .ZN(n7338) );
  XNOR2_X1 U6889 ( .A(n5807), .B(n5806), .ZN(n7239) );
  NAND2_X1 U6890 ( .A1(n6041), .A2(n7239), .ZN(n5809) );
  INV_X1 U6891 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n7241) );
  OR2_X1 U6892 ( .A1(n5771), .A2(n7241), .ZN(n5808) );
  OAI211_X1 U6893 ( .C1(n5745), .C2(n7338), .A(n5809), .B(n5808), .ZN(n7929)
         );
  NAND2_X1 U6894 ( .A1(n8011), .A2(n7929), .ZN(n6162) );
  INV_X1 U6895 ( .A(n8011), .ZN(n7994) );
  NAND2_X1 U6896 ( .A1(n7994), .A2(n10502), .ZN(n6160) );
  AND2_X1 U6897 ( .A1(n6162), .A2(n6160), .ZN(n10487) );
  NAND2_X1 U6898 ( .A1(n5810), .A2(n10487), .ZN(n5811) );
  NAND2_X1 U6899 ( .A1(n5734), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5818) );
  NAND2_X1 U6900 ( .A1(n5956), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5817) );
  INV_X1 U6901 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5812) );
  NAND2_X1 U6902 ( .A1(n5813), .A2(n5812), .ZN(n5814) );
  AND2_X1 U6903 ( .A1(n5827), .A2(n5814), .ZN(n8015) );
  NAND2_X1 U6904 ( .A1(n6047), .A2(n8015), .ZN(n5816) );
  NAND2_X1 U6905 ( .A1(n6032), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5815) );
  INV_X1 U6906 ( .A(n10490), .ZN(n10541) );
  OR2_X1 U6907 ( .A1(n5819), .A2(n5970), .ZN(n5821) );
  XNOR2_X1 U6908 ( .A(n5821), .B(n5820), .ZN(n7359) );
  OR2_X1 U6909 ( .A1(n7247), .A2(n5774), .ZN(n5825) );
  OR2_X1 U6910 ( .A1(n5771), .A2(n7246), .ZN(n5824) );
  OAI211_X1 U6911 ( .C1(n4854), .C2(n7359), .A(n5825), .B(n5824), .ZN(n7914)
         );
  NAND2_X1 U6912 ( .A1(n10541), .A2(n10518), .ZN(n6163) );
  NAND2_X1 U6913 ( .A1(n6163), .A2(n6160), .ZN(n6129) );
  NAND2_X1 U6914 ( .A1(n10490), .A2(n7914), .ZN(n10542) );
  NAND2_X1 U6915 ( .A1(n10542), .A2(n6162), .ZN(n5826) );
  MUX2_X1 U6916 ( .A(n6129), .B(n5826), .S(n7064), .Z(n5840) );
  NAND2_X1 U6917 ( .A1(n6031), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5833) );
  NAND2_X1 U6918 ( .A1(n5956), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5832) );
  INV_X1 U6919 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n7334) );
  NAND2_X1 U6920 ( .A1(n5827), .A2(n7334), .ZN(n5828) );
  AND2_X1 U6921 ( .A1(n5829), .A2(n5828), .ZN(n10562) );
  NAND2_X1 U6922 ( .A1(n6047), .A2(n10562), .ZN(n5831) );
  NAND2_X1 U6923 ( .A1(n6032), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5830) );
  XNOR2_X1 U6924 ( .A(n5835), .B(n5834), .ZN(n7251) );
  NAND2_X1 U6925 ( .A1(n7251), .A2(n6041), .ZN(n5838) );
  XNOR2_X1 U6926 ( .A(n5836), .B(P1_IR_REG_8__SCAN_IN), .ZN(n7341) );
  AOI22_X1 U6927 ( .A1(n6008), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n6007), .B2(
        n7341), .ZN(n5837) );
  NAND2_X1 U6928 ( .A1(n5838), .A2(n5837), .ZN(n8109) );
  NAND2_X1 U6929 ( .A1(n8098), .A2(n8109), .ZN(n7025) );
  INV_X1 U6930 ( .A(n8109), .ZN(n10566) );
  INV_X1 U6931 ( .A(n8098), .ZN(n9790) );
  NAND2_X1 U6932 ( .A1(n10566), .A2(n9790), .ZN(n8076) );
  MUX2_X1 U6933 ( .A(n6163), .B(n10542), .S(n4850), .Z(n5839) );
  MUX2_X1 U6934 ( .A(n8076), .B(n7025), .S(n7064), .Z(n5841) );
  OR2_X1 U6935 ( .A1(n10580), .A2(n8107), .ZN(n6098) );
  MUX2_X1 U6936 ( .A(n4850), .B(n5842), .S(n6098), .Z(n5858) );
  XNOR2_X1 U6937 ( .A(n5843), .B(n5390), .ZN(n7290) );
  NAND2_X1 U6938 ( .A1(n7290), .A2(n6041), .ZN(n5850) );
  NAND2_X1 U6939 ( .A1(n5846), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5845) );
  MUX2_X1 U6940 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5845), .S(
        P1_IR_REG_10__SCAN_IN), .Z(n5848) );
  INV_X1 U6941 ( .A(n5876), .ZN(n5847) );
  NAND2_X1 U6942 ( .A1(n5848), .A2(n5847), .ZN(n7579) );
  INV_X1 U6943 ( .A(n7579), .ZN(n10293) );
  AOI22_X1 U6944 ( .A1(n6008), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6007), .B2(
        n10293), .ZN(n5849) );
  NAND2_X1 U6945 ( .A1(n5850), .A2(n5849), .ZN(n8276) );
  NAND2_X1 U6946 ( .A1(n5956), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5857) );
  NAND2_X1 U6947 ( .A1(n6032), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5856) );
  NAND2_X1 U6948 ( .A1(n5852), .A2(n5851), .ZN(n5853) );
  AND2_X1 U6949 ( .A1(n5865), .A2(n5853), .ZN(n8270) );
  NAND2_X1 U6950 ( .A1(n6047), .A2(n8270), .ZN(n5855) );
  NAND2_X1 U6951 ( .A1(n6031), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5854) );
  OR2_X1 U6952 ( .A1(n8276), .A2(n8267), .ZN(n6100) );
  NAND2_X1 U6953 ( .A1(n8276), .A2(n8267), .ZN(n7030) );
  OAI211_X1 U6954 ( .C1(n7064), .C2(n7028), .A(n5858), .B(n8192), .ZN(n5872)
         );
  XNOR2_X1 U6955 ( .A(n5859), .B(n5860), .ZN(n7260) );
  NAND2_X1 U6956 ( .A1(n7260), .A2(n6041), .ZN(n5863) );
  INV_X1 U6957 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5970) );
  OR2_X1 U6958 ( .A1(n5876), .A2(n5970), .ZN(n5861) );
  XNOR2_X1 U6959 ( .A(n5861), .B(P1_IR_REG_11__SCAN_IN), .ZN(n7711) );
  AOI22_X1 U6960 ( .A1(n6008), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n6007), .B2(
        n7711), .ZN(n5862) );
  NAND2_X1 U6961 ( .A1(n5863), .A2(n5862), .ZN(n10168) );
  NAND2_X1 U6962 ( .A1(n6031), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5870) );
  NAND2_X1 U6963 ( .A1(n5956), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5869) );
  INV_X1 U6964 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5864) );
  NAND2_X1 U6965 ( .A1(n5865), .A2(n5864), .ZN(n5866) );
  AND2_X1 U6966 ( .A1(n5883), .A2(n5866), .ZN(n8334) );
  NAND2_X1 U6967 ( .A1(n6047), .A2(n8334), .ZN(n5868) );
  NAND2_X1 U6968 ( .A1(n6032), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5867) );
  OR2_X1 U6969 ( .A1(n10168), .A2(n8363), .ZN(n6102) );
  NAND2_X1 U6970 ( .A1(n10168), .A2(n8363), .ZN(n7032) );
  MUX2_X1 U6971 ( .A(n6100), .B(n7030), .S(n7064), .Z(n5871) );
  NAND2_X1 U6972 ( .A1(n4891), .A2(SI_12_), .ZN(n5873) );
  NAND2_X1 U6973 ( .A1(n5874), .A2(n5873), .ZN(n7422) );
  NAND2_X1 U6974 ( .A1(n7422), .A2(n6041), .ZN(n5882) );
  INV_X1 U6975 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n5875) );
  INV_X1 U6976 ( .A(n5879), .ZN(n5877) );
  NAND2_X1 U6977 ( .A1(n5877), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n5880) );
  INV_X1 U6978 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5878) );
  NAND2_X1 U6979 ( .A1(n5879), .A2(n5878), .ZN(n5896) );
  AOI22_X1 U6980 ( .A1(n6008), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n6007), .B2(
        n7836), .ZN(n5881) );
  NAND2_X1 U6981 ( .A1(n5956), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5888) );
  NAND2_X1 U6982 ( .A1(n6031), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5887) );
  INV_X1 U6983 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n7719) );
  NAND2_X1 U6984 ( .A1(n5883), .A2(n7719), .ZN(n5884) );
  AND2_X1 U6985 ( .A1(n5901), .A2(n5884), .ZN(n8359) );
  NAND2_X1 U6986 ( .A1(n6047), .A2(n8359), .ZN(n5886) );
  NAND2_X1 U6987 ( .A1(n6032), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5885) );
  OR2_X1 U6988 ( .A1(n10163), .A2(n8486), .ZN(n6103) );
  NAND2_X1 U6989 ( .A1(n10163), .A2(n8486), .ZN(n7033) );
  MUX2_X1 U6990 ( .A(n7032), .B(n6102), .S(n7064), .Z(n5889) );
  AND2_X1 U6991 ( .A1(n8295), .A2(n5889), .ZN(n5890) );
  INV_X1 U6992 ( .A(n5891), .ZN(n5893) );
  NAND2_X1 U6993 ( .A1(n5893), .A2(n5892), .ZN(n5895) );
  NAND2_X1 U6994 ( .A1(n5895), .A2(n5894), .ZN(n7547) );
  NAND2_X1 U6995 ( .A1(n7547), .A2(n6041), .ZN(n5899) );
  NAND2_X1 U6996 ( .A1(n5896), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5897) );
  XNOR2_X1 U6997 ( .A(n5897), .B(P1_IR_REG_13__SCAN_IN), .ZN(n8038) );
  AOI22_X1 U6998 ( .A1(n6008), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n6007), .B2(
        n8038), .ZN(n5898) );
  NAND2_X1 U6999 ( .A1(n6031), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5906) );
  NAND2_X1 U7000 ( .A1(n5956), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5905) );
  NAND2_X1 U7001 ( .A1(n5901), .A2(n5900), .ZN(n5902) );
  AND2_X1 U7002 ( .A1(n5919), .A2(n5902), .ZN(n8488) );
  NAND2_X1 U7003 ( .A1(n6047), .A2(n8488), .ZN(n5904) );
  NAND2_X1 U7004 ( .A1(n6032), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5903) );
  NAND2_X1 U7005 ( .A1(n10157), .A2(n8472), .ZN(n7035) );
  INV_X1 U7006 ( .A(n7035), .ZN(n5947) );
  AOI21_X1 U7007 ( .B1(n5925), .B2(n6103), .A(n5947), .ZN(n5932) );
  XNOR2_X1 U7008 ( .A(n5908), .B(n5907), .ZN(n7680) );
  NAND2_X1 U7009 ( .A1(n7680), .A2(n6041), .ZN(n5917) );
  NOR2_X1 U7010 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n5909) );
  NOR2_X1 U7011 ( .A1(n5914), .A2(n5970), .ZN(n5911) );
  MUX2_X1 U7012 ( .A(n5970), .B(n5911), .S(P1_IR_REG_14__SCAN_IN), .Z(n5912)
         );
  INV_X1 U7013 ( .A(n5912), .ZN(n5915) );
  INV_X1 U7014 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5913) );
  NAND2_X1 U7015 ( .A1(n5914), .A2(n5913), .ZN(n5952) );
  AOI22_X1 U7016 ( .A1(n6008), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n9798), .B2(
        n6007), .ZN(n5916) );
  NAND2_X1 U7017 ( .A1(n5956), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5924) );
  NAND2_X1 U7018 ( .A1(n6031), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5923) );
  INV_X1 U7019 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n5918) );
  NAND2_X1 U7020 ( .A1(n5919), .A2(n5918), .ZN(n5920) );
  AND2_X1 U7021 ( .A1(n5941), .A2(n5920), .ZN(n9410) );
  NAND2_X1 U7022 ( .A1(n6047), .A2(n9410), .ZN(n5922) );
  NAND2_X1 U7023 ( .A1(n6032), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5921) );
  NAND4_X1 U7024 ( .A1(n5924), .A2(n5923), .A3(n5922), .A4(n5921), .ZN(n9786)
         );
  INV_X1 U7025 ( .A(n9786), .ZN(n8525) );
  OR2_X1 U7026 ( .A1(n10157), .A2(n8472), .ZN(n6106) );
  NAND3_X1 U7027 ( .A1(n7037), .A2(n4850), .A3(n6106), .ZN(n5931) );
  NAND2_X1 U7028 ( .A1(n10152), .A2(n8525), .ZN(n6097) );
  NAND3_X1 U7029 ( .A1(n5926), .A2(n6097), .A3(n7064), .ZN(n5930) );
  AND2_X1 U7030 ( .A1(n9786), .A2(n7064), .ZN(n5928) );
  OAI21_X1 U7031 ( .B1(n9786), .B2(n7064), .A(n10152), .ZN(n5927) );
  OAI21_X1 U7032 ( .B1(n5928), .B2(n10152), .A(n5927), .ZN(n5929) );
  OAI211_X1 U7033 ( .C1(n5932), .C2(n5931), .A(n5930), .B(n5929), .ZN(n5949)
         );
  INV_X1 U7034 ( .A(n5933), .ZN(n5935) );
  NAND2_X1 U7035 ( .A1(n5935), .A2(n5934), .ZN(n5936) );
  NAND2_X1 U7036 ( .A1(n5937), .A2(n5936), .ZN(n7818) );
  NAND2_X1 U7037 ( .A1(n7818), .A2(n6041), .ZN(n5940) );
  NAND2_X1 U7038 ( .A1(n5952), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5938) );
  XNOR2_X1 U7039 ( .A(n5938), .B(P1_IR_REG_15__SCAN_IN), .ZN(n9810) );
  AOI22_X1 U7040 ( .A1(n6008), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n6007), .B2(
        n9810), .ZN(n5939) );
  NAND2_X1 U7041 ( .A1(n6031), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5946) );
  NAND2_X1 U7042 ( .A1(n5956), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5945) );
  NAND2_X1 U7043 ( .A1(n5941), .A2(n9557), .ZN(n5942) );
  AND2_X1 U7044 ( .A1(n5957), .A2(n5942), .ZN(n9555) );
  NAND2_X1 U7045 ( .A1(n6047), .A2(n9555), .ZN(n5944) );
  NAND2_X1 U7046 ( .A1(n6032), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n5943) );
  NAND2_X1 U7047 ( .A1(n10146), .A2(n9465), .ZN(n7039) );
  NAND3_X1 U7048 ( .A1(n7037), .A2(n5947), .A3(n7064), .ZN(n5948) );
  NAND3_X1 U7049 ( .A1(n5949), .A2(n8518), .A3(n5948), .ZN(n5967) );
  XNOR2_X1 U7050 ( .A(n5951), .B(n5950), .ZN(n7846) );
  NAND2_X1 U7051 ( .A1(n7846), .A2(n6041), .ZN(n5955) );
  NAND2_X1 U7052 ( .A1(n5953), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5972) );
  XNOR2_X1 U7053 ( .A(n5972), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9840) );
  AOI22_X1 U7054 ( .A1(n6008), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n9840), .B2(
        n6007), .ZN(n5954) );
  NAND2_X1 U7055 ( .A1(n5956), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n5962) );
  NAND2_X1 U7056 ( .A1(n6032), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n5961) );
  INV_X1 U7057 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n9815) );
  NAND2_X1 U7058 ( .A1(n5957), .A2(n9815), .ZN(n5958) );
  AND2_X1 U7059 ( .A1(n5998), .A2(n5958), .ZN(n9462) );
  NAND2_X1 U7060 ( .A1(n6047), .A2(n9462), .ZN(n5960) );
  NAND2_X1 U7061 ( .A1(n6031), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5959) );
  NAND2_X1 U7062 ( .A1(n10141), .A2(n9562), .ZN(n7040) );
  NAND2_X1 U7063 ( .A1(n7041), .A2(n7040), .ZN(n8556) );
  INV_X1 U7064 ( .A(n7039), .ZN(n5964) );
  INV_X1 U7065 ( .A(n6109), .ZN(n5963) );
  MUX2_X1 U7066 ( .A(n5964), .B(n5963), .S(n7064), .Z(n5965) );
  NOR2_X1 U7067 ( .A1(n8556), .A2(n5965), .ZN(n5966) );
  NAND2_X1 U7068 ( .A1(n5967), .A2(n5966), .ZN(n5985) );
  NAND2_X1 U7069 ( .A1(n5985), .A2(n7041), .ZN(n5984) );
  XNOR2_X1 U7070 ( .A(n5969), .B(n5968), .ZN(n7888) );
  NAND2_X1 U7071 ( .A1(n7888), .A2(n6041), .ZN(n5978) );
  INV_X1 U7072 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5971) );
  AOI21_X1 U7073 ( .B1(n5972), .B2(n5971), .A(n5970), .ZN(n5973) );
  NAND2_X1 U7074 ( .A1(n5973), .A2(P1_IR_REG_17__SCAN_IN), .ZN(n5976) );
  INV_X1 U7075 ( .A(n5973), .ZN(n5975) );
  INV_X1 U7076 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5974) );
  NAND2_X1 U7077 ( .A1(n5975), .A2(n5974), .ZN(n5992) );
  AOI22_X1 U7078 ( .A1(n9849), .A2(n6007), .B1(n6008), .B2(
        P2_DATAO_REG_17__SCAN_IN), .ZN(n5977) );
  NAND2_X1 U7079 ( .A1(n5956), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n5982) );
  NAND2_X1 U7080 ( .A1(n6032), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n5981) );
  XNOR2_X1 U7081 ( .A(n5998), .B(P1_REG3_REG_17__SCAN_IN), .ZN(n10060) );
  NAND2_X1 U7082 ( .A1(n6047), .A2(n10060), .ZN(n5980) );
  NAND2_X1 U7083 ( .A1(n6031), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5979) );
  NAND4_X1 U7084 ( .A1(n5982), .A2(n5981), .A3(n5980), .A4(n5979), .ZN(n9573)
         );
  INV_X1 U7085 ( .A(n9573), .ZN(n10035) );
  NAND2_X1 U7086 ( .A1(n10135), .A2(n10035), .ZN(n6095) );
  INV_X1 U7087 ( .A(n7043), .ZN(n5983) );
  AOI21_X1 U7088 ( .B1(n5984), .B2(n10050), .A(n5983), .ZN(n5989) );
  NAND2_X1 U7089 ( .A1(n5985), .A2(n7040), .ZN(n5987) );
  INV_X1 U7090 ( .A(n6095), .ZN(n5986) );
  AOI21_X1 U7091 ( .B1(n5987), .B2(n10050), .A(n5986), .ZN(n5988) );
  XNOR2_X1 U7092 ( .A(n5991), .B(n5990), .ZN(n8003) );
  NAND2_X1 U7093 ( .A1(n8003), .A2(n6041), .ZN(n5995) );
  NAND2_X1 U7094 ( .A1(n5992), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5993) );
  XNOR2_X1 U7095 ( .A(n5993), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9872) );
  AOI22_X1 U7096 ( .A1(n9872), .A2(n6007), .B1(n6008), .B2(
        P2_DATAO_REG_18__SCAN_IN), .ZN(n5994) );
  NAND2_X1 U7097 ( .A1(n6031), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n6003) );
  NAND2_X1 U7098 ( .A1(n5956), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n6002) );
  INV_X1 U7099 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n5997) );
  INV_X1 U7100 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n5996) );
  OAI21_X1 U7101 ( .B1(n5998), .B2(n5997), .A(n5996), .ZN(n5999) );
  AND2_X1 U7102 ( .A1(n5999), .A2(n6012), .ZN(n10041) );
  NAND2_X1 U7103 ( .A1(n6047), .A2(n10041), .ZN(n6001) );
  NAND2_X1 U7104 ( .A1(n6032), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n6000) );
  OR2_X1 U7105 ( .A1(n10043), .A2(n9474), .ZN(n6111) );
  NAND2_X1 U7106 ( .A1(n10043), .A2(n9474), .ZN(n7044) );
  INV_X1 U7107 ( .A(n10032), .ZN(n10030) );
  NAND2_X1 U7108 ( .A1(n4890), .A2(n6004), .ZN(n6005) );
  NAND2_X1 U7109 ( .A1(n6006), .A2(n6005), .ZN(n8112) );
  NAND2_X1 U7110 ( .A1(n8112), .A2(n6041), .ZN(n6010) );
  AOI22_X1 U7111 ( .A1(n6008), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9991), .B2(
        n6007), .ZN(n6009) );
  NAND2_X1 U7112 ( .A1(n5956), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n6018) );
  NAND2_X1 U7113 ( .A1(n6032), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n6017) );
  INV_X1 U7114 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n6011) );
  NAND2_X1 U7115 ( .A1(n6012), .A2(n6011), .ZN(n6013) );
  AND2_X1 U7116 ( .A1(n6014), .A2(n6013), .ZN(n10016) );
  NAND2_X1 U7117 ( .A1(n6047), .A2(n10016), .ZN(n6016) );
  NAND2_X1 U7118 ( .A1(n6031), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n6015) );
  NAND4_X1 U7119 ( .A1(n6018), .A2(n6017), .A3(n6016), .A4(n6015), .ZN(n9572)
         );
  INV_X1 U7120 ( .A(n9572), .ZN(n10036) );
  OR2_X1 U7121 ( .A1(n10123), .A2(n10036), .ZN(n6114) );
  NAND2_X1 U7122 ( .A1(n10123), .A2(n10036), .ZN(n7045) );
  MUX2_X1 U7123 ( .A(n7044), .B(n6111), .S(n7064), .Z(n6019) );
  MUX2_X1 U7124 ( .A(n6114), .B(n7045), .S(n7064), .Z(n6020) );
  NAND2_X1 U7125 ( .A1(n6021), .A2(n7047), .ZN(n9983) );
  INV_X1 U7126 ( .A(n9983), .ZN(n6022) );
  XNOR2_X1 U7127 ( .A(n10117), .B(n10022), .ZN(n9997) );
  NAND3_X1 U7128 ( .A1(n6023), .A2(n6022), .A3(n9997), .ZN(n6036) );
  XNOR2_X1 U7129 ( .A(n6025), .B(n6024), .ZN(n8306) );
  NAND2_X1 U7130 ( .A1(n8306), .A2(n6041), .ZN(n6027) );
  OR2_X1 U7131 ( .A1(n5771), .A2(n8309), .ZN(n6026) );
  NAND2_X1 U7132 ( .A1(n6028), .A2(n9513), .ZN(n6029) );
  NAND2_X1 U7133 ( .A1(n6030), .A2(n6029), .ZN(n9963) );
  AOI22_X1 U7134 ( .A1(n5956), .A2(P1_REG1_REG_22__SCAN_IN), .B1(n6031), .B2(
        P1_REG0_REG_22__SCAN_IN), .ZN(n6034) );
  NAND2_X1 U7135 ( .A1(n6032), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n6033) );
  OAI211_X1 U7136 ( .C1(n9963), .C2(n6035), .A(n6034), .B(n6033), .ZN(n9955)
         );
  INV_X1 U7137 ( .A(n9955), .ZN(n9987) );
  OR2_X1 U7138 ( .A1(n10106), .A2(n9987), .ZN(n7049) );
  NAND2_X1 U7139 ( .A1(n10106), .A2(n9987), .ZN(n7050) );
  XNOR2_X1 U7140 ( .A(n10102), .B(n9969), .ZN(n9952) );
  MUX2_X1 U7141 ( .A(n7049), .B(n7050), .S(n4850), .Z(n6038) );
  NAND2_X1 U7142 ( .A1(n8574), .A2(n6041), .ZN(n6043) );
  OR2_X1 U7143 ( .A1(n5771), .A2(n8575), .ZN(n6042) );
  NAND2_X1 U7144 ( .A1(n6044), .A2(n9447), .ZN(n6045) );
  NAND2_X1 U7145 ( .A1(n9917), .A2(n6047), .ZN(n6054) );
  INV_X1 U7146 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n6051) );
  NAND2_X1 U7147 ( .A1(n5734), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n6049) );
  NAND2_X1 U7148 ( .A1(n5760), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n6048) );
  OAI211_X1 U7149 ( .C1(n6051), .C2(n6050), .A(n6049), .B(n6048), .ZN(n6052)
         );
  INV_X1 U7150 ( .A(n6052), .ZN(n6053) );
  NAND2_X1 U7151 ( .A1(n10092), .A2(n9543), .ZN(n7056) );
  MUX2_X1 U7152 ( .A(n7054), .B(n6131), .S(n4850), .Z(n6055) );
  MUX2_X1 U7153 ( .A(n6133), .B(n7056), .S(n7064), .Z(n6057) );
  NAND3_X1 U7154 ( .A1(n8792), .A2(n6059), .A3(n6058), .ZN(n6060) );
  NAND3_X1 U7155 ( .A1(n9896), .A2(n6061), .A3(n6060), .ZN(n6062) );
  OAI211_X1 U7156 ( .C1(n8811), .C2(n7064), .A(n6181), .B(n6062), .ZN(n6063)
         );
  NOR2_X1 U7157 ( .A1(n10072), .A2(n9899), .ZN(n6073) );
  INV_X1 U7158 ( .A(n8810), .ZN(n6064) );
  OR2_X1 U7159 ( .A1(n6073), .A2(n6064), .ZN(n6183) );
  NAND2_X1 U7160 ( .A1(n6183), .A2(n7064), .ZN(n6065) );
  OR2_X1 U7161 ( .A1(n6069), .A2(n6068), .ZN(n6070) );
  INV_X1 U7162 ( .A(n7385), .ZN(n7138) );
  INV_X1 U7163 ( .A(n9921), .ZN(n7055) );
  INV_X1 U7164 ( .A(n8586), .ZN(n6086) );
  INV_X1 U7165 ( .A(n8556), .ZN(n8550) );
  INV_X1 U7166 ( .A(n8518), .ZN(n8522) );
  NAND2_X1 U7167 ( .A1(n7037), .A2(n6097), .ZN(n8419) );
  NAND2_X1 U7168 ( .A1(n6106), .A2(n7035), .ZN(n8343) );
  INV_X1 U7169 ( .A(n7761), .ZN(n6074) );
  NAND2_X1 U7170 ( .A1(n7380), .A2(n7759), .ZN(n6152) );
  NAND2_X1 U7171 ( .A1(n6074), .A2(n6152), .ZN(n7415) );
  NOR4_X1 U7172 ( .A1(n7415), .A2(n7743), .A3(n10406), .A4(n7087), .ZN(n6078)
         );
  NAND4_X1 U7173 ( .A1(n6078), .A2(n7993), .A3(n10487), .A4(n6077), .ZN(n6079)
         );
  NAND2_X1 U7174 ( .A1(n6098), .A2(n7028), .ZN(n8078) );
  NOR4_X1 U7175 ( .A1(n6079), .A2(n7101), .A3(n8078), .A4(n8013), .ZN(n6080)
         );
  NAND4_X1 U7176 ( .A1(n8295), .A2(n8192), .A3(n7031), .A4(n6080), .ZN(n6081)
         );
  NOR4_X1 U7177 ( .A1(n8522), .A2(n8419), .A3(n8343), .A4(n6081), .ZN(n6082)
         );
  NAND4_X1 U7178 ( .A1(n10021), .A2(n8550), .A3(n10050), .A4(n6082), .ZN(n6083) );
  NOR4_X1 U7179 ( .A1(n9983), .A2(n5197), .A3(n10032), .A4(n6083), .ZN(n6084)
         );
  NAND4_X1 U7180 ( .A1(n9928), .A2(n9967), .A3(n6084), .A4(n9952), .ZN(n6085)
         );
  NOR4_X1 U7181 ( .A1(n5366), .A2(n7055), .A3(n6086), .A4(n6085), .ZN(n6088)
         );
  NAND2_X1 U7182 ( .A1(n10067), .A2(n6087), .ZN(n6180) );
  NAND2_X1 U7183 ( .A1(n6090), .A2(n6089), .ZN(n6150) );
  INV_X1 U7184 ( .A(n6144), .ZN(n6092) );
  INV_X1 U7185 ( .A(n6137), .ZN(n8807) );
  INV_X1 U7186 ( .A(n7050), .ZN(n6094) );
  OR3_X1 U7187 ( .A1(n7053), .A2(n6094), .A3(n6093), .ZN(n6128) );
  AND2_X1 U7188 ( .A1(n6095), .A2(n7040), .ZN(n6096) );
  AND2_X1 U7189 ( .A1(n7044), .A2(n6096), .ZN(n6120) );
  AND2_X1 U7190 ( .A1(n7039), .A2(n6097), .ZN(n6121) );
  AND2_X1 U7191 ( .A1(n6098), .A2(n8076), .ZN(n7027) );
  AND2_X1 U7192 ( .A1(n6100), .A2(n7027), .ZN(n6104) );
  INV_X1 U7193 ( .A(n7028), .ZN(n6099) );
  NAND2_X1 U7194 ( .A1(n6100), .A2(n6099), .ZN(n6101) );
  NAND3_X1 U7195 ( .A1(n7032), .A2(n6101), .A3(n7030), .ZN(n6122) );
  OAI211_X1 U7196 ( .C1(n6104), .C2(n6122), .A(n6103), .B(n6102), .ZN(n6105)
         );
  NAND3_X1 U7197 ( .A1(n7035), .A2(n7033), .A3(n6105), .ZN(n6107) );
  NAND3_X1 U7198 ( .A1(n7037), .A2(n6107), .A3(n6106), .ZN(n6108) );
  NAND2_X1 U7199 ( .A1(n6121), .A2(n6108), .ZN(n6110) );
  NAND3_X1 U7200 ( .A1(n7041), .A2(n6110), .A3(n6109), .ZN(n6113) );
  NAND2_X1 U7201 ( .A1(n6111), .A2(n7043), .ZN(n6112) );
  AOI22_X1 U7202 ( .A1(n6120), .A2(n6113), .B1(n6112), .B2(n7044), .ZN(n6115)
         );
  OAI211_X1 U7203 ( .C1(n5196), .C2(n6115), .A(n7046), .B(n6114), .ZN(n6116)
         );
  INV_X1 U7204 ( .A(n6116), .ZN(n6117) );
  OAI22_X1 U7205 ( .A1(n6128), .A2(n6117), .B1(n7053), .B2(n7049), .ZN(n6118)
         );
  NOR2_X1 U7206 ( .A1(n6119), .A2(n6118), .ZN(n6171) );
  NAND2_X1 U7207 ( .A1(n6162), .A2(n10483), .ZN(n7021) );
  AOI21_X1 U7208 ( .B1(n10486), .B2(n10485), .A(n7021), .ZN(n6130) );
  INV_X1 U7209 ( .A(n6120), .ZN(n6126) );
  INV_X1 U7210 ( .A(n6121), .ZN(n6125) );
  INV_X1 U7211 ( .A(n6122), .ZN(n6123) );
  NAND4_X1 U7212 ( .A1(n7035), .A2(n6123), .A3(n7033), .A4(n10542), .ZN(n6124)
         );
  OR3_X1 U7213 ( .A1(n6126), .A2(n6125), .A3(n6124), .ZN(n6127) );
  NOR2_X1 U7214 ( .A1(n6128), .A2(n6127), .ZN(n6168) );
  AND2_X1 U7215 ( .A1(n7045), .A2(n7025), .ZN(n6167) );
  OAI211_X1 U7216 ( .C1(n6130), .C2(n6129), .A(n6168), .B(n6167), .ZN(n6132)
         );
  NAND2_X1 U7217 ( .A1(n7056), .A2(n6131), .ZN(n6169) );
  AOI21_X1 U7218 ( .B1(n6171), .B2(n6132), .A(n6169), .ZN(n6135) );
  NAND2_X1 U7219 ( .A1(n6134), .A2(n6133), .ZN(n6173) );
  NOR3_X1 U7220 ( .A1(n8807), .A2(n6135), .A3(n6173), .ZN(n6138) );
  NAND2_X1 U7221 ( .A1(n8811), .A2(n6136), .ZN(n6178) );
  INV_X1 U7222 ( .A(n7057), .ZN(n8806) );
  AND2_X1 U7223 ( .A1(n6137), .A2(n8806), .ZN(n6175) );
  NOR3_X1 U7224 ( .A1(n6138), .A2(n6178), .A3(n6175), .ZN(n6140) );
  OAI211_X1 U7225 ( .C1(n6140), .C2(n6183), .A(n6139), .B(n6181), .ZN(n6141)
         );
  AOI211_X1 U7226 ( .C1(n6142), .C2(n6141), .A(n8185), .B(n6184), .ZN(n6143)
         );
  NOR2_X1 U7227 ( .A1(n6144), .A2(n6143), .ZN(n6145) );
  MUX2_X1 U7228 ( .A(n6146), .B(n6145), .S(n8116), .Z(n6194) );
  NAND2_X1 U7229 ( .A1(n5386), .A2(n7063), .ZN(n6193) );
  INV_X1 U7230 ( .A(n6150), .ZN(n6186) );
  NAND2_X1 U7231 ( .A1(n7491), .A2(n10357), .ZN(n6151) );
  NAND3_X1 U7232 ( .A1(n6152), .A2(n7130), .A3(n6151), .ZN(n6153) );
  NAND2_X1 U7233 ( .A1(n6154), .A2(n6153), .ZN(n6156) );
  OAI21_X1 U7234 ( .B1(n7665), .B2(n6156), .A(n6155), .ZN(n6158) );
  AOI21_X1 U7235 ( .B1(n6158), .B2(n10407), .A(n6157), .ZN(n6165) );
  NAND3_X1 U7236 ( .A1(n6162), .A2(n10483), .A3(n6159), .ZN(n6164) );
  NAND2_X1 U7237 ( .A1(n10485), .A2(n6160), .ZN(n6161) );
  NAND2_X1 U7238 ( .A1(n6162), .A2(n6161), .ZN(n7022) );
  OAI211_X1 U7239 ( .C1(n6165), .C2(n6164), .A(n7022), .B(n6163), .ZN(n6166)
         );
  NAND3_X1 U7240 ( .A1(n6168), .A2(n6167), .A3(n6166), .ZN(n6170) );
  AOI21_X1 U7241 ( .B1(n6171), .B2(n6170), .A(n6169), .ZN(n6172) );
  NOR2_X1 U7242 ( .A1(n6173), .A2(n6172), .ZN(n6174) );
  NAND2_X1 U7243 ( .A1(n8792), .A2(n6174), .ZN(n6177) );
  INV_X1 U7244 ( .A(n6175), .ZN(n6176) );
  NAND2_X1 U7245 ( .A1(n6177), .A2(n6176), .ZN(n6179) );
  NOR2_X1 U7246 ( .A1(n6179), .A2(n6178), .ZN(n6182) );
  OAI211_X1 U7247 ( .C1(n6183), .C2(n6182), .A(n6181), .B(n6180), .ZN(n6185)
         );
  AOI21_X1 U7248 ( .B1(n6186), .B2(n6185), .A(n6184), .ZN(n6187) );
  NAND2_X1 U7249 ( .A1(n8166), .A2(n8116), .ZN(n7668) );
  INV_X1 U7250 ( .A(n7668), .ZN(n7376) );
  NAND2_X1 U7251 ( .A1(n4912), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6189) );
  XNOR2_X1 U7252 ( .A(n6189), .B(n6188), .ZN(n7141) );
  OR2_X1 U7253 ( .A1(n7141), .A2(P1_U3084), .ZN(n8397) );
  INV_X1 U7254 ( .A(n8397), .ZN(n6190) );
  OAI211_X1 U7255 ( .C1(n5394), .C2(n7063), .A(n5393), .B(n6190), .ZN(n6191)
         );
  INV_X1 U7256 ( .A(n6191), .ZN(n6192) );
  NAND2_X1 U7257 ( .A1(n6195), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6199) );
  XNOR2_X1 U7258 ( .A(n6199), .B(P1_IR_REG_25__SCAN_IN), .ZN(n7080) );
  NAND2_X1 U7259 ( .A1(n6196), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6197) );
  XNOR2_X1 U7260 ( .A(n6197), .B(n5540), .ZN(n8452) );
  NAND2_X1 U7261 ( .A1(n6199), .A2(n6198), .ZN(n6200) );
  INV_X1 U7262 ( .A(n7066), .ZN(n6203) );
  AND2_X1 U7263 ( .A1(n7141), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6204) );
  OR2_X1 U7264 ( .A1(n7138), .A2(n7668), .ZN(n7670) );
  NOR4_X1 U7265 ( .A1(n7388), .A2(n6205), .A3(n7670), .A4(n10260), .ZN(n6207)
         );
  INV_X1 U7266 ( .A(P1_B_REG_SCAN_IN), .ZN(n8815) );
  NAND2_X1 U7267 ( .A1(n5383), .A2(P1_B_REG_SCAN_IN), .ZN(n6206) );
  OR2_X1 U7268 ( .A1(n6207), .A2(n6206), .ZN(n6208) );
  NAND3_X1 U7269 ( .A1(n6489), .A2(n6625), .A3(n6628), .ZN(n6212) );
  INV_X1 U7270 ( .A(n6236), .ZN(n6218) );
  INV_X1 U7271 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n6217) );
  NAND2_X1 U7272 ( .A1(n6218), .A2(n6217), .ZN(n6233) );
  NOR2_X2 U7273 ( .A1(n6233), .A2(P2_IR_REG_29__SCAN_IN), .ZN(n6221) );
  INV_X1 U7274 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n6219) );
  XNOR2_X2 U7275 ( .A(n6220), .B(n6219), .ZN(n6227) );
  INV_X1 U7276 ( .A(n6221), .ZN(n9371) );
  NAND2_X1 U7277 ( .A1(n6233), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6222) );
  MUX2_X1 U7278 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6222), .S(
        P2_IR_REG_29__SCAN_IN), .Z(n6223) );
  INV_X1 U7279 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n6224) );
  AND2_X4 U7280 ( .A1(n6227), .A2(n9379), .ZN(n6605) );
  NOR2_X1 U7281 ( .A1(n6226), .A2(n6225), .ZN(n6231) );
  INV_X1 U7282 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n7154) );
  OR2_X1 U7283 ( .A1(n6498), .A2(n7154), .ZN(n6230) );
  AND2_X4 U7284 ( .A1(n9375), .A2(n9379), .ZN(n6286) );
  NAND2_X1 U7285 ( .A1(n6286), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n6229) );
  NAND3_X1 U7286 ( .A1(n6231), .A2(n6230), .A3(n6229), .ZN(n6242) );
  NAND2_X1 U7287 ( .A1(n6236), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6232) );
  NAND2_X1 U7288 ( .A1(n6234), .A2(n6233), .ZN(n6841) );
  MUX2_X1 U7289 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6235), .S(
        P2_IR_REG_27__SCAN_IN), .Z(n6237) );
  NAND2_X1 U7290 ( .A1(n6259), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n6241) );
  OR2_X1 U7291 ( .A1(n6239), .A2(n9370), .ZN(n6261) );
  XNOR2_X1 U7292 ( .A(n6261), .B(P2_IR_REG_2__SCAN_IN), .ZN(n8950) );
  NAND2_X1 U7293 ( .A1(n7177), .A2(n8950), .ZN(n6240) );
  OAI211_X1 U7294 ( .C1(n6328), .C2(n7234), .A(n6241), .B(n6240), .ZN(n7707)
         );
  INV_X1 U7295 ( .A(n7707), .ZN(n10377) );
  NAND2_X1 U7296 ( .A1(n6242), .A2(n10377), .ZN(n6649) );
  NAND2_X1 U7297 ( .A1(n6860), .A2(n7707), .ZN(n6258) );
  NAND2_X1 U7298 ( .A1(n6286), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n6247) );
  NAND2_X1 U7299 ( .A1(n6605), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6246) );
  INV_X1 U7300 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6243) );
  OR2_X1 U7301 ( .A1(n6273), .A2(n7438), .ZN(n6244) );
  NAND2_X1 U7302 ( .A1(n5021), .A2(SI_0_), .ZN(n6249) );
  INV_X1 U7303 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n6248) );
  NAND2_X1 U7304 ( .A1(n6249), .A2(n6248), .ZN(n6251) );
  AND2_X1 U7305 ( .A1(n6251), .A2(n6250), .ZN(n9388) );
  MUX2_X1 U7306 ( .A(P2_IR_REG_0__SCAN_IN), .B(n9388), .S(n7172), .Z(n7565) );
  NAND2_X1 U7307 ( .A1(n7485), .A2(n7565), .ZN(n7562) );
  NAND2_X1 U7308 ( .A1(n6286), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n6256) );
  NAND2_X1 U7309 ( .A1(n6605), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6255) );
  INV_X1 U7310 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n7881) );
  OR2_X1 U7311 ( .A1(n6498), .A2(n7881), .ZN(n6254) );
  INV_X1 U7312 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n6252) );
  OR2_X1 U7313 ( .A1(n6273), .A2(n6252), .ZN(n6253) );
  NAND2_X1 U7314 ( .A1(n7562), .A2(n6797), .ZN(n6257) );
  NAND4_X1 U7315 ( .A1(n6256), .A2(n6255), .A3(n6254), .A4(n6253), .ZN(n8946)
         );
  INV_X1 U7316 ( .A(n7885), .ZN(n7686) );
  NAND2_X1 U7317 ( .A1(n8946), .A2(n7686), .ZN(n6796) );
  AND2_X1 U7318 ( .A1(n6257), .A2(n6796), .ZN(n7695) );
  NAND2_X1 U7319 ( .A1(n7694), .A2(n7695), .ZN(n7693) );
  NAND2_X1 U7320 ( .A1(n7693), .A2(n6258), .ZN(n6651) );
  NAND2_X1 U7321 ( .A1(n4852), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n6265) );
  INV_X1 U7322 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n6260) );
  NAND2_X1 U7323 ( .A1(n6261), .A2(n6260), .ZN(n6262) );
  NAND2_X1 U7324 ( .A1(n6262), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6263) );
  XNOR2_X1 U7325 ( .A(n6263), .B(P2_IR_REG_3__SCAN_IN), .ZN(n7475) );
  NAND2_X1 U7326 ( .A1(n7177), .A2(n7475), .ZN(n6264) );
  INV_X1 U7327 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6266) );
  OR2_X1 U7328 ( .A1(n6498), .A2(n6266), .ZN(n6271) );
  INV_X1 U7329 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n9745) );
  NAND2_X1 U7330 ( .A1(n6286), .A2(n9745), .ZN(n6270) );
  INV_X1 U7331 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n6267) );
  OR2_X1 U7332 ( .A1(n6273), .A2(n6267), .ZN(n6269) );
  NAND2_X1 U7333 ( .A1(n6605), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6268) );
  NAND2_X1 U7334 ( .A1(n6651), .A2(n7730), .ZN(n7729) );
  NAND2_X1 U7335 ( .A1(n6482), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6278) );
  NAND2_X1 U7336 ( .A1(n6605), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6277) );
  OAI21_X1 U7337 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(P2_REG3_REG_4__SCAN_IN), 
        .A(n6288), .ZN(n10447) );
  INV_X1 U7338 ( .A(n10447), .ZN(n6272) );
  NAND2_X1 U7339 ( .A1(n6286), .A2(n6272), .ZN(n6276) );
  INV_X1 U7340 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n6274) );
  NAND4_X1 U7341 ( .A1(n6278), .A2(n6277), .A3(n6276), .A4(n6275), .ZN(n8943)
         );
  NAND2_X1 U7342 ( .A1(n5250), .A2(n6279), .ZN(n6284) );
  NAND2_X1 U7343 ( .A1(n4851), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n6283) );
  NAND2_X1 U7344 ( .A1(n6280), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6281) );
  XNOR2_X1 U7345 ( .A(n6281), .B(P2_IR_REG_4__SCAN_IN), .ZN(n7218) );
  NAND2_X1 U7346 ( .A1(n7177), .A2(n7218), .ZN(n6282) );
  NAND2_X1 U7347 ( .A1(n8943), .A2(n10434), .ZN(n8050) );
  NAND2_X1 U7348 ( .A1(n6605), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6295) );
  INV_X1 U7349 ( .A(n6288), .ZN(n6287) );
  NAND2_X1 U7350 ( .A1(n6287), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n6304) );
  INV_X1 U7351 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n9754) );
  NAND2_X1 U7352 ( .A1(n6288), .A2(n9754), .ZN(n6289) );
  AND2_X1 U7353 ( .A1(n6304), .A2(n6289), .ZN(n8054) );
  NAND2_X1 U7354 ( .A1(n6286), .A2(n8054), .ZN(n6294) );
  INV_X1 U7355 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n6290) );
  OR2_X1 U7356 ( .A1(n6498), .A2(n6290), .ZN(n6293) );
  INV_X1 U7357 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n6291) );
  OR2_X1 U7358 ( .A1(n6273), .A2(n6291), .ZN(n6292) );
  NAND2_X1 U7359 ( .A1(n4851), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n6299) );
  NAND2_X1 U7360 ( .A1(n6296), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6297) );
  XNOR2_X1 U7361 ( .A(n6297), .B(P2_IR_REG_5__SCAN_IN), .ZN(n7191) );
  NAND2_X1 U7362 ( .A1(n7177), .A2(n7191), .ZN(n6298) );
  INV_X1 U7363 ( .A(n10473), .ZN(n8059) );
  NAND2_X1 U7364 ( .A1(n8942), .A2(n8059), .ZN(n6665) );
  AND2_X1 U7365 ( .A1(n8050), .A2(n6665), .ZN(n6301) );
  NAND2_X1 U7366 ( .A1(n10439), .A2(n10473), .ZN(n6666) );
  INV_X1 U7367 ( .A(n6666), .ZN(n6300) );
  NAND2_X1 U7368 ( .A1(n6612), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n6309) );
  NAND2_X1 U7369 ( .A1(n6482), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6308) );
  INV_X1 U7370 ( .A(n6304), .ZN(n6302) );
  INV_X1 U7371 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n6303) );
  NAND2_X1 U7372 ( .A1(n6304), .A2(n6303), .ZN(n6305) );
  AND2_X1 U7373 ( .A1(n6316), .A2(n6305), .ZN(n7868) );
  NAND2_X1 U7374 ( .A1(n6286), .A2(n7868), .ZN(n6307) );
  NAND2_X1 U7375 ( .A1(n6605), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6306) );
  NAND4_X1 U7376 ( .A1(n6309), .A2(n6308), .A3(n6307), .A4(n6306), .ZN(n8941)
         );
  NAND2_X1 U7377 ( .A1(n5250), .A2(n7239), .ZN(n6313) );
  NAND2_X1 U7378 ( .A1(n4851), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n6312) );
  NOR2_X1 U7379 ( .A1(n6296), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n6324) );
  OR2_X1 U7380 ( .A1(n6324), .A2(n9370), .ZN(n6310) );
  XNOR2_X1 U7381 ( .A(n6310), .B(P2_IR_REG_6__SCAN_IN), .ZN(n7205) );
  NAND2_X1 U7382 ( .A1(n7177), .A2(n7205), .ZN(n6311) );
  AND2_X1 U7383 ( .A1(n8941), .A2(n10509), .ZN(n6314) );
  INV_X1 U7384 ( .A(n7978), .ZN(n6330) );
  NAND2_X1 U7385 ( .A1(n6605), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6322) );
  INV_X1 U7386 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n7147) );
  NAND2_X1 U7387 ( .A1(n6316), .A2(n7147), .ZN(n6317) );
  AND2_X1 U7388 ( .A1(n6331), .A2(n6317), .ZN(n7146) );
  NAND2_X1 U7389 ( .A1(n6286), .A2(n7146), .ZN(n6321) );
  INV_X1 U7390 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n7980) );
  OR2_X1 U7391 ( .A1(n6498), .A2(n7980), .ZN(n6320) );
  INV_X1 U7392 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n6318) );
  OR2_X1 U7393 ( .A1(n6273), .A2(n6318), .ZN(n6319) );
  NAND2_X1 U7394 ( .A1(n4851), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n6327) );
  NAND2_X1 U7395 ( .A1(n6324), .A2(n6323), .ZN(n6339) );
  NAND2_X1 U7396 ( .A1(n6339), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6325) );
  XNOR2_X1 U7397 ( .A(n6325), .B(P2_IR_REG_7__SCAN_IN), .ZN(n7524) );
  NAND2_X1 U7398 ( .A1(n7177), .A2(n7524), .ZN(n6326) );
  NAND2_X1 U7399 ( .A1(n8065), .A2(n10525), .ZN(n6673) );
  INV_X1 U7400 ( .A(n8065), .ZN(n8940) );
  NAND2_X1 U7401 ( .A1(n8940), .A2(n7985), .ZN(n7949) );
  NAND2_X1 U7402 ( .A1(n6673), .A2(n7949), .ZN(n7963) );
  NAND2_X1 U7403 ( .A1(n6330), .A2(n6329), .ZN(n7950) );
  NAND2_X1 U7404 ( .A1(n6331), .A2(n8068), .ZN(n6332) );
  AND2_X1 U7405 ( .A1(n6346), .A2(n6332), .ZN(n8071) );
  NAND2_X1 U7406 ( .A1(n6286), .A2(n8071), .ZN(n6338) );
  NAND2_X1 U7407 ( .A1(n6605), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n6337) );
  INV_X1 U7408 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n6333) );
  OR2_X1 U7409 ( .A1(n6273), .A2(n6333), .ZN(n6336) );
  INV_X1 U7410 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n6334) );
  OR2_X1 U7411 ( .A1(n6498), .A2(n6334), .ZN(n6335) );
  NAND2_X1 U7412 ( .A1(n5250), .A2(n7251), .ZN(n6342) );
  NAND2_X1 U7413 ( .A1(n6354), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6340) );
  XNOR2_X1 U7414 ( .A(n6340), .B(P2_IR_REG_8__SCAN_IN), .ZN(n7545) );
  NAND2_X1 U7415 ( .A1(n7177), .A2(n7545), .ZN(n6341) );
  OAI211_X1 U7416 ( .C1(n6504), .C2(n7254), .A(n6342), .B(n6341), .ZN(n8131)
         );
  NAND2_X1 U7417 ( .A1(n8175), .A2(n8131), .ZN(n6676) );
  INV_X1 U7418 ( .A(n8131), .ZN(n10575) );
  NAND2_X1 U7419 ( .A1(n8135), .A2(n10575), .ZN(n6675) );
  NAND2_X1 U7420 ( .A1(n6676), .A2(n6675), .ZN(n6802) );
  INV_X1 U7421 ( .A(n7949), .ZN(n6343) );
  NOR2_X1 U7422 ( .A1(n6802), .A2(n6343), .ZN(n6344) );
  NAND2_X1 U7423 ( .A1(n7950), .A2(n6344), .ZN(n7948) );
  INV_X1 U7424 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n9669) );
  NAND2_X1 U7425 ( .A1(n6346), .A2(n9669), .ZN(n6347) );
  AND2_X1 U7426 ( .A1(n6357), .A2(n6347), .ZN(n8171) );
  NAND2_X1 U7427 ( .A1(n6286), .A2(n8171), .ZN(n6353) );
  NAND2_X1 U7428 ( .A1(n6605), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n6352) );
  INV_X1 U7429 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n6348) );
  OR2_X1 U7430 ( .A1(n6498), .A2(n6348), .ZN(n6351) );
  INV_X1 U7431 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n6349) );
  OR2_X1 U7432 ( .A1(n6273), .A2(n6349), .ZN(n6350) );
  NAND2_X1 U7433 ( .A1(n6388), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6365) );
  XNOR2_X1 U7434 ( .A(n6365), .B(P2_IR_REG_9__SCAN_IN), .ZN(n7613) );
  AOI22_X1 U7435 ( .A1(n4852), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n7177), .B2(
        n7613), .ZN(n6355) );
  NAND2_X1 U7436 ( .A1(n10612), .A2(n8179), .ZN(n6686) );
  NAND2_X1 U7437 ( .A1(n6686), .A2(n6680), .ZN(n8136) );
  NAND2_X1 U7438 ( .A1(n6357), .A2(n6356), .ZN(n6358) );
  AND2_X1 U7439 ( .A1(n6376), .A2(n6358), .ZN(n10630) );
  NAND2_X1 U7440 ( .A1(n6286), .A2(n10630), .ZN(n6364) );
  NAND2_X1 U7441 ( .A1(n6605), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n6363) );
  INV_X1 U7442 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n6359) );
  OR2_X1 U7443 ( .A1(n6273), .A2(n6359), .ZN(n6362) );
  INV_X1 U7444 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n6360) );
  OR2_X1 U7445 ( .A1(n6498), .A2(n6360), .ZN(n6361) );
  NAND2_X1 U7446 ( .A1(n7290), .A2(n5250), .ZN(n6370) );
  AOI21_X1 U7447 ( .B1(n6365), .B2(n6386), .A(n9370), .ZN(n6366) );
  NAND2_X1 U7448 ( .A1(n6366), .A2(P2_IR_REG_10__SCAN_IN), .ZN(n6368) );
  INV_X1 U7449 ( .A(n6366), .ZN(n6367) );
  NAND2_X1 U7450 ( .A1(n6367), .A2(n6385), .ZN(n6371) );
  AOI22_X1 U7451 ( .A1(n4852), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n7177), .B2(
        n7940), .ZN(n6369) );
  NAND2_X1 U7452 ( .A1(n6370), .A2(n6369), .ZN(n10606) );
  OR2_X1 U7453 ( .A1(n8246), .A2(n10606), .ZN(n6688) );
  NAND2_X1 U7454 ( .A1(n10606), .A2(n8246), .ZN(n6685) );
  NAND2_X1 U7455 ( .A1(n7260), .A2(n5250), .ZN(n6374) );
  NAND2_X1 U7456 ( .A1(n6371), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6372) );
  XNOR2_X1 U7457 ( .A(n6372), .B(P2_IR_REG_11__SCAN_IN), .ZN(n8963) );
  AOI22_X1 U7458 ( .A1(n4852), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n7177), .B2(
        n8963), .ZN(n6373) );
  NAND2_X1 U7459 ( .A1(n6605), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n6383) );
  INV_X1 U7460 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n9767) );
  NAND2_X1 U7461 ( .A1(n6376), .A2(n9767), .ZN(n6377) );
  AND2_X1 U7462 ( .A1(n6393), .A2(n6377), .ZN(n8253) );
  NAND2_X1 U7463 ( .A1(n6286), .A2(n8253), .ZN(n6382) );
  INV_X1 U7464 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n6378) );
  OR2_X1 U7465 ( .A1(n6498), .A2(n6378), .ZN(n6381) );
  INV_X1 U7466 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n6379) );
  OR2_X1 U7467 ( .A1(n6273), .A2(n6379), .ZN(n6380) );
  AND2_X1 U7468 ( .A1(n10640), .A2(n10614), .ZN(n6694) );
  OR2_X1 U7469 ( .A1(n10640), .A2(n10614), .ZN(n6794) );
  OAI21_X1 U7470 ( .B1(n8227), .B2(n6694), .A(n6794), .ZN(n8279) );
  NAND2_X1 U7471 ( .A1(n7422), .A2(n5250), .ZN(n6391) );
  INV_X1 U7472 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n6384) );
  NAND3_X1 U7473 ( .A1(n6386), .A2(n6385), .A3(n6384), .ZN(n6387) );
  NOR2_X1 U7474 ( .A1(n6388), .A2(n6387), .ZN(n6402) );
  OR2_X1 U7475 ( .A1(n6402), .A2(n9370), .ZN(n6389) );
  XNOR2_X1 U7476 ( .A(n6389), .B(P2_IR_REG_12__SCAN_IN), .ZN(n8026) );
  AOI22_X1 U7477 ( .A1(n4852), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n7177), .B2(
        n8026), .ZN(n6390) );
  NAND2_X1 U7478 ( .A1(n6605), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n6400) );
  INV_X1 U7479 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n6392) );
  NAND2_X1 U7480 ( .A1(n6393), .A2(n6392), .ZN(n6394) );
  AND2_X1 U7481 ( .A1(n6406), .A2(n6394), .ZN(n8404) );
  NAND2_X1 U7482 ( .A1(n6286), .A2(n8404), .ZN(n6399) );
  INV_X1 U7483 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n6395) );
  OR2_X1 U7484 ( .A1(n6498), .A2(n6395), .ZN(n6398) );
  INV_X1 U7485 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n6396) );
  OR2_X1 U7486 ( .A1(n6273), .A2(n6396), .ZN(n6397) );
  OR2_X1 U7487 ( .A1(n8411), .A2(n8374), .ZN(n6698) );
  NAND2_X1 U7488 ( .A1(n8411), .A2(n8374), .ZN(n6697) );
  NAND2_X1 U7489 ( .A1(n6698), .A2(n6697), .ZN(n8284) );
  NAND2_X1 U7490 ( .A1(n7547), .A2(n5250), .ZN(n6405) );
  NAND2_X1 U7491 ( .A1(n6402), .A2(n6401), .ZN(n6403) );
  NAND2_X1 U7492 ( .A1(n6403), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6416) );
  XNOR2_X1 U7493 ( .A(n6416), .B(P2_IR_REG_13__SCAN_IN), .ZN(n8122) );
  AOI22_X1 U7494 ( .A1(n4851), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n7177), .B2(
        n8122), .ZN(n6404) );
  NAND2_X1 U7495 ( .A1(n6406), .A2(n9667), .ZN(n6407) );
  AND2_X1 U7496 ( .A1(n6422), .A2(n6407), .ZN(n8370) );
  NAND2_X1 U7497 ( .A1(n6286), .A2(n8370), .ZN(n6413) );
  NAND2_X1 U7498 ( .A1(n6605), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n6412) );
  INV_X1 U7499 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n6408) );
  OR2_X1 U7500 ( .A1(n6498), .A2(n6408), .ZN(n6411) );
  INV_X1 U7501 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n6409) );
  OR2_X1 U7502 ( .A1(n6273), .A2(n6409), .ZN(n6410) );
  OR2_X1 U7503 ( .A1(n8371), .A2(n8504), .ZN(n6705) );
  NAND2_X1 U7504 ( .A1(n8371), .A2(n8504), .ZN(n6704) );
  NAND2_X1 U7505 ( .A1(n8367), .A2(n6805), .ZN(n6414) );
  NAND2_X1 U7506 ( .A1(n7680), .A2(n5250), .ZN(n6419) );
  NAND2_X1 U7507 ( .A1(n6416), .A2(n6415), .ZN(n6417) );
  NAND2_X1 U7508 ( .A1(n6417), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6432) );
  XNOR2_X1 U7509 ( .A(n6432), .B(P2_IR_REG_14__SCAN_IN), .ZN(n8436) );
  AOI22_X1 U7510 ( .A1(n4851), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n7177), .B2(
        n8436), .ZN(n6418) );
  NAND2_X1 U7511 ( .A1(n6605), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n6429) );
  INV_X1 U7512 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n6421) );
  NAND2_X1 U7513 ( .A1(n6422), .A2(n6421), .ZN(n6423) );
  AND2_X1 U7514 ( .A1(n6438), .A2(n6423), .ZN(n8509) );
  NAND2_X1 U7515 ( .A1(n6286), .A2(n8509), .ZN(n6428) );
  INV_X1 U7516 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n6424) );
  OR2_X1 U7517 ( .A1(n6498), .A2(n6424), .ZN(n6427) );
  INV_X1 U7518 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n6425) );
  OR2_X1 U7519 ( .A1(n6273), .A2(n6425), .ZN(n6426) );
  NAND2_X1 U7520 ( .A1(n10661), .A2(n8783), .ZN(n6711) );
  NAND2_X1 U7521 ( .A1(n6712), .A2(n6711), .ZN(n8493) );
  INV_X1 U7522 ( .A(n8493), .ZN(n6430) );
  NAND2_X1 U7523 ( .A1(n7818), .A2(n5250), .ZN(n6436) );
  NAND2_X1 U7524 ( .A1(n6432), .A2(n6431), .ZN(n6433) );
  NAND2_X1 U7525 ( .A1(n6433), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6434) );
  XNOR2_X1 U7526 ( .A(n6434), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8978) );
  AOI22_X1 U7527 ( .A1(n4851), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n7177), .B2(
        n8978), .ZN(n6435) );
  NAND2_X1 U7528 ( .A1(n6605), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n6445) );
  INV_X1 U7529 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n9775) );
  NAND2_X1 U7530 ( .A1(n6438), .A2(n9775), .ZN(n6439) );
  AND2_X1 U7531 ( .A1(n6450), .A2(n6439), .ZN(n8776) );
  NAND2_X1 U7532 ( .A1(n6286), .A2(n8776), .ZN(n6444) );
  INV_X1 U7533 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n6440) );
  OR2_X1 U7534 ( .A1(n6498), .A2(n6440), .ZN(n6443) );
  INV_X1 U7535 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n6441) );
  OR2_X1 U7536 ( .A1(n6273), .A2(n6441), .ZN(n6442) );
  NAND2_X1 U7537 ( .A1(n8781), .A2(n8505), .ZN(n6715) );
  NAND2_X1 U7538 ( .A1(n7846), .A2(n5250), .ZN(n6448) );
  OR2_X1 U7539 ( .A1(n6459), .A2(n9370), .ZN(n6446) );
  XNOR2_X1 U7540 ( .A(n6446), .B(P2_IR_REG_16__SCAN_IN), .ZN(n8989) );
  AOI22_X1 U7541 ( .A1(n4851), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n7177), .B2(
        n8989), .ZN(n6447) );
  INV_X1 U7542 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n6449) );
  NAND2_X1 U7543 ( .A1(n6450), .A2(n6449), .ZN(n6451) );
  AND2_X1 U7544 ( .A1(n6464), .A2(n6451), .ZN(n8545) );
  NAND2_X1 U7545 ( .A1(n6286), .A2(n8545), .ZN(n6457) );
  NAND2_X1 U7546 ( .A1(n6605), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n6456) );
  INV_X1 U7547 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n6452) );
  OR2_X1 U7548 ( .A1(n6273), .A2(n6452), .ZN(n6455) );
  INV_X1 U7549 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n6453) );
  OR2_X1 U7550 ( .A1(n6498), .A2(n6453), .ZN(n6454) );
  NAND2_X1 U7551 ( .A1(n9349), .A2(n8775), .ZN(n9256) );
  NAND2_X1 U7552 ( .A1(n7888), .A2(n5250), .ZN(n6462) );
  OR2_X1 U7553 ( .A1(n6479), .A2(n9370), .ZN(n6460) );
  XNOR2_X1 U7554 ( .A(n6460), .B(P2_IR_REG_17__SCAN_IN), .ZN(n9004) );
  AOI22_X1 U7555 ( .A1(n4852), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n7177), .B2(
        n9004), .ZN(n6461) );
  NAND2_X1 U7556 ( .A1(n6612), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n6469) );
  NAND2_X1 U7557 ( .A1(n6482), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n6468) );
  INV_X1 U7558 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n9758) );
  NAND2_X1 U7559 ( .A1(n6464), .A2(n9758), .ZN(n6465) );
  AND2_X1 U7560 ( .A1(n6483), .A2(n6465), .ZN(n9267) );
  NAND2_X1 U7561 ( .A1(n6286), .A2(n9267), .ZN(n6467) );
  NAND2_X1 U7562 ( .A1(n6605), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n6466) );
  NAND4_X1 U7563 ( .A1(n6469), .A2(n6468), .A3(n6467), .A4(n6466), .ZN(n8933)
         );
  INV_X1 U7564 ( .A(n8933), .ZN(n9249) );
  OR2_X1 U7565 ( .A1(n9343), .A2(n9249), .ZN(n6473) );
  INV_X1 U7566 ( .A(n6473), .ZN(n6470) );
  NAND2_X1 U7567 ( .A1(n9343), .A2(n8933), .ZN(n6725) );
  NAND2_X1 U7568 ( .A1(n9046), .A2(n6725), .ZN(n9045) );
  OR2_X1 U7569 ( .A1(n6470), .A2(n9045), .ZN(n6472) );
  AND2_X1 U7570 ( .A1(n9256), .A2(n6472), .ZN(n6471) );
  INV_X1 U7571 ( .A(n6472), .ZN(n6475) );
  AND2_X1 U7572 ( .A1(n9257), .A2(n6473), .ZN(n6474) );
  OR2_X1 U7573 ( .A1(n6475), .A2(n6474), .ZN(n6476) );
  NAND2_X1 U7574 ( .A1(n6477), .A2(n6476), .ZN(n9245) );
  NAND2_X1 U7575 ( .A1(n8003), .A2(n5250), .ZN(n6481) );
  INV_X1 U7576 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n6478) );
  XNOR2_X1 U7577 ( .A(n6490), .B(P2_IR_REG_18__SCAN_IN), .ZN(n9017) );
  AOI22_X1 U7578 ( .A1(n4852), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n7177), .B2(
        n9017), .ZN(n6480) );
  NAND2_X1 U7579 ( .A1(n6612), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n6488) );
  NAND2_X1 U7580 ( .A1(n6482), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n6487) );
  INV_X1 U7581 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n9773) );
  NAND2_X1 U7582 ( .A1(n6483), .A2(n9773), .ZN(n6484) );
  AND2_X1 U7583 ( .A1(n6496), .A2(n6484), .ZN(n9242) );
  NAND2_X1 U7584 ( .A1(n6286), .A2(n9242), .ZN(n6486) );
  NAND2_X1 U7585 ( .A1(n6605), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n6485) );
  NAND4_X1 U7586 ( .A1(n6488), .A2(n6487), .A3(n6486), .A4(n6485), .ZN(n8932)
         );
  XNOR2_X1 U7587 ( .A(n9336), .B(n8932), .ZN(n9237) );
  INV_X1 U7588 ( .A(n8932), .ZN(n9047) );
  OR2_X1 U7589 ( .A1(n9336), .A2(n9047), .ZN(n9225) );
  NAND2_X1 U7590 ( .A1(n8112), .A2(n5250), .ZN(n6493) );
  AOI22_X1 U7591 ( .A1(n4851), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n7177), .B2(
        n4849), .ZN(n6492) );
  INV_X1 U7592 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n6495) );
  NAND2_X1 U7593 ( .A1(n6496), .A2(n6495), .ZN(n6497) );
  AND2_X1 U7594 ( .A1(n6509), .A2(n6497), .ZN(n9231) );
  NAND2_X1 U7595 ( .A1(n9231), .A2(n6286), .ZN(n6503) );
  NAND2_X1 U7596 ( .A1(n6605), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n6502) );
  INV_X1 U7597 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n9023) );
  OR2_X1 U7598 ( .A1(n6498), .A2(n9023), .ZN(n6501) );
  INV_X1 U7599 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n6499) );
  OR2_X1 U7600 ( .A1(n6273), .A2(n6499), .ZN(n6500) );
  NAND2_X1 U7601 ( .A1(n9333), .A2(n9248), .ZN(n6732) );
  NAND2_X1 U7602 ( .A1(n8164), .A2(n5250), .ZN(n6506) );
  NAND2_X1 U7603 ( .A1(n4852), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n6505) );
  NAND2_X1 U7604 ( .A1(n6482), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n6508) );
  NAND2_X1 U7605 ( .A1(n6605), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n6507) );
  AND2_X1 U7606 ( .A1(n6508), .A2(n6507), .ZN(n6513) );
  INV_X1 U7607 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n9661) );
  NAND2_X1 U7608 ( .A1(n6509), .A2(n9661), .ZN(n6510) );
  AND2_X1 U7609 ( .A1(n6517), .A2(n6510), .ZN(n9208) );
  NAND2_X1 U7610 ( .A1(n9208), .A2(n6286), .ZN(n6512) );
  NAND2_X1 U7611 ( .A1(n6612), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n6511) );
  NAND2_X1 U7612 ( .A1(n9326), .A2(n9196), .ZN(n6742) );
  NAND2_X1 U7613 ( .A1(n9216), .A2(n6743), .ZN(n9194) );
  NAND2_X1 U7614 ( .A1(n8183), .A2(n5250), .ZN(n6515) );
  NAND2_X1 U7615 ( .A1(n4851), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n6514) );
  INV_X1 U7616 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n9644) );
  NAND2_X1 U7617 ( .A1(n6517), .A2(n9644), .ZN(n6518) );
  NAND2_X1 U7618 ( .A1(n6524), .A2(n6518), .ZN(n9190) );
  OR2_X1 U7619 ( .A1(n9190), .A2(n6574), .ZN(n6521) );
  AOI22_X1 U7620 ( .A1(n6482), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n6612), .B2(
        P2_REG0_REG_21__SCAN_IN), .ZN(n6520) );
  NAND2_X1 U7621 ( .A1(n6605), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n6519) );
  NAND2_X1 U7622 ( .A1(n9321), .A2(n9214), .ZN(n6644) );
  NAND2_X1 U7623 ( .A1(n9194), .A2(n9188), .ZN(n9199) );
  NAND2_X1 U7624 ( .A1(n9199), .A2(n6645), .ZN(n9175) );
  NAND2_X1 U7625 ( .A1(n8306), .A2(n5250), .ZN(n6523) );
  NAND2_X1 U7626 ( .A1(n4852), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n6522) );
  INV_X1 U7627 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n8895) );
  NAND2_X1 U7628 ( .A1(n6524), .A2(n8895), .ZN(n6525) );
  AND2_X1 U7629 ( .A1(n6532), .A2(n6525), .ZN(n9170) );
  NAND2_X1 U7630 ( .A1(n9170), .A2(n6286), .ZN(n6528) );
  AOI22_X1 U7631 ( .A1(n6482), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n6612), .B2(
        P2_REG0_REG_22__SCAN_IN), .ZN(n6527) );
  NAND2_X1 U7632 ( .A1(n6605), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n6526) );
  NAND2_X1 U7633 ( .A1(n9316), .A2(n9197), .ZN(n6750) );
  NAND2_X1 U7634 ( .A1(n8396), .A2(n5250), .ZN(n6530) );
  NAND2_X1 U7635 ( .A1(n4851), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n6529) );
  INV_X1 U7636 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n9582) );
  NAND2_X1 U7637 ( .A1(n6532), .A2(n9582), .ZN(n6533) );
  NAND2_X1 U7638 ( .A1(n6542), .A2(n6533), .ZN(n9156) );
  OR2_X1 U7639 ( .A1(n9156), .A2(n6574), .ZN(n6539) );
  INV_X1 U7640 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n6536) );
  NAND2_X1 U7641 ( .A1(n6482), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n6535) );
  NAND2_X1 U7642 ( .A1(n6612), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n6534) );
  OAI211_X1 U7643 ( .C1(n6616), .C2(n6536), .A(n6535), .B(n6534), .ZN(n6537)
         );
  INV_X1 U7644 ( .A(n6537), .ZN(n6538) );
  NAND2_X1 U7645 ( .A1(n8447), .A2(n5250), .ZN(n6541) );
  NAND2_X1 U7646 ( .A1(n4852), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n6540) );
  INV_X1 U7647 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n9761) );
  NAND2_X1 U7648 ( .A1(n6542), .A2(n9761), .ZN(n6543) );
  NAND2_X1 U7649 ( .A1(n6552), .A2(n6543), .ZN(n9138) );
  OR2_X1 U7650 ( .A1(n9138), .A2(n6574), .ZN(n6549) );
  INV_X1 U7651 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n6546) );
  NAND2_X1 U7652 ( .A1(n6612), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n6545) );
  NAND2_X1 U7653 ( .A1(n6482), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n6544) );
  OAI211_X1 U7654 ( .C1(n6546), .C2(n6616), .A(n6545), .B(n6544), .ZN(n6547)
         );
  INV_X1 U7655 ( .A(n6547), .ZN(n6548) );
  NAND2_X1 U7656 ( .A1(n9304), .A2(n8868), .ZN(n6640) );
  NAND2_X1 U7657 ( .A1(n6763), .A2(n6640), .ZN(n9141) );
  NAND2_X1 U7658 ( .A1(n4851), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n6551) );
  INV_X1 U7659 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n9672) );
  NAND2_X1 U7660 ( .A1(n6552), .A2(n9672), .ZN(n6553) );
  INV_X1 U7661 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n6556) );
  NAND2_X1 U7662 ( .A1(n6612), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n6555) );
  NAND2_X1 U7663 ( .A1(n6482), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n6554) );
  OAI211_X1 U7664 ( .C1(n6556), .C2(n6616), .A(n6555), .B(n6554), .ZN(n6557)
         );
  NAND2_X1 U7665 ( .A1(n9301), .A2(n9144), .ZN(n6762) );
  NAND2_X1 U7666 ( .A1(n8579), .A2(n5250), .ZN(n6559) );
  NAND2_X1 U7667 ( .A1(n4852), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n6558) );
  INV_X1 U7668 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n9779) );
  NAND2_X1 U7669 ( .A1(n6561), .A2(n9779), .ZN(n6562) );
  NAND2_X1 U7670 ( .A1(n6572), .A2(n6562), .ZN(n9108) );
  INV_X1 U7671 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n6565) );
  NAND2_X1 U7672 ( .A1(n6482), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n6564) );
  NAND2_X1 U7673 ( .A1(n6612), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n6563) );
  OAI211_X1 U7674 ( .C1(n6616), .C2(n6565), .A(n6564), .B(n6563), .ZN(n6566)
         );
  INV_X1 U7675 ( .A(n6566), .ZN(n6567) );
  NAND2_X1 U7676 ( .A1(n9295), .A2(n8829), .ZN(n6791) );
  NAND2_X1 U7677 ( .A1(n10205), .A2(n5250), .ZN(n6570) );
  NAND2_X1 U7678 ( .A1(n4851), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n6569) );
  INV_X1 U7679 ( .A(n6572), .ZN(n6571) );
  NAND2_X1 U7680 ( .A1(n6571), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6586) );
  INV_X1 U7681 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n9735) );
  NAND2_X1 U7682 ( .A1(n6572), .A2(n9735), .ZN(n6573) );
  NAND2_X1 U7683 ( .A1(n6586), .A2(n6573), .ZN(n8830) );
  INV_X1 U7684 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n6577) );
  NAND2_X1 U7685 ( .A1(n6482), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n6576) );
  NAND2_X1 U7686 ( .A1(n6612), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n6575) );
  OAI211_X1 U7687 ( .C1(n6577), .C2(n6616), .A(n6576), .B(n6575), .ZN(n6578)
         );
  INV_X1 U7688 ( .A(n6578), .ZN(n6579) );
  NAND2_X1 U7689 ( .A1(n9289), .A2(n9059), .ZN(n6769) );
  INV_X1 U7690 ( .A(n6768), .ZN(n6581) );
  NAND2_X1 U7691 ( .A1(n4852), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n6583) );
  INV_X1 U7692 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n6585) );
  NAND2_X1 U7693 ( .A1(n6586), .A2(n6585), .ZN(n6587) );
  NAND2_X1 U7694 ( .A1(n9082), .A2(n6286), .ZN(n6593) );
  INV_X1 U7695 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n6590) );
  NAND2_X1 U7696 ( .A1(n6612), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6589) );
  NAND2_X1 U7697 ( .A1(n6482), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n6588) );
  OAI211_X1 U7698 ( .C1(n6590), .C2(n6616), .A(n6589), .B(n6588), .ZN(n6591)
         );
  INV_X1 U7699 ( .A(n6591), .ZN(n6592) );
  NAND2_X1 U7700 ( .A1(n9085), .A2(n6594), .ZN(n9084) );
  NAND2_X1 U7701 ( .A1(n9284), .A2(n9069), .ZN(n6595) );
  NAND2_X1 U7702 ( .A1(n8824), .A2(n5250), .ZN(n6597) );
  NAND2_X1 U7703 ( .A1(n4851), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n6596) );
  INV_X1 U7704 ( .A(n6598), .ZN(n9075) );
  INV_X1 U7705 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n6601) );
  NAND2_X1 U7706 ( .A1(n6612), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6600) );
  NAND2_X1 U7707 ( .A1(n6482), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n6599) );
  OAI211_X1 U7708 ( .C1(n6601), .C2(n6616), .A(n6600), .B(n6599), .ZN(n6602)
         );
  AOI21_X1 U7709 ( .B1(n9075), .B2(n6286), .A(n6602), .ZN(n7876) );
  AND2_X1 U7710 ( .A1(n9280), .A2(n7876), .ZN(n6637) );
  NAND2_X1 U7711 ( .A1(n8790), .A2(n5250), .ZN(n6604) );
  NAND2_X1 U7712 ( .A1(n4851), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n6603) );
  NAND2_X1 U7713 ( .A1(n6612), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n6608) );
  NAND2_X1 U7714 ( .A1(n6482), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n6607) );
  NAND2_X1 U7715 ( .A1(n6605), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n6606) );
  AND3_X1 U7716 ( .A1(n6608), .A2(n6607), .A3(n6606), .ZN(n9067) );
  NOR2_X1 U7717 ( .A1(n9039), .A2(n9067), .ZN(n6634) );
  NAND2_X1 U7718 ( .A1(n6609), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6611) );
  INV_X1 U7719 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n6610) );
  INV_X1 U7720 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n6615) );
  NAND2_X1 U7721 ( .A1(n6482), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n6614) );
  NAND2_X1 U7722 ( .A1(n6612), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n6613) );
  OAI211_X1 U7723 ( .C1(n6616), .C2(n6615), .A(n6614), .B(n6613), .ZN(n8929)
         );
  NAND2_X1 U7724 ( .A1(n6617), .A2(n5151), .ZN(n6618) );
  NAND2_X1 U7725 ( .A1(n6619), .A2(n6618), .ZN(n6623) );
  NAND2_X1 U7726 ( .A1(n9369), .A2(n5250), .ZN(n6621) );
  NAND2_X1 U7727 ( .A1(n4852), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n6620) );
  NAND2_X1 U7728 ( .A1(n6621), .A2(n6620), .ZN(n6781) );
  INV_X1 U7729 ( .A(n8929), .ZN(n6622) );
  NAND2_X1 U7730 ( .A1(n9039), .A2(n9067), .ZN(n6779) );
  AND2_X1 U7731 ( .A1(n6781), .A2(n6622), .ZN(n6633) );
  XNOR2_X1 U7732 ( .A(n6630), .B(n9029), .ZN(n6825) );
  NAND2_X1 U7733 ( .A1(n6626), .A2(n6625), .ZN(n6627) );
  XNOR2_X2 U7734 ( .A(n6629), .B(n6628), .ZN(n6849) );
  INV_X1 U7735 ( .A(n6630), .ZN(n6823) );
  NAND2_X1 U7736 ( .A1(n6632), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6827) );
  NAND2_X1 U7737 ( .A1(n8307), .A2(n8203), .ZN(n7435) );
  INV_X1 U7738 ( .A(n6633), .ZN(n6635) );
  INV_X1 U7739 ( .A(n6634), .ZN(n6780) );
  NAND2_X1 U7740 ( .A1(n6635), .A2(n6780), .ZN(n6789) );
  AND2_X1 U7741 ( .A1(n4849), .A2(n6842), .ZN(n7692) );
  AND2_X1 U7742 ( .A1(n8307), .A2(n7692), .ZN(n6775) );
  INV_X2 U7743 ( .A(n6775), .ZN(n6782) );
  INV_X1 U7744 ( .A(n6637), .ZN(n6777) );
  NAND2_X1 U7745 ( .A1(n6791), .A2(n6762), .ZN(n6638) );
  MUX2_X1 U7746 ( .A(n6638), .B(n4898), .S(n6782), .Z(n6639) );
  INV_X1 U7747 ( .A(n6639), .ZN(n6765) );
  NAND2_X1 U7748 ( .A1(n6763), .A2(n6752), .ZN(n6642) );
  NAND2_X1 U7749 ( .A1(n6640), .A2(n6755), .ZN(n6641) );
  MUX2_X1 U7750 ( .A(n6642), .B(n6641), .S(n6782), .Z(n6643) );
  INV_X1 U7751 ( .A(n6643), .ZN(n6761) );
  NAND2_X1 U7752 ( .A1(n6750), .A2(n6644), .ZN(n6647) );
  NAND2_X1 U7753 ( .A1(n6751), .A2(n6645), .ZN(n6646) );
  MUX2_X1 U7754 ( .A(n6647), .B(n6646), .S(n6775), .Z(n6759) );
  INV_X1 U7755 ( .A(n7565), .ZN(n7852) );
  NAND2_X1 U7756 ( .A1(n6847), .A2(n7852), .ZN(n6795) );
  AND2_X1 U7757 ( .A1(n6796), .A2(n6795), .ZN(n6652) );
  INV_X1 U7758 ( .A(n6652), .ZN(n6648) );
  NAND2_X1 U7759 ( .A1(n6648), .A2(n6797), .ZN(n6650) );
  OAI21_X1 U7760 ( .B1(n7725), .B2(n6650), .A(n6649), .ZN(n6656) );
  INV_X1 U7761 ( .A(n6651), .ZN(n6654) );
  INV_X1 U7762 ( .A(n7725), .ZN(n7694) );
  NAND3_X1 U7763 ( .A1(n7694), .A2(n6842), .A3(n6652), .ZN(n6653) );
  NAND2_X1 U7764 ( .A1(n6654), .A2(n6653), .ZN(n6655) );
  MUX2_X1 U7765 ( .A(n6656), .B(n6655), .S(n6782), .Z(n6660) );
  MUX2_X1 U7766 ( .A(n6658), .B(n6657), .S(n6782), .Z(n6659) );
  OAI21_X1 U7767 ( .B1(n6660), .B2(n7860), .A(n6659), .ZN(n6664) );
  INV_X1 U7768 ( .A(n8943), .ZN(n7777) );
  INV_X1 U7769 ( .A(n10434), .ZN(n10450) );
  NAND2_X1 U7770 ( .A1(n7777), .A2(n10450), .ZN(n6661) );
  MUX2_X1 U7771 ( .A(n6661), .B(n8050), .S(n6782), .Z(n6662) );
  NAND2_X1 U7772 ( .A1(n6662), .A2(n8058), .ZN(n6663) );
  AOI21_X1 U7773 ( .B1(n6664), .B2(n6285), .A(n6663), .ZN(n6669) );
  INV_X1 U7774 ( .A(n6665), .ZN(n6667) );
  MUX2_X1 U7775 ( .A(n6667), .B(n6300), .S(n6782), .Z(n6668) );
  INV_X1 U7776 ( .A(n10509), .ZN(n7871) );
  NOR2_X1 U7777 ( .A1(n8941), .A2(n7871), .ZN(n6800) );
  MUX2_X1 U7778 ( .A(n8941), .B(n7871), .S(n6782), .Z(n6670) );
  OAI22_X1 U7779 ( .A1(n6669), .A2(n6668), .B1(n6800), .B2(n6670), .ZN(n6672)
         );
  NAND2_X1 U7780 ( .A1(n8941), .A2(n7871), .ZN(n7962) );
  NAND2_X1 U7781 ( .A1(n6670), .A2(n7962), .ZN(n6671) );
  AOI21_X1 U7782 ( .B1(n6672), .B2(n6671), .A(n7963), .ZN(n6679) );
  MUX2_X1 U7783 ( .A(n6673), .B(n7949), .S(n6775), .Z(n6674) );
  NAND2_X1 U7784 ( .A1(n6674), .A2(n4975), .ZN(n6678) );
  MUX2_X1 U7785 ( .A(n6676), .B(n6675), .S(n6782), .Z(n6677) );
  OAI211_X1 U7786 ( .C1(n6679), .C2(n6678), .A(n6680), .B(n6677), .ZN(n6693)
         );
  NAND2_X1 U7787 ( .A1(n6688), .A2(n6680), .ZN(n6682) );
  INV_X1 U7788 ( .A(n6686), .ZN(n6681) );
  MUX2_X1 U7789 ( .A(n6682), .B(n6681), .S(n6782), .Z(n6683) );
  INV_X1 U7790 ( .A(n6683), .ZN(n6684) );
  NAND2_X1 U7791 ( .A1(n6684), .A2(n6685), .ZN(n6687) );
  INV_X1 U7792 ( .A(n6687), .ZN(n6692) );
  INV_X1 U7793 ( .A(n6694), .ZN(n6793) );
  OAI211_X1 U7794 ( .C1(n6687), .C2(n6686), .A(n6793), .B(n6685), .ZN(n6690)
         );
  NAND2_X1 U7795 ( .A1(n6794), .A2(n6688), .ZN(n6689) );
  MUX2_X1 U7796 ( .A(n6690), .B(n6689), .S(n6782), .Z(n6691) );
  AOI211_X1 U7797 ( .C1(n6693), .C2(n6692), .A(n6691), .B(n8284), .ZN(n6703)
         );
  NAND2_X1 U7798 ( .A1(n6698), .A2(n6694), .ZN(n6695) );
  NAND2_X1 U7799 ( .A1(n6695), .A2(n6697), .ZN(n6701) );
  INV_X1 U7800 ( .A(n6794), .ZN(n6696) );
  NAND2_X1 U7801 ( .A1(n6697), .A2(n6696), .ZN(n6699) );
  NAND2_X1 U7802 ( .A1(n6699), .A2(n6698), .ZN(n6700) );
  MUX2_X1 U7803 ( .A(n6701), .B(n6700), .S(n6775), .Z(n6702) );
  INV_X1 U7804 ( .A(n6704), .ZN(n6707) );
  INV_X1 U7805 ( .A(n6705), .ZN(n6706) );
  MUX2_X1 U7806 ( .A(n6707), .B(n6706), .S(n6782), .Z(n6708) );
  NOR2_X1 U7807 ( .A1(n8493), .A2(n6708), .ZN(n6709) );
  NAND2_X1 U7808 ( .A1(n6710), .A2(n6709), .ZN(n6714) );
  MUX2_X1 U7809 ( .A(n6712), .B(n6711), .S(n6782), .Z(n6713) );
  NAND3_X1 U7810 ( .A1(n6714), .A2(n8538), .A3(n6713), .ZN(n6721) );
  INV_X1 U7811 ( .A(n6715), .ZN(n6718) );
  INV_X1 U7812 ( .A(n6716), .ZN(n6717) );
  MUX2_X1 U7813 ( .A(n6718), .B(n6717), .S(n6782), .Z(n6719) );
  INV_X1 U7814 ( .A(n6719), .ZN(n6720) );
  NAND3_X1 U7815 ( .A1(n6721), .A2(n8541), .A3(n6720), .ZN(n6723) );
  MUX2_X1 U7816 ( .A(n9257), .B(n9256), .S(n6782), .Z(n6722) );
  NAND2_X1 U7817 ( .A1(n6723), .A2(n6722), .ZN(n6726) );
  MUX2_X1 U7818 ( .A(n8933), .B(n9343), .S(n6782), .Z(n6724) );
  OAI21_X1 U7819 ( .B1(n6726), .B2(n6725), .A(n6724), .ZN(n6728) );
  NAND2_X1 U7820 ( .A1(n6726), .A2(n5338), .ZN(n6727) );
  NAND2_X1 U7821 ( .A1(n6728), .A2(n6727), .ZN(n6741) );
  MUX2_X1 U7822 ( .A(n9336), .B(n8932), .S(n6782), .Z(n6739) );
  INV_X1 U7823 ( .A(n6739), .ZN(n6729) );
  OR2_X1 U7824 ( .A1(n6741), .A2(n6729), .ZN(n6735) );
  AND2_X1 U7825 ( .A1(n6732), .A2(n8932), .ZN(n6730) );
  AOI21_X1 U7826 ( .B1(n6735), .B2(n6730), .A(n5213), .ZN(n6737) );
  AND2_X1 U7827 ( .A1(n6731), .A2(n9336), .ZN(n6734) );
  INV_X1 U7828 ( .A(n6732), .ZN(n6733) );
  AOI21_X1 U7829 ( .B1(n6735), .B2(n6734), .A(n6733), .ZN(n6736) );
  MUX2_X1 U7830 ( .A(n6737), .B(n6736), .S(n6782), .Z(n6749) );
  NOR2_X1 U7831 ( .A1(n9224), .A2(n6739), .ZN(n6740) );
  AOI21_X1 U7832 ( .B1(n6741), .B2(n6740), .A(n9212), .ZN(n6748) );
  INV_X1 U7833 ( .A(n6742), .ZN(n6745) );
  INV_X1 U7834 ( .A(n6743), .ZN(n6744) );
  MUX2_X1 U7835 ( .A(n6745), .B(n6744), .S(n6782), .Z(n6746) );
  OR2_X1 U7836 ( .A1(n9051), .A2(n6746), .ZN(n6747) );
  AOI21_X1 U7837 ( .B1(n6749), .B2(n6748), .A(n6747), .ZN(n6758) );
  INV_X1 U7838 ( .A(n6750), .ZN(n6754) );
  NAND2_X1 U7839 ( .A1(n6752), .A2(n6751), .ZN(n6753) );
  MUX2_X1 U7840 ( .A(n6754), .B(n6753), .S(n6782), .Z(n6756) );
  NOR2_X1 U7841 ( .A1(n6756), .A2(n5224), .ZN(n6757) );
  OAI21_X1 U7842 ( .B1(n6759), .B2(n6758), .A(n6757), .ZN(n6760) );
  NAND2_X1 U7843 ( .A1(n6761), .A2(n6760), .ZN(n6764) );
  MUX2_X1 U7844 ( .A(n6792), .B(n6791), .S(n6782), .Z(n6766) );
  NAND2_X1 U7845 ( .A1(n6767), .A2(n9099), .ZN(n6771) );
  MUX2_X1 U7846 ( .A(n6769), .B(n6768), .S(n6775), .Z(n6770) );
  NAND3_X1 U7847 ( .A1(n6771), .A2(n6594), .A3(n6770), .ZN(n6774) );
  OR3_X1 U7848 ( .A1(n9284), .A2(n9069), .A3(n6775), .ZN(n6773) );
  NAND3_X1 U7849 ( .A1(n9284), .A2(n9069), .A3(n6775), .ZN(n6772) );
  MUX2_X1 U7850 ( .A(n6777), .B(n6776), .S(n6775), .Z(n6778) );
  MUX2_X1 U7851 ( .A(n8929), .B(n6781), .S(n6782), .Z(n6784) );
  NOR2_X1 U7852 ( .A1(n6781), .A2(n8929), .ZN(n6783) );
  OR2_X1 U7853 ( .A1(n6784), .A2(n6783), .ZN(n6785) );
  NAND2_X1 U7854 ( .A1(n6848), .A2(n4849), .ZN(n7429) );
  XNOR2_X1 U7855 ( .A(n6788), .B(n7429), .ZN(n6787) );
  NAND3_X1 U7856 ( .A1(n6787), .A2(n6849), .A3(n7435), .ZN(n6822) );
  NAND2_X1 U7857 ( .A1(n6788), .A2(n6849), .ZN(n6820) );
  INV_X1 U7858 ( .A(n6789), .ZN(n6817) );
  INV_X1 U7859 ( .A(n9237), .ZN(n9246) );
  INV_X1 U7860 ( .A(n8538), .ZN(n6807) );
  INV_X1 U7861 ( .A(n8284), .ZN(n8283) );
  NAND3_X1 U7862 ( .A1(n7694), .A2(n7730), .A3(n8058), .ZN(n6799) );
  AND2_X1 U7863 ( .A1(n7562), .A2(n6795), .ZN(n7857) );
  AND2_X1 U7864 ( .A1(n6797), .A2(n6796), .ZN(n7561) );
  NOR2_X1 U7865 ( .A1(n6799), .A2(n6798), .ZN(n6801) );
  INV_X1 U7866 ( .A(n6800), .ZN(n7975) );
  NAND2_X1 U7867 ( .A1(n7975), .A2(n7962), .ZN(n7866) );
  NAND4_X1 U7868 ( .A1(n6801), .A2(n6329), .A3(n6285), .A4(n7866), .ZN(n6803)
         );
  INV_X1 U7869 ( .A(n10610), .ZN(n10601) );
  NOR4_X1 U7870 ( .A1(n6803), .A2(n6802), .A3(n8136), .A4(n10601), .ZN(n6804)
         );
  NAND4_X1 U7871 ( .A1(n6805), .A2(n8283), .A3(n8236), .A4(n6804), .ZN(n6806)
         );
  NOR3_X1 U7872 ( .A1(n6807), .A2(n8493), .A3(n6806), .ZN(n6808) );
  NAND3_X1 U7873 ( .A1(n9045), .A2(n8541), .A3(n6808), .ZN(n6809) );
  NOR3_X1 U7874 ( .A1(n9224), .A2(n9246), .A3(n6809), .ZN(n6810) );
  NAND2_X1 U7875 ( .A1(n6811), .A2(n6810), .ZN(n6812) );
  NOR4_X1 U7876 ( .A1(n9162), .A2(n5225), .A3(n9051), .A4(n6812), .ZN(n6813)
         );
  NAND4_X1 U7877 ( .A1(n9115), .A2(n6550), .A3(n9124), .A4(n6813), .ZN(n6814)
         );
  NOR4_X1 U7878 ( .A1(n9064), .A2(n6814), .A3(n9060), .A4(n9058), .ZN(n6815)
         );
  NAND3_X1 U7879 ( .A1(n6817), .A2(n6816), .A3(n6815), .ZN(n6818) );
  XNOR2_X1 U7880 ( .A(n6818), .B(n4849), .ZN(n6819) );
  NAND3_X1 U7881 ( .A1(n6820), .A2(n6819), .A3(n8203), .ZN(n6821) );
  OAI211_X1 U7882 ( .C1(n6823), .C2(n6975), .A(n6822), .B(n6821), .ZN(n6824)
         );
  AOI21_X1 U7883 ( .B1(n6825), .B2(n7431), .A(n6824), .ZN(n6846) );
  NAND2_X1 U7884 ( .A1(n6827), .A2(n6826), .ZN(n6828) );
  NAND2_X1 U7885 ( .A1(n6828), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6835) );
  XNOR2_X1 U7886 ( .A(n6835), .B(n6834), .ZN(n7010) );
  OR2_X1 U7887 ( .A1(n7010), .A2(P2_U3152), .ZN(n8383) );
  NOR2_X1 U7888 ( .A1(n6829), .A2(n9370), .ZN(n6830) );
  MUX2_X1 U7889 ( .A(n9370), .B(n6830), .S(P2_IR_REG_25__SCAN_IN), .Z(n6831)
         );
  INV_X1 U7890 ( .A(n6831), .ZN(n6833) );
  NAND2_X1 U7891 ( .A1(n6833), .A2(n6832), .ZN(n8576) );
  INV_X1 U7892 ( .A(n8576), .ZN(n6839) );
  NAND2_X1 U7893 ( .A1(n6835), .A2(n6834), .ZN(n6836) );
  NAND2_X1 U7894 ( .A1(n6836), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6837) );
  NAND2_X1 U7895 ( .A1(n6832), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6838) );
  INV_X1 U7896 ( .A(n10312), .ZN(n6840) );
  NOR4_X1 U7897 ( .A1(n7442), .A2(n10611), .A3(n9385), .A4(n7009), .ZN(n6844)
         );
  OAI21_X1 U7898 ( .B1(n8383), .B2(n6848), .A(P2_B_REG_SCAN_IN), .ZN(n6843) );
  OR2_X1 U7899 ( .A1(n6844), .A2(n6843), .ZN(n6845) );
  OAI21_X1 U7900 ( .B1(n6846), .B2(n8383), .A(n6845), .ZN(P2_U3244) );
  INV_X1 U7901 ( .A(n7485), .ZN(n6847) );
  NAND2_X1 U7902 ( .A1(n6851), .A2(n6850), .ZN(n6853) );
  AND2_X1 U7903 ( .A1(n7435), .A2(n9029), .ZN(n6852) );
  NAND2_X1 U7904 ( .A1(n7852), .A2(n6976), .ZN(n6855) );
  NAND2_X1 U7905 ( .A1(n8946), .A2(n6975), .ZN(n6858) );
  XNOR2_X1 U7906 ( .A(n6858), .B(n6856), .ZN(n7483) );
  INV_X1 U7907 ( .A(n6856), .ZN(n6857) );
  NAND2_X1 U7908 ( .A1(n6858), .A2(n6857), .ZN(n6859) );
  NAND2_X1 U7909 ( .A1(n6861), .A2(n6862), .ZN(n6865) );
  INV_X1 U7910 ( .A(n6861), .ZN(n6863) );
  INV_X1 U7911 ( .A(n6862), .ZN(n7605) );
  NAND2_X1 U7912 ( .A1(n6863), .A2(n7605), .ZN(n6864) );
  NOR2_X1 U7913 ( .A1(n10438), .A2(n7701), .ZN(n6866) );
  XNOR2_X1 U7914 ( .A(n7738), .B(n6960), .ZN(n6867) );
  NAND2_X1 U7915 ( .A1(n6866), .A2(n6867), .ZN(n6870) );
  INV_X1 U7916 ( .A(n6866), .ZN(n6868) );
  INV_X1 U7917 ( .A(n6867), .ZN(n7783) );
  NAND2_X1 U7918 ( .A1(n6868), .A2(n7783), .ZN(n6869) );
  NAND2_X1 U7919 ( .A1(n8943), .A2(n6975), .ZN(n6873) );
  XNOR2_X1 U7920 ( .A(n6872), .B(n6873), .ZN(n7784) );
  AND2_X1 U7921 ( .A1(n7784), .A2(n6870), .ZN(n6871) );
  INV_X1 U7922 ( .A(n6872), .ZN(n7776) );
  NAND2_X1 U7923 ( .A1(n7776), .A2(n6873), .ZN(n6874) );
  NAND2_X1 U7924 ( .A1(n8942), .A2(n6975), .ZN(n6876) );
  XNOR2_X1 U7925 ( .A(n10473), .B(n6960), .ZN(n6875) );
  XNOR2_X1 U7926 ( .A(n6876), .B(n6875), .ZN(n7775) );
  INV_X1 U7927 ( .A(n6875), .ZN(n7825) );
  NAND2_X1 U7928 ( .A1(n6876), .A2(n7825), .ZN(n6877) );
  XNOR2_X1 U7929 ( .A(n10509), .B(n6976), .ZN(n6878) );
  NAND2_X1 U7930 ( .A1(n8941), .A2(n6975), .ZN(n6879) );
  INV_X1 U7931 ( .A(n6878), .ZN(n6880) );
  NAND2_X1 U7932 ( .A1(n6880), .A2(n6879), .ZN(n6881) );
  NOR2_X1 U7933 ( .A1(n8065), .A2(n7701), .ZN(n6882) );
  XNOR2_X1 U7934 ( .A(n10525), .B(n6960), .ZN(n6883) );
  NAND2_X1 U7935 ( .A1(n6882), .A2(n6883), .ZN(n6887) );
  INV_X1 U7936 ( .A(n6882), .ZN(n6884) );
  INV_X1 U7937 ( .A(n6883), .ZN(n8064) );
  NAND2_X1 U7938 ( .A1(n6884), .A2(n8064), .ZN(n6885) );
  NAND2_X1 U7939 ( .A1(n6887), .A2(n6885), .ZN(n7145) );
  NOR2_X1 U7940 ( .A1(n8175), .A2(n7701), .ZN(n6888) );
  XNOR2_X1 U7941 ( .A(n8131), .B(n6960), .ZN(n6889) );
  NAND2_X1 U7942 ( .A1(n6888), .A2(n6889), .ZN(n6892) );
  INV_X1 U7943 ( .A(n6888), .ZN(n6890) );
  INV_X1 U7944 ( .A(n6889), .ZN(n8168) );
  NAND2_X1 U7945 ( .A1(n6890), .A2(n8168), .ZN(n6891) );
  AND2_X1 U7946 ( .A1(n6892), .A2(n6891), .ZN(n8062) );
  NAND2_X1 U7947 ( .A1(n8939), .A2(n6975), .ZN(n6896) );
  XNOR2_X1 U7948 ( .A(n8179), .B(n6960), .ZN(n6894) );
  XNOR2_X1 U7949 ( .A(n6896), .B(n6894), .ZN(n8182) );
  AND2_X1 U7950 ( .A1(n8182), .A2(n6892), .ZN(n6893) );
  INV_X1 U7951 ( .A(n6894), .ZN(n6895) );
  NAND2_X1 U7952 ( .A1(n6896), .A2(n6895), .ZN(n6897) );
  XNOR2_X1 U7953 ( .A(n10606), .B(n6960), .ZN(n6898) );
  NOR2_X1 U7954 ( .A1(n8246), .A2(n7701), .ZN(n6899) );
  NAND2_X1 U7955 ( .A1(n6898), .A2(n6899), .ZN(n6902) );
  INV_X1 U7956 ( .A(n6898), .ZN(n8247) );
  INV_X1 U7957 ( .A(n6899), .ZN(n6900) );
  NAND2_X1 U7958 ( .A1(n8247), .A2(n6900), .ZN(n6901) );
  NAND2_X1 U7959 ( .A1(n6902), .A2(n6901), .ZN(n8843) );
  XNOR2_X1 U7960 ( .A(n10640), .B(n6960), .ZN(n6903) );
  NOR2_X1 U7961 ( .A1(n10614), .A2(n7701), .ZN(n6904) );
  NAND2_X1 U7962 ( .A1(n6903), .A2(n6904), .ZN(n6907) );
  INV_X1 U7963 ( .A(n6903), .ZN(n8401) );
  INV_X1 U7964 ( .A(n6904), .ZN(n6905) );
  NAND2_X1 U7965 ( .A1(n8401), .A2(n6905), .ZN(n6906) );
  AND2_X1 U7966 ( .A1(n6907), .A2(n6906), .ZN(n8245) );
  XNOR2_X1 U7967 ( .A(n8411), .B(n6976), .ZN(n8317) );
  NOR2_X1 U7968 ( .A1(n8374), .A2(n7701), .ZN(n6909) );
  XNOR2_X1 U7969 ( .A(n8317), .B(n6909), .ZN(n8414) );
  AND2_X1 U7970 ( .A1(n8414), .A2(n6907), .ZN(n6908) );
  INV_X1 U7971 ( .A(n6909), .ZN(n6910) );
  XNOR2_X1 U7972 ( .A(n8371), .B(n6976), .ZN(n8391) );
  NOR2_X1 U7973 ( .A1(n8504), .A2(n7701), .ZN(n6911) );
  XNOR2_X1 U7974 ( .A(n8391), .B(n6911), .ZN(n8316) );
  INV_X1 U7975 ( .A(n6911), .ZN(n6912) );
  XNOR2_X1 U7976 ( .A(n10661), .B(n6976), .ZN(n8784) );
  NOR2_X1 U7977 ( .A1(n8783), .A2(n7701), .ZN(n6914) );
  XNOR2_X1 U7978 ( .A(n8784), .B(n6914), .ZN(n8390) );
  INV_X1 U7979 ( .A(n6914), .ZN(n6915) );
  NAND2_X1 U7980 ( .A1(n8784), .A2(n6915), .ZN(n6916) );
  NAND2_X1 U7981 ( .A1(n8386), .A2(n6916), .ZN(n6917) );
  XNOR2_X1 U7982 ( .A(n8781), .B(n6976), .ZN(n8457) );
  NOR2_X1 U7983 ( .A1(n8505), .A2(n7701), .ZN(n6918) );
  XNOR2_X1 U7984 ( .A(n8457), .B(n6918), .ZN(n8782) );
  INV_X1 U7985 ( .A(n6918), .ZN(n6919) );
  NAND2_X1 U7986 ( .A1(n8457), .A2(n6919), .ZN(n6920) );
  NAND2_X1 U7987 ( .A1(n8789), .A2(n6920), .ZN(n6921) );
  XNOR2_X1 U7988 ( .A(n9349), .B(n6976), .ZN(n6924) );
  NOR2_X1 U7989 ( .A1(n8775), .A2(n7701), .ZN(n6922) );
  XNOR2_X1 U7990 ( .A(n6924), .B(n6922), .ZN(n8456) );
  INV_X1 U7991 ( .A(n6922), .ZN(n6923) );
  NAND2_X1 U7992 ( .A1(n6924), .A2(n6923), .ZN(n6925) );
  XNOR2_X1 U7993 ( .A(n9343), .B(n6976), .ZN(n6927) );
  NAND2_X1 U7994 ( .A1(n8933), .A2(n6975), .ZN(n6928) );
  AND2_X1 U7995 ( .A1(n6927), .A2(n6928), .ZN(n8565) );
  INV_X1 U7996 ( .A(n8565), .ZN(n6926) );
  INV_X1 U7997 ( .A(n6927), .ZN(n6930) );
  INV_X1 U7998 ( .A(n6928), .ZN(n6929) );
  NAND2_X1 U7999 ( .A1(n6930), .A2(n6929), .ZN(n8566) );
  XNOR2_X1 U8000 ( .A(n9336), .B(n6976), .ZN(n8903) );
  NAND2_X1 U8001 ( .A1(n8932), .A2(n6975), .ZN(n6931) );
  NAND2_X1 U8002 ( .A1(n8903), .A2(n6931), .ZN(n8908) );
  INV_X1 U8003 ( .A(n8903), .ZN(n6933) );
  INV_X1 U8004 ( .A(n6931), .ZN(n6932) );
  NAND2_X1 U8005 ( .A1(n6933), .A2(n6932), .ZN(n8909) );
  NAND2_X1 U8006 ( .A1(n8906), .A2(n8909), .ZN(n8853) );
  XNOR2_X1 U8007 ( .A(n9333), .B(n6976), .ZN(n6934) );
  NOR2_X1 U8008 ( .A1(n9248), .A2(n7701), .ZN(n6935) );
  XNOR2_X1 U8009 ( .A(n6934), .B(n6935), .ZN(n8852) );
  NAND2_X1 U8010 ( .A1(n8853), .A2(n8852), .ZN(n6938) );
  INV_X1 U8011 ( .A(n6934), .ZN(n6936) );
  NAND2_X1 U8012 ( .A1(n6936), .A2(n6935), .ZN(n6937) );
  NAND2_X1 U8013 ( .A1(n6938), .A2(n6937), .ZN(n8884) );
  XNOR2_X1 U8014 ( .A(n9326), .B(n6976), .ZN(n6939) );
  NOR2_X1 U8015 ( .A1(n9196), .A2(n7701), .ZN(n6940) );
  XNOR2_X1 U8016 ( .A(n6939), .B(n6940), .ZN(n8885) );
  NAND2_X1 U8017 ( .A1(n8884), .A2(n8885), .ZN(n6943) );
  INV_X1 U8018 ( .A(n6939), .ZN(n6941) );
  NAND2_X1 U8019 ( .A1(n6941), .A2(n6940), .ZN(n6942) );
  NAND2_X1 U8020 ( .A1(n6943), .A2(n6942), .ZN(n8858) );
  XNOR2_X1 U8021 ( .A(n9321), .B(n6976), .ZN(n6944) );
  NOR2_X1 U8022 ( .A1(n9214), .A2(n7701), .ZN(n6945) );
  XNOR2_X1 U8023 ( .A(n6944), .B(n6945), .ZN(n8859) );
  INV_X1 U8024 ( .A(n6944), .ZN(n6946) );
  NAND2_X1 U8025 ( .A1(n6946), .A2(n6945), .ZN(n6947) );
  XNOR2_X1 U8026 ( .A(n9316), .B(n6976), .ZN(n6948) );
  OR2_X1 U8027 ( .A1(n9197), .A2(n7701), .ZN(n6949) );
  NAND2_X1 U8028 ( .A1(n6948), .A2(n6949), .ZN(n6954) );
  INV_X1 U8029 ( .A(n6948), .ZN(n6951) );
  INV_X1 U8030 ( .A(n6949), .ZN(n6950) );
  NAND2_X1 U8031 ( .A1(n6951), .A2(n6950), .ZN(n6952) );
  NAND2_X1 U8032 ( .A1(n6954), .A2(n6952), .ZN(n8893) );
  NAND2_X1 U8033 ( .A1(n8891), .A2(n6954), .ZN(n6958) );
  XNOR2_X1 U8034 ( .A(n9159), .B(n6960), .ZN(n6956) );
  NAND2_X1 U8035 ( .A1(n9179), .A2(n6975), .ZN(n6955) );
  INV_X1 U8036 ( .A(n6956), .ZN(n6957) );
  NAND2_X1 U8037 ( .A1(n6958), .A2(n6957), .ZN(n6959) );
  NAND2_X1 U8038 ( .A1(n8842), .A2(n6959), .ZN(n6963) );
  XNOR2_X1 U8039 ( .A(n9304), .B(n6960), .ZN(n6961) );
  XNOR2_X1 U8040 ( .A(n6963), .B(n6961), .ZN(n8877) );
  NOR2_X1 U8041 ( .A1(n8868), .A2(n7701), .ZN(n8876) );
  INV_X1 U8042 ( .A(n6961), .ZN(n6962) );
  OR2_X1 U8043 ( .A1(n6963), .A2(n6962), .ZN(n6964) );
  XNOR2_X1 U8044 ( .A(n9301), .B(n6976), .ZN(n6965) );
  OR2_X1 U8045 ( .A1(n9144), .A2(n7701), .ZN(n6966) );
  NAND2_X1 U8046 ( .A1(n6965), .A2(n6966), .ZN(n8865) );
  INV_X1 U8047 ( .A(n6965), .ZN(n6968) );
  INV_X1 U8048 ( .A(n6966), .ZN(n6967) );
  NAND2_X1 U8049 ( .A1(n6968), .A2(n6967), .ZN(n8864) );
  XNOR2_X1 U8050 ( .A(n9295), .B(n6976), .ZN(n6969) );
  NOR2_X1 U8051 ( .A1(n8829), .A2(n7701), .ZN(n6970) );
  XNOR2_X1 U8052 ( .A(n6969), .B(n6970), .ZN(n8919) );
  INV_X1 U8053 ( .A(n6969), .ZN(n6971) );
  XNOR2_X1 U8054 ( .A(n9289), .B(n6976), .ZN(n6972) );
  NOR2_X1 U8055 ( .A1(n9059), .A2(n7701), .ZN(n6973) );
  XNOR2_X1 U8056 ( .A(n6972), .B(n6973), .ZN(n8827) );
  INV_X1 U8057 ( .A(n6972), .ZN(n6974) );
  NAND2_X1 U8058 ( .A1(n9100), .A2(n6975), .ZN(n6977) );
  MUX2_X1 U8059 ( .A(n9100), .B(n6977), .S(n6976), .Z(n6999) );
  NOR4_X1 U8060 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n6981) );
  NOR4_X1 U8061 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n6980) );
  NOR4_X1 U8062 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6979) );
  NOR4_X1 U8063 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n6978) );
  NAND4_X1 U8064 ( .A1(n6981), .A2(n6980), .A3(n6979), .A4(n6978), .ZN(n6989)
         );
  NOR2_X1 U8065 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .ZN(
        n6985) );
  NOR4_X1 U8066 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n6984) );
  NOR4_X1 U8067 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n6983) );
  NOR4_X1 U8068 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n6982) );
  NAND4_X1 U8069 ( .A1(n6985), .A2(n6984), .A3(n6983), .A4(n6982), .ZN(n6988)
         );
  INV_X1 U8070 ( .A(n10308), .ZN(n8449) );
  INV_X1 U8071 ( .A(P2_B_REG_SCAN_IN), .ZN(n6986) );
  OAI221_X1 U8072 ( .B1(n10308), .B2(P2_B_REG_SCAN_IN), .C1(n8449), .C2(n6986), 
        .A(n8576), .ZN(n6987) );
  OAI21_X1 U8073 ( .B1(n6989), .B2(n6988), .A(n10212), .ZN(n7427) );
  INV_X1 U8074 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n10310) );
  NAND2_X1 U8075 ( .A1(n10212), .A2(n10310), .ZN(n6991) );
  OR2_X1 U8076 ( .A1(n10308), .A2(n10307), .ZN(n6990) );
  INV_X1 U8077 ( .A(n10307), .ZN(n8581) );
  AND2_X1 U8078 ( .A1(n8581), .A2(n8576), .ZN(n10215) );
  INV_X1 U8079 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n10216) );
  AND2_X1 U8080 ( .A1(n10212), .A2(n10216), .ZN(n6992) );
  INV_X1 U8081 ( .A(n7441), .ZN(n7690) );
  INV_X1 U8082 ( .A(n7435), .ZN(n7567) );
  NOR2_X1 U8083 ( .A1(n7442), .A2(n7699), .ZN(n6993) );
  NAND2_X1 U8084 ( .A1(n7007), .A2(n6993), .ZN(n6996) );
  AND2_X1 U8085 ( .A1(n8307), .A2(n4849), .ZN(n6994) );
  NAND2_X1 U8086 ( .A1(n10622), .A2(n8203), .ZN(n7440) );
  INV_X1 U8087 ( .A(n7440), .ZN(n6995) );
  NOR3_X1 U8088 ( .A1(n5155), .A2(n6999), .A3(n8915), .ZN(n6997) );
  AOI21_X1 U8089 ( .B1(n5155), .B2(n6999), .A(n6997), .ZN(n7005) );
  NAND3_X1 U8090 ( .A1(n9284), .A2(n8922), .A3(n6999), .ZN(n6998) );
  OAI21_X1 U8091 ( .B1(n6999), .B2(n9284), .A(n6998), .ZN(n7000) );
  NAND2_X1 U8092 ( .A1(n9284), .A2(n8915), .ZN(n7003) );
  INV_X1 U8093 ( .A(n7180), .ZN(n7159) );
  OR2_X1 U8094 ( .A1(n10662), .A2(n7159), .ZN(n7001) );
  NOR2_X1 U8095 ( .A1(n7442), .A2(n7001), .ZN(n7002) );
  INV_X2 U8096 ( .A(n8905), .ZN(n8927) );
  NAND2_X1 U8097 ( .A1(n7003), .A2(n8927), .ZN(n7004) );
  OAI22_X1 U8098 ( .A1(n7876), .A2(n10613), .B1(n9059), .B2(n10611), .ZN(n9086) );
  INV_X1 U8099 ( .A(n9086), .ZN(n7015) );
  NOR2_X1 U8100 ( .A1(n7442), .A2(n7009), .ZN(n7006) );
  NAND2_X1 U8101 ( .A1(n7007), .A2(n7006), .ZN(n8871) );
  INV_X1 U8102 ( .A(n7007), .ZN(n7008) );
  NAND2_X1 U8103 ( .A1(n7008), .A2(n7440), .ZN(n7013) );
  NAND2_X1 U8104 ( .A1(n7159), .A2(n7009), .ZN(n7439) );
  NAND2_X1 U8105 ( .A1(n7439), .A2(n7010), .ZN(n7011) );
  NOR2_X1 U8106 ( .A1(n7157), .A2(n7011), .ZN(n7012) );
  NAND2_X1 U8107 ( .A1(n7013), .A2(n7012), .ZN(n7397) );
  AOI22_X1 U8108 ( .A1(n9082), .A2(n8910), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        n4846), .ZN(n7014) );
  INV_X1 U8109 ( .A(n7016), .ZN(n7017) );
  NAND2_X1 U8110 ( .A1(n7018), .A2(n7017), .ZN(P2_U3222) );
  NAND2_X1 U8111 ( .A1(n7129), .A2(n9991), .ZN(n7020) );
  OR2_X1 U8112 ( .A1(n8185), .A2(n8166), .ZN(n7019) );
  NAND2_X1 U8113 ( .A1(n7020), .A2(n7019), .ZN(n10546) );
  INV_X1 U8114 ( .A(n10546), .ZN(n7060) );
  INV_X1 U8115 ( .A(n8009), .ZN(n7024) );
  AND2_X1 U8116 ( .A1(n10542), .A2(n7025), .ZN(n7026) );
  NAND2_X1 U8117 ( .A1(n10543), .A2(n7026), .ZN(n8077) );
  NAND2_X1 U8118 ( .A1(n8077), .A2(n7027), .ZN(n7029) );
  NAND2_X1 U8119 ( .A1(n7029), .A2(n7028), .ZN(n8187) );
  NAND2_X1 U8120 ( .A1(n8293), .A2(n8295), .ZN(n7034) );
  NAND2_X1 U8121 ( .A1(n7034), .A2(n7033), .ZN(n8339) );
  INV_X1 U8122 ( .A(n8343), .ZN(n8338) );
  NAND2_X1 U8123 ( .A1(n8339), .A2(n8338), .ZN(n7036) );
  INV_X1 U8124 ( .A(n8521), .ZN(n7038) );
  NAND2_X1 U8125 ( .A1(n7038), .A2(n8518), .ZN(n8524) );
  INV_X1 U8126 ( .A(n7040), .ZN(n7042) );
  NAND2_X1 U8127 ( .A1(n10034), .A2(n7044), .ZN(n10020) );
  NAND2_X1 U8128 ( .A1(n7048), .A2(n7047), .ZN(n9968) );
  NAND2_X1 U8129 ( .A1(n9968), .A2(n7049), .ZN(n7051) );
  NAND2_X1 U8130 ( .A1(n8809), .A2(n7057), .ZN(n7058) );
  NAND2_X1 U8131 ( .A1(n6205), .A2(n7385), .ZN(n10489) );
  INV_X1 U8132 ( .A(n6205), .ZN(n7465) );
  INV_X1 U8133 ( .A(n10540), .ZN(n7059) );
  NAND2_X1 U8134 ( .A1(n10357), .A2(n7759), .ZN(n7758) );
  NAND2_X1 U8135 ( .A1(n7749), .A2(n7633), .ZN(n10400) );
  OR2_X1 U8136 ( .A1(n10400), .A2(n9496), .ZN(n10401) );
  INV_X1 U8137 ( .A(n8276), .ZN(n8198) );
  INV_X1 U8138 ( .A(n10168), .ZN(n8337) );
  NAND2_X1 U8139 ( .A1(n8212), .A2(n8337), .ZN(n8298) );
  INV_X1 U8140 ( .A(n10152), .ZN(n9407) );
  INV_X1 U8141 ( .A(n10146), .ZN(n8532) );
  INV_X1 U8142 ( .A(n10123), .ZN(n10018) );
  NAND2_X1 U8143 ( .A1(n10039), .A2(n10018), .ZN(n10013) );
  INV_X1 U8144 ( .A(n10113), .ZN(n7062) );
  INV_X1 U8145 ( .A(n10097), .ZN(n9489) );
  NAND2_X1 U8146 ( .A1(n9549), .A2(n9916), .ZN(n8595) );
  NAND2_X1 U8147 ( .A1(n8311), .A2(n8185), .ZN(n7627) );
  AOI211_X1 U8148 ( .C1(n10082), .C2(n8595), .A(n10582), .B(n8801), .ZN(n10081) );
  INV_X2 U8149 ( .A(n10005), .ZN(n10561) );
  AOI22_X1 U8150 ( .A1(n10081), .A2(n8116), .B1(n10561), .B2(n9393), .ZN(n7083) );
  NAND2_X1 U8151 ( .A1(n8452), .A2(P1_B_REG_SCAN_IN), .ZN(n7065) );
  OAI22_X1 U8152 ( .A1(n7080), .A2(n7065), .B1(P1_B_REG_SCAN_IN), .B2(n8452), 
        .ZN(n7067) );
  INV_X1 U8153 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n7068) );
  NAND2_X1 U8154 ( .A1(n7405), .A2(n7068), .ZN(n7069) );
  NAND2_X1 U8155 ( .A1(n7066), .A2(n8452), .ZN(n10194) );
  AND2_X1 U8156 ( .A1(n7385), .A2(n7668), .ZN(n7650) );
  INV_X1 U8157 ( .A(n7409), .ZN(n7391) );
  NOR4_X1 U8158 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n7073) );
  NOR4_X1 U8159 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n7072) );
  NOR4_X1 U8160 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n7071) );
  NOR4_X1 U8161 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n7070) );
  AND4_X1 U8162 ( .A1(n7073), .A2(n7072), .A3(n7071), .A4(n7070), .ZN(n7079)
         );
  NOR2_X1 U8163 ( .A1(P1_D_REG_31__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .ZN(
        n7077) );
  NOR4_X1 U8164 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_29__SCAN_IN), .A4(P1_D_REG_28__SCAN_IN), .ZN(n7076) );
  NOR4_X1 U8165 ( .A1(P1_D_REG_23__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_21__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n7075) );
  NOR4_X1 U8166 ( .A1(P1_D_REG_27__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_25__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n7074) );
  AND4_X1 U8167 ( .A1(n7077), .A2(n7076), .A3(n7075), .A4(n7074), .ZN(n7078)
         );
  NAND2_X1 U8168 ( .A1(n7079), .A2(n7078), .ZN(n7404) );
  INV_X1 U8169 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n7250) );
  NOR2_X1 U8170 ( .A1(n7404), .A2(n7250), .ZN(n7081) );
  NAND2_X1 U8171 ( .A1(n7066), .A2(n5026), .ZN(n7402) );
  OAI21_X1 U8172 ( .B1(n7403), .B2(n7081), .A(n7402), .ZN(n7082) );
  INV_X1 U8173 ( .A(n7082), .ZN(n7373) );
  NAND3_X1 U8174 ( .A1(n7417), .A2(n7391), .A3(n7373), .ZN(n8014) );
  AOI21_X1 U8175 ( .B1(n10084), .B2(n7083), .A(n9977), .ZN(n7137) );
  NAND2_X1 U8176 ( .A1(n7380), .A2(n7629), .ZN(n7756) );
  NAND2_X1 U8177 ( .A1(n7491), .A2(n7766), .ZN(n7084) );
  NAND2_X1 U8178 ( .A1(n7756), .A2(n7084), .ZN(n7085) );
  NAND2_X1 U8179 ( .A1(n7086), .A2(n7085), .ZN(n7662) );
  NAND2_X1 U8180 ( .A1(n7087), .A2(n7662), .ZN(n7089) );
  NAND2_X1 U8181 ( .A1(n7763), .A2(n7676), .ZN(n7088) );
  NAND2_X1 U8182 ( .A1(n7089), .A2(n7088), .ZN(n7742) );
  NAND2_X1 U8183 ( .A1(n7742), .A2(n7743), .ZN(n7091) );
  NAND2_X1 U8184 ( .A1(n10403), .A2(n7633), .ZN(n7090) );
  NAND2_X1 U8185 ( .A1(n7091), .A2(n7090), .ZN(n10399) );
  NAND2_X1 U8186 ( .A1(n10399), .A2(n10406), .ZN(n7093) );
  NAND2_X1 U8187 ( .A1(n7794), .A2(n10423), .ZN(n7092) );
  NAND2_X1 U8188 ( .A1(n7093), .A2(n7092), .ZN(n7991) );
  INV_X1 U8189 ( .A(n7991), .ZN(n7095) );
  INV_X1 U8190 ( .A(n7993), .ZN(n7094) );
  NAND2_X1 U8191 ( .A1(n9791), .A2(n7997), .ZN(n7096) );
  NAND2_X1 U8192 ( .A1(n8011), .A2(n10502), .ZN(n7099) );
  NAND2_X1 U8193 ( .A1(n10479), .A2(n7099), .ZN(n8012) );
  NAND2_X1 U8194 ( .A1(n10490), .A2(n10518), .ZN(n7100) );
  NAND2_X1 U8195 ( .A1(n9790), .A2(n8109), .ZN(n7102) );
  INV_X1 U8196 ( .A(n8267), .ZN(n9789) );
  OR2_X1 U8197 ( .A1(n8276), .A2(n9789), .ZN(n7104) );
  NAND2_X1 U8198 ( .A1(n8189), .A2(n7104), .ZN(n8206) );
  NAND2_X1 U8199 ( .A1(n8206), .A2(n8207), .ZN(n8205) );
  INV_X1 U8200 ( .A(n8363), .ZN(n9788) );
  OR2_X1 U8201 ( .A1(n10168), .A2(n9788), .ZN(n7105) );
  AND2_X2 U8202 ( .A1(n8205), .A2(n7105), .ZN(n8297) );
  INV_X1 U8203 ( .A(n8486), .ZN(n9787) );
  NAND2_X1 U8204 ( .A1(n10163), .A2(n9787), .ZN(n7107) );
  INV_X1 U8205 ( .A(n8472), .ZN(n9404) );
  OR2_X1 U8206 ( .A1(n10157), .A2(n9404), .ZN(n7108) );
  NAND2_X1 U8207 ( .A1(n10152), .A2(n9786), .ZN(n7109) );
  OR2_X1 U8208 ( .A1(n10152), .A2(n9786), .ZN(n7110) );
  NAND2_X1 U8209 ( .A1(n7111), .A2(n7110), .ZN(n8517) );
  INV_X1 U8210 ( .A(n9465), .ZN(n8552) );
  NAND2_X1 U8211 ( .A1(n10146), .A2(n8552), .ZN(n7112) );
  INV_X1 U8212 ( .A(n9562), .ZN(n10053) );
  NAND2_X1 U8213 ( .A1(n10141), .A2(n10053), .ZN(n7113) );
  NAND2_X1 U8214 ( .A1(n8555), .A2(n7113), .ZN(n10049) );
  OR2_X1 U8215 ( .A1(n10135), .A2(n9573), .ZN(n7114) );
  NAND2_X1 U8216 ( .A1(n10049), .A2(n7114), .ZN(n7116) );
  NAND2_X1 U8217 ( .A1(n10135), .A2(n9573), .ZN(n7115) );
  NAND2_X1 U8218 ( .A1(n7116), .A2(n7115), .ZN(n10029) );
  NAND2_X1 U8219 ( .A1(n10029), .A2(n10032), .ZN(n7118) );
  INV_X1 U8220 ( .A(n9474), .ZN(n10052) );
  NAND2_X1 U8221 ( .A1(n10043), .A2(n10052), .ZN(n7117) );
  NAND2_X1 U8222 ( .A1(n7118), .A2(n7117), .ZN(n10012) );
  OR2_X1 U8223 ( .A1(n10123), .A2(n9572), .ZN(n7119) );
  INV_X1 U8224 ( .A(n10117), .ZN(n7120) );
  NAND2_X1 U8225 ( .A1(n9976), .A2(n9983), .ZN(n9975) );
  NAND2_X1 U8226 ( .A1(n10113), .A2(n9970), .ZN(n7121) );
  NAND2_X1 U8227 ( .A1(n9975), .A2(n7121), .ZN(n9960) );
  OR2_X1 U8228 ( .A1(n10106), .A2(n9955), .ZN(n7122) );
  NAND2_X1 U8229 ( .A1(n9960), .A2(n7122), .ZN(n7124) );
  NAND2_X1 U8230 ( .A1(n10106), .A2(n9955), .ZN(n7123) );
  INV_X1 U8231 ( .A(n9928), .ZN(n9935) );
  OR2_X1 U8232 ( .A1(n10102), .A2(n9969), .ZN(n9932) );
  AND2_X1 U8233 ( .A1(n9935), .A2(n9932), .ZN(n7125) );
  NAND2_X1 U8234 ( .A1(n10097), .A2(n9954), .ZN(n7126) );
  NAND2_X1 U8235 ( .A1(n9934), .A2(n7126), .ZN(n9915) );
  INV_X1 U8236 ( .A(n9915), .ZN(n7127) );
  OR2_X1 U8237 ( .A1(n10092), .A2(n9930), .ZN(n7128) );
  XNOR2_X1 U8238 ( .A(n8793), .B(n5366), .ZN(n10085) );
  INV_X1 U8239 ( .A(n7670), .ZN(n7413) );
  NAND2_X1 U8240 ( .A1(n7129), .A2(n8116), .ZN(n7667) );
  NOR2_X1 U8241 ( .A1(n7413), .A2(n8711), .ZN(n7131) );
  NAND2_X1 U8242 ( .A1(n10568), .A2(n7131), .ZN(n10028) );
  OR2_X1 U8243 ( .A1(n7627), .A2(n8166), .ZN(n7387) );
  INV_X1 U8244 ( .A(n7387), .ZN(n7132) );
  NOR2_X1 U8245 ( .A1(n10568), .A2(n7133), .ZN(n7134) );
  NAND2_X1 U8246 ( .A1(n7377), .A2(n7138), .ZN(n7139) );
  NAND2_X1 U8247 ( .A1(n7139), .A2(n7141), .ZN(n10256) );
  NAND2_X1 U8248 ( .A1(n10256), .A2(n5745), .ZN(n7140) );
  NAND2_X1 U8249 ( .A1(n7140), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  NAND2_X2 U8250 ( .A1(n7157), .A2(n10312), .ZN(n8945) );
  INV_X1 U8251 ( .A(n7141), .ZN(n7649) );
  NOR2_X1 U8252 ( .A1(n7377), .A2(n7649), .ZN(n7262) );
  INV_X1 U8253 ( .A(n7142), .ZN(n7143) );
  AOI211_X1 U8254 ( .C1(n7145), .C2(n7144), .A(n8927), .B(n7143), .ZN(n7151)
         );
  NOR2_X1 U8255 ( .A1(n8922), .A2(n7985), .ZN(n7150) );
  NOR2_X1 U8256 ( .A1(n8871), .A2(n10611), .ZN(n8911) );
  INV_X1 U8257 ( .A(n8911), .ZN(n8897) );
  INV_X1 U8258 ( .A(n8941), .ZN(n7772) );
  INV_X1 U8259 ( .A(n8910), .ZN(n8921) );
  INV_X1 U8260 ( .A(n7146), .ZN(n7984) );
  OAI22_X1 U8261 ( .A1(n8897), .A2(n7772), .B1(n8921), .B2(n7984), .ZN(n7149)
         );
  OAI22_X1 U8262 ( .A1(n8913), .A2(n8175), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7147), .ZN(n7148) );
  OR4_X1 U8263 ( .A1(n7151), .A2(n7150), .A3(n7149), .A4(n7148), .ZN(P2_U3215)
         );
  INV_X1 U8264 ( .A(n8950), .ZN(n7226) );
  XOR2_X1 U8265 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n8950), .Z(n8949) );
  INV_X1 U8266 ( .A(n10319), .ZN(n7228) );
  OR2_X1 U8267 ( .A1(n10319), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n7152) );
  NAND2_X1 U8268 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n10321) );
  NOR2_X1 U8269 ( .A1(n10322), .A2(n10321), .ZN(n10324) );
  INV_X1 U8270 ( .A(n10324), .ZN(n7153) );
  OAI21_X1 U8271 ( .B1(n7228), .B2(n7881), .A(n7153), .ZN(n8948) );
  NAND2_X1 U8272 ( .A1(n8949), .A2(n8948), .ZN(n8947) );
  OAI21_X1 U8273 ( .B1(n7154), .B2(n7226), .A(n8947), .ZN(n7477) );
  MUX2_X1 U8274 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n6266), .S(n7475), .Z(n7478)
         );
  INV_X1 U8275 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n7155) );
  MUX2_X1 U8276 ( .A(n7155), .B(P2_REG2_REG_4__SCAN_IN), .S(n7218), .Z(n7216)
         );
  AOI21_X1 U8277 ( .B1(n7218), .B2(P2_REG2_REG_4__SCAN_IN), .A(n7215), .ZN(
        n7163) );
  MUX2_X1 U8278 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n6290), .S(n7191), .Z(n7156)
         );
  INV_X1 U8279 ( .A(n7156), .ZN(n7162) );
  NOR2_X1 U8280 ( .A1(n7163), .A2(n7162), .ZN(n7186) );
  NAND2_X1 U8281 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7157), .ZN(n7158) );
  OAI211_X1 U8282 ( .C1(n7442), .C2(n7159), .A(n7158), .B(n8383), .ZN(n7174)
         );
  NAND2_X1 U8283 ( .A1(n7174), .A2(n7172), .ZN(n7160) );
  NAND2_X1 U8284 ( .A1(n7160), .A2(n8945), .ZN(n7164) );
  NOR2_X1 U8285 ( .A1(n6841), .A2(n9385), .ZN(n7161) );
  NAND2_X1 U8286 ( .A1(n7164), .A2(n7161), .ZN(n10325) );
  AOI211_X1 U8287 ( .C1(n7163), .C2(n7162), .A(n7186), .B(n10325), .ZN(n7185)
         );
  INV_X1 U8288 ( .A(n10320), .ZN(n8998) );
  INV_X1 U8289 ( .A(n7191), .ZN(n7232) );
  NOR2_X1 U8290 ( .A1(n8998), .A2(n7232), .ZN(n7184) );
  INV_X1 U8291 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n7168) );
  XOR2_X1 U8292 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n8950), .Z(n8953) );
  INV_X1 U8293 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n7167) );
  NAND2_X1 U8294 ( .A1(n10319), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n7165) );
  OAI21_X1 U8295 ( .B1(n10319), .B2(P2_REG1_REG_1__SCAN_IN), .A(n7165), .ZN(
        n10316) );
  INV_X1 U8296 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n7448) );
  INV_X1 U8297 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n7166) );
  OR3_X1 U8298 ( .A1(n10316), .A2(n7448), .A3(n7166), .ZN(n10318) );
  OAI21_X1 U8299 ( .B1(n7228), .B2(n7167), .A(n10318), .ZN(n8952) );
  NAND2_X1 U8300 ( .A1(n8953), .A2(n8952), .ZN(n8951) );
  OAI21_X1 U8301 ( .B1(n7168), .B2(n7226), .A(n8951), .ZN(n7470) );
  INV_X1 U8302 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10397) );
  MUX2_X1 U8303 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n10397), .S(n7475), .Z(n7471)
         );
  NAND2_X1 U8304 ( .A1(n7470), .A2(n7471), .ZN(n7469) );
  INV_X1 U8305 ( .A(n7469), .ZN(n7169) );
  AOI21_X1 U8306 ( .B1(P2_REG1_REG_3__SCAN_IN), .B2(n7475), .A(n7169), .ZN(
        n7221) );
  INV_X1 U8307 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n7170) );
  MUX2_X1 U8308 ( .A(n7170), .B(P2_REG1_REG_4__SCAN_IN), .S(n7218), .Z(n7220)
         );
  NOR2_X1 U8309 ( .A1(n7221), .A2(n7220), .ZN(n7219) );
  AOI21_X1 U8310 ( .B1(n7218), .B2(P2_REG1_REG_4__SCAN_IN), .A(n7219), .ZN(
        n7176) );
  INV_X1 U8311 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n7171) );
  MUX2_X1 U8312 ( .A(n7171), .B(P2_REG1_REG_5__SCAN_IN), .S(n7191), .Z(n7175)
         );
  NOR2_X1 U8313 ( .A1(n7176), .A2(n7175), .ZN(n7190) );
  AND2_X1 U8314 ( .A1(n7172), .A2(n9385), .ZN(n7173) );
  NAND2_X1 U8315 ( .A1(n7174), .A2(n7173), .ZN(n10329) );
  AOI211_X1 U8316 ( .C1(n7176), .C2(n7175), .A(n7190), .B(n10329), .ZN(n7183)
         );
  NAND2_X1 U8317 ( .A1(n7442), .A2(n8383), .ZN(n7178) );
  NAND2_X1 U8318 ( .A1(n7178), .A2(n7177), .ZN(n7179) );
  OAI21_X2 U8319 ( .B1(n7442), .B2(n7180), .A(n7179), .ZN(n10314) );
  INV_X1 U8320 ( .A(n10314), .ZN(n8126) );
  INV_X1 U8321 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n7181) );
  NAND2_X1 U8322 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3152), .ZN(n7771) );
  OAI21_X1 U8323 ( .B1(n8126), .B2(n7181), .A(n7771), .ZN(n7182) );
  OR4_X1 U8324 ( .A1(n7185), .A2(n7184), .A3(n7183), .A4(n7182), .ZN(P2_U3250)
         );
  INV_X1 U8325 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7187) );
  MUX2_X1 U8326 ( .A(n7187), .B(P2_REG2_REG_6__SCAN_IN), .S(n7205), .Z(n7188)
         );
  AOI211_X1 U8327 ( .C1(n7189), .C2(n7188), .A(n7200), .B(n10325), .ZN(n7199)
         );
  INV_X1 U8328 ( .A(n7205), .ZN(n7240) );
  NOR2_X1 U8329 ( .A1(n8998), .A2(n7240), .ZN(n7198) );
  AOI21_X1 U8330 ( .B1(n7191), .B2(P2_REG1_REG_5__SCAN_IN), .A(n7190), .ZN(
        n7194) );
  INV_X1 U8331 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n7192) );
  MUX2_X1 U8332 ( .A(n7192), .B(P2_REG1_REG_6__SCAN_IN), .S(n7205), .Z(n7193)
         );
  NOR2_X1 U8333 ( .A1(n7194), .A2(n7193), .ZN(n7204) );
  AOI211_X1 U8334 ( .C1(n7194), .C2(n7193), .A(n7204), .B(n10329), .ZN(n7197)
         );
  INV_X1 U8335 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n7195) );
  NAND2_X1 U8336 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(n4846), .ZN(n7822) );
  OAI21_X1 U8337 ( .B1(n8126), .B2(n7195), .A(n7822), .ZN(n7196) );
  OR4_X1 U8338 ( .A1(n7199), .A2(n7198), .A3(n7197), .A4(n7196), .ZN(P2_U3251)
         );
  MUX2_X1 U8339 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n7980), .S(n7524), .Z(n7201)
         );
  INV_X1 U8340 ( .A(n7201), .ZN(n7202) );
  AOI211_X1 U8341 ( .C1(n7203), .C2(n7202), .A(n7518), .B(n10325), .ZN(n7214)
         );
  INV_X1 U8342 ( .A(n7524), .ZN(n7245) );
  NOR2_X1 U8343 ( .A1(n8998), .A2(n7245), .ZN(n7213) );
  AOI21_X1 U8344 ( .B1(n7205), .B2(P2_REG1_REG_6__SCAN_IN), .A(n7204), .ZN(
        n7208) );
  INV_X1 U8345 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n7206) );
  MUX2_X1 U8346 ( .A(n7206), .B(P2_REG1_REG_7__SCAN_IN), .S(n7524), .Z(n7207)
         );
  NOR2_X1 U8347 ( .A1(n7208), .A2(n7207), .ZN(n7523) );
  AOI211_X1 U8348 ( .C1(n7208), .C2(n7207), .A(n7523), .B(n10329), .ZN(n7212)
         );
  INV_X1 U8349 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n7210) );
  NAND2_X1 U8350 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(n4846), .ZN(n7209) );
  OAI21_X1 U8351 ( .B1(n8126), .B2(n7210), .A(n7209), .ZN(n7211) );
  OR4_X1 U8352 ( .A1(n7214), .A2(n7213), .A3(n7212), .A4(n7211), .ZN(P2_U3252)
         );
  AOI211_X1 U8353 ( .C1(n7217), .C2(n7216), .A(n7215), .B(n10325), .ZN(n7225)
         );
  INV_X1 U8354 ( .A(n7218), .ZN(n7231) );
  NOR2_X1 U8355 ( .A1(n8998), .A2(n7231), .ZN(n7224) );
  AOI211_X1 U8356 ( .C1(n7221), .C2(n7220), .A(n7219), .B(n10329), .ZN(n7223)
         );
  INV_X1 U8357 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n8730) );
  NAND2_X1 U8358 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(n4846), .ZN(n7786) );
  OAI21_X1 U8359 ( .B1(n8126), .B2(n8730), .A(n7786), .ZN(n7222) );
  OR4_X1 U8360 ( .A1(n7225), .A2(n7224), .A3(n7223), .A4(n7222), .ZN(P2_U3249)
         );
  NOR2_X1 U8361 ( .A1(n5021), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9378) );
  INV_X1 U8362 ( .A(n9378), .ZN(n9387) );
  OAI222_X1 U8363 ( .A1(n4846), .A2(n7226), .B1(n8243), .B2(n7234), .C1(n5415), 
        .C2(n9387), .ZN(P2_U3356) );
  INV_X1 U8364 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n7227) );
  OAI222_X1 U8365 ( .A1(P2_U3152), .A2(n7228), .B1(n8243), .B2(n7237), .C1(
        n7227), .C2(n9387), .ZN(P2_U3357) );
  INV_X1 U8366 ( .A(n7475), .ZN(n7229) );
  OAI222_X1 U8367 ( .A1(n4846), .A2(n7229), .B1(n8243), .B2(n7235), .C1(n9387), 
        .C2(n5420), .ZN(P2_U3355) );
  NOR2_X1 U8368 ( .A1(n5021), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10204) );
  INV_X2 U8369 ( .A(n10204), .ZN(n8826) );
  NAND2_X1 U8370 ( .A1(n5021), .A2(P1_U3084), .ZN(n10209) );
  OAI222_X1 U8371 ( .A1(n7304), .A2(P1_U3084), .B1(n8826), .B2(n7230), .C1(
        n4986), .C2(n10209), .ZN(P1_U3349) );
  INV_X1 U8372 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n7366) );
  OAI222_X1 U8373 ( .A1(P2_U3152), .A2(n7231), .B1(n8243), .B2(n7230), .C1(
        n9387), .C2(n7366), .ZN(P2_U3354) );
  INV_X1 U8374 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n7233) );
  OAI222_X1 U8375 ( .A1(n9387), .A2(n7233), .B1(n8243), .B2(n7244), .C1(
        P2_U3152), .C2(n7232), .ZN(P2_U3353) );
  INV_X1 U8376 ( .A(n10209), .ZN(n8004) );
  INV_X1 U8377 ( .A(n8004), .ZN(n10196) );
  OAI222_X1 U8378 ( .A1(n10196), .A2(n5746), .B1(n8826), .B2(n7234), .C1(n7460), .C2(P1_U3084), .ZN(P1_U3351) );
  OAI222_X1 U8379 ( .A1(n10196), .A2(n7236), .B1(n8826), .B2(n7235), .C1(n7300), .C2(P1_U3084), .ZN(P1_U3350) );
  OAI222_X1 U8380 ( .A1(n10196), .A2(n7238), .B1(n8826), .B2(n7237), .C1(n7323), .C2(P1_U3084), .ZN(P1_U3352) );
  INV_X1 U8381 ( .A(n7239), .ZN(n7242) );
  INV_X1 U8382 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n7370) );
  OAI222_X1 U8383 ( .A1(n4846), .A2(n7240), .B1(n8243), .B2(n7242), .C1(n9387), 
        .C2(n7370), .ZN(P2_U3352) );
  OAI222_X1 U8384 ( .A1(n7338), .A2(P1_U3084), .B1(n8826), .B2(n7242), .C1(
        n7241), .C2(n10196), .ZN(P1_U3347) );
  OAI222_X1 U8385 ( .A1(n7307), .A2(P1_U3084), .B1(n8826), .B2(n7244), .C1(
        n7243), .C2(n10196), .ZN(P1_U3348) );
  INV_X1 U8386 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n7372) );
  OAI222_X1 U8387 ( .A1(P2_U3152), .A2(n7245), .B1(n8243), .B2(n7247), .C1(
        n9387), .C2(n7372), .ZN(P2_U3351) );
  OAI222_X1 U8388 ( .A1(n7359), .A2(P1_U3084), .B1(n8826), .B2(n7247), .C1(
        n7246), .C2(n10209), .ZN(P1_U3346) );
  NOR2_X1 U8389 ( .A1(n10314), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U8390 ( .A(n7388), .ZN(n7249) );
  INV_X1 U8391 ( .A(n7402), .ZN(n7248) );
  AOI22_X1 U8392 ( .A1(n10211), .A2(n7250), .B1(n7249), .B2(n7248), .ZN(
        P1_U3441) );
  INV_X1 U8393 ( .A(n7341), .ZN(n7585) );
  INV_X1 U8394 ( .A(n7251), .ZN(n7253) );
  OAI222_X1 U8395 ( .A1(n7585), .A2(P1_U3084), .B1(n8826), .B2(n7253), .C1(
        n10196), .C2(n5435), .ZN(P1_U3345) );
  INV_X1 U8396 ( .A(n7545), .ZN(n7252) );
  OAI222_X1 U8397 ( .A1(n9387), .A2(n7254), .B1(n8243), .B2(n7253), .C1(n4846), 
        .C2(n7252), .ZN(P2_U3350) );
  INV_X1 U8398 ( .A(n7255), .ZN(n7257) );
  AOI22_X1 U8399 ( .A1(n10281), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n8004), .ZN(n7256) );
  OAI21_X1 U8400 ( .B1(n7257), .B2(n8826), .A(n7256), .ZN(P1_U3344) );
  INV_X1 U8401 ( .A(n7613), .ZN(n7619) );
  OAI222_X1 U8402 ( .A1(n9387), .A2(n7258), .B1(n8243), .B2(n7257), .C1(n7619), 
        .C2(P2_U3152), .ZN(P2_U3349) );
  NAND2_X1 U8403 ( .A1(n8552), .A2(P1_U4006), .ZN(n7259) );
  OAI21_X1 U8404 ( .B1(P1_U4006), .B2(n5467), .A(n7259), .ZN(P1_U3570) );
  INV_X1 U8405 ( .A(n7260), .ZN(n7316) );
  AOI22_X1 U8406 ( .A1(n8963), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n9378), .ZN(n7261) );
  OAI21_X1 U8407 ( .B1(n7316), .B2(n8243), .A(n7261), .ZN(P2_U3347) );
  INV_X1 U8408 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n7287) );
  OR2_X1 U8409 ( .A1(n10260), .A2(P1_U3084), .ZN(n10206) );
  INV_X1 U8410 ( .A(n10206), .ZN(n7263) );
  NAND2_X1 U8411 ( .A1(n10256), .A2(n7263), .ZN(n7588) );
  INV_X1 U8412 ( .A(n7588), .ZN(n7264) );
  AND2_X1 U8413 ( .A1(n7264), .A2(n6205), .ZN(n10339) );
  INV_X1 U8414 ( .A(n7300), .ZN(n7296) );
  AND2_X1 U8415 ( .A1(P1_U3084), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n7656) );
  OR2_X1 U8416 ( .A1(n6205), .A2(P1_U3084), .ZN(n10201) );
  INV_X1 U8417 ( .A(n10260), .ZN(n7265) );
  NOR2_X1 U8418 ( .A1(n10201), .A2(n7265), .ZN(n7266) );
  INV_X1 U8419 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10373) );
  MUX2_X1 U8420 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n10373), .S(n7460), .Z(n7456)
         );
  INV_X1 U8421 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n7267) );
  MUX2_X1 U8422 ( .A(n7267), .B(P1_REG1_REG_1__SCAN_IN), .S(n7323), .Z(n7269)
         );
  AND2_X1 U8423 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n7268) );
  NAND2_X1 U8424 ( .A1(n7269), .A2(n7268), .ZN(n7319) );
  OR2_X1 U8425 ( .A1(n7323), .A2(n7267), .ZN(n7270) );
  AND2_X1 U8426 ( .A1(n7319), .A2(n7270), .ZN(n7457) );
  NOR2_X1 U8427 ( .A1(n7456), .A2(n7457), .ZN(n7455) );
  INV_X1 U8428 ( .A(n7455), .ZN(n7273) );
  NAND2_X1 U8429 ( .A1(n5172), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n7272) );
  INV_X1 U8430 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n10388) );
  MUX2_X1 U8431 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n10388), .S(n7300), .Z(n7271)
         );
  AOI21_X1 U8432 ( .B1(n7273), .B2(n7272), .A(n7271), .ZN(n7295) );
  AND3_X1 U8433 ( .A1(n7273), .A2(n7272), .A3(n7271), .ZN(n7274) );
  NOR3_X1 U8434 ( .A1(n10299), .A2(n7295), .A3(n7274), .ZN(n7275) );
  AOI211_X1 U8435 ( .C1(n10339), .C2(n7296), .A(n7656), .B(n7275), .ZN(n7286)
         );
  INV_X1 U8436 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n7674) );
  MUX2_X1 U8437 ( .A(n7674), .B(P1_REG2_REG_2__SCAN_IN), .S(n7460), .Z(n7279)
         );
  INV_X1 U8438 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n7276) );
  MUX2_X1 U8439 ( .A(n7276), .B(P1_REG2_REG_1__SCAN_IN), .S(n7323), .Z(n7277)
         );
  AND2_X1 U8440 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n7322) );
  NAND2_X1 U8441 ( .A1(n7277), .A2(n7322), .ZN(n7324) );
  OR2_X1 U8442 ( .A1(n7323), .A2(n7276), .ZN(n7278) );
  NAND2_X1 U8443 ( .A1(n7324), .A2(n7278), .ZN(n7451) );
  AND2_X1 U8444 ( .A1(n7279), .A2(n7451), .ZN(n7452) );
  NOR2_X1 U8445 ( .A1(n7460), .A2(n7674), .ZN(n7283) );
  INV_X1 U8446 ( .A(n7283), .ZN(n7281) );
  INV_X1 U8447 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n7748) );
  MUX2_X1 U8448 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n7748), .S(n7300), .Z(n7280)
         );
  NAND2_X1 U8449 ( .A1(n7281), .A2(n7280), .ZN(n7284) );
  OR2_X1 U8450 ( .A1(n7588), .A2(n6205), .ZN(n10269) );
  INV_X1 U8451 ( .A(n10269), .ZN(n10335) );
  MUX2_X1 U8452 ( .A(n7748), .B(P1_REG2_REG_3__SCAN_IN), .S(n7300), .Z(n7282)
         );
  OAI21_X1 U8453 ( .B1(n7452), .B2(n7283), .A(n7282), .ZN(n7302) );
  OAI211_X1 U8454 ( .C1(n7452), .C2(n7284), .A(n10335), .B(n7302), .ZN(n7285)
         );
  OAI211_X1 U8455 ( .C1(n10342), .C2(n7287), .A(n7286), .B(n7285), .ZN(
        P1_U3244) );
  NAND2_X1 U8456 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(n8945), .ZN(n7288) );
  OAI21_X1 U8457 ( .B1(n9067), .B2(n8945), .A(n7288), .ZN(P2_U3582) );
  NAND2_X1 U8458 ( .A1(P2_DATAO_REG_19__SCAN_IN), .A2(n8945), .ZN(n7289) );
  OAI21_X1 U8459 ( .B1(n9248), .B2(n8945), .A(n7289), .ZN(P2_U3571) );
  INV_X1 U8460 ( .A(n7290), .ZN(n7292) );
  OAI222_X1 U8461 ( .A1(P1_U3084), .A2(n7579), .B1(n8826), .B2(n7292), .C1(
        n7291), .C2(n10209), .ZN(P1_U3343) );
  INV_X1 U8462 ( .A(n7940), .ZN(n7932) );
  OAI222_X1 U8463 ( .A1(n9387), .A2(n7293), .B1(n8243), .B2(n7292), .C1(n7932), 
        .C2(n4846), .ZN(P2_U3348) );
  NAND2_X1 U8464 ( .A1(n8135), .A2(P2_U3966), .ZN(n7294) );
  OAI21_X1 U8465 ( .B1(n5435), .B2(P2_U3966), .A(n7294), .ZN(P2_U3560) );
  INV_X1 U8466 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n7314) );
  INV_X1 U8467 ( .A(n7307), .ZN(n7337) );
  AND2_X1 U8468 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n7809) );
  INV_X1 U8469 ( .A(n7304), .ZN(n10338) );
  AOI21_X1 U8470 ( .B1(P1_REG1_REG_3__SCAN_IN), .B2(n7296), .A(n7295), .ZN(
        n10346) );
  INV_X1 U8471 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n10415) );
  MUX2_X1 U8472 ( .A(n10415), .B(P1_REG1_REG_4__SCAN_IN), .S(n7304), .Z(n10347) );
  NAND2_X1 U8473 ( .A1(n10346), .A2(n10347), .ZN(n10345) );
  OAI21_X1 U8474 ( .B1(n10338), .B2(P1_REG1_REG_4__SCAN_IN), .A(n10345), .ZN(
        n7298) );
  INV_X1 U8475 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n10469) );
  MUX2_X1 U8476 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n10469), .S(n7307), .Z(n7297)
         );
  NOR2_X1 U8477 ( .A1(n7298), .A2(n7297), .ZN(n7330) );
  AOI211_X1 U8478 ( .C1(n7298), .C2(n7297), .A(n7330), .B(n10299), .ZN(n7299)
         );
  AOI211_X1 U8479 ( .C1(n10339), .C2(n7337), .A(n7809), .B(n7299), .ZN(n7313)
         );
  OR2_X1 U8480 ( .A1(n7300), .A2(n7748), .ZN(n7301) );
  AND2_X1 U8481 ( .A1(n7302), .A2(n7301), .ZN(n10334) );
  INV_X1 U8482 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n7303) );
  OR2_X1 U8483 ( .A1(n7304), .A2(n7303), .ZN(n7305) );
  NAND2_X1 U8484 ( .A1(n7304), .A2(n7303), .ZN(n7306) );
  AND2_X1 U8485 ( .A1(n7305), .A2(n7306), .ZN(n10333) );
  AND2_X1 U8486 ( .A1(n10334), .A2(n10333), .ZN(n10337) );
  INV_X1 U8487 ( .A(n7306), .ZN(n7308) );
  INV_X1 U8488 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n7992) );
  MUX2_X1 U8489 ( .A(n7992), .B(P1_REG2_REG_5__SCAN_IN), .S(n7307), .Z(n7309)
         );
  OAI21_X1 U8490 ( .B1(n10337), .B2(n7308), .A(n7309), .ZN(n7336) );
  INV_X1 U8491 ( .A(n7336), .ZN(n7311) );
  NOR3_X1 U8492 ( .A1(n10337), .A2(n7309), .A3(n7308), .ZN(n7310) );
  OAI21_X1 U8493 ( .B1(n7311), .B2(n7310), .A(n10335), .ZN(n7312) );
  OAI211_X1 U8494 ( .C1(n10342), .C2(n7314), .A(n7313), .B(n7312), .ZN(
        P1_U3246) );
  INV_X1 U8495 ( .A(n7711), .ZN(n7594) );
  INV_X1 U8496 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n7315) );
  OAI222_X1 U8497 ( .A1(P1_U3084), .A2(n7594), .B1(n8826), .B2(n7316), .C1(
        n7315), .C2(n10196), .ZN(P1_U3342) );
  INV_X1 U8498 ( .A(n10342), .ZN(n10294) );
  INV_X1 U8499 ( .A(n10339), .ZN(n9836) );
  NAND2_X1 U8500 ( .A1(P1_REG3_REG_1__SCAN_IN), .A2(P1_U3084), .ZN(n7321) );
  INV_X1 U8501 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n10261) );
  INV_X1 U8502 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n10255) );
  MUX2_X1 U8503 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n7267), .S(n7323), .Z(n7317)
         );
  OAI21_X1 U8504 ( .B1(n10261), .B2(n10255), .A(n7317), .ZN(n7318) );
  NAND3_X1 U8505 ( .A1(n10349), .A2(n7319), .A3(n7318), .ZN(n7320) );
  OAI211_X1 U8506 ( .C1(n9836), .C2(n7323), .A(n7321), .B(n7320), .ZN(n7328)
         );
  INV_X1 U8507 ( .A(n7322), .ZN(n7464) );
  MUX2_X1 U8508 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n7276), .S(n7323), .Z(n7326)
         );
  INV_X1 U8509 ( .A(n7324), .ZN(n7325) );
  AOI211_X1 U8510 ( .C1(n7464), .C2(n7326), .A(n7325), .B(n10269), .ZN(n7327)
         );
  AOI211_X1 U8511 ( .C1(n10294), .C2(P1_ADDR_REG_1__SCAN_IN), .A(n7328), .B(
        n7327), .ZN(n7329) );
  INV_X1 U8512 ( .A(n7329), .ZN(P1_U3242) );
  INV_X1 U8513 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n7331) );
  INV_X1 U8514 ( .A(n7338), .ZN(n10267) );
  AOI21_X1 U8515 ( .B1(P1_REG1_REG_5__SCAN_IN), .B2(n7337), .A(n7330), .ZN(
        n10275) );
  INV_X1 U8516 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n10496) );
  MUX2_X1 U8517 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n10496), .S(n7338), .Z(n10274) );
  NOR2_X1 U8518 ( .A1(n10275), .A2(n10274), .ZN(n10273) );
  AOI21_X1 U8519 ( .B1(P1_REG1_REG_6__SCAN_IN), .B2(n10267), .A(n10273), .ZN(
        n7356) );
  MUX2_X1 U8520 ( .A(n7331), .B(P1_REG1_REG_7__SCAN_IN), .S(n7359), .Z(n7355)
         );
  AND2_X1 U8521 ( .A1(n7356), .A2(n7355), .ZN(n7357) );
  AOI21_X1 U8522 ( .B1(n7331), .B2(n7359), .A(n7357), .ZN(n7333) );
  INV_X1 U8523 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10553) );
  AOI22_X1 U8524 ( .A1(P1_REG1_REG_8__SCAN_IN), .A2(n7585), .B1(n7341), .B2(
        n10553), .ZN(n7332) );
  NOR2_X1 U8525 ( .A1(n7333), .A2(n7332), .ZN(n7572) );
  AOI21_X1 U8526 ( .B1(n7333), .B2(n7332), .A(n7572), .ZN(n7348) );
  NOR2_X1 U8527 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7334), .ZN(n8104) );
  NOR2_X1 U8528 ( .A1(n9836), .A2(n7585), .ZN(n7335) );
  AOI211_X1 U8529 ( .C1(n10294), .C2(P1_ADDR_REG_8__SCAN_IN), .A(n8104), .B(
        n7335), .ZN(n7347) );
  OAI21_X1 U8530 ( .B1(n7337), .B2(P1_REG2_REG_5__SCAN_IN), .A(n7336), .ZN(
        n10270) );
  INV_X1 U8531 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n7339) );
  MUX2_X1 U8532 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n7339), .S(n7338), .Z(n10271)
         );
  NOR2_X1 U8533 ( .A1(n10270), .A2(n10271), .ZN(n10268) );
  AOI21_X1 U8534 ( .B1(P1_REG2_REG_6__SCAN_IN), .B2(n10267), .A(n10268), .ZN(
        n7349) );
  INV_X1 U8535 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n7340) );
  MUX2_X1 U8536 ( .A(n7340), .B(P1_REG2_REG_7__SCAN_IN), .S(n7359), .Z(n7350)
         );
  NAND2_X1 U8537 ( .A1(n7349), .A2(n7350), .ZN(n7351) );
  NAND2_X1 U8538 ( .A1(n7359), .A2(n7340), .ZN(n7343) );
  INV_X1 U8539 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n7342) );
  MUX2_X1 U8540 ( .A(n7342), .B(P1_REG2_REG_8__SCAN_IN), .S(n7341), .Z(n7344)
         );
  AOI21_X1 U8541 ( .B1(n7351), .B2(n7343), .A(n7344), .ZN(n7584) );
  AND3_X1 U8542 ( .A1(n7351), .A2(n7344), .A3(n7343), .ZN(n7345) );
  OAI21_X1 U8543 ( .B1(n7584), .B2(n7345), .A(n10335), .ZN(n7346) );
  OAI211_X1 U8544 ( .C1(n7348), .C2(n10299), .A(n7347), .B(n7346), .ZN(
        P1_U3249) );
  INV_X1 U8545 ( .A(n7349), .ZN(n7354) );
  INV_X1 U8546 ( .A(n7350), .ZN(n7353) );
  INV_X1 U8547 ( .A(n7351), .ZN(n7352) );
  AOI21_X1 U8548 ( .B1(n7354), .B2(n7353), .A(n7352), .ZN(n7363) );
  NOR2_X1 U8549 ( .A1(n7356), .A2(n7355), .ZN(n7358) );
  OAI21_X1 U8550 ( .B1(n7358), .B2(n7357), .A(n10349), .ZN(n7362) );
  AND2_X1 U8551 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n7910) );
  NOR2_X1 U8552 ( .A1(n9836), .A2(n7359), .ZN(n7360) );
  AOI211_X1 U8553 ( .C1(n10294), .C2(P1_ADDR_REG_7__SCAN_IN), .A(n7910), .B(
        n7360), .ZN(n7361) );
  OAI211_X1 U8554 ( .C1(n7363), .C2(n10269), .A(n7362), .B(n7361), .ZN(
        P1_U3248) );
  NAND2_X1 U8555 ( .A1(n7364), .A2(P1_U4006), .ZN(n7365) );
  OAI21_X1 U8556 ( .B1(P1_U4006), .B2(n7366), .A(n7365), .ZN(P1_U3559) );
  NAND2_X1 U8557 ( .A1(n9404), .A2(P1_U4006), .ZN(n7367) );
  OAI21_X1 U8558 ( .B1(P1_U4006), .B2(n5457), .A(n7367), .ZN(P1_U3568) );
  NAND2_X1 U8559 ( .A1(n5777), .A2(P1_U4006), .ZN(n7368) );
  OAI21_X1 U8560 ( .B1(P1_U4006), .B2(n5420), .A(n7368), .ZN(P1_U3558) );
  NAND2_X1 U8561 ( .A1(n7994), .A2(P1_U4006), .ZN(n7369) );
  OAI21_X1 U8562 ( .B1(P1_U4006), .B2(n7370), .A(n7369), .ZN(P1_U3561) );
  NAND2_X1 U8563 ( .A1(n10541), .A2(P1_U4006), .ZN(n7371) );
  OAI21_X1 U8564 ( .B1(P1_U4006), .B2(n7372), .A(n7371), .ZN(P1_U3562) );
  NAND2_X1 U8565 ( .A1(n7373), .A2(n7411), .ZN(n7390) );
  OR2_X1 U8566 ( .A1(n7514), .A2(n7387), .ZN(n7374) );
  OAI21_X1 U8567 ( .B1(n10255), .B2(n7377), .A(n7378), .ZN(n7379) );
  INV_X4 U8568 ( .A(n8701), .ZN(n8721) );
  NAND2_X1 U8569 ( .A1(n7380), .A2(n8721), .ZN(n7383) );
  INV_X1 U8570 ( .A(n7377), .ZN(n7381) );
  AOI22_X1 U8571 ( .A1(n7629), .A2(n8718), .B1(n7381), .B2(
        P1_REG1_REG_0__SCAN_IN), .ZN(n7382) );
  NAND2_X1 U8572 ( .A1(n7384), .A2(n7495), .ZN(n7499) );
  OAI21_X1 U8573 ( .B1(n7384), .B2(n7495), .A(n7499), .ZN(n7463) );
  INV_X1 U8574 ( .A(n7627), .ZN(n7412) );
  OR2_X1 U8575 ( .A1(n10365), .A2(n7385), .ZN(n7386) );
  NAND2_X1 U8576 ( .A1(n7463), .A2(n9536), .ZN(n7395) );
  NOR2_X1 U8577 ( .A1(n7388), .A2(n7387), .ZN(n7389) );
  AND2_X1 U8578 ( .A1(n7390), .A2(n7389), .ZN(n7654) );
  INV_X1 U8579 ( .A(n7654), .ZN(n7392) );
  NAND2_X1 U8580 ( .A1(n7390), .A2(n10581), .ZN(n7652) );
  NAND3_X1 U8581 ( .A1(n7392), .A2(n7391), .A3(n7652), .ZN(n9523) );
  NAND2_X1 U8582 ( .A1(n6205), .A2(n7413), .ZN(n7393) );
  AOI22_X1 U8583 ( .A1(n9523), .A2(P1_REG3_REG_0__SCAN_IN), .B1(n9545), .B2(
        n7491), .ZN(n7394) );
  OAI211_X1 U8584 ( .C1(n9548), .C2(n7759), .A(n7395), .B(n7394), .ZN(P1_U3230) );
  INV_X1 U8585 ( .A(n7396), .ZN(n7401) );
  NOR2_X1 U8586 ( .A1(n8927), .A2(n7701), .ZN(n8875) );
  AOI22_X1 U8587 ( .A1(n8875), .A2(n6847), .B1(n7565), .B2(n8905), .ZN(n7400)
         );
  OR2_X1 U8588 ( .A1(n7397), .A2(P2_U3152), .ZN(n7557) );
  OAI22_X1 U8589 ( .A1(n8922), .A2(n7852), .B1(n8913), .B2(n7687), .ZN(n7398)
         );
  AOI21_X1 U8590 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(n7557), .A(n7398), .ZN(
        n7399) );
  OAI21_X1 U8591 ( .B1(n7401), .B2(n7400), .A(n7399), .ZN(P2_U3234) );
  OAI21_X1 U8592 ( .B1(n7403), .B2(P1_D_REG_1__SCAN_IN), .A(n7402), .ZN(n7408)
         );
  NAND2_X1 U8593 ( .A1(n7405), .A2(n7404), .ZN(n7407) );
  NAND3_X1 U8594 ( .A1(n7408), .A2(n7407), .A3(n7406), .ZN(n7410) );
  NOR2_X1 U8595 ( .A1(n7413), .A2(n7412), .ZN(n7414) );
  AOI22_X1 U8596 ( .A1(n7415), .A2(n7414), .B1(n10539), .B2(n7491), .ZN(n7632)
         );
  OAI21_X1 U8597 ( .B1(n7759), .B2(n7627), .A(n7632), .ZN(n7419) );
  NAND2_X1 U8598 ( .A1(n7419), .A2(n10590), .ZN(n7416) );
  OAI21_X1 U8599 ( .B1(n10590), .B2(n10261), .A(n7416), .ZN(P1_U3523) );
  INV_X1 U8600 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n7421) );
  NAND2_X1 U8601 ( .A1(n7419), .A2(n10594), .ZN(n7420) );
  OAI21_X1 U8602 ( .B1(n10594), .B2(n7421), .A(n7420), .ZN(P1_U3454) );
  INV_X1 U8603 ( .A(n7422), .ZN(n7449) );
  AOI22_X1 U8604 ( .A1(n7836), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n8004), .ZN(n7423) );
  OAI21_X1 U8605 ( .B1(n7449), .B2(n8826), .A(n7423), .ZN(P1_U3341) );
  INV_X1 U8606 ( .A(n7439), .ZN(n7424) );
  NOR3_X1 U8607 ( .A1(n7442), .A2(n7425), .A3(n7424), .ZN(n7426) );
  AND2_X1 U8608 ( .A1(n7441), .A2(n7440), .ZN(n7428) );
  INV_X1 U8609 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n7438) );
  INV_X1 U8610 ( .A(n7429), .ZN(n7430) );
  OR2_X1 U8611 ( .A1(n7857), .A2(n10436), .ZN(n7433) );
  NAND2_X1 U8612 ( .A1(n8946), .A2(n9178), .ZN(n7432) );
  NAND2_X1 U8613 ( .A1(n7433), .A2(n7432), .ZN(n7854) );
  INV_X1 U8614 ( .A(n10622), .ZN(n7434) );
  NAND2_X1 U8615 ( .A1(n10619), .A2(n7434), .ZN(n10677) );
  OAI22_X1 U8616 ( .A1(n7857), .A2(n10667), .B1(n7435), .B2(n7852), .ZN(n7436)
         );
  OR2_X1 U8617 ( .A1(n7854), .A2(n7436), .ZN(n7446) );
  NAND2_X1 U8618 ( .A1(n7446), .A2(n10684), .ZN(n7437) );
  OAI21_X1 U8619 ( .B1(n10684), .B2(n7438), .A(n7437), .ZN(P2_U3451) );
  NAND3_X1 U8620 ( .A1(n7441), .A2(n7440), .A3(n7439), .ZN(n7443) );
  NOR2_X1 U8621 ( .A1(n7443), .A2(n7442), .ZN(n7444) );
  NAND2_X1 U8622 ( .A1(n7446), .A2(n10681), .ZN(n7447) );
  OAI21_X1 U8623 ( .B1(n10681), .B2(n7448), .A(n7447), .ZN(P2_U3520) );
  INV_X1 U8624 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n7450) );
  INV_X1 U8625 ( .A(n8026), .ZN(n8022) );
  OAI222_X1 U8626 ( .A1(n9387), .A2(n7450), .B1(n8243), .B2(n7449), .C1(
        P2_U3152), .C2(n8022), .ZN(P2_U3346) );
  INV_X1 U8627 ( .A(n7451), .ZN(n7454) );
  MUX2_X1 U8628 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n7674), .S(n7460), .Z(n7453)
         );
  AOI211_X1 U8629 ( .C1(n7454), .C2(n7453), .A(n7452), .B(n10269), .ZN(n7462)
         );
  AOI211_X1 U8630 ( .C1(n7457), .C2(n7456), .A(n7455), .B(n10299), .ZN(n7458)
         );
  AOI21_X1 U8631 ( .B1(P1_REG3_REG_2__SCAN_IN), .B2(P1_U3084), .A(n7458), .ZN(
        n7459) );
  OAI21_X1 U8632 ( .B1(n7460), .B2(n9836), .A(n7459), .ZN(n7461) );
  AOI211_X1 U8633 ( .C1(n10294), .C2(P1_ADDR_REG_2__SCAN_IN), .A(n7462), .B(
        n7461), .ZN(n7468) );
  MUX2_X1 U8634 ( .A(n7464), .B(n7463), .S(n10260), .Z(n7467) );
  OAI21_X1 U8635 ( .B1(P1_REG2_REG_0__SCAN_IN), .B2(n10260), .A(n7465), .ZN(
        n10259) );
  NAND2_X1 U8636 ( .A1(n10259), .A2(n10255), .ZN(n7466) );
  OAI211_X1 U8637 ( .C1(n7467), .C2(n6205), .A(P1_U4006), .B(n7466), .ZN(
        n10351) );
  NAND2_X1 U8638 ( .A1(n7468), .A2(n10351), .ZN(P1_U3243) );
  INV_X1 U8639 ( .A(n10329), .ZN(n8993) );
  OAI211_X1 U8640 ( .C1(n7471), .C2(n7470), .A(n8993), .B(n7469), .ZN(n7473)
         );
  NAND2_X1 U8641 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_U3152), .ZN(n7472) );
  OAI211_X1 U8642 ( .C1(n8126), .C2(n8731), .A(n7473), .B(n7472), .ZN(n7474)
         );
  AOI21_X1 U8643 ( .B1(n7475), .B2(n10320), .A(n7474), .ZN(n7480) );
  INV_X1 U8644 ( .A(n10325), .ZN(n8976) );
  OAI211_X1 U8645 ( .C1(n7478), .C2(n7477), .A(n8976), .B(n7476), .ZN(n7479)
         );
  NAND2_X1 U8646 ( .A1(n7480), .A2(n7479), .ZN(P2_U3248) );
  INV_X1 U8647 ( .A(n7557), .ZN(n7490) );
  INV_X1 U8648 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n9747) );
  OAI21_X1 U8649 ( .B1(n7483), .B2(n7482), .A(n7481), .ZN(n7484) );
  NAND2_X1 U8650 ( .A1(n7484), .A2(n8905), .ZN(n7489) );
  NOR2_X1 U8651 ( .A1(n6860), .A2(n10613), .ZN(n7487) );
  NOR2_X1 U8652 ( .A1(n7485), .A2(n10611), .ZN(n7486) );
  OR2_X1 U8653 ( .A1(n7487), .A2(n7486), .ZN(n7563) );
  INV_X1 U8654 ( .A(n8871), .ZN(n8925) );
  AOI22_X1 U8655 ( .A1(n8915), .A2(n7885), .B1(n7563), .B2(n8925), .ZN(n7488)
         );
  OAI211_X1 U8656 ( .C1(n7490), .C2(n9747), .A(n7489), .B(n7488), .ZN(P2_U3224) );
  NAND2_X1 U8657 ( .A1(n7491), .A2(n8721), .ZN(n7493) );
  NAND2_X1 U8658 ( .A1(n7766), .A2(n8718), .ZN(n7492) );
  NAND2_X1 U8659 ( .A1(n7493), .A2(n7492), .ZN(n7494) );
  INV_X1 U8660 ( .A(n7495), .ZN(n7497) );
  XNOR2_X1 U8661 ( .A(n7506), .B(n7505), .ZN(n7503) );
  NAND2_X1 U8662 ( .A1(n7491), .A2(n8720), .ZN(n7501) );
  NAND2_X1 U8663 ( .A1(n7766), .A2(n8721), .ZN(n7500) );
  NAND2_X1 U8664 ( .A1(n7501), .A2(n7500), .ZN(n7509) );
  INV_X1 U8665 ( .A(n7509), .ZN(n7502) );
  NAND2_X1 U8666 ( .A1(n7503), .A2(n7502), .ZN(n7511) );
  NAND2_X1 U8667 ( .A1(n7505), .A2(n7506), .ZN(n7504) );
  NAND2_X1 U8668 ( .A1(n7504), .A2(n7509), .ZN(n7638) );
  NAND2_X1 U8669 ( .A1(n7508), .A2(n7507), .ZN(n7637) );
  INV_X1 U8670 ( .A(n7637), .ZN(n7510) );
  AOI22_X1 U8671 ( .A1(n7511), .A2(n7638), .B1(n7510), .B2(n7509), .ZN(n7517)
         );
  OR2_X1 U8672 ( .A1(n6205), .A2(n7670), .ZN(n7513) );
  AOI22_X1 U8673 ( .A1(n5029), .A2(n9545), .B1(n9558), .B2(n7380), .ZN(n7516)
         );
  AOI22_X1 U8674 ( .A1(n9523), .A2(P1_REG3_REG_1__SCAN_IN), .B1(n9564), .B2(
        n7766), .ZN(n7515) );
  OAI211_X1 U8675 ( .C1(n7517), .C2(n9566), .A(n7516), .B(n7515), .ZN(P1_U3220) );
  AOI21_X1 U8676 ( .B1(n7524), .B2(P2_REG2_REG_7__SCAN_IN), .A(n7518), .ZN(
        n7542) );
  NAND2_X1 U8677 ( .A1(n7545), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n7519) );
  OAI21_X1 U8678 ( .B1(n7545), .B2(P2_REG2_REG_8__SCAN_IN), .A(n7519), .ZN(
        n7541) );
  NOR2_X1 U8679 ( .A1(n7542), .A2(n7541), .ZN(n7540) );
  AOI21_X1 U8680 ( .B1(n7545), .B2(P2_REG2_REG_8__SCAN_IN), .A(n7540), .ZN(
        n7522) );
  MUX2_X1 U8681 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n6348), .S(n7613), .Z(n7520)
         );
  INV_X1 U8682 ( .A(n7520), .ZN(n7521) );
  NOR2_X1 U8683 ( .A1(n7522), .A2(n7521), .ZN(n7612) );
  AOI211_X1 U8684 ( .C1(n7522), .C2(n7521), .A(n7612), .B(n10325), .ZN(n7533)
         );
  NOR2_X1 U8685 ( .A1(n9669), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8172) );
  AOI21_X1 U8686 ( .B1(n10314), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n8172), .ZN(
        n7531) );
  AOI21_X1 U8687 ( .B1(n7524), .B2(P2_REG1_REG_7__SCAN_IN), .A(n7523), .ZN(
        n7535) );
  NAND2_X1 U8688 ( .A1(n7545), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n7534) );
  NAND2_X1 U8689 ( .A1(n7535), .A2(n7534), .ZN(n7526) );
  OR2_X1 U8690 ( .A1(n7545), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n7525) );
  AND2_X1 U8691 ( .A1(n7526), .A2(n7525), .ZN(n7529) );
  INV_X1 U8692 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n7527) );
  MUX2_X1 U8693 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n7527), .S(n7613), .Z(n7528)
         );
  NAND2_X1 U8694 ( .A1(n7529), .A2(n7528), .ZN(n7618) );
  OAI211_X1 U8695 ( .C1(n7529), .C2(n7528), .A(n8993), .B(n7618), .ZN(n7530)
         );
  OAI211_X1 U8696 ( .C1(n8998), .C2(n7619), .A(n7531), .B(n7530), .ZN(n7532)
         );
  OR2_X1 U8697 ( .A1(n7533), .A2(n7532), .ZN(P2_U3254) );
  OAI21_X1 U8698 ( .B1(n7545), .B2(P2_REG1_REG_8__SCAN_IN), .A(n7534), .ZN(
        n7536) );
  XNOR2_X1 U8699 ( .A(n7536), .B(n7535), .ZN(n7539) );
  NOR2_X1 U8700 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8068), .ZN(n7537) );
  AOI21_X1 U8701 ( .B1(n10314), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n7537), .ZN(
        n7538) );
  OAI21_X1 U8702 ( .B1(n10329), .B2(n7539), .A(n7538), .ZN(n7544) );
  AOI211_X1 U8703 ( .C1(n7542), .C2(n7541), .A(n7540), .B(n10325), .ZN(n7543)
         );
  AOI211_X1 U8704 ( .C1(n10320), .C2(n7545), .A(n7544), .B(n7543), .ZN(n7546)
         );
  INV_X1 U8705 ( .A(n7546), .ZN(P2_U3253) );
  INV_X1 U8706 ( .A(n7547), .ZN(n7601) );
  AOI22_X1 U8707 ( .A1(n8038), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n8004), .ZN(n7548) );
  OAI21_X1 U8708 ( .B1(n7601), .B2(n8826), .A(n7548), .ZN(P1_U3340) );
  AOI22_X1 U8709 ( .A1(n8976), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n8993), .ZN(n7552) );
  NOR2_X1 U8710 ( .A1(n10325), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n7550) );
  NOR2_X1 U8711 ( .A1(n10329), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n7549) );
  NOR3_X1 U8712 ( .A1(n7550), .A2(n10320), .A3(n7549), .ZN(n7551) );
  MUX2_X1 U8713 ( .A(n7552), .B(n7551), .S(P2_IR_REG_0__SCAN_IN), .Z(n7554) );
  AOI22_X1 U8714 ( .A1(n10314), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n7553) );
  NAND2_X1 U8715 ( .A1(n7554), .A2(n7553), .ZN(P2_U3245) );
  OAI22_X1 U8716 ( .A1(n10377), .A2(n8922), .B1(n8913), .B2(n10438), .ZN(n7556) );
  NOR2_X1 U8717 ( .A1(n8897), .A2(n7687), .ZN(n7555) );
  AOI211_X1 U8718 ( .C1(P2_REG3_REG_2__SCAN_IN), .C2(n7557), .A(n7556), .B(
        n7555), .ZN(n7560) );
  OAI211_X1 U8719 ( .C1(n4920), .C2(n7558), .A(n7604), .B(n8905), .ZN(n7559)
         );
  NAND2_X1 U8720 ( .A1(n7560), .A2(n7559), .ZN(P2_U3239) );
  XNOR2_X1 U8721 ( .A(n7561), .B(n7685), .ZN(n7882) );
  XOR2_X1 U8722 ( .A(n7562), .B(n7561), .Z(n7564) );
  AOI21_X1 U8723 ( .B1(n7564), .B2(n10616), .A(n7563), .ZN(n7887) );
  AND2_X1 U8724 ( .A1(n7885), .A2(n7565), .ZN(n7566) );
  NOR2_X1 U8725 ( .A1(n7703), .A2(n7566), .ZN(n7879) );
  NAND2_X1 U8726 ( .A1(n7567), .A2(n6849), .ZN(n10673) );
  AOI22_X1 U8727 ( .A1(n7879), .A2(n10663), .B1(n10662), .B2(n7885), .ZN(n7568) );
  OAI211_X1 U8728 ( .C1(n10667), .C2(n7882), .A(n7887), .B(n7568), .ZN(n7570)
         );
  NAND2_X1 U8729 ( .A1(n7570), .A2(n10684), .ZN(n7569) );
  OAI21_X1 U8730 ( .B1(n10684), .B2(n6252), .A(n7569), .ZN(P2_U3454) );
  NAND2_X1 U8731 ( .A1(n7570), .A2(n10681), .ZN(n7571) );
  OAI21_X1 U8732 ( .B1(n10681), .B2(n7167), .A(n7571), .ZN(P2_U3521) );
  INV_X1 U8733 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n8223) );
  OR2_X1 U8734 ( .A1(n10281), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n7575) );
  AOI21_X1 U8735 ( .B1(n7585), .B2(n10553), .A(n7572), .ZN(n10286) );
  INV_X1 U8736 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n7573) );
  MUX2_X1 U8737 ( .A(n7573), .B(P1_REG1_REG_9__SCAN_IN), .S(n10281), .Z(n10287) );
  NOR2_X1 U8738 ( .A1(n10286), .A2(n10287), .ZN(n10285) );
  INV_X1 U8739 ( .A(n10285), .ZN(n7574) );
  AND2_X1 U8740 ( .A1(n7575), .A2(n7574), .ZN(n10296) );
  MUX2_X1 U8741 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n8223), .S(n7579), .Z(n10297) );
  NOR2_X1 U8742 ( .A1(n10296), .A2(n10297), .ZN(n10295) );
  AOI21_X1 U8743 ( .B1(n8223), .B2(n7579), .A(n10295), .ZN(n7578) );
  INV_X1 U8744 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n7576) );
  AOI22_X1 U8745 ( .A1(n7711), .A2(n7576), .B1(P1_REG1_REG_11__SCAN_IN), .B2(
        n7594), .ZN(n7577) );
  NOR2_X1 U8746 ( .A1(n7578), .A2(n7577), .ZN(n7713) );
  AOI21_X1 U8747 ( .B1(n7578), .B2(n7577), .A(n7713), .ZN(n7600) );
  NAND2_X1 U8748 ( .A1(P1_REG2_REG_10__SCAN_IN), .A2(n10293), .ZN(n7587) );
  INV_X1 U8749 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7580) );
  MUX2_X1 U8750 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n7580), .S(n7579), .Z(n7581)
         );
  INV_X1 U8751 ( .A(n7581), .ZN(n10301) );
  NAND2_X1 U8752 ( .A1(n10281), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n7586) );
  INV_X1 U8753 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n7582) );
  MUX2_X1 U8754 ( .A(n7582), .B(P1_REG2_REG_9__SCAN_IN), .S(n10281), .Z(n7583)
         );
  INV_X1 U8755 ( .A(n7583), .ZN(n10283) );
  AOI21_X1 U8756 ( .B1(n7342), .B2(n7585), .A(n7584), .ZN(n10284) );
  NAND2_X1 U8757 ( .A1(n10283), .A2(n10284), .ZN(n10282) );
  NAND2_X1 U8758 ( .A1(n7586), .A2(n10282), .ZN(n10302) );
  NAND2_X1 U8759 ( .A1(n10301), .A2(n10302), .ZN(n10300) );
  NAND2_X1 U8760 ( .A1(n7587), .A2(n10300), .ZN(n7597) );
  NAND2_X1 U8761 ( .A1(P1_REG2_REG_11__SCAN_IN), .A2(n7597), .ZN(n7589) );
  OAI21_X1 U8762 ( .B1(n7589), .B2(n7588), .A(n9836), .ZN(n7592) );
  AND2_X1 U8763 ( .A1(P1_U3084), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n8331) );
  INV_X1 U8764 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n7590) );
  NOR2_X1 U8765 ( .A1(n10342), .A2(n7590), .ZN(n7591) );
  AOI211_X1 U8766 ( .C1(n7711), .C2(n7592), .A(n8331), .B(n7591), .ZN(n7599)
         );
  INV_X1 U8767 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7593) );
  NAND2_X1 U8768 ( .A1(n7594), .A2(n7593), .ZN(n7596) );
  OAI211_X1 U8769 ( .C1(n7597), .C2(n7596), .A(n7718), .B(n10335), .ZN(n7598)
         );
  OAI211_X1 U8770 ( .C1(n7600), .C2(n10299), .A(n7599), .B(n7598), .ZN(
        P1_U3252) );
  INV_X1 U8771 ( .A(n8122), .ZN(n8118) );
  OAI222_X1 U8772 ( .A1(n4846), .A2(n8118), .B1(n8243), .B2(n7601), .C1(n9387), 
        .C2(n5457), .ZN(P2_U3345) );
  INV_X1 U8773 ( .A(n7602), .ZN(n7603) );
  AOI21_X1 U8774 ( .B1(n7604), .B2(n7603), .A(n8927), .ZN(n7607) );
  NOR3_X1 U8775 ( .A1(n8902), .A2(n6860), .A3(n7605), .ZN(n7606) );
  OAI21_X1 U8776 ( .B1(n7607), .B2(n7606), .A(n7782), .ZN(n7611) );
  MUX2_X1 U8777 ( .A(n8910), .B(P2_U3152), .S(P2_REG3_REG_3__SCAN_IN), .Z(
        n7609) );
  OAI22_X1 U8778 ( .A1(n10392), .A2(n8922), .B1(n8913), .B2(n7777), .ZN(n7608)
         );
  AOI211_X1 U8779 ( .C1(n8911), .C2(n6242), .A(n7609), .B(n7608), .ZN(n7610)
         );
  NAND2_X1 U8780 ( .A1(n7611), .A2(n7610), .ZN(P2_U3220) );
  AOI21_X1 U8781 ( .B1(n7613), .B2(P2_REG2_REG_9__SCAN_IN), .A(n7612), .ZN(
        n7616) );
  NAND2_X1 U8782 ( .A1(n7940), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n7614) );
  OAI21_X1 U8783 ( .B1(n7940), .B2(P2_REG2_REG_10__SCAN_IN), .A(n7614), .ZN(
        n7615) );
  AOI211_X1 U8784 ( .C1(n7616), .C2(n7615), .A(n7939), .B(n10325), .ZN(n7626)
         );
  NOR2_X1 U8785 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6356), .ZN(n7617) );
  AOI21_X1 U8786 ( .B1(n10314), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n7617), .ZN(
        n7624) );
  OAI21_X1 U8787 ( .B1(n7619), .B2(n7527), .A(n7618), .ZN(n7622) );
  INV_X1 U8788 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n7620) );
  MUX2_X1 U8789 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n7620), .S(n7940), .Z(n7621)
         );
  NAND2_X1 U8790 ( .A1(n7621), .A2(n7622), .ZN(n7931) );
  OAI211_X1 U8791 ( .C1(n7622), .C2(n7621), .A(n8993), .B(n7931), .ZN(n7623)
         );
  OAI211_X1 U8792 ( .C1(n8998), .C2(n7932), .A(n7624), .B(n7623), .ZN(n7625)
         );
  OR2_X1 U8793 ( .A1(n7626), .A2(n7625), .ZN(P2_U3255) );
  AOI22_X1 U8794 ( .A1(n10563), .A2(P1_REG2_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(n10561), .ZN(n7631) );
  OR2_X1 U8795 ( .A1(n7627), .A2(n7668), .ZN(n7628) );
  OAI21_X1 U8796 ( .B1(n10558), .B2(n10042), .A(n7629), .ZN(n7630) );
  OAI211_X1 U8797 ( .C1(n7632), .C2(n10563), .A(n7631), .B(n7630), .ZN(
        P1_U3291) );
  OAI22_X1 U8798 ( .A1(n10403), .A2(n8701), .B1(n7633), .B2(n8702), .ZN(n7634)
         );
  XNOR2_X1 U8799 ( .A(n7634), .B(n8711), .ZN(n7799) );
  OR2_X1 U8800 ( .A1(n10403), .A2(n8713), .ZN(n7636) );
  NAND2_X1 U8801 ( .A1(n7753), .A2(n8721), .ZN(n7635) );
  NAND2_X1 U8802 ( .A1(n7636), .A2(n7635), .ZN(n7797) );
  XNOR2_X1 U8803 ( .A(n7799), .B(n7797), .ZN(n7648) );
  OAI22_X1 U8804 ( .A1(n7763), .A2(n8701), .B1(n7676), .B2(n8702), .ZN(n7639)
         );
  XNOR2_X1 U8805 ( .A(n7639), .B(n8711), .ZN(n7644) );
  INV_X1 U8806 ( .A(n7644), .ZN(n7642) );
  NAND2_X1 U8807 ( .A1(n10364), .A2(n8721), .ZN(n7640) );
  NAND2_X1 U8808 ( .A1(n7642), .A2(n7641), .ZN(n7645) );
  NAND2_X1 U8809 ( .A1(n7644), .A2(n7643), .ZN(n7646) );
  NAND2_X1 U8810 ( .A1(n9520), .A2(n7646), .ZN(n7647) );
  OAI21_X1 U8811 ( .B1(n7648), .B2(n7647), .A(n9491), .ZN(n7660) );
  NOR2_X1 U8812 ( .A1(n7650), .A2(n7649), .ZN(n7651) );
  AND2_X1 U8813 ( .A1(n7377), .A2(n7651), .ZN(n7653) );
  NAND2_X1 U8814 ( .A1(n7653), .A2(n7652), .ZN(n7655) );
  AOI21_X1 U8815 ( .B1(n7655), .B2(P1_STATE_REG_SCAN_IN), .A(n7654), .ZN(n9516) );
  AOI22_X1 U8816 ( .A1(n7364), .A2(n9545), .B1(n7753), .B2(n9564), .ZN(n7658)
         );
  AOI21_X1 U8817 ( .B1(n5029), .B2(n9558), .A(n7656), .ZN(n7657) );
  OAI211_X1 U8818 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n9516), .A(n7658), .B(
        n7657), .ZN(n7659) );
  AOI21_X1 U8819 ( .B1(n7660), .B2(n9536), .A(n7659), .ZN(n7661) );
  INV_X1 U8820 ( .A(n7661), .ZN(P1_U3216) );
  XNOR2_X1 U8821 ( .A(n7662), .B(n7666), .ZN(n10371) );
  NAND2_X1 U8822 ( .A1(n7663), .A2(n9991), .ZN(n9998) );
  OAI21_X1 U8823 ( .B1(n7666), .B2(n7665), .A(n7664), .ZN(n7673) );
  OAI21_X1 U8824 ( .B1(n8185), .B2(n7668), .A(n7667), .ZN(n7669) );
  NAND2_X1 U8825 ( .A1(n7670), .A2(n7669), .ZN(n10550) );
  AOI22_X1 U8826 ( .A1(n5777), .A2(n10539), .B1(n10540), .B2(n7491), .ZN(n7671) );
  OAI21_X1 U8827 ( .B1(n10371), .B2(n10550), .A(n7671), .ZN(n7672) );
  AOI21_X1 U8828 ( .B1(n10546), .B2(n7673), .A(n7672), .ZN(n10369) );
  MUX2_X1 U8829 ( .A(n7674), .B(n10369), .S(n10568), .Z(n7679) );
  AOI21_X1 U8830 ( .B1(n10364), .B2(n7758), .A(n7749), .ZN(n10367) );
  INV_X1 U8831 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n7675) );
  OAI22_X1 U8832 ( .A1(n10565), .A2(n7676), .B1(n10005), .B2(n7675), .ZN(n7677) );
  AOI21_X1 U8833 ( .B1(n10367), .B2(n10558), .A(n7677), .ZN(n7678) );
  OAI211_X1 U8834 ( .C1(n10371), .C2(n8598), .A(n7679), .B(n7678), .ZN(
        P1_U3289) );
  INV_X1 U8835 ( .A(n9798), .ZN(n9804) );
  INV_X1 U8836 ( .A(n7680), .ZN(n7683) );
  INV_X1 U8837 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n7681) );
  OAI222_X1 U8838 ( .A1(P1_U3084), .A2(n9804), .B1(n8826), .B2(n7683), .C1(
        n7681), .C2(n10209), .ZN(P1_U3339) );
  INV_X1 U8839 ( .A(n8436), .ZN(n8428) );
  INV_X1 U8840 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n7682) );
  OAI222_X1 U8841 ( .A1(P2_U3152), .A2(n8428), .B1(n8243), .B2(n7683), .C1(
        n7682), .C2(n9387), .ZN(P2_U3344) );
  NAND2_X1 U8842 ( .A1(n8946), .A2(n7885), .ZN(n7684) );
  NAND2_X1 U8843 ( .A1(n7685), .A2(n7684), .ZN(n7689) );
  NAND2_X1 U8844 ( .A1(n7687), .A2(n7686), .ZN(n7688) );
  NAND2_X1 U8845 ( .A1(n7689), .A2(n7688), .ZN(n7726) );
  XNOR2_X1 U8846 ( .A(n7726), .B(n7694), .ZN(n10376) );
  NAND2_X1 U8847 ( .A1(n7691), .A2(n7690), .ZN(n7700) );
  INV_X2 U8848 ( .A(n10448), .ZN(n9157) );
  NAND2_X1 U8849 ( .A1(n6849), .A2(n7692), .ZN(n7850) );
  NOR2_X1 U8850 ( .A1(n9157), .A2(n7850), .ZN(n10627) );
  INV_X1 U8851 ( .A(n10627), .ZN(n7741) );
  OAI21_X1 U8852 ( .B1(n7695), .B2(n7694), .A(n7693), .ZN(n7697) );
  OAI22_X1 U8853 ( .A1(n10438), .A2(n10613), .B1(n7687), .B2(n10611), .ZN(
        n7696) );
  AOI21_X1 U8854 ( .B1(n7697), .B2(n10616), .A(n7696), .ZN(n7698) );
  OAI21_X1 U8855 ( .B1(n10376), .B2(n10619), .A(n7698), .ZN(n10379) );
  NAND2_X1 U8856 ( .A1(n10379), .A2(n10448), .ZN(n7709) );
  NOR2_X2 U8857 ( .A1(n9157), .A2(n7699), .ZN(n10451) );
  INV_X1 U8858 ( .A(n7700), .ZN(n7702) );
  NAND2_X1 U8859 ( .A1(n7702), .A2(n7701), .ZN(n10454) );
  NAND2_X1 U8860 ( .A1(n7703), .A2(n10377), .ZN(n7734) );
  OR2_X1 U8861 ( .A1(n7703), .A2(n10377), .ZN(n7704) );
  NAND2_X1 U8862 ( .A1(n7734), .A2(n7704), .ZN(n10378) );
  INV_X2 U8863 ( .A(n10446), .ZN(n10629) );
  AOI22_X1 U8864 ( .A1(n9157), .A2(P2_REG2_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(n10629), .ZN(n7705) );
  OAI21_X1 U8865 ( .B1(n10454), .B2(n10378), .A(n7705), .ZN(n7706) );
  AOI21_X1 U8866 ( .B1(n10451), .B2(n7707), .A(n7706), .ZN(n7708) );
  OAI211_X1 U8867 ( .C1(n10376), .C2(n7741), .A(n7709), .B(n7708), .ZN(
        P2_U3294) );
  NAND2_X1 U8868 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(n8945), .ZN(n7710) );
  OAI21_X1 U8869 ( .B1(n9144), .B2(n8945), .A(n7710), .ZN(P2_U3577) );
  NOR2_X1 U8870 ( .A1(n7711), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n7712) );
  NOR2_X1 U8871 ( .A1(n7713), .A2(n7712), .ZN(n7715) );
  XNOR2_X1 U8872 ( .A(n7836), .B(P1_REG1_REG_12__SCAN_IN), .ZN(n7714) );
  NOR2_X1 U8873 ( .A1(n7715), .A2(n7714), .ZN(n7830) );
  AOI21_X1 U8874 ( .B1(n7715), .B2(n7714), .A(n7830), .ZN(n7724) );
  NAND2_X1 U8875 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n7836), .ZN(n7716) );
  OAI21_X1 U8876 ( .B1(n7836), .B2(P1_REG2_REG_12__SCAN_IN), .A(n7716), .ZN(
        n7717) );
  NOR2_X1 U8877 ( .A1(n7717), .A2(n7718), .ZN(n7835) );
  AOI211_X1 U8878 ( .C1(n7718), .C2(n7717), .A(n7835), .B(n10269), .ZN(n7722)
         );
  INV_X1 U8879 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n8756) );
  NOR2_X1 U8880 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7719), .ZN(n8360) );
  AOI21_X1 U8881 ( .B1(n10339), .B2(n7836), .A(n8360), .ZN(n7720) );
  OAI21_X1 U8882 ( .B1(n8756), .B2(n10342), .A(n7720), .ZN(n7721) );
  NOR2_X1 U8883 ( .A1(n7722), .A2(n7721), .ZN(n7723) );
  OAI21_X1 U8884 ( .B1(n7724), .B2(n10299), .A(n7723), .ZN(P1_U3253) );
  NAND2_X1 U8885 ( .A1(n7726), .A2(n7725), .ZN(n7728) );
  NAND2_X1 U8886 ( .A1(n6860), .A2(n10377), .ZN(n7727) );
  NAND2_X1 U8887 ( .A1(n7728), .A2(n7727), .ZN(n7861) );
  XNOR2_X1 U8888 ( .A(n7861), .B(n7730), .ZN(n10391) );
  OAI21_X1 U8889 ( .B1(n7730), .B2(n6651), .A(n7729), .ZN(n7732) );
  OAI22_X1 U8890 ( .A1(n7777), .A2(n10613), .B1(n6860), .B2(n10611), .ZN(n7731) );
  AOI21_X1 U8891 ( .B1(n7732), .B2(n10616), .A(n7731), .ZN(n7733) );
  OAI21_X1 U8892 ( .B1(n10391), .B2(n10619), .A(n7733), .ZN(n10394) );
  NAND2_X1 U8893 ( .A1(n10394), .A2(n10448), .ZN(n7740) );
  OAI22_X1 U8894 ( .A1(n10448), .A2(n6266), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n10446), .ZN(n7737) );
  NAND2_X1 U8895 ( .A1(n7734), .A2(n7738), .ZN(n7735) );
  NAND2_X1 U8896 ( .A1(n10431), .A2(n7735), .ZN(n10393) );
  NOR2_X1 U8897 ( .A1(n10393), .A2(n10454), .ZN(n7736) );
  AOI211_X1 U8898 ( .C1(n10451), .C2(n7738), .A(n7737), .B(n7736), .ZN(n7739)
         );
  OAI211_X1 U8899 ( .C1(n10391), .C2(n7741), .A(n7740), .B(n7739), .ZN(
        P2_U3293) );
  INV_X1 U8900 ( .A(n7743), .ZN(n7744) );
  XNOR2_X1 U8901 ( .A(n7742), .B(n7744), .ZN(n10383) );
  NAND2_X1 U8902 ( .A1(n7745), .A2(n10546), .ZN(n7747) );
  AOI22_X1 U8903 ( .A1(n10539), .A2(n7364), .B1(n5029), .B2(n10540), .ZN(n7746) );
  OAI211_X1 U8904 ( .C1(n10383), .C2(n10550), .A(n7747), .B(n7746), .ZN(n10385) );
  NAND2_X1 U8905 ( .A1(n10385), .A2(n10568), .ZN(n7755) );
  OAI22_X1 U8906 ( .A1(n10568), .A2(n7748), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n10005), .ZN(n7752) );
  OR2_X1 U8907 ( .A1(n7749), .A2(n7633), .ZN(n7750) );
  NAND2_X1 U8908 ( .A1(n10400), .A2(n7750), .ZN(n10384) );
  NOR2_X1 U8909 ( .A1(n10384), .A2(n10046), .ZN(n7751) );
  AOI211_X1 U8910 ( .C1(n10042), .C2(n7753), .A(n7752), .B(n7751), .ZN(n7754)
         );
  OAI211_X1 U8911 ( .C1(n10383), .C2(n8598), .A(n7755), .B(n7754), .ZN(
        P1_U3288) );
  INV_X1 U8912 ( .A(n7756), .ZN(n7757) );
  XNOR2_X1 U8913 ( .A(n6077), .B(n7757), .ZN(n10361) );
  INV_X1 U8914 ( .A(n10361), .ZN(n7769) );
  OAI211_X1 U8915 ( .C1(n10357), .C2(n7759), .A(n10366), .B(n7758), .ZN(n10355) );
  OAI21_X1 U8916 ( .B1(n7761), .B2(n6077), .A(n7760), .ZN(n7762) );
  INV_X1 U8917 ( .A(n10550), .ZN(n10522) );
  AOI222_X1 U8918 ( .A1(n7762), .A2(n10546), .B1(n10522), .B2(n10361), .C1(
        n7380), .C2(n10540), .ZN(n10358) );
  NOR2_X1 U8919 ( .A1(n7763), .A2(n10489), .ZN(n10354) );
  AOI21_X1 U8920 ( .B1(n10561), .B2(P1_REG3_REG_1__SCAN_IN), .A(n10354), .ZN(
        n7764) );
  OAI211_X1 U8921 ( .C1(n9991), .C2(n10355), .A(n10358), .B(n7764), .ZN(n7765)
         );
  NAND2_X1 U8922 ( .A1(n7765), .A2(n10568), .ZN(n7768) );
  AOI22_X1 U8923 ( .A1(n10042), .A2(n7766), .B1(n9977), .B2(
        P1_REG2_REG_1__SCAN_IN), .ZN(n7767) );
  OAI211_X1 U8924 ( .C1(n7769), .C2(n8598), .A(n7768), .B(n7767), .ZN(P1_U3290) );
  OAI21_X1 U8925 ( .B1(n8922), .B2(n8059), .A(n7771), .ZN(n7774) );
  OAI22_X1 U8926 ( .A1(n8897), .A2(n7777), .B1(n7772), .B2(n8913), .ZN(n7773)
         );
  AOI211_X1 U8927 ( .C1(n8054), .C2(n8910), .A(n7774), .B(n7773), .ZN(n7780)
         );
  OAI22_X1 U8928 ( .A1(n8902), .A2(n7777), .B1(n8927), .B2(n7776), .ZN(n7778)
         );
  NAND3_X1 U8929 ( .A1(n7781), .A2(n5317), .A3(n7778), .ZN(n7779) );
  OAI211_X1 U8930 ( .C1(n7770), .C2(n8927), .A(n7780), .B(n7779), .ZN(P2_U3229) );
  OAI21_X1 U8931 ( .B1(n7784), .B2(n7782), .A(n7781), .ZN(n7791) );
  NOR3_X1 U8932 ( .A1(n8902), .A2(n7784), .A3(n7783), .ZN(n7785) );
  OAI21_X1 U8933 ( .B1(n7785), .B2(n8911), .A(n8944), .ZN(n7789) );
  INV_X1 U8934 ( .A(n8913), .ZN(n8777) );
  OAI21_X1 U8935 ( .B1(n8922), .B2(n10434), .A(n7786), .ZN(n7787) );
  AOI21_X1 U8936 ( .B1(n8777), .B2(n8942), .A(n7787), .ZN(n7788) );
  OAI211_X1 U8937 ( .C1(n8921), .C2(n10447), .A(n7789), .B(n7788), .ZN(n7790)
         );
  AOI21_X1 U8938 ( .B1(n7791), .B2(n8905), .A(n7790), .ZN(n7792) );
  INV_X1 U8939 ( .A(n7792), .ZN(P2_U3232) );
  OAI22_X1 U8940 ( .A1(n7794), .A2(n8701), .B1(n10423), .B2(n8702), .ZN(n7793)
         );
  XNOR2_X1 U8941 ( .A(n7793), .B(n8711), .ZN(n7801) );
  OR2_X1 U8942 ( .A1(n7794), .A2(n8713), .ZN(n7796) );
  NAND2_X1 U8943 ( .A1(n9496), .A2(n8721), .ZN(n7795) );
  NAND2_X1 U8944 ( .A1(n7796), .A2(n7795), .ZN(n7802) );
  XNOR2_X1 U8945 ( .A(n7801), .B(n7802), .ZN(n9493) );
  INV_X1 U8946 ( .A(n7797), .ZN(n7798) );
  NAND2_X1 U8947 ( .A1(n7799), .A2(n7798), .ZN(n9490) );
  AND2_X1 U8948 ( .A1(n9493), .A2(n9490), .ZN(n7800) );
  NAND2_X1 U8949 ( .A1(n9491), .A2(n7800), .ZN(n9492) );
  INV_X1 U8950 ( .A(n7801), .ZN(n7803) );
  NAND2_X1 U8951 ( .A1(n7803), .A2(n7802), .ZN(n7804) );
  NAND2_X1 U8952 ( .A1(n9492), .A2(n7804), .ZN(n7893) );
  OAI22_X1 U8953 ( .A1(n10491), .A2(n8701), .B1(n10463), .B2(n8702), .ZN(n7805) );
  XNOR2_X1 U8954 ( .A(n7805), .B(n8711), .ZN(n7894) );
  OR2_X1 U8955 ( .A1(n10491), .A2(n8713), .ZN(n7807) );
  NAND2_X1 U8956 ( .A1(n7997), .A2(n8721), .ZN(n7806) );
  AND2_X1 U8957 ( .A1(n7807), .A2(n7806), .ZN(n7895) );
  XNOR2_X1 U8958 ( .A(n7894), .B(n7895), .ZN(n7808) );
  XNOR2_X1 U8959 ( .A(n7893), .B(n7808), .ZN(n7816) );
  AOI21_X1 U8960 ( .B1(n7364), .B2(n9558), .A(n7809), .ZN(n7814) );
  INV_X1 U8961 ( .A(n7998), .ZN(n7810) );
  OR2_X1 U8962 ( .A1(n9516), .A2(n7810), .ZN(n7813) );
  NAND2_X1 U8963 ( .A1(n9564), .A2(n7997), .ZN(n7812) );
  NAND2_X1 U8964 ( .A1(n7994), .A2(n9545), .ZN(n7811) );
  NAND4_X1 U8965 ( .A1(n7814), .A2(n7813), .A3(n7812), .A4(n7811), .ZN(n7815)
         );
  AOI21_X1 U8966 ( .B1(n7816), .B2(n9536), .A(n7815), .ZN(n7817) );
  INV_X1 U8967 ( .A(n7817), .ZN(P1_U3225) );
  INV_X1 U8968 ( .A(n8978), .ZN(n8437) );
  INV_X1 U8969 ( .A(n7818), .ZN(n7820) );
  OAI222_X1 U8970 ( .A1(n4846), .A2(n8437), .B1(n8243), .B2(n7820), .C1(n9387), 
        .C2(n5467), .ZN(P2_U3343) );
  INV_X1 U8971 ( .A(n9810), .ZN(n9820) );
  OAI222_X1 U8972 ( .A1(n9820), .A2(P1_U3084), .B1(n8826), .B2(n7820), .C1(
        n7819), .C2(n10196), .ZN(P1_U3338) );
  NAND2_X1 U8973 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(n8945), .ZN(n7821) );
  OAI21_X1 U8974 ( .B1(n9059), .B2(n8945), .A(n7821), .ZN(P2_U3579) );
  OAI21_X1 U8975 ( .B1(n8922), .B2(n10509), .A(n7822), .ZN(n7824) );
  OAI22_X1 U8976 ( .A1(n8897), .A2(n10439), .B1(n8065), .B2(n8913), .ZN(n7823)
         );
  AOI211_X1 U8977 ( .C1(n7868), .C2(n8910), .A(n7824), .B(n7823), .ZN(n7828)
         );
  OAI22_X1 U8978 ( .A1(n8902), .A2(n10439), .B1(n8927), .B2(n7825), .ZN(n7826)
         );
  NAND3_X1 U8979 ( .A1(n7770), .A2(n4918), .A3(n7826), .ZN(n7827) );
  OAI211_X1 U8980 ( .C1(n7829), .C2(n8927), .A(n7828), .B(n7827), .ZN(P2_U3241) );
  XNOR2_X1 U8981 ( .A(n8038), .B(P1_REG1_REG_13__SCAN_IN), .ZN(n7834) );
  INV_X1 U8982 ( .A(n7836), .ZN(n7832) );
  INV_X1 U8983 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n7831) );
  AOI21_X1 U8984 ( .B1(n7832), .B2(n7831), .A(n7830), .ZN(n7833) );
  NOR2_X1 U8985 ( .A1(n7833), .A2(n7834), .ZN(n8039) );
  AOI21_X1 U8986 ( .B1(n7834), .B2(n7833), .A(n8039), .ZN(n7845) );
  AND2_X1 U8987 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n8484) );
  INV_X1 U8988 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n7842) );
  AOI21_X1 U8989 ( .B1(n7836), .B2(P1_REG2_REG_12__SCAN_IN), .A(n7835), .ZN(
        n7839) );
  NAND2_X1 U8990 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n8038), .ZN(n7837) );
  OAI21_X1 U8991 ( .B1(n8038), .B2(P1_REG2_REG_13__SCAN_IN), .A(n7837), .ZN(
        n7838) );
  NOR2_X1 U8992 ( .A1(n7839), .A2(n7838), .ZN(n8034) );
  AOI211_X1 U8993 ( .C1(n7839), .C2(n7838), .A(n8034), .B(n10269), .ZN(n7840)
         );
  INV_X1 U8994 ( .A(n7840), .ZN(n7841) );
  OAI21_X1 U8995 ( .B1(n7842), .B2(n10342), .A(n7841), .ZN(n7843) );
  AOI211_X1 U8996 ( .C1(n8038), .C2(n10339), .A(n8484), .B(n7843), .ZN(n7844)
         );
  OAI21_X1 U8997 ( .B1(n7845), .B2(n10299), .A(n7844), .ZN(P1_U3254) );
  INV_X1 U8998 ( .A(n7846), .ZN(n7849) );
  AOI22_X1 U8999 ( .A1(n8989), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n9378), .ZN(n7847) );
  OAI21_X1 U9000 ( .B1(n7849), .B2(n8243), .A(n7847), .ZN(P2_U3342) );
  AOI22_X1 U9001 ( .A1(n9840), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n8004), .ZN(n7848) );
  OAI21_X1 U9002 ( .B1(n7849), .B2(n8826), .A(n7848), .ZN(P1_U3337) );
  AND2_X1 U9003 ( .A1(n10619), .A2(n7850), .ZN(n7851) );
  AOI21_X1 U9004 ( .B1(n10634), .B2(n10454), .A(n7852), .ZN(n7853) );
  AOI21_X1 U9005 ( .B1(n10448), .B2(n7854), .A(n7853), .ZN(n7856) );
  AOI22_X1 U9006 ( .A1(n9157), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(n10629), .ZN(n7855) );
  OAI211_X1 U9007 ( .C1(n7857), .C2(n9255), .A(n7856), .B(n7855), .ZN(P2_U3296) );
  XNOR2_X1 U9008 ( .A(n7858), .B(n7866), .ZN(n7859) );
  OAI222_X1 U9009 ( .A1(n10613), .A2(n8065), .B1(n10611), .B2(n10439), .C1(
        n7859), .C2(n10436), .ZN(n10511) );
  INV_X1 U9010 ( .A(n10511), .ZN(n7875) );
  NAND2_X1 U9011 ( .A1(n10438), .A2(n10392), .ZN(n7862) );
  NAND2_X1 U9012 ( .A1(n10450), .A2(n8943), .ZN(n7863) );
  NAND2_X1 U9013 ( .A1(n10428), .A2(n7863), .ZN(n8057) );
  NAND2_X1 U9014 ( .A1(n10439), .A2(n8059), .ZN(n7864) );
  NAND2_X1 U9015 ( .A1(n8058), .A2(n8942), .ZN(n7865) );
  XNOR2_X1 U9016 ( .A(n7961), .B(n7866), .ZN(n10513) );
  INV_X1 U9017 ( .A(n9255), .ZN(n10456) );
  OR2_X1 U9018 ( .A1(n8053), .A2(n10509), .ZN(n7867) );
  NAND2_X1 U9019 ( .A1(n7983), .A2(n7867), .ZN(n10510) );
  INV_X1 U9020 ( .A(n7868), .ZN(n7869) );
  OAI22_X1 U9021 ( .A1(n10448), .A2(n7187), .B1(n7869), .B2(n10446), .ZN(n7870) );
  AOI21_X1 U9022 ( .B1(n10451), .B2(n7871), .A(n7870), .ZN(n7872) );
  OAI21_X1 U9023 ( .B1(n10510), .B2(n10454), .A(n7872), .ZN(n7873) );
  AOI21_X1 U9024 ( .B1(n10513), .B2(n10456), .A(n7873), .ZN(n7874) );
  OAI21_X1 U9025 ( .B1(n7875), .B2(n10631), .A(n7874), .ZN(P2_U3290) );
  INV_X1 U9026 ( .A(n7876), .ZN(n7877) );
  NAND2_X1 U9027 ( .A1(n7877), .A2(P2_U3966), .ZN(n7878) );
  OAI21_X1 U9028 ( .B1(n5585), .B2(P2_U3966), .A(n7878), .ZN(P2_U3581) );
  AOI22_X1 U9029 ( .A1(n10626), .A2(n7879), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n10629), .ZN(n7880) );
  OAI21_X1 U9030 ( .B1(n7881), .B2(n10448), .A(n7880), .ZN(n7884) );
  NOR2_X1 U9031 ( .A1(n7882), .A2(n9255), .ZN(n7883) );
  AOI211_X1 U9032 ( .C1(n10451), .C2(n7885), .A(n7884), .B(n7883), .ZN(n7886)
         );
  OAI21_X1 U9033 ( .B1(n9157), .B2(n7887), .A(n7886), .ZN(P2_U3295) );
  INV_X1 U9034 ( .A(n7888), .ZN(n7890) );
  AOI22_X1 U9035 ( .A1(n9849), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n8004), .ZN(n7889) );
  OAI21_X1 U9036 ( .B1(n7890), .B2(n8826), .A(n7889), .ZN(P1_U3336) );
  INV_X1 U9037 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7891) );
  INV_X1 U9038 ( .A(n9004), .ZN(n9008) );
  OAI222_X1 U9039 ( .A1(n9387), .A2(n7891), .B1(n8243), .B2(n7890), .C1(n9008), 
        .C2(n4846), .ZN(P2_U3341) );
  NAND2_X1 U9040 ( .A1(n7894), .A2(n7895), .ZN(n7892) );
  NAND2_X1 U9041 ( .A1(n7893), .A2(n7892), .ZN(n7899) );
  INV_X1 U9042 ( .A(n7894), .ZN(n7897) );
  INV_X1 U9043 ( .A(n7895), .ZN(n7896) );
  NAND2_X1 U9044 ( .A1(n7897), .A2(n7896), .ZN(n7898) );
  NAND2_X1 U9045 ( .A1(n7899), .A2(n7898), .ZN(n7925) );
  OAI22_X1 U9046 ( .A1(n8011), .A2(n8701), .B1(n10502), .B2(n8702), .ZN(n7900)
         );
  XNOR2_X1 U9047 ( .A(n7900), .B(n7496), .ZN(n7903) );
  OR2_X1 U9048 ( .A1(n8011), .A2(n8713), .ZN(n7902) );
  NAND2_X1 U9049 ( .A1(n7929), .A2(n8721), .ZN(n7901) );
  NAND2_X1 U9050 ( .A1(n7902), .A2(n7901), .ZN(n7904) );
  AND2_X1 U9051 ( .A1(n7903), .A2(n7904), .ZN(n7922) );
  INV_X1 U9052 ( .A(n7903), .ZN(n7906) );
  INV_X1 U9053 ( .A(n7904), .ZN(n7905) );
  NAND2_X1 U9054 ( .A1(n7906), .A2(n7905), .ZN(n7921) );
  OAI22_X1 U9055 ( .A1(n10490), .A2(n8701), .B1(n10518), .B2(n8702), .ZN(n7907) );
  XNOR2_X1 U9056 ( .A(n7907), .B(n8711), .ZN(n8095) );
  OR2_X1 U9057 ( .A1(n10490), .A2(n8713), .ZN(n7909) );
  NAND2_X1 U9058 ( .A1(n7914), .A2(n8721), .ZN(n7908) );
  NAND2_X1 U9059 ( .A1(n7909), .A2(n7908), .ZN(n8093) );
  XNOR2_X1 U9060 ( .A(n8095), .B(n8093), .ZN(n8091) );
  XOR2_X1 U9061 ( .A(n8092), .B(n8091), .Z(n7916) );
  NAND2_X1 U9062 ( .A1(n9556), .A2(n8015), .ZN(n7912) );
  AOI21_X1 U9063 ( .B1(n7994), .B2(n9558), .A(n7910), .ZN(n7911) );
  OAI211_X1 U9064 ( .C1(n8098), .C2(n9561), .A(n7912), .B(n7911), .ZN(n7913)
         );
  AOI21_X1 U9065 ( .B1(n7914), .B2(n9564), .A(n7913), .ZN(n7915) );
  OAI21_X1 U9066 ( .B1(n7916), .B2(n9566), .A(n7915), .ZN(P1_U3211) );
  INV_X1 U9067 ( .A(n10506), .ZN(n7920) );
  NAND2_X1 U9068 ( .A1(P1_U3084), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n10279) );
  INV_X1 U9069 ( .A(n10279), .ZN(n7917) );
  AOI21_X1 U9070 ( .B1(n9791), .B2(n9558), .A(n7917), .ZN(n7919) );
  NAND2_X1 U9071 ( .A1(n10541), .A2(n9545), .ZN(n7918) );
  OAI211_X1 U9072 ( .C1(n9516), .C2(n7920), .A(n7919), .B(n7918), .ZN(n7928)
         );
  INV_X1 U9073 ( .A(n7921), .ZN(n7923) );
  NOR2_X1 U9074 ( .A1(n7923), .A2(n7922), .ZN(n7924) );
  XNOR2_X1 U9075 ( .A(n7925), .B(n7924), .ZN(n7926) );
  NOR2_X1 U9076 ( .A1(n7926), .A2(n9566), .ZN(n7927) );
  AOI211_X1 U9077 ( .C1(n7929), .C2(n9564), .A(n7928), .B(n7927), .ZN(n7930)
         );
  INV_X1 U9078 ( .A(n7930), .ZN(P1_U3237) );
  INV_X1 U9079 ( .A(n8963), .ZN(n7933) );
  INV_X1 U9080 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n10645) );
  MUX2_X1 U9081 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n10645), .S(n8963), .Z(n8965) );
  OAI21_X1 U9082 ( .B1(n7932), .B2(n7620), .A(n7931), .ZN(n8966) );
  NAND2_X1 U9083 ( .A1(n8965), .A2(n8966), .ZN(n8964) );
  OAI21_X1 U9084 ( .B1(n7933), .B2(n10645), .A(n8964), .ZN(n7936) );
  INV_X1 U9085 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7934) );
  MUX2_X1 U9086 ( .A(n7934), .B(P2_REG1_REG_12__SCAN_IN), .S(n8026), .Z(n7935)
         );
  NOR2_X1 U9087 ( .A1(n7935), .A2(n7936), .ZN(n8021) );
  AOI21_X1 U9088 ( .B1(n7936), .B2(n7935), .A(n8021), .ZN(n7938) );
  NOR2_X1 U9089 ( .A1(n6392), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8405) );
  AOI21_X1 U9090 ( .B1(n10314), .B2(P2_ADDR_REG_12__SCAN_IN), .A(n8405), .ZN(
        n7937) );
  OAI21_X1 U9091 ( .B1(n10329), .B2(n7938), .A(n7937), .ZN(n7946) );
  MUX2_X1 U9092 ( .A(n6378), .B(P2_REG2_REG_11__SCAN_IN), .S(n8963), .Z(n7941)
         );
  INV_X1 U9093 ( .A(n7941), .ZN(n8960) );
  MUX2_X1 U9094 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n6395), .S(n8026), .Z(n7942)
         );
  INV_X1 U9095 ( .A(n7942), .ZN(n7943) );
  NOR2_X1 U9096 ( .A1(n7943), .A2(n7944), .ZN(n8025) );
  AOI211_X1 U9097 ( .C1(n7944), .C2(n7943), .A(n8025), .B(n10325), .ZN(n7945)
         );
  AOI211_X1 U9098 ( .C1(n10320), .C2(n8026), .A(n7946), .B(n7945), .ZN(n7947)
         );
  INV_X1 U9099 ( .A(n7947), .ZN(P2_U3257) );
  INV_X1 U9100 ( .A(n7948), .ZN(n7952) );
  AOI21_X1 U9101 ( .B1(n7950), .B2(n7949), .A(n4975), .ZN(n7951) );
  OAI21_X1 U9102 ( .B1(n7952), .B2(n7951), .A(n10616), .ZN(n7955) );
  NAND2_X1 U9103 ( .A1(n8939), .A2(n9178), .ZN(n7954) );
  NAND2_X1 U9104 ( .A1(n8940), .A2(n9177), .ZN(n7953) );
  AND2_X1 U9105 ( .A1(n7954), .A2(n7953), .ZN(n8069) );
  NAND2_X1 U9106 ( .A1(n7955), .A2(n8069), .ZN(n10577) );
  NAND2_X1 U9107 ( .A1(n7981), .A2(n8131), .ZN(n7956) );
  NAND2_X1 U9108 ( .A1(n7956), .A2(n10663), .ZN(n7957) );
  OR2_X1 U9109 ( .A1(n7957), .A2(n8142), .ZN(n10573) );
  NOR2_X1 U9110 ( .A1(n9157), .A2(n4849), .ZN(n9266) );
  INV_X1 U9111 ( .A(n9266), .ZN(n7960) );
  AOI22_X1 U9112 ( .A1(n9157), .A2(P2_REG2_REG_8__SCAN_IN), .B1(n8071), .B2(
        n10629), .ZN(n7959) );
  NAND2_X1 U9113 ( .A1(n10451), .A2(n8131), .ZN(n7958) );
  OAI211_X1 U9114 ( .C1(n10573), .C2(n7960), .A(n7959), .B(n7958), .ZN(n7972)
         );
  INV_X1 U9115 ( .A(n7962), .ZN(n7974) );
  NAND2_X1 U9116 ( .A1(n8065), .A2(n7985), .ZN(n7965) );
  INV_X1 U9117 ( .A(n7965), .ZN(n7964) );
  AND2_X1 U9118 ( .A1(n7975), .A2(n7965), .ZN(n7966) );
  OR2_X1 U9119 ( .A1(n7967), .A2(n7966), .ZN(n7968) );
  NAND2_X1 U9120 ( .A1(n7969), .A2(n7968), .ZN(n7970) );
  NAND2_X1 U9121 ( .A1(n7970), .A2(n4975), .ZN(n10572) );
  AND3_X1 U9122 ( .A1(n8133), .A2(n10456), .A3(n10572), .ZN(n7971) );
  AOI211_X1 U9123 ( .C1(n10577), .C2(n10448), .A(n7972), .B(n7971), .ZN(n7973)
         );
  INV_X1 U9124 ( .A(n7973), .ZN(P2_U3288) );
  OR2_X1 U9125 ( .A1(n7961), .A2(n7974), .ZN(n7976) );
  NAND2_X1 U9126 ( .A1(n7976), .A2(n7975), .ZN(n7977) );
  XNOR2_X1 U9127 ( .A(n7977), .B(n6329), .ZN(n10529) );
  XNOR2_X1 U9128 ( .A(n7978), .B(n6329), .ZN(n7979) );
  AOI222_X1 U9129 ( .A1(n10616), .A2(n7979), .B1(n8941), .B2(n9177), .C1(n8135), .C2(n9178), .ZN(n10528) );
  MUX2_X1 U9130 ( .A(n7980), .B(n10528), .S(n10448), .Z(n7988) );
  INV_X1 U9131 ( .A(n7981), .ZN(n7982) );
  AOI21_X1 U9132 ( .B1(n10525), .B2(n7983), .A(n7982), .ZN(n10526) );
  OAI22_X1 U9133 ( .A1(n10634), .A2(n7985), .B1(n10446), .B2(n7984), .ZN(n7986) );
  AOI21_X1 U9134 ( .B1(n10526), .B2(n10626), .A(n7986), .ZN(n7987) );
  OAI211_X1 U9135 ( .C1(n10529), .C2(n9255), .A(n7988), .B(n7987), .ZN(
        P2_U3289) );
  INV_X1 U9136 ( .A(n7989), .ZN(n7990) );
  AOI21_X1 U9137 ( .B1(n7993), .B2(n7991), .A(n7990), .ZN(n10468) );
  INV_X1 U9138 ( .A(n10028), .ZN(n9911) );
  OAI22_X1 U9139 ( .A1(n10568), .A2(n7992), .B1(n10565), .B2(n10463), .ZN(
        n8001) );
  XNOR2_X1 U9140 ( .A(n7993), .B(n10486), .ZN(n7995) );
  AOI222_X1 U9141 ( .A1(n10546), .A2(n7995), .B1(n7364), .B2(n10540), .C1(
        n7994), .C2(n10539), .ZN(n10464) );
  INV_X1 U9142 ( .A(n7996), .ZN(n10482) );
  AOI211_X1 U9143 ( .C1(n7997), .C2(n10401), .A(n10582), .B(n10482), .ZN(
        n10461) );
  AOI22_X1 U9144 ( .A1(n10461), .A2(n8116), .B1(n10561), .B2(n7998), .ZN(n7999) );
  AOI21_X1 U9145 ( .B1(n10464), .B2(n7999), .A(n10563), .ZN(n8000) );
  AOI211_X1 U9146 ( .C1(n10468), .C2(n9911), .A(n8001), .B(n8000), .ZN(n8002)
         );
  INV_X1 U9147 ( .A(n8002), .ZN(P1_U3286) );
  INV_X1 U9148 ( .A(n8003), .ZN(n8007) );
  AOI22_X1 U9149 ( .A1(n9872), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n8004), .ZN(n8005) );
  OAI21_X1 U9150 ( .B1(n8007), .B2(n8826), .A(n8005), .ZN(P1_U3335) );
  AOI22_X1 U9151 ( .A1(n9017), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n9378), .ZN(n8006) );
  OAI21_X1 U9152 ( .B1(n8007), .B2(n8243), .A(n8006), .ZN(P2_U3340) );
  INV_X1 U9153 ( .A(n10543), .ZN(n8008) );
  AOI21_X1 U9154 ( .B1(n8013), .B2(n8009), .A(n8008), .ZN(n8010) );
  OAI222_X1 U9155 ( .A1(n7059), .A2(n8011), .B1(n10489), .B2(n8098), .C1(n7060), .C2(n8010), .ZN(n10519) );
  INV_X1 U9156 ( .A(n10519), .ZN(n8020) );
  XNOR2_X1 U9157 ( .A(n8012), .B(n8013), .ZN(n10521) );
  OAI211_X1 U9158 ( .C1(n10480), .C2(n10518), .A(n10366), .B(n10535), .ZN(
        n10516) );
  OR2_X1 U9159 ( .A1(n8014), .A2(n9991), .ZN(n8195) );
  AOI22_X1 U9160 ( .A1(n9977), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n8015), .B2(
        n10561), .ZN(n8017) );
  OR2_X1 U9161 ( .A1(n10565), .A2(n10518), .ZN(n8016) );
  OAI211_X1 U9162 ( .C1(n10516), .C2(n8195), .A(n8017), .B(n8016), .ZN(n8018)
         );
  AOI21_X1 U9163 ( .B1(n10521), .B2(n9911), .A(n8018), .ZN(n8019) );
  OAI21_X1 U9164 ( .B1(n8020), .B2(n9977), .A(n8019), .ZN(P1_U3284) );
  AOI21_X1 U9165 ( .B1(n8022), .B2(n7934), .A(n8021), .ZN(n8024) );
  INV_X1 U9166 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n10659) );
  AOI22_X1 U9167 ( .A1(n8122), .A2(n10659), .B1(P2_REG1_REG_13__SCAN_IN), .B2(
        n8118), .ZN(n8023) );
  NOR2_X1 U9168 ( .A1(n8024), .A2(n8023), .ZN(n8117) );
  AOI21_X1 U9169 ( .B1(n8024), .B2(n8023), .A(n8117), .ZN(n8033) );
  AOI22_X1 U9170 ( .A1(n8122), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n6408), .B2(
        n8118), .ZN(n8027) );
  OAI21_X1 U9171 ( .B1(n8028), .B2(n8027), .A(n8121), .ZN(n8031) );
  INV_X1 U9172 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n8759) );
  NAND2_X1 U9173 ( .A1(n10320), .A2(n8122), .ZN(n8029) );
  NAND2_X1 U9174 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_U3152), .ZN(n8313) );
  OAI211_X1 U9175 ( .C1(n8126), .C2(n8759), .A(n8029), .B(n8313), .ZN(n8030)
         );
  AOI21_X1 U9176 ( .B1(n8031), .B2(n8976), .A(n8030), .ZN(n8032) );
  OAI21_X1 U9177 ( .B1(n8033), .B2(n10329), .A(n8032), .ZN(P2_U3258) );
  AOI21_X1 U9178 ( .B1(n8038), .B2(P1_REG2_REG_13__SCAN_IN), .A(n8034), .ZN(
        n8037) );
  NAND2_X1 U9179 ( .A1(n9798), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n8035) );
  OAI21_X1 U9180 ( .B1(n9798), .B2(P1_REG2_REG_14__SCAN_IN), .A(n8035), .ZN(
        n8036) );
  NOR2_X1 U9181 ( .A1(n8037), .A2(n8036), .ZN(n9797) );
  AOI211_X1 U9182 ( .C1(n8037), .C2(n8036), .A(n9797), .B(n10269), .ZN(n8049)
         );
  XNOR2_X1 U9183 ( .A(n9798), .B(P1_REG1_REG_14__SCAN_IN), .ZN(n8043) );
  OR2_X1 U9184 ( .A1(n8038), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n8041) );
  INV_X1 U9185 ( .A(n8039), .ZN(n8040) );
  NOR2_X1 U9186 ( .A1(n8042), .A2(n8043), .ZN(n9802) );
  AOI21_X1 U9187 ( .B1(n8043), .B2(n8042), .A(n9802), .ZN(n8044) );
  NOR2_X1 U9188 ( .A1(n8044), .A2(n10299), .ZN(n8048) );
  INV_X1 U9189 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n8046) );
  NAND2_X1 U9190 ( .A1(n10339), .A2(n9798), .ZN(n8045) );
  NAND2_X1 U9191 ( .A1(P1_U3084), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n9405) );
  OAI211_X1 U9192 ( .C1(n10342), .C2(n8046), .A(n8045), .B(n9405), .ZN(n8047)
         );
  OR3_X1 U9193 ( .A1(n8049), .A2(n8048), .A3(n8047), .ZN(P1_U3255) );
  NAND2_X1 U9194 ( .A1(n10441), .A2(n8050), .ZN(n8051) );
  XOR2_X1 U9195 ( .A(n8051), .B(n8058), .Z(n8052) );
  AOI222_X1 U9196 ( .A1(n10616), .A2(n8052), .B1(n8941), .B2(n9178), .C1(n8943), .C2(n9177), .ZN(n10475) );
  AOI211_X1 U9197 ( .C1(n10473), .C2(n10432), .A(n10673), .B(n8053), .ZN(
        n10472) );
  AOI22_X1 U9198 ( .A1(n10472), .A2(n9029), .B1(n10629), .B2(n8054), .ZN(n8055) );
  NAND2_X1 U9199 ( .A1(n10475), .A2(n8055), .ZN(n8056) );
  MUX2_X1 U9200 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n8056), .S(n10448), .Z(n8061)
         );
  XOR2_X1 U9201 ( .A(n8057), .B(n8058), .Z(n10476) );
  OAI22_X1 U9202 ( .A1(n10476), .A2(n9255), .B1(n8059), .B2(n10634), .ZN(n8060) );
  OR2_X1 U9203 ( .A1(n8061), .A2(n8060), .ZN(P2_U3291) );
  INV_X1 U9204 ( .A(n8062), .ZN(n8063) );
  AOI21_X1 U9205 ( .B1(n7142), .B2(n8063), .A(n8927), .ZN(n8067) );
  NOR3_X1 U9206 ( .A1(n8902), .A2(n8065), .A3(n8064), .ZN(n8066) );
  OAI21_X1 U9207 ( .B1(n8067), .B2(n8066), .A(n8167), .ZN(n8073) );
  OAI22_X1 U9208 ( .A1(n8069), .A2(n8871), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8068), .ZN(n8070) );
  AOI21_X1 U9209 ( .B1(n8071), .B2(n8910), .A(n8070), .ZN(n8072) );
  OAI211_X1 U9210 ( .C1(n10575), .C2(n8922), .A(n8073), .B(n8072), .ZN(
        P2_U3223) );
  INV_X1 U9211 ( .A(n8078), .ZN(n8074) );
  XNOR2_X1 U9212 ( .A(n8075), .B(n8074), .ZN(n10586) );
  NAND2_X1 U9213 ( .A1(n10586), .A2(n10522), .ZN(n8083) );
  NAND2_X1 U9214 ( .A1(n8077), .A2(n8076), .ZN(n8079) );
  XNOR2_X1 U9215 ( .A(n8079), .B(n8078), .ZN(n8081) );
  OAI22_X1 U9216 ( .A1(n8098), .A2(n7059), .B1(n8267), .B2(n10489), .ZN(n8080)
         );
  AOI21_X1 U9217 ( .B1(n8081), .B2(n10546), .A(n8080), .ZN(n8082) );
  AND2_X1 U9218 ( .A1(n10536), .A2(n10580), .ZN(n8084) );
  OR2_X1 U9219 ( .A1(n8084), .A2(n8193), .ZN(n10583) );
  AOI22_X1 U9220 ( .A1(n9977), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n8158), .B2(
        n10561), .ZN(n8086) );
  NAND2_X1 U9221 ( .A1(n10580), .A2(n10042), .ZN(n8085) );
  OAI211_X1 U9222 ( .C1(n10583), .C2(n10046), .A(n8086), .B(n8085), .ZN(n8087)
         );
  AOI21_X1 U9223 ( .B1(n10586), .B2(n10559), .A(n8087), .ZN(n8088) );
  OAI21_X1 U9224 ( .B1(n10588), .B2(n9977), .A(n8088), .ZN(P1_U3282) );
  NAND2_X1 U9225 ( .A1(n8109), .A2(n8718), .ZN(n8089) );
  OAI21_X1 U9226 ( .B1(n8098), .B2(n8701), .A(n8089), .ZN(n8090) );
  XNOR2_X1 U9227 ( .A(n8090), .B(n7496), .ZN(n8152) );
  NAND2_X1 U9228 ( .A1(n8092), .A2(n8091), .ZN(n8097) );
  INV_X1 U9229 ( .A(n8093), .ZN(n8094) );
  NAND2_X1 U9230 ( .A1(n8095), .A2(n8094), .ZN(n8096) );
  OR2_X1 U9231 ( .A1(n8098), .A2(n8713), .ZN(n8100) );
  NAND2_X1 U9232 ( .A1(n8109), .A2(n8721), .ZN(n8099) );
  AND2_X1 U9233 ( .A1(n8100), .A2(n8099), .ZN(n8102) );
  INV_X1 U9234 ( .A(n8102), .ZN(n8101) );
  NAND2_X1 U9235 ( .A1(n8154), .A2(n8153), .ZN(n8103) );
  XOR2_X1 U9236 ( .A(n8152), .B(n8103), .Z(n8111) );
  NAND2_X1 U9237 ( .A1(n9556), .A2(n10562), .ZN(n8106) );
  AOI21_X1 U9238 ( .B1(n10541), .B2(n9558), .A(n8104), .ZN(n8105) );
  OAI211_X1 U9239 ( .C1(n8107), .C2(n9561), .A(n8106), .B(n8105), .ZN(n8108)
         );
  AOI21_X1 U9240 ( .B1(n8109), .B2(n9564), .A(n8108), .ZN(n8110) );
  OAI21_X1 U9241 ( .B1(n8111), .B2(n9566), .A(n8110), .ZN(P1_U3219) );
  INV_X1 U9242 ( .A(n8112), .ZN(n8115) );
  OAI222_X1 U9243 ( .A1(n9387), .A2(n8113), .B1(n8243), .B2(n8115), .C1(n9029), 
        .C2(P2_U3152), .ZN(P2_U3339) );
  OAI222_X1 U9244 ( .A1(n8116), .A2(P1_U3084), .B1(n8826), .B2(n8115), .C1(
        n8114), .C2(n10209), .ZN(P1_U3334) );
  AOI21_X1 U9245 ( .B1(n8118), .B2(n10659), .A(n8117), .ZN(n8120) );
  INV_X1 U9246 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n10670) );
  AOI22_X1 U9247 ( .A1(n8436), .A2(n10670), .B1(P2_REG1_REG_14__SCAN_IN), .B2(
        n8428), .ZN(n8119) );
  NOR2_X1 U9248 ( .A1(n8120), .A2(n8119), .ZN(n8427) );
  AOI21_X1 U9249 ( .B1(n8120), .B2(n8119), .A(n8427), .ZN(n8130) );
  AOI22_X1 U9250 ( .A1(n8436), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n6424), .B2(
        n8428), .ZN(n8124) );
  OAI21_X1 U9251 ( .B1(n8124), .B2(n8123), .A(n8435), .ZN(n8128) );
  INV_X1 U9252 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n8762) );
  NAND2_X1 U9253 ( .A1(n10320), .A2(n8436), .ZN(n8125) );
  NAND2_X1 U9254 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(n4846), .ZN(n8387) );
  OAI211_X1 U9255 ( .C1(n8126), .C2(n8762), .A(n8125), .B(n8387), .ZN(n8127)
         );
  AOI21_X1 U9256 ( .B1(n8128), .B2(n8976), .A(n8127), .ZN(n8129) );
  OAI21_X1 U9257 ( .B1(n8130), .B2(n10329), .A(n8129), .ZN(P2_U3259) );
  NAND2_X1 U9258 ( .A1(n8135), .A2(n8131), .ZN(n8132) );
  OAI21_X1 U9259 ( .B1(n8134), .B2(n8136), .A(n8234), .ZN(n10599) );
  INV_X1 U9260 ( .A(n10599), .ZN(n8141) );
  INV_X1 U9261 ( .A(n8246), .ZN(n8938) );
  AOI22_X1 U9262 ( .A1(n9177), .A2(n8135), .B1(n8938), .B2(n9178), .ZN(n8140)
         );
  OAI211_X1 U9263 ( .C1(n8138), .C2(n5343), .A(n10616), .B(n8137), .ZN(n8139)
         );
  OAI211_X1 U9264 ( .C1(n8141), .C2(n10619), .A(n8140), .B(n8139), .ZN(n10597)
         );
  INV_X1 U9265 ( .A(n10597), .ZN(n8148) );
  NAND2_X1 U9266 ( .A1(n8142), .A2(n10595), .ZN(n10605) );
  OR2_X1 U9267 ( .A1(n8142), .A2(n10595), .ZN(n8143) );
  NAND2_X1 U9268 ( .A1(n10605), .A2(n8143), .ZN(n10596) );
  AOI22_X1 U9269 ( .A1(n9157), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n8171), .B2(
        n10629), .ZN(n8145) );
  NAND2_X1 U9270 ( .A1(n10451), .A2(n8179), .ZN(n8144) );
  OAI211_X1 U9271 ( .C1(n10596), .C2(n10454), .A(n8145), .B(n8144), .ZN(n8146)
         );
  AOI21_X1 U9272 ( .B1(n10599), .B2(n10627), .A(n8146), .ZN(n8147) );
  OAI21_X1 U9273 ( .B1(n8148), .B2(n10631), .A(n8147), .ZN(P2_U3287) );
  NAND2_X1 U9274 ( .A1(n10580), .A2(n8718), .ZN(n8150) );
  NAND2_X1 U9275 ( .A1(n10538), .A2(n8721), .ZN(n8149) );
  NAND2_X1 U9276 ( .A1(n8150), .A2(n8149), .ZN(n8151) );
  XNOR2_X1 U9277 ( .A(n8151), .B(n8711), .ZN(n8258) );
  AOI22_X1 U9278 ( .A1(n10580), .A2(n8721), .B1(n8720), .B2(n10538), .ZN(n8257) );
  XNOR2_X1 U9279 ( .A(n8258), .B(n8257), .ZN(n8157) );
  INV_X1 U9280 ( .A(n8260), .ZN(n8156) );
  AOI21_X1 U9281 ( .B1(n8157), .B2(n8155), .A(n8156), .ZN(n8163) );
  AOI22_X1 U9282 ( .A1(n9790), .A2(n9558), .B1(P1_REG3_REG_9__SCAN_IN), .B2(
        P1_U3084), .ZN(n8160) );
  NAND2_X1 U9283 ( .A1(n9556), .A2(n8158), .ZN(n8159) );
  OAI211_X1 U9284 ( .C1(n8267), .C2(n9561), .A(n8160), .B(n8159), .ZN(n8161)
         );
  AOI21_X1 U9285 ( .B1(n10580), .B2(n9564), .A(n8161), .ZN(n8162) );
  OAI21_X1 U9286 ( .B1(n8163), .B2(n9566), .A(n8162), .ZN(P1_U3229) );
  INV_X1 U9287 ( .A(n8164), .ZN(n8242) );
  OAI222_X1 U9288 ( .A1(P1_U3084), .A2(n8166), .B1(n8826), .B2(n8242), .C1(
        n8165), .C2(n10209), .ZN(P1_U3333) );
  INV_X1 U9289 ( .A(n8167), .ZN(n8170) );
  NOR3_X1 U9290 ( .A1(n8902), .A2(n8175), .A3(n8168), .ZN(n8169) );
  AOI21_X1 U9291 ( .B1(n8170), .B2(n8905), .A(n8169), .ZN(n8181) );
  AOI22_X1 U9292 ( .A1(n8777), .A2(n8938), .B1(n8910), .B2(n8171), .ZN(n8174)
         );
  INV_X1 U9293 ( .A(n8172), .ZN(n8173) );
  OAI211_X1 U9294 ( .C1(n8175), .C2(n8897), .A(n8174), .B(n8173), .ZN(n8178)
         );
  NOR2_X1 U9295 ( .A1(n8176), .A2(n8927), .ZN(n8177) );
  AOI211_X1 U9296 ( .C1(n8179), .C2(n8915), .A(n8178), .B(n8177), .ZN(n8180)
         );
  OAI21_X1 U9297 ( .B1(n8182), .B2(n8181), .A(n8180), .ZN(P2_U3233) );
  INV_X1 U9298 ( .A(n8183), .ZN(n8202) );
  OAI222_X1 U9299 ( .A1(P1_U3084), .A2(n8185), .B1(n8826), .B2(n8202), .C1(
        n8184), .C2(n10209), .ZN(P1_U3332) );
  OAI21_X1 U9300 ( .B1(n8192), .B2(n8187), .A(n8186), .ZN(n8188) );
  AOI222_X1 U9301 ( .A1(n10546), .A2(n8188), .B1(n9788), .B2(n10539), .C1(
        n10538), .C2(n10540), .ZN(n8220) );
  INV_X1 U9302 ( .A(n8189), .ZN(n8190) );
  AOI21_X1 U9303 ( .B1(n8192), .B2(n8191), .A(n8190), .ZN(n8221) );
  INV_X1 U9304 ( .A(n8221), .ZN(n8200) );
  OAI21_X1 U9305 ( .B1(n8193), .B2(n8198), .A(n10366), .ZN(n8194) );
  NOR2_X1 U9306 ( .A1(n8194), .A2(n8212), .ZN(n8218) );
  INV_X1 U9307 ( .A(n8195), .ZN(n10026) );
  NAND2_X1 U9308 ( .A1(n8218), .A2(n10026), .ZN(n8197) );
  AOI22_X1 U9309 ( .A1(n9977), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n8270), .B2(
        n10561), .ZN(n8196) );
  OAI211_X1 U9310 ( .C1(n8198), .C2(n10565), .A(n8197), .B(n8196), .ZN(n8199)
         );
  AOI21_X1 U9311 ( .B1(n8200), .B2(n9911), .A(n8199), .ZN(n8201) );
  OAI21_X1 U9312 ( .B1(n9977), .B2(n8220), .A(n8201), .ZN(P1_U3281) );
  OAI222_X1 U9313 ( .A1(n9387), .A2(n8204), .B1(n4846), .B2(n8203), .C1(n8243), 
        .C2(n8202), .ZN(P2_U3337) );
  OAI21_X1 U9314 ( .B1(n8206), .B2(n8207), .A(n8205), .ZN(n10167) );
  XNOR2_X1 U9315 ( .A(n8208), .B(n8207), .ZN(n8209) );
  NOR2_X1 U9316 ( .A1(n8209), .A2(n7060), .ZN(n8211) );
  OAI22_X1 U9317 ( .A1(n8267), .A2(n7059), .B1(n8486), .B2(n10489), .ZN(n8210)
         );
  AOI211_X1 U9318 ( .C1(n10167), .C2(n10522), .A(n8211), .B(n8210), .ZN(n10171) );
  OR2_X1 U9319 ( .A1(n8212), .A2(n8337), .ZN(n8213) );
  AND2_X1 U9320 ( .A1(n8298), .A2(n8213), .ZN(n10169) );
  NAND2_X1 U9321 ( .A1(n10169), .A2(n10558), .ZN(n8215) );
  AOI22_X1 U9322 ( .A1(n10563), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n8334), .B2(
        n10561), .ZN(n8214) );
  OAI211_X1 U9323 ( .C1(n8337), .C2(n10565), .A(n8215), .B(n8214), .ZN(n8216)
         );
  AOI21_X1 U9324 ( .B1(n10167), .B2(n10559), .A(n8216), .ZN(n8217) );
  OAI21_X1 U9325 ( .B1(n10171), .B2(n9977), .A(n8217), .ZN(P1_U3280) );
  AOI21_X1 U9326 ( .B1(n10365), .B2(n8276), .A(n8218), .ZN(n8219) );
  OAI211_X1 U9327 ( .C1(n8221), .C2(n10460), .A(n8220), .B(n8219), .ZN(n8224)
         );
  NAND2_X1 U9328 ( .A1(n8224), .A2(n10590), .ZN(n8222) );
  OAI21_X1 U9329 ( .B1(n10590), .B2(n8223), .A(n8222), .ZN(P1_U3533) );
  INV_X1 U9330 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n8226) );
  NAND2_X1 U9331 ( .A1(n8224), .A2(n10594), .ZN(n8225) );
  OAI21_X1 U9332 ( .B1(n10594), .B2(n8226), .A(n8225), .ZN(P1_U3484) );
  XNOR2_X1 U9333 ( .A(n8227), .B(n8236), .ZN(n8230) );
  NOR2_X1 U9334 ( .A1(n8374), .A2(n10613), .ZN(n8229) );
  NOR2_X1 U9335 ( .A1(n8246), .A2(n10611), .ZN(n8228) );
  OR2_X1 U9336 ( .A1(n8229), .A2(n8228), .ZN(n8250) );
  AOI21_X1 U9337 ( .B1(n8230), .B2(n10616), .A(n8250), .ZN(n10642) );
  XNOR2_X1 U9338 ( .A(n10607), .B(n10640), .ZN(n8231) );
  NOR2_X1 U9339 ( .A1(n8231), .A2(n10673), .ZN(n10639) );
  INV_X1 U9340 ( .A(n10640), .ZN(n8256) );
  AOI22_X1 U9341 ( .A1(n9157), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n8253), .B2(
        n10629), .ZN(n8232) );
  OAI21_X1 U9342 ( .B1(n10634), .B2(n8256), .A(n8232), .ZN(n8240) );
  NAND2_X1 U9343 ( .A1(n10612), .A2(n10595), .ZN(n8233) );
  NAND2_X1 U9344 ( .A1(n8938), .A2(n10606), .ZN(n8235) );
  NAND2_X1 U9345 ( .A1(n10604), .A2(n8235), .ZN(n8238) );
  INV_X1 U9346 ( .A(n8236), .ZN(n8237) );
  NAND2_X1 U9347 ( .A1(n8238), .A2(n8237), .ZN(n8282) );
  OAI21_X1 U9348 ( .B1(n8238), .B2(n8237), .A(n8282), .ZN(n10643) );
  NOR2_X1 U9349 ( .A1(n10643), .A2(n9255), .ZN(n8239) );
  AOI211_X1 U9350 ( .C1(n9266), .C2(n10639), .A(n8240), .B(n8239), .ZN(n8241)
         );
  OAI21_X1 U9351 ( .B1(n9157), .B2(n10642), .A(n8241), .ZN(P2_U3285) );
  OAI222_X1 U9352 ( .A1(n9387), .A2(n8244), .B1(P2_U3152), .B2(n6849), .C1(
        n8243), .C2(n8242), .ZN(P2_U3338) );
  AOI21_X1 U9353 ( .B1(n8845), .B2(n5147), .A(n8927), .ZN(n8249) );
  NOR3_X1 U9354 ( .A1(n8902), .A2(n8247), .A3(n8246), .ZN(n8248) );
  OAI21_X1 U9355 ( .B1(n8249), .B2(n8248), .A(n8400), .ZN(n8255) );
  INV_X1 U9356 ( .A(n8250), .ZN(n8251) );
  OAI22_X1 U9357 ( .A1(n8251), .A2(n8871), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9767), .ZN(n8252) );
  AOI21_X1 U9358 ( .B1(n8253), .B2(n8910), .A(n8252), .ZN(n8254) );
  OAI211_X1 U9359 ( .C1(n8256), .C2(n8922), .A(n8255), .B(n8254), .ZN(P2_U3238) );
  NAND2_X1 U9360 ( .A1(n8258), .A2(n8257), .ZN(n8259) );
  NAND2_X1 U9361 ( .A1(n8260), .A2(n8259), .ZN(n8266) );
  NAND2_X1 U9362 ( .A1(n8276), .A2(n8718), .ZN(n8262) );
  OR2_X1 U9363 ( .A1(n8267), .A2(n8701), .ZN(n8261) );
  NAND2_X1 U9364 ( .A1(n8262), .A2(n8261), .ZN(n8263) );
  XNOR2_X1 U9365 ( .A(n8263), .B(n7496), .ZN(n8264) );
  INV_X1 U9366 ( .A(n8264), .ZN(n8265) );
  NAND2_X1 U9367 ( .A1(n8324), .A2(n5244), .ZN(n8269) );
  NOR2_X1 U9368 ( .A1(n8267), .A2(n8713), .ZN(n8268) );
  AOI21_X1 U9369 ( .B1(n8276), .B2(n8721), .A(n8268), .ZN(n8323) );
  XNOR2_X1 U9370 ( .A(n8269), .B(n8323), .ZN(n8278) );
  INV_X1 U9371 ( .A(n8270), .ZN(n8274) );
  NAND2_X1 U9372 ( .A1(P1_U3084), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n10305) );
  INV_X1 U9373 ( .A(n10305), .ZN(n8271) );
  AOI21_X1 U9374 ( .B1(n9558), .B2(n10538), .A(n8271), .ZN(n8273) );
  NAND2_X1 U9375 ( .A1(n9788), .A2(n9545), .ZN(n8272) );
  OAI211_X1 U9376 ( .C1(n9516), .C2(n8274), .A(n8273), .B(n8272), .ZN(n8275)
         );
  AOI21_X1 U9377 ( .B1(n8276), .B2(n9564), .A(n8275), .ZN(n8277) );
  OAI21_X1 U9378 ( .B1(n8278), .B2(n9566), .A(n8277), .ZN(P1_U3215) );
  XNOR2_X1 U9379 ( .A(n8279), .B(n8283), .ZN(n8280) );
  OAI222_X1 U9380 ( .A1(n10611), .A2(n10614), .B1(n10613), .B2(n8504), .C1(
        n10436), .C2(n8280), .ZN(n10649) );
  INV_X1 U9381 ( .A(n10649), .ZN(n8292) );
  INV_X1 U9382 ( .A(n10614), .ZN(n8937) );
  NAND2_X1 U9383 ( .A1(n10640), .A2(n8937), .ZN(n8281) );
  OAI21_X1 U9384 ( .B1(n8285), .B2(n8284), .A(n8376), .ZN(n10651) );
  INV_X1 U9385 ( .A(n8411), .ZN(n10647) );
  NOR2_X1 U9386 ( .A1(n8286), .A2(n10647), .ZN(n8287) );
  OR2_X1 U9387 ( .A1(n8369), .A2(n8287), .ZN(n10648) );
  AOI22_X1 U9388 ( .A1(n9157), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n8404), .B2(
        n10629), .ZN(n8289) );
  NAND2_X1 U9389 ( .A1(n8411), .A2(n10451), .ZN(n8288) );
  OAI211_X1 U9390 ( .C1(n10648), .C2(n10454), .A(n8289), .B(n8288), .ZN(n8290)
         );
  AOI21_X1 U9391 ( .B1(n10651), .B2(n10456), .A(n8290), .ZN(n8291) );
  OAI21_X1 U9392 ( .B1(n8292), .B2(n10631), .A(n8291), .ZN(P2_U3284) );
  XNOR2_X1 U9393 ( .A(n8293), .B(n8295), .ZN(n8294) );
  AOI222_X1 U9394 ( .A1(n10546), .A2(n8294), .B1(n9404), .B2(n10539), .C1(
        n9788), .C2(n10540), .ZN(n10165) );
  OAI21_X1 U9395 ( .B1(n8297), .B2(n7106), .A(n8296), .ZN(n10166) );
  INV_X1 U9396 ( .A(n10166), .ZN(n8304) );
  INV_X1 U9397 ( .A(n10163), .ZN(n8302) );
  AOI21_X1 U9398 ( .B1(n8298), .B2(n10163), .A(n10582), .ZN(n8299) );
  AND2_X1 U9399 ( .A1(n8299), .A2(n8344), .ZN(n10162) );
  NAND2_X1 U9400 ( .A1(n10162), .A2(n10026), .ZN(n8301) );
  AOI22_X1 U9401 ( .A1(n9977), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n8359), .B2(
        n10561), .ZN(n8300) );
  OAI211_X1 U9402 ( .C1(n8302), .C2(n10565), .A(n8301), .B(n8300), .ZN(n8303)
         );
  AOI21_X1 U9403 ( .B1(n8304), .B2(n9911), .A(n8303), .ZN(n8305) );
  OAI21_X1 U9404 ( .B1(n9977), .B2(n10165), .A(n8305), .ZN(P1_U3279) );
  INV_X1 U9405 ( .A(n8306), .ZN(n8310) );
  OAI222_X1 U9406 ( .A1(n9387), .A2(n8308), .B1(n8243), .B2(n8310), .C1(n8307), 
        .C2(P2_U3152), .ZN(P2_U3336) );
  OAI222_X1 U9407 ( .A1(n8311), .A2(P1_U3084), .B1(n8826), .B2(n8310), .C1(
        n8309), .C2(n10209), .ZN(P1_U3331) );
  AOI22_X1 U9408 ( .A1(n8777), .A2(n8494), .B1(n8910), .B2(n8370), .ZN(n8314)
         );
  OAI211_X1 U9409 ( .C1(n8374), .C2(n8897), .A(n8314), .B(n8313), .ZN(n8315)
         );
  AOI21_X1 U9410 ( .B1(n8371), .B2(n8915), .A(n8315), .ZN(n8321) );
  INV_X1 U9411 ( .A(n8316), .ZN(n8319) );
  OAI22_X1 U9412 ( .A1(n8317), .A2(n8927), .B1(n8374), .B2(n8902), .ZN(n8318)
         );
  NAND3_X1 U9413 ( .A1(n8408), .A2(n8319), .A3(n8318), .ZN(n8320) );
  OAI211_X1 U9414 ( .C1(n8312), .C2(n8927), .A(n8321), .B(n8320), .ZN(P2_U3236) );
  NAND2_X1 U9415 ( .A1(n10168), .A2(n8718), .ZN(n8326) );
  OR2_X1 U9416 ( .A1(n8363), .A2(n8701), .ZN(n8325) );
  NAND2_X1 U9417 ( .A1(n8326), .A2(n8325), .ZN(n8327) );
  XNOR2_X1 U9418 ( .A(n8327), .B(n7496), .ZN(n8349) );
  NOR2_X1 U9419 ( .A1(n8363), .A2(n8713), .ZN(n8328) );
  AOI21_X1 U9420 ( .B1(n10168), .B2(n8721), .A(n8328), .ZN(n8350) );
  XNOR2_X1 U9421 ( .A(n8349), .B(n8350), .ZN(n8329) );
  OAI211_X1 U9422 ( .C1(n8330), .C2(n8329), .A(n8353), .B(n9536), .ZN(n8336)
         );
  AOI21_X1 U9423 ( .B1(n9789), .B2(n9558), .A(n8331), .ZN(n8332) );
  OAI21_X1 U9424 ( .B1(n8486), .B2(n9561), .A(n8332), .ZN(n8333) );
  AOI21_X1 U9425 ( .B1(n8334), .B2(n9556), .A(n8333), .ZN(n8335) );
  OAI211_X1 U9426 ( .C1(n8337), .C2(n9548), .A(n8336), .B(n8335), .ZN(P1_U3234) );
  XNOR2_X1 U9427 ( .A(n8339), .B(n8338), .ZN(n8340) );
  AOI222_X1 U9428 ( .A1(n10546), .A2(n8340), .B1(n9786), .B2(n10539), .C1(
        n9787), .C2(n10540), .ZN(n10160) );
  OAI21_X1 U9429 ( .B1(n8341), .B2(n8343), .A(n8342), .ZN(n10156) );
  AOI21_X1 U9430 ( .B1(n10157), .B2(n8344), .A(n8416), .ZN(n10158) );
  NAND2_X1 U9431 ( .A1(n10158), .A2(n10558), .ZN(n8346) );
  AOI22_X1 U9432 ( .A1(n9977), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n8488), .B2(
        n10561), .ZN(n8345) );
  OAI211_X1 U9433 ( .C1(n5012), .C2(n10565), .A(n8346), .B(n8345), .ZN(n8347)
         );
  AOI21_X1 U9434 ( .B1(n10156), .B2(n9911), .A(n8347), .ZN(n8348) );
  OAI21_X1 U9435 ( .B1(n9977), .B2(n10160), .A(n8348), .ZN(P1_U3278) );
  INV_X1 U9436 ( .A(n8349), .ZN(n8351) );
  OR2_X1 U9437 ( .A1(n8351), .A2(n8350), .ZN(n8352) );
  NAND2_X1 U9438 ( .A1(n10163), .A2(n8718), .ZN(n8355) );
  OR2_X1 U9439 ( .A1(n8486), .A2(n8701), .ZN(n8354) );
  NAND2_X1 U9440 ( .A1(n8355), .A2(n8354), .ZN(n8356) );
  XNOR2_X1 U9441 ( .A(n8356), .B(n8711), .ZN(n8465) );
  NOR2_X1 U9442 ( .A1(n8486), .A2(n8713), .ZN(n8357) );
  AOI21_X1 U9443 ( .B1(n10163), .B2(n8721), .A(n8357), .ZN(n8462) );
  INV_X1 U9444 ( .A(n8462), .ZN(n8466) );
  XNOR2_X1 U9445 ( .A(n8465), .B(n8466), .ZN(n8358) );
  XNOR2_X1 U9446 ( .A(n8464), .B(n8358), .ZN(n8366) );
  NAND2_X1 U9447 ( .A1(n9556), .A2(n8359), .ZN(n8362) );
  AOI21_X1 U9448 ( .B1(n9404), .B2(n9545), .A(n8360), .ZN(n8361) );
  OAI211_X1 U9449 ( .C1(n8363), .C2(n9542), .A(n8362), .B(n8361), .ZN(n8364)
         );
  AOI21_X1 U9450 ( .B1(n10163), .B2(n9564), .A(n8364), .ZN(n8365) );
  OAI21_X1 U9451 ( .B1(n8366), .B2(n9566), .A(n8365), .ZN(P1_U3222) );
  XNOR2_X1 U9452 ( .A(n8367), .B(n8377), .ZN(n8368) );
  OAI222_X1 U9453 ( .A1(n10611), .A2(n8374), .B1(n10613), .B2(n8783), .C1(
        n8368), .C2(n10436), .ZN(n10656) );
  OAI21_X1 U9454 ( .B1(n8369), .B2(n10654), .A(n8508), .ZN(n10655) );
  AOI22_X1 U9455 ( .A1(n10631), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n8370), .B2(
        n10629), .ZN(n8373) );
  NAND2_X1 U9456 ( .A1(n8371), .A2(n10451), .ZN(n8372) );
  OAI211_X1 U9457 ( .C1(n10655), .C2(n10454), .A(n8373), .B(n8372), .ZN(n8381)
         );
  INV_X1 U9458 ( .A(n8374), .ZN(n8936) );
  OR2_X1 U9459 ( .A1(n8411), .A2(n8936), .ZN(n8375) );
  NOR2_X1 U9460 ( .A1(n8378), .A2(n8377), .ZN(n10653) );
  INV_X1 U9461 ( .A(n8492), .ZN(n8379) );
  NOR3_X1 U9462 ( .A1(n10653), .A2(n8379), .A3(n9255), .ZN(n8380) );
  AOI211_X1 U9463 ( .C1(n10448), .C2(n10656), .A(n8381), .B(n8380), .ZN(n8382)
         );
  INV_X1 U9464 ( .A(n8382), .ZN(P2_U3283) );
  INV_X1 U9465 ( .A(n8396), .ZN(n8385) );
  NAND2_X1 U9466 ( .A1(n9378), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n8384) );
  OAI211_X1 U9467 ( .C1(n8385), .C2(n8243), .A(n8384), .B(n8383), .ZN(P2_U3335) );
  INV_X1 U9468 ( .A(n8505), .ZN(n8934) );
  AOI22_X1 U9469 ( .A1(n8777), .A2(n8934), .B1(n8910), .B2(n8509), .ZN(n8388)
         );
  OAI211_X1 U9470 ( .C1(n8504), .C2(n8897), .A(n8388), .B(n8387), .ZN(n8389)
         );
  AOI21_X1 U9471 ( .B1(n10661), .B2(n8915), .A(n8389), .ZN(n8395) );
  INV_X1 U9472 ( .A(n8390), .ZN(n8393) );
  OAI22_X1 U9473 ( .A1(n8391), .A2(n8927), .B1(n8504), .B2(n8902), .ZN(n8392)
         );
  NAND3_X1 U9474 ( .A1(n8312), .A2(n8393), .A3(n8392), .ZN(n8394) );
  OAI211_X1 U9475 ( .C1(n8386), .C2(n8927), .A(n8395), .B(n8394), .ZN(P2_U3217) );
  NAND2_X1 U9476 ( .A1(n8396), .A2(n10204), .ZN(n8398) );
  OAI211_X1 U9477 ( .C1(n8399), .C2(n10196), .A(n8398), .B(n8397), .ZN(
        P1_U3330) );
  INV_X1 U9478 ( .A(n8400), .ZN(n8403) );
  NOR3_X1 U9479 ( .A1(n8401), .A2(n10614), .A3(n8902), .ZN(n8402) );
  AOI21_X1 U9480 ( .B1(n8403), .B2(n8905), .A(n8402), .ZN(n8413) );
  INV_X1 U9481 ( .A(n8504), .ZN(n8935) );
  AOI22_X1 U9482 ( .A1(n8777), .A2(n8935), .B1(n8910), .B2(n8404), .ZN(n8407)
         );
  INV_X1 U9483 ( .A(n8405), .ZN(n8406) );
  OAI211_X1 U9484 ( .C1(n10614), .C2(n8897), .A(n8407), .B(n8406), .ZN(n8410)
         );
  NOR2_X1 U9485 ( .A1(n8408), .A2(n8927), .ZN(n8409) );
  AOI211_X1 U9486 ( .C1(n8411), .C2(n8915), .A(n8410), .B(n8409), .ZN(n8412)
         );
  OAI21_X1 U9487 ( .B1(n8414), .B2(n8413), .A(n8412), .ZN(P2_U3226) );
  XOR2_X1 U9488 ( .A(n8415), .B(n8419), .Z(n10155) );
  INV_X1 U9489 ( .A(n8416), .ZN(n8417) );
  AOI211_X1 U9490 ( .C1(n10152), .C2(n8417), .A(n10582), .B(n8528), .ZN(n10151) );
  AOI22_X1 U9491 ( .A1(n10563), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n9410), .B2(
        n10561), .ZN(n8418) );
  OAI21_X1 U9492 ( .B1(n9407), .B2(n10565), .A(n8418), .ZN(n8425) );
  AOI21_X1 U9493 ( .B1(n8420), .B2(n8419), .A(n7060), .ZN(n8423) );
  OAI22_X1 U9494 ( .A1(n8472), .A2(n7059), .B1(n9465), .B2(n10489), .ZN(n8421)
         );
  AOI21_X1 U9495 ( .B1(n8423), .B2(n8422), .A(n8421), .ZN(n10154) );
  NOR2_X1 U9496 ( .A1(n10154), .A2(n10563), .ZN(n8424) );
  AOI211_X1 U9497 ( .C1(n10026), .C2(n10151), .A(n8425), .B(n8424), .ZN(n8426)
         );
  OAI21_X1 U9498 ( .B1(n10155), .B2(n10028), .A(n8426), .ZN(P1_U3277) );
  AOI21_X1 U9499 ( .B1(n8428), .B2(n10670), .A(n8427), .ZN(n8429) );
  NAND2_X1 U9500 ( .A1(n8978), .A2(n8429), .ZN(n8430) );
  XNOR2_X1 U9501 ( .A(n8429), .B(n8437), .ZN(n8972) );
  NAND2_X1 U9502 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n8972), .ZN(n8971) );
  NAND2_X1 U9503 ( .A1(n8430), .A2(n8971), .ZN(n8432) );
  XNOR2_X1 U9504 ( .A(n8989), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n8431) );
  NOR2_X1 U9505 ( .A1(n8432), .A2(n8431), .ZN(n8990) );
  AOI21_X1 U9506 ( .B1(n8432), .B2(n8431), .A(n8990), .ZN(n8446) );
  NOR2_X1 U9507 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6449), .ZN(n8433) );
  AOI21_X1 U9508 ( .B1(n10314), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n8433), .ZN(
        n8434) );
  INV_X1 U9509 ( .A(n8434), .ZN(n8444) );
  OAI21_X1 U9510 ( .B1(n8436), .B2(P2_REG2_REG_14__SCAN_IN), .A(n8435), .ZN(
        n8438) );
  NAND2_X1 U9511 ( .A1(n8437), .A2(n8438), .ZN(n8439) );
  XNOR2_X1 U9512 ( .A(n8438), .B(n8978), .ZN(n8975) );
  NAND2_X1 U9513 ( .A1(n8975), .A2(n6440), .ZN(n8974) );
  NAND2_X1 U9514 ( .A1(n8439), .A2(n8974), .ZN(n8442) );
  NAND2_X1 U9515 ( .A1(n8989), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n8440) );
  OAI21_X1 U9516 ( .B1(n8989), .B2(P2_REG2_REG_16__SCAN_IN), .A(n8440), .ZN(
        n8441) );
  NOR2_X1 U9517 ( .A1(n8442), .A2(n8441), .ZN(n8983) );
  AOI211_X1 U9518 ( .C1(n8442), .C2(n8441), .A(n8983), .B(n10325), .ZN(n8443)
         );
  AOI211_X1 U9519 ( .C1(n10320), .C2(n8989), .A(n8444), .B(n8443), .ZN(n8445)
         );
  OAI21_X1 U9520 ( .B1(n8446), .B2(n10329), .A(n8445), .ZN(P2_U3261) );
  INV_X1 U9521 ( .A(n8447), .ZN(n8451) );
  INV_X1 U9522 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n8448) );
  OAI222_X1 U9523 ( .A1(P2_U3152), .A2(n8449), .B1(n8243), .B2(n8451), .C1(
        n8448), .C2(n9387), .ZN(P2_U3334) );
  OAI222_X1 U9524 ( .A1(n8452), .A2(P1_U3084), .B1(n8826), .B2(n8451), .C1(
        n8450), .C2(n10209), .ZN(P1_U3329) );
  INV_X1 U9525 ( .A(n8545), .ZN(n8454) );
  OAI22_X1 U9526 ( .A1(n9249), .A2(n10613), .B1(n8505), .B2(n10611), .ZN(n8536) );
  AOI22_X1 U9527 ( .A1(n8536), .A2(n8925), .B1(P2_REG3_REG_16__SCAN_IN), .B2(
        P2_U3152), .ZN(n8453) );
  OAI21_X1 U9528 ( .B1(n8454), .B2(n8921), .A(n8453), .ZN(n8455) );
  AOI21_X1 U9529 ( .B1(n9349), .B2(n8915), .A(n8455), .ZN(n8460) );
  OAI22_X1 U9530 ( .A1(n8457), .A2(n8927), .B1(n8505), .B2(n8902), .ZN(n8458)
         );
  NAND3_X1 U9531 ( .A1(n8789), .A2(n4946), .A3(n8458), .ZN(n8459) );
  OAI211_X1 U9532 ( .C1(n8461), .C2(n8927), .A(n8460), .B(n8459), .ZN(P2_U3228) );
  NAND2_X1 U9533 ( .A1(n8465), .A2(n8462), .ZN(n8463) );
  INV_X1 U9534 ( .A(n8465), .ZN(n8467) );
  NAND2_X1 U9535 ( .A1(n8467), .A2(n8466), .ZN(n8468) );
  NAND2_X1 U9536 ( .A1(n10157), .A2(n8718), .ZN(n8470) );
  OR2_X1 U9537 ( .A1(n8472), .A2(n8701), .ZN(n8469) );
  NAND2_X1 U9538 ( .A1(n8470), .A2(n8469), .ZN(n8471) );
  XNOR2_X1 U9539 ( .A(n8471), .B(n7496), .ZN(n8476) );
  NAND2_X1 U9540 ( .A1(n10157), .A2(n8721), .ZN(n8474) );
  OR2_X1 U9541 ( .A1(n8472), .A2(n8713), .ZN(n8473) );
  NAND2_X1 U9542 ( .A1(n8474), .A2(n8473), .ZN(n8477) );
  AND2_X1 U9543 ( .A1(n8476), .A2(n8477), .ZN(n8481) );
  INV_X1 U9544 ( .A(n8481), .ZN(n8475) );
  INV_X1 U9545 ( .A(n8476), .ZN(n8479) );
  INV_X1 U9546 ( .A(n8477), .ZN(n8478) );
  NAND2_X1 U9547 ( .A1(n8479), .A2(n8478), .ZN(n8609) );
  OAI21_X1 U9548 ( .B1(n5207), .B2(n8481), .A(n8480), .ZN(n8482) );
  OAI21_X1 U9549 ( .B1(n8610), .B2(n5207), .A(n8482), .ZN(n8483) );
  NAND2_X1 U9550 ( .A1(n8483), .A2(n9536), .ZN(n8490) );
  AOI21_X1 U9551 ( .B1(n9545), .B2(n9786), .A(n8484), .ZN(n8485) );
  OAI21_X1 U9552 ( .B1(n8486), .B2(n9542), .A(n8485), .ZN(n8487) );
  AOI21_X1 U9553 ( .B1(n8488), .B2(n9556), .A(n8487), .ZN(n8489) );
  OAI211_X1 U9554 ( .C1(n5012), .C2(n9548), .A(n8490), .B(n8489), .ZN(P1_U3232) );
  NAND2_X1 U9555 ( .A1(n8371), .A2(n8935), .ZN(n8491) );
  NAND2_X1 U9556 ( .A1(n8492), .A2(n8491), .ZN(n8513) );
  INV_X1 U9557 ( .A(n10661), .ZN(n8511) );
  NOR2_X1 U9558 ( .A1(n10661), .A2(n8494), .ZN(n8495) );
  NOR2_X1 U9559 ( .A1(n8512), .A2(n8495), .ZN(n8539) );
  XNOR2_X1 U9560 ( .A(n8539), .B(n8538), .ZN(n10678) );
  INV_X1 U9561 ( .A(n10678), .ZN(n8502) );
  XNOR2_X1 U9562 ( .A(n8496), .B(n8538), .ZN(n8497) );
  OAI222_X1 U9563 ( .A1(n10613), .A2(n8775), .B1(n10611), .B2(n8783), .C1(
        n10436), .C2(n8497), .ZN(n10675) );
  OAI21_X1 U9564 ( .B1(n4917), .B2(n5164), .A(n8542), .ZN(n10674) );
  AOI22_X1 U9565 ( .A1(n10631), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n8776), .B2(
        n10629), .ZN(n8499) );
  NAND2_X1 U9566 ( .A1(n8781), .A2(n10451), .ZN(n8498) );
  OAI211_X1 U9567 ( .C1(n10674), .C2(n10454), .A(n8499), .B(n8498), .ZN(n8500)
         );
  AOI21_X1 U9568 ( .B1(n10675), .B2(n10448), .A(n8500), .ZN(n8501) );
  OAI21_X1 U9569 ( .B1(n8502), .B2(n9255), .A(n8501), .ZN(P2_U3281) );
  XNOR2_X1 U9570 ( .A(n8503), .B(n6430), .ZN(n8507) );
  OAI22_X1 U9571 ( .A1(n8505), .A2(n10613), .B1(n8504), .B2(n10611), .ZN(n8506) );
  AOI21_X1 U9572 ( .B1(n8507), .B2(n10616), .A(n8506), .ZN(n10666) );
  XNOR2_X1 U9573 ( .A(n8508), .B(n8511), .ZN(n10664) );
  AOI22_X1 U9574 ( .A1(n10631), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n8509), .B2(
        n10629), .ZN(n8510) );
  OAI21_X1 U9575 ( .B1(n8511), .B2(n10634), .A(n8510), .ZN(n8515) );
  AOI21_X1 U9576 ( .B1(n6430), .B2(n8513), .A(n8512), .ZN(n10668) );
  NOR2_X1 U9577 ( .A1(n10668), .A2(n9255), .ZN(n8514) );
  AOI211_X1 U9578 ( .C1(n10626), .C2(n10664), .A(n8515), .B(n8514), .ZN(n8516)
         );
  OAI21_X1 U9579 ( .B1(n9157), .B2(n10666), .A(n8516), .ZN(P2_U3282) );
  NAND2_X1 U9580 ( .A1(n8517), .A2(n8518), .ZN(n8519) );
  NAND2_X1 U9581 ( .A1(n8521), .A2(n8522), .ZN(n8523) );
  AOI21_X1 U9582 ( .B1(n8524), .B2(n8523), .A(n7060), .ZN(n8527) );
  OAI22_X1 U9583 ( .A1(n8525), .A2(n7059), .B1(n9562), .B2(n10489), .ZN(n8526)
         );
  AOI211_X1 U9584 ( .C1(n10145), .C2(n10522), .A(n8527), .B(n8526), .ZN(n10149) );
  OR2_X1 U9585 ( .A1(n8528), .A2(n8532), .ZN(n8529) );
  AND2_X1 U9586 ( .A1(n4916), .A2(n8529), .ZN(n10147) );
  NAND2_X1 U9587 ( .A1(n10147), .A2(n10558), .ZN(n8531) );
  AOI22_X1 U9588 ( .A1(n10563), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n9555), .B2(
        n10561), .ZN(n8530) );
  OAI211_X1 U9589 ( .C1(n8532), .C2(n10565), .A(n8531), .B(n8530), .ZN(n8533)
         );
  AOI21_X1 U9590 ( .B1(n10145), .B2(n10559), .A(n8533), .ZN(n8534) );
  OAI21_X1 U9591 ( .B1(n10149), .B2(n9977), .A(n8534), .ZN(P1_U3276) );
  XOR2_X1 U9592 ( .A(n8535), .B(n8541), .Z(n8537) );
  AOI21_X1 U9593 ( .B1(n8537), .B2(n10616), .A(n8536), .ZN(n9351) );
  OAI22_X1 U9594 ( .A1(n8539), .A2(n8538), .B1(n8934), .B2(n8781), .ZN(n8540)
         );
  AOI21_X1 U9595 ( .B1(n8541), .B2(n8540), .A(n9044), .ZN(n9347) );
  NAND2_X1 U9596 ( .A1(n8542), .A2(n9349), .ZN(n8543) );
  NAND2_X1 U9597 ( .A1(n8543), .A2(n10663), .ZN(n8544) );
  NOR2_X1 U9598 ( .A1(n9264), .A2(n8544), .ZN(n9348) );
  NAND2_X1 U9599 ( .A1(n9348), .A2(n9266), .ZN(n8547) );
  AOI22_X1 U9600 ( .A1(n10631), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n8545), .B2(
        n10629), .ZN(n8546) );
  OAI211_X1 U9601 ( .C1(n5162), .C2(n10634), .A(n8547), .B(n8546), .ZN(n8548)
         );
  AOI21_X1 U9602 ( .B1(n9347), .B2(n10456), .A(n8548), .ZN(n8549) );
  OAI21_X1 U9603 ( .B1(n9157), .B2(n9351), .A(n8549), .ZN(P2_U3280) );
  XNOR2_X1 U9604 ( .A(n8551), .B(n8550), .ZN(n8553) );
  AOI222_X1 U9605 ( .A1(n10546), .A2(n8553), .B1(n9573), .B2(n10539), .C1(
        n8552), .C2(n10540), .ZN(n10143) );
  OAI21_X1 U9606 ( .B1(n8554), .B2(n8556), .A(n8555), .ZN(n10144) );
  INV_X1 U9607 ( .A(n10144), .ZN(n8563) );
  INV_X1 U9608 ( .A(n10141), .ZN(n8561) );
  AOI21_X1 U9609 ( .B1(n4916), .B2(n10141), .A(n10582), .ZN(n8558) );
  INV_X1 U9610 ( .A(n8557), .ZN(n10059) );
  AND2_X1 U9611 ( .A1(n8558), .A2(n10059), .ZN(n10140) );
  NAND2_X1 U9612 ( .A1(n10140), .A2(n10026), .ZN(n8560) );
  AOI22_X1 U9613 ( .A1(n10563), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9462), .B2(
        n10561), .ZN(n8559) );
  OAI211_X1 U9614 ( .C1(n8561), .C2(n10565), .A(n8560), .B(n8559), .ZN(n8562)
         );
  AOI21_X1 U9615 ( .B1(n8563), .B2(n9911), .A(n8562), .ZN(n8564) );
  OAI21_X1 U9616 ( .B1(n9977), .B2(n10143), .A(n8564), .ZN(P1_U3275) );
  NAND2_X1 U9617 ( .A1(n6926), .A2(n8566), .ZN(n8567) );
  XNOR2_X1 U9618 ( .A(n8568), .B(n8567), .ZN(n8573) );
  INV_X1 U9619 ( .A(n9267), .ZN(n8570) );
  OAI22_X1 U9620 ( .A1(n9047), .A2(n10613), .B1(n8775), .B2(n10611), .ZN(n9260) );
  AOI22_X1 U9621 ( .A1(n9260), .A2(n8925), .B1(P2_REG3_REG_17__SCAN_IN), .B2(
        n4846), .ZN(n8569) );
  OAI21_X1 U9622 ( .B1(n8570), .B2(n8921), .A(n8569), .ZN(n8571) );
  AOI21_X1 U9623 ( .B1(n9343), .B2(n8915), .A(n8571), .ZN(n8572) );
  OAI21_X1 U9624 ( .B1(n8573), .B2(n8927), .A(n8572), .ZN(P2_U3230) );
  INV_X1 U9625 ( .A(n8574), .ZN(n8577) );
  OAI222_X1 U9626 ( .A1(P1_U3084), .A2(n5026), .B1(n8826), .B2(n8577), .C1(
        n8575), .C2(n10196), .ZN(P1_U3328) );
  OAI222_X1 U9627 ( .A1(n9387), .A2(n8578), .B1(n8243), .B2(n8577), .C1(n4846), 
        .C2(n8576), .ZN(P2_U3333) );
  INV_X1 U9628 ( .A(n8579), .ZN(n8583) );
  OAI222_X1 U9629 ( .A1(n4846), .A2(n8581), .B1(n8243), .B2(n8583), .C1(n8580), 
        .C2(n9387), .ZN(P2_U3332) );
  OAI222_X1 U9630 ( .A1(n7066), .A2(P1_U3084), .B1(n8826), .B2(n8583), .C1(
        n8582), .C2(n10196), .ZN(P1_U3327) );
  OAI21_X1 U9631 ( .B1(n8586), .B2(n8585), .A(n8809), .ZN(n8587) );
  OAI22_X1 U9632 ( .A1(n9898), .A2(n10489), .B1(n9543), .B2(n7059), .ZN(n8588)
         );
  INV_X1 U9633 ( .A(n8588), .ZN(n8589) );
  INV_X1 U9634 ( .A(n9916), .ZN(n8593) );
  NAND2_X1 U9635 ( .A1(n8593), .A2(n10086), .ZN(n8594) );
  AND2_X1 U9636 ( .A1(n8595), .A2(n8594), .ZN(n10087) );
  INV_X1 U9637 ( .A(n8596), .ZN(n9540) );
  AOI22_X1 U9638 ( .A1(n9540), .A2(n10561), .B1(P1_REG2_REG_26__SCAN_IN), .B2(
        n10563), .ZN(n8597) );
  OAI21_X1 U9639 ( .B1(n9549), .B2(n10565), .A(n8597), .ZN(n8600) );
  NOR2_X1 U9640 ( .A1(n10090), .A2(n8598), .ZN(n8599) );
  AOI211_X1 U9641 ( .C1(n10558), .C2(n10087), .A(n8600), .B(n8599), .ZN(n8601)
         );
  OAI21_X1 U9642 ( .B1(n10089), .B2(n9977), .A(n8601), .ZN(P1_U3265) );
  INV_X1 U9643 ( .A(n9289), .ZN(n9097) );
  INV_X1 U9644 ( .A(n9343), .ZN(n9270) );
  NAND2_X1 U9645 ( .A1(n9264), .A2(n9270), .ZN(n9241) );
  INV_X1 U9646 ( .A(n9326), .ZN(n9210) );
  XOR2_X1 U9647 ( .A(n6781), .B(n9038), .Z(n9274) );
  INV_X1 U9648 ( .A(n9385), .ZN(n8604) );
  NAND2_X1 U9649 ( .A1(n8604), .A2(P2_B_REG_SCAN_IN), .ZN(n8605) );
  NAND2_X1 U9650 ( .A1(n9178), .A2(n8605), .ZN(n9068) );
  INV_X1 U9651 ( .A(n9068), .ZN(n8606) );
  NAND2_X1 U9652 ( .A1(n8929), .A2(n8606), .ZN(n9277) );
  NOR2_X1 U9653 ( .A1(n9157), .A2(n9277), .ZN(n9040) );
  AOI21_X1 U9654 ( .B1(n9157), .B2(P2_REG2_REG_31__SCAN_IN), .A(n9040), .ZN(
        n8608) );
  NAND2_X1 U9655 ( .A1(n6781), .A2(n10451), .ZN(n8607) );
  OAI211_X1 U9656 ( .C1(n9274), .C2(n10454), .A(n8608), .B(n8607), .ZN(
        P2_U3265) );
  NAND2_X1 U9657 ( .A1(n10152), .A2(n8718), .ZN(n8612) );
  NAND2_X1 U9658 ( .A1(n9786), .A2(n8721), .ZN(n8611) );
  NAND2_X1 U9659 ( .A1(n8612), .A2(n8611), .ZN(n8613) );
  XNOR2_X1 U9660 ( .A(n8613), .B(n8711), .ZN(n8616) );
  NAND2_X1 U9661 ( .A1(n10152), .A2(n8721), .ZN(n8615) );
  NAND2_X1 U9662 ( .A1(n9786), .A2(n8720), .ZN(n8614) );
  NAND2_X1 U9663 ( .A1(n8615), .A2(n8614), .ZN(n9403) );
  NAND2_X1 U9664 ( .A1(n10141), .A2(n8718), .ZN(n8618) );
  OR2_X1 U9665 ( .A1(n9562), .A2(n8701), .ZN(n8617) );
  NAND2_X1 U9666 ( .A1(n8618), .A2(n8617), .ZN(n8619) );
  XNOR2_X1 U9667 ( .A(n8619), .B(n8711), .ZN(n9459) );
  NOR2_X1 U9668 ( .A1(n9562), .A2(n8713), .ZN(n8620) );
  AOI21_X1 U9669 ( .B1(n10141), .B2(n8721), .A(n8620), .ZN(n8627) );
  NOR2_X1 U9670 ( .A1(n9465), .A2(n8713), .ZN(n8621) );
  AOI21_X1 U9671 ( .B1(n10146), .B2(n8721), .A(n8621), .ZN(n9553) );
  NAND2_X1 U9672 ( .A1(n10146), .A2(n8718), .ZN(n8623) );
  OR2_X1 U9673 ( .A1(n9465), .A2(n8701), .ZN(n8622) );
  NAND2_X1 U9674 ( .A1(n8623), .A2(n8622), .ZN(n8624) );
  XNOR2_X1 U9675 ( .A(n8624), .B(n8711), .ZN(n9456) );
  OAI22_X1 U9676 ( .A1(n9459), .A2(n8627), .B1(n9553), .B2(n9456), .ZN(n8630)
         );
  NAND2_X1 U9677 ( .A1(n9456), .A2(n9553), .ZN(n8625) );
  INV_X1 U9678 ( .A(n8627), .ZN(n9458) );
  NAND2_X1 U9679 ( .A1(n8625), .A2(n9458), .ZN(n8628) );
  INV_X1 U9680 ( .A(n8625), .ZN(n8626) );
  AOI22_X1 U9681 ( .A1(n9459), .A2(n8628), .B1(n8627), .B2(n8626), .ZN(n8629)
         );
  NAND2_X1 U9682 ( .A1(n10135), .A2(n8718), .ZN(n8632) );
  NAND2_X1 U9683 ( .A1(n9573), .A2(n8721), .ZN(n8631) );
  NAND2_X1 U9684 ( .A1(n8632), .A2(n8631), .ZN(n8633) );
  XNOR2_X1 U9685 ( .A(n8633), .B(n8711), .ZN(n9471) );
  AND2_X1 U9686 ( .A1(n9573), .A2(n8720), .ZN(n8634) );
  AOI21_X1 U9687 ( .B1(n10135), .B2(n8721), .A(n8634), .ZN(n9470) );
  AND2_X1 U9688 ( .A1(n9471), .A2(n9470), .ZN(n8635) );
  NAND2_X1 U9689 ( .A1(n10043), .A2(n8721), .ZN(n8637) );
  OR2_X1 U9690 ( .A1(n9474), .A2(n8713), .ZN(n8636) );
  NAND2_X1 U9691 ( .A1(n8637), .A2(n8636), .ZN(n9528) );
  NAND2_X1 U9692 ( .A1(n10043), .A2(n8718), .ZN(n8639) );
  OR2_X1 U9693 ( .A1(n9474), .A2(n8701), .ZN(n8638) );
  NAND2_X1 U9694 ( .A1(n8639), .A2(n8638), .ZN(n8640) );
  XNOR2_X1 U9695 ( .A(n8640), .B(n7496), .ZN(n9527) );
  NAND2_X1 U9696 ( .A1(n10123), .A2(n8718), .ZN(n8642) );
  NAND2_X1 U9697 ( .A1(n9572), .A2(n8721), .ZN(n8641) );
  NAND2_X1 U9698 ( .A1(n8642), .A2(n8641), .ZN(n8643) );
  XNOR2_X1 U9699 ( .A(n8643), .B(n8711), .ZN(n8645) );
  AND2_X1 U9700 ( .A1(n9572), .A2(n8720), .ZN(n8644) );
  AOI21_X1 U9701 ( .B1(n10123), .B2(n8721), .A(n8644), .ZN(n8646) );
  NAND2_X1 U9702 ( .A1(n8645), .A2(n8646), .ZN(n8650) );
  INV_X1 U9703 ( .A(n8645), .ZN(n8648) );
  INV_X1 U9704 ( .A(n8646), .ZN(n8647) );
  NAND2_X1 U9705 ( .A1(n8648), .A2(n8647), .ZN(n8649) );
  NAND2_X1 U9706 ( .A1(n8650), .A2(n8649), .ZN(n9424) );
  NAND2_X1 U9707 ( .A1(n10117), .A2(n8718), .ZN(n8652) );
  NAND2_X1 U9708 ( .A1(n10022), .A2(n8721), .ZN(n8651) );
  NAND2_X1 U9709 ( .A1(n8652), .A2(n8651), .ZN(n8653) );
  XNOR2_X1 U9710 ( .A(n8653), .B(n8711), .ZN(n8656) );
  AND2_X1 U9711 ( .A1(n10022), .A2(n8720), .ZN(n8654) );
  AOI21_X1 U9712 ( .B1(n10117), .B2(n8721), .A(n8654), .ZN(n8657) );
  AND2_X1 U9713 ( .A1(n8656), .A2(n8657), .ZN(n9502) );
  INV_X1 U9714 ( .A(n9502), .ZN(n8655) );
  INV_X1 U9715 ( .A(n8656), .ZN(n8659) );
  INV_X1 U9716 ( .A(n8657), .ZN(n8658) );
  NAND2_X1 U9717 ( .A1(n8659), .A2(n8658), .ZN(n9503) );
  NAND2_X1 U9718 ( .A1(n10113), .A2(n8718), .ZN(n8661) );
  NAND2_X1 U9719 ( .A1(n9970), .A2(n8721), .ZN(n8660) );
  NAND2_X1 U9720 ( .A1(n8661), .A2(n8660), .ZN(n8662) );
  XNOR2_X1 U9721 ( .A(n8662), .B(n7496), .ZN(n8665) );
  NAND2_X1 U9722 ( .A1(n10113), .A2(n8721), .ZN(n8664) );
  NAND2_X1 U9723 ( .A1(n9970), .A2(n8720), .ZN(n8663) );
  NAND2_X1 U9724 ( .A1(n8664), .A2(n8663), .ZN(n8666) );
  AND2_X1 U9725 ( .A1(n8665), .A2(n8666), .ZN(n9431) );
  INV_X1 U9726 ( .A(n8665), .ZN(n8668) );
  INV_X1 U9727 ( .A(n8666), .ZN(n8667) );
  NAND2_X1 U9728 ( .A1(n8668), .A2(n8667), .ZN(n9430) );
  NAND2_X1 U9729 ( .A1(n10106), .A2(n8718), .ZN(n8670) );
  NAND2_X1 U9730 ( .A1(n9955), .A2(n8721), .ZN(n8669) );
  NAND2_X1 U9731 ( .A1(n8670), .A2(n8669), .ZN(n8671) );
  XNOR2_X1 U9732 ( .A(n8671), .B(n7496), .ZN(n8673) );
  AND2_X1 U9733 ( .A1(n9955), .A2(n8720), .ZN(n8672) );
  AOI21_X1 U9734 ( .B1(n10106), .B2(n8721), .A(n8672), .ZN(n8674) );
  XNOR2_X1 U9735 ( .A(n8673), .B(n8674), .ZN(n9512) );
  INV_X1 U9736 ( .A(n8673), .ZN(n8675) );
  NAND2_X1 U9737 ( .A1(n8675), .A2(n8674), .ZN(n8676) );
  NAND2_X1 U9738 ( .A1(n8677), .A2(n8676), .ZN(n8682) );
  NAND2_X1 U9739 ( .A1(n10102), .A2(n8718), .ZN(n8679) );
  NAND2_X1 U9740 ( .A1(n9969), .A2(n8721), .ZN(n8678) );
  NAND2_X1 U9741 ( .A1(n8679), .A2(n8678), .ZN(n8680) );
  XNOR2_X1 U9742 ( .A(n8680), .B(n8711), .ZN(n8683) );
  INV_X1 U9743 ( .A(n10102), .ZN(n9951) );
  OAI22_X1 U9744 ( .A1(n9951), .A2(n8701), .B1(n8681), .B2(n8713), .ZN(n9415)
         );
  INV_X1 U9745 ( .A(n8682), .ZN(n8685) );
  INV_X1 U9746 ( .A(n8683), .ZN(n8684) );
  NAND2_X1 U9747 ( .A1(n10097), .A2(n8718), .ZN(n8687) );
  NAND2_X1 U9748 ( .A1(n9954), .A2(n8721), .ZN(n8686) );
  NAND2_X1 U9749 ( .A1(n8687), .A2(n8686), .ZN(n8688) );
  XNOR2_X1 U9750 ( .A(n8688), .B(n7496), .ZN(n8692) );
  NOR2_X1 U9751 ( .A1(n9448), .A2(n8713), .ZN(n8689) );
  AOI21_X1 U9752 ( .B1(n10097), .B2(n8721), .A(n8689), .ZN(n8690) );
  XNOR2_X1 U9753 ( .A(n8692), .B(n8690), .ZN(n9480) );
  INV_X1 U9754 ( .A(n8690), .ZN(n8691) );
  NAND2_X1 U9755 ( .A1(n10092), .A2(n8718), .ZN(n8695) );
  NAND2_X1 U9756 ( .A1(n9930), .A2(n8721), .ZN(n8694) );
  NAND2_X1 U9757 ( .A1(n8695), .A2(n8694), .ZN(n8696) );
  XNOR2_X1 U9758 ( .A(n8696), .B(n7496), .ZN(n8700) );
  NAND2_X1 U9759 ( .A1(n10092), .A2(n8721), .ZN(n8698) );
  NAND2_X1 U9760 ( .A1(n9930), .A2(n8720), .ZN(n8697) );
  NAND2_X1 U9761 ( .A1(n8698), .A2(n8697), .ZN(n8699) );
  NOR2_X1 U9762 ( .A1(n8700), .A2(n8699), .ZN(n9442) );
  NAND2_X1 U9763 ( .A1(n8700), .A2(n8699), .ZN(n9443) );
  OAI22_X1 U9764 ( .A1(n9549), .A2(n8702), .B1(n9451), .B2(n8701), .ZN(n8703)
         );
  XNOR2_X1 U9765 ( .A(n8703), .B(n7496), .ZN(n8705) );
  AND2_X1 U9766 ( .A1(n9923), .A2(n8720), .ZN(n8704) );
  AOI21_X1 U9767 ( .B1(n10086), .B2(n8721), .A(n8704), .ZN(n8706) );
  XNOR2_X1 U9768 ( .A(n8705), .B(n8706), .ZN(n9538) );
  INV_X1 U9769 ( .A(n8706), .ZN(n8707) );
  NAND2_X1 U9770 ( .A1(n10082), .A2(n8718), .ZN(n8710) );
  NAND2_X1 U9771 ( .A1(n9571), .A2(n8721), .ZN(n8709) );
  NAND2_X1 U9772 ( .A1(n8710), .A2(n8709), .ZN(n8712) );
  XNOR2_X1 U9773 ( .A(n8712), .B(n8711), .ZN(n9390) );
  NOR2_X1 U9774 ( .A1(n9898), .A2(n8713), .ZN(n8714) );
  AOI21_X1 U9775 ( .B1(n10082), .B2(n8721), .A(n8714), .ZN(n8715) );
  NAND2_X1 U9776 ( .A1(n9390), .A2(n8715), .ZN(n8717) );
  INV_X1 U9777 ( .A(n9390), .ZN(n8716) );
  INV_X1 U9778 ( .A(n8715), .ZN(n9389) );
  AOI22_X1 U9779 ( .A1(n10076), .A2(n8718), .B1(n8721), .B2(n9570), .ZN(n8719)
         );
  XNOR2_X1 U9780 ( .A(n8719), .B(n7496), .ZN(n8723) );
  AOI22_X1 U9781 ( .A1(n10076), .A2(n8721), .B1(n8720), .B2(n9570), .ZN(n8722)
         );
  OAI22_X1 U9782 ( .A1(n9903), .A2(n9516), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8724), .ZN(n8725) );
  AOI21_X1 U9783 ( .B1(n9571), .B2(n9558), .A(n8725), .ZN(n8726) );
  OAI21_X1 U9784 ( .B1(n9899), .B2(n9561), .A(n8726), .ZN(n8727) );
  AOI21_X1 U9785 ( .B1(n10076), .B2(n9564), .A(n8727), .ZN(n8728) );
  OAI21_X1 U9786 ( .B1(n8729), .B2(n9566), .A(n8728), .ZN(P1_U3218) );
  NOR2_X1 U9787 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n8770) );
  NOR2_X1 U9788 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n8768) );
  NOR2_X1 U9789 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n8766) );
  NOR2_X1 U9790 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n8764) );
  NOR2_X1 U9791 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n8761) );
  NOR2_X1 U9792 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n8758) );
  NAND2_X1 U9793 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n8755) );
  XOR2_X1 U9794 ( .A(P2_ADDR_REG_11__SCAN_IN), .B(P1_ADDR_REG_11__SCAN_IN), 
        .Z(n10238) );
  NAND2_X1 U9795 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n8753) );
  XOR2_X1 U9796 ( .A(P2_ADDR_REG_10__SCAN_IN), .B(P1_ADDR_REG_10__SCAN_IN), 
        .Z(n10236) );
  NOR2_X1 U9797 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n8737) );
  XOR2_X1 U9798 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(n8730), .Z(n10227) );
  NAND2_X1 U9799 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(P1_ADDR_REG_3__SCAN_IN), 
        .ZN(n8735) );
  XNOR2_X1 U9800 ( .A(n8731), .B(P1_ADDR_REG_3__SCAN_IN), .ZN(n10225) );
  NAND2_X1 U9801 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n8733) );
  XOR2_X1 U9802 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P2_ADDR_REG_2__SCAN_IN), .Z(
        n10223) );
  AOI21_X1 U9803 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10217) );
  INV_X1 U9804 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10221) );
  NAND3_X1 U9805 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_0__SCAN_IN), .ZN(n10219) );
  OAI21_X1 U9806 ( .B1(n10217), .B2(n10221), .A(n10219), .ZN(n10222) );
  NAND2_X1 U9807 ( .A1(n10223), .A2(n10222), .ZN(n8732) );
  NAND2_X1 U9808 ( .A1(n8733), .A2(n8732), .ZN(n10224) );
  NAND2_X1 U9809 ( .A1(n10225), .A2(n10224), .ZN(n8734) );
  NAND2_X1 U9810 ( .A1(n8735), .A2(n8734), .ZN(n10226) );
  NOR2_X1 U9811 ( .A1(n10227), .A2(n10226), .ZN(n8736) );
  NOR2_X1 U9812 ( .A1(n8737), .A2(n8736), .ZN(n8738) );
  NOR2_X1 U9813 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n8738), .ZN(n10228) );
  AND2_X1 U9814 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n8738), .ZN(n10229) );
  NOR2_X1 U9815 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n10229), .ZN(n8739) );
  NAND2_X1 U9816 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(n8740), .ZN(n8742) );
  XOR2_X1 U9817 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(n8740), .Z(n10231) );
  NAND2_X1 U9818 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(n10231), .ZN(n8741) );
  NAND2_X1 U9819 ( .A1(n8742), .A2(n8741), .ZN(n8743) );
  NAND2_X1 U9820 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n8743), .ZN(n8745) );
  XOR2_X1 U9821 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n8743), .Z(n10232) );
  NAND2_X1 U9822 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n10232), .ZN(n8744) );
  NAND2_X1 U9823 ( .A1(n8745), .A2(n8744), .ZN(n8746) );
  NAND2_X1 U9824 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n8746), .ZN(n8748) );
  XOR2_X1 U9825 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n8746), .Z(n10233) );
  NAND2_X1 U9826 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n10233), .ZN(n8747) );
  NAND2_X1 U9827 ( .A1(n8748), .A2(n8747), .ZN(n8749) );
  NAND2_X1 U9828 ( .A1(P1_ADDR_REG_9__SCAN_IN), .A2(n8749), .ZN(n8751) );
  XOR2_X1 U9829 ( .A(P1_ADDR_REG_9__SCAN_IN), .B(n8749), .Z(n10234) );
  NAND2_X1 U9830 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n10234), .ZN(n8750) );
  NAND2_X1 U9831 ( .A1(n8751), .A2(n8750), .ZN(n10235) );
  NAND2_X1 U9832 ( .A1(n10236), .A2(n10235), .ZN(n8752) );
  NAND2_X1 U9833 ( .A1(n8753), .A2(n8752), .ZN(n10237) );
  NAND2_X1 U9834 ( .A1(n10238), .A2(n10237), .ZN(n8754) );
  NAND2_X1 U9835 ( .A1(n8755), .A2(n8754), .ZN(n10240) );
  XOR2_X1 U9836 ( .A(P2_ADDR_REG_12__SCAN_IN), .B(n8756), .Z(n10239) );
  XOR2_X1 U9837 ( .A(n8759), .B(P1_ADDR_REG_13__SCAN_IN), .Z(n10241) );
  XOR2_X1 U9838 ( .A(n8762), .B(P1_ADDR_REG_14__SCAN_IN), .Z(n10243) );
  INV_X1 U9839 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n9794) );
  XOR2_X1 U9840 ( .A(P2_ADDR_REG_15__SCAN_IN), .B(n9794), .Z(n10245) );
  NOR2_X1 U9841 ( .A1(n10246), .A2(n10245), .ZN(n8765) );
  NOR2_X1 U9842 ( .A1(n8766), .A2(n8765), .ZN(n10248) );
  INV_X1 U9843 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n9819) );
  XOR2_X1 U9844 ( .A(P2_ADDR_REG_16__SCAN_IN), .B(n9819), .Z(n10247) );
  NOR2_X1 U9845 ( .A1(n10248), .A2(n10247), .ZN(n8767) );
  NOR2_X1 U9846 ( .A1(n8768), .A2(n8767), .ZN(n10250) );
  INV_X1 U9847 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9837) );
  XOR2_X1 U9848 ( .A(P2_ADDR_REG_17__SCAN_IN), .B(n9837), .Z(n10249) );
  NOR2_X1 U9849 ( .A1(n10250), .A2(n10249), .ZN(n8769) );
  NOR2_X1 U9850 ( .A1(n8770), .A2(n8769), .ZN(n8771) );
  AND2_X1 U9851 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(n8771), .ZN(n10251) );
  NOR2_X1 U9852 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n10251), .ZN(n8772) );
  NOR2_X1 U9853 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(n8771), .ZN(n10252) );
  NOR2_X1 U9854 ( .A1(n8772), .A2(n10252), .ZN(n8774) );
  XNOR2_X1 U9855 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n8773) );
  XNOR2_X1 U9856 ( .A(n8774), .B(n8773), .ZN(ADD_1071_U4) );
  INV_X1 U9857 ( .A(n8775), .ZN(n9043) );
  AOI22_X1 U9858 ( .A1(n8777), .A2(n9043), .B1(n8910), .B2(n8776), .ZN(n8779)
         );
  NOR2_X1 U9859 ( .A1(n9775), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8973) );
  INV_X1 U9860 ( .A(n8973), .ZN(n8778) );
  OAI211_X1 U9861 ( .C1(n8783), .C2(n8897), .A(n8779), .B(n8778), .ZN(n8780)
         );
  AOI21_X1 U9862 ( .B1(n8781), .B2(n8915), .A(n8780), .ZN(n8788) );
  INV_X1 U9863 ( .A(n8782), .ZN(n8786) );
  OAI22_X1 U9864 ( .A1(n8784), .A2(n8927), .B1(n8783), .B2(n8902), .ZN(n8785)
         );
  NAND3_X1 U9865 ( .A1(n8386), .A2(n8786), .A3(n8785), .ZN(n8787) );
  OAI211_X1 U9866 ( .C1(n8789), .C2(n8927), .A(n8788), .B(n8787), .ZN(P2_U3243) );
  INV_X1 U9867 ( .A(n8790), .ZN(n9377) );
  OAI222_X1 U9868 ( .A1(n8826), .A2(n9377), .B1(n5562), .B2(P1_U3084), .C1(
        n8791), .C2(n10196), .ZN(P1_U3323) );
  NOR2_X1 U9869 ( .A1(n9895), .A2(n9896), .ZN(n9894) );
  NOR2_X1 U9870 ( .A1(n9894), .A2(n8794), .ZN(n8797) );
  INV_X1 U9871 ( .A(n8797), .ZN(n8796) );
  INV_X1 U9872 ( .A(n8813), .ZN(n8795) );
  NAND2_X1 U9873 ( .A1(n8796), .A2(n8795), .ZN(n8799) );
  NAND2_X1 U9874 ( .A1(n8797), .A2(n8813), .ZN(n8798) );
  NAND2_X1 U9875 ( .A1(n8799), .A2(n8798), .ZN(n10074) );
  NOR2_X2 U9876 ( .A1(n10072), .A2(n9907), .ZN(n9888) );
  INV_X1 U9877 ( .A(n8802), .ZN(n8803) );
  AOI22_X1 U9878 ( .A1(n8803), .A2(n10561), .B1(P1_REG2_REG_29__SCAN_IN), .B2(
        n10563), .ZN(n8804) );
  OAI21_X1 U9879 ( .B1(n8805), .B2(n10565), .A(n8804), .ZN(n8822) );
  NOR2_X1 U9880 ( .A1(n5366), .A2(n8806), .ZN(n8808) );
  NAND2_X1 U9881 ( .A1(n8812), .A2(n8811), .ZN(n8814) );
  XNOR2_X1 U9882 ( .A(n8814), .B(n8813), .ZN(n8820) );
  NOR2_X1 U9883 ( .A1(n10260), .A2(n8815), .ZN(n8816) );
  NOR2_X1 U9884 ( .A1(n10489), .A2(n8816), .ZN(n9883) );
  NAND2_X1 U9885 ( .A1(n9568), .A2(n9883), .ZN(n8817) );
  AOI21_X2 U9886 ( .B1(n8820), .B2(n10546), .A(n8819), .ZN(n10073) );
  NOR2_X1 U9887 ( .A1(n10073), .A2(n10563), .ZN(n8821) );
  OAI21_X1 U9888 ( .B1(n10074), .B2(n10028), .A(n8823), .ZN(P1_U3355) );
  INV_X1 U9889 ( .A(n8824), .ZN(n9381) );
  OAI222_X1 U9890 ( .A1(n8826), .A2(n9381), .B1(n10209), .B2(n5585), .C1(
        P1_U3084), .C2(n8825), .ZN(P1_U3324) );
  XNOR2_X1 U9891 ( .A(n8828), .B(n8827), .ZN(n8835) );
  AOI22_X1 U9892 ( .A1(n9101), .A2(n8911), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        n4846), .ZN(n8832) );
  INV_X1 U9893 ( .A(n8830), .ZN(n9095) );
  NAND2_X1 U9894 ( .A1(n9095), .A2(n8910), .ZN(n8831) );
  OAI211_X1 U9895 ( .C1(n9069), .C2(n8913), .A(n8832), .B(n8831), .ZN(n8833)
         );
  AOI21_X1 U9896 ( .B1(n9289), .B2(n8915), .A(n8833), .ZN(n8834) );
  OAI21_X1 U9897 ( .B1(n8835), .B2(n8927), .A(n8834), .ZN(P2_U3216) );
  INV_X1 U9898 ( .A(n8836), .ZN(n8837) );
  NAND3_X1 U9899 ( .A1(n8837), .A2(n8875), .A3(n9179), .ZN(n8841) );
  NOR2_X1 U9900 ( .A1(n8921), .A2(n9156), .ZN(n8839) );
  INV_X1 U9901 ( .A(n9197), .ZN(n8930) );
  AOI22_X1 U9902 ( .A1(n9054), .A2(n9178), .B1(n9177), .B2(n8930), .ZN(n9152)
         );
  OAI22_X1 U9903 ( .A1(n9152), .A2(n8871), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9582), .ZN(n8838) );
  AOI211_X1 U9904 ( .C1(n9159), .C2(n8915), .A(n8839), .B(n8838), .ZN(n8840)
         );
  OAI211_X1 U9905 ( .C1(n8842), .C2(n8927), .A(n8841), .B(n8840), .ZN(P2_U3218) );
  AOI21_X1 U9906 ( .B1(n8844), .B2(n8843), .A(n8927), .ZN(n8846) );
  NAND2_X1 U9907 ( .A1(n8846), .A2(n8845), .ZN(n8851) );
  OAI22_X1 U9908 ( .A1(n8913), .A2(n10614), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6356), .ZN(n8847) );
  INV_X1 U9909 ( .A(n8847), .ZN(n8850) );
  AOI22_X1 U9910 ( .A1(n8911), .A2(n8939), .B1(n8910), .B2(n10630), .ZN(n8849)
         );
  NAND2_X1 U9911 ( .A1(n8915), .A2(n10606), .ZN(n8848) );
  NAND4_X1 U9912 ( .A1(n8851), .A2(n8850), .A3(n8849), .A4(n8848), .ZN(
        P2_U3219) );
  XNOR2_X1 U9913 ( .A(n8853), .B(n8852), .ZN(n8857) );
  INV_X1 U9914 ( .A(n9196), .ZN(n8931) );
  AOI22_X1 U9915 ( .A1(n8931), .A2(n9178), .B1(n9177), .B2(n8932), .ZN(n9228)
         );
  NAND2_X1 U9916 ( .A1(P2_U3152), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n9033) );
  NAND2_X1 U9917 ( .A1(n8910), .A2(n9231), .ZN(n8854) );
  OAI211_X1 U9918 ( .C1(n9228), .C2(n8871), .A(n9033), .B(n8854), .ZN(n8855)
         );
  AOI21_X1 U9919 ( .B1(n9333), .B2(n8915), .A(n8855), .ZN(n8856) );
  OAI21_X1 U9920 ( .B1(n8857), .B2(n8927), .A(n8856), .ZN(P2_U3221) );
  XNOR2_X1 U9921 ( .A(n8858), .B(n8859), .ZN(n8863) );
  OAI22_X1 U9922 ( .A1(n9197), .A2(n8913), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9644), .ZN(n8861) );
  OAI22_X1 U9923 ( .A1(n8897), .A2(n9196), .B1(n8921), .B2(n9190), .ZN(n8860)
         );
  AOI211_X1 U9924 ( .C1(n9321), .C2(n8915), .A(n8861), .B(n8860), .ZN(n8862)
         );
  OAI21_X1 U9925 ( .B1(n8863), .B2(n8927), .A(n8862), .ZN(P2_U3225) );
  NAND2_X1 U9926 ( .A1(n8865), .A2(n8864), .ZN(n8867) );
  XOR2_X1 U9927 ( .A(n8867), .B(n8866), .Z(n8874) );
  NOR2_X1 U9928 ( .A1(n8868), .A2(n10611), .ZN(n8869) );
  AOI21_X1 U9929 ( .B1(n9101), .B2(n9178), .A(n8869), .ZN(n9125) );
  AOI22_X1 U9930 ( .A1(n9129), .A2(n8910), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3152), .ZN(n8870) );
  OAI21_X1 U9931 ( .B1(n9125), .B2(n8871), .A(n8870), .ZN(n8872) );
  AOI21_X1 U9932 ( .B1(n9301), .B2(n8915), .A(n8872), .ZN(n8873) );
  OAI21_X1 U9933 ( .B1(n8874), .B2(n8927), .A(n8873), .ZN(P2_U3227) );
  NAND2_X1 U9934 ( .A1(n9054), .A2(n8875), .ZN(n8879) );
  OR2_X1 U9935 ( .A1(n8876), .A2(n8927), .ZN(n8878) );
  MUX2_X1 U9936 ( .A(n8879), .B(n8878), .S(n8877), .Z(n8883) );
  NOR2_X1 U9937 ( .A1(n9761), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8881) );
  OAI22_X1 U9938 ( .A1(n9144), .A2(n8913), .B1(n9138), .B2(n8921), .ZN(n8880)
         );
  AOI211_X1 U9939 ( .C1(n8911), .C2(n9179), .A(n8881), .B(n8880), .ZN(n8882)
         );
  OAI211_X1 U9940 ( .C1(n9055), .C2(n8922), .A(n8883), .B(n8882), .ZN(P2_U3231) );
  XNOR2_X1 U9941 ( .A(n8884), .B(n8885), .ZN(n8890) );
  OAI22_X1 U9942 ( .A1(n8913), .A2(n9214), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9661), .ZN(n8888) );
  INV_X1 U9943 ( .A(n9208), .ZN(n8886) );
  OAI22_X1 U9944 ( .A1(n8897), .A2(n9248), .B1(n8921), .B2(n8886), .ZN(n8887)
         );
  AOI211_X1 U9945 ( .C1(n9326), .C2(n8915), .A(n8888), .B(n8887), .ZN(n8889)
         );
  OAI21_X1 U9946 ( .B1(n8890), .B2(n8927), .A(n8889), .ZN(P2_U3235) );
  INV_X1 U9947 ( .A(n8891), .ZN(n8892) );
  AOI21_X1 U9948 ( .B1(n8894), .B2(n8893), .A(n8892), .ZN(n8901) );
  OAI22_X1 U9949 ( .A1(n9143), .A2(n8913), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8895), .ZN(n8899) );
  INV_X1 U9950 ( .A(n9170), .ZN(n8896) );
  OAI22_X1 U9951 ( .A1(n8897), .A2(n9214), .B1(n8921), .B2(n8896), .ZN(n8898)
         );
  AOI211_X1 U9952 ( .C1(n9316), .C2(n8915), .A(n8899), .B(n8898), .ZN(n8900)
         );
  OAI21_X1 U9953 ( .B1(n8901), .B2(n8927), .A(n8900), .ZN(P2_U3237) );
  NOR3_X1 U9954 ( .A1(n8903), .A2(n9047), .A3(n8902), .ZN(n8904) );
  AOI21_X1 U9955 ( .B1(n8906), .B2(n8905), .A(n8904), .ZN(n8918) );
  AOI21_X1 U9956 ( .B1(n8909), .B2(n8908), .A(n8907), .ZN(n8917) );
  AOI22_X1 U9957 ( .A1(n8911), .A2(n8933), .B1(n8910), .B2(n9242), .ZN(n8912)
         );
  NAND2_X1 U9958 ( .A1(n4846), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n9014) );
  OAI211_X1 U9959 ( .C1(n9248), .C2(n8913), .A(n8912), .B(n9014), .ZN(n8914)
         );
  AOI21_X1 U9960 ( .B1(n9336), .B2(n8915), .A(n8914), .ZN(n8916) );
  OAI21_X1 U9961 ( .B1(n8918), .B2(n8917), .A(n8916), .ZN(P2_U3240) );
  XNOR2_X1 U9962 ( .A(n8920), .B(n8919), .ZN(n8928) );
  OAI22_X1 U9963 ( .A1(n9059), .A2(n10613), .B1(n9144), .B2(n10611), .ZN(n9116) );
  OAI22_X1 U9964 ( .A1(n9108), .A2(n8921), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9779), .ZN(n8924) );
  INV_X1 U9965 ( .A(n9295), .ZN(n9111) );
  NOR2_X1 U9966 ( .A1(n9111), .A2(n8922), .ZN(n8923) );
  AOI211_X1 U9967 ( .C1(n8925), .C2(n9116), .A(n8924), .B(n8923), .ZN(n8926)
         );
  OAI21_X1 U9968 ( .B1(n8928), .B2(n8927), .A(n8926), .ZN(P2_U3242) );
  MUX2_X1 U9969 ( .A(n8929), .B(P2_DATAO_REG_31__SCAN_IN), .S(n8945), .Z(
        P2_U3583) );
  MUX2_X1 U9970 ( .A(n9100), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8945), .Z(
        P2_U3580) );
  MUX2_X1 U9971 ( .A(n9101), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8945), .Z(
        P2_U3578) );
  MUX2_X1 U9972 ( .A(n9054), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8945), .Z(
        P2_U3576) );
  MUX2_X1 U9973 ( .A(n9179), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8945), .Z(
        P2_U3575) );
  MUX2_X1 U9974 ( .A(n8930), .B(P2_DATAO_REG_22__SCAN_IN), .S(n8945), .Z(
        P2_U3574) );
  INV_X1 U9975 ( .A(n9214), .ZN(n9176) );
  MUX2_X1 U9976 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n9176), .S(P2_U3966), .Z(
        P2_U3573) );
  MUX2_X1 U9977 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8931), .S(P2_U3966), .Z(
        P2_U3572) );
  MUX2_X1 U9978 ( .A(n8932), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8945), .Z(
        P2_U3570) );
  MUX2_X1 U9979 ( .A(n8933), .B(P2_DATAO_REG_17__SCAN_IN), .S(n8945), .Z(
        P2_U3569) );
  MUX2_X1 U9980 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n9043), .S(P2_U3966), .Z(
        P2_U3568) );
  MUX2_X1 U9981 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8934), .S(P2_U3966), .Z(
        P2_U3567) );
  MUX2_X1 U9982 ( .A(n8494), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8945), .Z(
        P2_U3566) );
  MUX2_X1 U9983 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n8935), .S(P2_U3966), .Z(
        P2_U3565) );
  MUX2_X1 U9984 ( .A(n8936), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8945), .Z(
        P2_U3564) );
  MUX2_X1 U9985 ( .A(n8937), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8945), .Z(
        P2_U3563) );
  MUX2_X1 U9986 ( .A(n8938), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8945), .Z(
        P2_U3562) );
  MUX2_X1 U9987 ( .A(n8939), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8945), .Z(
        P2_U3561) );
  MUX2_X1 U9988 ( .A(n8940), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8945), .Z(
        P2_U3559) );
  MUX2_X1 U9989 ( .A(n8941), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8945), .Z(
        P2_U3558) );
  MUX2_X1 U9990 ( .A(n8942), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8945), .Z(
        P2_U3557) );
  MUX2_X1 U9991 ( .A(n8943), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8945), .Z(
        P2_U3556) );
  MUX2_X1 U9992 ( .A(n8944), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8945), .Z(
        P2_U3555) );
  MUX2_X1 U9993 ( .A(n6242), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8945), .Z(
        P2_U3554) );
  MUX2_X1 U9994 ( .A(n8946), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8945), .Z(
        P2_U3553) );
  MUX2_X1 U9995 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n6847), .S(P2_U3966), .Z(
        P2_U3552) );
  OAI211_X1 U9996 ( .C1(n8949), .C2(n8948), .A(n8976), .B(n8947), .ZN(n8957)
         );
  AOI22_X1 U9997 ( .A1(n10314), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(n4846), .ZN(n8956) );
  NAND2_X1 U9998 ( .A1(n10320), .A2(n8950), .ZN(n8955) );
  OAI211_X1 U9999 ( .C1(n8953), .C2(n8952), .A(n8993), .B(n8951), .ZN(n8954)
         );
  NAND4_X1 U10000 ( .A1(n8957), .A2(n8956), .A3(n8955), .A4(n8954), .ZN(
        P2_U3247) );
  OAI21_X1 U10001 ( .B1(n8960), .B2(n8959), .A(n8958), .ZN(n8961) );
  NAND2_X1 U10002 ( .A1(n8976), .A2(n8961), .ZN(n8970) );
  NOR2_X1 U10003 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9767), .ZN(n8962) );
  AOI21_X1 U10004 ( .B1(n10314), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n8962), .ZN(
        n8969) );
  NAND2_X1 U10005 ( .A1(n10320), .A2(n8963), .ZN(n8968) );
  OAI211_X1 U10006 ( .C1(n8966), .C2(n8965), .A(n8993), .B(n8964), .ZN(n8967)
         );
  NAND4_X1 U10007 ( .A1(n8970), .A2(n8969), .A3(n8968), .A4(n8967), .ZN(
        P2_U3256) );
  OAI211_X1 U10008 ( .C1(n8972), .C2(P2_REG1_REG_15__SCAN_IN), .A(n8993), .B(
        n8971), .ZN(n8982) );
  AOI21_X1 U10009 ( .B1(n10314), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n8973), .ZN(
        n8981) );
  OAI21_X1 U10010 ( .B1(n8975), .B2(n6440), .A(n8974), .ZN(n8977) );
  NAND2_X1 U10011 ( .A1(n8977), .A2(n8976), .ZN(n8980) );
  NAND2_X1 U10012 ( .A1(n10320), .A2(n8978), .ZN(n8979) );
  NAND4_X1 U10013 ( .A1(n8982), .A2(n8981), .A3(n8980), .A4(n8979), .ZN(
        P2_U3260) );
  AOI21_X1 U10014 ( .B1(n8989), .B2(P2_REG2_REG_16__SCAN_IN), .A(n8983), .ZN(
        n8987) );
  INV_X1 U10015 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8985) );
  NOR2_X1 U10016 ( .A1(n9004), .A2(n8985), .ZN(n8984) );
  AOI21_X1 U10017 ( .B1(n9004), .B2(n8985), .A(n8984), .ZN(n8986) );
  AOI211_X1 U10018 ( .C1(n8987), .C2(n8986), .A(n9003), .B(n10325), .ZN(n9000)
         );
  NOR2_X1 U10019 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9758), .ZN(n8988) );
  AOI21_X1 U10020 ( .B1(n10314), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n8988), .ZN(
        n8997) );
  INV_X1 U10021 ( .A(n8989), .ZN(n8992) );
  INV_X1 U10022 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8991) );
  AOI21_X1 U10023 ( .B1(n8992), .B2(n8991), .A(n8990), .ZN(n8995) );
  XNOR2_X1 U10024 ( .A(n9008), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n8994) );
  NAND2_X1 U10025 ( .A1(n8994), .A2(n8995), .ZN(n9007) );
  OAI211_X1 U10026 ( .C1(n8995), .C2(n8994), .A(n8993), .B(n9007), .ZN(n8996)
         );
  OAI211_X1 U10027 ( .C1(n8998), .C2(n9008), .A(n8997), .B(n8996), .ZN(n8999)
         );
  OR2_X1 U10028 ( .A1(n9000), .A2(n8999), .ZN(P2_U3262) );
  OR2_X1 U10029 ( .A1(n9017), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n9002) );
  NAND2_X1 U10030 ( .A1(n9017), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n9001) );
  NAND2_X1 U10031 ( .A1(n9002), .A2(n9001), .ZN(n9006) );
  AOI21_X1 U10032 ( .B1(n9006), .B2(n9005), .A(n9020), .ZN(n9019) );
  INV_X1 U10033 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n9009) );
  OAI21_X1 U10034 ( .B1(n9009), .B2(n9008), .A(n9007), .ZN(n9012) );
  INV_X1 U10035 ( .A(n9017), .ZN(n9022) );
  INV_X1 U10036 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n9010) );
  NAND2_X1 U10037 ( .A1(n9022), .A2(n9010), .ZN(n9026) );
  OAI21_X1 U10038 ( .B1(n9022), .B2(n9010), .A(n9026), .ZN(n9011) );
  NOR2_X1 U10039 ( .A1(n9011), .A2(n9012), .ZN(n9028) );
  AOI21_X1 U10040 ( .B1(n9012), .B2(n9011), .A(n9028), .ZN(n9015) );
  NAND2_X1 U10041 ( .A1(n10314), .A2(P2_ADDR_REG_18__SCAN_IN), .ZN(n9013) );
  OAI211_X1 U10042 ( .C1(n10329), .C2(n9015), .A(n9014), .B(n9013), .ZN(n9016)
         );
  AOI21_X1 U10043 ( .B1(n9017), .B2(n10320), .A(n9016), .ZN(n9018) );
  OAI21_X1 U10044 ( .B1(n9019), .B2(n10325), .A(n9018), .ZN(P2_U3263) );
  INV_X1 U10045 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n9021) );
  AOI21_X1 U10046 ( .B1(n9022), .B2(n9021), .A(n9020), .ZN(n9025) );
  XNOR2_X1 U10047 ( .A(n4849), .B(n9023), .ZN(n9024) );
  XNOR2_X1 U10048 ( .A(n9025), .B(n9024), .ZN(n9037) );
  INV_X1 U10049 ( .A(n9026), .ZN(n9027) );
  NOR2_X1 U10050 ( .A1(n9028), .A2(n9027), .ZN(n9031) );
  XNOR2_X1 U10051 ( .A(n9029), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n9030) );
  XNOR2_X1 U10052 ( .A(n9031), .B(n9030), .ZN(n9034) );
  NAND2_X1 U10053 ( .A1(n10314), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n9032) );
  OAI211_X1 U10054 ( .C1(n10329), .C2(n9034), .A(n9033), .B(n9032), .ZN(n9035)
         );
  AOI21_X1 U10055 ( .B1(n4849), .B2(n10320), .A(n9035), .ZN(n9036) );
  OAI21_X1 U10056 ( .B1(n10325), .B2(n9037), .A(n9036), .ZN(P2_U3264) );
  INV_X1 U10057 ( .A(n9038), .ZN(n9276) );
  NAND2_X1 U10058 ( .A1(n9074), .A2(n9039), .ZN(n9275) );
  NAND3_X1 U10059 ( .A1(n9276), .A2(n10626), .A3(n9275), .ZN(n9042) );
  AOI21_X1 U10060 ( .B1(n9157), .B2(P2_REG2_REG_30__SCAN_IN), .A(n9040), .ZN(
        n9041) );
  OAI211_X1 U10061 ( .C1(n5151), .C2(n10634), .A(n9042), .B(n9041), .ZN(
        P2_U3266) );
  INV_X1 U10062 ( .A(n9045), .ZN(n9263) );
  INV_X1 U10063 ( .A(n9336), .ZN(n9244) );
  INV_X1 U10064 ( .A(n9248), .ZN(n9049) );
  NAND2_X1 U10065 ( .A1(n9333), .A2(n9049), .ZN(n9050) );
  NAND2_X1 U10066 ( .A1(n9185), .A2(n9052), .ZN(n9168) );
  INV_X1 U10067 ( .A(n9316), .ZN(n9172) );
  NAND2_X1 U10068 ( .A1(n9159), .A2(n9179), .ZN(n9053) );
  INV_X1 U10069 ( .A(n9301), .ZN(n9132) );
  NAND2_X1 U10070 ( .A1(n9081), .A2(n9060), .ZN(n9062) );
  NAND2_X1 U10071 ( .A1(n9062), .A2(n9061), .ZN(n9063) );
  XNOR2_X1 U10072 ( .A(n9063), .B(n9064), .ZN(n9279) );
  INV_X1 U10073 ( .A(n9279), .ZN(n9080) );
  XNOR2_X1 U10074 ( .A(n9065), .B(n6790), .ZN(n9066) );
  NAND2_X1 U10075 ( .A1(n9066), .A2(n10616), .ZN(n9072) );
  OAI22_X1 U10076 ( .A1(n9069), .A2(n10611), .B1(n9068), .B2(n9067), .ZN(n9070) );
  INV_X1 U10077 ( .A(n9070), .ZN(n9071) );
  NAND2_X1 U10078 ( .A1(n9072), .A2(n9071), .ZN(n9282) );
  OAI21_X1 U10079 ( .B1(n8603), .B2(n9073), .A(n9074), .ZN(n9281) );
  AOI22_X1 U10080 ( .A1(n9075), .A2(n10629), .B1(P2_REG2_REG_29__SCAN_IN), 
        .B2(n10631), .ZN(n9077) );
  NAND2_X1 U10081 ( .A1(n9280), .A2(n10451), .ZN(n9076) );
  OAI211_X1 U10082 ( .C1(n9281), .C2(n10454), .A(n9077), .B(n9076), .ZN(n9078)
         );
  AOI21_X1 U10083 ( .B1(n9282), .B2(n10448), .A(n9078), .ZN(n9079) );
  OAI21_X1 U10084 ( .B1(n9080), .B2(n9255), .A(n9079), .ZN(P2_U3267) );
  XNOR2_X1 U10085 ( .A(n9081), .B(n6594), .ZN(n9288) );
  AOI21_X1 U10086 ( .B1(n9284), .B2(n9092), .A(n9073), .ZN(n9285) );
  AOI22_X1 U10087 ( .A1(n9082), .A2(n10629), .B1(P2_REG2_REG_28__SCAN_IN), 
        .B2(n9157), .ZN(n9083) );
  OAI21_X1 U10088 ( .B1(n5155), .B2(n10634), .A(n9083), .ZN(n9089) );
  OAI21_X1 U10089 ( .B1(n9085), .B2(n6594), .A(n9084), .ZN(n9087) );
  AOI21_X1 U10090 ( .B1(n9087), .B2(n10616), .A(n9086), .ZN(n9287) );
  NOR2_X1 U10091 ( .A1(n9287), .A2(n10631), .ZN(n9088) );
  AOI211_X1 U10092 ( .C1(n10626), .C2(n9285), .A(n9089), .B(n9088), .ZN(n9090)
         );
  OAI21_X1 U10093 ( .B1(n9288), .B2(n9255), .A(n9090), .ZN(P2_U3268) );
  XNOR2_X1 U10094 ( .A(n9091), .B(n9099), .ZN(n9293) );
  INV_X1 U10095 ( .A(n9107), .ZN(n9094) );
  INV_X1 U10096 ( .A(n9092), .ZN(n9093) );
  AOI21_X1 U10097 ( .B1(n9289), .B2(n9094), .A(n9093), .ZN(n9290) );
  AOI22_X1 U10098 ( .A1(n9095), .A2(n10629), .B1(P2_REG2_REG_27__SCAN_IN), 
        .B2(n9157), .ZN(n9096) );
  OAI21_X1 U10099 ( .B1(n9097), .B2(n10634), .A(n9096), .ZN(n9104) );
  XNOR2_X1 U10100 ( .A(n9098), .B(n9099), .ZN(n9102) );
  AOI222_X1 U10101 ( .A1(n10616), .A2(n9102), .B1(n9101), .B2(n9177), .C1(
        n9100), .C2(n9178), .ZN(n9292) );
  NOR2_X1 U10102 ( .A1(n9292), .A2(n10631), .ZN(n9103) );
  AOI211_X1 U10103 ( .C1(n10626), .C2(n9290), .A(n9104), .B(n9103), .ZN(n9105)
         );
  OAI21_X1 U10104 ( .B1(n9293), .B2(n9255), .A(n9105), .ZN(P2_U3269) );
  XOR2_X1 U10105 ( .A(n9115), .B(n9106), .Z(n9298) );
  AOI211_X1 U10106 ( .C1(n9295), .C2(n9127), .A(n10673), .B(n9107), .ZN(n9294)
         );
  INV_X1 U10107 ( .A(n9108), .ZN(n9109) );
  AOI22_X1 U10108 ( .A1(n9109), .A2(n10629), .B1(P2_REG2_REG_26__SCAN_IN), 
        .B2(n9157), .ZN(n9110) );
  OAI21_X1 U10109 ( .B1(n9111), .B2(n10634), .A(n9110), .ZN(n9119) );
  NAND2_X1 U10110 ( .A1(n9122), .A2(n9113), .ZN(n9114) );
  XOR2_X1 U10111 ( .A(n9115), .B(n9114), .Z(n9117) );
  AOI21_X1 U10112 ( .B1(n9117), .B2(n10616), .A(n9116), .ZN(n9297) );
  NOR2_X1 U10113 ( .A1(n9297), .A2(n10631), .ZN(n9118) );
  AOI211_X1 U10114 ( .C1(n9294), .C2(n9266), .A(n9119), .B(n9118), .ZN(n9120)
         );
  OAI21_X1 U10115 ( .B1(n9298), .B2(n9255), .A(n9120), .ZN(P2_U3270) );
  XNOR2_X1 U10116 ( .A(n9121), .B(n9124), .ZN(n9303) );
  OAI211_X1 U10117 ( .C1(n9124), .C2(n9123), .A(n9122), .B(n10616), .ZN(n9126)
         );
  NAND2_X1 U10118 ( .A1(n9126), .A2(n9125), .ZN(n9299) );
  AOI211_X1 U10119 ( .C1(n9301), .C2(n9128), .A(n10673), .B(n8602), .ZN(n9300)
         );
  NAND2_X1 U10120 ( .A1(n9300), .A2(n9266), .ZN(n9131) );
  AOI22_X1 U10121 ( .A1(n9129), .A2(n10629), .B1(P2_REG2_REG_25__SCAN_IN), 
        .B2(n10631), .ZN(n9130) );
  OAI211_X1 U10122 ( .C1(n9132), .C2(n10634), .A(n9131), .B(n9130), .ZN(n9133)
         );
  AOI21_X1 U10123 ( .B1(n9299), .B2(n10448), .A(n9133), .ZN(n9134) );
  OAI21_X1 U10124 ( .B1(n9303), .B2(n9255), .A(n9134), .ZN(P2_U3271) );
  INV_X1 U10125 ( .A(n9135), .ZN(n9136) );
  AOI21_X1 U10126 ( .B1(n6550), .B2(n9137), .A(n9136), .ZN(n9308) );
  XNOR2_X1 U10127 ( .A(n9155), .B(n9304), .ZN(n9305) );
  INV_X1 U10128 ( .A(n9138), .ZN(n9139) );
  AOI22_X1 U10129 ( .A1(n9139), .A2(n10629), .B1(P2_REG2_REG_24__SCAN_IN), 
        .B2(n9157), .ZN(n9140) );
  OAI21_X1 U10130 ( .B1(n9055), .B2(n10634), .A(n9140), .ZN(n9149) );
  AOI21_X1 U10131 ( .B1(n9142), .B2(n9141), .A(n10436), .ZN(n9147) );
  OAI22_X1 U10132 ( .A1(n9144), .A2(n10613), .B1(n9143), .B2(n10611), .ZN(
        n9145) );
  AOI21_X1 U10133 ( .B1(n9147), .B2(n9146), .A(n9145), .ZN(n9307) );
  NOR2_X1 U10134 ( .A1(n9307), .A2(n10631), .ZN(n9148) );
  AOI211_X1 U10135 ( .C1(n9305), .C2(n10626), .A(n9149), .B(n9148), .ZN(n9150)
         );
  OAI21_X1 U10136 ( .B1(n9308), .B2(n9255), .A(n9150), .ZN(P2_U3272) );
  XOR2_X1 U10137 ( .A(n9151), .B(n9162), .Z(n9153) );
  OAI21_X1 U10138 ( .B1(n9153), .B2(n10436), .A(n9152), .ZN(n9314) );
  NOR2_X1 U10139 ( .A1(n9169), .A2(n9311), .ZN(n9154) );
  OR2_X1 U10140 ( .A1(n9155), .A2(n9154), .ZN(n9312) );
  INV_X1 U10141 ( .A(n9156), .ZN(n9158) );
  AOI22_X1 U10142 ( .A1(n9158), .A2(n10629), .B1(P2_REG2_REG_23__SCAN_IN), 
        .B2(n9157), .ZN(n9161) );
  NAND2_X1 U10143 ( .A1(n9159), .A2(n10451), .ZN(n9160) );
  OAI211_X1 U10144 ( .C1(n9312), .C2(n10454), .A(n9161), .B(n9160), .ZN(n9166)
         );
  NOR2_X1 U10145 ( .A1(n9163), .A2(n9162), .ZN(n9310) );
  INV_X1 U10146 ( .A(n9164), .ZN(n9309) );
  NOR3_X1 U10147 ( .A1(n9310), .A2(n9309), .A3(n9255), .ZN(n9165) );
  AOI211_X1 U10148 ( .C1(n10448), .C2(n9314), .A(n9166), .B(n9165), .ZN(n9167)
         );
  INV_X1 U10149 ( .A(n9167), .ZN(P2_U3273) );
  XNOR2_X1 U10150 ( .A(n9168), .B(n9174), .ZN(n9320) );
  AOI21_X1 U10151 ( .B1(n9316), .B2(n9189), .A(n9169), .ZN(n9317) );
  AOI22_X1 U10152 ( .A1(n10631), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n9170), 
        .B2(n10629), .ZN(n9171) );
  OAI21_X1 U10153 ( .B1(n9172), .B2(n10634), .A(n9171), .ZN(n9183) );
  OAI211_X1 U10154 ( .C1(n9175), .C2(n9174), .A(n9173), .B(n10616), .ZN(n9181)
         );
  AOI22_X1 U10155 ( .A1(n9179), .A2(n9178), .B1(n9177), .B2(n9176), .ZN(n9180)
         );
  NOR2_X1 U10156 ( .A1(n9319), .A2(n10631), .ZN(n9182) );
  AOI211_X1 U10157 ( .C1(n9317), .C2(n10626), .A(n9183), .B(n9182), .ZN(n9184)
         );
  OAI21_X1 U10158 ( .B1(n9320), .B2(n9255), .A(n9184), .ZN(P2_U3274) );
  INV_X1 U10159 ( .A(n9185), .ZN(n9186) );
  AOI21_X1 U10160 ( .B1(n9188), .B2(n9187), .A(n9186), .ZN(n9325) );
  AOI21_X1 U10161 ( .B1(n9321), .B2(n9206), .A(n5161), .ZN(n9322) );
  INV_X1 U10162 ( .A(n9321), .ZN(n9193) );
  INV_X1 U10163 ( .A(n9190), .ZN(n9191) );
  AOI22_X1 U10164 ( .A1(n10631), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n9191), 
        .B2(n10629), .ZN(n9192) );
  OAI21_X1 U10165 ( .B1(n9193), .B2(n10634), .A(n9192), .ZN(n9202) );
  INV_X1 U10166 ( .A(n9194), .ZN(n9195) );
  AOI21_X1 U10167 ( .B1(n9195), .B2(n9051), .A(n10436), .ZN(n9200) );
  OAI22_X1 U10168 ( .A1(n9197), .A2(n10613), .B1(n9196), .B2(n10611), .ZN(
        n9198) );
  AOI21_X1 U10169 ( .B1(n9200), .B2(n9199), .A(n9198), .ZN(n9324) );
  NOR2_X1 U10170 ( .A1(n9324), .A2(n10631), .ZN(n9201) );
  AOI211_X1 U10171 ( .C1(n9322), .C2(n10626), .A(n9202), .B(n9201), .ZN(n9203)
         );
  OAI21_X1 U10172 ( .B1(n9325), .B2(n9255), .A(n9203), .ZN(P2_U3275) );
  OAI21_X1 U10173 ( .B1(n9205), .B2(n9212), .A(n9204), .ZN(n9330) );
  INV_X1 U10174 ( .A(n9230), .ZN(n9207) );
  AOI21_X1 U10175 ( .B1(n9326), .B2(n9207), .A(n5159), .ZN(n9327) );
  AOI22_X1 U10176 ( .A1(n10631), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n9208), 
        .B2(n10629), .ZN(n9209) );
  OAI21_X1 U10177 ( .B1(n9210), .B2(n10634), .A(n9209), .ZN(n9219) );
  INV_X1 U10178 ( .A(n9211), .ZN(n9213) );
  AOI21_X1 U10179 ( .B1(n9213), .B2(n9212), .A(n10436), .ZN(n9217) );
  OAI22_X1 U10180 ( .A1(n9214), .A2(n10613), .B1(n9248), .B2(n10611), .ZN(
        n9215) );
  AOI21_X1 U10181 ( .B1(n9217), .B2(n9216), .A(n9215), .ZN(n9329) );
  NOR2_X1 U10182 ( .A1(n9329), .A2(n10631), .ZN(n9218) );
  AOI211_X1 U10183 ( .C1(n9327), .C2(n10626), .A(n9219), .B(n9218), .ZN(n9220)
         );
  OAI21_X1 U10184 ( .B1(n9330), .B2(n9255), .A(n9220), .ZN(P2_U3276) );
  OAI21_X1 U10185 ( .B1(n9221), .B2(n9224), .A(n9222), .ZN(n9335) );
  AOI22_X1 U10186 ( .A1(n9333), .A2(n10451), .B1(n9157), .B2(
        P2_REG2_REG_19__SCAN_IN), .ZN(n9236) );
  NAND3_X1 U10187 ( .A1(n9223), .A2(n9225), .A3(n9224), .ZN(n9226) );
  NAND3_X1 U10188 ( .A1(n9227), .A2(n10616), .A3(n9226), .ZN(n9229) );
  NAND2_X1 U10189 ( .A1(n9229), .A2(n9228), .ZN(n9331) );
  AOI211_X1 U10190 ( .C1(n9333), .C2(n9239), .A(n10673), .B(n9230), .ZN(n9332)
         );
  INV_X1 U10191 ( .A(n9332), .ZN(n9233) );
  INV_X1 U10192 ( .A(n9231), .ZN(n9232) );
  OAI22_X1 U10193 ( .A1(n9233), .A2(n4849), .B1(n10446), .B2(n9232), .ZN(n9234) );
  OAI21_X1 U10194 ( .B1(n9331), .B2(n9234), .A(n10448), .ZN(n9235) );
  OAI211_X1 U10195 ( .C1(n9335), .C2(n9255), .A(n9236), .B(n9235), .ZN(
        P2_U3277) );
  XNOR2_X1 U10196 ( .A(n9238), .B(n9237), .ZN(n9340) );
  INV_X1 U10197 ( .A(n9239), .ZN(n9240) );
  AOI21_X1 U10198 ( .B1(n9336), .B2(n9241), .A(n9240), .ZN(n9337) );
  AOI22_X1 U10199 ( .A1(n10631), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n9242), 
        .B2(n10629), .ZN(n9243) );
  OAI21_X1 U10200 ( .B1(n9244), .B2(n10634), .A(n9243), .ZN(n9253) );
  INV_X1 U10201 ( .A(n9245), .ZN(n9247) );
  AOI21_X1 U10202 ( .B1(n9247), .B2(n9246), .A(n10436), .ZN(n9251) );
  OAI22_X1 U10203 ( .A1(n9249), .A2(n10611), .B1(n9248), .B2(n10613), .ZN(
        n9250) );
  AOI21_X1 U10204 ( .B1(n9251), .B2(n9223), .A(n9250), .ZN(n9339) );
  NOR2_X1 U10205 ( .A1(n9339), .A2(n10631), .ZN(n9252) );
  AOI211_X1 U10206 ( .C1(n9337), .C2(n10626), .A(n9253), .B(n9252), .ZN(n9254)
         );
  OAI21_X1 U10207 ( .B1(n9340), .B2(n9255), .A(n9254), .ZN(P2_U3278) );
  NAND2_X1 U10208 ( .A1(n8535), .A2(n9256), .ZN(n9258) );
  NAND2_X1 U10209 ( .A1(n9258), .A2(n9257), .ZN(n9259) );
  XNOR2_X1 U10210 ( .A(n9259), .B(n9263), .ZN(n9261) );
  AOI21_X1 U10211 ( .B1(n9261), .B2(n10616), .A(n9260), .ZN(n9345) );
  OAI21_X1 U10212 ( .B1(n4915), .B2(n9263), .A(n9262), .ZN(n9341) );
  XNOR2_X1 U10213 ( .A(n9264), .B(n9343), .ZN(n9265) );
  AND2_X1 U10214 ( .A1(n9265), .A2(n10663), .ZN(n9342) );
  NAND2_X1 U10215 ( .A1(n9342), .A2(n9266), .ZN(n9269) );
  AOI22_X1 U10216 ( .A1(n10631), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n9267), 
        .B2(n10629), .ZN(n9268) );
  OAI211_X1 U10217 ( .C1(n9270), .C2(n10634), .A(n9269), .B(n9268), .ZN(n9271)
         );
  AOI21_X1 U10218 ( .B1(n9341), .B2(n10456), .A(n9271), .ZN(n9272) );
  OAI21_X1 U10219 ( .B1(n9157), .B2(n9345), .A(n9272), .ZN(P2_U3279) );
  NAND2_X1 U10220 ( .A1(n6781), .A2(n10662), .ZN(n9273) );
  OAI211_X1 U10221 ( .C1(n9274), .C2(n10673), .A(n9273), .B(n9277), .ZN(n9353)
         );
  MUX2_X1 U10222 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n9353), .S(n10681), .Z(
        P2_U3551) );
  NAND3_X1 U10223 ( .A1(n9276), .A2(n10663), .A3(n9275), .ZN(n9278) );
  OAI211_X1 U10224 ( .C1(n5151), .C2(n10672), .A(n9278), .B(n9277), .ZN(n9354)
         );
  MUX2_X1 U10225 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n9354), .S(n10681), .Z(
        P2_U3550) );
  NAND2_X1 U10226 ( .A1(n9279), .A2(n10677), .ZN(n9283) );
  MUX2_X1 U10227 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n9355), .S(n10681), .Z(
        P2_U3549) );
  AOI22_X1 U10228 ( .A1(n9285), .A2(n10663), .B1(n10662), .B2(n9284), .ZN(
        n9286) );
  OAI211_X1 U10229 ( .C1(n9288), .C2(n10667), .A(n9287), .B(n9286), .ZN(n9356)
         );
  MUX2_X1 U10230 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n9356), .S(n10681), .Z(
        P2_U3548) );
  AOI22_X1 U10231 ( .A1(n9290), .A2(n10663), .B1(n10662), .B2(n9289), .ZN(
        n9291) );
  OAI211_X1 U10232 ( .C1(n9293), .C2(n10667), .A(n9292), .B(n9291), .ZN(n9357)
         );
  MUX2_X1 U10233 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n9357), .S(n10681), .Z(
        P2_U3547) );
  AOI21_X1 U10234 ( .B1(n10662), .B2(n9295), .A(n9294), .ZN(n9296) );
  OAI211_X1 U10235 ( .C1(n9298), .C2(n10667), .A(n9297), .B(n9296), .ZN(n9358)
         );
  MUX2_X1 U10236 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n9358), .S(n10681), .Z(
        P2_U3546) );
  AOI211_X1 U10237 ( .C1(n10662), .C2(n9301), .A(n9300), .B(n9299), .ZN(n9302)
         );
  OAI21_X1 U10238 ( .B1(n9303), .B2(n10667), .A(n9302), .ZN(n9359) );
  MUX2_X1 U10239 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n9359), .S(n10681), .Z(
        P2_U3545) );
  AOI22_X1 U10240 ( .A1(n9305), .A2(n10663), .B1(n10662), .B2(n9304), .ZN(
        n9306) );
  OAI211_X1 U10241 ( .C1(n9308), .C2(n10667), .A(n9307), .B(n9306), .ZN(n9360)
         );
  MUX2_X1 U10242 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n9360), .S(n10681), .Z(
        P2_U3544) );
  NOR3_X1 U10243 ( .A1(n9310), .A2(n9309), .A3(n10667), .ZN(n9315) );
  OAI22_X1 U10244 ( .A1(n9312), .A2(n10673), .B1(n9311), .B2(n10672), .ZN(
        n9313) );
  MUX2_X1 U10245 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n9361), .S(n10681), .Z(
        P2_U3543) );
  AOI22_X1 U10246 ( .A1(n9317), .A2(n10663), .B1(n10662), .B2(n9316), .ZN(
        n9318) );
  OAI211_X1 U10247 ( .C1(n9320), .C2(n10667), .A(n9319), .B(n9318), .ZN(n9362)
         );
  MUX2_X1 U10248 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n9362), .S(n10681), .Z(
        P2_U3542) );
  AOI22_X1 U10249 ( .A1(n9322), .A2(n10663), .B1(n10662), .B2(n9321), .ZN(
        n9323) );
  OAI211_X1 U10250 ( .C1(n9325), .C2(n10667), .A(n9324), .B(n9323), .ZN(n9363)
         );
  MUX2_X1 U10251 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n9363), .S(n10681), .Z(
        P2_U3541) );
  AOI22_X1 U10252 ( .A1(n9327), .A2(n10663), .B1(n10662), .B2(n9326), .ZN(
        n9328) );
  OAI211_X1 U10253 ( .C1(n9330), .C2(n10667), .A(n9329), .B(n9328), .ZN(n9364)
         );
  MUX2_X1 U10254 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n9364), .S(n10681), .Z(
        P2_U3540) );
  AOI211_X1 U10255 ( .C1(n10662), .C2(n9333), .A(n9332), .B(n9331), .ZN(n9334)
         );
  OAI21_X1 U10256 ( .B1(n9335), .B2(n10667), .A(n9334), .ZN(n9365) );
  MUX2_X1 U10257 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n9365), .S(n10681), .Z(
        P2_U3539) );
  AOI22_X1 U10258 ( .A1(n9337), .A2(n10663), .B1(n10662), .B2(n9336), .ZN(
        n9338) );
  OAI211_X1 U10259 ( .C1(n9340), .C2(n10667), .A(n9339), .B(n9338), .ZN(n9366)
         );
  MUX2_X1 U10260 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n9366), .S(n10681), .Z(
        P2_U3538) );
  INV_X1 U10261 ( .A(n9341), .ZN(n9346) );
  AOI21_X1 U10262 ( .B1(n10662), .B2(n9343), .A(n9342), .ZN(n9344) );
  OAI211_X1 U10263 ( .C1(n9346), .C2(n10667), .A(n9345), .B(n9344), .ZN(n9367)
         );
  MUX2_X1 U10264 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n9367), .S(n10681), .Z(
        P2_U3537) );
  INV_X1 U10265 ( .A(n9347), .ZN(n9352) );
  AOI21_X1 U10266 ( .B1(n10662), .B2(n9349), .A(n9348), .ZN(n9350) );
  OAI211_X1 U10267 ( .C1(n9352), .C2(n10667), .A(n9351), .B(n9350), .ZN(n9368)
         );
  MUX2_X1 U10268 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n9368), .S(n10681), .Z(
        P2_U3536) );
  MUX2_X1 U10269 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n9353), .S(n10684), .Z(
        P2_U3519) );
  MUX2_X1 U10270 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n9354), .S(n10684), .Z(
        P2_U3518) );
  MUX2_X1 U10271 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n9355), .S(n10684), .Z(
        P2_U3517) );
  MUX2_X1 U10272 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n9356), .S(n10684), .Z(
        P2_U3516) );
  MUX2_X1 U10273 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n9357), .S(n10684), .Z(
        P2_U3515) );
  MUX2_X1 U10274 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n9358), .S(n10684), .Z(
        P2_U3514) );
  MUX2_X1 U10275 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n9359), .S(n10684), .Z(
        P2_U3513) );
  MUX2_X1 U10276 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n9360), .S(n10684), .Z(
        P2_U3512) );
  MUX2_X1 U10277 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n9361), .S(n10684), .Z(
        P2_U3511) );
  MUX2_X1 U10278 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n9362), .S(n10684), .Z(
        P2_U3510) );
  MUX2_X1 U10279 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n9363), .S(n10684), .Z(
        P2_U3509) );
  MUX2_X1 U10280 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n9364), .S(n10684), .Z(
        P2_U3508) );
  MUX2_X1 U10281 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n9365), .S(n10684), .Z(
        P2_U3507) );
  MUX2_X1 U10282 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n9366), .S(n10684), .Z(
        P2_U3505) );
  MUX2_X1 U10283 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n9367), .S(n10684), .Z(
        P2_U3502) );
  MUX2_X1 U10284 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n9368), .S(n10684), .Z(
        P2_U3499) );
  INV_X1 U10285 ( .A(n9369), .ZN(n9374) );
  NOR4_X1 U10286 ( .A1(n9371), .A2(P2_IR_REG_30__SCAN_IN), .A3(n9370), .A4(
        n4846), .ZN(n9372) );
  AOI21_X1 U10287 ( .B1(P1_DATAO_REG_31__SCAN_IN), .B2(n9378), .A(n9372), .ZN(
        n9373) );
  OAI21_X1 U10288 ( .B1(n9374), .B2(n8243), .A(n9373), .ZN(P2_U3327) );
  AOI22_X1 U10289 ( .A1(n9375), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n9378), .ZN(n9376) );
  OAI21_X1 U10290 ( .B1(n9377), .B2(n8243), .A(n9376), .ZN(P2_U3328) );
  AOI22_X1 U10291 ( .A1(n9379), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n9378), .ZN(n9380) );
  OAI21_X1 U10292 ( .B1(n9381), .B2(n8243), .A(n9380), .ZN(P2_U3329) );
  INV_X1 U10293 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n9383) );
  INV_X1 U10294 ( .A(n6582), .ZN(n9382) );
  OAI222_X1 U10295 ( .A1(n9387), .A2(n9383), .B1(P2_U3152), .B2(n6841), .C1(
        n8243), .C2(n9382), .ZN(P2_U3330) );
  INV_X1 U10296 ( .A(n10205), .ZN(n9384) );
  OAI222_X1 U10297 ( .A1(n9387), .A2(n9386), .B1(n4846), .B2(n9385), .C1(n8243), .C2(n9384), .ZN(P2_U3331) );
  MUX2_X1 U10298 ( .A(n9388), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  XNOR2_X1 U10299 ( .A(n9390), .B(n9389), .ZN(n9391) );
  XNOR2_X1 U10300 ( .A(n9392), .B(n9391), .ZN(n9399) );
  AOI22_X1 U10301 ( .A1(n9393), .A2(n9556), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3084), .ZN(n9395) );
  NAND2_X1 U10302 ( .A1(n9923), .A2(n9558), .ZN(n9394) );
  OAI211_X1 U10303 ( .C1(n9396), .C2(n9561), .A(n9395), .B(n9394), .ZN(n9397)
         );
  AOI21_X1 U10304 ( .B1(n10082), .B2(n9564), .A(n9397), .ZN(n9398) );
  OAI21_X1 U10305 ( .B1(n9399), .B2(n9566), .A(n9398), .ZN(P1_U3212) );
  NAND2_X1 U10306 ( .A1(n9401), .A2(n9400), .ZN(n9402) );
  XOR2_X1 U10307 ( .A(n9403), .B(n9402), .Z(n9412) );
  NAND2_X1 U10308 ( .A1(n9404), .A2(n9558), .ZN(n9406) );
  OAI211_X1 U10309 ( .C1(n9465), .C2(n9561), .A(n9406), .B(n9405), .ZN(n9409)
         );
  NOR2_X1 U10310 ( .A1(n9407), .A2(n9548), .ZN(n9408) );
  AOI211_X1 U10311 ( .C1(n9410), .C2(n9556), .A(n9409), .B(n9408), .ZN(n9411)
         );
  OAI21_X1 U10312 ( .B1(n9412), .B2(n9566), .A(n9411), .ZN(P1_U3213) );
  NAND2_X1 U10313 ( .A1(n9481), .A2(n9413), .ZN(n9414) );
  XOR2_X1 U10314 ( .A(n9415), .B(n9414), .Z(n9420) );
  NAND2_X1 U10315 ( .A1(n9954), .A2(n9545), .ZN(n9417) );
  AOI22_X1 U10316 ( .A1(n9955), .A2(n9558), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3084), .ZN(n9416) );
  OAI211_X1 U10317 ( .C1(n9516), .C2(n9948), .A(n9417), .B(n9416), .ZN(n9418)
         );
  AOI21_X1 U10318 ( .B1(n10102), .B2(n9564), .A(n9418), .ZN(n9419) );
  OAI21_X1 U10319 ( .B1(n9420), .B2(n9566), .A(n9419), .ZN(P1_U3214) );
  INV_X1 U10320 ( .A(n9422), .ZN(n9423) );
  AOI21_X1 U10321 ( .B1(n9424), .B2(n9421), .A(n9423), .ZN(n9429) );
  NAND2_X1 U10322 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9875) );
  NAND2_X1 U10323 ( .A1(n10022), .A2(n9545), .ZN(n9425) );
  OAI211_X1 U10324 ( .C1(n9474), .C2(n9542), .A(n9875), .B(n9425), .ZN(n9427)
         );
  NOR2_X1 U10325 ( .A1(n10018), .A2(n9548), .ZN(n9426) );
  AOI211_X1 U10326 ( .C1(n10016), .C2(n9556), .A(n9427), .B(n9426), .ZN(n9428)
         );
  OAI21_X1 U10327 ( .B1(n9429), .B2(n9566), .A(n9428), .ZN(P1_U3217) );
  INV_X1 U10328 ( .A(n9430), .ZN(n9432) );
  NOR2_X1 U10329 ( .A1(n9432), .A2(n9431), .ZN(n9433) );
  XNOR2_X1 U10330 ( .A(n9434), .B(n9433), .ZN(n9441) );
  OAI22_X1 U10331 ( .A1(n9436), .A2(n9542), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9435), .ZN(n9437) );
  AOI21_X1 U10332 ( .B1(n9545), .B2(n9955), .A(n9437), .ZN(n9438) );
  OAI21_X1 U10333 ( .B1(n9516), .B2(n9986), .A(n9438), .ZN(n9439) );
  AOI21_X1 U10334 ( .B1(n10113), .B2(n9564), .A(n9439), .ZN(n9440) );
  OAI21_X1 U10335 ( .B1(n9441), .B2(n9566), .A(n9440), .ZN(P1_U3221) );
  INV_X1 U10336 ( .A(n9442), .ZN(n9444) );
  NAND2_X1 U10337 ( .A1(n9444), .A2(n9443), .ZN(n9445) );
  XNOR2_X1 U10338 ( .A(n9446), .B(n9445), .ZN(n9454) );
  OAI22_X1 U10339 ( .A1(n9448), .A2(n9542), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9447), .ZN(n9449) );
  AOI21_X1 U10340 ( .B1(n9917), .B2(n9556), .A(n9449), .ZN(n9450) );
  OAI21_X1 U10341 ( .B1(n9451), .B2(n9561), .A(n9450), .ZN(n9452) );
  AOI21_X1 U10342 ( .B1(n10092), .B2(n9564), .A(n9452), .ZN(n9453) );
  OAI21_X1 U10343 ( .B1(n9454), .B2(n9566), .A(n9453), .ZN(P1_U3223) );
  INV_X1 U10344 ( .A(n9456), .ZN(n9457) );
  NOR2_X1 U10345 ( .A1(n9455), .A2(n9457), .ZN(n9550) );
  NAND2_X1 U10346 ( .A1(n9455), .A2(n9457), .ZN(n9551) );
  OAI21_X1 U10347 ( .B1(n9550), .B2(n9553), .A(n9551), .ZN(n9461) );
  XNOR2_X1 U10348 ( .A(n9459), .B(n9458), .ZN(n9460) );
  XNOR2_X1 U10349 ( .A(n9461), .B(n9460), .ZN(n9468) );
  NAND2_X1 U10350 ( .A1(n9556), .A2(n9462), .ZN(n9464) );
  AOI22_X1 U10351 ( .A1(n9545), .A2(n9573), .B1(P1_REG3_REG_16__SCAN_IN), .B2(
        P1_U3084), .ZN(n9463) );
  OAI211_X1 U10352 ( .C1(n9465), .C2(n9542), .A(n9464), .B(n9463), .ZN(n9466)
         );
  AOI21_X1 U10353 ( .B1(n10141), .B2(n9564), .A(n9466), .ZN(n9467) );
  OAI21_X1 U10354 ( .B1(n9468), .B2(n9566), .A(n9467), .ZN(P1_U3224) );
  XNOR2_X1 U10355 ( .A(n9471), .B(n9470), .ZN(n9472) );
  XNOR2_X1 U10356 ( .A(n9469), .B(n9472), .ZN(n9478) );
  NAND2_X1 U10357 ( .A1(n10053), .A2(n9558), .ZN(n9473) );
  NAND2_X1 U10358 ( .A1(P1_U3084), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9834) );
  OAI211_X1 U10359 ( .C1(n9474), .C2(n9561), .A(n9473), .B(n9834), .ZN(n9476)
         );
  NOR2_X1 U10360 ( .A1(n7061), .A2(n9548), .ZN(n9475) );
  AOI211_X1 U10361 ( .C1(n10060), .C2(n9556), .A(n9476), .B(n9475), .ZN(n9477)
         );
  OAI21_X1 U10362 ( .B1(n9478), .B2(n9566), .A(n9477), .ZN(P1_U3226) );
  INV_X1 U10363 ( .A(n9479), .ZN(n9484) );
  AOI21_X1 U10364 ( .B1(n9482), .B2(n9481), .A(n9480), .ZN(n9483) );
  OAI21_X1 U10365 ( .B1(n9484), .B2(n9483), .A(n9536), .ZN(n9488) );
  AOI22_X1 U10366 ( .A1(n9969), .A2(n9558), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3084), .ZN(n9485) );
  OAI21_X1 U10367 ( .B1(n9516), .B2(n9938), .A(n9485), .ZN(n9486) );
  AOI21_X1 U10368 ( .B1(n9930), .B2(n9545), .A(n9486), .ZN(n9487) );
  OAI211_X1 U10369 ( .C1(n9489), .C2(n9548), .A(n9488), .B(n9487), .ZN(
        P1_U3227) );
  AND2_X1 U10370 ( .A1(n9491), .A2(n9490), .ZN(n9494) );
  OAI211_X1 U10371 ( .C1(n9494), .C2(n9493), .A(n9536), .B(n9492), .ZN(n9501)
         );
  NAND2_X1 U10372 ( .A1(P1_U3084), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n10352) );
  INV_X1 U10373 ( .A(n10352), .ZN(n9495) );
  AOI21_X1 U10374 ( .B1(n5777), .B2(n9558), .A(n9495), .ZN(n9500) );
  AOI22_X1 U10375 ( .A1(n9791), .A2(n9545), .B1(n9496), .B2(n9564), .ZN(n9499)
         );
  INV_X1 U10376 ( .A(n10421), .ZN(n9497) );
  OR2_X1 U10377 ( .A1(n9516), .A2(n9497), .ZN(n9498) );
  NAND4_X1 U10378 ( .A1(n9501), .A2(n9500), .A3(n9499), .A4(n9498), .ZN(
        P1_U3228) );
  NAND2_X1 U10379 ( .A1(n8655), .A2(n9503), .ZN(n9504) );
  XNOR2_X1 U10380 ( .A(n9505), .B(n9504), .ZN(n9510) );
  NAND2_X1 U10381 ( .A1(n9970), .A2(n9545), .ZN(n9507) );
  AOI22_X1 U10382 ( .A1(n9558), .A2(n9572), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3084), .ZN(n9506) );
  OAI211_X1 U10383 ( .C1(n9516), .C2(n10006), .A(n9507), .B(n9506), .ZN(n9508)
         );
  AOI21_X1 U10384 ( .B1(n10117), .B2(n9564), .A(n9508), .ZN(n9509) );
  OAI21_X1 U10385 ( .B1(n9510), .B2(n9566), .A(n9509), .ZN(P1_U3231) );
  XOR2_X1 U10386 ( .A(n9512), .B(n9511), .Z(n9519) );
  OAI22_X1 U10387 ( .A1(n10000), .A2(n9542), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9513), .ZN(n9514) );
  AOI21_X1 U10388 ( .B1(n9545), .B2(n9969), .A(n9514), .ZN(n9515) );
  OAI21_X1 U10389 ( .B1(n9516), .B2(n9963), .A(n9515), .ZN(n9517) );
  AOI21_X1 U10390 ( .B1(n10106), .B2(n9564), .A(n9517), .ZN(n9518) );
  OAI21_X1 U10391 ( .B1(n9519), .B2(n9566), .A(n9518), .ZN(P1_U3233) );
  NAND2_X1 U10392 ( .A1(n9522), .A2(n9536), .ZN(n9526) );
  AOI22_X1 U10393 ( .A1(n5777), .A2(n9545), .B1(n9558), .B2(n7491), .ZN(n9525)
         );
  AOI22_X1 U10394 ( .A1(n9523), .A2(P1_REG3_REG_2__SCAN_IN), .B1(n9564), .B2(
        n10364), .ZN(n9524) );
  NAND3_X1 U10395 ( .A1(n9526), .A2(n9525), .A3(n9524), .ZN(P1_U3235) );
  XOR2_X1 U10396 ( .A(n9528), .B(n9527), .Z(n9529) );
  XNOR2_X1 U10397 ( .A(n9530), .B(n9529), .ZN(n9535) );
  NAND2_X1 U10398 ( .A1(n9545), .A2(n9572), .ZN(n9531) );
  NAND2_X1 U10399 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9860) );
  OAI211_X1 U10400 ( .C1(n10035), .C2(n9542), .A(n9531), .B(n9860), .ZN(n9533)
         );
  INV_X1 U10401 ( .A(n10043), .ZN(n10128) );
  NOR2_X1 U10402 ( .A1(n10128), .A2(n9548), .ZN(n9532) );
  AOI211_X1 U10403 ( .C1(n10041), .C2(n9556), .A(n9533), .B(n9532), .ZN(n9534)
         );
  OAI21_X1 U10404 ( .B1(n9535), .B2(n9566), .A(n9534), .ZN(P1_U3236) );
  OAI211_X1 U10405 ( .C1(n9539), .C2(n9538), .A(n9537), .B(n9536), .ZN(n9547)
         );
  AOI22_X1 U10406 ( .A1(n9540), .A2(n9556), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3084), .ZN(n9541) );
  OAI21_X1 U10407 ( .B1(n9543), .B2(n9542), .A(n9541), .ZN(n9544) );
  AOI21_X1 U10408 ( .B1(n9571), .B2(n9545), .A(n9544), .ZN(n9546) );
  OAI211_X1 U10409 ( .C1(n9549), .C2(n9548), .A(n9547), .B(n9546), .ZN(
        P1_U3238) );
  INV_X1 U10410 ( .A(n9550), .ZN(n9552) );
  NAND2_X1 U10411 ( .A1(n9552), .A2(n9551), .ZN(n9554) );
  XNOR2_X1 U10412 ( .A(n9554), .B(n9553), .ZN(n9567) );
  NAND2_X1 U10413 ( .A1(n9556), .A2(n9555), .ZN(n9560) );
  NOR2_X1 U10414 ( .A1(n9557), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9796) );
  AOI21_X1 U10415 ( .B1(n9558), .B2(n9786), .A(n9796), .ZN(n9559) );
  OAI211_X1 U10416 ( .C1(n9562), .C2(n9561), .A(n9560), .B(n9559), .ZN(n9563)
         );
  AOI21_X1 U10417 ( .B1(n10146), .B2(n9564), .A(n9563), .ZN(n9565) );
  OAI21_X1 U10418 ( .B1(n9567), .B2(n9566), .A(n9565), .ZN(P1_U3239) );
  MUX2_X1 U10419 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n9884), .S(P1_U4006), .Z(
        P1_U3586) );
  MUX2_X1 U10420 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9568), .S(P1_U4006), .Z(
        P1_U3585) );
  MUX2_X1 U10421 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9569), .S(P1_U4006), .Z(
        P1_U3584) );
  MUX2_X1 U10422 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9570), .S(P1_U4006), .Z(
        P1_U3583) );
  MUX2_X1 U10423 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9571), .S(P1_U4006), .Z(
        P1_U3582) );
  MUX2_X1 U10424 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9923), .S(P1_U4006), .Z(
        P1_U3581) );
  MUX2_X1 U10425 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9930), .S(P1_U4006), .Z(
        P1_U3580) );
  MUX2_X1 U10426 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9954), .S(P1_U4006), .Z(
        P1_U3579) );
  MUX2_X1 U10427 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9969), .S(P1_U4006), .Z(
        P1_U3578) );
  MUX2_X1 U10428 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9955), .S(P1_U4006), .Z(
        P1_U3577) );
  MUX2_X1 U10429 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9970), .S(P1_U4006), .Z(
        P1_U3576) );
  MUX2_X1 U10430 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n10022), .S(P1_U4006), .Z(
        P1_U3575) );
  MUX2_X1 U10431 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9572), .S(P1_U4006), .Z(
        P1_U3574) );
  MUX2_X1 U10432 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n10052), .S(P1_U4006), .Z(
        P1_U3573) );
  MUX2_X1 U10433 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9573), .S(P1_U4006), .Z(
        n9785) );
  INV_X1 U10434 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n9772) );
  OAI22_X1 U10435 ( .A1(n9772), .A2(keyinput_59), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(keyinput_62), .ZN(n9574) );
  AOI221_X1 U10436 ( .B1(n9772), .B2(keyinput_59), .C1(keyinput_62), .C2(
        P2_REG3_REG_26__SCAN_IN), .A(n9574), .ZN(n9577) );
  OAI22_X1 U10437 ( .A1(n9775), .A2(keyinput_63), .B1(keyinput_61), .B2(
        P2_REG3_REG_6__SCAN_IN), .ZN(n9575) );
  AOI221_X1 U10438 ( .B1(n9775), .B2(keyinput_63), .C1(P2_REG3_REG_6__SCAN_IN), 
        .C2(keyinput_61), .A(n9575), .ZN(n9576) );
  OAI211_X1 U10439 ( .C1(P2_REG3_REG_18__SCAN_IN), .C2(keyinput_60), .A(n9577), 
        .B(n9576), .ZN(n9578) );
  AOI21_X1 U10440 ( .B1(P2_REG3_REG_18__SCAN_IN), .B2(keyinput_60), .A(n9578), 
        .ZN(n9783) );
  INV_X1 U10441 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n9659) );
  AOI22_X1 U10442 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(keyinput_52), .B1(n9669), 
        .B2(keyinput_53), .ZN(n9579) );
  OAI221_X1 U10443 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(keyinput_52), .C1(n9669), 
        .C2(keyinput_53), .A(n9579), .ZN(n9657) );
  INV_X1 U10444 ( .A(keyinput_51), .ZN(n9655) );
  INV_X1 U10445 ( .A(keyinput_50), .ZN(n9653) );
  AOI22_X1 U10446 ( .A1(P2_REG3_REG_25__SCAN_IN), .A2(keyinput_47), .B1(n6449), 
        .B2(keyinput_48), .ZN(n9580) );
  OAI221_X1 U10447 ( .B1(P2_REG3_REG_25__SCAN_IN), .B2(keyinput_47), .C1(n6449), .C2(keyinput_48), .A(n9580), .ZN(n9650) );
  AOI22_X1 U10448 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(keyinput_39), .B1(n9582), 
        .B2(keyinput_38), .ZN(n9581) );
  OAI221_X1 U10449 ( .B1(P2_REG3_REG_10__SCAN_IN), .B2(keyinput_39), .C1(n9582), .C2(keyinput_38), .A(n9581), .ZN(n9639) );
  OAI22_X1 U10450 ( .A1(n9716), .A2(keyinput_22), .B1(keyinput_23), .B2(SI_9_), 
        .ZN(n9583) );
  AOI221_X1 U10451 ( .B1(n9716), .B2(keyinput_22), .C1(SI_9_), .C2(keyinput_23), .A(n9583), .ZN(n9621) );
  INV_X1 U10452 ( .A(SI_6_), .ZN(n9714) );
  OAI22_X1 U10453 ( .A1(n9714), .A2(keyinput_26), .B1(keyinput_27), .B2(SI_5_), 
        .ZN(n9584) );
  AOI221_X1 U10454 ( .B1(n9714), .B2(keyinput_26), .C1(SI_5_), .C2(keyinput_27), .A(n9584), .ZN(n9620) );
  INV_X1 U10455 ( .A(SI_7_), .ZN(n9717) );
  OAI22_X1 U10456 ( .A1(n9586), .A2(keyinput_24), .B1(n9717), .B2(keyinput_25), 
        .ZN(n9585) );
  AOI221_X1 U10457 ( .B1(n9586), .B2(keyinput_24), .C1(keyinput_25), .C2(n9717), .A(n9585), .ZN(n9619) );
  INV_X1 U10458 ( .A(keyinput_17), .ZN(n9611) );
  INV_X1 U10459 ( .A(keyinput_16), .ZN(n9609) );
  INV_X1 U10460 ( .A(keyinput_15), .ZN(n9607) );
  AOI22_X1 U10461 ( .A1(SI_31_), .A2(keyinput_1), .B1(SI_29_), .B2(keyinput_3), 
        .ZN(n9587) );
  OAI221_X1 U10462 ( .B1(SI_31_), .B2(keyinput_1), .C1(SI_29_), .C2(keyinput_3), .A(n9587), .ZN(n9590) );
  AOI22_X1 U10463 ( .A1(P2_WR_REG_SCAN_IN), .A2(keyinput_0), .B1(SI_30_), .B2(
        keyinput_2), .ZN(n9588) );
  OAI221_X1 U10464 ( .B1(P2_WR_REG_SCAN_IN), .B2(keyinput_0), .C1(SI_30_), 
        .C2(keyinput_2), .A(n9588), .ZN(n9589) );
  OAI22_X1 U10465 ( .A1(n9590), .A2(n9589), .B1(n5530), .B2(keyinput_4), .ZN(
        n9591) );
  AOI21_X1 U10466 ( .B1(n5530), .B2(keyinput_4), .A(n9591), .ZN(n9600) );
  OAI22_X1 U10467 ( .A1(n9593), .A2(keyinput_5), .B1(keyinput_6), .B2(SI_26_), 
        .ZN(n9592) );
  AOI221_X1 U10468 ( .B1(n9593), .B2(keyinput_5), .C1(SI_26_), .C2(keyinput_6), 
        .A(n9592), .ZN(n9599) );
  AOI22_X1 U10469 ( .A1(SI_24_), .A2(keyinput_8), .B1(n9595), .B2(keyinput_10), 
        .ZN(n9594) );
  OAI221_X1 U10470 ( .B1(SI_24_), .B2(keyinput_8), .C1(n9595), .C2(keyinput_10), .A(n9594), .ZN(n9598) );
  AOI22_X1 U10471 ( .A1(SI_23_), .A2(keyinput_9), .B1(SI_25_), .B2(keyinput_7), 
        .ZN(n9596) );
  OAI221_X1 U10472 ( .B1(SI_23_), .B2(keyinput_9), .C1(SI_25_), .C2(keyinput_7), .A(n9596), .ZN(n9597) );
  AOI211_X1 U10473 ( .C1(n9600), .C2(n9599), .A(n9598), .B(n9597), .ZN(n9605)
         );
  INV_X1 U10474 ( .A(SI_21_), .ZN(n9678) );
  AOI22_X1 U10475 ( .A1(n9678), .A2(keyinput_11), .B1(keyinput_14), .B2(n9677), 
        .ZN(n9601) );
  OAI221_X1 U10476 ( .B1(n9678), .B2(keyinput_11), .C1(n9677), .C2(keyinput_14), .A(n9601), .ZN(n9604) );
  AOI22_X1 U10477 ( .A1(SI_19_), .A2(keyinput_13), .B1(SI_20_), .B2(
        keyinput_12), .ZN(n9602) );
  OAI221_X1 U10478 ( .B1(SI_19_), .B2(keyinput_13), .C1(SI_20_), .C2(
        keyinput_12), .A(n9602), .ZN(n9603) );
  NOR3_X1 U10479 ( .A1(n9605), .A2(n9604), .A3(n9603), .ZN(n9606) );
  AOI221_X1 U10480 ( .B1(SI_17_), .B2(n9607), .C1(n9700), .C2(keyinput_15), 
        .A(n9606), .ZN(n9608) );
  AOI221_X1 U10481 ( .B1(SI_16_), .B2(keyinput_16), .C1(n9703), .C2(n9609), 
        .A(n9608), .ZN(n9610) );
  AOI221_X1 U10482 ( .B1(SI_15_), .B2(keyinput_17), .C1(n9705), .C2(n9611), 
        .A(n9610), .ZN(n9617) );
  AOI22_X1 U10483 ( .A1(SI_13_), .A2(keyinput_19), .B1(SI_14_), .B2(
        keyinput_18), .ZN(n9612) );
  OAI221_X1 U10484 ( .B1(SI_13_), .B2(keyinput_19), .C1(SI_14_), .C2(
        keyinput_18), .A(n9612), .ZN(n9616) );
  OAI22_X1 U10485 ( .A1(n9614), .A2(keyinput_20), .B1(keyinput_21), .B2(SI_11_), .ZN(n9613) );
  AOI221_X1 U10486 ( .B1(n9614), .B2(keyinput_20), .C1(SI_11_), .C2(
        keyinput_21), .A(n9613), .ZN(n9615) );
  OAI21_X1 U10487 ( .B1(n9617), .B2(n9616), .A(n9615), .ZN(n9618) );
  NAND4_X1 U10488 ( .A1(n9621), .A2(n9620), .A3(n9619), .A4(n9618), .ZN(n9624)
         );
  INV_X1 U10489 ( .A(keyinput_28), .ZN(n9622) );
  MUX2_X1 U10490 ( .A(n9622), .B(keyinput_28), .S(SI_4_), .Z(n9623) );
  NAND2_X1 U10491 ( .A1(n9624), .A2(n9623), .ZN(n9627) );
  INV_X1 U10492 ( .A(keyinput_29), .ZN(n9625) );
  MUX2_X1 U10493 ( .A(keyinput_29), .B(n9625), .S(SI_3_), .Z(n9626) );
  NAND2_X1 U10494 ( .A1(n9627), .A2(n9626), .ZN(n9630) );
  OAI22_X1 U10495 ( .A1(SI_2_), .A2(keyinput_30), .B1(SI_0_), .B2(keyinput_32), 
        .ZN(n9628) );
  AOI221_X1 U10496 ( .B1(SI_2_), .B2(keyinput_30), .C1(keyinput_32), .C2(SI_0_), .A(n9628), .ZN(n9629) );
  OAI211_X1 U10497 ( .C1(SI_1_), .C2(keyinput_31), .A(n9630), .B(n9629), .ZN(
        n9631) );
  AOI21_X1 U10498 ( .B1(SI_1_), .B2(keyinput_31), .A(n9631), .ZN(n9637) );
  XNOR2_X1 U10499 ( .A(P2_RD_REG_SCAN_IN), .B(keyinput_33), .ZN(n9636) );
  AOI22_X1 U10500 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(keyinput_35), .B1(
        P2_U3152), .B2(keyinput_34), .ZN(n9632) );
  OAI221_X1 U10501 ( .B1(P2_REG3_REG_7__SCAN_IN), .B2(keyinput_35), .C1(n4846), 
        .C2(keyinput_34), .A(n9632), .ZN(n9635) );
  AOI22_X1 U10502 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(keyinput_37), .B1(n9735), 
        .B2(keyinput_36), .ZN(n9633) );
  OAI221_X1 U10503 ( .B1(P2_REG3_REG_14__SCAN_IN), .B2(keyinput_37), .C1(n9735), .C2(keyinput_36), .A(n9633), .ZN(n9634) );
  NOR4_X1 U10504 ( .A1(n9637), .A2(n9636), .A3(n9635), .A4(n9634), .ZN(n9638)
         );
  OAI22_X1 U10505 ( .A1(n9639), .A2(n9638), .B1(n6585), .B2(keyinput_42), .ZN(
        n9640) );
  AOI21_X1 U10506 ( .B1(n6585), .B2(keyinput_42), .A(n9640), .ZN(n9648) );
  OAI22_X1 U10507 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(keyinput_40), .B1(
        P2_REG3_REG_19__SCAN_IN), .B2(keyinput_41), .ZN(n9641) );
  AOI221_X1 U10508 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(keyinput_40), .C1(
        keyinput_41), .C2(P2_REG3_REG_19__SCAN_IN), .A(n9641), .ZN(n9647) );
  AOI22_X1 U10509 ( .A1(n6392), .A2(keyinput_46), .B1(n8068), .B2(keyinput_43), 
        .ZN(n9642) );
  OAI221_X1 U10510 ( .B1(n6392), .B2(keyinput_46), .C1(n8068), .C2(keyinput_43), .A(n9642), .ZN(n9646) );
  AOI22_X1 U10511 ( .A1(P2_REG3_REG_1__SCAN_IN), .A2(keyinput_44), .B1(n9644), 
        .B2(keyinput_45), .ZN(n9643) );
  OAI221_X1 U10512 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(keyinput_44), .C1(n9644), 
        .C2(keyinput_45), .A(n9643), .ZN(n9645) );
  AOI211_X1 U10513 ( .C1(n9648), .C2(n9647), .A(n9646), .B(n9645), .ZN(n9649)
         );
  OAI22_X1 U10514 ( .A1(n9650), .A2(n9649), .B1(keyinput_49), .B2(
        P2_REG3_REG_5__SCAN_IN), .ZN(n9651) );
  AOI21_X1 U10515 ( .B1(keyinput_49), .B2(P2_REG3_REG_5__SCAN_IN), .A(n9651), 
        .ZN(n9652) );
  AOI221_X1 U10516 ( .B1(P2_REG3_REG_17__SCAN_IN), .B2(keyinput_50), .C1(n9758), .C2(n9653), .A(n9652), .ZN(n9654) );
  AOI221_X1 U10517 ( .B1(P2_REG3_REG_24__SCAN_IN), .B2(keyinput_51), .C1(n9761), .C2(n9655), .A(n9654), .ZN(n9656) );
  OAI22_X1 U10518 ( .A1(keyinput_54), .A2(n9659), .B1(n9657), .B2(n9656), .ZN(
        n9658) );
  AOI21_X1 U10519 ( .B1(keyinput_54), .B2(n9659), .A(n9658), .ZN(n9665) );
  AOI22_X1 U10520 ( .A1(n9661), .A2(keyinput_55), .B1(n9667), .B2(keyinput_56), 
        .ZN(n9660) );
  OAI221_X1 U10521 ( .B1(n9661), .B2(keyinput_55), .C1(n9667), .C2(keyinput_56), .A(n9660), .ZN(n9664) );
  OAI22_X1 U10522 ( .A1(n9767), .A2(keyinput_58), .B1(keyinput_57), .B2(
        P2_REG3_REG_22__SCAN_IN), .ZN(n9662) );
  AOI221_X1 U10523 ( .B1(n9767), .B2(keyinput_58), .C1(P2_REG3_REG_22__SCAN_IN), .C2(keyinput_57), .A(n9662), .ZN(n9663) );
  OAI21_X1 U10524 ( .B1(n9665), .B2(n9664), .A(n9663), .ZN(n9782) );
  OAI22_X1 U10525 ( .A1(n9667), .A2(keyinput_120), .B1(P2_REG3_REG_20__SCAN_IN), .B2(keyinput_119), .ZN(n9666) );
  AOI221_X1 U10526 ( .B1(n9667), .B2(keyinput_120), .C1(keyinput_119), .C2(
        P2_REG3_REG_20__SCAN_IN), .A(n9666), .ZN(n9770) );
  INV_X1 U10527 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n9670) );
  OAI22_X1 U10528 ( .A1(n9670), .A2(keyinput_116), .B1(n9669), .B2(
        keyinput_117), .ZN(n9668) );
  AOI221_X1 U10529 ( .B1(n9670), .B2(keyinput_116), .C1(keyinput_117), .C2(
        n9669), .A(n9668), .ZN(n9764) );
  INV_X1 U10530 ( .A(keyinput_115), .ZN(n9762) );
  INV_X1 U10531 ( .A(keyinput_114), .ZN(n9759) );
  AOI22_X1 U10532 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(keyinput_112), .B1(n9672), .B2(keyinput_111), .ZN(n9671) );
  OAI221_X1 U10533 ( .B1(P2_REG3_REG_16__SCAN_IN), .B2(keyinput_112), .C1(
        n9672), .C2(keyinput_111), .A(n9671), .ZN(n9756) );
  AOI22_X1 U10534 ( .A1(P2_REG3_REG_23__SCAN_IN), .A2(keyinput_102), .B1(n6356), .B2(keyinput_103), .ZN(n9673) );
  OAI221_X1 U10535 ( .B1(P2_REG3_REG_23__SCAN_IN), .B2(keyinput_102), .C1(
        n6356), .C2(keyinput_103), .A(n9673), .ZN(n9742) );
  OAI22_X1 U10536 ( .A1(n9675), .A2(keyinput_83), .B1(keyinput_82), .B2(SI_14_), .ZN(n9674) );
  AOI221_X1 U10537 ( .B1(n9675), .B2(keyinput_83), .C1(SI_14_), .C2(
        keyinput_82), .A(n9674), .ZN(n9710) );
  INV_X1 U10538 ( .A(keyinput_81), .ZN(n9706) );
  INV_X1 U10539 ( .A(keyinput_80), .ZN(n9702) );
  INV_X1 U10540 ( .A(keyinput_79), .ZN(n9699) );
  OAI22_X1 U10541 ( .A1(n9678), .A2(keyinput_75), .B1(n9677), .B2(keyinput_78), 
        .ZN(n9676) );
  AOI221_X1 U10542 ( .B1(n9678), .B2(keyinput_75), .C1(keyinput_78), .C2(n9677), .A(n9676), .ZN(n9697) );
  OAI22_X1 U10543 ( .A1(SI_20_), .A2(keyinput_76), .B1(keyinput_77), .B2(
        SI_19_), .ZN(n9679) );
  AOI221_X1 U10544 ( .B1(SI_20_), .B2(keyinput_76), .C1(SI_19_), .C2(
        keyinput_77), .A(n9679), .ZN(n9696) );
  OAI22_X1 U10545 ( .A1(SI_29_), .A2(keyinput_67), .B1(P2_WR_REG_SCAN_IN), 
        .B2(keyinput_64), .ZN(n9680) );
  AOI221_X1 U10546 ( .B1(SI_29_), .B2(keyinput_67), .C1(keyinput_64), .C2(
        P2_WR_REG_SCAN_IN), .A(n9680), .ZN(n9684) );
  OAI22_X1 U10547 ( .A1(n9682), .A2(keyinput_66), .B1(keyinput_65), .B2(SI_31_), .ZN(n9681) );
  AOI221_X1 U10548 ( .B1(n9682), .B2(keyinput_66), .C1(SI_31_), .C2(
        keyinput_65), .A(n9681), .ZN(n9683) );
  AOI22_X1 U10549 ( .A1(n9684), .A2(n9683), .B1(keyinput_68), .B2(n5530), .ZN(
        n9685) );
  OAI21_X1 U10550 ( .B1(keyinput_68), .B2(n5530), .A(n9685), .ZN(n9694) );
  AOI22_X1 U10551 ( .A1(SI_27_), .A2(keyinput_69), .B1(n9687), .B2(keyinput_70), .ZN(n9686) );
  OAI221_X1 U10552 ( .B1(SI_27_), .B2(keyinput_69), .C1(n9687), .C2(
        keyinput_70), .A(n9686), .ZN(n9693) );
  OAI22_X1 U10553 ( .A1(n9689), .A2(keyinput_71), .B1(keyinput_74), .B2(SI_22_), .ZN(n9688) );
  AOI221_X1 U10554 ( .B1(n9689), .B2(keyinput_71), .C1(SI_22_), .C2(
        keyinput_74), .A(n9688), .ZN(n9692) );
  OAI22_X1 U10555 ( .A1(SI_24_), .A2(keyinput_72), .B1(keyinput_73), .B2(
        SI_23_), .ZN(n9690) );
  AOI221_X1 U10556 ( .B1(SI_24_), .B2(keyinput_72), .C1(SI_23_), .C2(
        keyinput_73), .A(n9690), .ZN(n9691) );
  OAI211_X1 U10557 ( .C1(n9694), .C2(n9693), .A(n9692), .B(n9691), .ZN(n9695)
         );
  NAND3_X1 U10558 ( .A1(n9697), .A2(n9696), .A3(n9695), .ZN(n9698) );
  OAI221_X1 U10559 ( .B1(SI_17_), .B2(keyinput_79), .C1(n9700), .C2(n9699), 
        .A(n9698), .ZN(n9701) );
  OAI221_X1 U10560 ( .B1(SI_16_), .B2(keyinput_80), .C1(n9703), .C2(n9702), 
        .A(n9701), .ZN(n9704) );
  OAI221_X1 U10561 ( .B1(SI_15_), .B2(n9706), .C1(n9705), .C2(keyinput_81), 
        .A(n9704), .ZN(n9709) );
  AOI22_X1 U10562 ( .A1(SI_12_), .A2(keyinput_84), .B1(SI_11_), .B2(
        keyinput_85), .ZN(n9707) );
  OAI221_X1 U10563 ( .B1(SI_12_), .B2(keyinput_84), .C1(SI_11_), .C2(
        keyinput_85), .A(n9707), .ZN(n9708) );
  AOI21_X1 U10564 ( .B1(n9710), .B2(n9709), .A(n9708), .ZN(n9721) );
  AOI22_X1 U10565 ( .A1(SI_8_), .A2(keyinput_88), .B1(n9712), .B2(keyinput_87), 
        .ZN(n9711) );
  OAI221_X1 U10566 ( .B1(SI_8_), .B2(keyinput_88), .C1(n9712), .C2(keyinput_87), .A(n9711), .ZN(n9720) );
  AOI22_X1 U10567 ( .A1(SI_5_), .A2(keyinput_91), .B1(n9714), .B2(keyinput_90), 
        .ZN(n9713) );
  OAI221_X1 U10568 ( .B1(SI_5_), .B2(keyinput_91), .C1(n9714), .C2(keyinput_90), .A(n9713), .ZN(n9719) );
  AOI22_X1 U10569 ( .A1(n9717), .A2(keyinput_89), .B1(n9716), .B2(keyinput_86), 
        .ZN(n9715) );
  OAI221_X1 U10570 ( .B1(n9717), .B2(keyinput_89), .C1(n9716), .C2(keyinput_86), .A(n9715), .ZN(n9718) );
  NOR4_X1 U10571 ( .A1(n9721), .A2(n9720), .A3(n9719), .A4(n9718), .ZN(n9724)
         );
  INV_X1 U10572 ( .A(keyinput_92), .ZN(n9722) );
  MUX2_X1 U10573 ( .A(n9722), .B(keyinput_92), .S(SI_4_), .Z(n9723) );
  NOR2_X1 U10574 ( .A1(n9724), .A2(n9723), .ZN(n9727) );
  INV_X1 U10575 ( .A(keyinput_93), .ZN(n9725) );
  MUX2_X1 U10576 ( .A(n9725), .B(keyinput_93), .S(SI_3_), .Z(n9726) );
  NOR2_X1 U10577 ( .A1(n9727), .A2(n9726), .ZN(n9733) );
  XNOR2_X1 U10578 ( .A(n9728), .B(keyinput_95), .ZN(n9732) );
  XOR2_X1 U10579 ( .A(SI_0_), .B(keyinput_96), .Z(n9731) );
  XNOR2_X1 U10580 ( .A(n9729), .B(keyinput_94), .ZN(n9730) );
  NOR4_X1 U10581 ( .A1(n9733), .A2(n9732), .A3(n9731), .A4(n9730), .ZN(n9740)
         );
  AOI22_X1 U10582 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(keyinput_99), .B1(n9735), 
        .B2(keyinput_100), .ZN(n9734) );
  OAI221_X1 U10583 ( .B1(P2_REG3_REG_7__SCAN_IN), .B2(keyinput_99), .C1(n9735), 
        .C2(keyinput_100), .A(n9734), .ZN(n9739) );
  AOI22_X1 U10584 ( .A1(P2_STATE_REG_SCAN_IN), .A2(keyinput_98), .B1(
        P2_RD_REG_SCAN_IN), .B2(keyinput_97), .ZN(n9736) );
  OAI221_X1 U10585 ( .B1(P2_STATE_REG_SCAN_IN), .B2(keyinput_98), .C1(
        P2_RD_REG_SCAN_IN), .C2(keyinput_97), .A(n9736), .ZN(n9738) );
  XNOR2_X1 U10586 ( .A(P2_REG3_REG_14__SCAN_IN), .B(keyinput_101), .ZN(n9737)
         );
  NOR4_X1 U10587 ( .A1(n9740), .A2(n9739), .A3(n9738), .A4(n9737), .ZN(n9741)
         );
  OAI22_X1 U10588 ( .A1(n9742), .A2(n9741), .B1(P2_REG3_REG_19__SCAN_IN), .B2(
        keyinput_105), .ZN(n9743) );
  AOI21_X1 U10589 ( .B1(P2_REG3_REG_19__SCAN_IN), .B2(keyinput_105), .A(n9743), 
        .ZN(n9752) );
  OAI22_X1 U10590 ( .A1(n9745), .A2(keyinput_104), .B1(n6585), .B2(
        keyinput_106), .ZN(n9744) );
  AOI221_X1 U10591 ( .B1(n9745), .B2(keyinput_104), .C1(keyinput_106), .C2(
        n6585), .A(n9744), .ZN(n9751) );
  AOI22_X1 U10592 ( .A1(n9747), .A2(keyinput_108), .B1(n6392), .B2(
        keyinput_110), .ZN(n9746) );
  OAI221_X1 U10593 ( .B1(n9747), .B2(keyinput_108), .C1(n6392), .C2(
        keyinput_110), .A(n9746), .ZN(n9750) );
  AOI22_X1 U10594 ( .A1(P2_REG3_REG_21__SCAN_IN), .A2(keyinput_109), .B1(n8068), .B2(keyinput_107), .ZN(n9748) );
  OAI221_X1 U10595 ( .B1(P2_REG3_REG_21__SCAN_IN), .B2(keyinput_109), .C1(
        n8068), .C2(keyinput_107), .A(n9748), .ZN(n9749) );
  AOI211_X1 U10596 ( .C1(n9752), .C2(n9751), .A(n9750), .B(n9749), .ZN(n9755)
         );
  NAND2_X1 U10597 ( .A1(n9754), .A2(keyinput_113), .ZN(n9753) );
  OAI221_X1 U10598 ( .B1(n9756), .B2(n9755), .C1(n9754), .C2(keyinput_113), 
        .A(n9753), .ZN(n9757) );
  OAI221_X1 U10599 ( .B1(P2_REG3_REG_17__SCAN_IN), .B2(n9759), .C1(n9758), 
        .C2(keyinput_114), .A(n9757), .ZN(n9760) );
  OAI221_X1 U10600 ( .B1(P2_REG3_REG_24__SCAN_IN), .B2(n9762), .C1(n9761), 
        .C2(keyinput_115), .A(n9760), .ZN(n9763) );
  AOI22_X1 U10601 ( .A1(n9764), .A2(n9763), .B1(keyinput_118), .B2(
        P2_REG3_REG_0__SCAN_IN), .ZN(n9765) );
  OAI21_X1 U10602 ( .B1(keyinput_118), .B2(P2_REG3_REG_0__SCAN_IN), .A(n9765), 
        .ZN(n9769) );
  AOI22_X1 U10603 ( .A1(P2_REG3_REG_22__SCAN_IN), .A2(keyinput_121), .B1(n9767), .B2(keyinput_122), .ZN(n9766) );
  OAI221_X1 U10604 ( .B1(P2_REG3_REG_22__SCAN_IN), .B2(keyinput_121), .C1(
        n9767), .C2(keyinput_122), .A(n9766), .ZN(n9768) );
  AOI21_X1 U10605 ( .B1(n9770), .B2(n9769), .A(n9768), .ZN(n9781) );
  OAI22_X1 U10606 ( .A1(n9773), .A2(keyinput_124), .B1(n9772), .B2(
        keyinput_123), .ZN(n9771) );
  AOI221_X1 U10607 ( .B1(n9773), .B2(keyinput_124), .C1(keyinput_123), .C2(
        n9772), .A(n9771), .ZN(n9778) );
  AOI22_X1 U10608 ( .A1(n6303), .A2(keyinput_125), .B1(keyinput_127), .B2(
        n9775), .ZN(n9774) );
  OAI221_X1 U10609 ( .B1(n6303), .B2(keyinput_125), .C1(n9775), .C2(
        keyinput_127), .A(n9774), .ZN(n9776) );
  AOI21_X1 U10610 ( .B1(keyinput_126), .B2(n9779), .A(n9776), .ZN(n9777) );
  OAI211_X1 U10611 ( .C1(keyinput_126), .C2(n9779), .A(n9778), .B(n9777), .ZN(
        n9780) );
  AOI211_X1 U10612 ( .C1(n9783), .C2(n9782), .A(n9781), .B(n9780), .ZN(n9784)
         );
  XOR2_X1 U10613 ( .A(n9785), .B(n9784), .Z(P1_U3572) );
  MUX2_X1 U10614 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n10053), .S(P1_U4006), .Z(
        P1_U3571) );
  MUX2_X1 U10615 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9786), .S(P1_U4006), .Z(
        P1_U3569) );
  MUX2_X1 U10616 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9787), .S(P1_U4006), .Z(
        P1_U3567) );
  MUX2_X1 U10617 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9788), .S(P1_U4006), .Z(
        P1_U3566) );
  MUX2_X1 U10618 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9789), .S(P1_U4006), .Z(
        P1_U3565) );
  MUX2_X1 U10619 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n10538), .S(P1_U4006), .Z(
        P1_U3564) );
  MUX2_X1 U10620 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9790), .S(P1_U4006), .Z(
        P1_U3563) );
  MUX2_X1 U10621 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9791), .S(P1_U4006), .Z(
        P1_U3560) );
  MUX2_X1 U10622 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n5029), .S(P1_U4006), .Z(
        P1_U3557) );
  MUX2_X1 U10623 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n7491), .S(P1_U4006), .Z(
        P1_U3556) );
  MUX2_X1 U10624 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n7380), .S(P1_U4006), .Z(
        P1_U3555) );
  NOR2_X1 U10625 ( .A1(n10342), .A2(n9794), .ZN(n9795) );
  AOI211_X1 U10626 ( .C1(n9810), .C2(n10339), .A(n9796), .B(n9795), .ZN(n9808)
         );
  AOI21_X1 U10627 ( .B1(P1_REG2_REG_14__SCAN_IN), .B2(n9798), .A(n9797), .ZN(
        n9821) );
  XNOR2_X1 U10628 ( .A(n9820), .B(n9821), .ZN(n9800) );
  INV_X1 U10629 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9799) );
  NOR2_X1 U10630 ( .A1(n9799), .A2(n9800), .ZN(n9822) );
  AOI211_X1 U10631 ( .C1(n9800), .C2(n9799), .A(n9822), .B(n10269), .ZN(n9801)
         );
  INV_X1 U10632 ( .A(n9801), .ZN(n9807) );
  INV_X1 U10633 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n9803) );
  AOI21_X1 U10634 ( .B1(n9804), .B2(n9803), .A(n9802), .ZN(n9809) );
  XNOR2_X1 U10635 ( .A(n9820), .B(n9809), .ZN(n9805) );
  NAND2_X1 U10636 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n9805), .ZN(n9811) );
  OAI211_X1 U10637 ( .C1(n9805), .C2(P1_REG1_REG_15__SCAN_IN), .A(n10349), .B(
        n9811), .ZN(n9806) );
  NAND3_X1 U10638 ( .A1(n9808), .A2(n9807), .A3(n9806), .ZN(P1_U3256) );
  NAND2_X1 U10639 ( .A1(n9810), .A2(n9809), .ZN(n9812) );
  NAND2_X1 U10640 ( .A1(n9812), .A2(n9811), .ZN(n9814) );
  XOR2_X1 U10641 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9840), .Z(n9813) );
  NAND2_X1 U10642 ( .A1(n9813), .A2(n9814), .ZN(n9829) );
  OAI211_X1 U10643 ( .C1(n9814), .C2(n9813), .A(n10349), .B(n9829), .ZN(n9818)
         );
  NOR2_X1 U10644 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9815), .ZN(n9816) );
  AOI21_X1 U10645 ( .B1(n10339), .B2(n9840), .A(n9816), .ZN(n9817) );
  OAI211_X1 U10646 ( .C1(n9819), .C2(n10342), .A(n9818), .B(n9817), .ZN(n9828)
         );
  NOR2_X1 U10647 ( .A1(n9821), .A2(n9820), .ZN(n9823) );
  NOR2_X1 U10648 ( .A1(n9823), .A2(n9822), .ZN(n9826) );
  NAND2_X1 U10649 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n9840), .ZN(n9824) );
  OAI21_X1 U10650 ( .B1(n9840), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9824), .ZN(
        n9825) );
  NOR2_X1 U10651 ( .A1(n9826), .A2(n9825), .ZN(n9839) );
  AOI211_X1 U10652 ( .C1(n9826), .C2(n9825), .A(n9839), .B(n10269), .ZN(n9827)
         );
  OR2_X1 U10653 ( .A1(n9828), .A2(n9827), .ZN(P1_U3257) );
  INV_X1 U10654 ( .A(n9849), .ZN(n9856) );
  XNOR2_X1 U10655 ( .A(n9856), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n9833) );
  INV_X1 U10656 ( .A(n9840), .ZN(n9831) );
  INV_X1 U10657 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9830) );
  OAI21_X1 U10658 ( .B1(n9831), .B2(n9830), .A(n9829), .ZN(n9832) );
  NAND2_X1 U10659 ( .A1(n9833), .A2(n9832), .ZN(n9854) );
  OAI211_X1 U10660 ( .C1(n9833), .C2(n9832), .A(n9854), .B(n10349), .ZN(n9835)
         );
  OAI211_X1 U10661 ( .C1(n9856), .C2(n9836), .A(n9835), .B(n9834), .ZN(n9845)
         );
  NOR2_X1 U10662 ( .A1(n10342), .A2(n9837), .ZN(n9844) );
  NAND2_X1 U10663 ( .A1(n9849), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9838) );
  OAI21_X1 U10664 ( .B1(n9849), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9838), .ZN(
        n9842) );
  AOI21_X1 U10665 ( .B1(n9840), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9839), .ZN(
        n9841) );
  NOR2_X1 U10666 ( .A1(n9841), .A2(n9842), .ZN(n9848) );
  AOI211_X1 U10667 ( .C1(n9842), .C2(n9841), .A(n9848), .B(n10269), .ZN(n9843)
         );
  OR3_X1 U10668 ( .A1(n9845), .A2(n9844), .A3(n9843), .ZN(P1_U3258) );
  INV_X1 U10669 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9846) );
  MUX2_X1 U10670 ( .A(P1_REG2_REG_18__SCAN_IN), .B(n9846), .S(n9872), .Z(n9847) );
  INV_X1 U10671 ( .A(n9847), .ZN(n9851) );
  AOI21_X1 U10672 ( .B1(n9849), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9848), .ZN(
        n9850) );
  NOR2_X1 U10673 ( .A1(n9850), .A2(n9851), .ZN(n9871) );
  AOI211_X1 U10674 ( .C1(n9851), .C2(n9850), .A(n9871), .B(n10269), .ZN(n9864)
         );
  INV_X1 U10675 ( .A(n9872), .ZN(n9853) );
  INV_X1 U10676 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9852) );
  NAND2_X1 U10677 ( .A1(n9853), .A2(n9852), .ZN(n9867) );
  OAI21_X1 U10678 ( .B1(n9853), .B2(n9852), .A(n9867), .ZN(n9858) );
  INV_X1 U10679 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9855) );
  OAI21_X1 U10680 ( .B1(n9856), .B2(n9855), .A(n9854), .ZN(n9857) );
  NOR2_X1 U10681 ( .A1(n9857), .A2(n9858), .ZN(n9865) );
  AOI21_X1 U10682 ( .B1(n9858), .B2(n9857), .A(n9865), .ZN(n9859) );
  NOR2_X1 U10683 ( .A1(n9859), .A2(n10299), .ZN(n9863) );
  INV_X1 U10684 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10254) );
  NAND2_X1 U10685 ( .A1(n9872), .A2(n10339), .ZN(n9861) );
  OAI211_X1 U10686 ( .C1(n10254), .C2(n10342), .A(n9861), .B(n9860), .ZN(n9862) );
  OR3_X1 U10687 ( .A1(n9864), .A2(n9863), .A3(n9862), .ZN(P1_U3259) );
  INV_X1 U10688 ( .A(n9865), .ZN(n9866) );
  NAND2_X1 U10689 ( .A1(n9867), .A2(n9866), .ZN(n9869) );
  XNOR2_X1 U10690 ( .A(n9991), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n9868) );
  XNOR2_X1 U10691 ( .A(n9869), .B(n9868), .ZN(n9881) );
  INV_X1 U10692 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n9870) );
  MUX2_X1 U10693 ( .A(n9870), .B(P1_REG2_REG_19__SCAN_IN), .S(n9991), .Z(n9874) );
  AOI21_X1 U10694 ( .B1(n9872), .B2(P1_REG2_REG_18__SCAN_IN), .A(n9871), .ZN(
        n9873) );
  XOR2_X1 U10695 ( .A(n9874), .B(n9873), .Z(n9879) );
  NAND2_X1 U10696 ( .A1(n10339), .A2(n9991), .ZN(n9876) );
  OAI211_X1 U10697 ( .C1(n10342), .C2(n9877), .A(n9876), .B(n9875), .ZN(n9878)
         );
  AOI21_X1 U10698 ( .B1(n9879), .B2(n10335), .A(n9878), .ZN(n9880) );
  OAI21_X1 U10699 ( .B1(n10299), .B2(n9881), .A(n9880), .ZN(P1_U3260) );
  NAND2_X1 U10700 ( .A1(n9889), .A2(n9888), .ZN(n9887) );
  XNOR2_X1 U10701 ( .A(n5579), .B(n9887), .ZN(n10065) );
  NAND2_X1 U10702 ( .A1(n10065), .A2(n10558), .ZN(n9886) );
  NAND2_X1 U10703 ( .A1(n9884), .A2(n9883), .ZN(n10069) );
  NOR2_X1 U10704 ( .A1(n10069), .A2(n10563), .ZN(n9891) );
  AOI21_X1 U10705 ( .B1(n9977), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9891), .ZN(
        n9885) );
  OAI211_X1 U10706 ( .C1(n5579), .C2(n10565), .A(n9886), .B(n9885), .ZN(
        P1_U3261) );
  OAI21_X1 U10707 ( .B1(n9889), .B2(n9888), .A(n9887), .ZN(n10070) );
  NOR2_X1 U10708 ( .A1(n10568), .A2(n9890), .ZN(n9892) );
  AOI211_X1 U10709 ( .C1(n10067), .C2(n10042), .A(n9892), .B(n9891), .ZN(n9893) );
  OAI21_X1 U10710 ( .B1(n10070), .B2(n10046), .A(n9893), .ZN(P1_U3262) );
  AOI21_X1 U10711 ( .B1(n9896), .B2(n9895), .A(n9894), .ZN(n10075) );
  XNOR2_X1 U10712 ( .A(n9897), .B(n9896), .ZN(n9901) );
  OAI22_X1 U10713 ( .A1(n9899), .A2(n10489), .B1(n9898), .B2(n7059), .ZN(n9900) );
  AOI21_X1 U10714 ( .B1(n9901), .B2(n10546), .A(n9900), .ZN(n10079) );
  OAI22_X1 U10715 ( .A1(n9903), .A2(n10005), .B1(n9902), .B2(n10568), .ZN(
        n9904) );
  AOI21_X1 U10716 ( .B1(n10076), .B2(n10042), .A(n9904), .ZN(n9909) );
  NAND2_X1 U10717 ( .A1(n10076), .A2(n9905), .ZN(n9906) );
  AND2_X1 U10718 ( .A1(n9907), .A2(n9906), .ZN(n10077) );
  NAND2_X1 U10719 ( .A1(n10077), .A2(n10558), .ZN(n9908) );
  OAI211_X1 U10720 ( .C1(n10079), .C2(n9977), .A(n9909), .B(n9908), .ZN(n9910)
         );
  AOI21_X1 U10721 ( .B1(n10075), .B2(n9911), .A(n9910), .ZN(n9912) );
  INV_X1 U10722 ( .A(n9912), .ZN(P1_U3263) );
  INV_X1 U10723 ( .A(n9913), .ZN(n9914) );
  AOI21_X1 U10724 ( .B1(n9921), .B2(n9915), .A(n9914), .ZN(n10095) );
  AOI211_X1 U10725 ( .C1(n10092), .C2(n9941), .A(n10582), .B(n9916), .ZN(
        n10091) );
  INV_X1 U10726 ( .A(n10092), .ZN(n9919) );
  AOI22_X1 U10727 ( .A1(n9917), .A2(n10561), .B1(P1_REG2_REG_25__SCAN_IN), 
        .B2(n10563), .ZN(n9918) );
  OAI21_X1 U10728 ( .B1(n9919), .B2(n10565), .A(n9918), .ZN(n9926) );
  OAI21_X1 U10729 ( .B1(n9922), .B2(n9921), .A(n9920), .ZN(n9924) );
  AOI222_X1 U10730 ( .A1(n10546), .A2(n9924), .B1(n9954), .B2(n10540), .C1(
        n9923), .C2(n10539), .ZN(n10094) );
  NOR2_X1 U10731 ( .A1(n10094), .A2(n10563), .ZN(n9925) );
  AOI211_X1 U10732 ( .C1(n10091), .C2(n10026), .A(n9926), .B(n9925), .ZN(n9927) );
  OAI21_X1 U10733 ( .B1(n10095), .B2(n10028), .A(n9927), .ZN(P1_U3266) );
  XOR2_X1 U10734 ( .A(n9929), .B(n9928), .Z(n9931) );
  AOI222_X1 U10735 ( .A1(n10546), .A2(n9931), .B1(n9969), .B2(n10540), .C1(
        n9930), .C2(n10539), .ZN(n10099) );
  AND2_X1 U10736 ( .A1(n9933), .A2(n9932), .ZN(n9936) );
  OAI21_X1 U10737 ( .B1(n9936), .B2(n9935), .A(n9934), .ZN(n10100) );
  OAI22_X1 U10738 ( .A1(n9938), .A2(n10005), .B1(n9937), .B2(n10568), .ZN(
        n9939) );
  AOI21_X1 U10739 ( .B1(n10097), .B2(n10042), .A(n9939), .ZN(n9943) );
  NAND2_X1 U10740 ( .A1(n5008), .A2(n10097), .ZN(n9940) );
  AND3_X1 U10741 ( .A1(n9941), .A2(n9940), .A3(n10366), .ZN(n10096) );
  NAND2_X1 U10742 ( .A1(n10096), .A2(n10026), .ZN(n9942) );
  OAI211_X1 U10743 ( .C1(n10100), .C2(n10028), .A(n9943), .B(n9942), .ZN(n9944) );
  INV_X1 U10744 ( .A(n9944), .ZN(n9945) );
  OAI21_X1 U10745 ( .B1(n9977), .B2(n10099), .A(n9945), .ZN(P1_U3267) );
  XOR2_X1 U10746 ( .A(n9946), .B(n9952), .Z(n10105) );
  AOI211_X1 U10747 ( .C1(n10102), .C2(n9961), .A(n10582), .B(n9947), .ZN(
        n10101) );
  INV_X1 U10748 ( .A(n9948), .ZN(n9949) );
  AOI22_X1 U10749 ( .A1(n9949), .A2(n10561), .B1(P1_REG2_REG_23__SCAN_IN), 
        .B2(n10563), .ZN(n9950) );
  OAI21_X1 U10750 ( .B1(n9951), .B2(n10565), .A(n9950), .ZN(n9958) );
  XNOR2_X1 U10751 ( .A(n9953), .B(n9952), .ZN(n9956) );
  AOI222_X1 U10752 ( .A1(n10546), .A2(n9956), .B1(n9955), .B2(n10540), .C1(
        n9954), .C2(n10539), .ZN(n10104) );
  NOR2_X1 U10753 ( .A1(n10104), .A2(n10563), .ZN(n9957) );
  AOI211_X1 U10754 ( .C1(n10101), .C2(n10026), .A(n9958), .B(n9957), .ZN(n9959) );
  OAI21_X1 U10755 ( .B1(n10105), .B2(n10028), .A(n9959), .ZN(P1_U3268) );
  XOR2_X1 U10756 ( .A(n9960), .B(n9967), .Z(n10110) );
  INV_X1 U10757 ( .A(n9961), .ZN(n9962) );
  AOI21_X1 U10758 ( .B1(n10106), .B2(n9978), .A(n9962), .ZN(n10107) );
  INV_X1 U10759 ( .A(n10106), .ZN(n9966) );
  INV_X1 U10760 ( .A(n9963), .ZN(n9964) );
  AOI22_X1 U10761 ( .A1(n9964), .A2(n10561), .B1(P1_REG2_REG_22__SCAN_IN), 
        .B2(n10563), .ZN(n9965) );
  OAI21_X1 U10762 ( .B1(n9966), .B2(n10565), .A(n9965), .ZN(n9973) );
  XNOR2_X1 U10763 ( .A(n9968), .B(n9967), .ZN(n9971) );
  AOI222_X1 U10764 ( .A1(n10546), .A2(n9971), .B1(n9970), .B2(n10540), .C1(
        n9969), .C2(n10539), .ZN(n10109) );
  NOR2_X1 U10765 ( .A1(n10109), .A2(n9977), .ZN(n9972) );
  AOI211_X1 U10766 ( .C1(n10107), .C2(n10558), .A(n9973), .B(n9972), .ZN(n9974) );
  OAI21_X1 U10767 ( .B1(n10028), .B2(n10110), .A(n9974), .ZN(P1_U3269) );
  OAI21_X1 U10768 ( .B1(n9976), .B2(n9983), .A(n9975), .ZN(n10116) );
  AOI22_X1 U10769 ( .A1(n10113), .A2(n10042), .B1(n9977), .B2(
        P1_REG2_REG_21__SCAN_IN), .ZN(n9994) );
  INV_X1 U10770 ( .A(n9995), .ZN(n9980) );
  INV_X1 U10771 ( .A(n9978), .ZN(n9979) );
  AOI211_X1 U10772 ( .C1(n10113), .C2(n9980), .A(n10582), .B(n9979), .ZN(
        n10111) );
  INV_X1 U10773 ( .A(n10111), .ZN(n9990) );
  NAND2_X1 U10774 ( .A1(n9982), .A2(n9981), .ZN(n9984) );
  XNOR2_X1 U10775 ( .A(n9984), .B(n9983), .ZN(n9985) );
  AOI22_X1 U10776 ( .A1(n9985), .A2(n10546), .B1(n10540), .B2(n10022), .ZN(
        n10115) );
  INV_X1 U10777 ( .A(n9986), .ZN(n9988) );
  NOR2_X1 U10778 ( .A1(n9987), .A2(n10489), .ZN(n10112) );
  AOI21_X1 U10779 ( .B1(n10561), .B2(n9988), .A(n10112), .ZN(n9989) );
  OAI211_X1 U10780 ( .C1(n9991), .C2(n9990), .A(n10115), .B(n9989), .ZN(n9992)
         );
  NAND2_X1 U10781 ( .A1(n9992), .A2(n10568), .ZN(n9993) );
  OAI211_X1 U10782 ( .C1(n10116), .C2(n10028), .A(n9994), .B(n9993), .ZN(
        P1_U3270) );
  AOI21_X1 U10783 ( .B1(n10117), .B2(n10013), .A(n9995), .ZN(n10118) );
  INV_X1 U10784 ( .A(n10118), .ZN(n10011) );
  XNOR2_X1 U10785 ( .A(n9996), .B(n9997), .ZN(n10121) );
  AOI21_X1 U10786 ( .B1(n10550), .B2(n9998), .A(n10121), .ZN(n10004) );
  XNOR2_X1 U10787 ( .A(n9999), .B(n5197), .ZN(n10002) );
  OAI22_X1 U10788 ( .A1(n10000), .A2(n10489), .B1(n10036), .B2(n7059), .ZN(
        n10001) );
  AOI21_X1 U10789 ( .B1(n10002), .B2(n10546), .A(n10001), .ZN(n10120) );
  INV_X1 U10790 ( .A(n10120), .ZN(n10003) );
  OAI21_X1 U10791 ( .B1(n10004), .B2(n10003), .A(n10568), .ZN(n10010) );
  OAI22_X1 U10792 ( .A1(n10568), .A2(n10007), .B1(n10006), .B2(n10005), .ZN(
        n10008) );
  AOI21_X1 U10793 ( .B1(n10117), .B2(n10042), .A(n10008), .ZN(n10009) );
  OAI211_X1 U10794 ( .C1(n10011), .C2(n10046), .A(n10010), .B(n10009), .ZN(
        P1_U3271) );
  XOR2_X1 U10795 ( .A(n10012), .B(n10021), .Z(n10126) );
  INV_X1 U10796 ( .A(n10039), .ZN(n10015) );
  INV_X1 U10797 ( .A(n10013), .ZN(n10014) );
  AOI211_X1 U10798 ( .C1(n10123), .C2(n10015), .A(n10582), .B(n10014), .ZN(
        n10122) );
  AOI22_X1 U10799 ( .A1(n10563), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n10016), 
        .B2(n10561), .ZN(n10017) );
  OAI21_X1 U10800 ( .B1(n10018), .B2(n10565), .A(n10017), .ZN(n10025) );
  OAI21_X1 U10801 ( .B1(n10021), .B2(n10020), .A(n10019), .ZN(n10023) );
  AOI222_X1 U10802 ( .A1(n10546), .A2(n10023), .B1(n10022), .B2(n10539), .C1(
        n10052), .C2(n10540), .ZN(n10125) );
  NOR2_X1 U10803 ( .A1(n10125), .A2(n10563), .ZN(n10024) );
  AOI211_X1 U10804 ( .C1(n10122), .C2(n10026), .A(n10025), .B(n10024), .ZN(
        n10027) );
  OAI21_X1 U10805 ( .B1(n10028), .B2(n10126), .A(n10027), .ZN(P1_U3272) );
  XNOR2_X1 U10806 ( .A(n10029), .B(n10030), .ZN(n10127) );
  NAND2_X1 U10807 ( .A1(n10031), .A2(n10032), .ZN(n10033) );
  AOI21_X1 U10808 ( .B1(n10034), .B2(n10033), .A(n7060), .ZN(n10038) );
  OAI22_X1 U10809 ( .A1(n10036), .A2(n10489), .B1(n10035), .B2(n7059), .ZN(
        n10037) );
  AOI211_X1 U10810 ( .C1(n10127), .C2(n10522), .A(n10038), .B(n10037), .ZN(
        n10132) );
  AND2_X1 U10811 ( .A1(n10057), .A2(n10043), .ZN(n10040) );
  OR2_X1 U10812 ( .A1(n10040), .A2(n10039), .ZN(n10129) );
  AOI22_X1 U10813 ( .A1(n10563), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n10041), 
        .B2(n10561), .ZN(n10045) );
  NAND2_X1 U10814 ( .A1(n10043), .A2(n10042), .ZN(n10044) );
  OAI211_X1 U10815 ( .C1(n10129), .C2(n10046), .A(n10045), .B(n10044), .ZN(
        n10047) );
  AOI21_X1 U10816 ( .B1(n10127), .B2(n10559), .A(n10047), .ZN(n10048) );
  OAI21_X1 U10817 ( .B1(n10132), .B2(n9977), .A(n10048), .ZN(P1_U3273) );
  XNOR2_X1 U10818 ( .A(n10049), .B(n10050), .ZN(n10134) );
  XNOR2_X1 U10819 ( .A(n10051), .B(n10050), .ZN(n10055) );
  AOI22_X1 U10820 ( .A1(n10540), .A2(n10053), .B1(n10052), .B2(n10539), .ZN(
        n10054) );
  OAI21_X1 U10821 ( .B1(n10055), .B2(n7060), .A(n10054), .ZN(n10056) );
  AOI21_X1 U10822 ( .B1(n10134), .B2(n10522), .A(n10056), .ZN(n10138) );
  INV_X1 U10823 ( .A(n10057), .ZN(n10058) );
  AOI21_X1 U10824 ( .B1(n10135), .B2(n10059), .A(n10058), .ZN(n10136) );
  NAND2_X1 U10825 ( .A1(n10136), .A2(n10558), .ZN(n10062) );
  AOI22_X1 U10826 ( .A1(n10563), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n10060), 
        .B2(n10561), .ZN(n10061) );
  OAI211_X1 U10827 ( .C1(n7061), .C2(n10565), .A(n10062), .B(n10061), .ZN(
        n10063) );
  AOI21_X1 U10828 ( .B1(n10134), .B2(n10559), .A(n10063), .ZN(n10064) );
  OAI21_X1 U10829 ( .B1(n10138), .B2(n9977), .A(n10064), .ZN(P1_U3274) );
  NAND2_X1 U10830 ( .A1(n10065), .A2(n10366), .ZN(n10066) );
  OAI211_X1 U10831 ( .C1(n5579), .C2(n10581), .A(n10066), .B(n10069), .ZN(
        n10173) );
  MUX2_X1 U10832 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n10173), .S(n10590), .Z(
        P1_U3554) );
  NAND2_X1 U10833 ( .A1(n10067), .A2(n10365), .ZN(n10068) );
  OAI211_X1 U10834 ( .C1(n10070), .C2(n10582), .A(n10069), .B(n10068), .ZN(
        n10174) );
  MUX2_X1 U10835 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n10174), .S(n10590), .Z(
        P1_U3553) );
  MUX2_X1 U10836 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n10175), .S(n10590), .Z(
        P1_U3552) );
  INV_X1 U10837 ( .A(n10075), .ZN(n10080) );
  AOI22_X1 U10838 ( .A1(n10077), .A2(n10366), .B1(n10365), .B2(n10076), .ZN(
        n10078) );
  OAI211_X1 U10839 ( .C1(n10080), .C2(n10460), .A(n10079), .B(n10078), .ZN(
        n10176) );
  MUX2_X1 U10840 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n10176), .S(n10590), .Z(
        P1_U3551) );
  AOI21_X1 U10841 ( .B1(n10365), .B2(n10082), .A(n10081), .ZN(n10083) );
  MUX2_X1 U10842 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n10177), .S(n10590), .Z(
        P1_U3550) );
  AOI22_X1 U10843 ( .A1(n10087), .A2(n10366), .B1(n10365), .B2(n10086), .ZN(
        n10088) );
  OAI211_X1 U10844 ( .C1(n10090), .C2(n10370), .A(n10089), .B(n10088), .ZN(
        n10178) );
  MUX2_X1 U10845 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n10178), .S(n10590), .Z(
        P1_U3549) );
  AOI21_X1 U10846 ( .B1(n10365), .B2(n10092), .A(n10091), .ZN(n10093) );
  OAI211_X1 U10847 ( .C1(n10095), .C2(n10460), .A(n10094), .B(n10093), .ZN(
        n10179) );
  MUX2_X1 U10848 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n10179), .S(n10590), .Z(
        P1_U3548) );
  AOI21_X1 U10849 ( .B1(n10365), .B2(n10097), .A(n10096), .ZN(n10098) );
  OAI211_X1 U10850 ( .C1(n10100), .C2(n10460), .A(n10099), .B(n10098), .ZN(
        n10180) );
  MUX2_X1 U10851 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n10180), .S(n10590), .Z(
        P1_U3547) );
  AOI21_X1 U10852 ( .B1(n10365), .B2(n10102), .A(n10101), .ZN(n10103) );
  OAI211_X1 U10853 ( .C1(n10105), .C2(n10460), .A(n10104), .B(n10103), .ZN(
        n10181) );
  MUX2_X1 U10854 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n10181), .S(n10590), .Z(
        P1_U3546) );
  AOI22_X1 U10855 ( .A1(n10107), .A2(n10366), .B1(n10365), .B2(n10106), .ZN(
        n10108) );
  OAI211_X1 U10856 ( .C1(n10110), .C2(n10460), .A(n10109), .B(n10108), .ZN(
        n10182) );
  MUX2_X1 U10857 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n10182), .S(n10590), .Z(
        P1_U3545) );
  AOI211_X1 U10858 ( .C1(n10365), .C2(n10113), .A(n10112), .B(n10111), .ZN(
        n10114) );
  OAI211_X1 U10859 ( .C1(n10116), .C2(n10460), .A(n10115), .B(n10114), .ZN(
        n10183) );
  MUX2_X1 U10860 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n10183), .S(n10590), .Z(
        P1_U3544) );
  AOI22_X1 U10861 ( .A1(n10118), .A2(n10366), .B1(n10365), .B2(n10117), .ZN(
        n10119) );
  OAI211_X1 U10862 ( .C1(n10121), .C2(n10460), .A(n10120), .B(n10119), .ZN(
        n10184) );
  MUX2_X1 U10863 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n10184), .S(n10590), .Z(
        P1_U3543) );
  AOI21_X1 U10864 ( .B1(n10365), .B2(n10123), .A(n10122), .ZN(n10124) );
  OAI211_X1 U10865 ( .C1(n10126), .C2(n10460), .A(n10125), .B(n10124), .ZN(
        n10185) );
  MUX2_X1 U10866 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n10185), .S(n10590), .Z(
        P1_U3542) );
  INV_X1 U10867 ( .A(n10127), .ZN(n10133) );
  OAI22_X1 U10868 ( .A1(n10129), .A2(n10582), .B1(n10128), .B2(n10581), .ZN(
        n10130) );
  INV_X1 U10869 ( .A(n10130), .ZN(n10131) );
  OAI211_X1 U10870 ( .C1(n10370), .C2(n10133), .A(n10132), .B(n10131), .ZN(
        n10186) );
  MUX2_X1 U10871 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n10186), .S(n10590), .Z(
        P1_U3541) );
  INV_X1 U10872 ( .A(n10134), .ZN(n10139) );
  AOI22_X1 U10873 ( .A1(n10136), .A2(n10366), .B1(n10365), .B2(n10135), .ZN(
        n10137) );
  OAI211_X1 U10874 ( .C1(n10370), .C2(n10139), .A(n10138), .B(n10137), .ZN(
        n10187) );
  MUX2_X1 U10875 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n10187), .S(n10590), .Z(
        P1_U3540) );
  AOI21_X1 U10876 ( .B1(n10365), .B2(n10141), .A(n10140), .ZN(n10142) );
  OAI211_X1 U10877 ( .C1(n10144), .C2(n10460), .A(n10143), .B(n10142), .ZN(
        n10188) );
  MUX2_X1 U10878 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n10188), .S(n10590), .Z(
        P1_U3539) );
  INV_X1 U10879 ( .A(n10145), .ZN(n10150) );
  AOI22_X1 U10880 ( .A1(n10147), .A2(n10366), .B1(n10365), .B2(n10146), .ZN(
        n10148) );
  OAI211_X1 U10881 ( .C1(n10370), .C2(n10150), .A(n10149), .B(n10148), .ZN(
        n10189) );
  MUX2_X1 U10882 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n10189), .S(n10590), .Z(
        P1_U3538) );
  AOI21_X1 U10883 ( .B1(n10365), .B2(n10152), .A(n10151), .ZN(n10153) );
  OAI211_X1 U10884 ( .C1(n10155), .C2(n10460), .A(n10154), .B(n10153), .ZN(
        n10190) );
  MUX2_X1 U10885 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n10190), .S(n10590), .Z(
        P1_U3537) );
  INV_X1 U10886 ( .A(n10156), .ZN(n10161) );
  AOI22_X1 U10887 ( .A1(n10158), .A2(n10366), .B1(n10365), .B2(n10157), .ZN(
        n10159) );
  OAI211_X1 U10888 ( .C1(n10161), .C2(n10460), .A(n10160), .B(n10159), .ZN(
        n10191) );
  MUX2_X1 U10889 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n10191), .S(n10590), .Z(
        P1_U3536) );
  AOI21_X1 U10890 ( .B1(n10365), .B2(n10163), .A(n10162), .ZN(n10164) );
  OAI211_X1 U10891 ( .C1(n10166), .C2(n10460), .A(n10165), .B(n10164), .ZN(
        n10192) );
  MUX2_X1 U10892 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n10192), .S(n10590), .Z(
        P1_U3535) );
  INV_X1 U10893 ( .A(n10167), .ZN(n10172) );
  AOI22_X1 U10894 ( .A1(n10169), .A2(n10366), .B1(n10365), .B2(n10168), .ZN(
        n10170) );
  OAI211_X1 U10895 ( .C1(n10172), .C2(n10370), .A(n10171), .B(n10170), .ZN(
        n10193) );
  MUX2_X1 U10896 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n10193), .S(n10590), .Z(
        P1_U3534) );
  MUX2_X1 U10897 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n10173), .S(n10594), .Z(
        P1_U3522) );
  MUX2_X1 U10898 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n10174), .S(n10594), .Z(
        P1_U3521) );
  MUX2_X1 U10899 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n10175), .S(n10594), .Z(
        P1_U3520) );
  MUX2_X1 U10900 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n10176), .S(n10594), .Z(
        P1_U3519) );
  MUX2_X1 U10901 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n10177), .S(n10594), .Z(
        P1_U3518) );
  MUX2_X1 U10902 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n10178), .S(n10594), .Z(
        P1_U3517) );
  MUX2_X1 U10903 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n10179), .S(n10594), .Z(
        P1_U3516) );
  MUX2_X1 U10904 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n10180), .S(n10594), .Z(
        P1_U3515) );
  MUX2_X1 U10905 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n10181), .S(n10594), .Z(
        P1_U3514) );
  MUX2_X1 U10906 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n10182), .S(n10594), .Z(
        P1_U3513) );
  MUX2_X1 U10907 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n10183), .S(n10594), .Z(
        P1_U3512) );
  MUX2_X1 U10908 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n10184), .S(n10594), .Z(
        P1_U3511) );
  MUX2_X1 U10909 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n10185), .S(n10594), .Z(
        P1_U3510) );
  MUX2_X1 U10910 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n10186), .S(n10594), .Z(
        P1_U3508) );
  MUX2_X1 U10911 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n10187), .S(n10594), .Z(
        P1_U3505) );
  MUX2_X1 U10912 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n10188), .S(n10594), .Z(
        P1_U3502) );
  MUX2_X1 U10913 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n10189), .S(n10594), .Z(
        P1_U3499) );
  MUX2_X1 U10914 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n10190), .S(n10594), .Z(
        P1_U3496) );
  MUX2_X1 U10915 ( .A(P1_REG0_REG_13__SCAN_IN), .B(n10191), .S(n10594), .Z(
        P1_U3493) );
  MUX2_X1 U10916 ( .A(P1_REG0_REG_12__SCAN_IN), .B(n10192), .S(n10594), .Z(
        P1_U3490) );
  MUX2_X1 U10917 ( .A(P1_REG0_REG_11__SCAN_IN), .B(n10193), .S(n10594), .Z(
        P1_U3487) );
  MUX2_X1 U10918 ( .A(n10194), .B(P1_D_REG_0__SCAN_IN), .S(n10211), .Z(
        P1_U3440) );
  NAND3_X1 U10919 ( .A1(n10195), .A2(P1_STATE_REG_SCAN_IN), .A3(
        P1_IR_REG_31__SCAN_IN), .ZN(n10198) );
  OAI22_X1 U10920 ( .A1(n5560), .A2(n10198), .B1(n10197), .B2(n10196), .ZN(
        n10199) );
  AOI21_X1 U10921 ( .B1(n9369), .B2(n10204), .A(n10199), .ZN(n10200) );
  INV_X1 U10922 ( .A(n10200), .ZN(P1_U3322) );
  NAND2_X1 U10923 ( .A1(n6582), .A2(n10204), .ZN(n10202) );
  OAI211_X1 U10924 ( .C1(n10209), .C2(n10203), .A(n10202), .B(n10201), .ZN(
        P1_U3325) );
  NAND2_X1 U10925 ( .A1(n10205), .A2(n10204), .ZN(n10207) );
  OAI211_X1 U10926 ( .C1(n10209), .C2(n10208), .A(n10207), .B(n10206), .ZN(
        P1_U3326) );
  MUX2_X1 U10927 ( .A(n10210), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  AND2_X1 U10928 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n10211), .ZN(P1_U3321) );
  AND2_X1 U10929 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n10211), .ZN(P1_U3320) );
  AND2_X1 U10930 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n10211), .ZN(P1_U3319) );
  AND2_X1 U10931 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n10211), .ZN(P1_U3318) );
  AND2_X1 U10932 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n10211), .ZN(P1_U3317) );
  AND2_X1 U10933 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n10211), .ZN(P1_U3316) );
  AND2_X1 U10934 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n10211), .ZN(P1_U3315) );
  AND2_X1 U10935 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n10211), .ZN(P1_U3314) );
  AND2_X1 U10936 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n10211), .ZN(P1_U3313) );
  AND2_X1 U10937 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n10211), .ZN(P1_U3312) );
  AND2_X1 U10938 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n10211), .ZN(P1_U3311) );
  AND2_X1 U10939 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n10211), .ZN(P1_U3310) );
  AND2_X1 U10940 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n10211), .ZN(P1_U3309) );
  AND2_X1 U10941 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n10211), .ZN(P1_U3308) );
  AND2_X1 U10942 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n10211), .ZN(P1_U3307) );
  AND2_X1 U10943 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n10211), .ZN(P1_U3306) );
  AND2_X1 U10944 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n10211), .ZN(P1_U3305) );
  AND2_X1 U10945 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n10211), .ZN(P1_U3304) );
  AND2_X1 U10946 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n10211), .ZN(P1_U3303) );
  AND2_X1 U10947 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n10211), .ZN(P1_U3302) );
  AND2_X1 U10948 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n10211), .ZN(P1_U3301) );
  AND2_X1 U10949 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n10211), .ZN(P1_U3300) );
  AND2_X1 U10950 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n10211), .ZN(P1_U3299) );
  AND2_X1 U10951 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n10211), .ZN(P1_U3298) );
  AND2_X1 U10952 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n10211), .ZN(P1_U3297) );
  AND2_X1 U10953 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n10211), .ZN(P1_U3296) );
  AND2_X1 U10954 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n10211), .ZN(P1_U3295) );
  AND2_X1 U10955 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n10211), .ZN(P1_U3294) );
  AND2_X1 U10956 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n10211), .ZN(P1_U3293) );
  AND2_X1 U10957 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n10211), .ZN(P1_U3292) );
  INV_X1 U10958 ( .A(n10212), .ZN(n10214) );
  AOI22_X1 U10959 ( .A1(n10216), .A2(n10309), .B1(n10312), .B2(n10215), .ZN(
        P2_U3438) );
  AND2_X1 U10960 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n10309), .ZN(P2_U3326) );
  AND2_X1 U10961 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n10309), .ZN(P2_U3325) );
  AND2_X1 U10962 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n10309), .ZN(P2_U3324) );
  AND2_X1 U10963 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n10309), .ZN(P2_U3323) );
  AND2_X1 U10964 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n10309), .ZN(P2_U3322) );
  AND2_X1 U10965 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n10309), .ZN(P2_U3321) );
  AND2_X1 U10966 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n10309), .ZN(P2_U3320) );
  AND2_X1 U10967 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n10309), .ZN(P2_U3319) );
  AND2_X1 U10968 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n10309), .ZN(P2_U3318) );
  AND2_X1 U10969 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n10309), .ZN(P2_U3317) );
  AND2_X1 U10970 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n10309), .ZN(P2_U3316) );
  AND2_X1 U10971 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n10309), .ZN(P2_U3315) );
  AND2_X1 U10972 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n10309), .ZN(P2_U3314) );
  AND2_X1 U10973 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n10309), .ZN(P2_U3313) );
  AND2_X1 U10974 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n10309), .ZN(P2_U3312) );
  AND2_X1 U10975 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n10309), .ZN(P2_U3311) );
  AND2_X1 U10976 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n10309), .ZN(P2_U3310) );
  AND2_X1 U10977 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n10309), .ZN(P2_U3309) );
  AND2_X1 U10978 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n10309), .ZN(P2_U3308) );
  AND2_X1 U10979 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n10309), .ZN(P2_U3307) );
  AND2_X1 U10980 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n10309), .ZN(P2_U3306) );
  AND2_X1 U10981 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n10309), .ZN(P2_U3305) );
  AND2_X1 U10982 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n10309), .ZN(P2_U3304) );
  AND2_X1 U10983 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n10309), .ZN(P2_U3303) );
  AND2_X1 U10984 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n10309), .ZN(P2_U3302) );
  AND2_X1 U10985 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n10309), .ZN(P2_U3301) );
  AND2_X1 U10986 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n10309), .ZN(P2_U3300) );
  AND2_X1 U10987 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n10309), .ZN(P2_U3299) );
  AND2_X1 U10988 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n10309), .ZN(P2_U3298) );
  AND2_X1 U10989 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n10309), .ZN(P2_U3297) );
  XOR2_X1 U10990 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(P1_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  INV_X1 U10991 ( .A(n10217), .ZN(n10218) );
  NAND2_X1 U10992 ( .A1(n10219), .A2(n10218), .ZN(n10220) );
  XOR2_X1 U10993 ( .A(n10221), .B(n10220), .Z(ADD_1071_U5) );
  XOR2_X1 U10994 ( .A(n10223), .B(n10222), .Z(ADD_1071_U54) );
  XOR2_X1 U10995 ( .A(n10225), .B(n10224), .Z(ADD_1071_U53) );
  XNOR2_X1 U10996 ( .A(n10227), .B(n10226), .ZN(ADD_1071_U52) );
  NOR2_X1 U10997 ( .A1(n10229), .A2(n10228), .ZN(n10230) );
  XOR2_X1 U10998 ( .A(n10230), .B(P2_ADDR_REG_5__SCAN_IN), .Z(ADD_1071_U51) );
  XOR2_X1 U10999 ( .A(n10231), .B(P2_ADDR_REG_6__SCAN_IN), .Z(ADD_1071_U50) );
  XOR2_X1 U11000 ( .A(n10232), .B(P2_ADDR_REG_7__SCAN_IN), .Z(ADD_1071_U49) );
  XOR2_X1 U11001 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n10233), .Z(ADD_1071_U48) );
  XOR2_X1 U11002 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n10234), .Z(ADD_1071_U47) );
  XOR2_X1 U11003 ( .A(n10236), .B(n10235), .Z(ADD_1071_U63) );
  XOR2_X1 U11004 ( .A(n10238), .B(n10237), .Z(ADD_1071_U62) );
  XNOR2_X1 U11005 ( .A(n10240), .B(n10239), .ZN(ADD_1071_U61) );
  XNOR2_X1 U11006 ( .A(n10242), .B(n10241), .ZN(ADD_1071_U60) );
  XNOR2_X1 U11007 ( .A(n10244), .B(n10243), .ZN(ADD_1071_U59) );
  XNOR2_X1 U11008 ( .A(n10246), .B(n10245), .ZN(ADD_1071_U58) );
  XNOR2_X1 U11009 ( .A(n10248), .B(n10247), .ZN(ADD_1071_U57) );
  XNOR2_X1 U11010 ( .A(n10250), .B(n10249), .ZN(ADD_1071_U56) );
  NOR2_X1 U11011 ( .A1(n10252), .A2(n10251), .ZN(n10253) );
  XNOR2_X1 U11012 ( .A(n10254), .B(n10253), .ZN(ADD_1071_U55) );
  INV_X1 U11013 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n10266) );
  OAI211_X1 U11014 ( .C1(n10259), .C2(n10255), .A(P1_STATE_REG_SCAN_IN), .B(
        n4854), .ZN(n10258) );
  INV_X1 U11015 ( .A(n10256), .ZN(n10257) );
  OAI22_X1 U11016 ( .A1(n10299), .A2(P1_REG1_REG_0__SCAN_IN), .B1(n10258), 
        .B2(n10257), .ZN(n10264) );
  AOI21_X1 U11017 ( .B1(n10261), .B2(n10260), .A(n10259), .ZN(n10262) );
  OR2_X1 U11018 ( .A1(n10262), .A2(P1_IR_REG_0__SCAN_IN), .ZN(n10263) );
  AOI22_X1 U11019 ( .A1(n10264), .A2(n10263), .B1(n10294), .B2(
        P1_ADDR_REG_0__SCAN_IN), .ZN(n10265) );
  OAI21_X1 U11020 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n10266), .A(n10265), .ZN(
        P1_U3241) );
  AOI22_X1 U11021 ( .A1(n10294), .A2(P1_ADDR_REG_6__SCAN_IN), .B1(n10339), 
        .B2(n10267), .ZN(n10280) );
  AOI211_X1 U11022 ( .C1(n10271), .C2(n10270), .A(n10269), .B(n10268), .ZN(
        n10272) );
  INV_X1 U11023 ( .A(n10272), .ZN(n10278) );
  AOI211_X1 U11024 ( .C1(n10275), .C2(n10274), .A(n10299), .B(n10273), .ZN(
        n10276) );
  INV_X1 U11025 ( .A(n10276), .ZN(n10277) );
  NAND4_X1 U11026 ( .A1(n10280), .A2(n10279), .A3(n10278), .A4(n10277), .ZN(
        P1_U3247) );
  AOI22_X1 U11027 ( .A1(n10294), .A2(P1_ADDR_REG_9__SCAN_IN), .B1(n10339), 
        .B2(n10281), .ZN(n10292) );
  NAND2_X1 U11028 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3084), .ZN(n10291) );
  OAI211_X1 U11029 ( .C1(n10284), .C2(n10283), .A(n10335), .B(n10282), .ZN(
        n10290) );
  AOI21_X1 U11030 ( .B1(n10287), .B2(n10286), .A(n10285), .ZN(n10288) );
  OR2_X1 U11031 ( .A1(n10299), .A2(n10288), .ZN(n10289) );
  NAND4_X1 U11032 ( .A1(n10292), .A2(n10291), .A3(n10290), .A4(n10289), .ZN(
        P1_U3250) );
  AOI22_X1 U11033 ( .A1(n10294), .A2(P1_ADDR_REG_10__SCAN_IN), .B1(n10339), 
        .B2(n10293), .ZN(n10306) );
  AOI21_X1 U11034 ( .B1(n10297), .B2(n10296), .A(n10295), .ZN(n10298) );
  OR2_X1 U11035 ( .A1(n10299), .A2(n10298), .ZN(n10304) );
  OAI211_X1 U11036 ( .C1(n10302), .C2(n10301), .A(n10335), .B(n10300), .ZN(
        n10303) );
  NAND4_X1 U11037 ( .A1(n10306), .A2(n10305), .A3(n10304), .A4(n10303), .ZN(
        P1_U3251) );
  NOR2_X1 U11038 ( .A1(n10308), .A2(n10307), .ZN(n10311) );
  AOI22_X1 U11039 ( .A1(n10312), .A2(n10311), .B1(n10310), .B2(n10309), .ZN(
        P2_U3437) );
  AOI22_X1 U11040 ( .A1(n10314), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(n4846), .ZN(n10332) );
  NAND2_X1 U11041 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n10315) );
  NAND2_X1 U11042 ( .A1(n10316), .A2(n10315), .ZN(n10317) );
  NAND2_X1 U11043 ( .A1(n10318), .A2(n10317), .ZN(n10328) );
  NAND2_X1 U11044 ( .A1(n10320), .A2(n10319), .ZN(n10327) );
  AND2_X1 U11045 ( .A1(n10322), .A2(n10321), .ZN(n10323) );
  OR3_X1 U11046 ( .A1(n10325), .A2(n10324), .A3(n10323), .ZN(n10326) );
  OAI211_X1 U11047 ( .C1(n10329), .C2(n10328), .A(n10327), .B(n10326), .ZN(
        n10330) );
  INV_X1 U11048 ( .A(n10330), .ZN(n10331) );
  NAND2_X1 U11049 ( .A1(n10332), .A2(n10331), .ZN(P2_U3246) );
  XNOR2_X1 U11050 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  INV_X1 U11051 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n10343) );
  NOR2_X1 U11052 ( .A1(n10334), .A2(n10333), .ZN(n10336) );
  OAI21_X1 U11053 ( .B1(n10337), .B2(n10336), .A(n10335), .ZN(n10341) );
  NAND2_X1 U11054 ( .A1(n10339), .A2(n10338), .ZN(n10340) );
  OAI211_X1 U11055 ( .C1(n10343), .C2(n10342), .A(n10341), .B(n10340), .ZN(
        n10344) );
  INV_X1 U11056 ( .A(n10344), .ZN(n10353) );
  OAI21_X1 U11057 ( .B1(n10347), .B2(n10346), .A(n10345), .ZN(n10348) );
  NAND2_X1 U11058 ( .A1(n10349), .A2(n10348), .ZN(n10350) );
  NAND4_X1 U11059 ( .A1(n10353), .A2(n10352), .A3(n10351), .A4(n10350), .ZN(
        P1_U3245) );
  INV_X1 U11060 ( .A(n10370), .ZN(n10585) );
  INV_X1 U11061 ( .A(n10354), .ZN(n10356) );
  OAI211_X1 U11062 ( .C1(n10357), .C2(n10581), .A(n10356), .B(n10355), .ZN(
        n10360) );
  INV_X1 U11063 ( .A(n10358), .ZN(n10359) );
  AOI211_X1 U11064 ( .C1(n10585), .C2(n10361), .A(n10360), .B(n10359), .ZN(
        n10363) );
  AOI22_X1 U11065 ( .A1(n10590), .A2(n10363), .B1(n7267), .B2(n10589), .ZN(
        P1_U3524) );
  INV_X1 U11066 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n10362) );
  AOI22_X1 U11067 ( .A1(n10594), .A2(n10363), .B1(n10362), .B2(n10591), .ZN(
        P1_U3457) );
  AOI22_X1 U11068 ( .A1(n10367), .A2(n10366), .B1(n10365), .B2(n10364), .ZN(
        n10368) );
  OAI211_X1 U11069 ( .C1(n10371), .C2(n10370), .A(n10369), .B(n10368), .ZN(
        n10372) );
  INV_X1 U11070 ( .A(n10372), .ZN(n10375) );
  AOI22_X1 U11071 ( .A1(n10590), .A2(n10375), .B1(n10373), .B2(n10589), .ZN(
        P1_U3525) );
  INV_X1 U11072 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n10374) );
  AOI22_X1 U11073 ( .A1(n10594), .A2(n10375), .B1(n10374), .B2(n10591), .ZN(
        P1_U3460) );
  INV_X1 U11074 ( .A(n10376), .ZN(n10381) );
  OAI22_X1 U11075 ( .A1(n10378), .A2(n10673), .B1(n10377), .B2(n10672), .ZN(
        n10380) );
  AOI211_X1 U11076 ( .C1(n10622), .C2(n10381), .A(n10380), .B(n10379), .ZN(
        n10382) );
  AOI22_X1 U11077 ( .A1(n10681), .A2(n10382), .B1(n7168), .B2(n10679), .ZN(
        P2_U3522) );
  AOI22_X1 U11078 ( .A1(n10684), .A2(n10382), .B1(n6224), .B2(n10682), .ZN(
        P2_U3457) );
  INV_X1 U11079 ( .A(n10383), .ZN(n10387) );
  OAI22_X1 U11080 ( .A1(n10384), .A2(n10582), .B1(n7633), .B2(n10581), .ZN(
        n10386) );
  AOI211_X1 U11081 ( .C1(n10585), .C2(n10387), .A(n10386), .B(n10385), .ZN(
        n10390) );
  AOI22_X1 U11082 ( .A1(n10590), .A2(n10390), .B1(n10388), .B2(n10589), .ZN(
        P1_U3526) );
  INV_X1 U11083 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n10389) );
  AOI22_X1 U11084 ( .A1(n10594), .A2(n10390), .B1(n10389), .B2(n10591), .ZN(
        P1_U3463) );
  INV_X1 U11085 ( .A(n10391), .ZN(n10396) );
  OAI22_X1 U11086 ( .A1(n10393), .A2(n10673), .B1(n10392), .B2(n10672), .ZN(
        n10395) );
  AOI211_X1 U11087 ( .C1(n10622), .C2(n10396), .A(n10395), .B(n10394), .ZN(
        n10398) );
  AOI22_X1 U11088 ( .A1(n10681), .A2(n10398), .B1(n10397), .B2(n10679), .ZN(
        P2_U3523) );
  AOI22_X1 U11089 ( .A1(n10684), .A2(n10398), .B1(n6267), .B2(n10682), .ZN(
        P2_U3460) );
  XNOR2_X1 U11090 ( .A(n10406), .B(n10399), .ZN(n10420) );
  INV_X1 U11091 ( .A(n10400), .ZN(n10402) );
  OAI21_X1 U11092 ( .B1(n10402), .B2(n10423), .A(n10401), .ZN(n10418) );
  OAI22_X1 U11093 ( .A1(n10418), .A2(n10582), .B1(n10423), .B2(n10581), .ZN(
        n10414) );
  OAI22_X1 U11094 ( .A1(n10491), .A2(n10489), .B1(n10403), .B2(n7059), .ZN(
        n10412) );
  NAND2_X1 U11095 ( .A1(n10408), .A2(n10407), .ZN(n10405) );
  INV_X1 U11096 ( .A(n10406), .ZN(n10404) );
  NAND2_X1 U11097 ( .A1(n10405), .A2(n10404), .ZN(n10410) );
  NAND3_X1 U11098 ( .A1(n10408), .A2(n10407), .A3(n10406), .ZN(n10409) );
  AOI21_X1 U11099 ( .B1(n10410), .B2(n10409), .A(n7060), .ZN(n10411) );
  AOI211_X1 U11100 ( .C1(n10522), .C2(n10420), .A(n10412), .B(n10411), .ZN(
        n10413) );
  INV_X1 U11101 ( .A(n10413), .ZN(n10425) );
  AOI211_X1 U11102 ( .C1(n10585), .C2(n10420), .A(n10414), .B(n10425), .ZN(
        n10417) );
  AOI22_X1 U11103 ( .A1(n10590), .A2(n10417), .B1(n10415), .B2(n10589), .ZN(
        P1_U3527) );
  INV_X1 U11104 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10416) );
  AOI22_X1 U11105 ( .A1(n10594), .A2(n10417), .B1(n10416), .B2(n10591), .ZN(
        P1_U3466) );
  INV_X1 U11106 ( .A(n10418), .ZN(n10419) );
  AOI22_X1 U11107 ( .A1(n10420), .A2(n10559), .B1(n10558), .B2(n10419), .ZN(
        n10427) );
  AOI22_X1 U11108 ( .A1(n10563), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n10421), 
        .B2(n10561), .ZN(n10422) );
  OAI21_X1 U11109 ( .B1(n10423), .B2(n10565), .A(n10422), .ZN(n10424) );
  AOI21_X1 U11110 ( .B1(n10425), .B2(n10568), .A(n10424), .ZN(n10426) );
  NAND2_X1 U11111 ( .A1(n10427), .A2(n10426), .ZN(P1_U3287) );
  INV_X1 U11112 ( .A(n10428), .ZN(n10429) );
  AOI21_X1 U11113 ( .B1(n6285), .B2(n10430), .A(n10429), .ZN(n10457) );
  INV_X1 U11114 ( .A(n10431), .ZN(n10433) );
  OAI21_X1 U11115 ( .B1(n10433), .B2(n10434), .A(n10432), .ZN(n10453) );
  OAI22_X1 U11116 ( .A1(n10453), .A2(n10673), .B1(n10434), .B2(n10672), .ZN(
        n10444) );
  AOI21_X1 U11117 ( .B1(n10435), .B2(n10437), .A(n10436), .ZN(n10442) );
  OAI22_X1 U11118 ( .A1(n10439), .A2(n10613), .B1(n10438), .B2(n10611), .ZN(
        n10440) );
  AOI21_X1 U11119 ( .B1(n10442), .B2(n10441), .A(n10440), .ZN(n10459) );
  INV_X1 U11120 ( .A(n10459), .ZN(n10443) );
  AOI211_X1 U11121 ( .C1(n10457), .C2(n10677), .A(n10444), .B(n10443), .ZN(
        n10445) );
  AOI22_X1 U11122 ( .A1(n10681), .A2(n10445), .B1(n7170), .B2(n10679), .ZN(
        P2_U3524) );
  AOI22_X1 U11123 ( .A1(n10684), .A2(n10445), .B1(n6274), .B2(n10682), .ZN(
        P2_U3463) );
  OAI22_X1 U11124 ( .A1(n10448), .A2(n7155), .B1(n10447), .B2(n10446), .ZN(
        n10449) );
  AOI21_X1 U11125 ( .B1(n10451), .B2(n10450), .A(n10449), .ZN(n10452) );
  OAI21_X1 U11126 ( .B1(n10454), .B2(n10453), .A(n10452), .ZN(n10455) );
  AOI21_X1 U11127 ( .B1(n10457), .B2(n10456), .A(n10455), .ZN(n10458) );
  OAI21_X1 U11128 ( .B1(n9157), .B2(n10459), .A(n10458), .ZN(P2_U3292) );
  INV_X1 U11129 ( .A(n10460), .ZN(n10467) );
  INV_X1 U11130 ( .A(n10461), .ZN(n10462) );
  OAI21_X1 U11131 ( .B1(n10463), .B2(n10581), .A(n10462), .ZN(n10466) );
  INV_X1 U11132 ( .A(n10464), .ZN(n10465) );
  AOI211_X1 U11133 ( .C1(n10468), .C2(n10467), .A(n10466), .B(n10465), .ZN(
        n10471) );
  AOI22_X1 U11134 ( .A1(n10590), .A2(n10471), .B1(n10469), .B2(n10589), .ZN(
        P1_U3528) );
  INV_X1 U11135 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n10470) );
  AOI22_X1 U11136 ( .A1(n10594), .A2(n10471), .B1(n10470), .B2(n10591), .ZN(
        P1_U3469) );
  AOI21_X1 U11137 ( .B1(n10662), .B2(n10473), .A(n10472), .ZN(n10474) );
  OAI211_X1 U11138 ( .C1(n10667), .C2(n10476), .A(n10475), .B(n10474), .ZN(
        n10477) );
  INV_X1 U11139 ( .A(n10477), .ZN(n10478) );
  AOI22_X1 U11140 ( .A1(n10681), .A2(n10478), .B1(n7171), .B2(n10679), .ZN(
        P2_U3525) );
  AOI22_X1 U11141 ( .A1(n10684), .A2(n10478), .B1(n6291), .B2(n10682), .ZN(
        P2_U3466) );
  OAI21_X1 U11142 ( .B1(n7098), .B2(n7097), .A(n10479), .ZN(n10501) );
  INV_X1 U11143 ( .A(n10480), .ZN(n10481) );
  OAI21_X1 U11144 ( .B1(n10502), .B2(n10482), .A(n10481), .ZN(n10499) );
  OAI22_X1 U11145 ( .A1(n10499), .A2(n10582), .B1(n10502), .B2(n10581), .ZN(
        n10495) );
  INV_X1 U11146 ( .A(n10483), .ZN(n10484) );
  AOI21_X1 U11147 ( .B1(n10486), .B2(n10485), .A(n10484), .ZN(n10488) );
  XNOR2_X1 U11148 ( .A(n10488), .B(n10487), .ZN(n10494) );
  OAI22_X1 U11149 ( .A1(n10491), .A2(n7059), .B1(n10490), .B2(n10489), .ZN(
        n10492) );
  AOI21_X1 U11150 ( .B1(n10501), .B2(n10522), .A(n10492), .ZN(n10493) );
  OAI21_X1 U11151 ( .B1(n10494), .B2(n7060), .A(n10493), .ZN(n10503) );
  AOI211_X1 U11152 ( .C1(n10585), .C2(n10501), .A(n10495), .B(n10503), .ZN(
        n10498) );
  AOI22_X1 U11153 ( .A1(n10590), .A2(n10498), .B1(n10496), .B2(n10589), .ZN(
        P1_U3529) );
  INV_X1 U11154 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10497) );
  AOI22_X1 U11155 ( .A1(n10594), .A2(n10498), .B1(n10497), .B2(n10591), .ZN(
        P1_U3472) );
  INV_X1 U11156 ( .A(n10499), .ZN(n10500) );
  AOI22_X1 U11157 ( .A1(n10501), .A2(n10559), .B1(n10558), .B2(n10500), .ZN(
        n10508) );
  NOR2_X1 U11158 ( .A1(n10565), .A2(n10502), .ZN(n10505) );
  MUX2_X1 U11159 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n10503), .S(n10568), .Z(
        n10504) );
  AOI211_X1 U11160 ( .C1(n10561), .C2(n10506), .A(n10505), .B(n10504), .ZN(
        n10507) );
  NAND2_X1 U11161 ( .A1(n10508), .A2(n10507), .ZN(P1_U3285) );
  OAI22_X1 U11162 ( .A1(n10510), .A2(n10673), .B1(n10509), .B2(n10672), .ZN(
        n10512) );
  AOI211_X1 U11163 ( .C1(n10677), .C2(n10513), .A(n10512), .B(n10511), .ZN(
        n10515) );
  AOI22_X1 U11164 ( .A1(n10681), .A2(n10515), .B1(n7192), .B2(n10679), .ZN(
        P2_U3526) );
  INV_X1 U11165 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10514) );
  AOI22_X1 U11166 ( .A1(n10684), .A2(n10515), .B1(n10514), .B2(n10682), .ZN(
        P2_U3469) );
  NAND2_X1 U11167 ( .A1(n10521), .A2(n10585), .ZN(n10517) );
  OAI211_X1 U11168 ( .C1(n10518), .C2(n10581), .A(n10517), .B(n10516), .ZN(
        n10520) );
  AOI211_X1 U11169 ( .C1(n10522), .C2(n10521), .A(n10520), .B(n10519), .ZN(
        n10524) );
  AOI22_X1 U11170 ( .A1(n10590), .A2(n10524), .B1(n7331), .B2(n10589), .ZN(
        P1_U3530) );
  INV_X1 U11171 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n10523) );
  AOI22_X1 U11172 ( .A1(n10594), .A2(n10524), .B1(n10523), .B2(n10591), .ZN(
        P1_U3475) );
  AOI22_X1 U11173 ( .A1(n10526), .A2(n10663), .B1(n10662), .B2(n10525), .ZN(
        n10527) );
  OAI211_X1 U11174 ( .C1(n10667), .C2(n10529), .A(n10528), .B(n10527), .ZN(
        n10530) );
  INV_X1 U11175 ( .A(n10530), .ZN(n10531) );
  AOI22_X1 U11176 ( .A1(n10681), .A2(n10531), .B1(n7206), .B2(n10679), .ZN(
        P2_U3527) );
  AOI22_X1 U11177 ( .A1(n10684), .A2(n10531), .B1(n6318), .B2(n10682), .ZN(
        P2_U3472) );
  NAND2_X1 U11178 ( .A1(n10533), .A2(n10544), .ZN(n10534) );
  NAND2_X1 U11179 ( .A1(n10532), .A2(n10534), .ZN(n10551) );
  INV_X1 U11180 ( .A(n10551), .ZN(n10560) );
  INV_X1 U11181 ( .A(n10535), .ZN(n10537) );
  OAI21_X1 U11182 ( .B1(n10537), .B2(n10566), .A(n10536), .ZN(n10556) );
  OAI22_X1 U11183 ( .A1(n10556), .A2(n10582), .B1(n10566), .B2(n10581), .ZN(
        n10552) );
  AOI22_X1 U11184 ( .A1(n10541), .A2(n10540), .B1(n10539), .B2(n10538), .ZN(
        n10549) );
  NAND2_X1 U11185 ( .A1(n10543), .A2(n10542), .ZN(n10545) );
  XNOR2_X1 U11186 ( .A(n10545), .B(n10544), .ZN(n10547) );
  NAND2_X1 U11187 ( .A1(n10547), .A2(n10546), .ZN(n10548) );
  OAI211_X1 U11188 ( .C1(n10551), .C2(n10550), .A(n10549), .B(n10548), .ZN(
        n10569) );
  AOI211_X1 U11189 ( .C1(n10585), .C2(n10560), .A(n10552), .B(n10569), .ZN(
        n10555) );
  AOI22_X1 U11190 ( .A1(n10590), .A2(n10555), .B1(n10553), .B2(n10589), .ZN(
        P1_U3531) );
  INV_X1 U11191 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n10554) );
  AOI22_X1 U11192 ( .A1(n10594), .A2(n10555), .B1(n10554), .B2(n10591), .ZN(
        P1_U3478) );
  INV_X1 U11193 ( .A(n10556), .ZN(n10557) );
  AOI22_X1 U11194 ( .A1(n10560), .A2(n10559), .B1(n10558), .B2(n10557), .ZN(
        n10571) );
  AOI22_X1 U11195 ( .A1(n10563), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n10562), 
        .B2(n10561), .ZN(n10564) );
  OAI21_X1 U11196 ( .B1(n10566), .B2(n10565), .A(n10564), .ZN(n10567) );
  AOI21_X1 U11197 ( .B1(n10569), .B2(n10568), .A(n10567), .ZN(n10570) );
  NAND2_X1 U11198 ( .A1(n10571), .A2(n10570), .ZN(P1_U3283) );
  NAND3_X1 U11199 ( .A1(n8133), .A2(n10572), .A3(n10677), .ZN(n10574) );
  OAI211_X1 U11200 ( .C1(n10575), .C2(n10672), .A(n10574), .B(n10573), .ZN(
        n10576) );
  NOR2_X1 U11201 ( .A1(n10577), .A2(n10576), .ZN(n10579) );
  INV_X1 U11202 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n10578) );
  AOI22_X1 U11203 ( .A1(n10681), .A2(n10579), .B1(n10578), .B2(n10679), .ZN(
        P2_U3528) );
  AOI22_X1 U11204 ( .A1(n10684), .A2(n10579), .B1(n6333), .B2(n10682), .ZN(
        P2_U3475) );
  OAI22_X1 U11205 ( .A1(n10583), .A2(n10582), .B1(n5000), .B2(n10581), .ZN(
        n10584) );
  AOI21_X1 U11206 ( .B1(n10586), .B2(n10585), .A(n10584), .ZN(n10587) );
  AOI22_X1 U11207 ( .A1(n10590), .A2(n10593), .B1(n7573), .B2(n10589), .ZN(
        P1_U3532) );
  INV_X1 U11208 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n10592) );
  AOI22_X1 U11209 ( .A1(n10594), .A2(n10593), .B1(n10592), .B2(n10591), .ZN(
        P1_U3481) );
  OAI22_X1 U11210 ( .A1(n10596), .A2(n10673), .B1(n10595), .B2(n10672), .ZN(
        n10598) );
  AOI211_X1 U11211 ( .C1(n10622), .C2(n10599), .A(n10598), .B(n10597), .ZN(
        n10600) );
  AOI22_X1 U11212 ( .A1(n10681), .A2(n10600), .B1(n7527), .B2(n10679), .ZN(
        P2_U3529) );
  AOI22_X1 U11213 ( .A1(n10684), .A2(n10600), .B1(n6349), .B2(n10682), .ZN(
        P2_U3478) );
  OR2_X1 U11214 ( .A1(n10602), .A2(n10601), .ZN(n10603) );
  NAND2_X1 U11215 ( .A1(n10604), .A2(n10603), .ZN(n10620) );
  INV_X1 U11216 ( .A(n10620), .ZN(n10628) );
  INV_X1 U11217 ( .A(n10605), .ZN(n10608) );
  INV_X1 U11218 ( .A(n10606), .ZN(n10633) );
  OAI21_X1 U11219 ( .B1(n10608), .B2(n10633), .A(n10607), .ZN(n10624) );
  OAI22_X1 U11220 ( .A1(n10624), .A2(n10673), .B1(n10633), .B2(n10672), .ZN(
        n10621) );
  OAI21_X1 U11221 ( .B1(n4914), .B2(n10610), .A(n10609), .ZN(n10617) );
  OAI22_X1 U11222 ( .A1(n10614), .A2(n10613), .B1(n10612), .B2(n10611), .ZN(
        n10615) );
  AOI21_X1 U11223 ( .B1(n10617), .B2(n10616), .A(n10615), .ZN(n10618) );
  OAI21_X1 U11224 ( .B1(n10620), .B2(n10619), .A(n10618), .ZN(n10636) );
  AOI211_X1 U11225 ( .C1(n10622), .C2(n10628), .A(n10621), .B(n10636), .ZN(
        n10623) );
  AOI22_X1 U11226 ( .A1(n10681), .A2(n10623), .B1(n7620), .B2(n10679), .ZN(
        P2_U3530) );
  AOI22_X1 U11227 ( .A1(n10684), .A2(n10623), .B1(n6359), .B2(n10682), .ZN(
        P2_U3481) );
  INV_X1 U11228 ( .A(n10624), .ZN(n10625) );
  AOI22_X1 U11229 ( .A1(n10628), .A2(n10627), .B1(n10626), .B2(n10625), .ZN(
        n10638) );
  AOI22_X1 U11230 ( .A1(n10631), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n10630), 
        .B2(n10629), .ZN(n10632) );
  OAI21_X1 U11231 ( .B1(n10634), .B2(n10633), .A(n10632), .ZN(n10635) );
  AOI21_X1 U11232 ( .B1(n10636), .B2(n10448), .A(n10635), .ZN(n10637) );
  NAND2_X1 U11233 ( .A1(n10638), .A2(n10637), .ZN(P2_U3286) );
  AOI21_X1 U11234 ( .B1(n10662), .B2(n10640), .A(n10639), .ZN(n10641) );
  OAI211_X1 U11235 ( .C1(n10643), .C2(n10667), .A(n10642), .B(n10641), .ZN(
        n10644) );
  INV_X1 U11236 ( .A(n10644), .ZN(n10646) );
  AOI22_X1 U11237 ( .A1(n10681), .A2(n10646), .B1(n10645), .B2(n10679), .ZN(
        P2_U3531) );
  AOI22_X1 U11238 ( .A1(n10684), .A2(n10646), .B1(n6379), .B2(n10682), .ZN(
        P2_U3484) );
  OAI22_X1 U11239 ( .A1(n10648), .A2(n10673), .B1(n10647), .B2(n10672), .ZN(
        n10650) );
  AOI211_X1 U11240 ( .C1(n10677), .C2(n10651), .A(n10650), .B(n10649), .ZN(
        n10652) );
  AOI22_X1 U11241 ( .A1(n10681), .A2(n10652), .B1(n7934), .B2(n10679), .ZN(
        P2_U3532) );
  AOI22_X1 U11242 ( .A1(n10684), .A2(n10652), .B1(n6396), .B2(n10682), .ZN(
        P2_U3487) );
  NOR2_X1 U11243 ( .A1(n10653), .A2(n10667), .ZN(n10658) );
  OAI22_X1 U11244 ( .A1(n10655), .A2(n10673), .B1(n10654), .B2(n10672), .ZN(
        n10657) );
  AOI211_X1 U11245 ( .C1(n10658), .C2(n8492), .A(n10657), .B(n10656), .ZN(
        n10660) );
  AOI22_X1 U11246 ( .A1(n10681), .A2(n10660), .B1(n10659), .B2(n10679), .ZN(
        P2_U3533) );
  AOI22_X1 U11247 ( .A1(n10684), .A2(n10660), .B1(n6409), .B2(n10682), .ZN(
        P2_U3490) );
  AOI22_X1 U11248 ( .A1(n10664), .A2(n10663), .B1(n10662), .B2(n10661), .ZN(
        n10665) );
  OAI211_X1 U11249 ( .C1(n10668), .C2(n10667), .A(n10666), .B(n10665), .ZN(
        n10669) );
  INV_X1 U11250 ( .A(n10669), .ZN(n10671) );
  AOI22_X1 U11251 ( .A1(n10681), .A2(n10671), .B1(n10670), .B2(n10679), .ZN(
        P2_U3534) );
  AOI22_X1 U11252 ( .A1(n10684), .A2(n10671), .B1(n6425), .B2(n10682), .ZN(
        P2_U3493) );
  OAI22_X1 U11253 ( .A1(n10674), .A2(n10673), .B1(n5164), .B2(n10672), .ZN(
        n10676) );
  AOI211_X1 U11254 ( .C1(n10678), .C2(n10677), .A(n10676), .B(n10675), .ZN(
        n10683) );
  INV_X1 U11255 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n10680) );
  AOI22_X1 U11256 ( .A1(n10681), .A2(n10683), .B1(n10680), .B2(n10679), .ZN(
        P2_U3535) );
  AOI22_X1 U11257 ( .A1(n10684), .A2(n10683), .B1(n6441), .B2(n10682), .ZN(
        P2_U3496) );
  XNOR2_X1 U11258 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  BUF_X1 U4962 ( .A(n5734), .Z(n6031) );
  BUF_X1 U4961 ( .A(n5760), .Z(n5956) );
  CLKBUF_X1 U4919 ( .A(n6259), .Z(n4851) );
  CLKBUF_X3 U4920 ( .A(n5763), .Z(n6032) );
  CLKBUF_X1 U4922 ( .A(n6624), .Z(n4849) );
endmodule

