

module b22_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, keyinput_128, keyinput_129, 
        keyinput_130, keyinput_131, keyinput_132, keyinput_133, keyinput_134, 
        keyinput_135, keyinput_136, keyinput_137, keyinput_138, keyinput_139, 
        keyinput_140, keyinput_141, keyinput_142, keyinput_143, keyinput_144, 
        keyinput_145, keyinput_146, keyinput_147, keyinput_148, keyinput_149, 
        keyinput_150, keyinput_151, keyinput_152, keyinput_153, keyinput_154, 
        keyinput_155, keyinput_156, keyinput_157, keyinput_158, keyinput_159, 
        keyinput_160, keyinput_161, keyinput_162, keyinput_163, keyinput_164, 
        keyinput_165, keyinput_166, keyinput_167, keyinput_168, keyinput_169, 
        keyinput_170, keyinput_171, keyinput_172, keyinput_173, keyinput_174, 
        keyinput_175, keyinput_176, keyinput_177, keyinput_178, keyinput_179, 
        keyinput_180, keyinput_181, keyinput_182, keyinput_183, keyinput_184, 
        keyinput_185, keyinput_186, keyinput_187, keyinput_188, keyinput_189, 
        keyinput_190, keyinput_191, keyinput_192, keyinput_193, keyinput_194, 
        keyinput_195, keyinput_196, keyinput_197, keyinput_198, keyinput_199, 
        keyinput_200, keyinput_201, keyinput_202, keyinput_203, keyinput_204, 
        keyinput_205, keyinput_206, keyinput_207, keyinput_208, keyinput_209, 
        keyinput_210, keyinput_211, keyinput_212, keyinput_213, keyinput_214, 
        keyinput_215, keyinput_216, keyinput_217, keyinput_218, keyinput_219, 
        keyinput_220, keyinput_221, keyinput_222, keyinput_223, keyinput_224, 
        keyinput_225, keyinput_226, keyinput_227, keyinput_228, keyinput_229, 
        keyinput_230, keyinput_231, keyinput_232, keyinput_233, keyinput_234, 
        keyinput_235, keyinput_236, keyinput_237, keyinput_238, keyinput_239, 
        keyinput_240, keyinput_241, keyinput_242, keyinput_243, keyinput_244, 
        keyinput_245, keyinput_246, keyinput_247, keyinput_248, keyinput_249, 
        keyinput_250, keyinput_251, keyinput_252, keyinput_253, keyinput_254, 
        keyinput_255, P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, 
        SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, 
        SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, 
        SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_, 
        P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, SUB_1596_U4, 
        SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, 
        SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, 
        SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, 
        SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, U29, U28, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, 
        P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, 
        P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, P1_U3515, 
        P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, 
        P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, 
        P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, 
        P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, 
        P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, 
        P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, P1_U3557, 
        P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, P1_U3561, 
        P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, 
        P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, 
        P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, 
        P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, P1_U3589, 
        P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U4016, 
        P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, 
        P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, 
        P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, 
        P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, 
        P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, P2_U3295, 
        P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, 
        P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, 
        P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, 
        P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, 
        P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, P2_U3445, 
        P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, 
        P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3486, 
        P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, P2_U3493, 
        P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, 
        P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, 
        P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, 
        P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, 
        P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, 
        P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, 
        P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, P2_U3532, 
        P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, 
        P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, 
        P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, P2_U3553, 
        P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, 
        P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, P2_U3210, 
        P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, 
        P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, 
        P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, 
        P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, P2_U3947, 
        P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, P3_U3289, 
        P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, P3_U3282, 
        P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, P3_U3275, 
        P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, P3_U3268, 
        P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, P3_U3263, 
        P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, P3_U3256, 
        P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, P3_U3249, 
        P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, P3_U3242, 
        P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, P3_U3235, 
        P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, P3_U3405, 
        P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, P3_U3426, 
        P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, P3_U3446, 
        P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, P3_U3453, 
        P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, P3_U3460, 
        P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, P3_U3467, 
        P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, P3_U3474, 
        P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, P3_U3481, 
        P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, P3_U3488, 
        P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, P3_U3229, 
        P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, P3_U3222, 
        P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, P3_U3215, 
        P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, P3_U3208, 
        P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, P3_U3201, 
        P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, P3_U3194, 
        P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, P3_U3187, 
        P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, P3_U3492, 
        P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, P3_U3499, 
        P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, P3_U3506, 
        P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, P3_U3513, 
        P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, P3_U3520, 
        P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, P3_U3178, 
        P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, P3_U3171, 
        P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, P3_U3164, 
        P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, P3_U3157, 
        P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, P3_U3897
 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, keyinput_128, keyinput_129, keyinput_130,
         keyinput_131, keyinput_132, keyinput_133, keyinput_134, keyinput_135,
         keyinput_136, keyinput_137, keyinput_138, keyinput_139, keyinput_140,
         keyinput_141, keyinput_142, keyinput_143, keyinput_144, keyinput_145,
         keyinput_146, keyinput_147, keyinput_148, keyinput_149, keyinput_150,
         keyinput_151, keyinput_152, keyinput_153, keyinput_154, keyinput_155,
         keyinput_156, keyinput_157, keyinput_158, keyinput_159, keyinput_160,
         keyinput_161, keyinput_162, keyinput_163, keyinput_164, keyinput_165,
         keyinput_166, keyinput_167, keyinput_168, keyinput_169, keyinput_170,
         keyinput_171, keyinput_172, keyinput_173, keyinput_174, keyinput_175,
         keyinput_176, keyinput_177, keyinput_178, keyinput_179, keyinput_180,
         keyinput_181, keyinput_182, keyinput_183, keyinput_184, keyinput_185,
         keyinput_186, keyinput_187, keyinput_188, keyinput_189, keyinput_190,
         keyinput_191, keyinput_192, keyinput_193, keyinput_194, keyinput_195,
         keyinput_196, keyinput_197, keyinput_198, keyinput_199, keyinput_200,
         keyinput_201, keyinput_202, keyinput_203, keyinput_204, keyinput_205,
         keyinput_206, keyinput_207, keyinput_208, keyinput_209, keyinput_210,
         keyinput_211, keyinput_212, keyinput_213, keyinput_214, keyinput_215,
         keyinput_216, keyinput_217, keyinput_218, keyinput_219, keyinput_220,
         keyinput_221, keyinput_222, keyinput_223, keyinput_224, keyinput_225,
         keyinput_226, keyinput_227, keyinput_228, keyinput_229, keyinput_230,
         keyinput_231, keyinput_232, keyinput_233, keyinput_234, keyinput_235,
         keyinput_236, keyinput_237, keyinput_238, keyinput_239, keyinput_240,
         keyinput_241, keyinput_242, keyinput_243, keyinput_244, keyinput_245,
         keyinput_246, keyinput_247, keyinput_248, keyinput_249, keyinput_250,
         keyinput_251, keyinput_252, keyinput_253, keyinput_254, keyinput_255,
         P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n7410, n7411, n7412, n7413, n7414, n7416, n7417, n7418, n7419, n7420,
         n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430,
         n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440,
         n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450,
         n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460,
         n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470,
         n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480,
         n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490,
         n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500,
         n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510,
         n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520,
         n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530,
         n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540,
         n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550,
         n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560,
         n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570,
         n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580,
         n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590,
         n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600,
         n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610,
         n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620,
         n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630,
         n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640,
         n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650,
         n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660,
         n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670,
         n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680,
         n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690,
         n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700,
         n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710,
         n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720,
         n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730,
         n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740,
         n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750,
         n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760,
         n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770,
         n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780,
         n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790,
         n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800,
         n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810,
         n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820,
         n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830,
         n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840,
         n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850,
         n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860,
         n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870,
         n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880,
         n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890,
         n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900,
         n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910,
         n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920,
         n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930,
         n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940,
         n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950,
         n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960,
         n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970,
         n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980,
         n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990,
         n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000,
         n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010,
         n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020,
         n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030,
         n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040,
         n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050,
         n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060,
         n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070,
         n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080,
         n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090,
         n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100,
         n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110,
         n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120,
         n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130,
         n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140,
         n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150,
         n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160,
         n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170,
         n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180,
         n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190,
         n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200,
         n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210,
         n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220,
         n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230,
         n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240,
         n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250,
         n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260,
         n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270,
         n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280,
         n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290,
         n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300,
         n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310,
         n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320,
         n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330,
         n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340,
         n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350,
         n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360,
         n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370,
         n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380,
         n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390,
         n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400,
         n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410,
         n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420,
         n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430,
         n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440,
         n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450,
         n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460,
         n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470,
         n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480,
         n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490,
         n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500,
         n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510,
         n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520,
         n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530,
         n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540,
         n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550,
         n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560,
         n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570,
         n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580,
         n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590,
         n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600,
         n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610,
         n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620,
         n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630,
         n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640,
         n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650,
         n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660,
         n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670,
         n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680,
         n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690,
         n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700,
         n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710,
         n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720,
         n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730,
         n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740,
         n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750,
         n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760,
         n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770,
         n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780,
         n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790,
         n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800,
         n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810,
         n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820,
         n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830,
         n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840,
         n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850,
         n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860,
         n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870,
         n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880,
         n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890,
         n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900,
         n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910,
         n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920,
         n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930,
         n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940,
         n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950,
         n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960,
         n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970,
         n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980,
         n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990,
         n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000,
         n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010,
         n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020,
         n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030,
         n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040,
         n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050,
         n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060,
         n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070,
         n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080,
         n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090,
         n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100,
         n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110,
         n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120,
         n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130,
         n9131, n9132, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141,
         n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151,
         n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161,
         n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171,
         n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181,
         n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191,
         n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201,
         n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211,
         n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221,
         n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231,
         n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241,
         n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251,
         n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261,
         n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271,
         n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281,
         n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291,
         n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301,
         n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311,
         n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321,
         n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331,
         n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341,
         n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351,
         n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361,
         n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371,
         n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381,
         n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391,
         n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401,
         n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411,
         n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421,
         n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431,
         n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441,
         n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451,
         n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461,
         n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471,
         n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481,
         n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491,
         n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501,
         n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511,
         n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521,
         n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531,
         n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541,
         n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551,
         n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561,
         n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571,
         n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581,
         n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591,
         n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601,
         n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611,
         n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621,
         n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631,
         n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641,
         n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651,
         n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661,
         n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671,
         n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681,
         n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691,
         n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701,
         n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711,
         n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721,
         n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731,
         n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741,
         n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751,
         n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761,
         n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771,
         n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781,
         n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791,
         n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801,
         n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811,
         n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821,
         n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831,
         n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841,
         n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851,
         n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861,
         n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871,
         n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881,
         n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891,
         n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901,
         n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911,
         n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921,
         n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931,
         n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941,
         n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951,
         n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961,
         n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971,
         n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981,
         n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991,
         n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
         n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
         n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
         n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
         n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
         n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,
         n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
         n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
         n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656,
         n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664,
         n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672,
         n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680,
         n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688,
         n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696,
         n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704,
         n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712,
         n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720,
         n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728,
         n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736,
         n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744,
         n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752,
         n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760,
         n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768,
         n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776,
         n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784,
         n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792,
         n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800,
         n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808,
         n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816,
         n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824,
         n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832,
         n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840,
         n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848,
         n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856,
         n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864,
         n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872,
         n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880,
         n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888,
         n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896,
         n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904,
         n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912,
         n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920,
         n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928,
         n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936,
         n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944,
         n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952,
         n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960,
         n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968,
         n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976,
         n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984,
         n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992,
         n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000,
         n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008,
         n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016,
         n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024,
         n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032,
         n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040,
         n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048,
         n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056,
         n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064,
         n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072,
         n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080,
         n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088,
         n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096,
         n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104,
         n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112,
         n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120,
         n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128,
         n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136,
         n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144,
         n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152,
         n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160,
         n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168,
         n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176,
         n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184,
         n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192,
         n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200,
         n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208,
         n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216,
         n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224,
         n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232,
         n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240,
         n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248,
         n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256,
         n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264,
         n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272,
         n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280,
         n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288,
         n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296,
         n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304,
         n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312,
         n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320,
         n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328,
         n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336,
         n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344,
         n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352,
         n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360,
         n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368,
         n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376,
         n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384,
         n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392,
         n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400,
         n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408,
         n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416,
         n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424,
         n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432,
         n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440,
         n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448,
         n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456,
         n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464,
         n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472,
         n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480,
         n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488,
         n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496,
         n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504,
         n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512,
         n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520,
         n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528,
         n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536,
         n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544,
         n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552,
         n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560,
         n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568,
         n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576,
         n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584,
         n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592,
         n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600,
         n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608,
         n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616,
         n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624,
         n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632,
         n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640,
         n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648,
         n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656,
         n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664,
         n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672,
         n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680,
         n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688,
         n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696,
         n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704,
         n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712,
         n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720,
         n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728,
         n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736,
         n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744,
         n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752,
         n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760,
         n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768,
         n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776,
         n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784,
         n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792,
         n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800,
         n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808,
         n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816,
         n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824,
         n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832,
         n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840,
         n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848,
         n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856,
         n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864,
         n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872,
         n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880,
         n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888,
         n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896,
         n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904,
         n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912,
         n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920,
         n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928,
         n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936,
         n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944,
         n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952,
         n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960,
         n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968,
         n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976,
         n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984,
         n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992,
         n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000,
         n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008,
         n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016,
         n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024,
         n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032,
         n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040,
         n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048,
         n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056,
         n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064,
         n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072,
         n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080,
         n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088,
         n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096,
         n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104,
         n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112,
         n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120,
         n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128,
         n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136,
         n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144,
         n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152,
         n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160,
         n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168,
         n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176,
         n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184,
         n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192,
         n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200,
         n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208,
         n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216,
         n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224,
         n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232,
         n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240,
         n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248,
         n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256,
         n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264,
         n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272,
         n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280,
         n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288,
         n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296,
         n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304,
         n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312,
         n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320,
         n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328,
         n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336,
         n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344,
         n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352,
         n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360,
         n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368,
         n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376,
         n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384,
         n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392,
         n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400,
         n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408,
         n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416,
         n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424,
         n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432,
         n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440,
         n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448,
         n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456,
         n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464,
         n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472,
         n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480,
         n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488,
         n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496,
         n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504,
         n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512,
         n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520,
         n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528,
         n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536,
         n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544,
         n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552,
         n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560,
         n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568,
         n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576,
         n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584,
         n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592,
         n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600,
         n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608,
         n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616,
         n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624,
         n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632,
         n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640,
         n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648,
         n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656,
         n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664,
         n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672,
         n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680,
         n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688,
         n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696,
         n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704,
         n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712,
         n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720,
         n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728,
         n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736,
         n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744,
         n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752,
         n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760,
         n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768,
         n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776,
         n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784,
         n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792,
         n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800,
         n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808,
         n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816,
         n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824,
         n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832,
         n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840,
         n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848,
         n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856,
         n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864,
         n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872,
         n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880,
         n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888,
         n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896,
         n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904,
         n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912,
         n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920,
         n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928,
         n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936,
         n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944,
         n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952,
         n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960,
         n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968,
         n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976,
         n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984,
         n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992,
         n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000,
         n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008,
         n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016,
         n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024,
         n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032,
         n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040,
         n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048,
         n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056,
         n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064,
         n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072,
         n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080,
         n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088,
         n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096,
         n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104,
         n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112,
         n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120,
         n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128,
         n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136,
         n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144,
         n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152,
         n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160,
         n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168,
         n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176,
         n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184,
         n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192,
         n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200,
         n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208,
         n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216,
         n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224,
         n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232,
         n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240,
         n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248,
         n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256,
         n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264,
         n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272,
         n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280,
         n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288,
         n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296,
         n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304,
         n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312,
         n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320,
         n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328,
         n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336,
         n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344,
         n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352,
         n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360,
         n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368,
         n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376,
         n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384,
         n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392,
         n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400,
         n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408,
         n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416,
         n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424,
         n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432,
         n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440,
         n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448,
         n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456,
         n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464,
         n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472,
         n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480,
         n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488,
         n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496,
         n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504,
         n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512,
         n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520,
         n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528,
         n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536,
         n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544,
         n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552,
         n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560,
         n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568,
         n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576,
         n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584,
         n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592,
         n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600,
         n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608,
         n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616,
         n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624,
         n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632,
         n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640,
         n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648,
         n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656,
         n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664,
         n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672,
         n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680,
         n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688,
         n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696,
         n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704,
         n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712,
         n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720,
         n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728,
         n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736,
         n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744,
         n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752,
         n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760,
         n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768,
         n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776,
         n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784,
         n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792,
         n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800,
         n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808,
         n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816,
         n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824,
         n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832,
         n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840,
         n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848,
         n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856,
         n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864,
         n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872,
         n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880,
         n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888,
         n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896,
         n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904,
         n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912,
         n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920,
         n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928,
         n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936,
         n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944,
         n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952,
         n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960,
         n13961, n13962, n13963, n13964, n13965, n13966, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
         n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
         n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
         n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
         n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
         n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
         n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
         n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897,
         n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
         n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913,
         n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
         n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929,
         n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937,
         n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
         n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
         n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
         n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
         n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
         n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
         n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009,
         n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
         n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
         n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
         n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041,
         n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
         n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
         n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
         n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073,
         n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081,
         n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089,
         n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097,
         n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105,
         n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113,
         n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121,
         n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
         n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
         n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145,
         n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153,
         n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161,
         n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169,
         n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177,
         n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185,
         n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
         n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
         n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
         n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217,
         n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225,
         n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
         n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241,
         n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249,
         n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257,
         n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265,
         n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273,
         n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281,
         n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289,
         n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297,
         n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305,
         n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313,
         n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321,
         n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329,
         n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
         n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345,
         n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353,
         n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361,
         n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369,
         n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377,
         n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385,
         n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393,
         n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401,
         n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409,
         n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417,
         n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425,
         n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433,
         n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441,
         n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449,
         n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457,
         n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465,
         n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473,
         n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481,
         n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489,
         n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497,
         n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505,
         n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513,
         n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521,
         n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529,
         n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537,
         n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545,
         n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553,
         n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561,
         n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569,
         n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577,
         n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585,
         n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593,
         n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601,
         n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609,
         n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617,
         n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625,
         n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633,
         n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641,
         n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649,
         n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657,
         n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665,
         n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673,
         n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681,
         n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689,
         n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697,
         n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705,
         n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713,
         n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721,
         n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729,
         n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737,
         n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745,
         n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753,
         n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761,
         n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769,
         n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777,
         n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785,
         n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793,
         n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801,
         n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809,
         n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817,
         n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825,
         n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833,
         n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841,
         n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849,
         n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857,
         n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865,
         n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873,
         n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881,
         n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889,
         n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897,
         n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905,
         n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913,
         n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921,
         n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929,
         n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937,
         n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945,
         n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953,
         n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961,
         n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969,
         n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977,
         n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985,
         n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993,
         n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001,
         n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009,
         n16010, n16011, n16012, n16013, n16014, n16015, n16016, n16017,
         n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16025,
         n16026, n16027, n16028, n16029, n16030, n16031, n16032, n16033,
         n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16041,
         n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049,
         n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057,
         n16058, n16059, n16060, n16061, n16062, n16063, n16064, n16065,
         n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073,
         n16074, n16075, n16076, n16077, n16078, n16079, n16080, n16081,
         n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089,
         n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097,
         n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105,
         n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113,
         n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121,
         n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129,
         n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137,
         n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145,
         n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153,
         n16154, n16156, n16157, n16158, n16159, n16160, n16161, n16162,
         n16163, n16164, n16165, n16166, n16167, n16168, n16169, n16170,
         n16171, n16172, n16173, n16174, n16175, n16176, n16177, n16178,
         n16179, n16180, n16181, n16182, n16183, n16184, n16185, n16186,
         n16187, n16188, n16189, n16190, n16191, n16192, n16193, n16194,
         n16195, n16196, n16197, n16198, n16199, n16200, n16201, n16202,
         n16203, n16204, n16205, n16206, n16207, n16208, n16209, n16210,
         n16211, n16212, n16213, n16214, n16215, n16216, n16217, n16218,
         n16219, n16220, n16221, n16222, n16223, n16224, n16225, n16226,
         n16227, n16228, n16229, n16230, n16231, n16232, n16233, n16234,
         n16235, n16236, n16237, n16238, n16239, n16240, n16241, n16242,
         n16243, n16244, n16245, n16246, n16247, n16248, n16249, n16250,
         n16251, n16252, n16253, n16254, n16255, n16256, n16257, n16258,
         n16259, n16260, n16261, n16262, n16263, n16264, n16265, n16266,
         n16267, n16268, n16269, n16270, n16271, n16272, n16273, n16274,
         n16275, n16276, n16277, n16278, n16279, n16280, n16281, n16282,
         n16283, n16284, n16285, n16286, n16287, n16288, n16289, n16290,
         n16291, n16292, n16293, n16294, n16295, n16296, n16297, n16298,
         n16299, n16300, n16301, n16302, n16303, n16304, n16305, n16306,
         n16307, n16308, n16309, n16310, n16311, n16312, n16313, n16314,
         n16315, n16316, n16317, n16318, n16319, n16320, n16321, n16322,
         n16323, n16324, n16325, n16326, n16327, n16328, n16329, n16330,
         n16331, n16332, n16333, n16334, n16335, n16336, n16337, n16338,
         n16339, n16340, n16341, n16342, n16343, n16344, n16345, n16346,
         n16347, n16348, n16349, n16350, n16351, n16352, n16353, n16354,
         n16355, n16356, n16357, n16358, n16359, n16360, n16361, n16362,
         n16363, n16364, n16365, n16366, n16367, n16368, n16369, n16370,
         n16371, n16372, n16373, n16374, n16375, n16376, n16377, n16378,
         n16379, n16380, n16381, n16382, n16383, n16384, n16385, n16386,
         n16387, n16388, n16389, n16390, n16391, n16392, n16393, n16394,
         n16395, n16396, n16397, n16398, n16399, n16400, n16401, n16402,
         n16403, n16404, n16405, n16406, n16407, n16408, n16409, n16410,
         n16411, n16412, n16413, n16414, n16415, n16416, n16417, n16418,
         n16419, n16420, n16421, n16422, n16423, n16424, n16425, n16426,
         n16427, n16428, n16429, n16430, n16431, n16432, n16433, n16434,
         n16435, n16436, n16437, n16438, n16439, n16440, n16441, n16442,
         n16443, n16444, n16445, n16446, n16447, n16448, n16449, n16450,
         n16451, n16452, n16453, n16454, n16455, n16456, n16457, n16458,
         n16459, n16460, n16461, n16462, n16463, n16464, n16465, n16466,
         n16467, n16468, n16469, n16470, n16471, n16472, n16473, n16474,
         n16475, n16476, n16477, n16478, n16479, n16480, n16481, n16482,
         n16483, n16484, n16485, n16486, n16487, n16488, n16489, n16490,
         n16491, n16492, n16493, n16494, n16495, n16496, n16497, n16498,
         n16499, n16500, n16501, n16502, n16503, n16504, n16505, n16506,
         n16507, n16508, n16509, n16510, n16511, n16512, n16513, n16514,
         n16515, n16516, n16517, n16518, n16519, n16520, n16521, n16522,
         n16523, n16524, n16525, n16526, n16527, n16528, n16529, n16530,
         n16531, n16532, n16533, n16534, n16535, n16536, n16537, n16538,
         n16539, n16540, n16541, n16542, n16543, n16544, n16545, n16546,
         n16547, n16548, n16549, n16550, n16551, n16552, n16553, n16554,
         n16555, n16556, n16557, n16558, n16559, n16560, n16561, n16562,
         n16563, n16564, n16565, n16566, n16567, n16568, n16569, n16570,
         n16571, n16572, n16573, n16574, n16575, n16576, n16577, n16578,
         n16579, n16580, n16581, n16582, n16583, n16584, n16585, n16586,
         n16587, n16588, n16589, n16590, n16591, n16592, n16593, n16594,
         n16595, n16596, n16597, n16598, n16599, n16600, n16601, n16602,
         n16603, n16604, n16605, n16606, n16607, n16608, n16609, n16610,
         n16611, n16612, n16613, n16614, n16615, n16616, n16617, n16618,
         n16619, n16620, n16621, n16622, n16623, n16624, n16625, n16626,
         n16627, n16628, n16629, n16630, n16631, n16632, n16633, n16634,
         n16635, n16636, n16637, n16638, n16639, n16640, n16641, n16642,
         n16643, n16644, n16645, n16646, n16647, n16648, n16649, n16650,
         n16651, n16652, n16653, n16654, n16655, n16656, n16657, n16658,
         n16659, n16660, n16661, n16662, n16663, n16664, n16665, n16666,
         n16667, n16668, n16669, n16670, n16671, n16672, n16673, n16674,
         n16675, n16676, n16677, n16678, n16679, n16680, n16681, n16682,
         n16683, n16684, n16685, n16686, n16687, n16688, n16689, n16690,
         n16691, n16692, n16693, n16694, n16695, n16696, n16697, n16698,
         n16699, n16700, n16701, n16702, n16703, n16704, n16705, n16706,
         n16707, n16708, n16709, n16710, n16711, n16712, n16713, n16714,
         n16715, n16716, n16717, n16718, n16719, n16720, n16721, n16722,
         n16723, n16724, n16725, n16726, n16727, n16728, n16729, n16730,
         n16731, n16732, n16733, n16734, n16735, n16736, n16737, n16738,
         n16739, n16740, n16741, n16742, n16743, n16744, n16745, n16746,
         n16747, n16748, n16749, n16750, n16751, n16752;

  NAND2_X1 U7511 ( .A1(n10429), .A2(n15988), .ZN(n16464) );
  CLKBUF_X2 U7512 ( .A(n11068), .Z(n14936) );
  INV_X1 U7513 ( .A(n13555), .ZN(n14139) );
  NAND2_X1 U7515 ( .A1(n8984), .A2(n9844), .ZN(n13494) );
  BUF_X2 U7516 ( .A(n9253), .Z(n7411) );
  CLKBUF_X2 U7517 ( .A(n9788), .Z(n10847) );
  INV_X1 U7518 ( .A(n10418), .ZN(n13566) );
  AND2_X1 U7519 ( .A1(n9758), .A2(n9759), .ZN(n9884) );
  INV_X1 U7520 ( .A(n13612), .ZN(n13782) );
  INV_X1 U7521 ( .A(n13782), .ZN(n13735) );
  NOR2_X1 U7522 ( .A1(n15339), .A2(n8752), .ZN(n8751) );
  NAND2_X1 U7523 ( .A1(n14112), .A2(n14921), .ZN(n8984) );
  AND4_X1 U7524 ( .A1(n8881), .A2(n8880), .A3(n8879), .A4(n8352), .ZN(n7462)
         );
  AOI22_X1 U7525 ( .A1(n15190), .A2(n15164), .B1(n15163), .B2(n15195), .ZN(
        n15180) );
  INV_X2 U7526 ( .A(n10271), .ZN(n7413) );
  INV_X2 U7527 ( .A(n12940), .ZN(n7412) );
  INV_X1 U7528 ( .A(n9874), .ZN(n9844) );
  INV_X1 U7529 ( .A(n13491), .ZN(n13480) );
  INV_X2 U7530 ( .A(n8976), .ZN(n13247) );
  INV_X1 U7531 ( .A(n14929), .ZN(n14959) );
  OAI21_X1 U7532 ( .B1(n12499), .B2(n7540), .A(n7970), .ZN(n15316) );
  NAND2_X2 U7533 ( .A1(n10090), .A2(n10089), .ZN(n11062) );
  NAND2_X1 U7534 ( .A1(n10626), .A2(n10625), .ZN(n10870) );
  AOI21_X1 U7535 ( .B1(n9399), .B2(n11935), .A(n12294), .ZN(n10319) );
  NAND2_X1 U7536 ( .A1(n8045), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8924) );
  CLKBUF_X3 U7537 ( .A(n13247), .Z(n7416) );
  INV_X1 U7538 ( .A(n15362), .ZN(n15353) );
  INV_X1 U7539 ( .A(n10817), .ZN(n12720) );
  NAND2_X1 U7540 ( .A1(n15408), .A2(n15161), .ZN(n7410) );
  BUF_X4 U7541 ( .A(n8995), .Z(n9335) );
  INV_X1 U7542 ( .A(n10998), .ZN(n9354) );
  NAND2_X2 U7543 ( .A1(n10053), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9996) );
  OAI21_X2 U7544 ( .B1(n10554), .B2(n9459), .A(n11503), .ZN(n11661) );
  NOR2_X2 U7545 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n9758) );
  NOR2_X2 U7546 ( .A1(n15148), .A2(n8758), .ZN(n8757) );
  OR2_X2 U7547 ( .A1(n10430), .A2(n16466), .ZN(n13669) );
  NAND2_X1 U7548 ( .A1(n8890), .A2(n8891), .ZN(n9253) );
  XNOR2_X2 U7549 ( .A(n8924), .B(n8923), .ZN(n14921) );
  AOI21_X1 U7550 ( .B1(n15911), .B2(n15774), .A(n15773), .ZN(n15889) );
  NAND2_X1 U7551 ( .A1(n13258), .A2(n13257), .ZN(n15184) );
  AND2_X1 U7552 ( .A1(n8292), .A2(n8295), .ZN(n15001) );
  NAND2_X1 U7553 ( .A1(n12781), .A2(n12780), .ZN(n16059) );
  NAND2_X1 U7554 ( .A1(n12972), .A2(n12971), .ZN(n15304) );
  NAND2_X1 U7555 ( .A1(n12730), .A2(n12729), .ZN(n16078) );
  NAND2_X1 U7556 ( .A1(n12542), .A2(n12541), .ZN(n16085) );
  AND4_X2 U7557 ( .A1(n9257), .A2(n9256), .A3(n9255), .A4(n9254), .ZN(n14264)
         );
  AOI21_X1 U7558 ( .B1(n8006), .B2(n8663), .A(n8004), .ZN(n8003) );
  INV_X2 U7559 ( .A(n13048), .ZN(n11284) );
  NAND2_X1 U7560 ( .A1(n10379), .A2(n9565), .ZN(n10392) );
  NAND4_X1 U7561 ( .A1(n10361), .A2(n10360), .A3(n10359), .A4(n10358), .ZN(
        n10430) );
  NAND2_X1 U7562 ( .A1(n15043), .A2(n14937), .ZN(n9745) );
  INV_X2 U7563 ( .A(n13035), .ZN(n10581) );
  CLKBUF_X2 U7564 ( .A(n10396), .Z(n12862) );
  INV_X1 U7565 ( .A(n12946), .ZN(n12802) );
  INV_X4 U7566 ( .A(n10463), .ZN(n12053) );
  NAND4_X2 U7567 ( .A1(n9864), .A2(n9543), .A3(n8830), .A4(n8829), .ZN(n9929)
         );
  INV_X2 U7568 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n8829) );
  INV_X2 U7569 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  AOI211_X1 U7570 ( .C1(n13337), .C2(n13345), .A(n13342), .B(n13336), .ZN(
        n13349) );
  OR2_X1 U7571 ( .A1(n13346), .A2(n8013), .ZN(n8012) );
  AOI21_X1 U7572 ( .B1(n8559), .B2(n16561), .A(n8556), .ZN(n16014) );
  NAND2_X1 U7573 ( .A1(n7999), .A2(n7997), .ZN(n15799) );
  OR2_X1 U7574 ( .A1(n16036), .A2(n16035), .ZN(n16104) );
  AOI21_X1 U7575 ( .B1(n8098), .B2(n16561), .A(n8095), .ZN(n16023) );
  NAND2_X1 U7576 ( .A1(n7922), .A2(n7921), .ZN(n8503) );
  NAND2_X1 U7577 ( .A1(n8613), .A2(n8612), .ZN(n15801) );
  OR2_X1 U7578 ( .A1(n8841), .A2(n13803), .ZN(n8653) );
  AND2_X1 U7579 ( .A1(n13646), .A2(n13644), .ZN(n13636) );
  AOI21_X1 U7580 ( .B1(n7794), .B2(n7796), .A(n7793), .ZN(n7792) );
  NAND2_X1 U7581 ( .A1(n7525), .A2(n8689), .ZN(n8688) );
  NAND2_X1 U7582 ( .A1(n15613), .A2(n15614), .ZN(n15612) );
  NOR2_X1 U7583 ( .A1(n13604), .A2(n8402), .ZN(n13605) );
  NAND2_X1 U7584 ( .A1(n14162), .A2(n13355), .ZN(n13513) );
  INV_X1 U7585 ( .A(n8811), .ZN(n7793) );
  OAI22_X1 U7586 ( .A1(n15205), .A2(n15209), .B1(n15485), .B2(n15162), .ZN(
        n15190) );
  OAI21_X1 U7587 ( .B1(n15210), .B2(n7444), .A(n7548), .ZN(n7972) );
  OAI21_X1 U7588 ( .B1(n15168), .B2(n15166), .A(n15346), .ZN(n7863) );
  AOI21_X1 U7589 ( .B1(n8812), .B2(n8814), .A(n7529), .ZN(n8811) );
  AND2_X1 U7590 ( .A1(n8812), .A2(n7795), .ZN(n7794) );
  AND2_X1 U7591 ( .A1(n8614), .A2(n8406), .ZN(n8612) );
  AND2_X1 U7592 ( .A1(n15804), .A2(n7998), .ZN(n7997) );
  NOR4_X1 U7593 ( .A1(n15165), .A2(n15193), .A3(n15209), .A4(n13333), .ZN(
        n13335) );
  NAND2_X1 U7594 ( .A1(n15131), .A2(n7431), .ZN(n15240) );
  AOI21_X1 U7595 ( .B1(n7428), .B2(n15577), .A(n7544), .ZN(n7797) );
  OR2_X1 U7596 ( .A1(n15184), .A2(n15172), .ZN(n15166) );
  NAND2_X1 U7597 ( .A1(n13230), .A2(n13229), .ZN(n15386) );
  NAND2_X1 U7598 ( .A1(n13602), .A2(n13601), .ZN(n15786) );
  AOI211_X1 U7599 ( .C1(n16040), .C2(n16606), .A(n16039), .B(n16038), .ZN(
        n16041) );
  NAND2_X1 U7600 ( .A1(n15864), .A2(n16027), .ZN(n15848) );
  AOI21_X1 U7601 ( .B1(n15524), .B2(n11544), .A(n7632), .ZN(n16002) );
  OAI21_X1 U7602 ( .B1(n14192), .B2(n8138), .A(n8137), .ZN(n14172) );
  AND2_X1 U7603 ( .A1(n7952), .A2(n7435), .ZN(n7957) );
  XNOR2_X1 U7604 ( .A(n13250), .B(n13249), .ZN(n15519) );
  AOI21_X2 U7605 ( .B1(n13255), .B2(n11544), .A(n7612), .ZN(n15808) );
  XNOR2_X1 U7606 ( .A(n13246), .B(n13243), .ZN(n15524) );
  NAND2_X1 U7607 ( .A1(n13255), .A2(n12053), .ZN(n13258) );
  NAND2_X1 U7608 ( .A1(n8671), .A2(n8668), .ZN(n13250) );
  AND2_X1 U7609 ( .A1(n8296), .A2(n15763), .ZN(n15864) );
  NOR2_X1 U7610 ( .A1(n8634), .A2(n15872), .ZN(n8633) );
  NAND2_X1 U7611 ( .A1(n14970), .A2(n14969), .ZN(n14968) );
  AOI211_X1 U7612 ( .C1(n16040), .C2(n15894), .A(n16464), .B(n8296), .ZN(
        n16038) );
  AND2_X1 U7613 ( .A1(n8608), .A2(n7706), .ZN(n15890) );
  OR2_X1 U7614 ( .A1(n7960), .A2(n13768), .ZN(n7952) );
  NAND2_X1 U7615 ( .A1(n12917), .A2(n12916), .ZN(n15819) );
  NOR2_X1 U7616 ( .A1(n7443), .A2(n7708), .ZN(n7704) );
  NAND2_X1 U7617 ( .A1(n13194), .A2(n13193), .ZN(n15195) );
  OAI21_X1 U7618 ( .B1(n12653), .B2(n8677), .A(n8674), .ZN(n13246) );
  XNOR2_X1 U7619 ( .A(n12653), .B(n12652), .ZN(n13255) );
  NAND2_X1 U7620 ( .A1(n13199), .A2(n13198), .ZN(n15211) );
  NAND2_X1 U7621 ( .A1(n12638), .A2(n12637), .ZN(n12653) );
  NAND2_X1 U7622 ( .A1(n12894), .A2(n12893), .ZN(n16021) );
  AND2_X1 U7623 ( .A1(n15156), .A2(n7565), .ZN(n7877) );
  OR2_X1 U7624 ( .A1(n7726), .A2(n7725), .ZN(n15894) );
  NAND2_X1 U7625 ( .A1(n12878), .A2(n12877), .ZN(n15738) );
  XNOR2_X1 U7626 ( .A(n12915), .B(n12914), .ZN(n15531) );
  XNOR2_X1 U7627 ( .A(n16046), .B(n15761), .ZN(n15891) );
  NAND2_X1 U7628 ( .A1(n12857), .A2(n12856), .ZN(n15869) );
  NAND2_X1 U7629 ( .A1(n8034), .A2(n8022), .ZN(n12915) );
  XNOR2_X1 U7630 ( .A(n15424), .B(n15286), .ZN(n15269) );
  NAND2_X1 U7631 ( .A1(n15322), .A2(n15151), .ZN(n15305) );
  NAND2_X1 U7632 ( .A1(n13156), .A2(n13155), .ZN(n15256) );
  NOR2_X1 U7633 ( .A1(n8391), .A2(n7620), .ZN(n8022) );
  XNOR2_X1 U7634 ( .A(n12876), .B(n12875), .ZN(n15535) );
  NAND2_X1 U7635 ( .A1(n12629), .A2(n12628), .ZN(n12876) );
  XNOR2_X1 U7636 ( .A(n12855), .B(n12854), .ZN(n15538) );
  XNOR2_X1 U7637 ( .A(n12813), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n16141) );
  AND2_X1 U7638 ( .A1(n14294), .A2(n14293), .ZN(n14296) );
  OAI21_X1 U7639 ( .B1(n8751), .B2(n7465), .A(n15317), .ZN(n7971) );
  OAI21_X1 U7640 ( .B1(n12829), .B2(n12622), .A(n7432), .ZN(n8084) );
  NAND2_X1 U7641 ( .A1(n12196), .A2(n12209), .ZN(n12449) );
  XNOR2_X1 U7642 ( .A(n12830), .B(SI_22_), .ZN(n12829) );
  OAI21_X1 U7643 ( .B1(n12471), .B2(n8710), .A(n8708), .ZN(n15149) );
  XNOR2_X1 U7644 ( .A(n15304), .B(n14936), .ZN(n12975) );
  NAND2_X1 U7645 ( .A1(n12798), .A2(n12797), .ZN(n15906) );
  NAND2_X1 U7646 ( .A1(n12960), .A2(n12959), .ZN(n15291) );
  NAND2_X1 U7647 ( .A1(n7932), .A2(n12175), .ZN(n12212) );
  AOI21_X1 U7648 ( .B1(n7429), .B2(n8602), .A(n7499), .ZN(n7718) );
  NAND2_X1 U7649 ( .A1(n7672), .A2(n12003), .ZN(n12315) );
  OAI21_X1 U7650 ( .B1(n13876), .B2(n10505), .A(n13874), .ZN(n8726) );
  NAND2_X1 U7651 ( .A1(n12076), .A2(n12075), .ZN(n12175) );
  NAND2_X1 U7652 ( .A1(n13876), .A2(n10505), .ZN(n8725) );
  OR2_X1 U7653 ( .A1(n12716), .A2(n12715), .ZN(n8855) );
  XNOR2_X1 U7654 ( .A(n16068), .B(n15954), .ZN(n15933) );
  NAND2_X1 U7655 ( .A1(n12337), .A2(n12336), .ZN(n12555) );
  AND2_X1 U7656 ( .A1(n12696), .A2(n12065), .ZN(n12076) );
  NAND2_X1 U7657 ( .A1(n12599), .A2(n12598), .ZN(n15329) );
  NAND2_X1 U7658 ( .A1(n11999), .A2(n11998), .ZN(n12090) );
  NAND2_X1 U7659 ( .A1(n8844), .A2(n12370), .ZN(n12511) );
  NAND2_X1 U7660 ( .A1(n12497), .A2(n12496), .ZN(n12499) );
  XNOR2_X1 U7661 ( .A(n12369), .B(n12153), .ZN(n12969) );
  NAND2_X1 U7662 ( .A1(n7801), .A2(n7799), .ZN(n12711) );
  NAND2_X1 U7663 ( .A1(n7993), .A2(n12150), .ZN(n12369) );
  NAND2_X1 U7664 ( .A1(n8033), .A2(n11722), .ZN(n11764) );
  OAI211_X1 U7665 ( .C1(n8684), .C2(n8682), .A(n8680), .B(n14664), .ZN(n12368)
         );
  XNOR2_X1 U7666 ( .A(n12152), .B(n12151), .ZN(n12758) );
  XNOR2_X1 U7667 ( .A(n16078), .B(n15755), .ZN(n15981) );
  NAND2_X1 U7668 ( .A1(n8681), .A2(n12150), .ZN(n8680) );
  NAND2_X1 U7669 ( .A1(n12440), .A2(n12439), .ZN(n15444) );
  NAND2_X1 U7670 ( .A1(n8015), .A2(n12195), .ZN(n15146) );
  NOR2_X1 U7671 ( .A1(n12561), .A2(n16085), .ZN(n8310) );
  NAND2_X1 U7672 ( .A1(n12743), .A2(n12742), .ZN(n16074) );
  NAND2_X1 U7673 ( .A1(n8375), .A2(n11880), .ZN(n8684) );
  NOR2_X1 U7674 ( .A1(n12327), .A2(n13736), .ZN(n12347) );
  XNOR2_X1 U7675 ( .A(n8106), .B(n11742), .ZN(n12728) );
  NAND2_X1 U7676 ( .A1(n11574), .A2(n13585), .ZN(n11869) );
  OAI211_X1 U7677 ( .C1(n8816), .C2(n7780), .A(n7779), .B(n8064), .ZN(n12128)
         );
  NAND2_X1 U7678 ( .A1(n12539), .A2(n12053), .ZN(n8251) );
  OAI21_X1 U7679 ( .B1(n11158), .B2(n8661), .A(n8388), .ZN(n8106) );
  NAND2_X1 U7680 ( .A1(n7731), .A2(n7730), .ZN(n12327) );
  AND2_X1 U7681 ( .A1(n8382), .A2(SI_18_), .ZN(n8381) );
  INV_X1 U7682 ( .A(n12094), .ZN(n7731) );
  NAND2_X1 U7683 ( .A1(n8380), .A2(n8384), .ZN(n8063) );
  XNOR2_X1 U7684 ( .A(n11158), .B(n11159), .ZN(n12539) );
  NAND2_X1 U7685 ( .A1(n8383), .A2(SI_16_), .ZN(n8388) );
  NAND2_X1 U7686 ( .A1(n7728), .A2(n7727), .ZN(n12094) );
  XNOR2_X1 U7687 ( .A(n11161), .B(n11160), .ZN(n11158) );
  NAND2_X1 U7688 ( .A1(n11786), .A2(n11785), .ZN(n13102) );
  NAND2_X1 U7689 ( .A1(n11762), .A2(n11761), .ZN(n16700) );
  NAND2_X1 U7690 ( .A1(n11363), .A2(n11362), .ZN(n15368) );
  NAND2_X1 U7691 ( .A1(n11438), .A2(n11144), .ZN(n11345) );
  NAND2_X1 U7692 ( .A1(n11093), .A2(n11092), .ZN(n13083) );
  NAND2_X1 U7693 ( .A1(n8005), .A2(n8003), .ZN(n10617) );
  NOR2_X1 U7694 ( .A1(n9197), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n9217) );
  INV_X2 U7695 ( .A(n16625), .ZN(n7414) );
  NOR2_X2 U7696 ( .A1(n10095), .A2(P2_U3088), .ZN(n10096) );
  AND2_X1 U7697 ( .A1(n8289), .A2(n8007), .ZN(n8006) );
  INV_X1 U7698 ( .A(n12846), .ZN(n12921) );
  INV_X1 U7699 ( .A(n11828), .ZN(n16496) );
  NAND2_X1 U7700 ( .A1(n10655), .A2(n10654), .ZN(n16586) );
  INV_X1 U7701 ( .A(n16554), .ZN(n13677) );
  INV_X2 U7702 ( .A(n15677), .ZN(P1_U4016) );
  NAND4_X1 U7703 ( .A1(n8972), .A2(n8971), .A3(n8970), .A4(n8969), .ZN(n11534)
         );
  NAND2_X1 U7704 ( .A1(n8961), .A2(n8960), .ZN(n16497) );
  OAI211_X1 U7705 ( .C1(n10702), .C2(n9893), .A(n10363), .B(n7522), .ZN(n16466) );
  NAND2_X1 U7706 ( .A1(n7430), .A2(n9741), .ZN(n13024) );
  NAND2_X2 U7707 ( .A1(n10392), .A2(n10432), .ZN(n10271) );
  NAND2_X1 U7708 ( .A1(n10392), .A2(n13660), .ZN(n12940) );
  OAI211_X1 U7709 ( .C1(n10687), .C2(n12814), .A(n10686), .B(n10685), .ZN(
        n16527) );
  NAND2_X1 U7710 ( .A1(n7986), .A2(n7984), .ZN(n9917) );
  NAND4_X1 U7711 ( .A1(n10423), .A2(n10422), .A3(n10421), .A4(n10420), .ZN(
        n15690) );
  INV_X1 U7712 ( .A(n8980), .ZN(n9157) );
  NOR2_X1 U7713 ( .A1(n10447), .A2(n8397), .ZN(n8396) );
  NAND2_X2 U7714 ( .A1(n14911), .A2(n14915), .ZN(n10998) );
  NOR2_X2 U7715 ( .A1(n13624), .A2(n10401), .ZN(n16462) );
  NAND2_X1 U7716 ( .A1(n8112), .A2(n7512), .ZN(n9870) );
  AND2_X1 U7717 ( .A1(n9561), .A2(n9560), .ZN(n10379) );
  OAI211_X1 U7718 ( .C1(n10463), .C2(n10683), .A(n9785), .B(n9784), .ZN(n13035) );
  NAND2_X1 U7719 ( .A1(n9349), .A2(n9348), .ZN(n10835) );
  INV_X1 U7720 ( .A(n9783), .ZN(n12597) );
  INV_X1 U7721 ( .A(n8891), .ZN(n14915) );
  NOR2_X1 U7722 ( .A1(n7988), .A2(n9896), .ZN(n7987) );
  OAI21_X1 U7723 ( .B1(n13247), .B2(n9923), .A(n8109), .ZN(n9939) );
  XNOR2_X1 U7724 ( .A(n9956), .B(SI_8_), .ZN(n9953) );
  INV_X1 U7725 ( .A(n8890), .ZN(n14911) );
  INV_X1 U7726 ( .A(n13606), .ZN(n15733) );
  NAND2_X2 U7727 ( .A1(n10356), .A2(n10355), .ZN(n12946) );
  AND2_X2 U7728 ( .A1(n9720), .A2(n7460), .ZN(n8082) );
  AND2_X1 U7729 ( .A1(n10380), .A2(n16128), .ZN(n9565) );
  INV_X1 U7730 ( .A(n10355), .ZN(n12655) );
  AND2_X2 U7731 ( .A1(n9704), .A2(n9705), .ZN(n9786) );
  INV_X1 U7732 ( .A(n13555), .ZN(n14112) );
  CLKBUF_X3 U7733 ( .A(n9730), .Z(n13342) );
  NAND2_X2 U7734 ( .A1(n9729), .A2(n9728), .ZN(n13345) );
  XNOR2_X1 U7735 ( .A(n7719), .B(P1_IR_REG_29__SCAN_IN), .ZN(n10355) );
  NAND3_X1 U7736 ( .A1(n8637), .A2(n8636), .A3(n8638), .ZN(n13607) );
  XNOR2_X1 U7737 ( .A(n8297), .B(n9995), .ZN(n16240) );
  XNOR2_X1 U7738 ( .A(n9898), .B(SI_5_), .ZN(n9896) );
  XNOR2_X1 U7739 ( .A(n10249), .B(P1_IR_REG_19__SCAN_IN), .ZN(n13606) );
  NAND2_X1 U7740 ( .A1(n10246), .A2(n10245), .ZN(n13610) );
  NAND2_X1 U7741 ( .A1(n7720), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7719) );
  NAND2_X1 U7742 ( .A1(n9997), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8297) );
  NAND2_X1 U7743 ( .A1(n16117), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10250) );
  OAI21_X1 U7744 ( .B1(n9563), .B2(P1_IR_REG_25__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9562) );
  XNOR2_X1 U7745 ( .A(n8527), .B(n9702), .ZN(n15526) );
  INV_X2 U7746 ( .A(n15528), .ZN(n15545) );
  OR2_X1 U7747 ( .A1(n9553), .A2(n8642), .ZN(n8637) );
  XNOR2_X1 U7748 ( .A(n9717), .B(n9716), .ZN(n10090) );
  OAI21_X1 U7749 ( .B1(n9874), .B2(n9878), .A(n8107), .ZN(n9898) );
  NAND2_X1 U7750 ( .A1(n9727), .A2(P2_IR_REG_20__SCAN_IN), .ZN(n9728) );
  NAND2_X1 U7751 ( .A1(n7461), .A2(n9713), .ZN(n10089) );
  INV_X1 U7752 ( .A(n9554), .ZN(n9553) );
  NAND2_X1 U7753 ( .A1(n15520), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8527) );
  OR2_X1 U7754 ( .A1(n9714), .A2(n9715), .ZN(n9717) );
  OR2_X1 U7755 ( .A1(n9554), .A2(n9993), .ZN(n9563) );
  CLKBUF_X1 U7756 ( .A(n8877), .Z(n8044) );
  AND2_X1 U7757 ( .A1(n9994), .A2(n9995), .ZN(n8839) );
  AND2_X1 U7758 ( .A1(n8743), .A2(n8876), .ZN(n8742) );
  AND2_X1 U7759 ( .A1(n8354), .A2(n8882), .ZN(n8353) );
  AND2_X1 U7760 ( .A1(n7468), .A2(n9578), .ZN(n8693) );
  AND4_X1 U7761 ( .A1(n9701), .A2(n9884), .A3(n10147), .A4(n9716), .ZN(n8692)
         );
  AND4_X1 U7762 ( .A1(n9579), .A2(n9698), .A3(n9697), .A4(n9696), .ZN(n9701)
         );
  INV_X1 U7763 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n8926) );
  INV_X2 U7764 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n9543) );
  INV_X1 U7765 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n8352) );
  NOR2_X1 U7766 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n10635) );
  INV_X1 U7767 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n9883) );
  INV_X1 U7768 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n14617) );
  INV_X1 U7769 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n9552) );
  INV_X1 U7770 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n9991) );
  INV_X1 U7771 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n16405) );
  INV_X1 U7772 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n9556) );
  NOR2_X1 U7773 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n9545) );
  INV_X1 U7774 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n9697) );
  OAI21_X2 U7775 ( .B1(n7983), .B2(n7980), .A(n7491), .ZN(n12497) );
  NAND2_X1 U7776 ( .A1(n8376), .A2(n8684), .ZN(n7993) );
  INV_X1 U7777 ( .A(n7972), .ZN(n15194) );
  OR2_X2 U7778 ( .A1(n15885), .A2(n15884), .ZN(n7680) );
  AOI21_X2 U7779 ( .B1(n15889), .B2(n15891), .A(n15776), .ZN(n15885) );
  NAND2_X1 U7780 ( .A1(n15799), .A2(n15782), .ZN(n15784) );
  AND2_X1 U7781 ( .A1(n8755), .A2(n8756), .ZN(n8752) );
  OAI22_X2 U7782 ( .A1(n11161), .A2(n7608), .B1(n8385), .B2(n8386), .ZN(n8384)
         );
  XNOR2_X1 U7783 ( .A(n16040), .B(n15777), .ZN(n15884) );
  OR2_X2 U7784 ( .A1(n9371), .A2(n14264), .ZN(n13447) );
  NOR2_X2 U7785 ( .A1(n9929), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n9875) );
  AOI211_X1 U7786 ( .C1(n16466), .C2(n16606), .A(n16482), .B(n16485), .ZN(
        n16473) );
  INV_X1 U7787 ( .A(n16466), .ZN(n16480) );
  XNOR2_X2 U7788 ( .A(n15146), .B(n15342), .ZN(n15148) );
  NAND2_X2 U7789 ( .A1(n10352), .A2(n13660), .ZN(n10817) );
  XNOR2_X2 U7790 ( .A(n9974), .B(SI_9_), .ZN(n9972) );
  XNOR2_X2 U7791 ( .A(n9996), .B(n7965), .ZN(n10019) );
  CLKBUF_X1 U7792 ( .A(n16240), .Z(n7417) );
  NAND2_X1 U7793 ( .A1(n16120), .A2(n12655), .ZN(n7418) );
  NAND2_X1 U7794 ( .A1(n16053), .A2(n15772), .ZN(n8609) );
  INV_X1 U7795 ( .A(n13485), .ZN(n13545) );
  NOR2_X1 U7796 ( .A1(n13325), .A2(n8705), .ZN(n8704) );
  AND2_X1 U7797 ( .A1(n13324), .A2(n12135), .ZN(n8705) );
  NAND2_X1 U7798 ( .A1(n11882), .A2(n8683), .ZN(n8681) );
  INV_X1 U7799 ( .A(n12151), .ZN(n8683) );
  AND4_X2 U7800 ( .A1(n8742), .A2(n8353), .A3(n8883), .A4(n8877), .ZN(n8171)
         );
  NOR2_X1 U7801 ( .A1(n9987), .A2(P1_IR_REG_22__SCAN_IN), .ZN(n9566) );
  NAND2_X1 U7802 ( .A1(n9553), .A2(n7593), .ZN(n9987) );
  NAND2_X1 U7803 ( .A1(n14911), .A2(n8891), .ZN(n8979) );
  INV_X1 U7804 ( .A(n13494), .ZN(n13504) );
  AOI21_X1 U7805 ( .B1(n7927), .B2(n7925), .A(n7538), .ZN(n7924) );
  INV_X1 U7806 ( .A(n7927), .ZN(n7926) );
  NAND2_X1 U7807 ( .A1(n15916), .A2(n7528), .ZN(n8608) );
  AND2_X1 U7808 ( .A1(n13020), .A2(n13019), .ZN(n13029) );
  OAI21_X1 U7809 ( .B1(n8651), .B2(n13687), .A(n13686), .ZN(n13696) );
  NAND2_X1 U7810 ( .A1(n7748), .A2(n7747), .ZN(n7746) );
  NAND2_X1 U7811 ( .A1(n13056), .A2(n13055), .ZN(n7747) );
  OAI21_X1 U7812 ( .B1(n13055), .B2(n13056), .A(n8797), .ZN(n7748) );
  AND2_X1 U7813 ( .A1(n7754), .A2(n8032), .ZN(n7753) );
  INV_X1 U7814 ( .A(n13103), .ZN(n8032) );
  NAND2_X1 U7815 ( .A1(n7755), .A2(n13104), .ZN(n7754) );
  OAI21_X1 U7816 ( .B1(n7766), .B2(n7765), .A(n7546), .ZN(n13127) );
  OAI21_X1 U7817 ( .B1(n13116), .B2(n13115), .A(n7515), .ZN(n7766) );
  AOI21_X1 U7818 ( .B1(n13116), .B2(n13115), .A(n13114), .ZN(n7765) );
  NAND2_X1 U7819 ( .A1(n7944), .A2(n13755), .ZN(n7943) );
  INV_X1 U7820 ( .A(n13768), .ZN(n7955) );
  INV_X1 U7821 ( .A(n13177), .ZN(n8796) );
  INV_X1 U7822 ( .A(n10215), .ZN(n8397) );
  AND2_X1 U7823 ( .A1(n13479), .A2(n13478), .ZN(n13482) );
  INV_X1 U7824 ( .A(n9940), .ZN(n7991) );
  INV_X1 U7825 ( .A(n11950), .ZN(n8197) );
  NAND2_X1 U7826 ( .A1(n8884), .A2(n8749), .ZN(n8748) );
  INV_X1 U7827 ( .A(n8998), .ZN(n8877) );
  INV_X1 U7828 ( .A(n13254), .ZN(n8689) );
  NOR2_X1 U7829 ( .A1(n11248), .A2(n7868), .ZN(n7867) );
  NAND2_X1 U7830 ( .A1(n11161), .A2(n7454), .ZN(n8382) );
  NOR2_X1 U7831 ( .A1(n11742), .A2(n11159), .ZN(n8386) );
  INV_X1 U7832 ( .A(n11741), .ZN(n8385) );
  NAND2_X2 U7833 ( .A1(n10870), .A2(n10869), .ZN(n11161) );
  NAND2_X1 U7834 ( .A1(n13544), .A2(n13515), .ZN(n8359) );
  AND2_X1 U7835 ( .A1(n13545), .A2(n8577), .ZN(n8576) );
  AND2_X1 U7836 ( .A1(n14205), .A2(n7493), .ZN(n8577) );
  AND2_X1 U7837 ( .A1(n8580), .A2(n8579), .ZN(n13521) );
  NAND2_X1 U7838 ( .A1(n14840), .A2(n14151), .ZN(n8580) );
  NAND2_X1 U7839 ( .A1(n13510), .A2(n13507), .ZN(n8579) );
  OR2_X1 U7840 ( .A1(n9657), .A2(n11524), .ZN(n8191) );
  OAI21_X1 U7841 ( .B1(n11516), .B2(n7848), .A(n7847), .ZN(n8184) );
  NAND2_X1 U7842 ( .A1(n7849), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n7848) );
  NAND2_X1 U7843 ( .A1(n9658), .A2(n7849), .ZN(n7847) );
  INV_X1 U7844 ( .A(n8185), .ZN(n7849) );
  NAND2_X1 U7845 ( .A1(n16428), .A2(n8186), .ZN(n8185) );
  NAND2_X1 U7846 ( .A1(n7605), .A2(n11613), .ZN(n8186) );
  AND2_X1 U7847 ( .A1(n9662), .A2(n7814), .ZN(n7810) );
  NAND2_X1 U7848 ( .A1(n7549), .A2(n9498), .ZN(n8144) );
  INV_X1 U7849 ( .A(n8149), .ZN(n8147) );
  INV_X1 U7850 ( .A(n10835), .ZN(n13357) );
  INV_X1 U7851 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n8884) );
  AND2_X1 U7852 ( .A1(n9191), .A2(n9168), .ZN(n8354) );
  INV_X1 U7853 ( .A(n8570), .ZN(n8569) );
  OAI21_X1 U7854 ( .B1(n9118), .B2(n8571), .A(n9134), .ZN(n8570) );
  AND2_X1 U7855 ( .A1(n8745), .A2(n8878), .ZN(n8743) );
  INV_X1 U7856 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n8878) );
  INV_X1 U7857 ( .A(n15526), .ZN(n9705) );
  NOR2_X1 U7858 ( .A1(n15386), .A2(n15184), .ZN(n8317) );
  NAND2_X1 U7859 ( .A1(n8696), .A2(n7410), .ZN(n8695) );
  INV_X1 U7860 ( .A(n12587), .ZN(n8758) );
  INV_X1 U7861 ( .A(n13345), .ZN(n13307) );
  INV_X1 U7862 ( .A(n7971), .ZN(n7970) );
  OR2_X1 U7863 ( .A1(n8779), .A2(n8777), .ZN(n8776) );
  INV_X1 U7864 ( .A(n12465), .ZN(n8777) );
  NOR2_X1 U7865 ( .A1(n8778), .A2(n7982), .ZN(n7981) );
  INV_X1 U7866 ( .A(n12134), .ZN(n7982) );
  NAND2_X1 U7867 ( .A1(n13325), .A2(n12465), .ZN(n8778) );
  NOR2_X1 U7868 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n8312) );
  AND3_X1 U7869 ( .A1(n9577), .A2(n9576), .A3(n9575), .ZN(n10147) );
  NOR2_X1 U7870 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n9577) );
  NOR2_X1 U7871 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n9575) );
  NOR2_X1 U7872 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n9576) );
  AND4_X1 U7873 ( .A1(n9574), .A2(n9573), .A3(n9572), .A4(n9883), .ZN(n9578)
         );
  NOR2_X1 U7874 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n9573) );
  NOR2_X1 U7875 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n9572) );
  INV_X1 U7876 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n9696) );
  INV_X1 U7877 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n9698) );
  NOR2_X1 U7878 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n9724) );
  INV_X1 U7879 ( .A(n8813), .ZN(n8812) );
  OAI21_X1 U7880 ( .B1(n15614), .B2(n8814), .A(n15585), .ZN(n8813) );
  OR2_X1 U7881 ( .A1(n13637), .A2(n13639), .ZN(n13800) );
  AOI21_X1 U7882 ( .B1(n15814), .B2(n8002), .A(n8001), .ZN(n8000) );
  INV_X1 U7883 ( .A(n15780), .ZN(n8001) );
  INV_X1 U7884 ( .A(n15779), .ZN(n8002) );
  NOR2_X1 U7885 ( .A1(n15933), .A2(n8548), .ZN(n8547) );
  INV_X1 U7886 ( .A(n15769), .ZN(n8548) );
  OR2_X1 U7887 ( .A1(n16090), .A2(n12713), .ZN(n12538) );
  AND2_X1 U7888 ( .A1(n13587), .A2(n11868), .ZN(n8635) );
  INV_X1 U7889 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n8644) );
  NAND2_X1 U7890 ( .A1(n16345), .A2(n16346), .ZN(n16347) );
  NAND2_X1 U7891 ( .A1(n12296), .A2(n8088), .ZN(n12416) );
  NAND2_X1 U7892 ( .A1(n9464), .A2(n12420), .ZN(n8088) );
  XNOR2_X1 U7893 ( .A(n9450), .B(n16524), .ZN(n9456) );
  AND2_X1 U7894 ( .A1(n8725), .A2(n7892), .ZN(n7887) );
  AND2_X1 U7895 ( .A1(n13835), .A2(n7895), .ZN(n7892) );
  AOI21_X1 U7896 ( .B1(n14165), .B2(n9326), .A(n8896), .ZN(n11040) );
  NOR2_X1 U7897 ( .A1(n10920), .A2(n9024), .ZN(n10919) );
  AND2_X1 U7898 ( .A1(n7818), .A2(n7817), .ZN(n10904) );
  INV_X1 U7899 ( .A(n10905), .ZN(n7817) );
  OR2_X1 U7900 ( .A1(n11952), .A2(n7740), .ZN(n7737) );
  INV_X1 U7901 ( .A(n12157), .ZN(n7740) );
  NOR2_X1 U7902 ( .A1(n13993), .A2(n14024), .ZN(n14010) );
  INV_X1 U7903 ( .A(n14132), .ZN(n14147) );
  NAND2_X1 U7904 ( .A1(n8422), .A2(n14117), .ZN(n14131) );
  OR2_X1 U7905 ( .A1(n14157), .A2(n14163), .ZN(n14160) );
  AOI21_X1 U7906 ( .B1(n14187), .B2(n9326), .A(n9317), .ZN(n14198) );
  AOI21_X1 U7907 ( .B1(n14217), .B2(n14216), .A(n7899), .ZN(n14206) );
  AND2_X1 U7908 ( .A1(n13847), .A2(n14232), .ZN(n7899) );
  INV_X1 U7909 ( .A(n8139), .ZN(n8138) );
  AOI21_X1 U7910 ( .B1(n8141), .B2(n8139), .A(n7851), .ZN(n8137) );
  NAND2_X1 U7911 ( .A1(n14903), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8886) );
  XNOR2_X1 U7912 ( .A(n8889), .B(P3_IR_REG_29__SCAN_IN), .ZN(n8891) );
  AOI21_X1 U7913 ( .B1(n8122), .B2(n9319), .A(n8121), .ZN(n9334) );
  AND2_X1 U7914 ( .A1(n16123), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n8121) );
  NOR2_X1 U7915 ( .A1(n11798), .A2(n8524), .ZN(n8523) );
  INV_X1 U7916 ( .A(n11796), .ZN(n8524) );
  AOI21_X1 U7917 ( .B1(n7924), .B2(n7926), .A(n8508), .ZN(n7921) );
  NAND2_X1 U7918 ( .A1(n14977), .A2(n7924), .ZN(n7922) );
  NAND2_X1 U7919 ( .A1(n14968), .A2(n7471), .ZN(n8277) );
  NAND2_X1 U7920 ( .A1(n12449), .A2(n12448), .ZN(n12450) );
  NAND2_X1 U7921 ( .A1(n8499), .A2(n8497), .ZN(n11058) );
  NOR2_X1 U7922 ( .A1(n8498), .A2(n10660), .ZN(n8497) );
  AND2_X1 U7923 ( .A1(n8082), .A2(n13342), .ZN(n10077) );
  AND2_X1 U7924 ( .A1(n13350), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9818) );
  OR2_X1 U7925 ( .A1(n8315), .A2(n15468), .ZN(n8314) );
  NAND2_X1 U7926 ( .A1(n15240), .A2(n8768), .ZN(n15224) );
  NOR2_X1 U7927 ( .A1(n15220), .A2(n8769), .ZN(n8768) );
  INV_X1 U7928 ( .A(n15133), .ZN(n8769) );
  AND2_X1 U7929 ( .A1(n15281), .A2(n15154), .ZN(n15265) );
  AOI21_X1 U7930 ( .B1(n15149), .B2(n15148), .A(n15147), .ZN(n15340) );
  NAND2_X1 U7931 ( .A1(n7879), .A2(n7506), .ZN(n12470) );
  INV_X1 U7932 ( .A(n13327), .ZN(n7878) );
  AND2_X1 U7933 ( .A1(n16704), .A2(n12371), .ZN(n9829) );
  NAND2_X2 U7934 ( .A1(n11062), .A2(n9844), .ZN(n9783) );
  NAND2_X1 U7935 ( .A1(n11062), .A2(n7416), .ZN(n10463) );
  OR2_X1 U7936 ( .A1(n15534), .A2(n9810), .ZN(n16147) );
  XNOR2_X1 U7937 ( .A(n9703), .B(P2_IR_REG_29__SCAN_IN), .ZN(n9704) );
  NAND2_X1 U7938 ( .A1(n7461), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9703) );
  AND2_X1 U7939 ( .A1(n8821), .A2(n8819), .ZN(n8818) );
  INV_X1 U7940 ( .A(n11713), .ZN(n8819) );
  INV_X1 U7941 ( .A(n12757), .ZN(n7790) );
  NOR2_X1 U7942 ( .A1(n15891), .A2(n7707), .ZN(n7706) );
  INV_X1 U7943 ( .A(n8606), .ZN(n7707) );
  NAND2_X1 U7944 ( .A1(n8605), .A2(n12713), .ZN(n8604) );
  NAND2_X1 U7945 ( .A1(n12543), .A2(n15766), .ZN(n12556) );
  AOI21_X1 U7946 ( .B1(n12344), .B2(n8534), .A(n8533), .ZN(n8532) );
  INV_X1 U7947 ( .A(n12538), .ZN(n8533) );
  NAND2_X1 U7948 ( .A1(n12345), .A2(n8534), .ZN(n8531) );
  NAND2_X1 U7949 ( .A1(n7673), .A2(n11557), .ZN(n11848) );
  NOR2_X1 U7950 ( .A1(n11751), .A2(n8625), .ZN(n8624) );
  INV_X1 U7951 ( .A(n8627), .ZN(n8625) );
  AND2_X1 U7952 ( .A1(n13580), .A2(n11342), .ZN(n8553) );
  INV_X1 U7953 ( .A(n10704), .ZN(n12760) );
  NAND2_X1 U7954 ( .A1(n9844), .A2(n12814), .ZN(n10702) );
  AND2_X1 U7955 ( .A1(n10389), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9969) );
  OR2_X1 U7956 ( .A1(n16128), .A2(n15739), .ZN(n9968) );
  NAND2_X1 U7957 ( .A1(n8643), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8642) );
  INV_X1 U7958 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n8643) );
  NAND2_X1 U7959 ( .A1(n7662), .A2(n16344), .ZN(n16349) );
  OAI21_X1 U7960 ( .B1(n16342), .B2(n16343), .A(P2_ADDR_REG_10__SCAN_IN), .ZN(
        n7662) );
  NAND2_X1 U7961 ( .A1(n7638), .A2(n7636), .ZN(n16367) );
  NAND2_X1 U7962 ( .A1(P3_ADDR_REG_12__SCAN_IN), .A2(n7637), .ZN(n7636) );
  NAND2_X1 U7963 ( .A1(n16359), .A2(n16358), .ZN(n7638) );
  XNOR2_X1 U7964 ( .A(n16393), .B(P3_ADDR_REG_17__SCAN_IN), .ZN(n16398) );
  NOR2_X1 U7965 ( .A1(n16380), .A2(n16381), .ZN(n16383) );
  AND3_X1 U7966 ( .A1(n7846), .A2(n14056), .A3(P3_REG1_REG_15__SCAN_IN), .ZN(
        n14057) );
  OR2_X1 U7967 ( .A1(n14061), .A2(n14060), .ZN(n8188) );
  AOI21_X1 U7968 ( .B1(n14912), .B2(n13504), .A(n9336), .ZN(n13810) );
  NAND2_X1 U7969 ( .A1(n14957), .A2(n14929), .ZN(n8507) );
  OAI21_X1 U7970 ( .B1(n14977), .B2(n14935), .A(n14978), .ZN(n15010) );
  OAI211_X1 U7971 ( .C1(n7679), .C2(n16726), .A(n7678), .B(n7677), .ZN(n16015)
         );
  INV_X1 U7972 ( .A(n15817), .ZN(n7678) );
  NAND2_X1 U7973 ( .A1(n16017), .A2(n16472), .ZN(n7677) );
  XNOR2_X1 U7974 ( .A(n15813), .B(n8405), .ZN(n7679) );
  INV_X1 U7975 ( .A(n13049), .ZN(n8801) );
  AOI22_X1 U7976 ( .A1(SI_29_), .A2(keyinput_3), .B1(n14910), .B2(keyinput_2), 
        .ZN(n14478) );
  NAND2_X1 U7977 ( .A1(n8482), .A2(n8481), .ZN(n8480) );
  NOR2_X1 U7978 ( .A1(n14487), .A2(n14486), .ZN(n8481) );
  NAND2_X1 U7979 ( .A1(n8476), .A2(n8475), .ZN(n8474) );
  NAND2_X1 U7980 ( .A1(n14490), .A2(SI_20_), .ZN(n8475) );
  NAND2_X1 U7981 ( .A1(n14664), .A2(keyinput_12), .ZN(n8476) );
  AND2_X1 U7982 ( .A1(n8479), .A2(n8478), .ZN(n8477) );
  NAND2_X1 U7983 ( .A1(n14489), .A2(SI_21_), .ZN(n8478) );
  NAND2_X1 U7984 ( .A1(n14662), .A2(keyinput_11), .ZN(n8479) );
  NAND2_X1 U7985 ( .A1(n8207), .A2(n14686), .ZN(n8206) );
  NAND2_X1 U7986 ( .A1(n8210), .A2(n8208), .ZN(n8207) );
  INV_X1 U7987 ( .A(n8209), .ZN(n8208) );
  NOR2_X1 U7988 ( .A1(n14685), .A2(n14684), .ZN(n8205) );
  NAND2_X1 U7989 ( .A1(n13712), .A2(n13714), .ZN(n7962) );
  AOI21_X1 U7990 ( .B1(n14694), .B2(n14695), .A(n8202), .ZN(n8201) );
  XNOR2_X1 U7991 ( .A(keyinput_162), .B(P3_STATE_REG_SCAN_IN), .ZN(n8202) );
  OAI22_X1 U7992 ( .A1(n8861), .A2(n14696), .B1(P3_REG3_REG_7__SCAN_IN), .B2(
        keyinput_163), .ZN(n8200) );
  NAND2_X1 U7993 ( .A1(n7597), .A2(n7455), .ZN(n8466) );
  NAND2_X1 U7994 ( .A1(keyinput_34), .A2(P3_STATE_REG_SCAN_IN), .ZN(n8464) );
  NAND2_X1 U7995 ( .A1(n13080), .A2(n7509), .ZN(n8809) );
  NAND2_X1 U7996 ( .A1(n13729), .A2(n13731), .ZN(n8113) );
  NAND2_X1 U7997 ( .A1(n7949), .A2(n13732), .ZN(n7948) );
  AND2_X1 U7998 ( .A1(n13734), .A2(n7951), .ZN(n7950) );
  INV_X1 U7999 ( .A(n13732), .ZN(n7951) );
  NAND2_X1 U8000 ( .A1(n7751), .A2(n7531), .ZN(n7750) );
  AOI21_X1 U8001 ( .B1(n7753), .B2(n7756), .A(n7557), .ZN(n7752) );
  INV_X1 U8002 ( .A(n13750), .ZN(n7939) );
  AOI21_X1 U8003 ( .B1(n8217), .B2(n8216), .A(n8213), .ZN(n14749) );
  NAND2_X1 U8004 ( .A1(n8215), .A2(n8214), .ZN(n8213) );
  INV_X1 U8005 ( .A(n14721), .ZN(n8216) );
  NAND2_X1 U8006 ( .A1(n8218), .A2(n14722), .ZN(n8217) );
  INV_X1 U8007 ( .A(keyinput_210), .ZN(n8232) );
  AOI21_X1 U8008 ( .B1(n13137), .B2(n13138), .A(n7554), .ZN(n7762) );
  INV_X1 U8009 ( .A(n13131), .ZN(n8806) );
  INV_X1 U8010 ( .A(n13755), .ZN(n7945) );
  NAND2_X1 U8011 ( .A1(n13752), .A2(n13754), .ZN(n8056) );
  OAI21_X1 U8012 ( .B1(n7423), .B2(n7555), .A(n7445), .ZN(n8057) );
  NAND2_X1 U8013 ( .A1(n8062), .A2(n8061), .ZN(n13769) );
  NAND2_X1 U8014 ( .A1(n15777), .A2(n13652), .ZN(n8061) );
  NAND2_X1 U8015 ( .A1(n15882), .A2(n13735), .ZN(n8062) );
  AOI21_X1 U8016 ( .B1(n8230), .B2(n8227), .A(n8224), .ZN(n14772) );
  NAND2_X1 U8017 ( .A1(n13766), .A2(n13765), .ZN(n7958) );
  NOR2_X1 U8018 ( .A1(n8791), .A2(n7511), .ZN(n8790) );
  INV_X1 U8019 ( .A(n13148), .ZN(n8053) );
  OAI21_X1 U8020 ( .B1(n13154), .B2(n8790), .A(n8080), .ZN(n8102) );
  AND2_X1 U8021 ( .A1(n8789), .A2(n8081), .ZN(n8080) );
  INV_X1 U8022 ( .A(n13163), .ZN(n8081) );
  NAND2_X1 U8023 ( .A1(n13780), .A2(n8659), .ZN(n8658) );
  INV_X1 U8024 ( .A(n13652), .ZN(n13612) );
  NAND2_X1 U8025 ( .A1(n12621), .A2(n8667), .ZN(n8666) );
  INV_X1 U8026 ( .A(n12513), .ZN(n8667) );
  AOI21_X1 U8027 ( .B1(n8394), .B2(n8396), .A(n7552), .ZN(n8393) );
  INV_X1 U8028 ( .A(n8856), .ZN(n8394) );
  NAND2_X1 U8029 ( .A1(n8662), .A2(n9999), .ZN(n8007) );
  INV_X1 U8030 ( .A(n10139), .ZN(n8290) );
  OAI21_X1 U8031 ( .B1(n13868), .B2(n13866), .A(n13864), .ZN(n9500) );
  NAND2_X1 U8032 ( .A1(n7851), .A2(n7850), .ZN(n13485) );
  AND2_X1 U8033 ( .A1(n14186), .A2(n8347), .ZN(n7850) );
  AND2_X1 U8034 ( .A1(n13483), .A2(n13491), .ZN(n8076) );
  NOR2_X1 U8035 ( .A1(n14262), .A2(n7543), .ZN(n8151) );
  INV_X1 U8036 ( .A(n9259), .ZN(n8152) );
  NAND2_X1 U8037 ( .A1(n13011), .A2(n13342), .ZN(n13302) );
  INV_X1 U8038 ( .A(n16059), .ZN(n7724) );
  NAND2_X1 U8039 ( .A1(n13247), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n8109) );
  NAND2_X1 U8040 ( .A1(n9874), .A2(n10464), .ZN(n8118) );
  OAI21_X1 U8041 ( .B1(n16283), .B2(P1_ADDR_REG_2__SCAN_IN), .A(n7476), .ZN(
        n7641) );
  NAND2_X1 U8042 ( .A1(n9500), .A2(n9499), .ZN(n9503) );
  NAND2_X1 U8043 ( .A1(n9501), .A2(n9503), .ZN(n13943) );
  OR2_X1 U8044 ( .A1(n9500), .A2(n9499), .ZN(n9501) );
  INV_X1 U8045 ( .A(n8191), .ZN(n9658) );
  OR2_X1 U8046 ( .A1(n9677), .A2(n11524), .ZN(n8420) );
  NAND2_X1 U8047 ( .A1(n9630), .A2(n7605), .ZN(n8187) );
  INV_X1 U8048 ( .A(n11613), .ZN(n8183) );
  INV_X1 U8049 ( .A(n8187), .ZN(n8180) );
  OR2_X1 U8050 ( .A1(n11605), .A2(n9680), .ZN(n9682) );
  AOI21_X1 U8051 ( .B1(n8178), .B2(n8197), .A(n9661), .ZN(n8195) );
  NAND2_X1 U8052 ( .A1(n16425), .A2(n8197), .ZN(n8196) );
  NAND2_X1 U8053 ( .A1(n7690), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n8414) );
  INV_X1 U8054 ( .A(n12161), .ZN(n7690) );
  NAND2_X1 U8055 ( .A1(n9685), .A2(n9684), .ZN(n8415) );
  NAND2_X1 U8056 ( .A1(n7478), .A2(n8429), .ZN(n14039) );
  NAND2_X1 U8057 ( .A1(n8431), .A2(n8430), .ZN(n8429) );
  NOR2_X1 U8058 ( .A1(n8433), .A2(n14017), .ZN(n8430) );
  NOR2_X1 U8059 ( .A1(n14039), .A2(n7699), .ZN(n14040) );
  AND2_X1 U8060 ( .A1(n14046), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n7699) );
  OR2_X1 U8061 ( .A1(n9384), .A2(n14198), .ZN(n13474) );
  NOR2_X1 U8062 ( .A1(n8165), .A2(n8157), .ZN(n8156) );
  INV_X1 U8063 ( .A(n9124), .ZN(n8157) );
  AOI21_X1 U8064 ( .B1(n8161), .B2(n8164), .A(n8160), .ZN(n8159) );
  INV_X1 U8065 ( .A(n8162), .ZN(n8161) );
  NOR2_X1 U8066 ( .A1(n13537), .A2(n8163), .ZN(n8162) );
  INV_X1 U8067 ( .A(n9139), .ZN(n8163) );
  INV_X1 U8068 ( .A(n13379), .ZN(n8338) );
  NOR2_X1 U8069 ( .A1(n8339), .A2(n8336), .ZN(n8335) );
  OR2_X1 U8070 ( .A1(n9448), .A2(n14184), .ZN(n13478) );
  AND2_X1 U8071 ( .A1(n8747), .A2(n8374), .ZN(n8373) );
  NOR2_X1 U8072 ( .A1(P3_IR_REG_28__SCAN_IN), .A2(n8885), .ZN(n8374) );
  NOR2_X1 U8073 ( .A1(P3_IR_REG_22__SCAN_IN), .A2(P3_IR_REG_23__SCAN_IN), .ZN(
        n8741) );
  NAND2_X1 U8074 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(n8582), .ZN(n8581) );
  INV_X1 U8075 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n9423) );
  AND2_X1 U8076 ( .A1(n8945), .A2(n8746), .ZN(n9344) );
  INV_X1 U8077 ( .A(n8748), .ZN(n8746) );
  NOR2_X1 U8078 ( .A1(n9346), .A2(P3_IR_REG_21__SCAN_IN), .ZN(n9389) );
  NAND2_X1 U8079 ( .A1(n8910), .A2(n8077), .ZN(n8911) );
  NAND2_X1 U8080 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n8078), .ZN(n8077) );
  INV_X1 U8081 ( .A(n8909), .ZN(n8571) );
  NAND2_X1 U8082 ( .A1(n7833), .A2(n8908), .ZN(n7832) );
  NAND2_X1 U8083 ( .A1(n7489), .A2(n7834), .ZN(n7830) );
  INV_X1 U8084 ( .A(n8908), .ZN(n7834) );
  INV_X1 U8085 ( .A(n8903), .ZN(n7840) );
  INV_X1 U8086 ( .A(n7839), .ZN(n7838) );
  OAI21_X1 U8087 ( .B1(n9012), .B2(n7840), .A(n9029), .ZN(n7839) );
  NOR2_X1 U8088 ( .A1(P3_IR_REG_4__SCAN_IN), .A2(P3_IR_REG_3__SCAN_IN), .ZN(
        n8876) );
  INV_X1 U8089 ( .A(n11360), .ZN(n8279) );
  INV_X1 U8090 ( .A(n7471), .ZN(n8273) );
  NAND2_X1 U8091 ( .A1(n8688), .A2(n8686), .ZN(n8685) );
  CLKBUF_X1 U8092 ( .A(n13302), .Z(n8104) );
  NAND2_X1 U8093 ( .A1(n7410), .A2(n15160), .ZN(n8697) );
  INV_X1 U8094 ( .A(n15158), .ZN(n7875) );
  NAND2_X1 U8095 ( .A1(n12584), .A2(n8711), .ZN(n8710) );
  NAND2_X1 U8096 ( .A1(n13328), .A2(n12492), .ZN(n8711) );
  AOI21_X1 U8097 ( .B1(n8704), .B2(n8702), .A(n7537), .ZN(n8701) );
  INV_X1 U8098 ( .A(n12135), .ZN(n8702) );
  NAND2_X1 U8099 ( .A1(n11764), .A2(n7880), .ZN(n7879) );
  NOR2_X1 U8100 ( .A1(n8703), .A2(n7881), .ZN(n7880) );
  INV_X1 U8101 ( .A(n11763), .ZN(n7881) );
  INV_X1 U8102 ( .A(n8704), .ZN(n8703) );
  NAND2_X1 U8103 ( .A1(n11764), .A2(n11763), .ZN(n11765) );
  AND2_X1 U8104 ( .A1(n8764), .A2(n8762), .ZN(n11264) );
  INV_X1 U8105 ( .A(n8765), .ZN(n8762) );
  OR2_X1 U8106 ( .A1(n7981), .A2(n7980), .ZN(n7979) );
  INV_X1 U8107 ( .A(n8776), .ZN(n7980) );
  NAND2_X1 U8108 ( .A1(n9715), .A2(P2_IR_REG_28__SCAN_IN), .ZN(n7857) );
  NAND2_X1 U8109 ( .A1(n7977), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7859) );
  NOR2_X1 U8110 ( .A1(n10990), .A2(n7545), .ZN(n9721) );
  AND2_X1 U8111 ( .A1(n7446), .A2(n16529), .ZN(n7422) );
  OR2_X1 U8112 ( .A1(n13719), .A2(n13715), .ZN(n7729) );
  NAND2_X1 U8113 ( .A1(n15689), .A2(n13677), .ZN(n8544) );
  NAND2_X1 U8114 ( .A1(n15955), .A2(n8547), .ZN(n8549) );
  AND2_X1 U8115 ( .A1(n13217), .A2(n12645), .ZN(n13215) );
  NAND2_X1 U8116 ( .A1(n12915), .A2(n12635), .ZN(n12638) );
  INV_X1 U8117 ( .A(n12875), .ZN(n8023) );
  NAND2_X1 U8118 ( .A1(n12627), .A2(SI_24_), .ZN(n12628) );
  NAND2_X1 U8119 ( .A1(n7993), .A2(n7457), .ZN(n8844) );
  NAND2_X1 U8120 ( .A1(n11883), .A2(n14666), .ZN(n12150) );
  XNOR2_X1 U8121 ( .A(n8063), .B(n14492), .ZN(n11881) );
  NAND2_X1 U8122 ( .A1(n11161), .A2(n7454), .ZN(n8380) );
  INV_X1 U8123 ( .A(n11161), .ZN(n8383) );
  INV_X1 U8124 ( .A(n10619), .ZN(n8660) );
  NAND2_X1 U8125 ( .A1(n10140), .A2(n10139), .ZN(n10214) );
  NAND2_X1 U8126 ( .A1(n8664), .A2(n8662), .ZN(n10140) );
  INV_X1 U8127 ( .A(n9973), .ZN(n8399) );
  XNOR2_X1 U8128 ( .A(n16284), .B(n8009), .ZN(n16285) );
  OAI21_X1 U8129 ( .B1(n16313), .B2(n16314), .A(n16312), .ZN(n16315) );
  NAND2_X1 U8130 ( .A1(n7643), .A2(n16330), .ZN(n16335) );
  NAND2_X1 U8131 ( .A1(n16328), .A2(n16329), .ZN(n7643) );
  AND2_X1 U8132 ( .A1(n7640), .A2(n7639), .ZN(n16359) );
  NAND2_X1 U8133 ( .A1(n16354), .A2(P1_ADDR_REG_11__SCAN_IN), .ZN(n7639) );
  OR2_X1 U8134 ( .A1(n16352), .A2(n16353), .ZN(n7640) );
  OAI21_X1 U8135 ( .B1(P3_ADDR_REG_15__SCAN_IN), .B2(n16379), .A(n7645), .ZN(
        n16385) );
  NAND2_X1 U8136 ( .A1(n16378), .A2(n16377), .ZN(n7645) );
  INV_X1 U8137 ( .A(n9468), .ZN(n7895) );
  NAND2_X1 U8138 ( .A1(n7894), .A2(n7895), .ZN(n7893) );
  INV_X1 U8139 ( .A(n13932), .ZN(n7894) );
  OR2_X1 U8140 ( .A1(n9454), .A2(n9455), .ZN(n8733) );
  INV_X1 U8141 ( .A(n8732), .ZN(n8728) );
  NOR2_X1 U8142 ( .A1(n12299), .A2(n7885), .ZN(n7884) );
  INV_X1 U8143 ( .A(n7886), .ZN(n7885) );
  AND3_X1 U8144 ( .A1(n8988), .A2(n8987), .A3(n8986), .ZN(n9449) );
  NAND2_X1 U8145 ( .A1(n11661), .A2(n11660), .ZN(n8724) );
  OR2_X1 U8146 ( .A1(n7893), .A2(n7891), .ZN(n7890) );
  INV_X1 U8147 ( .A(n13835), .ZN(n7891) );
  AND2_X1 U8148 ( .A1(n7888), .A2(n7890), .ZN(n13974) );
  NAND2_X1 U8149 ( .A1(n8359), .A2(n8358), .ZN(n8357) );
  INV_X1 U8150 ( .A(n13512), .ZN(n8360) );
  NAND2_X1 U8151 ( .A1(n13513), .A2(n13514), .ZN(n8361) );
  AND3_X1 U8152 ( .A1(n8358), .A2(n13520), .A3(n7576), .ZN(n13548) );
  AND2_X1 U8153 ( .A1(n14163), .A2(n8576), .ZN(n8575) );
  OAI211_X1 U8154 ( .C1(n13490), .C2(n7845), .A(n7844), .B(n8578), .ZN(n13508)
         );
  NAND2_X1 U8155 ( .A1(n13511), .A2(n13480), .ZN(n7845) );
  OAI21_X1 U8156 ( .B1(n13490), .B2(n13509), .A(n13491), .ZN(n7844) );
  NAND2_X1 U8157 ( .A1(n9422), .A2(n9421), .ZN(n9589) );
  NOR2_X1 U8158 ( .A1(n13831), .A2(n12294), .ZN(n9421) );
  OR2_X1 U8160 ( .A1(n10995), .A2(n9597), .ZN(n8969) );
  OR2_X1 U8161 ( .A1(n10919), .A2(n7819), .ZN(n7818) );
  AND2_X1 U8162 ( .A1(n9655), .A2(n9675), .ZN(n7819) );
  NAND2_X1 U8163 ( .A1(n8191), .A2(n8190), .ZN(n11516) );
  NOR2_X1 U8164 ( .A1(n11516), .A2(n9620), .ZN(n11515) );
  NAND2_X1 U8165 ( .A1(n8420), .A2(n8419), .ZN(n11518) );
  NAND2_X1 U8166 ( .A1(n9677), .A2(n11524), .ZN(n8419) );
  NAND2_X1 U8167 ( .A1(n11511), .A2(n9623), .ZN(n11608) );
  NAND2_X1 U8168 ( .A1(n7689), .A2(n9630), .ZN(n8417) );
  INV_X1 U8169 ( .A(n9682), .ZN(n7689) );
  NAND2_X1 U8170 ( .A1(n7688), .A2(n7687), .ZN(n11956) );
  INV_X1 U8171 ( .A(n11959), .ZN(n7687) );
  INV_X1 U8172 ( .A(n11958), .ZN(n7688) );
  NOR2_X1 U8173 ( .A1(n16426), .A2(n9628), .ZN(n16425) );
  NAND2_X1 U8174 ( .A1(n7811), .A2(n7809), .ZN(n13992) );
  NAND2_X1 U8175 ( .A1(n9664), .A2(n7814), .ZN(n7811) );
  NAND2_X1 U8176 ( .A1(n7812), .A2(n7810), .ZN(n7809) );
  NOR2_X1 U8177 ( .A1(n9640), .A2(n7736), .ZN(n7735) );
  INV_X1 U8178 ( .A(n7738), .ZN(n7736) );
  OR2_X1 U8179 ( .A1(n14014), .A2(n8433), .ZN(n8432) );
  NOR2_X1 U8180 ( .A1(n13994), .A2(n9155), .ZN(n14009) );
  NAND2_X1 U8181 ( .A1(n7843), .A2(n7842), .ZN(n8177) );
  INV_X1 U8182 ( .A(n14011), .ZN(n7842) );
  NAND2_X1 U8183 ( .A1(n14040), .A2(n14063), .ZN(n8436) );
  OR2_X1 U8184 ( .A1(n14040), .A2(n14063), .ZN(n8437) );
  OR2_X1 U8185 ( .A1(n14094), .A2(n14095), .ZN(n14111) );
  INV_X1 U8186 ( .A(n8423), .ZN(n14118) );
  NOR2_X1 U8187 ( .A1(n14118), .A2(n8424), .ZN(n14119) );
  XNOR2_X1 U8188 ( .A(n14138), .B(n7757), .ZN(n14115) );
  INV_X1 U8189 ( .A(n14137), .ZN(n7757) );
  OAI21_X1 U8190 ( .B1(n14105), .B2(n14104), .A(n14103), .ZN(n14129) );
  NAND2_X1 U8191 ( .A1(n14115), .A2(n14114), .ZN(n14136) );
  XNOR2_X1 U8192 ( .A(n7914), .B(n14186), .ZN(n7913) );
  NAND2_X1 U8193 ( .A1(n14192), .A2(n8142), .ZN(n7914) );
  NOR2_X1 U8194 ( .A1(n14184), .A2(n14314), .ZN(n7911) );
  AOI21_X1 U8195 ( .B1(n8347), .B2(n13484), .A(n7559), .ZN(n8346) );
  AND2_X1 U8196 ( .A1(n13474), .A2(n13473), .ZN(n14186) );
  NOR2_X1 U8197 ( .A1(n14193), .A2(n8349), .ZN(n8348) );
  OAI22_X1 U8198 ( .A1(n14222), .A2(n14216), .B1(n13847), .B2(n14208), .ZN(
        n14210) );
  NAND2_X1 U8199 ( .A1(n7896), .A2(n7897), .ZN(n14217) );
  NAND2_X1 U8200 ( .A1(n7563), .A2(n7900), .ZN(n7897) );
  OR3_X1 U8201 ( .A1(n14296), .A2(n13459), .A3(n8145), .ZN(n7896) );
  AOI21_X1 U8202 ( .B1(n14327), .B2(n14326), .A(n9224), .ZN(n14308) );
  NAND2_X1 U8203 ( .A1(n8356), .A2(n13427), .ZN(n14315) );
  OR2_X1 U8204 ( .A1(n14367), .A2(n9366), .ZN(n8356) );
  AOI21_X1 U8205 ( .B1(n12392), .B2(n8162), .A(n8165), .ZN(n8158) );
  NOR2_X1 U8207 ( .A1(n8370), .A2(n12282), .ZN(n8369) );
  INV_X1 U8208 ( .A(n13403), .ZN(n8370) );
  NAND2_X1 U8209 ( .A1(n9361), .A2(n13392), .ZN(n12234) );
  NAND2_X1 U8210 ( .A1(n9360), .A2(n13374), .ZN(n11920) );
  OR2_X1 U8211 ( .A1(n16493), .A2(n16499), .ZN(n16491) );
  AND4_X1 U8212 ( .A1(n9011), .A2(n9010), .A3(n9009), .A4(n9008), .ZN(n11925)
         );
  INV_X1 U8213 ( .A(n16498), .ZN(n14312) );
  NAND2_X1 U8214 ( .A1(n7434), .A2(n7495), .ZN(n8139) );
  AND2_X1 U8215 ( .A1(n9535), .A2(n13480), .ZN(n16495) );
  OAI21_X1 U8216 ( .B1(n8447), .B2(n8446), .A(n8452), .ZN(n8445) );
  NAND2_X1 U8217 ( .A1(n13496), .A2(n13495), .ZN(n13510) );
  NAND2_X1 U8218 ( .A1(n10787), .A2(n14147), .ZN(n13550) );
  AND2_X1 U8219 ( .A1(n9589), .A2(n14899), .ZN(n11012) );
  INV_X1 U8220 ( .A(n16497), .ZN(n11333) );
  INV_X1 U8221 ( .A(n16495), .ZN(n14314) );
  INV_X1 U8222 ( .A(n8590), .ZN(n8589) );
  OAI21_X1 U8223 ( .B1(n13492), .B2(n8592), .A(n8591), .ZN(n8590) );
  NAND2_X1 U8224 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n13600), .ZN(n8591) );
  NAND2_X1 U8225 ( .A1(n8171), .A2(n7505), .ZN(n9395) );
  NAND2_X1 U8226 ( .A1(n7828), .A2(n7826), .ZN(n9293) );
  NAND2_X1 U8227 ( .A1(P2_DATAO_REG_22__SCAN_IN), .A2(n7827), .ZN(n7826) );
  NAND2_X1 U8228 ( .A1(n9282), .A2(n9281), .ZN(n7828) );
  AOI21_X1 U8229 ( .B1(n9261), .B2(n9260), .A(n8574), .ZN(n8573) );
  NOR2_X1 U8230 ( .A1(n12779), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8574) );
  NAND2_X1 U8231 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n8120), .ZN(n8119) );
  AOI21_X1 U8232 ( .B1(n7823), .B2(n7825), .A(n7610), .ZN(n7821) );
  XNOR2_X1 U8233 ( .A(n8911), .B(P2_DATAO_REG_13__SCAN_IN), .ZN(n9164) );
  AND2_X1 U8234 ( .A1(n9170), .A2(n9190), .ZN(n14024) );
  NAND2_X1 U8235 ( .A1(n7831), .A2(n8908), .ZN(n9120) );
  NAND2_X1 U8236 ( .A1(n9076), .A2(n9075), .ZN(n7831) );
  XNOR2_X1 U8237 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .ZN(n9118) );
  OAI22_X1 U8238 ( .A1(n9067), .A2(n9065), .B1(P2_DATAO_REG_7__SCAN_IN), .B2(
        n9928), .ZN(n9096) );
  XNOR2_X1 U8239 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .ZN(n9095) );
  XNOR2_X1 U8240 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .ZN(n9029) );
  OAI21_X1 U8241 ( .B1(n8997), .B2(n8901), .A(n8902), .ZN(n9014) );
  XNOR2_X1 U8242 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .ZN(n9012) );
  INV_X1 U8243 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n8413) );
  NAND2_X1 U8244 ( .A1(n7930), .A2(n11135), .ZN(n10647) );
  NOR2_X1 U8245 ( .A1(n9822), .A2(n7931), .ZN(n7930) );
  INV_X1 U8246 ( .A(n9769), .ZN(n7931) );
  NOR2_X1 U8247 ( .A1(n7483), .A2(n8286), .ZN(n8285) );
  INV_X1 U8248 ( .A(n11061), .ZN(n8286) );
  NOR2_X1 U8249 ( .A1(n14999), .A2(n12974), .ZN(n8295) );
  NAND2_X1 U8250 ( .A1(n14923), .A2(n8273), .ZN(n8270) );
  NAND2_X1 U8251 ( .A1(n14968), .A2(n8272), .ZN(n8271) );
  NOR2_X1 U8252 ( .A1(n14923), .A2(n8273), .ZN(n8272) );
  NAND2_X1 U8253 ( .A1(n7918), .A2(n11102), .ZN(n11361) );
  NAND2_X1 U8254 ( .A1(n11101), .A2(n11090), .ZN(n7918) );
  NAND2_X1 U8255 ( .A1(n8291), .A2(n7472), .ZN(n8498) );
  NAND2_X1 U8256 ( .A1(n8502), .A2(n11047), .ZN(n8291) );
  AND2_X1 U8257 ( .A1(n7929), .A2(n7928), .ZN(n7927) );
  AND2_X1 U8258 ( .A1(n15025), .A2(n14938), .ZN(n7929) );
  NAND2_X1 U8259 ( .A1(n14978), .A2(n14935), .ZN(n7928) );
  NOR2_X1 U8260 ( .A1(n8316), .A2(n15110), .ZN(n8315) );
  NAND2_X1 U8261 ( .A1(n7975), .A2(n7973), .ZN(n15131) );
  NOR2_X1 U8262 ( .A1(n15129), .A2(n7974), .ZN(n7973) );
  INV_X1 U8263 ( .A(n15128), .ZN(n7974) );
  NAND2_X1 U8264 ( .A1(n7876), .A2(n15158), .ZN(n15236) );
  NAND2_X1 U8265 ( .A1(n8690), .A2(n7877), .ZN(n7876) );
  NAND2_X1 U8266 ( .A1(n15270), .A2(n15269), .ZN(n7975) );
  NOR2_X1 U8267 ( .A1(n15284), .A2(n7871), .ZN(n7870) );
  INV_X1 U8268 ( .A(n15152), .ZN(n7871) );
  NAND2_X1 U8269 ( .A1(n15305), .A2(n15306), .ZN(n7872) );
  NAND2_X1 U8270 ( .A1(n12499), .A2(n8757), .ZN(n8754) );
  OAI21_X1 U8271 ( .B1(n12499), .B2(n8753), .A(n8751), .ZN(n15347) );
  NAND2_X1 U8272 ( .A1(n8759), .A2(n13329), .ZN(n12588) );
  INV_X1 U8273 ( .A(n12499), .ZN(n8759) );
  NAND2_X1 U8274 ( .A1(n8713), .A2(n8712), .ZN(n12493) );
  AND2_X1 U8275 ( .A1(n13327), .A2(n12223), .ZN(n8779) );
  NAND2_X1 U8276 ( .A1(n7602), .A2(n13325), .ZN(n12224) );
  NAND2_X1 U8277 ( .A1(n11719), .A2(n8773), .ZN(n11760) );
  NOR2_X1 U8278 ( .A1(n11722), .A2(n8774), .ZN(n8773) );
  INV_X1 U8279 ( .A(n11718), .ZN(n8774) );
  NAND2_X1 U8280 ( .A1(n11590), .A2(n13320), .ZN(n11592) );
  NAND2_X1 U8281 ( .A1(n11592), .A2(n8775), .ZN(n11719) );
  AND2_X1 U8282 ( .A1(n13321), .A2(n11591), .ZN(n8775) );
  AND2_X1 U8283 ( .A1(n10077), .A2(n10089), .ZN(n15343) );
  NAND2_X1 U8284 ( .A1(n11383), .A2(n8771), .ZN(n11638) );
  NOR2_X1 U8285 ( .A1(n13317), .A2(n8772), .ZN(n8771) );
  INV_X1 U8286 ( .A(n11382), .ZN(n8772) );
  OR2_X1 U8287 ( .A1(n11264), .A2(n7669), .ZN(n11238) );
  NOR2_X1 U8288 ( .A1(n8765), .A2(n16586), .ZN(n8763) );
  NAND3_X1 U8289 ( .A1(n11239), .A2(n11238), .A3(n13319), .ZN(n11383) );
  NAND2_X1 U8290 ( .A1(n10520), .A2(n13312), .ZN(n10519) );
  NAND2_X1 U8291 ( .A1(n13345), .A2(n9824), .ZN(n11246) );
  OR2_X1 U8292 ( .A1(n9893), .A2(n10463), .ZN(n9741) );
  NAND2_X1 U8293 ( .A1(n12728), .A2(n12053), .ZN(n8015) );
  NAND2_X1 U8294 ( .A1(n12056), .A2(n12055), .ZN(n13113) );
  INV_X1 U8295 ( .A(n13011), .ZN(n16590) );
  AND2_X1 U8296 ( .A1(n9817), .A2(n9816), .ZN(n11242) );
  INV_X1 U8297 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n9699) );
  NAND2_X1 U8298 ( .A1(n9582), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9585) );
  XNOR2_X1 U8299 ( .A(n9587), .B(n9698), .ZN(n13350) );
  OAI21_X1 U8300 ( .B1(n11327), .B2(n9725), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n9731) );
  INV_X1 U8301 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n9726) );
  INV_X1 U8302 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n9722) );
  INV_X1 U8303 ( .A(n8832), .ZN(n8831) );
  OAI22_X1 U8304 ( .A1(n12526), .A2(n8836), .B1(n12524), .B2(n12525), .ZN(
        n8832) );
  NAND2_X1 U8305 ( .A1(n12377), .A2(n7802), .ZN(n7801) );
  INV_X1 U8306 ( .A(n8834), .ZN(n8833) );
  NAND2_X1 U8307 ( .A1(n8066), .A2(n8065), .ZN(n8064) );
  NAND2_X1 U8308 ( .A1(n11022), .A2(n7532), .ZN(n7779) );
  NOR2_X1 U8309 ( .A1(n11690), .A2(n8824), .ZN(n8823) );
  INV_X1 U8310 ( .A(n11021), .ZN(n8824) );
  INV_X1 U8311 ( .A(n8822), .ZN(n8821) );
  OAI21_X1 U8312 ( .B1(n11690), .B2(n8828), .A(n8827), .ZN(n8822) );
  INV_X1 U8313 ( .A(n10730), .ZN(n7772) );
  NAND2_X1 U8314 ( .A1(n10694), .A2(n7777), .ZN(n7774) );
  NAND2_X1 U8315 ( .A1(n7776), .A2(n7422), .ZN(n7775) );
  NAND3_X1 U8316 ( .A1(n7422), .A2(n7776), .A3(n7777), .ZN(n7773) );
  OR2_X1 U8317 ( .A1(n8818), .A2(n8817), .ZN(n8816) );
  INV_X1 U8318 ( .A(n8826), .ZN(n8817) );
  NAND2_X1 U8319 ( .A1(n10354), .A2(n7767), .ZN(n10353) );
  OR2_X1 U8320 ( .A1(n15646), .A2(n7790), .ZN(n7789) );
  OR2_X1 U8321 ( .A1(n15576), .A2(n15577), .ZN(n15574) );
  NAND2_X1 U8322 ( .A1(n15560), .A2(n12853), .ZN(n7795) );
  INV_X1 U8323 ( .A(n13800), .ZN(n8073) );
  NOR3_X2 U8324 ( .A1(n15848), .A2(n15786), .A3(n8305), .ZN(n15785) );
  NOR2_X1 U8325 ( .A1(n15848), .A2(n8304), .ZN(n15818) );
  INV_X1 U8326 ( .A(n8306), .ZN(n8304) );
  NAND2_X1 U8327 ( .A1(n15838), .A2(n16462), .ZN(n8097) );
  NOR2_X1 U8328 ( .A1(n15843), .A2(n7996), .ZN(n7994) );
  INV_X1 U8329 ( .A(n8538), .ZN(n7996) );
  NAND2_X1 U8330 ( .A1(n7487), .A2(n8632), .ZN(n8631) );
  NAND2_X1 U8331 ( .A1(n7705), .A2(n7704), .ZN(n8630) );
  OR2_X1 U8332 ( .A1(n15774), .A2(n15760), .ZN(n8607) );
  AND4_X1 U8333 ( .A1(n12822), .A2(n12821), .A3(n12820), .A4(n12819), .ZN(
        n15761) );
  NAND2_X1 U8334 ( .A1(n7479), .A2(n8546), .ZN(n8021) );
  NAND2_X1 U8335 ( .A1(n15956), .A2(n7479), .ZN(n7681) );
  AOI21_X1 U8336 ( .B1(n15934), .B2(n15933), .A(n7551), .ZN(n15916) );
  OR2_X1 U8337 ( .A1(n15757), .A2(n15758), .ZN(n8611) );
  INV_X1 U8338 ( .A(n15916), .ZN(n15757) );
  INV_X1 U8339 ( .A(n15956), .ZN(n15955) );
  NAND2_X1 U8340 ( .A1(n7718), .A2(n7717), .ZN(n15948) );
  NAND2_X1 U8341 ( .A1(n8310), .A2(n8309), .ZN(n15975) );
  NAND2_X1 U8342 ( .A1(n8599), .A2(n7601), .ZN(n15753) );
  NAND2_X1 U8343 ( .A1(n12555), .A2(n8604), .ZN(n8599) );
  NAND2_X1 U8344 ( .A1(n12554), .A2(n8604), .ZN(n8598) );
  INV_X1 U8345 ( .A(n12345), .ZN(n8537) );
  INV_X1 U8346 ( .A(n12343), .ZN(n8535) );
  AOI21_X1 U8347 ( .B1(n7712), .B2(n7713), .A(n7536), .ZN(n7711) );
  OR2_X1 U8348 ( .A1(n11869), .A2(n7714), .ZN(n7710) );
  NAND2_X1 U8349 ( .A1(n12021), .A2(n12020), .ZN(n12324) );
  NAND2_X1 U8350 ( .A1(n8621), .A2(n8619), .ZN(n11906) );
  NOR2_X1 U8351 ( .A1(n8622), .A2(n8620), .ZN(n8619) );
  NOR2_X1 U8352 ( .A1(n8552), .A2(n13582), .ZN(n8550) );
  INV_X1 U8353 ( .A(n7675), .ZN(n7674) );
  OAI21_X1 U8354 ( .B1(n10704), .B2(n9878), .A(n7676), .ZN(n7675) );
  OAI21_X1 U8355 ( .B1(n10932), .B2(n7703), .A(n10947), .ZN(n7702) );
  NOR2_X1 U8356 ( .A1(n10933), .A2(n7703), .ZN(n7700) );
  OR2_X1 U8357 ( .A1(n16464), .A2(n15733), .ZN(n10876) );
  INV_X1 U8358 ( .A(n15690), .ZN(n13655) );
  NAND2_X1 U8359 ( .A1(n10876), .A2(n10879), .ZN(n16606) );
  OAI21_X1 U8360 ( .B1(n10381), .B2(P1_D_REG_0__SCAN_IN), .A(n16114), .ZN(
        n11137) );
  INV_X1 U8361 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n9990) );
  NAND2_X1 U8362 ( .A1(n9569), .A2(n8845), .ZN(n9561) );
  AND2_X1 U8363 ( .A1(n7593), .A2(P1_IR_REG_22__SCAN_IN), .ZN(n8641) );
  OAI21_X1 U8364 ( .B1(n7593), .B2(n8642), .A(n8640), .ZN(n8639) );
  NAND2_X1 U8365 ( .A1(n10054), .A2(P1_IR_REG_22__SCAN_IN), .ZN(n8640) );
  INV_X1 U8366 ( .A(n9551), .ZN(n7803) );
  INV_X1 U8367 ( .A(n9550), .ZN(n7806) );
  NOR2_X1 U8368 ( .A1(n9929), .A2(n7805), .ZN(n7804) );
  NOR2_X1 U8369 ( .A1(n16278), .A2(P2_ADDR_REG_2__SCAN_IN), .ZN(n16279) );
  NOR2_X1 U8370 ( .A1(n16294), .A2(n16293), .ZN(n16308) );
  NOR2_X1 U8371 ( .A1(n7648), .A2(P1_ADDR_REG_4__SCAN_IN), .ZN(n16293) );
  AOI21_X1 U8372 ( .B1(n16414), .B2(n16310), .A(n16411), .ZN(n16321) );
  INV_X1 U8373 ( .A(n7663), .ZN(n16338) );
  OAI21_X1 U8374 ( .B1(n16351), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n7498), .ZN(
        n8518) );
  AOI22_X1 U8375 ( .A1(P3_ADDR_REG_13__SCAN_IN), .A2(n16368), .B1(n16367), 
        .B2(n16366), .ZN(n16374) );
  NAND2_X1 U8376 ( .A1(n7649), .A2(n16401), .ZN(n7656) );
  AOI21_X1 U8377 ( .B1(n16382), .B2(n8512), .A(n7651), .ZN(n7650) );
  OR2_X1 U8378 ( .A1(n11661), .A2(n8722), .ZN(n8720) );
  AOI21_X1 U8379 ( .B1(n13975), .B2(n9492), .A(n8851), .ZN(n13925) );
  INV_X1 U8380 ( .A(n9449), .ZN(n16494) );
  AND4_X1 U8381 ( .A1(n9028), .A2(n9027), .A3(n9026), .A4(n9025), .ZN(n11829)
         );
  NAND2_X1 U8382 ( .A1(n9397), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7764) );
  NAND2_X1 U8383 ( .A1(n7562), .A2(n7442), .ZN(n10517) );
  OR2_X1 U8384 ( .A1(n14009), .A2(n14010), .ZN(n7843) );
  INV_X1 U8385 ( .A(n8177), .ZN(n14036) );
  NOR2_X1 U8386 ( .A1(n14057), .A2(n14058), .ZN(n14061) );
  NOR2_X1 U8387 ( .A1(n14081), .A2(n14439), .ZN(n14105) );
  OAI21_X1 U8388 ( .B1(n16438), .B2(n16404), .A(n14123), .ZN(n7696) );
  INV_X1 U8389 ( .A(n8443), .ZN(n8442) );
  AOI21_X1 U8390 ( .B1(n14146), .B2(n14147), .A(n8444), .ZN(n8443) );
  NAND2_X1 U8391 ( .A1(n14134), .A2(n14135), .ZN(n8444) );
  XNOR2_X1 U8392 ( .A(n14133), .B(n8440), .ZN(n8439) );
  INV_X1 U8393 ( .A(n14141), .ZN(n8440) );
  OR2_X1 U8394 ( .A1(n11212), .A2(n13555), .ZN(n16429) );
  NAND2_X1 U8395 ( .A1(n8125), .A2(n7503), .ZN(n8126) );
  INV_X1 U8396 ( .A(n14160), .ZN(n8125) );
  NAND2_X1 U8397 ( .A1(n8132), .A2(n13547), .ZN(n8131) );
  NAND2_X1 U8398 ( .A1(n14160), .A2(n8129), .ZN(n8128) );
  NOR2_X1 U8399 ( .A1(n8130), .A2(n14310), .ZN(n8129) );
  AND2_X1 U8400 ( .A1(n7583), .A2(n8132), .ZN(n8130) );
  OR2_X1 U8401 ( .A1(n11014), .A2(n11013), .ZN(n14384) );
  AND2_X1 U8402 ( .A1(n14352), .A2(n11814), .ZN(n14372) );
  AND3_X1 U8403 ( .A1(n9038), .A2(n9037), .A3(n9036), .ZN(n11931) );
  NAND2_X1 U8404 ( .A1(n9181), .A2(n9180), .ZN(n14895) );
  XNOR2_X1 U8405 ( .A(n8043), .B(n13492), .ZN(n14912) );
  NAND2_X1 U8406 ( .A1(n8945), .A2(n8371), .ZN(n8045) );
  NAND2_X1 U8407 ( .A1(n9244), .A2(n9247), .ZN(n14132) );
  NAND2_X1 U8408 ( .A1(n14945), .A2(n14944), .ZN(n8101) );
  NAND2_X1 U8409 ( .A1(n12059), .A2(n12058), .ZN(n16741) );
  NAND2_X1 U8410 ( .A1(n8263), .A2(n8262), .ZN(n8261) );
  NAND2_X1 U8411 ( .A1(n15184), .A2(n8849), .ZN(n8262) );
  NAND2_X1 U8412 ( .A1(n15165), .A2(n14961), .ZN(n8263) );
  NOR2_X1 U8413 ( .A1(n8506), .A2(n8264), .ZN(n8256) );
  INV_X1 U8414 ( .A(n8265), .ZN(n8264) );
  OAI21_X1 U8415 ( .B1(n15165), .B2(n15011), .A(n8266), .ZN(n8265) );
  OAI21_X1 U8416 ( .B1(n11101), .B2(n7920), .A(n7915), .ZN(n7917) );
  NAND2_X1 U8417 ( .A1(n10469), .A2(n10468), .ZN(n13054) );
  NAND2_X1 U8418 ( .A1(n14927), .A2(n14926), .ZN(n14928) );
  NAND2_X1 U8419 ( .A1(n7923), .A2(n7927), .ZN(n15022) );
  NAND2_X1 U8420 ( .A1(n14977), .A2(n14978), .ZN(n7923) );
  NAND2_X1 U8421 ( .A1(n9830), .A2(n15364), .ZN(n15024) );
  CLKBUF_X1 U8422 ( .A(n15014), .Z(n15000) );
  XNOR2_X1 U8423 ( .A(n8071), .B(n13338), .ZN(n13336) );
  NAND2_X1 U8424 ( .A1(n13345), .A2(n13338), .ZN(n13351) );
  NAND2_X1 U8425 ( .A1(n10077), .A2(n9837), .ZN(n15289) );
  NAND2_X1 U8426 ( .A1(n13174), .A2(n13173), .ZN(n15132) );
  OR2_X1 U8427 ( .A1(n15242), .A2(n13262), .ZN(n13174) );
  NAND2_X1 U8428 ( .A1(n9786), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n9744) );
  NAND2_X1 U8429 ( .A1(n9788), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n8691) );
  NAND2_X1 U8430 ( .A1(n7862), .A2(n15168), .ZN(n7861) );
  AND2_X1 U8431 ( .A1(n15184), .A2(n15137), .ZN(n8016) );
  INV_X1 U8432 ( .A(n15359), .ZN(n15369) );
  NAND2_X1 U8433 ( .A1(n16148), .A2(n9829), .ZN(n15364) );
  INV_X1 U8434 ( .A(n7854), .ZN(n7853) );
  OR2_X1 U8435 ( .A1(n10408), .A2(n10463), .ZN(n7855) );
  NAND3_X1 U8436 ( .A1(n8692), .A2(n8693), .A3(n7976), .ZN(n15520) );
  NOR2_X1 U8437 ( .A1(P2_IR_REG_28__SCAN_IN), .A2(P2_IR_REG_29__SCAN_IN), .ZN(
        n7976) );
  NAND2_X1 U8438 ( .A1(n15549), .A2(n15550), .ZN(n15548) );
  NAND2_X1 U8439 ( .A1(n12321), .A2(n12320), .ZN(n13736) );
  NAND2_X1 U8440 ( .A1(n7798), .A2(n7797), .ZN(n15559) );
  OAI21_X1 U8441 ( .B1(n12913), .B2(n7784), .A(n7782), .ZN(n7785) );
  AOI21_X1 U8442 ( .B1(n15550), .B2(n7783), .A(n12926), .ZN(n7782) );
  INV_X1 U8443 ( .A(n15550), .ZN(n7784) );
  INV_X1 U8444 ( .A(n15656), .ZN(n7783) );
  OR2_X1 U8445 ( .A1(n10393), .A2(n10386), .ZN(n15673) );
  XNOR2_X1 U8446 ( .A(n8050), .B(n15783), .ZN(n16003) );
  NAND2_X1 U8447 ( .A1(n15801), .A2(n8051), .ZN(n8050) );
  NAND2_X1 U8448 ( .A1(n16011), .A2(n15791), .ZN(n8051) );
  NAND2_X1 U8449 ( .A1(n8613), .A2(n8614), .ZN(n15803) );
  NAND2_X1 U8450 ( .A1(n8558), .A2(n8557), .ZN(n8556) );
  OAI21_X1 U8451 ( .B1(n8560), .B2(n15804), .A(n15799), .ZN(n8559) );
  NAND2_X1 U8452 ( .A1(n15800), .A2(n16462), .ZN(n8557) );
  NAND2_X1 U8453 ( .A1(n8617), .A2(n8616), .ZN(n15812) );
  NAND2_X1 U8454 ( .A1(n7716), .A2(n15814), .ZN(n7715) );
  NAND2_X1 U8455 ( .A1(n8617), .A2(n7482), .ZN(n7716) );
  NAND2_X1 U8456 ( .A1(n8626), .A2(n8627), .ZN(n11747) );
  OR2_X1 U8457 ( .A1(n11572), .A2(n13580), .ZN(n8626) );
  NAND2_X1 U8458 ( .A1(n7658), .A2(n16299), .ZN(n16301) );
  NAND2_X1 U8459 ( .A1(n16297), .A2(n16298), .ZN(n7658) );
  XNOR2_X1 U8460 ( .A(n16338), .B(n8520), .ZN(n16339) );
  INV_X1 U8461 ( .A(n16337), .ZN(n8520) );
  XNOR2_X1 U8462 ( .A(n16349), .B(n16350), .ZN(n16351) );
  XNOR2_X1 U8463 ( .A(n8518), .B(n7666), .ZN(n16357) );
  INV_X1 U8464 ( .A(n16355), .ZN(n7666) );
  OR2_X1 U8465 ( .A1(n16388), .A2(P2_ADDR_REG_16__SCAN_IN), .ZN(n8516) );
  NAND2_X1 U8466 ( .A1(n7655), .A2(n7654), .ZN(n7653) );
  INV_X1 U8467 ( .A(n16408), .ZN(n7654) );
  INV_X1 U8468 ( .A(n7656), .ZN(n7655) );
  XNOR2_X1 U8469 ( .A(n7656), .B(n16408), .ZN(n16409) );
  NAND2_X1 U8470 ( .A1(n8059), .A2(n8058), .ZN(n13664) );
  NAND2_X1 U8471 ( .A1(n13663), .A2(n13612), .ZN(n8058) );
  NAND2_X1 U8472 ( .A1(n8060), .A2(n13779), .ZN(n8059) );
  NAND2_X1 U8473 ( .A1(n13662), .A2(n13661), .ZN(n8060) );
  OR2_X1 U8474 ( .A1(n13612), .A2(n16466), .ZN(n8055) );
  INV_X1 U8475 ( .A(n13665), .ZN(n13654) );
  NAND2_X1 U8476 ( .A1(n14660), .A2(n8240), .ZN(n8239) );
  NAND2_X1 U8477 ( .A1(keyinput_134), .A2(SI_26_), .ZN(n8240) );
  AOI22_X1 U8478 ( .A1(n14914), .A2(keyinput_131), .B1(SI_30_), .B2(
        keyinput_130), .ZN(n14648) );
  NOR2_X1 U8479 ( .A1(n14658), .A2(n14659), .ZN(n8238) );
  NAND2_X1 U8480 ( .A1(n14663), .A2(n14664), .ZN(n8235) );
  NAND2_X1 U8481 ( .A1(keyinput_140), .A2(SI_20_), .ZN(n8234) );
  AOI21_X1 U8482 ( .B1(n8237), .B2(n8236), .A(n8233), .ZN(n14670) );
  AOI22_X1 U8483 ( .A1(n14662), .A2(n14661), .B1(keyinput_139), .B2(SI_21_), 
        .ZN(n8236) );
  NAND2_X1 U8484 ( .A1(n8235), .A2(n8234), .ZN(n8233) );
  OAI21_X1 U8485 ( .B1(n14652), .B2(n8239), .A(n8238), .ZN(n8237) );
  NAND2_X1 U8486 ( .A1(n8800), .A2(n8801), .ZN(n8798) );
  INV_X1 U8487 ( .A(n14482), .ZN(n8484) );
  AOI221_X1 U8488 ( .B1(SI_31_), .B2(keyinput_1), .C1(keyinput_0), .C2(
        P3_WR_REG_SCAN_IN), .A(n14479), .ZN(n14480) );
  NAND2_X1 U8489 ( .A1(n14483), .A2(keyinput_6), .ZN(n8483) );
  OAI22_X1 U8490 ( .A1(n13700), .A2(n7967), .B1(n13701), .B2(n7966), .ZN(
        n13705) );
  INV_X1 U8491 ( .A(n13699), .ZN(n7966) );
  NOR2_X1 U8492 ( .A1(n13702), .A2(n13699), .ZN(n7967) );
  OAI22_X1 U8493 ( .A1(n14678), .A2(n14679), .B1(SI_11_), .B2(keyinput_149), 
        .ZN(n8209) );
  NAND2_X1 U8494 ( .A1(n14675), .A2(n8211), .ZN(n8210) );
  INV_X1 U8495 ( .A(n8212), .ZN(n8211) );
  OAI22_X1 U8496 ( .A1(SI_12_), .A2(n14677), .B1(n14676), .B2(keyinput_148), 
        .ZN(n8212) );
  NAND2_X1 U8497 ( .A1(n7746), .A2(n13059), .ZN(n7744) );
  OAI21_X1 U8498 ( .B1(n7746), .B2(n13059), .A(n13060), .ZN(n7745) );
  INV_X1 U8499 ( .A(n13712), .ZN(n7963) );
  AOI21_X1 U8500 ( .B1(n8480), .B2(n8477), .A(n8474), .ZN(n14496) );
  NAND2_X1 U8501 ( .A1(n8204), .A2(n8203), .ZN(n14693) );
  INV_X1 U8502 ( .A(n14688), .ZN(n8203) );
  NAND2_X1 U8503 ( .A1(n8206), .A2(n8205), .ZN(n8204) );
  NOR2_X1 U8504 ( .A1(n13080), .A2(n7509), .ZN(n8810) );
  INV_X1 U8505 ( .A(n13072), .ZN(n8025) );
  NAND2_X1 U8506 ( .A1(n13716), .A2(n13718), .ZN(n8115) );
  AND2_X1 U8507 ( .A1(n8199), .A2(n8198), .ZN(n14708) );
  INV_X1 U8508 ( .A(n14700), .ZN(n8198) );
  OAI21_X1 U8509 ( .B1(n8201), .B2(n8200), .A(n14701), .ZN(n8199) );
  AOI21_X1 U8510 ( .B1(n8465), .B2(n7615), .A(n8463), .ZN(n14517) );
  NAND2_X1 U8511 ( .A1(n7625), .A2(n8464), .ZN(n8463) );
  OAI21_X1 U8512 ( .B1(n14511), .B2(n8466), .A(n7598), .ZN(n8465) );
  NAND2_X1 U8513 ( .A1(n7595), .A2(n8105), .ZN(n7742) );
  NOR2_X1 U8514 ( .A1(n7595), .A2(n8105), .ZN(n7743) );
  INV_X1 U8515 ( .A(n13099), .ZN(n8804) );
  INV_X1 U8516 ( .A(n8803), .ZN(n7755) );
  INV_X1 U8517 ( .A(n8167), .ZN(n13360) );
  INV_X1 U8518 ( .A(n8223), .ZN(n8222) );
  OAI22_X1 U8519 ( .A1(n14715), .A2(n14714), .B1(P3_REG3_REG_16__SCAN_IN), 
        .B2(keyinput_176), .ZN(n8223) );
  NAND2_X1 U8520 ( .A1(n8804), .A2(n7510), .ZN(n8803) );
  INV_X1 U8521 ( .A(n7753), .ZN(n7751) );
  NAND2_X1 U8522 ( .A1(n7947), .A2(n7946), .ZN(n13742) );
  AOI21_X1 U8523 ( .B1(n7488), .B2(n7950), .A(n7427), .ZN(n7946) );
  NAND2_X1 U8524 ( .A1(n8221), .A2(n8219), .ZN(n8218) );
  INV_X1 U8525 ( .A(n8220), .ZN(n8219) );
  NAND2_X1 U8526 ( .A1(n14713), .A2(n8222), .ZN(n8221) );
  OAI22_X1 U8527 ( .A1(n14716), .A2(keyinput_177), .B1(n14717), .B2(
        P3_REG3_REG_5__SCAN_IN), .ZN(n8220) );
  NAND2_X1 U8528 ( .A1(n16509), .A2(keyinput_187), .ZN(n8215) );
  NAND2_X1 U8529 ( .A1(n14723), .A2(P3_REG3_REG_2__SCAN_IN), .ZN(n8214) );
  OR2_X1 U8530 ( .A1(n14530), .A2(n14531), .ZN(n8473) );
  XNOR2_X1 U8531 ( .A(n14712), .B(keyinput_47), .ZN(n8472) );
  NAND2_X1 U8532 ( .A1(n14716), .A2(keyinput_49), .ZN(n8469) );
  NAND2_X1 U8533 ( .A1(n14533), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n8468) );
  AOI21_X1 U8534 ( .B1(n8471), .B2(n8470), .A(n8467), .ZN(n14546) );
  AOI22_X1 U8535 ( .A1(n14715), .A2(n14532), .B1(keyinput_48), .B2(
        P3_REG3_REG_16__SCAN_IN), .ZN(n8470) );
  NAND2_X1 U8536 ( .A1(n8469), .A2(n8468), .ZN(n8467) );
  NAND2_X1 U8537 ( .A1(n8473), .A2(n8472), .ZN(n8471) );
  INV_X1 U8538 ( .A(n13109), .ZN(n8784) );
  INV_X1 U8539 ( .A(n13121), .ZN(n8792) );
  OR2_X1 U8540 ( .A1(n7939), .A2(n13751), .ZN(n7938) );
  XNOR2_X1 U8541 ( .A(n14762), .B(n8232), .ZN(n8231) );
  NAND2_X1 U8542 ( .A1(n8226), .A2(n8225), .ZN(n8224) );
  INV_X1 U8543 ( .A(n14770), .ZN(n8225) );
  NOR2_X1 U8544 ( .A1(n14769), .A2(n14771), .ZN(n8226) );
  AND2_X1 U8545 ( .A1(n8229), .A2(n8228), .ZN(n8227) );
  NAND2_X1 U8546 ( .A1(n14764), .A2(P3_DATAO_REG_12__SCAN_IN), .ZN(n8228) );
  NAND2_X1 U8547 ( .A1(n14763), .A2(keyinput_212), .ZN(n8229) );
  NOR2_X1 U8548 ( .A1(n13137), .A2(n13138), .ZN(n7761) );
  NAND2_X1 U8549 ( .A1(n8805), .A2(n7762), .ZN(n7758) );
  OAI21_X1 U8550 ( .B1(n13127), .B2(n13126), .A(n7550), .ZN(n8805) );
  INV_X1 U8551 ( .A(n13134), .ZN(n8807) );
  NAND2_X1 U8552 ( .A1(n7941), .A2(n7940), .ZN(n13763) );
  AOI21_X1 U8553 ( .B1(n7419), .B2(n7441), .A(n7426), .ZN(n7940) );
  AND2_X1 U8554 ( .A1(n7419), .A2(n7943), .ZN(n7942) );
  INV_X1 U8555 ( .A(n14571), .ZN(n8461) );
  XNOR2_X1 U8556 ( .A(n14762), .B(n8460), .ZN(n8459) );
  INV_X1 U8557 ( .A(keyinput_82), .ZN(n8460) );
  OAI22_X1 U8558 ( .A1(n14763), .A2(n14572), .B1(P3_DATAO_REG_12__SCAN_IN), 
        .B2(keyinput_84), .ZN(n8457) );
  NAND2_X1 U8559 ( .A1(n14791), .A2(n16311), .ZN(n8250) );
  OAI21_X1 U8560 ( .B1(n8462), .B2(n8458), .A(n8456), .ZN(n14573) );
  INV_X1 U8561 ( .A(n8457), .ZN(n8456) );
  NAND2_X1 U8562 ( .A1(n8461), .A2(n8459), .ZN(n8458) );
  AOI211_X1 U8563 ( .C1(n14568), .C2(n14569), .A(n14567), .B(n14566), .ZN(
        n8462) );
  INV_X1 U8564 ( .A(n13153), .ZN(n8791) );
  OAI21_X1 U8565 ( .B1(n7954), .B2(n7541), .A(n7435), .ZN(n7953) );
  NOR2_X1 U8566 ( .A1(n13767), .A2(n7955), .ZN(n7954) );
  OR2_X1 U8567 ( .A1(n14790), .A2(n8248), .ZN(n8247) );
  NAND2_X1 U8568 ( .A1(n8250), .A2(n8249), .ZN(n8248) );
  NAND2_X1 U8569 ( .A1(keyinput_231), .A2(P3_ADDR_REG_6__SCAN_IN), .ZN(n8249)
         );
  AOI22_X1 U8570 ( .A1(n16316), .A2(n14792), .B1(keyinput_232), .B2(
        P3_ADDR_REG_7__SCAN_IN), .ZN(n8246) );
  NAND2_X1 U8571 ( .A1(n14794), .A2(n16439), .ZN(n8243) );
  NAND2_X1 U8572 ( .A1(keyinput_234), .A2(P3_ADDR_REG_9__SCAN_IN), .ZN(n8242)
         );
  AND2_X1 U8573 ( .A1(n8788), .A2(n13163), .ZN(n8787) );
  NAND2_X1 U8574 ( .A1(n8790), .A2(n8789), .ZN(n8788) );
  NAND2_X1 U8575 ( .A1(n8791), .A2(n7511), .ZN(n8789) );
  AOI21_X1 U8576 ( .B1(n8245), .B2(n8244), .A(n8241), .ZN(n14795) );
  AOI22_X1 U8577 ( .A1(n11611), .A2(n14793), .B1(keyinput_233), .B2(
        P3_ADDR_REG_8__SCAN_IN), .ZN(n8244) );
  NAND2_X1 U8578 ( .A1(n8243), .A2(n8242), .ZN(n8241) );
  NAND2_X1 U8579 ( .A1(n8247), .A2(n8246), .ZN(n8245) );
  NAND2_X1 U8580 ( .A1(n14595), .A2(n16311), .ZN(n8494) );
  INV_X1 U8581 ( .A(n8396), .ZN(n8395) );
  OR2_X1 U8582 ( .A1(n14594), .A2(n8492), .ZN(n8491) );
  NAND2_X1 U8583 ( .A1(n8494), .A2(n8493), .ZN(n8492) );
  NAND2_X1 U8584 ( .A1(keyinput_103), .A2(P3_ADDR_REG_6__SCAN_IN), .ZN(n8493)
         );
  AOI22_X1 U8585 ( .A1(n16316), .A2(n14596), .B1(keyinput_104), .B2(
        P3_ADDR_REG_7__SCAN_IN), .ZN(n8490) );
  NAND2_X1 U8586 ( .A1(n14598), .A2(n16439), .ZN(n8487) );
  NAND2_X1 U8587 ( .A1(keyinput_106), .A2(P3_ADDR_REG_9__SCAN_IN), .ZN(n8486)
         );
  NAND2_X1 U8588 ( .A1(n7539), .A2(n8796), .ZN(n8795) );
  OAI22_X1 U8589 ( .A1(n13784), .A2(n7936), .B1(n13785), .B2(n7937), .ZN(
        n13788) );
  AND2_X1 U8590 ( .A1(n13785), .A2(n7937), .ZN(n7936) );
  INV_X1 U8591 ( .A(n13783), .ZN(n7937) );
  NAND2_X1 U8592 ( .A1(n7613), .A2(n12633), .ZN(n8392) );
  AND2_X1 U8593 ( .A1(n14083), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n7691) );
  AOI21_X1 U8594 ( .B1(n8489), .B2(n8488), .A(n8485), .ZN(n14602) );
  AOI22_X1 U8595 ( .A1(n11611), .A2(n14597), .B1(keyinput_105), .B2(
        P3_ADDR_REG_8__SCAN_IN), .ZN(n8488) );
  NAND2_X1 U8596 ( .A1(n8487), .A2(n8486), .ZN(n8485) );
  NAND2_X1 U8597 ( .A1(n8491), .A2(n8490), .ZN(n8489) );
  INV_X1 U8598 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n8875) );
  NAND2_X1 U8599 ( .A1(n7525), .A2(n8687), .ZN(n8686) );
  NAND2_X1 U8600 ( .A1(n8074), .A2(n13615), .ZN(n13632) );
  INV_X1 U8601 ( .A(n12629), .ZN(n8036) );
  INV_X1 U8602 ( .A(n8392), .ZN(n8035) );
  AND2_X1 U8603 ( .A1(n8666), .A2(n12625), .ZN(n8665) );
  INV_X1 U8604 ( .A(n12150), .ZN(n8682) );
  INV_X1 U8605 ( .A(n11742), .ZN(n8387) );
  NAND2_X1 U8606 ( .A1(n10001), .A2(n8006), .ZN(n8005) );
  INV_X1 U8607 ( .A(n8393), .ZN(n8004) );
  NOR2_X1 U8608 ( .A1(n9957), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n10637) );
  AOI21_X1 U8609 ( .B1(n9954), .B2(n7991), .A(n7547), .ZN(n7989) );
  AND2_X1 U8610 ( .A1(n7519), .A2(n7642), .ZN(n16282) );
  NOR2_X1 U8611 ( .A1(n16274), .A2(P1_ADDR_REG_0__SCAN_IN), .ZN(n8525) );
  OAI21_X1 U8612 ( .B1(n13485), .B2(n13484), .A(n8076), .ZN(n8075) );
  NAND2_X1 U8613 ( .A1(n7683), .A2(n7682), .ZN(n7685) );
  AND2_X1 U8614 ( .A1(n7685), .A2(n9675), .ZN(n8852) );
  OAI21_X1 U8615 ( .B1(n10922), .B2(n8427), .A(n7684), .ZN(n10907) );
  NAND2_X1 U8616 ( .A1(n8428), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n8427) );
  NAND2_X1 U8617 ( .A1(n8852), .A2(n8428), .ZN(n7684) );
  INV_X1 U8618 ( .A(n10908), .ZN(n8428) );
  NOR2_X1 U8619 ( .A1(n10904), .A2(n7815), .ZN(n9657) );
  NOR2_X1 U8620 ( .A1(n7816), .A2(n9616), .ZN(n7815) );
  AOI21_X1 U8621 ( .B1(n9855), .B2(P3_REG2_REG_6__SCAN_IN), .A(n10907), .ZN(
        n9677) );
  INV_X1 U8622 ( .A(n9665), .ZN(n7814) );
  AND2_X1 U8623 ( .A1(n8192), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n7812) );
  AOI21_X1 U8624 ( .B1(n13997), .B2(P3_REG1_REG_12__SCAN_IN), .A(n13992), .ZN(
        n13993) );
  NAND2_X1 U8625 ( .A1(n14049), .A2(n14048), .ZN(n14062) );
  NAND2_X1 U8626 ( .A1(n8177), .A2(n7617), .ZN(n8176) );
  NAND2_X1 U8627 ( .A1(n7475), .A2(n14098), .ZN(n8425) );
  NAND2_X1 U8628 ( .A1(n8421), .A2(n14108), .ZN(n8423) );
  INV_X1 U8629 ( .A(n7475), .ZN(n8421) );
  NAND2_X1 U8630 ( .A1(n8425), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n8424) );
  NOR2_X1 U8631 ( .A1(n9343), .A2(n14158), .ZN(n13509) );
  NAND2_X1 U8632 ( .A1(n9510), .A2(n8350), .ZN(n8142) );
  NAND2_X1 U8633 ( .A1(n8146), .A2(n9498), .ZN(n8145) );
  AOI21_X1 U8634 ( .B1(n8151), .B2(n9258), .A(n7424), .ZN(n8149) );
  NOR2_X1 U8635 ( .A1(n8150), .A2(n7594), .ZN(n8146) );
  INV_X1 U8636 ( .A(n8151), .ZN(n8150) );
  INV_X1 U8637 ( .A(n8355), .ZN(n14258) );
  OAI21_X1 U8638 ( .B1(n14315), .B2(n9367), .A(n9370), .ZN(n8355) );
  OR2_X1 U8639 ( .A1(n9182), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n9197) );
  NOR2_X1 U8640 ( .A1(n7467), .A2(n11938), .ZN(n9103) );
  NAND2_X1 U8641 ( .A1(n13387), .A2(n8339), .ZN(n11938) );
  NAND2_X1 U8642 ( .A1(n10517), .A2(n16494), .ZN(n13364) );
  INV_X1 U8643 ( .A(n14619), .ZN(n8446) );
  AND2_X1 U8644 ( .A1(n8449), .A2(n8448), .ZN(n8447) );
  INV_X1 U8645 ( .A(n8453), .ZN(n8448) );
  OR2_X1 U8646 ( .A1(n8455), .A2(n8454), .ZN(n8449) );
  OAI22_X1 U8647 ( .A1(n10144), .A2(keyinput_118), .B1(n14615), .B2(
        P1_IR_REG_11__SCAN_IN), .ZN(n8453) );
  INV_X1 U8648 ( .A(n14618), .ZN(n8452) );
  INV_X1 U8649 ( .A(n8454), .ZN(n8450) );
  INV_X1 U8650 ( .A(n14613), .ZN(n8451) );
  OR2_X1 U8651 ( .A1(P3_IR_REG_26__SCAN_IN), .A2(P3_IR_REG_27__SCAN_IN), .ZN(
        n8885) );
  NOR2_X1 U8652 ( .A1(n8750), .A2(n8748), .ZN(n8747) );
  NOR2_X1 U8653 ( .A1(P3_IR_REG_22__SCAN_IN), .A2(P3_IR_REG_25__SCAN_IN), .ZN(
        n7763) );
  INV_X1 U8654 ( .A(n8914), .ZN(n7825) );
  INV_X1 U8655 ( .A(n7824), .ZN(n7823) );
  OAI21_X1 U8656 ( .B1(n9188), .B2(n7825), .A(n9207), .ZN(n7824) );
  AND3_X1 U8657 ( .A1(n8881), .A2(n8880), .A3(n8879), .ZN(n9165) );
  AND2_X1 U8658 ( .A1(n9176), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n8564) );
  INV_X1 U8659 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n9168) );
  INV_X1 U8660 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n8745) );
  INV_X1 U8661 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n11081) );
  INV_X1 U8662 ( .A(n10650), .ZN(n8502) );
  NOR2_X1 U8663 ( .A1(n15274), .A2(n15256), .ZN(n8323) );
  NOR2_X1 U8664 ( .A1(n8008), .A2(n15511), .ZN(n7667) );
  NOR2_X1 U8665 ( .A1(n11777), .A2(n16700), .ZN(n8320) );
  OR2_X1 U8666 ( .A1(n11082), .A2(n11081), .ZN(n11095) );
  NAND2_X1 U8667 ( .A1(n11642), .A2(n7671), .ZN(n11596) );
  NOR2_X1 U8668 ( .A1(n13077), .A2(n13071), .ZN(n7671) );
  OR2_X1 U8669 ( .A1(n11070), .A2(n11069), .ZN(n11082) );
  NOR2_X1 U8670 ( .A1(n11265), .A2(n11250), .ZN(n8765) );
  NAND2_X1 U8671 ( .A1(n10519), .A2(n8766), .ZN(n8764) );
  AND2_X1 U8672 ( .A1(n10467), .A2(n8767), .ZN(n8766) );
  NAND2_X1 U8673 ( .A1(n11265), .A2(n11250), .ZN(n8767) );
  AOI21_X1 U8674 ( .B1(n13312), .B2(n7867), .A(n7513), .ZN(n7866) );
  NAND2_X1 U8675 ( .A1(n7865), .A2(n7867), .ZN(n7864) );
  INV_X1 U8676 ( .A(n8323), .ZN(n15257) );
  XNOR2_X1 U8677 ( .A(n9723), .B(P2_IR_REG_21__SCAN_IN), .ZN(n9730) );
  INV_X1 U8678 ( .A(n11977), .ZN(n8066) );
  INV_X1 U8679 ( .A(n11978), .ZN(n8065) );
  NAND2_X1 U8680 ( .A1(n11694), .A2(n11695), .ZN(n8826) );
  AND2_X1 U8681 ( .A1(n11563), .A2(n10571), .ZN(n11859) );
  NOR2_X1 U8682 ( .A1(n12403), .A2(n8835), .ZN(n8834) );
  INV_X1 U8683 ( .A(n8838), .ZN(n8835) );
  INV_X1 U8684 ( .A(n12874), .ZN(n8814) );
  AND2_X1 U8685 ( .A1(n13603), .A2(n8404), .ZN(n8403) );
  NOR2_X1 U8686 ( .A1(n8406), .A2(n8405), .ZN(n8404) );
  NAND2_X1 U8687 ( .A1(n15808), .A2(n8306), .ZN(n8305) );
  NOR2_X1 U8688 ( .A1(n15819), .A2(n16021), .ZN(n8306) );
  NAND2_X1 U8689 ( .A1(n15819), .A2(n13570), .ZN(n15780) );
  INV_X1 U8690 ( .A(n15890), .ZN(n7705) );
  NAND2_X1 U8691 ( .A1(n8308), .A2(n7721), .ZN(n7725) );
  NOR2_X1 U8692 ( .A1(n7723), .A2(n15906), .ZN(n7721) );
  NOR2_X1 U8693 ( .A1(n12351), .A2(n12350), .ZN(n12349) );
  INV_X1 U8694 ( .A(n8635), .ZN(n7712) );
  INV_X1 U8695 ( .A(n15682), .ZN(n11997) );
  OR2_X1 U8696 ( .A1(n11550), .A2(n11704), .ZN(n11565) );
  NAND2_X1 U8697 ( .A1(n8545), .A2(n8544), .ZN(n8543) );
  NAND2_X1 U8698 ( .A1(n12759), .A2(n10731), .ZN(n7676) );
  NAND2_X1 U8699 ( .A1(n16463), .A2(n10934), .ZN(n13668) );
  NOR2_X1 U8700 ( .A1(n8046), .A2(n16527), .ZN(n7732) );
  NAND2_X1 U8701 ( .A1(n8308), .A2(n7722), .ZN(n15921) );
  INV_X1 U8702 ( .A(n13215), .ZN(n8679) );
  AOI21_X1 U8703 ( .B1(n8678), .B2(n8676), .A(n8675), .ZN(n8674) );
  INV_X1 U8704 ( .A(n13217), .ZN(n8675) );
  INV_X1 U8705 ( .A(n12642), .ZN(n8676) );
  INV_X1 U8706 ( .A(n9563), .ZN(n9559) );
  NAND2_X1 U8707 ( .A1(n12512), .A2(SI_21_), .ZN(n12513) );
  NAND2_X1 U8708 ( .A1(n9991), .A2(n9930), .ZN(n7805) );
  INV_X1 U8709 ( .A(n8681), .ZN(n8376) );
  INV_X1 U8710 ( .A(n10627), .ZN(n10625) );
  OR2_X1 U8711 ( .A1(n9941), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n9957) );
  INV_X1 U8712 ( .A(n7985), .ZN(n7984) );
  OAI21_X1 U8713 ( .B1(n9874), .B2(P2_DATAO_REG_3__SCAN_IN), .A(n9770), .ZN(
        n9867) );
  NAND2_X1 U8714 ( .A1(n9874), .A2(n9895), .ZN(n9770) );
  INV_X1 U8715 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n8379) );
  XNOR2_X1 U8716 ( .A(P1_ADDR_REG_1__SCAN_IN), .B(P3_ADDR_REG_1__SCAN_IN), 
        .ZN(n8526) );
  XNOR2_X1 U8717 ( .A(n16282), .B(n16281), .ZN(n16283) );
  NOR2_X1 U8718 ( .A1(n16286), .A2(n16287), .ZN(n16292) );
  XNOR2_X1 U8719 ( .A(n16292), .B(n8522), .ZN(n7648) );
  NOR2_X1 U8720 ( .A1(n16319), .A2(n16318), .ZN(n16328) );
  AOI21_X1 U8721 ( .B1(n16386), .B2(P3_ADDR_REG_16__SCAN_IN), .A(n16387), .ZN(
        n16392) );
  XNOR2_X1 U8722 ( .A(n16392), .B(n7644), .ZN(n16393) );
  INV_X1 U8723 ( .A(n8516), .ZN(n7651) );
  AOI21_X1 U8724 ( .B1(n8723), .B2(n8721), .A(n7481), .ZN(n7882) );
  INV_X1 U8725 ( .A(n11660), .ZN(n8721) );
  INV_X1 U8726 ( .A(n8723), .ZN(n8722) );
  NAND2_X1 U8727 ( .A1(n7906), .A2(n9519), .ZN(n7905) );
  INV_X1 U8728 ( .A(n9520), .ZN(n7906) );
  AOI21_X1 U8729 ( .B1(n7907), .B2(n9518), .A(n7904), .ZN(n7903) );
  NOR2_X1 U8730 ( .A1(n13965), .A2(n7905), .ZN(n7904) );
  NAND2_X1 U8731 ( .A1(n9453), .A2(n11817), .ZN(n8732) );
  INV_X1 U8732 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n14641) );
  AND2_X1 U8733 ( .A1(n9515), .A2(n9513), .ZN(n13886) );
  XNOR2_X1 U8734 ( .A(n9450), .B(n11931), .ZN(n9460) );
  INV_X1 U8735 ( .A(n9503), .ZN(n8737) );
  INV_X1 U8736 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n14535) );
  NAND2_X1 U8737 ( .A1(n9463), .A2(n13396), .ZN(n7886) );
  NOR2_X1 U8738 ( .A1(n9249), .A2(n8868), .ZN(n9264) );
  AND2_X1 U8739 ( .A1(n9264), .A2(n13926), .ZN(n9273) );
  AND2_X1 U8740 ( .A1(n13416), .A2(n13412), .ZN(n13533) );
  AND2_X1 U8741 ( .A1(n7501), .A2(n11680), .ZN(n8723) );
  NAND2_X1 U8742 ( .A1(n8870), .A2(n14712), .ZN(n9323) );
  INV_X1 U8743 ( .A(n7411), .ZN(n9326) );
  NAND2_X1 U8744 ( .A1(n9287), .A2(P3_REG3_REG_2__SCAN_IN), .ZN(n8365) );
  OR2_X1 U8745 ( .A1(n10998), .A2(n8363), .ZN(n8362) );
  NAND2_X1 U8746 ( .A1(n8980), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n8364) );
  INV_X1 U8747 ( .A(P3_ADDR_REG_1__SCAN_IN), .ZN(n16272) );
  NAND2_X1 U8748 ( .A1(n8409), .A2(n8407), .ZN(n10889) );
  OAI22_X1 U8749 ( .A1(n11221), .A2(n11222), .B1(P3_REG1_REG_2__SCAN_IN), .B2(
        n11234), .ZN(n11220) );
  INV_X1 U8750 ( .A(P3_ADDR_REG_2__SCAN_IN), .ZN(n16281) );
  NOR2_X1 U8751 ( .A1(n10855), .A2(n11820), .ZN(n11193) );
  NAND2_X1 U8752 ( .A1(n10854), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n11198) );
  XNOR2_X1 U8753 ( .A(n7685), .B(n9675), .ZN(n10922) );
  NOR2_X1 U8754 ( .A1(n10922), .A2(n11928), .ZN(n10921) );
  NOR2_X1 U8755 ( .A1(n11518), .A2(n9621), .ZN(n11517) );
  INV_X1 U8756 ( .A(n8420), .ZN(n9678) );
  OAI22_X1 U8757 ( .A1(n8185), .A2(n7605), .B1(n8187), .B2(n8183), .ZN(n8182)
         );
  AND2_X1 U8758 ( .A1(n8418), .A2(n9681), .ZN(n11958) );
  NAND2_X1 U8759 ( .A1(n8416), .A2(n8415), .ZN(n12161) );
  NAND2_X1 U8760 ( .A1(n8038), .A2(n12166), .ZN(n8416) );
  INV_X1 U8761 ( .A(n8414), .ZN(n12160) );
  NAND2_X1 U8762 ( .A1(n8196), .A2(n8195), .ZN(n9663) );
  AOI21_X1 U8763 ( .B1(n12157), .B2(n7739), .A(n7596), .ZN(n7738) );
  INV_X1 U8764 ( .A(n9635), .ZN(n7739) );
  AND2_X1 U8765 ( .A1(n8414), .A2(n8415), .ZN(n9686) );
  NOR2_X1 U8766 ( .A1(n9686), .A2(n9687), .ZN(n13996) );
  OR2_X1 U8767 ( .A1(n8189), .A2(n14010), .ZN(n13994) );
  AND2_X1 U8768 ( .A1(n13993), .A2(n14024), .ZN(n8189) );
  AND2_X1 U8769 ( .A1(n8432), .A2(n8431), .ZN(n14016) );
  OR2_X1 U8770 ( .A1(n14029), .A2(n14030), .ZN(n14049) );
  NAND2_X1 U8771 ( .A1(n7698), .A2(n7622), .ZN(n14070) );
  NAND2_X1 U8772 ( .A1(n14040), .A2(n8434), .ZN(n7698) );
  OR2_X1 U8773 ( .A1(n14063), .A2(n8435), .ZN(n8434) );
  NAND2_X1 U8774 ( .A1(n8188), .A2(n7630), .ZN(n7841) );
  NAND2_X1 U8775 ( .A1(n7841), .A2(n14108), .ZN(n14101) );
  NAND2_X1 U8776 ( .A1(n14111), .A2(n14110), .ZN(n14138) );
  NAND2_X1 U8777 ( .A1(n13520), .A2(n7470), .ZN(n8132) );
  AND2_X1 U8778 ( .A1(n13356), .A2(n13355), .ZN(n14163) );
  AOI21_X1 U8779 ( .B1(n8137), .B2(n8138), .A(n7526), .ZN(n8134) );
  NAND2_X1 U8780 ( .A1(n14186), .A2(n8345), .ZN(n8344) );
  INV_X1 U8781 ( .A(n14221), .ZN(n14216) );
  AND2_X1 U8782 ( .A1(n7898), .A2(n8144), .ZN(n14229) );
  OR2_X1 U8783 ( .A1(n14296), .A2(n8145), .ZN(n7898) );
  OR2_X1 U8784 ( .A1(n13459), .A2(n13458), .ZN(n14230) );
  NAND2_X1 U8785 ( .A1(n8148), .A2(n8149), .ZN(n14244) );
  OR2_X1 U8786 ( .A1(n14296), .A2(n8143), .ZN(n8148) );
  INV_X1 U8787 ( .A(n8146), .ZN(n8143) );
  AND2_X1 U8788 ( .A1(n13456), .A2(n13455), .ZN(n14245) );
  AOI21_X1 U8789 ( .B1(n14276), .B2(n9259), .A(n9258), .ZN(n14263) );
  AND2_X1 U8790 ( .A1(n13451), .A2(n13452), .ZN(n14262) );
  NOR2_X1 U8791 ( .A1(n14296), .A2(n7594), .ZN(n14276) );
  AND2_X1 U8792 ( .A1(n13447), .A2(n13446), .ZN(n14285) );
  OR2_X1 U8793 ( .A1(n9235), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n9249) );
  NAND2_X1 U8794 ( .A1(n7883), .A2(n9175), .ZN(n14359) );
  NAND2_X1 U8795 ( .A1(n8158), .A2(n8160), .ZN(n7883) );
  OR2_X1 U8796 ( .A1(n14359), .A2(n14366), .ZN(n14360) );
  NAND2_X1 U8797 ( .A1(n9365), .A2(n13425), .ZN(n14367) );
  AND2_X1 U8798 ( .A1(n13426), .A2(n13427), .ZN(n14366) );
  AND3_X1 U8799 ( .A1(n9153), .A2(n9152), .A3(n9151), .ZN(n13877) );
  AND2_X1 U8800 ( .A1(n8166), .A2(n7486), .ZN(n14377) );
  NAND2_X1 U8801 ( .A1(n12392), .A2(n9139), .ZN(n8166) );
  OR2_X1 U8802 ( .A1(n9126), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n9140) );
  NAND2_X1 U8803 ( .A1(n8368), .A2(n8366), .ZN(n12391) );
  AOI21_X1 U8804 ( .B1(n8369), .B2(n13395), .A(n8367), .ZN(n8366) );
  INV_X1 U8805 ( .A(n13407), .ZN(n8367) );
  OR2_X1 U8806 ( .A1(n9108), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n9126) );
  OR2_X1 U8807 ( .A1(n9087), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n9089) );
  AND2_X1 U8808 ( .A1(n12041), .A2(n9104), .ZN(n12233) );
  NAND2_X1 U8809 ( .A1(n13532), .A2(n8338), .ZN(n8337) );
  OR2_X1 U8810 ( .A1(n9041), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n9058) );
  NAND2_X1 U8811 ( .A1(n11923), .A2(n9040), .ZN(n12247) );
  AOI21_X1 U8812 ( .B1(n13527), .B2(n8332), .A(n8331), .ZN(n8330) );
  INV_X1 U8813 ( .A(n13370), .ZN(n8331) );
  INV_X1 U8814 ( .A(n13368), .ZN(n8332) );
  NAND2_X1 U8815 ( .A1(n8167), .A2(n13361), .ZN(n13525) );
  NAND2_X1 U8816 ( .A1(n9322), .A2(n9321), .ZN(n9448) );
  NAND2_X1 U8817 ( .A1(n8079), .A2(n7616), .ZN(n9384) );
  NAND2_X1 U8818 ( .A1(n12292), .A2(n13504), .ZN(n8079) );
  NAND2_X1 U8819 ( .A1(n9304), .A2(n9303), .ZN(n13470) );
  NAND2_X1 U8820 ( .A1(n9284), .A2(n9283), .ZN(n13942) );
  INV_X1 U8821 ( .A(n16711), .ZN(n16652) );
  INV_X1 U8822 ( .A(n14899), .ZN(n10318) );
  NAND2_X1 U8823 ( .A1(n9402), .A2(n9401), .ZN(n8739) );
  AOI21_X1 U8824 ( .B1(n8589), .B2(n9333), .A(n8585), .ZN(n8584) );
  INV_X1 U8825 ( .A(n8587), .ZN(n8585) );
  AOI21_X1 U8826 ( .B1(n8589), .B2(n13492), .A(n8588), .ZN(n8587) );
  INV_X1 U8827 ( .A(n13498), .ZN(n8588) );
  NAND2_X1 U8828 ( .A1(n12927), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n8592) );
  AND2_X1 U8829 ( .A1(n8747), .A2(n8372), .ZN(n8371) );
  INV_X1 U8830 ( .A(n8885), .ZN(n8372) );
  AOI21_X1 U8831 ( .B1(n8597), .B2(n8596), .A(n8595), .ZN(n9320) );
  AND2_X1 U8832 ( .A1(n16125), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n8595) );
  NAND2_X1 U8833 ( .A1(n8168), .A2(n8171), .ZN(n9397) );
  AND2_X1 U8834 ( .A1(n8169), .A2(n8747), .ZN(n8168) );
  AND2_X1 U8835 ( .A1(n7462), .A2(n8170), .ZN(n8169) );
  INV_X1 U8836 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n8170) );
  AOI21_X1 U8837 ( .B1(n9302), .B2(P1_DATAO_REG_24__SCAN_IN), .A(n8922), .ZN(
        n8931) );
  XNOR2_X1 U8838 ( .A(n8921), .B(n16134), .ZN(n9302) );
  XNOR2_X1 U8839 ( .A(n9424), .B(n9423), .ZN(n9642) );
  INV_X1 U8840 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n9388) );
  OAI22_X1 U8841 ( .A1(n8573), .A2(n8572), .B1(P1_DATAO_REG_21__SCAN_IN), .B2(
        n12796), .ZN(n9282) );
  INV_X1 U8842 ( .A(n9270), .ZN(n8572) );
  NAND2_X1 U8843 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n8040), .ZN(n8039) );
  NOR2_X1 U8844 ( .A1(n8172), .A2(n8173), .ZN(n9229) );
  INV_X1 U8845 ( .A(n7462), .ZN(n8172) );
  AOI21_X1 U8846 ( .B1(n8569), .B2(n8571), .A(n7609), .ZN(n8567) );
  OR2_X1 U8847 ( .A1(n9051), .A2(P3_IR_REG_7__SCAN_IN), .ZN(n9097) );
  AOI21_X1 U8848 ( .B1(n7838), .B2(n7840), .A(n7553), .ZN(n7836) );
  NAND2_X1 U8849 ( .A1(n8044), .A2(n8876), .ZN(n9032) );
  AND2_X1 U8850 ( .A1(n8044), .A2(n8744), .ZN(n9048) );
  AND2_X1 U8851 ( .A1(n8876), .A2(n8745), .ZN(n8744) );
  XNOR2_X1 U8852 ( .A(n8985), .B(P3_IR_REG_2__SCAN_IN), .ZN(n9671) );
  OR2_X1 U8853 ( .A1(n9668), .A2(n9077), .ZN(n8985) );
  XNOR2_X1 U8854 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(P1_DATAO_REG_1__SCAN_IN), 
        .ZN(n8964) );
  AND2_X1 U8855 ( .A1(n9710), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n8973) );
  NAND2_X1 U8856 ( .A1(n15477), .A2(n8849), .ZN(n8266) );
  INV_X1 U8857 ( .A(n11090), .ZN(n7919) );
  NAND2_X1 U8858 ( .A1(n10841), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n12179) );
  INV_X1 U8859 ( .A(n12079), .ZN(n10841) );
  AND2_X1 U8860 ( .A1(n13013), .A2(n10984), .ZN(n10460) );
  OR2_X1 U8861 ( .A1(n12179), .A2(n12178), .ZN(n12198) );
  NAND2_X1 U8862 ( .A1(n7734), .A2(n13304), .ZN(n13346) );
  NAND2_X1 U8863 ( .A1(n8024), .A2(n7521), .ZN(n7734) );
  INV_X1 U8864 ( .A(n9786), .ZN(n13262) );
  OR2_X1 U8865 ( .A1(n10449), .A2(P2_IR_REG_13__SCAN_IN), .ZN(n10630) );
  INV_X1 U8866 ( .A(n7863), .ZN(n7862) );
  OAI21_X1 U8867 ( .B1(n8690), .B2(n7474), .A(n7873), .ZN(n15205) );
  OAI21_X1 U8868 ( .B1(n7474), .B2(n7877), .A(n8695), .ZN(n7874) );
  NAND2_X1 U8869 ( .A1(n15224), .A2(n15135), .ZN(n15210) );
  AND2_X1 U8870 ( .A1(n8323), .A2(n8322), .ZN(n15246) );
  NAND2_X1 U8871 ( .A1(n15246), .A2(n15228), .ZN(n15227) );
  NAND2_X1 U8872 ( .A1(n8325), .A2(n8324), .ZN(n15274) );
  INV_X1 U8873 ( .A(n15424), .ZN(n8324) );
  NAND2_X1 U8874 ( .A1(n15316), .A2(n15123), .ZN(n15300) );
  OR2_X1 U8875 ( .A1(n12454), .A2(n12453), .ZN(n12608) );
  NAND2_X1 U8876 ( .A1(n15338), .A2(n7524), .ZN(n15322) );
  NOR2_X1 U8877 ( .A1(n15355), .A2(n15329), .ZN(n15328) );
  NOR2_X1 U8878 ( .A1(n7490), .A2(n8709), .ZN(n8708) );
  NOR2_X1 U8879 ( .A1(n8710), .A2(n12492), .ZN(n8709) );
  NAND2_X1 U8880 ( .A1(n8328), .A2(n8327), .ZN(n12589) );
  OR2_X1 U8881 ( .A1(n12067), .A2(n12066), .ZN(n12079) );
  OR2_X1 U8882 ( .A1(n16741), .A2(n12226), .ZN(n12474) );
  NAND2_X1 U8883 ( .A1(n7879), .A2(n8701), .ZN(n12218) );
  NAND2_X1 U8884 ( .A1(n12136), .A2(n12135), .ZN(n12217) );
  NAND2_X1 U8885 ( .A1(n8320), .A2(n8319), .ZN(n12226) );
  OR2_X1 U8886 ( .A1(n11369), .A2(n11368), .ZN(n11768) );
  INV_X1 U8887 ( .A(n8320), .ZN(n12143) );
  NAND2_X1 U8888 ( .A1(n8707), .A2(n8706), .ZN(n12136) );
  INV_X1 U8889 ( .A(n11765), .ZN(n8707) );
  INV_X1 U8890 ( .A(n11729), .ZN(n8033) );
  NAND2_X1 U8891 ( .A1(n11723), .A2(n11732), .ZN(n11777) );
  NAND2_X1 U8892 ( .A1(n11638), .A2(n11385), .ZN(n11590) );
  NAND2_X1 U8893 ( .A1(n11642), .A2(n16639), .ZN(n11641) );
  NAND2_X1 U8894 ( .A1(n7864), .A2(n7866), .ZN(n11267) );
  NAND2_X1 U8895 ( .A1(n10537), .A2(n11284), .ZN(n10522) );
  XNOR2_X1 U8896 ( .A(n8111), .B(n10581), .ZN(n10539) );
  INV_X1 U8897 ( .A(n10539), .ZN(n13311) );
  NOR2_X1 U8898 ( .A1(n10538), .A2(n13035), .ZN(n10537) );
  NAND2_X1 U8899 ( .A1(n7627), .A2(n8321), .ZN(n10538) );
  INV_X1 U8900 ( .A(n10460), .ZN(n10545) );
  NOR2_X1 U8901 ( .A1(n13342), .A2(n8082), .ZN(n10232) );
  NAND2_X1 U8902 ( .A1(n11062), .A2(n7439), .ZN(n8318) );
  NAND2_X1 U8903 ( .A1(n7969), .A2(n7968), .ZN(n15318) );
  NAND2_X1 U8904 ( .A1(n12499), .A2(n8751), .ZN(n7969) );
  AOI21_X1 U8905 ( .B1(n8751), .B2(n8753), .A(n7465), .ZN(n7968) );
  NAND2_X1 U8906 ( .A1(n7978), .A2(n8776), .ZN(n12467) );
  NAND2_X1 U8907 ( .A1(n7983), .A2(n7981), .ZN(n7978) );
  INV_X1 U8908 ( .A(n11062), .ZN(n12596) );
  CLKBUF_X1 U8909 ( .A(n13011), .Z(n16704) );
  INV_X1 U8910 ( .A(n16678), .ZN(n16740) );
  NOR2_X1 U8911 ( .A1(n11245), .A2(n10225), .ZN(n10240) );
  AND2_X1 U8912 ( .A1(n10076), .A2(n9818), .ZN(n16148) );
  NAND2_X1 U8913 ( .A1(n7858), .A2(n7856), .ZN(n9713) );
  AND2_X1 U8914 ( .A1(n7859), .A2(n7857), .ZN(n7856) );
  INV_X1 U8915 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n9581) );
  OR2_X1 U8916 ( .A1(n9944), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n9946) );
  OR2_X1 U8917 ( .A1(n9946), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n9979) );
  NOR2_X1 U8918 ( .A1(n9910), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n10148) );
  OR2_X1 U8919 ( .A1(n9890), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n9910) );
  INV_X1 U8920 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n9759) );
  INV_X1 U8921 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n9710) );
  AND2_X1 U8922 ( .A1(n8831), .A2(n7800), .ZN(n7799) );
  INV_X1 U8923 ( .A(n12530), .ZN(n7800) );
  NAND2_X1 U8924 ( .A1(n12848), .A2(n12847), .ZN(n15557) );
  NAND2_X1 U8925 ( .A1(n15557), .A2(n12853), .ZN(n15613) );
  INV_X1 U8926 ( .A(n10270), .ZN(n7768) );
  NAND2_X1 U8927 ( .A1(n10274), .A2(n8067), .ZN(n10354) );
  INV_X1 U8928 ( .A(n8068), .ZN(n8067) );
  OAI21_X1 U8929 ( .B1(n12940), .B2(n15990), .A(n10273), .ZN(n8068) );
  NAND2_X1 U8930 ( .A1(n12381), .A2(n12382), .ZN(n8836) );
  NAND2_X1 U8931 ( .A1(n12377), .A2(n8834), .ZN(n8837) );
  AOI22_X1 U8932 ( .A1(n12128), .A2(n12127), .B1(n11985), .B2(n11984), .ZN(
        n11986) );
  NAND2_X1 U8933 ( .A1(n15645), .A2(n15646), .ZN(n15644) );
  OR2_X1 U8934 ( .A1(n12308), .A2(n12307), .ZN(n12351) );
  AND4_X1 U8935 ( .A1(n10721), .A2(n10720), .A3(n10719), .A4(n10718), .ZN(
        n13684) );
  INV_X2 U8936 ( .A(n7420), .ZN(n12929) );
  NAND2_X1 U8937 ( .A1(n12945), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n10701) );
  AOI21_X1 U8938 ( .B1(P1_REG1_REG_4__SCAN_IN), .B2(n10041), .A(n10290), .ZN(
        n10063) );
  AOI21_X1 U8939 ( .B1(P1_REG1_REG_10__SCAN_IN), .B2(n11559), .A(n10755), .ZN(
        n10757) );
  XNOR2_X1 U8940 ( .A(n15718), .B(n15717), .ZN(n15712) );
  NOR2_X1 U8941 ( .A1(n15708), .A2(n8020), .ZN(n15718) );
  AND2_X1 U8942 ( .A1(n15709), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n8020) );
  NOR2_X1 U8943 ( .A1(n15808), .A2(n15791), .ZN(n15781) );
  AOI21_X1 U8944 ( .B1(n8616), .B2(n8615), .A(n7425), .ZN(n8614) );
  NAND2_X1 U8945 ( .A1(n8000), .A2(n8405), .ZN(n7998) );
  NAND2_X1 U8946 ( .A1(n15838), .A2(n15971), .ZN(n8558) );
  NAND2_X1 U8947 ( .A1(n15829), .A2(n15828), .ZN(n8617) );
  NAND2_X1 U8948 ( .A1(n15842), .A2(n15764), .ZN(n15829) );
  OR2_X1 U8949 ( .A1(n15869), .A2(n15778), .ZN(n8538) );
  INV_X1 U8950 ( .A(n8843), .ZN(n8634) );
  AND2_X1 U8951 ( .A1(n16040), .A2(n15777), .ZN(n8539) );
  NAND2_X1 U8952 ( .A1(n7680), .A2(n7995), .ZN(n15857) );
  NOR2_X1 U8953 ( .A1(n15762), .A2(n8539), .ZN(n7995) );
  INV_X1 U8954 ( .A(n7680), .ZN(n15883) );
  NAND2_X1 U8955 ( .A1(n7466), .A2(n15884), .ZN(n15876) );
  NAND2_X1 U8956 ( .A1(n8308), .A2(n8311), .ZN(n15936) );
  NAND2_X1 U8957 ( .A1(n12556), .A2(n8601), .ZN(n8600) );
  INV_X1 U8958 ( .A(n8604), .ZN(n8601) );
  NAND2_X1 U8959 ( .A1(n12556), .A2(n13592), .ZN(n8602) );
  INV_X1 U8960 ( .A(n8310), .ZN(n15977) );
  NOR2_X1 U8961 ( .A1(n12556), .A2(n8529), .ZN(n8530) );
  INV_X1 U8962 ( .A(n8532), .ZN(n8529) );
  INV_X1 U8963 ( .A(n12556), .ZN(n13595) );
  NOR2_X1 U8964 ( .A1(n13728), .A2(n7729), .ZN(n7727) );
  INV_X1 U8965 ( .A(n11909), .ZN(n7728) );
  NOR2_X1 U8966 ( .A1(n11909), .A2(n7729), .ZN(n12095) );
  NOR2_X1 U8967 ( .A1(n11909), .A2(n13715), .ZN(n11872) );
  NAND2_X1 U8968 ( .A1(n11750), .A2(n11543), .ZN(n11913) );
  NAND2_X1 U8969 ( .A1(n8629), .A2(n8628), .ZN(n8627) );
  INV_X1 U8970 ( .A(n16607), .ZN(n8628) );
  NOR2_X1 U8971 ( .A1(n11349), .A2(n16607), .ZN(n11748) );
  OR2_X1 U8972 ( .A1(n11440), .A2(n13689), .ZN(n11349) );
  NAND2_X1 U8973 ( .A1(n8542), .A2(n8544), .ZN(n11446) );
  OR2_X1 U8974 ( .A1(n11147), .A2(n8545), .ZN(n8542) );
  NAND2_X1 U8975 ( .A1(n8298), .A2(n16572), .ZN(n11440) );
  INV_X1 U8976 ( .A(n11439), .ZN(n8298) );
  XNOR2_X1 U8977 ( .A(n15689), .B(n16554), .ZN(n13675) );
  NAND2_X1 U8978 ( .A1(n7458), .A2(n10934), .ZN(n10940) );
  AND2_X1 U8979 ( .A1(n7458), .A2(n7732), .ZN(n10950) );
  INV_X1 U8980 ( .A(n10932), .ZN(n13575) );
  INV_X1 U8981 ( .A(n15738), .ZN(n16027) );
  INV_X1 U8982 ( .A(n15906), .ZN(n16053) );
  NAND2_X1 U8983 ( .A1(n7479), .A2(n8549), .ZN(n15928) );
  NAND2_X1 U8984 ( .A1(n8549), .A2(n15770), .ZN(n15926) );
  NAND2_X1 U8985 ( .A1(n12728), .A2(n11544), .ZN(n12730) );
  INV_X1 U8986 ( .A(n16606), .ZN(n16725) );
  NAND2_X1 U8987 ( .A1(n12653), .A2(n8672), .ZN(n8671) );
  NOR2_X1 U8988 ( .A1(n8673), .A2(n13245), .ZN(n8672) );
  INV_X1 U8989 ( .A(n8674), .ZN(n8673) );
  AOI21_X1 U8990 ( .B1(n8670), .B2(n8674), .A(n8669), .ZN(n8668) );
  NOR2_X1 U8991 ( .A1(n13244), .A2(n14910), .ZN(n8669) );
  NOR2_X1 U8992 ( .A1(n8678), .A2(n13245), .ZN(n8670) );
  OAI21_X1 U8993 ( .B1(n12653), .B2(n12652), .A(n12642), .ZN(n13216) );
  XNOR2_X1 U8994 ( .A(n9562), .B(P1_IR_REG_26__SCAN_IN), .ZN(n10380) );
  NAND2_X1 U8995 ( .A1(n8390), .A2(n12633), .ZN(n12892) );
  NAND2_X1 U8996 ( .A1(n7464), .A2(n12629), .ZN(n8390) );
  NAND2_X1 U8997 ( .A1(n9570), .A2(n9569), .ZN(n10389) );
  XNOR2_X1 U8998 ( .A(n9988), .B(P1_IR_REG_21__SCAN_IN), .ZN(n13608) );
  NAND2_X1 U8999 ( .A1(n9553), .A2(n9552), .ZN(n10245) );
  NAND2_X1 U9000 ( .A1(n8684), .A2(n11882), .ZN(n12152) );
  OR2_X1 U9001 ( .A1(n11166), .A2(P1_IR_REG_16__SCAN_IN), .ZN(n11744) );
  NAND2_X1 U9002 ( .A1(n8398), .A2(n10215), .ZN(n10448) );
  NAND2_X1 U9003 ( .A1(n10214), .A2(n8856), .ZN(n8398) );
  NAND2_X1 U9004 ( .A1(n8664), .A2(n10003), .ZN(n10136) );
  NAND2_X1 U9005 ( .A1(n7992), .A2(n9940), .ZN(n9955) );
  NAND2_X1 U9006 ( .A1(n9938), .A2(n9937), .ZN(n7992) );
  NAND2_X1 U9007 ( .A1(n8389), .A2(n9873), .ZN(n9897) );
  NAND2_X1 U9008 ( .A1(n9870), .A2(n9888), .ZN(n8389) );
  INV_X1 U9009 ( .A(n9870), .ZN(n9889) );
  XNOR2_X1 U9010 ( .A(n9867), .B(SI_3_), .ZN(n9869) );
  AND2_X1 U9011 ( .A1(n7661), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n16270) );
  INV_X1 U9012 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n7661) );
  INV_X1 U9013 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n16274) );
  XNOR2_X1 U9014 ( .A(n16273), .B(n7660), .ZN(n16271) );
  INV_X1 U9015 ( .A(n16270), .ZN(n7660) );
  INV_X1 U9016 ( .A(n8526), .ZN(n16273) );
  XNOR2_X1 U9017 ( .A(n7648), .B(P1_ADDR_REG_4__SCAN_IN), .ZN(n16296) );
  INV_X1 U9018 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n16306) );
  AOI22_X1 U9019 ( .A1(n16308), .A2(n16307), .B1(P1_ADDR_REG_5__SCAN_IN), .B2(
        n16306), .ZN(n16313) );
  OR2_X1 U9020 ( .A1(n16306), .A2(P1_ADDR_REG_5__SCAN_IN), .ZN(n16307) );
  INV_X1 U9021 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n16311) );
  INV_X1 U9022 ( .A(n16322), .ZN(n8510) );
  INV_X1 U9023 ( .A(n16323), .ZN(n8511) );
  OAI22_X1 U9024 ( .A1(n16335), .A2(n16336), .B1(P1_ADDR_REG_9__SCAN_IN), .B2(
        n16439), .ZN(n16345) );
  NOR2_X1 U9025 ( .A1(n7647), .A2(n7646), .ZN(n16378) );
  AND2_X1 U9026 ( .A1(n16375), .A2(P3_ADDR_REG_14__SCAN_IN), .ZN(n7646) );
  NOR2_X1 U9027 ( .A1(n16374), .A2(n16373), .ZN(n7647) );
  NAND2_X1 U9028 ( .A1(n7903), .A2(n7905), .ZN(n7902) );
  NAND2_X1 U9029 ( .A1(n7889), .A2(n7893), .ZN(n13834) );
  NAND2_X1 U9030 ( .A1(n8734), .A2(n13914), .ZN(n13843) );
  NAND2_X1 U9031 ( .A1(n9295), .A2(n9294), .ZN(n13847) );
  INV_X1 U9032 ( .A(n12415), .ZN(n8086) );
  NAND2_X1 U9033 ( .A1(n11334), .A2(n8732), .ZN(n11420) );
  NAND2_X1 U9034 ( .A1(n8928), .A2(n8927), .ZN(n14392) );
  NAND2_X1 U9035 ( .A1(n11839), .A2(n8037), .ZN(n11969) );
  INV_X1 U9036 ( .A(n11408), .ZN(n11530) );
  NAND2_X1 U9037 ( .A1(n13923), .A2(n9495), .ZN(n13868) );
  NAND2_X1 U9038 ( .A1(n12574), .A2(n8727), .ZN(n13876) );
  NAND2_X1 U9039 ( .A1(n7599), .A2(n14380), .ZN(n8727) );
  AND4_X1 U9040 ( .A1(n8955), .A2(n8954), .A3(n8953), .A4(n8952), .ZN(n14313)
         );
  OAI21_X1 U9041 ( .B1(n8730), .B2(n8731), .A(n8729), .ZN(n11504) );
  INV_X1 U9042 ( .A(n8731), .ZN(n8085) );
  AND2_X1 U9043 ( .A1(n9457), .A2(n16496), .ZN(n8731) );
  NAND2_X1 U9044 ( .A1(n11967), .A2(n7886), .ZN(n12298) );
  AND3_X1 U9045 ( .A1(n9085), .A2(n9084), .A3(n9083), .ZN(n16651) );
  NAND2_X1 U9046 ( .A1(n13925), .A2(n13924), .ZN(n13923) );
  NAND2_X1 U9047 ( .A1(n8726), .A2(n8725), .ZN(n13933) );
  AND2_X1 U9048 ( .A1(n9280), .A2(n9279), .ZN(n14265) );
  INV_X1 U9049 ( .A(n13406), .ZN(n12577) );
  NAND2_X1 U9050 ( .A1(n12576), .A2(n12575), .ZN(n12574) );
  NAND2_X1 U9051 ( .A1(n9536), .A2(n9534), .ZN(n13947) );
  AND2_X1 U9052 ( .A1(n8724), .A2(n7501), .ZN(n11681) );
  NAND2_X1 U9053 ( .A1(n8723), .A2(n8724), .ZN(n11679) );
  AND4_X1 U9054 ( .A1(n9223), .A2(n9222), .A3(n9221), .A4(n9220), .ZN(n14311)
         );
  NAND2_X1 U9055 ( .A1(n7888), .A2(n7530), .ZN(n13975) );
  AND2_X1 U9056 ( .A1(n13976), .A2(n13973), .ZN(n8092) );
  AND2_X1 U9057 ( .A1(n9522), .A2(n11012), .ZN(n16451) );
  AND2_X1 U9058 ( .A1(n13519), .A2(n13518), .ZN(n8124) );
  OAI21_X1 U9059 ( .B1(n13553), .B2(n13550), .A(n8042), .ZN(n8041) );
  NAND2_X1 U9060 ( .A1(n13551), .A2(n8738), .ZN(n8042) );
  INV_X1 U9061 ( .A(n14184), .ZN(n13821) );
  INV_X1 U9062 ( .A(n11925), .ZN(n10554) );
  NAND2_X1 U9063 ( .A1(n7808), .A2(n9649), .ZN(n10892) );
  NAND2_X1 U9064 ( .A1(n10898), .A2(n9650), .ZN(n7808) );
  NAND2_X1 U9065 ( .A1(n10889), .A2(n9669), .ZN(n11218) );
  INV_X1 U9066 ( .A(n7818), .ZN(n10906) );
  OR2_X1 U9067 ( .A1(n11513), .A2(n11514), .ZN(n11511) );
  OAI21_X1 U9068 ( .B1(n10903), .B2(n10899), .A(n10900), .ZN(n11513) );
  OAI21_X1 U9069 ( .B1(n11518), .B2(n7693), .A(n7692), .ZN(n11605) );
  NAND2_X1 U9070 ( .A1(n7694), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n7693) );
  NAND2_X1 U9071 ( .A1(n9678), .A2(n7694), .ZN(n7692) );
  INV_X1 U9072 ( .A(n11606), .ZN(n7694) );
  INV_X1 U9073 ( .A(P3_ADDR_REG_9__SCAN_IN), .ZN(n16439) );
  INV_X1 U9074 ( .A(n16150), .ZN(n16438) );
  NAND2_X1 U9075 ( .A1(n8417), .A2(n9681), .ZN(n16422) );
  NOR2_X1 U9076 ( .A1(n16425), .A2(n8178), .ZN(n11951) );
  NOR2_X1 U9077 ( .A1(n11951), .A2(n11950), .ZN(n11949) );
  NAND2_X1 U9078 ( .A1(n12158), .A2(n12157), .ZN(n12156) );
  NAND2_X1 U9079 ( .A1(n11952), .A2(n9635), .ZN(n12158) );
  INV_X1 U9080 ( .A(n7813), .ZN(n12154) );
  NAND2_X1 U9081 ( .A1(n7737), .A2(n7738), .ZN(n9639) );
  AND2_X1 U9082 ( .A1(n13988), .A2(n13987), .ZN(n13990) );
  INV_X1 U9083 ( .A(n8432), .ZN(n14015) );
  NAND2_X1 U9084 ( .A1(n8436), .A2(n8437), .ZN(n8857) );
  OAI21_X1 U9085 ( .B1(n7841), .B2(n14108), .A(n14101), .ZN(n14081) );
  NOR2_X1 U9086 ( .A1(n7911), .A2(n7910), .ZN(n7909) );
  NAND2_X1 U9087 ( .A1(n7913), .A2(n16501), .ZN(n7912) );
  NOR2_X1 U9088 ( .A1(n14209), .A2(n14312), .ZN(n7910) );
  NAND2_X1 U9089 ( .A1(n8342), .A2(n8346), .ZN(n14185) );
  NAND2_X1 U9090 ( .A1(n8341), .A2(n8348), .ZN(n8342) );
  AOI21_X1 U9091 ( .B1(n8341), .B2(n14205), .A(n13484), .ZN(n14199) );
  INV_X1 U9092 ( .A(n8158), .ZN(n12568) );
  NAND2_X1 U9093 ( .A1(n16648), .A2(n13403), .ZN(n12280) );
  OR2_X1 U9094 ( .A1(n12049), .A2(n13395), .ZN(n16648) );
  AND3_X1 U9095 ( .A1(n9102), .A2(n9101), .A3(n9100), .ZN(n16614) );
  NAND2_X1 U9096 ( .A1(n8340), .A2(n13379), .ZN(n12245) );
  NAND2_X1 U9097 ( .A1(n11920), .A2(n13526), .ZN(n8340) );
  AND3_X1 U9098 ( .A1(n9019), .A2(n9018), .A3(n9017), .ZN(n11836) );
  INV_X1 U9099 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n14474) );
  NAND2_X1 U9100 ( .A1(n16491), .A2(n13368), .ZN(n11815) );
  NAND2_X1 U9101 ( .A1(n8990), .A2(n8989), .ZN(n11816) );
  NAND2_X1 U9102 ( .A1(n11012), .A2(n11011), .ZN(n16508) );
  INV_X1 U9103 ( .A(n16508), .ZN(n14369) );
  NAND2_X1 U9104 ( .A1(n8136), .A2(n8139), .ZN(n14174) );
  AND2_X1 U9105 ( .A1(n13506), .A2(n13505), .ZN(n14840) );
  INV_X1 U9106 ( .A(n13510), .ZN(n14843) );
  NAND3_X1 U9107 ( .A1(n8128), .A2(n8126), .A3(n8127), .ZN(n9442) );
  NOR2_X1 U9108 ( .A1(n7438), .A2(n9358), .ZN(n8127) );
  INV_X1 U9109 ( .A(n9448), .ZN(n14850) );
  OR2_X1 U9110 ( .A1(n13557), .A2(n13550), .ZN(n16615) );
  INV_X1 U9111 ( .A(n9384), .ZN(n14854) );
  INV_X1 U9112 ( .A(n13470), .ZN(n14861) );
  INV_X1 U9113 ( .A(n13847), .ZN(n14865) );
  INV_X1 U9114 ( .A(n13942), .ZN(n14869) );
  AOI21_X1 U9115 ( .B1(n10675), .B2(n13504), .A(n9248), .ZN(n14881) );
  OR2_X1 U9116 ( .A1(n14436), .A2(n14435), .ZN(n14882) );
  NAND2_X1 U9117 ( .A1(n9234), .A2(n9233), .ZN(n14886) );
  INV_X1 U9118 ( .A(n8739), .ZN(n14900) );
  AND2_X1 U9119 ( .A1(n9642), .A2(P3_STATE_REG_SCAN_IN), .ZN(n14899) );
  INV_X1 U9120 ( .A(SI_30_), .ZN(n14910) );
  NAND2_X1 U9121 ( .A1(n8586), .A2(n8589), .ZN(n13497) );
  OR2_X1 U9122 ( .A1(n8593), .A2(n13492), .ZN(n8586) );
  INV_X1 U9123 ( .A(SI_29_), .ZN(n14914) );
  INV_X1 U9124 ( .A(SI_28_), .ZN(n14919) );
  NAND2_X1 U9125 ( .A1(n9394), .A2(n9395), .ZN(n11935) );
  MUX2_X1 U9126 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9393), .S(
        P3_IR_REG_25__SCAN_IN), .Z(n9394) );
  INV_X1 U9127 ( .A(SI_25_), .ZN(n14656) );
  NAND3_X1 U9128 ( .A1(n8089), .A2(n9392), .A3(n8090), .ZN(n13831) );
  NAND2_X1 U9129 ( .A1(n8091), .A2(n9077), .ZN(n8090) );
  OR2_X1 U9130 ( .A1(n9391), .A2(n8091), .ZN(n8089) );
  INV_X1 U9131 ( .A(SI_23_), .ZN(n12618) );
  XNOR2_X1 U9132 ( .A(n9345), .B(P3_IR_REG_22__SCAN_IN), .ZN(n13557) );
  NAND2_X1 U9133 ( .A1(n9348), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9345) );
  INV_X1 U9134 ( .A(n8573), .ZN(n9271) );
  XNOR2_X1 U9135 ( .A(n9350), .B(n8749), .ZN(n10787) );
  INV_X1 U9136 ( .A(SI_19_), .ZN(n14666) );
  INV_X1 U9137 ( .A(SI_17_), .ZN(n11162) );
  NAND2_X1 U9138 ( .A1(n7822), .A2(n8914), .ZN(n9209) );
  NAND2_X1 U9139 ( .A1(n9189), .A2(n9188), .ZN(n7822) );
  INV_X1 U9140 ( .A(SI_15_), .ZN(n10621) );
  INV_X1 U9141 ( .A(SI_14_), .ZN(n14647) );
  NAND2_X1 U9142 ( .A1(n9164), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n8565) );
  INV_X1 U9143 ( .A(SI_12_), .ZN(n14676) );
  INV_X1 U9144 ( .A(SI_11_), .ZN(n14679) );
  NAND2_X1 U9145 ( .A1(n8568), .A2(n8909), .ZN(n9136) );
  NAND2_X1 U9146 ( .A1(n9120), .A2(n9118), .ZN(n8568) );
  XNOR2_X1 U9147 ( .A(n9064), .B(P3_IR_REG_7__SCAN_IN), .ZN(n11524) );
  NAND2_X1 U9148 ( .A1(n7837), .A2(n8903), .ZN(n9031) );
  NAND2_X1 U9149 ( .A1(n9014), .A2(n9012), .ZN(n7837) );
  AND2_X1 U9150 ( .A1(n7416), .A2(P3_U3151), .ZN(n9852) );
  OR2_X1 U9151 ( .A1(n8412), .A2(n9668), .ZN(n10898) );
  NAND2_X1 U9152 ( .A1(n11135), .A2(n9769), .ZN(n9823) );
  INV_X1 U9153 ( .A(n12602), .ZN(n8293) );
  NAND2_X1 U9154 ( .A1(n12603), .A2(n12604), .ZN(n8294) );
  NAND2_X1 U9155 ( .A1(n8288), .A2(n12676), .ZN(n12682) );
  NAND2_X1 U9156 ( .A1(n11184), .A2(n11061), .ZN(n8288) );
  NOR2_X1 U9157 ( .A1(n12176), .A2(n7933), .ZN(n7932) );
  INV_X1 U9158 ( .A(n12172), .ZN(n7933) );
  CLKBUF_X1 U9159 ( .A(n15146), .Z(n8008) );
  AND2_X1 U9160 ( .A1(n12656), .A2(n8287), .ZN(n8283) );
  OR2_X1 U9161 ( .A1(n12676), .A2(n7483), .ZN(n8287) );
  NAND2_X1 U9162 ( .A1(n10460), .A2(n14937), .ZN(n10982) );
  NAND2_X1 U9163 ( .A1(n12709), .A2(n11796), .ZN(n11797) );
  INV_X1 U9164 ( .A(n8270), .ZN(n8269) );
  INV_X1 U9165 ( .A(n15032), .ZN(n12137) );
  NAND2_X1 U9166 ( .A1(n8282), .A2(n11365), .ZN(n12706) );
  NAND2_X1 U9167 ( .A1(n11361), .A2(n11360), .ZN(n8282) );
  NAND2_X1 U9168 ( .A1(n8499), .A2(n8501), .ZN(n10661) );
  INV_X1 U9169 ( .A(n15037), .ZN(n13064) );
  NAND4_X1 U9170 ( .A1(n9764), .A2(n9763), .A3(n9762), .A4(n9761), .ZN(n15042)
         );
  OR2_X2 U9171 ( .A1(n10076), .A2(n9588), .ZN(n15044) );
  NAND2_X1 U9172 ( .A1(n8313), .A2(n7436), .ZN(n15377) );
  NAND2_X1 U9173 ( .A1(n15198), .A2(n8315), .ZN(n15118) );
  AND2_X1 U9174 ( .A1(n15240), .A2(n15133), .ZN(n15226) );
  NAND2_X1 U9175 ( .A1(n8698), .A2(n15160), .ZN(n15221) );
  NAND2_X1 U9176 ( .A1(n15236), .A2(n15239), .ZN(n8698) );
  NAND2_X1 U9177 ( .A1(n8690), .A2(n15156), .ZN(n15251) );
  NAND2_X1 U9178 ( .A1(n7975), .A2(n15128), .ZN(n15255) );
  NAND2_X1 U9179 ( .A1(n7872), .A2(n15152), .ZN(n15283) );
  NAND2_X1 U9180 ( .A1(n8755), .A2(n8754), .ZN(n15349) );
  NAND2_X1 U9181 ( .A1(n12588), .A2(n12587), .ZN(n15122) );
  NAND2_X1 U9182 ( .A1(n12493), .A2(n12492), .ZN(n12585) );
  NAND2_X1 U9183 ( .A1(n12224), .A2(n8779), .ZN(n12466) );
  AND2_X1 U9184 ( .A1(n12224), .A2(n12223), .ZN(n12225) );
  NAND2_X1 U9185 ( .A1(n11719), .A2(n11718), .ZN(n11721) );
  NAND2_X1 U9186 ( .A1(n11383), .A2(n11382), .ZN(n11640) );
  NAND2_X1 U9187 ( .A1(n11239), .A2(n11238), .ZN(n11241) );
  NAND2_X1 U9188 ( .A1(n7869), .A2(n10486), .ZN(n11249) );
  NAND2_X1 U9189 ( .A1(n10523), .A2(n10484), .ZN(n7869) );
  NAND2_X1 U9190 ( .A1(n10519), .A2(n10467), .ZN(n11236) );
  INV_X1 U9191 ( .A(n15330), .ZN(n15367) );
  AND2_X1 U9192 ( .A1(n15353), .A2(n13338), .ZN(n15371) );
  NAND2_X1 U9193 ( .A1(n15353), .A2(n11280), .ZN(n15359) );
  NOR2_X1 U9194 ( .A1(n15385), .A2(n8715), .ZN(n8714) );
  AND2_X1 U9195 ( .A1(n15386), .A2(n16740), .ZN(n8715) );
  INV_X1 U9196 ( .A(n15195), .ZN(n15481) );
  INV_X1 U9197 ( .A(n15211), .ZN(n15485) );
  INV_X1 U9198 ( .A(n15304), .ZN(n15500) );
  INV_X1 U9199 ( .A(n13113), .ZN(n15518) );
  INV_X1 U9200 ( .A(n13024), .ZN(n11294) );
  AND2_X2 U9201 ( .A1(n10240), .A2(n10239), .ZN(n16751) );
  INV_X1 U9202 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n9702) );
  NOR2_X1 U9203 ( .A1(n7416), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15528) );
  NOR2_X1 U9204 ( .A1(n10990), .A2(n8694), .ZN(n9714) );
  XNOR2_X1 U9205 ( .A(n9584), .B(n9699), .ZN(n15534) );
  NAND2_X1 U9206 ( .A1(n9583), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9584) );
  XNOR2_X1 U9207 ( .A(n9585), .B(n9697), .ZN(n15536) );
  INV_X1 U9208 ( .A(n9807), .ZN(n15539) );
  AND2_X1 U9209 ( .A1(n7416), .A2(P2_U3088), .ZN(n15542) );
  INV_X1 U9210 ( .A(n13342), .ZN(n12371) );
  AOI21_X1 U9211 ( .B1(n9731), .B2(n9726), .A(n9715), .ZN(n9727) );
  INV_X1 U9212 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n11889) );
  INV_X1 U9213 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n10015) );
  INV_X1 U9214 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n9928) );
  INV_X1 U9215 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n9914) );
  AOI21_X1 U9216 ( .B1(n11022), .B2(n11021), .A(n8825), .ZN(n11691) );
  NAND2_X1 U9217 ( .A1(n7801), .A2(n8831), .ZN(n12529) );
  NAND2_X1 U9218 ( .A1(n15644), .A2(n12757), .ZN(n15568) );
  NAND2_X1 U9219 ( .A1(n11022), .A2(n8823), .ZN(n8820) );
  NAND2_X1 U9220 ( .A1(n12377), .A2(n8838), .ZN(n12402) );
  NAND2_X1 U9221 ( .A1(n15612), .A2(n12874), .ZN(n15584) );
  NAND2_X1 U9222 ( .A1(n12717), .A2(n8855), .ZN(n15592) );
  INV_X1 U9223 ( .A(n7769), .ZN(n10810) );
  OAI211_X1 U9224 ( .C1(n7775), .C2(n7772), .A(n7770), .B(n7773), .ZN(n7769)
         );
  INV_X1 U9225 ( .A(n7771), .ZN(n7770) );
  NAND2_X1 U9226 ( .A1(n7773), .A2(n7774), .ZN(n10729) );
  NAND2_X1 U9227 ( .A1(n7781), .A2(n8816), .ZN(n11700) );
  NAND2_X1 U9228 ( .A1(n11022), .A2(n7437), .ZN(n7781) );
  NAND2_X1 U9229 ( .A1(n11700), .A2(n11699), .ZN(n11976) );
  OAI21_X1 U9230 ( .B1(n10354), .B2(n7767), .A(n10353), .ZN(n12649) );
  NAND2_X1 U9231 ( .A1(n7556), .A2(n7788), .ZN(n7787) );
  NAND2_X1 U9232 ( .A1(n7463), .A2(n7790), .ZN(n7788) );
  NAND2_X1 U9233 ( .A1(n8815), .A2(n15565), .ZN(n15627) );
  OAI21_X1 U9234 ( .B1(n15645), .B2(n7790), .A(n7463), .ZN(n8815) );
  AND2_X1 U9235 ( .A1(n8837), .A2(n8836), .ZN(n12527) );
  NAND2_X1 U9236 ( .A1(n15574), .A2(n12812), .ZN(n15633) );
  NAND2_X1 U9237 ( .A1(n15574), .A2(n7428), .ZN(n15634) );
  INV_X1 U9238 ( .A(n12853), .ZN(n7796) );
  AND2_X1 U9239 ( .A1(n13651), .A2(n7571), .ZN(n13802) );
  NOR2_X1 U9240 ( .A1(n8654), .A2(n8854), .ZN(n8070) );
  NAND2_X1 U9241 ( .A1(n10402), .A2(n10401), .ZN(n15951) );
  OR2_X1 U9242 ( .A1(n10392), .A2(n9571), .ZN(n15677) );
  INV_X1 U9243 ( .A(n13684), .ZN(n15688) );
  NAND2_X1 U9244 ( .A1(n7420), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n10421) );
  NAND2_X1 U9245 ( .A1(n8019), .A2(n8018), .ZN(n15697) );
  OR2_X1 U9246 ( .A1(n10364), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n8019) );
  NAND2_X1 U9247 ( .A1(n10364), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n8018) );
  NAND2_X1 U9248 ( .A1(n15697), .A2(n15696), .ZN(n15695) );
  AOI21_X1 U9249 ( .B1(P1_REG1_REG_2__SCAN_IN), .B2(n10283), .A(n10021), .ZN(
        n10024) );
  AOI21_X1 U9250 ( .B1(n10812), .B2(P1_REG1_REG_6__SCAN_IN), .A(n10155), .ZN(
        n10157) );
  NOR2_X1 U9251 ( .A1(n11468), .A2(n11469), .ZN(n11890) );
  NAND2_X1 U9252 ( .A1(n8303), .A2(n16079), .ZN(n15999) );
  XNOR2_X1 U9253 ( .A(n15746), .B(n8074), .ZN(n8303) );
  NAND2_X1 U9254 ( .A1(n8097), .A2(n8096), .ZN(n8095) );
  NAND2_X1 U9255 ( .A1(n15859), .A2(n15971), .ZN(n8096) );
  NAND2_X1 U9256 ( .A1(n8608), .A2(n8606), .ZN(n15892) );
  AND2_X1 U9257 ( .A1(n8611), .A2(n8610), .ZN(n15901) );
  NAND2_X1 U9258 ( .A1(n12969), .A2(n11544), .ZN(n12781) );
  NAND2_X1 U9259 ( .A1(n15955), .A2(n15769), .ZN(n15932) );
  OR2_X1 U9260 ( .A1(n7414), .A2(n10879), .ZN(n16481) );
  OAI21_X1 U9261 ( .B1(n12555), .B2(n12554), .A(n8604), .ZN(n12557) );
  NAND2_X1 U9262 ( .A1(n8536), .A2(n12343), .ZN(n12346) );
  NAND2_X1 U9263 ( .A1(n8537), .A2(n13593), .ZN(n8536) );
  NAND2_X1 U9264 ( .A1(n12324), .A2(n12323), .ZN(n12326) );
  AND2_X1 U9265 ( .A1(n12019), .A2(n12018), .ZN(n12089) );
  NAND2_X1 U9266 ( .A1(n11869), .A2(n11868), .ZN(n11871) );
  AND2_X1 U9267 ( .A1(n8621), .A2(n8623), .ZN(n11907) );
  AND2_X1 U9268 ( .A1(n8551), .A2(n11538), .ZN(n11752) );
  NAND2_X1 U9269 ( .A1(n11343), .A2(n11342), .ZN(n11537) );
  INV_X1 U9270 ( .A(n16486), .ZN(n16631) );
  NAND2_X1 U9271 ( .A1(n10878), .A2(n10877), .ZN(n16622) );
  NOR2_X1 U9272 ( .A1(n7414), .A2(n16726), .ZN(n15855) );
  NAND2_X1 U9273 ( .A1(n15790), .A2(n16622), .ZN(n16625) );
  INV_X1 U9274 ( .A(n16481), .ZN(n16628) );
  NOR2_X1 U9275 ( .A1(n15790), .A2(n13606), .ZN(n16486) );
  AND2_X2 U9276 ( .A1(n11139), .A2(n10442), .ZN(n16734) );
  NAND2_X1 U9277 ( .A1(n15999), .A2(n8301), .ZN(n16097) );
  INV_X1 U9278 ( .A(n8302), .ZN(n8301) );
  OAI21_X1 U9279 ( .B1(n8074), .B2(n16725), .A(n16000), .ZN(n8302) );
  NAND2_X1 U9280 ( .A1(n16003), .A2(n16730), .ZN(n7733) );
  AOI21_X1 U9281 ( .B1(n16010), .B2(n16730), .A(n8555), .ZN(n8554) );
  NAND2_X1 U9282 ( .A1(n16013), .A2(n16012), .ZN(n8555) );
  NAND2_X1 U9283 ( .A1(n16019), .A2(n7504), .ZN(n16101) );
  AND2_X2 U9284 ( .A1(n11139), .A2(n11138), .ZN(n16737) );
  NOR2_X1 U9285 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_29__SCAN_IN), .ZN(
        n7964) );
  INV_X1 U9286 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n16125) );
  INV_X1 U9287 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n16131) );
  XNOR2_X1 U9288 ( .A(n9564), .B(P1_IR_REG_25__SCAN_IN), .ZN(n16128) );
  NOR2_X1 U9289 ( .A1(n7416), .A2(P1_STATE_REG_SCAN_IN), .ZN(n16135) );
  OR2_X1 U9290 ( .A1(n12829), .A2(n7416), .ZN(n12813) );
  INV_X1 U9291 ( .A(n8639), .ZN(n8638) );
  INV_X1 U9292 ( .A(n13608), .ZN(n15988) );
  INV_X1 U9293 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n12779) );
  INV_X1 U9294 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n11887) );
  INV_X1 U9295 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10644) );
  INV_X1 U9296 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10457) );
  INV_X1 U9297 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n12005) );
  INV_X1 U9298 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n10010) );
  INV_X1 U9299 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n9978) );
  INV_X1 U9300 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n9959) );
  INV_X1 U9301 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n9943) );
  INV_X1 U9302 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n10684) );
  OAI21_X1 U9303 ( .B1(n9874), .B2(n8094), .A(n8093), .ZN(n9739) );
  XNOR2_X1 U9304 ( .A(n9738), .B(n9861), .ZN(n9740) );
  NAND2_X1 U9305 ( .A1(n9874), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n8093) );
  INV_X1 U9306 ( .A(P2_RD_REG_SCAN_IN), .ZN(n8925) );
  NOR2_X1 U9307 ( .A1(n16276), .A2(n16275), .ZN(n16278) );
  XNOR2_X1 U9308 ( .A(n16296), .B(n8521), .ZN(n16298) );
  INV_X1 U9309 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n8521) );
  AND2_X1 U9310 ( .A1(n7659), .A2(n7566), .ZN(n16297) );
  OR2_X1 U9311 ( .A1(n16290), .A2(P2_ADDR_REG_3__SCAN_IN), .ZN(n7659) );
  AOI21_X1 U9312 ( .B1(n16305), .B2(n16304), .A(n16303), .ZN(n16413) );
  XNOR2_X1 U9313 ( .A(n16321), .B(P2_ADDR_REG_7__SCAN_IN), .ZN(n16323) );
  NAND2_X1 U9314 ( .A1(n8519), .A2(n16340), .ZN(n16342) );
  NAND2_X1 U9315 ( .A1(n16339), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n8519) );
  NAND2_X1 U9316 ( .A1(n16342), .A2(n16343), .ZN(n16344) );
  INV_X1 U9317 ( .A(n7665), .ZN(n16363) );
  OAI21_X1 U9318 ( .B1(n16357), .B2(P2_ADDR_REG_12__SCAN_IN), .A(n7517), .ZN(
        n7665) );
  INV_X1 U9319 ( .A(n8518), .ZN(n16356) );
  NAND2_X1 U9320 ( .A1(n16363), .A2(n16362), .ZN(n16364) );
  NAND2_X1 U9321 ( .A1(n8495), .A2(n16364), .ZN(n16371) );
  OAI21_X1 U9322 ( .B1(n16363), .B2(n16362), .A(P2_ADDR_REG_13__SCAN_IN), .ZN(
        n8495) );
  NAND2_X1 U9323 ( .A1(n16371), .A2(n16370), .ZN(n16372) );
  NAND2_X1 U9324 ( .A1(n7657), .A2(n16372), .ZN(n16380) );
  OAI21_X1 U9325 ( .B1(n16371), .B2(n16370), .A(P2_ADDR_REG_14__SCAN_IN), .ZN(
        n7657) );
  INV_X1 U9326 ( .A(n7843), .ZN(n14012) );
  INV_X1 U9327 ( .A(n8188), .ZN(n14080) );
  OAI211_X1 U9328 ( .C1(n14127), .C2(n16429), .A(n7697), .B(n7695), .ZN(
        P3_U3200) );
  AOI21_X1 U9329 ( .B1(n14126), .B2(n14125), .A(n7624), .ZN(n7695) );
  OAI21_X1 U9330 ( .B1(n14121), .B2(n14122), .A(n14120), .ZN(n7697) );
  NAND2_X1 U9331 ( .A1(n8439), .A2(n14120), .ZN(n8438) );
  NOR2_X1 U9332 ( .A1(n14145), .A2(n8442), .ZN(n8441) );
  XNOR2_X1 U9333 ( .A(n8174), .B(n14140), .ZN(n14148) );
  AND3_X1 U9334 ( .A1(n8128), .A2(n8133), .A3(n8126), .ZN(n13814) );
  OAI21_X1 U9335 ( .B1(n14830), .B2(n14829), .A(n14828), .ZN(n14837) );
  OAI21_X1 U9336 ( .B1(n14958), .B2(n8100), .A(n8099), .ZN(P2_U3186) );
  INV_X1 U9337 ( .A(n14948), .ZN(n8099) );
  NAND2_X1 U9338 ( .A1(n8101), .A2(n15000), .ZN(n8100) );
  AOI21_X1 U9339 ( .B1(n8506), .B2(n8261), .A(n7560), .ZN(n8258) );
  NAND2_X1 U9340 ( .A1(n8500), .A2(n11047), .ZN(n11052) );
  NAND2_X1 U9341 ( .A1(n11173), .A2(n10650), .ZN(n8500) );
  OAI211_X1 U9342 ( .C1(n15026), .C2(n15025), .A(n7477), .B(n8017), .ZN(
        P2_U3212) );
  AOI21_X1 U9343 ( .B1(n15211), .B2(n15024), .A(n15023), .ZN(n8017) );
  XNOR2_X1 U9344 ( .A(n7785), .B(n12944), .ZN(n12956) );
  MUX2_X1 U9345 ( .A(n15735), .B(n15734), .S(n15733), .Z(n15737) );
  OAI21_X1 U9346 ( .B1(n8300), .B2(n16735), .A(n8299), .ZN(P1_U3527) );
  NAND2_X1 U9347 ( .A1(n16735), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n8299) );
  INV_X1 U9348 ( .A(n16097), .ZN(n8300) );
  NOR2_X1 U9349 ( .A1(n16389), .A2(n16388), .ZN(n16390) );
  NAND2_X1 U9350 ( .A1(n8515), .A2(n8514), .ZN(n16399) );
  NAND2_X1 U9351 ( .A1(n16389), .A2(n8516), .ZN(n8515) );
  XNOR2_X1 U9352 ( .A(n16410), .B(P3_ADDR_REG_19__SCAN_IN), .ZN(n8528) );
  OAI21_X1 U9353 ( .B1(n16409), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n7653), .ZN(
        n7652) );
  NAND2_X1 U9354 ( .A1(n13759), .A2(n8646), .ZN(n7419) );
  AND2_X2 U9355 ( .A1(n12655), .A2(n10356), .ZN(n7420) );
  INV_X2 U9356 ( .A(n10702), .ZN(n11544) );
  AND3_X1 U9357 ( .A1(n11250), .A2(n10537), .A3(n7568), .ZN(n7421) );
  AND3_X1 U9358 ( .A1(n13747), .A2(n13746), .A3(n7588), .ZN(n7423) );
  AND2_X1 U9359 ( .A1(n14272), .A2(n8153), .ZN(n7424) );
  AND2_X1 U9360 ( .A1(n8618), .A2(n13570), .ZN(n7425) );
  AND2_X1 U9361 ( .A1(n13758), .A2(n13760), .ZN(n7426) );
  AND2_X1 U9362 ( .A1(n13737), .A2(n13739), .ZN(n7427) );
  NAND2_X1 U9363 ( .A1(n8509), .A2(n14929), .ZN(n8505) );
  NAND2_X1 U9364 ( .A1(n16141), .A2(n12814), .ZN(n16046) );
  NAND2_X2 U9365 ( .A1(n7412), .A2(n12329), .ZN(n12846) );
  XNOR2_X1 U9366 ( .A(n7764), .B(P3_IR_REG_27__SCAN_IN), .ZN(n13555) );
  INV_X1 U9367 ( .A(n9847), .ZN(n7686) );
  NOR2_X1 U9368 ( .A1(n13489), .A2(n13509), .ZN(n13520) );
  AND2_X1 U9369 ( .A1(n12824), .A2(n12812), .ZN(n7428) );
  XNOR2_X1 U9370 ( .A(n15043), .B(n13024), .ZN(n13309) );
  XNOR2_X1 U9371 ( .A(n13384), .B(n16580), .ZN(n13532) );
  INV_X1 U9372 ( .A(n13532), .ZN(n8339) );
  INV_X1 U9373 ( .A(n13021), .ZN(n8321) );
  INV_X1 U9374 ( .A(n16586), .ZN(n7669) );
  AND2_X1 U9375 ( .A1(n8603), .A2(n8600), .ZN(n7429) );
  AND2_X1 U9376 ( .A1(n7514), .A2(n8318), .ZN(n7430) );
  AND2_X1 U9377 ( .A1(n8770), .A2(n15130), .ZN(n7431) );
  OAI21_X1 U9378 ( .B1(n8508), .B2(n8509), .A(n8507), .ZN(n8506) );
  NAND2_X1 U9379 ( .A1(n12341), .A2(n12340), .ZN(n16090) );
  OR2_X1 U9380 ( .A1(n12830), .A2(SI_22_), .ZN(n7432) );
  INV_X1 U9381 ( .A(n13546), .ZN(n8358) );
  AND2_X1 U9382 ( .A1(n8761), .A2(n8760), .ZN(n7433) );
  NAND2_X1 U9383 ( .A1(n8742), .A2(n8044), .ZN(n9051) );
  OR2_X1 U9384 ( .A1(n14854), .A2(n14198), .ZN(n7434) );
  INV_X1 U9385 ( .A(n14978), .ZN(n7925) );
  OR2_X1 U9386 ( .A1(n13769), .A2(n13770), .ZN(n7435) );
  NAND2_X1 U9387 ( .A1(n13252), .A2(n13251), .ZN(n15111) );
  INV_X1 U9388 ( .A(n15111), .ZN(n15468) );
  AND3_X1 U9389 ( .A1(n8314), .A2(n14960), .A3(n7670), .ZN(n7436) );
  AND2_X1 U9390 ( .A1(n8823), .A2(n8826), .ZN(n7437) );
  INV_X1 U9391 ( .A(n10934), .ZN(n8046) );
  AND2_X1 U9392 ( .A1(n13812), .A2(n16647), .ZN(n7438) );
  INV_X1 U9393 ( .A(n14173), .ZN(n7851) );
  XNOR2_X1 U9394 ( .A(n15040), .B(n11284), .ZN(n13312) );
  AND2_X1 U9395 ( .A1(n9844), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n7439) );
  XNOR2_X1 U9396 ( .A(n15424), .B(n14959), .ZN(n14923) );
  XNOR2_X1 U9397 ( .A(n10652), .B(n10651), .ZN(n11047) );
  AND3_X1 U9398 ( .A1(n8436), .A2(P3_REG2_REG_15__SCAN_IN), .A3(n8437), .ZN(
        n7440) );
  AND2_X1 U9399 ( .A1(n7561), .A2(n7943), .ZN(n7441) );
  AND2_X1 U9400 ( .A1(n8365), .A2(n8362), .ZN(n7442) );
  INV_X1 U9401 ( .A(n9789), .ZN(n10470) );
  NAND2_X1 U9402 ( .A1(n15884), .A2(n7487), .ZN(n7443) );
  NAND2_X1 U9403 ( .A1(n13565), .A2(n13564), .ZN(n15743) );
  INV_X1 U9404 ( .A(n15743), .ZN(n8074) );
  AND2_X1 U9405 ( .A1(n15485), .A2(n15136), .ZN(n7444) );
  AND2_X1 U9406 ( .A1(n7564), .A2(n7938), .ZN(n7445) );
  INV_X1 U9407 ( .A(n14272), .ZN(n14877) );
  NAND2_X1 U9408 ( .A1(n9263), .A2(n9262), .ZN(n14272) );
  OR2_X1 U9409 ( .A1(n14957), .A2(n14929), .ZN(n8508) );
  INV_X1 U9410 ( .A(n13758), .ZN(n8646) );
  INV_X1 U9411 ( .A(n13737), .ZN(n8645) );
  INV_X1 U9412 ( .A(n13716), .ZN(n8647) );
  INV_X1 U9413 ( .A(n16017), .ZN(n15827) );
  NAND2_X1 U9414 ( .A1(n15812), .A2(n7715), .ZN(n16017) );
  NAND2_X1 U9415 ( .A1(n10679), .A2(n10680), .ZN(n7446) );
  AND2_X1 U9416 ( .A1(n9844), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n7447) );
  NAND2_X1 U9417 ( .A1(n16046), .A2(n15761), .ZN(n7709) );
  INV_X1 U9418 ( .A(n15444), .ZN(n8329) );
  AND2_X1 U9419 ( .A1(n9401), .A2(n8738), .ZN(n7448) );
  AND2_X1 U9420 ( .A1(n12344), .A2(n12323), .ZN(n7449) );
  INV_X1 U9421 ( .A(n8505), .ZN(n8504) );
  INV_X1 U9422 ( .A(n13749), .ZN(n8117) );
  AND2_X1 U9423 ( .A1(n7686), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n7450) );
  AND2_X1 U9424 ( .A1(n13748), .A2(n8117), .ZN(n7451) );
  NAND2_X1 U9425 ( .A1(n13738), .A2(n8645), .ZN(n7452) );
  NAND2_X1 U9426 ( .A1(n13717), .A2(n8647), .ZN(n7453) );
  AND2_X1 U9427 ( .A1(n8387), .A2(n11160), .ZN(n7454) );
  INV_X1 U9428 ( .A(n15838), .ZN(n13570) );
  XNOR2_X1 U9429 ( .A(SI_4_), .B(keyinput_28), .ZN(n7455) );
  NAND2_X1 U9430 ( .A1(n8820), .A2(n8821), .ZN(n11712) );
  AND2_X1 U9431 ( .A1(n9662), .A2(n7813), .ZN(n7456) );
  AND4_X1 U9432 ( .A1(n9131), .A2(n9130), .A3(n9129), .A4(n9128), .ZN(n12419)
         );
  INV_X1 U9433 ( .A(n12419), .ZN(n14380) );
  NAND2_X1 U9434 ( .A1(n8328), .A2(n7667), .ZN(n7668) );
  AND2_X1 U9435 ( .A1(n16388), .A2(P2_ADDR_REG_16__SCAN_IN), .ZN(n8517) );
  INV_X1 U9436 ( .A(n8517), .ZN(n8514) );
  AND2_X1 U9437 ( .A1(n12150), .A2(SI_20_), .ZN(n7457) );
  INV_X1 U9438 ( .A(n13328), .ZN(n8712) );
  INV_X1 U9439 ( .A(n11102), .ZN(n7920) );
  AND2_X1 U9440 ( .A1(n16480), .A2(n15990), .ZN(n7458) );
  AND2_X1 U9441 ( .A1(n14619), .A2(n7634), .ZN(n7459) );
  INV_X1 U9442 ( .A(n7411), .ZN(n9287) );
  INV_X1 U9443 ( .A(n8950), .ZN(n10995) );
  INV_X1 U9444 ( .A(n8979), .ZN(n8950) );
  OR2_X1 U9445 ( .A1(n9718), .A2(P2_IR_REG_22__SCAN_IN), .ZN(n7460) );
  NAND2_X1 U9446 ( .A1(n7855), .A2(n7853), .ZN(n13021) );
  NAND2_X1 U9447 ( .A1(n11530), .A2(n16497), .ZN(n8167) );
  NAND3_X1 U9448 ( .A1(n8692), .A2(n7977), .A3(n8693), .ZN(n7461) );
  INV_X1 U9449 ( .A(n15041), .ZN(n8111) );
  NAND2_X1 U9450 ( .A1(n8984), .A2(n7416), .ZN(n8995) );
  AND2_X1 U9451 ( .A1(n15566), .A2(n7789), .ZN(n7463) );
  NAND2_X1 U9452 ( .A1(n8945), .A2(n8884), .ZN(n9244) );
  AND2_X1 U9453 ( .A1(n12628), .A2(n8023), .ZN(n7464) );
  NOR2_X1 U9454 ( .A1(n15444), .A2(n15319), .ZN(n7465) );
  AND2_X1 U9455 ( .A1(n7705), .A2(n7709), .ZN(n7466) );
  NAND2_X1 U9456 ( .A1(n13395), .A2(n12041), .ZN(n7467) );
  NOR2_X1 U9457 ( .A1(n13013), .A2(n13012), .ZN(n13015) );
  NAND4_X1 U9458 ( .A1(n9709), .A2(n9708), .A3(n9707), .A4(n9706), .ZN(n13013)
         );
  AND4_X1 U9459 ( .A1(n9724), .A2(n8312), .A3(n9700), .A4(n9699), .ZN(n7468)
         );
  OR2_X1 U9460 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n7469) );
  NOR2_X1 U9461 ( .A1(n14167), .A2(n11040), .ZN(n7470) );
  OR2_X1 U9462 ( .A1(n12980), .A2(n12979), .ZN(n7471) );
  NAND2_X1 U9463 ( .A1(n10653), .A2(n10652), .ZN(n7472) );
  INV_X1 U9464 ( .A(n9258), .ZN(n8154) );
  INV_X1 U9465 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n8923) );
  XNOR2_X1 U9466 ( .A(n15869), .B(n15778), .ZN(n15762) );
  INV_X1 U9467 ( .A(n8165), .ZN(n8164) );
  OAI21_X1 U9468 ( .B1(n13537), .B2(n7486), .A(n9154), .ZN(n8165) );
  AND2_X1 U9469 ( .A1(n8741), .A2(n8740), .ZN(n7473) );
  INV_X1 U9470 ( .A(n15184), .ZN(n15477) );
  OR2_X1 U9471 ( .A1(n8697), .A2(n7875), .ZN(n7474) );
  NOR2_X1 U9472 ( .A1(n14082), .A2(n7691), .ZN(n7475) );
  OR2_X1 U9473 ( .A1(n16282), .A2(n16281), .ZN(n7476) );
  INV_X1 U9474 ( .A(n8578), .ZN(n13544) );
  OR2_X1 U9475 ( .A1(n13510), .A2(n13507), .ZN(n8578) );
  OR2_X1 U9476 ( .A1(n15022), .A2(n15021), .ZN(n7477) );
  OR2_X1 U9477 ( .A1(n8431), .A2(n14017), .ZN(n7478) );
  AND2_X1 U9478 ( .A1(n15758), .A2(n15770), .ZN(n7479) );
  INV_X1 U9479 ( .A(n13612), .ZN(n13779) );
  OR2_X1 U9480 ( .A1(n11220), .A2(n9652), .ZN(n7480) );
  XNOR2_X1 U9481 ( .A(n9450), .B(n9449), .ZN(n9453) );
  NOR2_X1 U9482 ( .A1(n9461), .A2(n11842), .ZN(n7481) );
  NAND4_X1 U9483 ( .A1(n10399), .A2(n10400), .A3(n10398), .A4(n10397), .ZN(
        n16463) );
  INV_X1 U9484 ( .A(n16463), .ZN(n8047) );
  NAND2_X1 U9485 ( .A1(n8933), .A2(n8932), .ZN(n9510) );
  INV_X1 U9486 ( .A(n9510), .ZN(n8351) );
  INV_X1 U9487 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n8078) );
  XNOR2_X1 U9488 ( .A(n8886), .B(P3_IR_REG_30__SCAN_IN), .ZN(n8890) );
  NAND2_X1 U9489 ( .A1(n16021), .A2(n15765), .ZN(n7482) );
  AND2_X1 U9490 ( .A1(n12658), .A2(n11077), .ZN(n7483) );
  AND2_X1 U9491 ( .A1(n12703), .A2(n11792), .ZN(n7484) );
  AND2_X1 U9492 ( .A1(n7778), .A2(n10709), .ZN(n7485) );
  NAND2_X1 U9493 ( .A1(n14380), .A2(n12580), .ZN(n7486) );
  INV_X1 U9494 ( .A(n15828), .ZN(n8615) );
  OR2_X1 U9495 ( .A1(n15869), .A2(n15675), .ZN(n7487) );
  AND2_X1 U9496 ( .A1(n7452), .A2(n7948), .ZN(n7488) );
  AND2_X1 U9497 ( .A1(n8569), .A2(n7832), .ZN(n7489) );
  AND2_X1 U9498 ( .A1(n13329), .A2(n15028), .ZN(n7490) );
  INV_X1 U9499 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n7965) );
  AND2_X1 U9500 ( .A1(n7979), .A2(n13328), .ZN(n7491) );
  OR2_X1 U9501 ( .A1(n15477), .A2(n15517), .ZN(n7492) );
  AND4_X1 U9502 ( .A1(n14245), .A2(n14221), .A3(n13543), .A4(n14230), .ZN(
        n7493) );
  AND2_X1 U9503 ( .A1(n15808), .A2(n15791), .ZN(n7494) );
  INV_X1 U9504 ( .A(n11699), .ZN(n7780) );
  AND2_X1 U9505 ( .A1(n14854), .A2(n14198), .ZN(n7495) );
  AND2_X1 U9506 ( .A1(n16627), .A2(n15685), .ZN(n7496) );
  NOR2_X1 U9507 ( .A1(n11246), .A2(n8082), .ZN(n13011) );
  INV_X1 U9508 ( .A(n13781), .ZN(n8659) );
  OR2_X1 U9509 ( .A1(n15848), .A2(n8305), .ZN(n7497) );
  NAND2_X1 U9510 ( .A1(n10733), .A2(n7674), .ZN(n13685) );
  INV_X1 U9511 ( .A(n13685), .ZN(n16572) );
  OR2_X1 U9512 ( .A1(n16349), .A2(n16350), .ZN(n7498) );
  AND2_X1 U9513 ( .A1(n16078), .A2(n15755), .ZN(n7499) );
  OR2_X1 U9514 ( .A1(n14608), .A2(n14607), .ZN(n7500) );
  NAND2_X1 U9515 ( .A1(n9460), .A2(n11829), .ZN(n7501) );
  AND2_X1 U9516 ( .A1(n8423), .A2(n8425), .ZN(n7502) );
  AND2_X1 U9517 ( .A1(n8131), .A2(n16501), .ZN(n7503) );
  AND3_X1 U9518 ( .A1(n8848), .A2(n8859), .A3(n16018), .ZN(n7504) );
  INV_X1 U9519 ( .A(n10709), .ZN(n7777) );
  AND2_X1 U9520 ( .A1(n8747), .A2(n7462), .ZN(n7505) );
  AND2_X1 U9521 ( .A1(n8701), .A2(n7878), .ZN(n7506) );
  AND3_X1 U9522 ( .A1(n8271), .A2(n8270), .A3(n8267), .ZN(n7507) );
  AND2_X1 U9523 ( .A1(n14186), .A2(n8348), .ZN(n7508) );
  AND2_X1 U9524 ( .A1(n13076), .A2(n13075), .ZN(n7509) );
  INV_X1 U9525 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n9716) );
  AND2_X1 U9526 ( .A1(n13098), .A2(n13097), .ZN(n7510) );
  NAND2_X1 U9527 ( .A1(n10138), .A2(n10003), .ZN(n8663) );
  INV_X1 U9528 ( .A(n8735), .ZN(n13914) );
  OAI21_X1 U9529 ( .B1(n13943), .B2(n9502), .A(n8736), .ZN(n8735) );
  NOR2_X1 U9530 ( .A1(n13592), .A2(n8535), .ZN(n8534) );
  INV_X1 U9531 ( .A(n13582), .ZN(n11751) );
  AND2_X1 U9532 ( .A1(n13152), .A2(n13151), .ZN(n7511) );
  OR2_X1 U9533 ( .A1(n9867), .A2(n9866), .ZN(n7512) );
  AND2_X1 U9534 ( .A1(n11250), .A2(n15039), .ZN(n7513) );
  OR2_X1 U9535 ( .A1(n11062), .A2(n10128), .ZN(n7514) );
  AOI21_X1 U9536 ( .B1(n15645), .B2(n7463), .A(n7787), .ZN(n7786) );
  OR2_X1 U9537 ( .A1(n13121), .A2(n8793), .ZN(n7515) );
  OR2_X1 U9538 ( .A1(n15477), .A2(n15464), .ZN(n7516) );
  INV_X1 U9539 ( .A(n8296), .ZN(n15877) );
  NOR2_X1 U9540 ( .A1(n15894), .A2(n16040), .ZN(n8296) );
  OR2_X1 U9541 ( .A1(n16356), .A2(n16355), .ZN(n7517) );
  AND2_X1 U9542 ( .A1(n15857), .A2(n8538), .ZN(n7518) );
  AND2_X1 U9543 ( .A1(n13379), .A2(n13380), .ZN(n13526) );
  INV_X1 U9544 ( .A(n13526), .ZN(n8336) );
  OR2_X1 U9545 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n16272), .ZN(n7519) );
  AND2_X1 U9546 ( .A1(n15131), .A2(n15130), .ZN(n7520) );
  OR2_X1 U9547 ( .A1(n9721), .A2(n9715), .ZN(n9723) );
  INV_X1 U9548 ( .A(n7908), .ZN(n7907) );
  OAI21_X1 U9549 ( .B1(n13965), .B2(n9518), .A(n9520), .ZN(n7908) );
  AND2_X1 U9550 ( .A1(n15780), .A2(n13571), .ZN(n15814) );
  INV_X1 U9551 ( .A(n15814), .ZN(n8405) );
  INV_X1 U9552 ( .A(n15160), .ZN(n8700) );
  INV_X1 U9553 ( .A(n13757), .ZN(n7944) );
  AND2_X1 U9554 ( .A1(n8685), .A2(n13297), .ZN(n7521) );
  OR2_X1 U9555 ( .A1(n12814), .A2(n10364), .ZN(n7522) );
  AND2_X1 U9556 ( .A1(n8855), .A2(n12726), .ZN(n7523) );
  INV_X1 U9557 ( .A(n8307), .ZN(n15830) );
  NOR2_X1 U9558 ( .A1(n15848), .A2(n16021), .ZN(n8307) );
  AND2_X1 U9559 ( .A1(n15324), .A2(n15321), .ZN(n7524) );
  AND2_X1 U9560 ( .A1(n13298), .A2(n13253), .ZN(n7525) );
  AND2_X1 U9561 ( .A1(n9383), .A2(n9382), .ZN(n14205) );
  INV_X1 U9562 ( .A(n14205), .ZN(n8349) );
  AND2_X1 U9563 ( .A1(n14850), .A2(n14184), .ZN(n7526) );
  AND2_X1 U9564 ( .A1(n8578), .A2(n8575), .ZN(n7527) );
  AND2_X1 U9565 ( .A1(n8609), .A2(n15925), .ZN(n7528) );
  AND2_X1 U9566 ( .A1(n12891), .A2(n12890), .ZN(n7529) );
  AND2_X1 U9567 ( .A1(n7890), .A2(n8092), .ZN(n7530) );
  INV_X1 U9568 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n8091) );
  INV_X1 U9569 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n8888) );
  NAND2_X1 U9570 ( .A1(n7756), .A2(n8803), .ZN(n7531) );
  AND2_X1 U9571 ( .A1(n11699), .A2(n7437), .ZN(n7532) );
  AND2_X1 U9572 ( .A1(n13751), .A2(n7939), .ZN(n7533) );
  AND2_X1 U9573 ( .A1(n15876), .A2(n8633), .ZN(n7534) );
  AND2_X1 U9574 ( .A1(n13370), .A2(n13363), .ZN(n13527) );
  INV_X1 U9575 ( .A(n13527), .ZN(n8333) );
  INV_X1 U9576 ( .A(n15511), .ZN(n8327) );
  INV_X1 U9577 ( .A(n15110), .ZN(n15472) );
  NAND2_X1 U9578 ( .A1(n13219), .A2(n13218), .ZN(n15110) );
  NOR2_X1 U9579 ( .A1(n8782), .A2(n8781), .ZN(n7535) );
  NOR2_X1 U9580 ( .A1(n13728), .A2(n15681), .ZN(n7536) );
  NOR2_X1 U9581 ( .A1(n13102), .A2(n12697), .ZN(n7537) );
  NOR2_X1 U9582 ( .A1(n14941), .A2(n14940), .ZN(n7538) );
  AND2_X1 U9583 ( .A1(n13176), .A2(n13175), .ZN(n7539) );
  OR2_X1 U9584 ( .A1(n8753), .A2(n7465), .ZN(n7540) );
  INV_X1 U9585 ( .A(n7723), .ZN(n7722) );
  NAND2_X1 U9586 ( .A1(n8311), .A2(n7724), .ZN(n7723) );
  AND2_X1 U9587 ( .A1(n13769), .A2(n13770), .ZN(n7541) );
  NAND2_X1 U9588 ( .A1(n15168), .A2(n15166), .ZN(n7542) );
  AND2_X1 U9589 ( .A1(n8152), .A2(n8154), .ZN(n7543) );
  NAND4_X1 U9590 ( .A1(n10701), .A2(n10700), .A3(n10699), .A4(n10698), .ZN(
        n15689) );
  NOR2_X1 U9591 ( .A1(n12828), .A2(n12827), .ZN(n7544) );
  OR2_X1 U9592 ( .A1(n9580), .A2(P2_IR_REG_16__SCAN_IN), .ZN(n7545) );
  OR2_X1 U9593 ( .A1(n8792), .A2(n13122), .ZN(n7546) );
  AND2_X1 U9594 ( .A1(n9956), .A2(SI_8_), .ZN(n7547) );
  INV_X1 U9595 ( .A(n7709), .ZN(n7708) );
  INV_X1 U9596 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n9923) );
  NAND2_X1 U9597 ( .A1(n15211), .A2(n15162), .ZN(n7548) );
  INV_X1 U9598 ( .A(n8828), .ZN(n8825) );
  OR2_X1 U9599 ( .A1(n9497), .A2(n8147), .ZN(n7549) );
  NAND2_X1 U9600 ( .A1(n8807), .A2(n13131), .ZN(n7550) );
  NOR2_X1 U9601 ( .A1(n16068), .A2(n15756), .ZN(n7551) );
  AND2_X1 U9602 ( .A1(n10446), .A2(SI_13_), .ZN(n7552) );
  AND2_X1 U9603 ( .A1(n9878), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n7553) );
  AND2_X1 U9604 ( .A1(n8806), .A2(n13134), .ZN(n7554) );
  OR2_X1 U9605 ( .A1(n7533), .A2(n7451), .ZN(n7555) );
  AND2_X1 U9606 ( .A1(n12790), .A2(n15565), .ZN(n7556) );
  NOR2_X1 U9607 ( .A1(n13109), .A2(n8785), .ZN(n7557) );
  INV_X1 U9608 ( .A(n8141), .ZN(n8140) );
  NAND2_X1 U9609 ( .A1(n7434), .A2(n8142), .ZN(n8141) );
  OR2_X1 U9610 ( .A1(n12846), .A2(n10265), .ZN(n7558) );
  AND2_X1 U9611 ( .A1(n8351), .A2(n8350), .ZN(n7559) );
  NAND2_X1 U9612 ( .A1(n14966), .A2(n14967), .ZN(n7560) );
  AND2_X1 U9613 ( .A1(n13757), .A2(n7945), .ZN(n7561) );
  AND2_X1 U9614 ( .A1(n8364), .A2(n8981), .ZN(n7562) );
  NAND2_X1 U9615 ( .A1(n8144), .A2(n13457), .ZN(n7563) );
  NAND2_X1 U9616 ( .A1(n13753), .A2(n8649), .ZN(n7564) );
  INV_X1 U9617 ( .A(n10694), .ZN(n7778) );
  INV_X1 U9618 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n7977) );
  INV_X1 U9619 ( .A(n13752), .ZN(n8649) );
  INV_X1 U9620 ( .A(n13748), .ZN(n8648) );
  XNOR2_X1 U9621 ( .A(n16607), .B(n15686), .ZN(n13580) );
  AND2_X1 U9622 ( .A1(n9015), .A2(n9001), .ZN(n9652) );
  OR2_X1 U9623 ( .A1(n15256), .A2(n15157), .ZN(n7565) );
  OR2_X1 U9624 ( .A1(n16289), .A2(n16288), .ZN(n7566) );
  INV_X1 U9625 ( .A(n13459), .ZN(n7900) );
  AND2_X1 U9626 ( .A1(n7903), .A2(n7908), .ZN(n7567) );
  AND2_X1 U9627 ( .A1(n11284), .A2(n7669), .ZN(n7568) );
  NOR2_X1 U9628 ( .A1(n16008), .A2(n16007), .ZN(n7569) );
  AND2_X1 U9629 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n16271), .ZN(n7570) );
  AND2_X1 U9630 ( .A1(n13650), .A2(n8072), .ZN(n7571) );
  AND2_X1 U9631 ( .A1(n8504), .A2(n8261), .ZN(n7572) );
  AND2_X1 U9632 ( .A1(n9503), .A2(n9504), .ZN(n7573) );
  XNOR2_X1 U9633 ( .A(n9453), .B(n10517), .ZN(n11331) );
  AND2_X1 U9634 ( .A1(n9103), .A2(n9040), .ZN(n7574) );
  AND2_X1 U9635 ( .A1(n7830), .A2(n8567), .ZN(n7575) );
  INV_X1 U9636 ( .A(n8406), .ZN(n15804) );
  OR2_X1 U9637 ( .A1(n7494), .A2(n15781), .ZN(n8406) );
  INV_X1 U9638 ( .A(n13734), .ZN(n7949) );
  AND2_X1 U9639 ( .A1(n13521), .A2(n7527), .ZN(n7576) );
  AND2_X1 U9640 ( .A1(n8337), .A2(n13385), .ZN(n7577) );
  OR2_X1 U9641 ( .A1(n8659), .A2(n13780), .ZN(n7578) );
  OR2_X1 U9642 ( .A1(n8784), .A2(n13110), .ZN(n7579) );
  OR2_X1 U9643 ( .A1(n13141), .A2(n13142), .ZN(n7580) );
  AND2_X1 U9644 ( .A1(n8333), .A2(n8989), .ZN(n7581) );
  AND2_X1 U9645 ( .A1(n7862), .A2(n7542), .ZN(n7582) );
  OR2_X1 U9646 ( .A1(n13520), .A2(n7470), .ZN(n7583) );
  AND2_X1 U9647 ( .A1(n8373), .A2(n8888), .ZN(n7584) );
  INV_X1 U9648 ( .A(n7714), .ZN(n7713) );
  NAND2_X1 U9649 ( .A1(n12088), .A2(n12018), .ZN(n7714) );
  AND2_X1 U9650 ( .A1(n7473), .A2(n8091), .ZN(n7585) );
  AND2_X1 U9651 ( .A1(n16059), .A2(n15759), .ZN(n15760) );
  NAND2_X1 U9652 ( .A1(n13713), .A2(n7963), .ZN(n7586) );
  NAND2_X1 U9653 ( .A1(n13730), .A2(n8650), .ZN(n7587) );
  NAND2_X1 U9654 ( .A1(n13749), .A2(n8648), .ZN(n7588) );
  AND2_X1 U9655 ( .A1(n8405), .A2(n7482), .ZN(n8616) );
  AND2_X1 U9656 ( .A1(n7453), .A2(n7962), .ZN(n7589) );
  NAND2_X1 U9657 ( .A1(n9898), .A2(SI_5_), .ZN(n7590) );
  OR2_X1 U9658 ( .A1(n8796), .A2(n7539), .ZN(n7591) );
  INV_X1 U9659 ( .A(n14923), .ZN(n8274) );
  OR2_X1 U9660 ( .A1(n8804), .A2(n7510), .ZN(n7592) );
  INV_X1 U9661 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n9579) );
  OR2_X1 U9662 ( .A1(n16059), .A2(n15939), .ZN(n15771) );
  INV_X1 U9663 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n8740) );
  INV_X2 U9664 ( .A(n15327), .ZN(n15362) );
  AND4_X1 U9665 ( .A1(n9269), .A2(n9268), .A3(n9267), .A4(n9266), .ZN(n14278)
         );
  INV_X1 U9666 ( .A(n14278), .ZN(n8153) );
  NAND2_X1 U9667 ( .A1(n12133), .A2(n13324), .ZN(n7983) );
  INV_X1 U9668 ( .A(n14379), .ZN(n8160) );
  INV_X1 U9669 ( .A(n9855), .ZN(n7816) );
  AND2_X1 U9670 ( .A1(n9552), .A2(n8644), .ZN(n7593) );
  NAND2_X1 U9671 ( .A1(n11986), .A2(n11987), .ZN(n12377) );
  INV_X1 U9672 ( .A(n15342), .ZN(n8760) );
  AND2_X1 U9673 ( .A1(n14433), .A2(n14313), .ZN(n7594) );
  INV_X1 U9674 ( .A(n9630), .ZN(n16428) );
  XNOR2_X1 U9675 ( .A(n15414), .B(n15132), .ZN(n15239) );
  AND2_X1 U9676 ( .A1(n13082), .A2(n13081), .ZN(n7595) );
  INV_X1 U9677 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n8830) );
  XNOR2_X1 U9678 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(P2_DATAO_REG_9__SCAN_IN), 
        .ZN(n9075) );
  INV_X1 U9679 ( .A(n9075), .ZN(n7833) );
  INV_X1 U9680 ( .A(n15819), .ZN(n8618) );
  INV_X1 U9681 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n8749) );
  AND2_X1 U9682 ( .A1(n9637), .A2(n12166), .ZN(n7596) );
  NAND2_X1 U9683 ( .A1(n12019), .A2(n7713), .ZN(n12087) );
  XNOR2_X1 U9684 ( .A(SI_5_), .B(keyinput_27), .ZN(n7597) );
  AND3_X1 U9685 ( .A1(n14514), .A2(n14513), .A3(n14512), .ZN(n7598) );
  INV_X1 U9686 ( .A(n8308), .ZN(n15961) );
  NOR2_X1 U9687 ( .A1(n15975), .A2(n16074), .ZN(n8308) );
  AND4_X1 U9688 ( .A1(n9145), .A2(n9144), .A3(n9143), .A4(n9142), .ZN(n13934)
         );
  XOR2_X1 U9689 ( .A(n9516), .B(n12580), .Z(n7599) );
  INV_X1 U9690 ( .A(n8328), .ZN(n12501) );
  NOR2_X1 U9691 ( .A1(n12474), .A2(n13113), .ZN(n8328) );
  AND2_X1 U9692 ( .A1(n8939), .A2(n8938), .ZN(n14209) );
  INV_X1 U9693 ( .A(n14209), .ZN(n8350) );
  AND4_X1 U9694 ( .A1(n9094), .A2(n9093), .A3(n9092), .A4(n9091), .ZN(n12300)
         );
  INV_X1 U9695 ( .A(n12300), .ZN(n13396) );
  OR2_X1 U9696 ( .A1(n13810), .A2(n14455), .ZN(n7600) );
  AND2_X1 U9697 ( .A1(n12556), .A2(n8598), .ZN(n7601) );
  AND2_X1 U9698 ( .A1(n7983), .A2(n12134), .ZN(n7602) );
  AND2_X1 U9699 ( .A1(n8531), .A2(n8532), .ZN(n7603) );
  NAND2_X1 U9700 ( .A1(n12236), .A2(n12235), .ZN(n7604) );
  NAND2_X1 U9701 ( .A1(n9881), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n7605) );
  INV_X1 U9702 ( .A(n12420), .ZN(n12287) );
  AND4_X1 U9703 ( .A1(n9074), .A2(n9073), .A3(n9072), .A4(n9071), .ZN(n12420)
         );
  INV_X1 U9704 ( .A(n8325), .ZN(n15290) );
  NOR2_X1 U9705 ( .A1(n15311), .A2(n15291), .ZN(n8325) );
  INV_X1 U9706 ( .A(n9358), .ZN(n8133) );
  INV_X1 U9707 ( .A(n15414), .ZN(n8322) );
  AND2_X1 U9708 ( .A1(n11592), .A2(n11591), .ZN(n7606) );
  AND2_X1 U9709 ( .A1(n8536), .A2(n8534), .ZN(n7607) );
  INV_X1 U9710 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n8009) );
  INV_X1 U9711 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n8522) );
  INV_X1 U9712 ( .A(n8292), .ZN(n14998) );
  NAND2_X1 U9713 ( .A1(n8294), .A2(n8293), .ZN(n8292) );
  INV_X1 U9714 ( .A(n8757), .ZN(n8756) );
  INV_X1 U9715 ( .A(n11159), .ZN(n8661) );
  OR2_X1 U9716 ( .A1(n8385), .A2(n11160), .ZN(n7608) );
  INV_X1 U9717 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n9878) );
  AND2_X1 U9718 ( .A1(n10010), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n7609) );
  NAND2_X1 U9719 ( .A1(n12470), .A2(n12469), .ZN(n12471) );
  INV_X1 U9720 ( .A(n12471), .ZN(n8713) );
  AND2_X1 U9721 ( .A1(n8915), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n7610) );
  INV_X1 U9722 ( .A(n13729), .ZN(n8650) );
  INV_X1 U9723 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n10153) );
  AND2_X1 U9724 ( .A1(n15753), .A2(n15752), .ZN(n7611) );
  INV_X1 U9725 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n10221) );
  INV_X1 U9726 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n8040) );
  INV_X2 U9727 ( .A(n16719), .ZN(n14891) );
  INV_X1 U9728 ( .A(n13324), .ZN(n8706) );
  INV_X1 U9729 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n8120) );
  INV_X1 U9730 ( .A(n15146), .ZN(n8761) );
  INV_X1 U9731 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n8582) );
  INV_X1 U9732 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7827) );
  AOI21_X1 U9733 ( .B1(n10810), .B2(n10809), .A(n10808), .ZN(n11022) );
  NAND2_X2 U9734 ( .A1(n11014), .A2(n16508), .ZN(n14352) );
  INV_X1 U9735 ( .A(n13583), .ZN(n8620) );
  INV_X1 U9736 ( .A(n13102), .ZN(n8319) );
  INV_X1 U9737 ( .A(n16078), .ZN(n8309) );
  NAND2_X1 U9738 ( .A1(n9682), .A2(n16428), .ZN(n9681) );
  NOR2_X1 U9739 ( .A1(n10704), .A2(n12927), .ZN(n7612) );
  NAND2_X1 U9740 ( .A1(n12762), .A2(n12761), .ZN(n16068) );
  INV_X1 U9741 ( .A(n16068), .ZN(n8311) );
  XOR2_X1 U9742 ( .A(n12634), .B(SI_26_), .Z(n7613) );
  NAND2_X1 U9743 ( .A1(n12009), .A2(n12008), .ZN(n16722) );
  INV_X1 U9744 ( .A(n16722), .ZN(n7730) );
  AND2_X1 U9745 ( .A1(n15000), .A2(n14937), .ZN(n14961) );
  XOR2_X1 U9746 ( .A(n12832), .B(SI_23_), .Z(n7614) );
  AND2_X1 U9747 ( .A1(n14516), .A2(n14515), .ZN(n7615) );
  INV_X1 U9748 ( .A(n8678), .ZN(n8677) );
  AOI21_X1 U9749 ( .B1(n12652), .B2(n12642), .A(n8679), .ZN(n8678) );
  INV_X1 U9750 ( .A(SI_16_), .ZN(n11160) );
  INV_X1 U9751 ( .A(SI_20_), .ZN(n14664) );
  OR2_X1 U9752 ( .A1(n9335), .A2(n14483), .ZN(n7616) );
  NAND2_X1 U9753 ( .A1(n14046), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n7617) );
  AND2_X1 U9754 ( .A1(n16648), .A2(n8369), .ZN(n7618) );
  AND2_X1 U9755 ( .A1(n8626), .A2(n8624), .ZN(n7619) );
  AND2_X1 U9756 ( .A1(n12634), .A2(SI_26_), .ZN(n7620) );
  AND2_X1 U9757 ( .A1(n8820), .A2(n8818), .ZN(n7621) );
  NAND2_X1 U9758 ( .A1(n11869), .A2(n8635), .ZN(n12019) );
  NAND2_X1 U9759 ( .A1(n14063), .A2(n8435), .ZN(n7622) );
  NAND2_X1 U9760 ( .A1(n9389), .A2(n9388), .ZN(n7623) );
  OR2_X1 U9761 ( .A1(n14124), .A2(n7696), .ZN(n7624) );
  INV_X1 U9762 ( .A(SI_18_), .ZN(n14492) );
  OR2_X1 U9763 ( .A1(P3_STATE_REG_SCAN_IN), .A2(keyinput_34), .ZN(n7625) );
  INV_X1 U9764 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n11329) );
  INV_X1 U9765 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n11743) );
  AND2_X1 U9766 ( .A1(n7776), .A2(n7446), .ZN(n7626) );
  INV_X1 U9767 ( .A(n8623), .ZN(n8622) );
  AOI21_X1 U9768 ( .B1(n8624), .B2(n13580), .A(n7496), .ZN(n8623) );
  INV_X1 U9769 ( .A(n11538), .ZN(n8552) );
  OR2_X1 U9770 ( .A1(n9589), .A2(n10318), .ZN(n10989) );
  NAND2_X1 U9771 ( .A1(n9425), .A2(n11012), .ZN(n16719) );
  AND3_X1 U9772 ( .A1(n7430), .A2(n13012), .A3(n9741), .ZN(n7627) );
  NAND2_X1 U9773 ( .A1(n13557), .A2(n13357), .ZN(n13491) );
  NAND2_X1 U9774 ( .A1(n9417), .A2(n13517), .ZN(n16501) );
  INV_X1 U9775 ( .A(n9312), .ZN(n8596) );
  NAND2_X1 U9776 ( .A1(n10647), .A2(n10646), .ZN(n11173) );
  INV_X1 U9777 ( .A(n11173), .ZN(n8496) );
  NOR2_X1 U9778 ( .A1(n10921), .A2(n8852), .ZN(n7628) );
  NOR2_X1 U9779 ( .A1(n11517), .A2(n9678), .ZN(n7629) );
  NAND2_X1 U9780 ( .A1(n14083), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n7630) );
  AND2_X1 U9781 ( .A1(n7775), .A2(n7485), .ZN(n7631) );
  NOR2_X1 U9782 ( .A1(n10704), .A2(n16121), .ZN(n7632) );
  INV_X1 U9783 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n13493) );
  NAND2_X1 U9784 ( .A1(n16131), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n7633) );
  INV_X1 U9785 ( .A(n13549), .ZN(n8738) );
  INV_X1 U9786 ( .A(n9824), .ZN(n13338) );
  INV_X1 U9787 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n8435) );
  NAND2_X1 U9788 ( .A1(n10388), .A2(n10387), .ZN(n16561) );
  AND2_X1 U9789 ( .A1(n8451), .A2(n8450), .ZN(n7634) );
  AND2_X1 U9790 ( .A1(n8409), .A2(n9669), .ZN(n7635) );
  INV_X1 U9791 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n8094) );
  INV_X1 U9792 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n7637) );
  INV_X1 U9793 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n8426) );
  INV_X1 U9794 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n7644) );
  INV_X1 U9795 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n8363) );
  NOR2_X1 U9796 ( .A1(n7416), .A2(P3_STATE_REG_SCAN_IN), .ZN(n14901) );
  INV_X1 U9797 ( .A(n7641), .ZN(n16284) );
  NAND2_X1 U9798 ( .A1(n8525), .A2(n8526), .ZN(n7642) );
  NAND3_X1 U9799 ( .A1(n8513), .A2(n16400), .A3(n7650), .ZN(n7649) );
  XNOR2_X1 U9800 ( .A(n7652), .B(n8528), .ZN(SUB_1596_U4) );
  OAI21_X1 U9801 ( .B1(n16333), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n7664), .ZN(
        n7663) );
  INV_X1 U9802 ( .A(n16334), .ZN(n7664) );
  AND2_X1 U9803 ( .A1(n16325), .A2(n16326), .ZN(n16333) );
  AOI21_X1 U9804 ( .B1(n8511), .B2(n8510), .A(n16324), .ZN(n16325) );
  AOI21_X1 U9805 ( .B1(n16416), .B2(n16417), .A(n7570), .ZN(n16276) );
  NAND3_X1 U9806 ( .A1(n8328), .A2(n7667), .A3(n8329), .ZN(n15355) );
  INV_X1 U9807 ( .A(n7668), .ZN(n8326) );
  NAND3_X1 U9808 ( .A1(n11250), .A2(n10537), .A3(n11284), .ZN(n11274) );
  NAND3_X1 U9809 ( .A1(n15198), .A2(n15468), .A3(n8315), .ZN(n7670) );
  NOR2_X2 U9810 ( .A1(n11596), .A2(n13083), .ZN(n11723) );
  NAND3_X1 U9811 ( .A1(n9578), .A2(n10147), .A3(n9884), .ZN(n10990) );
  MUX2_X1 U9812 ( .A(n10130), .B(n15546), .S(n11062), .Z(n13012) );
  NAND2_X1 U9813 ( .A1(n12315), .A2(n13590), .ZN(n12317) );
  NAND2_X1 U9814 ( .A1(n12090), .A2(n13588), .ZN(n7672) );
  NAND2_X1 U9815 ( .A1(n11848), .A2(n11847), .ZN(n11850) );
  NAND2_X1 U9816 ( .A1(n11913), .A2(n11556), .ZN(n7673) );
  AND2_X2 U9817 ( .A1(n15857), .A2(n7994), .ZN(n15845) );
  NAND3_X1 U9818 ( .A1(n7681), .A2(n8021), .A3(n15771), .ZN(n15911) );
  NOR2_X2 U9819 ( .A1(n15957), .A2(n15958), .ZN(n15956) );
  OAI21_X1 U9820 ( .B1(n11193), .B2(n11192), .A(n11191), .ZN(n11195) );
  AOI21_X1 U9821 ( .B1(n11192), .B2(n11191), .A(n7450), .ZN(n7682) );
  NAND2_X1 U9822 ( .A1(n11193), .A2(n11191), .ZN(n7683) );
  NAND3_X1 U9823 ( .A1(n9681), .A2(n8417), .A3(P3_REG2_REG_9__SCAN_IN), .ZN(
        n8418) );
  NAND2_X1 U9824 ( .A1(n9668), .A2(n8875), .ZN(n8998) );
  NOR2_X4 U9825 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .ZN(
        n9668) );
  OAI21_X1 U9826 ( .B1(n7702), .B2(n7700), .A(n10949), .ZN(n11142) );
  NAND2_X1 U9827 ( .A1(n7701), .A2(n10935), .ZN(n10948) );
  NAND2_X1 U9828 ( .A1(n10933), .A2(n10932), .ZN(n7701) );
  INV_X1 U9829 ( .A(n10935), .ZN(n7703) );
  NAND2_X1 U9830 ( .A1(n7710), .A2(n7711), .ZN(n12021) );
  NAND2_X1 U9831 ( .A1(n12555), .A2(n7429), .ZN(n7717) );
  NAND3_X1 U9832 ( .A1(n7717), .A2(n7718), .A3(n15958), .ZN(n15949) );
  AOI22_X1 U9833 ( .A1(n15949), .A2(n15973), .B1(n15948), .B2(n16074), .ZN(
        n15934) );
  OAI21_X1 U9834 ( .B1(n12555), .B2(n8602), .A(n7429), .ZN(n15982) );
  NAND3_X1 U9835 ( .A1(n10247), .A2(n8839), .A3(n7965), .ZN(n7720) );
  AND2_X2 U9836 ( .A1(n7807), .A2(n9875), .ZN(n10247) );
  XNOR2_X1 U9837 ( .A(n9740), .B(n9739), .ZN(n9893) );
  INV_X1 U9838 ( .A(n7725), .ZN(n15904) );
  INV_X1 U9839 ( .A(n16046), .ZN(n7726) );
  NAND3_X1 U9840 ( .A1(n7732), .A2(n7458), .A3(n13677), .ZN(n11439) );
  NAND3_X1 U9841 ( .A1(n7733), .A2(n8110), .A3(n7569), .ZN(n16099) );
  XNOR2_X1 U9842 ( .A(n14062), .B(n14063), .ZN(n14051) );
  NAND2_X1 U9843 ( .A1(n14027), .A2(n14026), .ZN(n14029) );
  INV_X2 U9844 ( .A(n13302), .ZN(n13160) );
  NAND2_X1 U9845 ( .A1(n7737), .A2(n7735), .ZN(n13988) );
  OR2_X1 U9846 ( .A1(n13085), .A2(n7743), .ZN(n7741) );
  NAND2_X1 U9847 ( .A1(n7741), .A2(n7742), .ZN(n13092) );
  INV_X1 U9848 ( .A(n13092), .ZN(n13095) );
  AND2_X1 U9849 ( .A1(n7745), .A2(n7744), .ZN(n13067) );
  NAND2_X1 U9850 ( .A1(n7749), .A2(n7752), .ZN(n8783) );
  NAND2_X1 U9851 ( .A1(n8802), .A2(n7750), .ZN(n7749) );
  INV_X1 U9852 ( .A(n13104), .ZN(n7756) );
  NAND4_X1 U9853 ( .A1(n9578), .A2(n10147), .A3(n9884), .A4(n9579), .ZN(n11327) );
  NAND2_X1 U9854 ( .A1(n13128), .A2(n7762), .ZN(n7759) );
  NAND3_X1 U9855 ( .A1(n7759), .A2(n7760), .A3(n7758), .ZN(n8780) );
  NOR2_X1 U9856 ( .A1(n7535), .A2(n7761), .ZN(n7760) );
  NAND4_X1 U9857 ( .A1(n7763), .A2(n8091), .A3(n8740), .A4(n9423), .ZN(n8750)
         );
  NAND2_X1 U9858 ( .A1(n7558), .A2(n7768), .ZN(n7767) );
  NAND2_X1 U9859 ( .A1(n10682), .A2(n10681), .ZN(n7776) );
  OAI21_X1 U9860 ( .B1(n7485), .B2(n7772), .A(n7774), .ZN(n7771) );
  NAND2_X1 U9861 ( .A1(n12913), .A2(n15656), .ZN(n15549) );
  INV_X1 U9862 ( .A(n7786), .ZN(n15626) );
  NAND2_X1 U9863 ( .A1(n12848), .A2(n7794), .ZN(n7791) );
  NAND2_X1 U9864 ( .A1(n7791), .A2(n7792), .ZN(n15654) );
  NAND2_X1 U9865 ( .A1(n15576), .A2(n7428), .ZN(n7798) );
  NOR2_X1 U9866 ( .A1(n8833), .A2(n12526), .ZN(n7802) );
  NOR2_X1 U9867 ( .A1(n9550), .A2(n9551), .ZN(n7807) );
  NAND3_X1 U9868 ( .A1(n7806), .A2(n7804), .A3(n7803), .ZN(n9554) );
  NAND2_X1 U9869 ( .A1(n8181), .A2(n8179), .ZN(n16426) );
  INV_X1 U9870 ( .A(n9668), .ZN(n8411) );
  INV_X1 U9871 ( .A(n8412), .ZN(n8410) );
  NAND2_X1 U9872 ( .A1(n7812), .A2(n9662), .ZN(n7813) );
  NAND2_X1 U9873 ( .A1(n9662), .A2(n8192), .ZN(n12155) );
  NAND2_X1 U9874 ( .A1(n9189), .A2(n7823), .ZN(n7820) );
  NAND2_X1 U9875 ( .A1(n7820), .A2(n7821), .ZN(n9226) );
  NAND2_X1 U9876 ( .A1(n9076), .A2(n7489), .ZN(n7829) );
  NAND2_X1 U9877 ( .A1(n7829), .A2(n7575), .ZN(n9148) );
  NAND2_X1 U9878 ( .A1(n9014), .A2(n7838), .ZN(n7835) );
  NAND2_X1 U9879 ( .A1(n7835), .A2(n7836), .ZN(n9055) );
  NAND2_X1 U9880 ( .A1(n7846), .A2(n14056), .ZN(n14038) );
  NAND2_X1 U9881 ( .A1(n8175), .A2(n14063), .ZN(n7846) );
  NOR2_X1 U9882 ( .A1(n11515), .A2(n9658), .ZN(n11614) );
  OAI21_X1 U9883 ( .B1(n11062), .B2(n15045), .A(n7852), .ZN(n7854) );
  NAND2_X1 U9884 ( .A1(n11062), .A2(n7447), .ZN(n7852) );
  XNOR2_X1 U9885 ( .A(n9757), .B(n9756), .ZN(n10408) );
  NAND3_X1 U9886 ( .A1(n8692), .A2(n8693), .A3(P2_IR_REG_28__SCAN_IN), .ZN(
        n7858) );
  NAND2_X1 U9887 ( .A1(n15178), .A2(n7582), .ZN(n7860) );
  OAI211_X1 U9888 ( .C1(n15178), .C2(n7861), .A(n7860), .B(n15174), .ZN(n15384) );
  INV_X1 U9889 ( .A(n10523), .ZN(n7865) );
  INV_X1 U9890 ( .A(n10486), .ZN(n7868) );
  NAND3_X1 U9891 ( .A1(n7864), .A2(n7866), .A3(n13315), .ZN(n11269) );
  NAND2_X1 U9892 ( .A1(n7872), .A2(n7870), .ZN(n15281) );
  INV_X1 U9893 ( .A(n7874), .ZN(n7873) );
  NAND2_X1 U9894 ( .A1(n7882), .A2(n11661), .ZN(n8719) );
  AOI21_X1 U9895 ( .B1(n7882), .B2(n8722), .A(n8718), .ZN(n8717) );
  NAND2_X1 U9896 ( .A1(n8720), .A2(n7882), .ZN(n11841) );
  NAND2_X1 U9897 ( .A1(n11967), .A2(n7884), .ZN(n12296) );
  NAND2_X1 U9898 ( .A1(n7887), .A2(n8726), .ZN(n7888) );
  NAND3_X1 U9899 ( .A1(n8726), .A2(n8725), .A3(n7895), .ZN(n7889) );
  NAND2_X1 U9900 ( .A1(n13964), .A2(n7567), .ZN(n7901) );
  OAI211_X1 U9901 ( .C1(n13964), .C2(n7902), .A(n16451), .B(n7901), .ZN(n9542)
         );
  NAND2_X1 U9902 ( .A1(n13964), .A2(n13965), .ZN(n13963) );
  OAI21_X1 U9903 ( .B1(n13964), .B2(n9518), .A(n7907), .ZN(n13828) );
  NAND2_X1 U9904 ( .A1(n9344), .A2(n7585), .ZN(n9392) );
  NAND2_X1 U9905 ( .A1(n9344), .A2(n7473), .ZN(n9390) );
  NAND2_X1 U9906 ( .A1(n9392), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9393) );
  NAND2_X1 U9907 ( .A1(n7912), .A2(n7909), .ZN(n14401) );
  NAND2_X1 U9908 ( .A1(n14194), .A2(n14193), .ZN(n14192) );
  INV_X2 U9909 ( .A(n9450), .ZN(n13815) );
  AND2_X1 U9910 ( .A1(n8278), .A2(n7916), .ZN(n7915) );
  NAND2_X1 U9911 ( .A1(n11102), .A2(n7919), .ZN(n7916) );
  NAND2_X1 U9912 ( .A1(n8280), .A2(n7917), .ZN(n12709) );
  OR2_X2 U9914 ( .A1(n12450), .A2(n12451), .ZN(n12603) );
  OR2_X2 U9915 ( .A1(n14968), .A2(n8274), .ZN(n8267) );
  NOR2_X2 U9916 ( .A1(n15001), .A2(n8847), .ZN(n14970) );
  NAND2_X1 U9917 ( .A1(n9721), .A2(n9581), .ZN(n9718) );
  NAND2_X2 U9918 ( .A1(n10232), .A2(n13345), .ZN(n14937) );
  NAND2_X1 U9919 ( .A1(n7934), .A2(n13669), .ZN(n13670) );
  NAND2_X1 U9920 ( .A1(n8055), .A2(n7935), .ZN(n7934) );
  NAND3_X1 U9921 ( .A1(n13667), .A2(n13612), .A3(n13668), .ZN(n7935) );
  INV_X1 U9922 ( .A(n10430), .ZN(n13667) );
  NAND2_X1 U9923 ( .A1(n13788), .A2(n13789), .ZN(n13787) );
  NAND2_X1 U9924 ( .A1(n13756), .A2(n7942), .ZN(n7941) );
  NAND2_X1 U9925 ( .A1(n13733), .A2(n7488), .ZN(n7947) );
  NAND2_X1 U9926 ( .A1(n13762), .A2(n13761), .ZN(n7959) );
  AND2_X1 U9927 ( .A1(n7956), .A2(n7953), .ZN(n13773) );
  NAND3_X1 U9928 ( .A1(n7959), .A2(n7958), .A3(n7957), .ZN(n7956) );
  INV_X1 U9929 ( .A(n13767), .ZN(n7960) );
  NAND3_X1 U9930 ( .A1(n13710), .A2(n13709), .A3(n7586), .ZN(n7961) );
  NAND2_X1 U9931 ( .A1(n7961), .A2(n7589), .ZN(n8116) );
  NAND2_X1 U9932 ( .A1(n8839), .A2(n10247), .ZN(n10053) );
  NAND3_X1 U9933 ( .A1(n8839), .A2(n10247), .A3(n7964), .ZN(n16117) );
  NAND2_X1 U9934 ( .A1(n13705), .A2(n13706), .ZN(n13704) );
  NAND2_X1 U9935 ( .A1(n9917), .A2(n9916), .ZN(n8014) );
  OAI21_X1 U9936 ( .B1(n9896), .B2(n9873), .A(n7590), .ZN(n7985) );
  NAND2_X1 U9937 ( .A1(n9870), .A2(n7987), .ZN(n7986) );
  INV_X1 U9938 ( .A(n9888), .ZN(n7988) );
  NAND2_X1 U9939 ( .A1(n7990), .A2(n7989), .ZN(n9974) );
  NAND3_X1 U9940 ( .A1(n9938), .A2(n9937), .A3(n9954), .ZN(n7990) );
  NOR2_X1 U9941 ( .A1(n15883), .A2(n8539), .ZN(n15858) );
  NAND2_X1 U9942 ( .A1(n15837), .A2(n15779), .ZN(n15813) );
  OAI21_X1 U9943 ( .B1(n15837), .B2(n8405), .A(n8000), .ZN(n8560) );
  NAND2_X1 U9944 ( .A1(n15837), .A2(n8000), .ZN(n7999) );
  NAND2_X1 U9945 ( .A1(n10001), .A2(n10000), .ZN(n8664) );
  INV_X1 U9946 ( .A(n8663), .ZN(n8662) );
  OAI21_X2 U9947 ( .B1(n15280), .B2(n15126), .A(n15127), .ZN(n15270) );
  OAI21_X1 U9948 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(n16348), .A(n16347), .ZN(
        n16352) );
  OAI21_X1 U9949 ( .B1(n13051), .B2(n8799), .A(n8798), .ZN(n8797) );
  NOR2_X1 U9950 ( .A1(n13349), .A2(n8010), .ZN(n13354) );
  NAND2_X1 U9951 ( .A1(n8012), .A2(n8011), .ZN(n8010) );
  NAND2_X1 U9952 ( .A1(n13346), .A2(n13347), .ZN(n8011) );
  INV_X1 U9953 ( .A(n13348), .ZN(n8013) );
  NAND3_X1 U9954 ( .A1(n13016), .A2(n8083), .A3(n13014), .ZN(n13027) );
  NAND2_X2 U9955 ( .A1(n8014), .A2(n9919), .ZN(n9938) );
  NAND2_X1 U9956 ( .A1(n15125), .A2(n15124), .ZN(n15280) );
  OAI22_X2 U9957 ( .A1(n15194), .A2(n15164), .B1(n15481), .B2(n15163), .ZN(
        n15177) );
  XNOR2_X2 U9958 ( .A(n9871), .B(SI_4_), .ZN(n9888) );
  INV_X1 U9959 ( .A(n15925), .ZN(n15758) );
  NAND2_X1 U9960 ( .A1(n8036), .A2(n8035), .ZN(n8034) );
  INV_X1 U9961 ( .A(n8317), .ZN(n8316) );
  AOI21_X1 U9962 ( .B1(n15177), .B2(n15165), .A(n8016), .ZN(n15138) );
  NAND2_X1 U9963 ( .A1(n15394), .A2(n7516), .ZN(P2_U3527) );
  NAND2_X1 U9964 ( .A1(n15476), .A2(n7492), .ZN(P2_U3495) );
  XNOR2_X1 U9965 ( .A(n12627), .B(n13832), .ZN(n12626) );
  INV_X1 U9966 ( .A(n8633), .ZN(n8632) );
  NOR2_X1 U9967 ( .A1(n8269), .A2(n12993), .ZN(n8268) );
  NAND2_X1 U9968 ( .A1(n8400), .A2(n8665), .ZN(n12627) );
  NAND2_X1 U9969 ( .A1(n8699), .A2(n15220), .ZN(n8696) );
  OAI21_X1 U9970 ( .B1(n13032), .B2(n13031), .A(n13030), .ZN(n13040) );
  NAND2_X1 U9971 ( .A1(n12514), .A2(n12513), .ZN(n12830) );
  OAI22_X1 U9972 ( .A1(n9243), .A2(n8918), .B1(P1_DATAO_REG_19__SCAN_IN), .B2(
        n11887), .ZN(n9261) );
  NAND2_X1 U9973 ( .A1(n8344), .A2(n13474), .ZN(n8343) );
  NAND2_X1 U9974 ( .A1(n14164), .A2(n14163), .ZN(n14162) );
  INV_X1 U9975 ( .A(n8346), .ZN(n8345) );
  NAND2_X1 U9976 ( .A1(n8916), .A2(n8039), .ZN(n8942) );
  INV_X1 U9977 ( .A(n14193), .ZN(n8347) );
  NAND2_X2 U9978 ( .A1(n12834), .A2(n12833), .ZN(n16040) );
  NAND2_X1 U9979 ( .A1(n8530), .A2(n8531), .ZN(n15767) );
  NAND2_X1 U9980 ( .A1(n11343), .A2(n8553), .ZN(n8551) );
  OAI21_X2 U9981 ( .B1(n15845), .B2(n15835), .A(n8615), .ZN(n15837) );
  INV_X1 U9982 ( .A(n11881), .ZN(n8375) );
  NAND2_X1 U9983 ( .A1(n13150), .A2(n8052), .ZN(n13154) );
  NAND2_X1 U9984 ( .A1(n8108), .A2(n8616), .ZN(n8613) );
  INV_X1 U9985 ( .A(n15801), .ZN(n15802) );
  NAND3_X1 U9986 ( .A1(n13164), .A2(n8102), .A3(n7591), .ZN(n8794) );
  NAND2_X1 U9987 ( .A1(n13074), .A2(n13073), .ZN(n8026) );
  INV_X1 U9988 ( .A(n13292), .ZN(n8687) );
  NAND2_X1 U9989 ( .A1(n8026), .A2(n8025), .ZN(n8027) );
  NAND3_X1 U9990 ( .A1(n13285), .A2(n8688), .A3(n13284), .ZN(n8024) );
  AOI21_X1 U9991 ( .B1(n8030), .B2(n8029), .A(n8810), .ZN(n8028) );
  INV_X1 U9992 ( .A(n13084), .ZN(n8105) );
  INV_X1 U9993 ( .A(n13073), .ZN(n8029) );
  INV_X1 U9994 ( .A(n13074), .ZN(n8030) );
  NAND2_X1 U9995 ( .A1(n8028), .A2(n8027), .ZN(n8808) );
  NAND2_X1 U9996 ( .A1(n8054), .A2(n8053), .ZN(n8052) );
  OAI21_X1 U9997 ( .B1(n13214), .B2(n13213), .A(n8858), .ZN(n13285) );
  NAND3_X1 U9998 ( .A1(n8031), .A2(n7592), .A3(n13096), .ZN(n8802) );
  NAND2_X1 U9999 ( .A1(n13091), .A2(n13090), .ZN(n8031) );
  NAND2_X1 U10000 ( .A1(n8808), .A2(n8809), .ZN(n13085) );
  NOR2_X1 U10001 ( .A1(n12620), .A2(n12509), .ZN(n8401) );
  NAND2_X1 U10002 ( .A1(n8073), .A2(n13797), .ZN(n8072) );
  NAND2_X1 U10003 ( .A1(n13944), .A2(n7573), .ZN(n8734) );
  INV_X1 U10004 ( .A(n11840), .ZN(n8718) );
  NAND2_X1 U10005 ( .A1(n11969), .A2(n11968), .ZN(n11967) );
  OR2_X1 U10006 ( .A1(n9462), .A2(n12240), .ZN(n8037) );
  NAND2_X1 U10007 ( .A1(n8087), .A2(n8086), .ZN(n12417) );
  INV_X1 U10008 ( .A(n15239), .ZN(n8770) );
  INV_X4 U10009 ( .A(n13815), .ZN(n9516) );
  NAND2_X1 U10010 ( .A1(n9673), .A2(n11215), .ZN(n11216) );
  INV_X1 U10011 ( .A(n9685), .ZN(n8038) );
  NAND2_X1 U10012 ( .A1(n8920), .A2(n8581), .ZN(n8921) );
  NAND2_X1 U10013 ( .A1(n8942), .A2(n8940), .ZN(n8917) );
  OAI21_X1 U10014 ( .B1(n9055), .B2(n9053), .A(n8905), .ZN(n9067) );
  OAI21_X1 U10015 ( .B1(n8931), .B2(n8929), .A(n7633), .ZN(n8597) );
  NAND2_X1 U10016 ( .A1(n8593), .A2(n8592), .ZN(n8043) );
  NAND2_X1 U10017 ( .A1(n13945), .A2(n14219), .ZN(n13944) );
  INV_X1 U10018 ( .A(n8041), .ZN(n13552) );
  INV_X1 U10019 ( .A(n12416), .ZN(n8087) );
  NAND2_X1 U10020 ( .A1(n8964), .A2(n8973), .ZN(n8963) );
  NAND2_X1 U10021 ( .A1(n9514), .A2(n13886), .ZN(n13888) );
  NOR2_X1 U10022 ( .A1(n11421), .A2(n8728), .ZN(n8730) );
  NAND2_X1 U10023 ( .A1(n8657), .A2(n8658), .ZN(n13784) );
  NAND2_X1 U10024 ( .A1(n8047), .A2(n8046), .ZN(n13665) );
  NAND2_X1 U10025 ( .A1(n13015), .A2(n13309), .ZN(n10546) );
  NAND2_X1 U10026 ( .A1(n8048), .A2(n11727), .ZN(n11729) );
  NAND2_X1 U10027 ( .A1(n11726), .A2(n11725), .ZN(n8048) );
  NOR2_X1 U10028 ( .A1(n8049), .A2(n8070), .ZN(n13807) );
  NAND3_X1 U10029 ( .A1(n13802), .A2(n8652), .A3(n8653), .ZN(n8049) );
  INV_X1 U10030 ( .A(n15384), .ZN(n8716) );
  NAND2_X1 U10031 ( .A1(n13796), .A2(n8655), .ZN(n8654) );
  NAND2_X1 U10032 ( .A1(n8057), .A2(n8056), .ZN(n13756) );
  NAND2_X1 U10033 ( .A1(n8114), .A2(n8113), .ZN(n13733) );
  NAND2_X1 U10034 ( .A1(n8116), .A2(n8115), .ZN(n13722) );
  INV_X1 U10035 ( .A(n15829), .ZN(n8108) );
  NAND2_X1 U10036 ( .A1(n15844), .A2(n15843), .ZN(n15842) );
  NAND2_X1 U10037 ( .A1(n8607), .A2(n8609), .ZN(n8606) );
  NAND2_X1 U10038 ( .A1(n16014), .A2(n8554), .ZN(n16100) );
  INV_X1 U10039 ( .A(n13149), .ZN(n8054) );
  NAND2_X4 U10040 ( .A1(n8251), .A2(n12171), .ZN(n15511) );
  NAND2_X1 U10041 ( .A1(n8069), .A2(n13683), .ZN(n8651) );
  INV_X1 U10042 ( .A(n10628), .ZN(n10626) );
  NAND2_X1 U10043 ( .A1(n15593), .A2(n12727), .ZN(n15604) );
  NAND3_X1 U10044 ( .A1(n13676), .A2(n13674), .A3(n13675), .ZN(n8069) );
  NAND4_X1 U10045 ( .A1(n13335), .A2(n7525), .A3(n13334), .A4(n15167), .ZN(
        n8071) );
  OAI22_X2 U10046 ( .A1(n10618), .A2(n8660), .B1(n10620), .B2(n14647), .ZN(
        n10628) );
  NOR2_X1 U10047 ( .A1(n7464), .A2(n8392), .ZN(n8391) );
  NAND2_X1 U10048 ( .A1(n15604), .A2(n15605), .ZN(n15603) );
  NAND2_X1 U10049 ( .A1(n15626), .A2(n12795), .ZN(n15576) );
  NAND2_X1 U10050 ( .A1(n12717), .A2(n7523), .ZN(n15593) );
  NAND3_X1 U10051 ( .A1(n8075), .A2(n13486), .A3(n14163), .ZN(n13487) );
  XNOR2_X1 U10052 ( .A(n15138), .B(n15167), .ZN(n15387) );
  NAND2_X1 U10053 ( .A1(n8780), .A2(n7580), .ZN(n13149) );
  NAND2_X1 U10054 ( .A1(n13149), .A2(n13148), .ZN(n13147) );
  NAND3_X1 U10055 ( .A1(n13160), .A2(n13013), .A3(n13012), .ZN(n8083) );
  NAND2_X1 U10056 ( .A1(n8103), .A2(n13068), .ZN(n13074) );
  NAND2_X1 U10057 ( .A1(n12511), .A2(n12510), .ZN(n12514) );
  NAND2_X1 U10058 ( .A1(n15767), .A2(n15766), .ZN(n15970) );
  INV_X1 U10059 ( .A(n8547), .ZN(n8546) );
  XNOR2_X2 U10060 ( .A(n8084), .B(n7614), .ZN(n16136) );
  NAND2_X1 U10061 ( .A1(n8737), .A2(n9505), .ZN(n8736) );
  NAND3_X1 U10062 ( .A1(n11331), .A2(n8733), .A3(n8085), .ZN(n8729) );
  NAND2_X1 U10063 ( .A1(n8717), .A2(n8719), .ZN(n11839) );
  NAND2_X1 U10064 ( .A1(n9226), .A2(n9225), .ZN(n8916) );
  INV_X1 U10065 ( .A(n8597), .ZN(n9313) );
  OAI22_X1 U10066 ( .A1(n11645), .A2(n11390), .B1(n11391), .B2(n13071), .ZN(
        n11587) );
  NOR2_X1 U10067 ( .A1(n8395), .A2(n8290), .ZN(n8289) );
  NAND2_X1 U10068 ( .A1(n16009), .A2(n16561), .ZN(n8110) );
  NAND2_X1 U10069 ( .A1(n15836), .A2(n15837), .ZN(n8098) );
  NAND2_X1 U10070 ( .A1(n9868), .A2(n9869), .ZN(n8112) );
  NAND2_X1 U10071 ( .A1(n15265), .A2(n15155), .ZN(n8690) );
  OAI21_X1 U10072 ( .B1(n13067), .B2(n13066), .A(n13065), .ZN(n8103) );
  INV_X1 U10073 ( .A(n13050), .ZN(n8800) );
  NAND2_X1 U10074 ( .A1(n9874), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n8107) );
  NAND3_X1 U10075 ( .A1(n8734), .A2(n13914), .A3(n14208), .ZN(n13842) );
  OAI21_X2 U10076 ( .B1(n8656), .B2(n13795), .A(n13794), .ZN(n13796) );
  NAND2_X1 U10077 ( .A1(n14129), .A2(n14128), .ZN(n8174) );
  OAI211_X1 U10078 ( .C1(n14148), .C2(n16429), .A(n8441), .B(n8438), .ZN(
        P3_U3201) );
  NAND2_X1 U10079 ( .A1(n9657), .A2(n11524), .ZN(n8190) );
  AND2_X1 U10080 ( .A1(n13552), .A2(n8123), .ZN(n13561) );
  INV_X1 U10081 ( .A(n9320), .ZN(n8122) );
  INV_X1 U10082 ( .A(n8562), .ZN(n8561) );
  NAND2_X1 U10083 ( .A1(n8917), .A2(n8119), .ZN(n9243) );
  OAI21_X1 U10084 ( .B1(n8912), .B2(n8566), .A(n8913), .ZN(n8562) );
  NAND2_X1 U10085 ( .A1(n15340), .A2(n15339), .ZN(n15338) );
  NAND2_X1 U10086 ( .A1(n10540), .A2(n10539), .ZN(n10483) );
  AND2_X1 U10087 ( .A1(n15754), .A2(n15752), .ZN(n8603) );
  NAND2_X1 U10088 ( .A1(n8377), .A2(n8926), .ZN(n8253) );
  NAND2_X1 U10089 ( .A1(n11389), .A2(n11388), .ZN(n11645) );
  OAI211_X1 U10090 ( .C1(n16738), .C2(n15387), .A(n8716), .B(n8714), .ZN(
        n15473) );
  NAND3_X1 U10091 ( .A1(n13727), .A2(n13726), .A3(n7587), .ZN(n8114) );
  AND2_X2 U10092 ( .A1(n13793), .A2(n13792), .ZN(n8656) );
  INV_X1 U10093 ( .A(n13679), .ZN(n13682) );
  NAND2_X1 U10094 ( .A1(n8378), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n8252) );
  OAI21_X2 U10095 ( .B1(n9874), .B2(P2_DATAO_REG_4__SCAN_IN), .A(n8118), .ZN(
        n9871) );
  NAND2_X1 U10096 ( .A1(n8900), .A2(n8899), .ZN(n8997) );
  AOI21_X1 U10097 ( .B1(n13553), .B2(n13554), .A(n8124), .ZN(n8123) );
  NAND2_X1 U10098 ( .A1(n14192), .A2(n8140), .ZN(n8136) );
  NAND2_X1 U10099 ( .A1(n8135), .A2(n8134), .ZN(n14157) );
  NAND2_X1 U10100 ( .A1(n14192), .A2(n8137), .ZN(n8135) );
  NAND2_X1 U10101 ( .A1(n11827), .A2(n11824), .ZN(n9020) );
  NAND2_X1 U10102 ( .A1(n7581), .A2(n8990), .ZN(n11827) );
  NAND2_X1 U10103 ( .A1(n12286), .A2(n8156), .ZN(n8155) );
  NAND2_X1 U10104 ( .A1(n12286), .A2(n9124), .ZN(n12392) );
  NAND2_X1 U10105 ( .A1(n8155), .A2(n8159), .ZN(n9174) );
  NAND2_X1 U10106 ( .A1(n8167), .A2(n9359), .ZN(n16493) );
  NAND3_X1 U10107 ( .A1(n8167), .A2(n13358), .A3(n13357), .ZN(n13359) );
  AND2_X2 U10108 ( .A1(n8171), .A2(n7462), .ZN(n8945) );
  NAND3_X1 U10109 ( .A1(n8742), .A2(n8353), .A3(n8044), .ZN(n8173) );
  NAND2_X1 U10110 ( .A1(n11923), .A2(n7574), .ZN(n12039) );
  NAND2_X1 U10111 ( .A1(n12039), .A2(n9106), .ZN(n9123) );
  INV_X1 U10112 ( .A(n8176), .ZN(n8175) );
  NAND2_X1 U10113 ( .A1(n8176), .A2(n14037), .ZN(n14056) );
  NOR2_X1 U10114 ( .A1(n11614), .A2(n11613), .ZN(n11612) );
  AOI21_X1 U10115 ( .B1(n11614), .B2(n7605), .A(n8185), .ZN(n8178) );
  NAND2_X1 U10116 ( .A1(n11614), .A2(n8180), .ZN(n8179) );
  NOR2_X1 U10117 ( .A1(n8184), .A2(n8182), .ZN(n8181) );
  AOI21_X1 U10118 ( .B1(n11198), .B2(n7480), .A(n11197), .ZN(n11201) );
  XNOR2_X1 U10119 ( .A(n11220), .B(n10868), .ZN(n10854) );
  NAND2_X1 U10120 ( .A1(n8196), .A2(n8193), .ZN(n8192) );
  NOR2_X1 U10121 ( .A1(n8194), .A2(n9684), .ZN(n8193) );
  INV_X1 U10122 ( .A(n8195), .ZN(n8194) );
  NAND3_X1 U10123 ( .A1(n14760), .A2(n14761), .A3(n8231), .ZN(n8230) );
  OAI21_X2 U10124 ( .B1(n9972), .B2(n8399), .A(n9975), .ZN(n10001) );
  NAND2_X4 U10125 ( .A1(n8253), .A2(n8252), .ZN(n9874) );
  NAND2_X1 U10126 ( .A1(n8254), .A2(n8261), .ZN(n8257) );
  INV_X1 U10127 ( .A(n8503), .ZN(n8254) );
  INV_X1 U10128 ( .A(n14945), .ZN(n8260) );
  OAI211_X1 U10129 ( .C1(n14945), .C2(n8505), .A(n8503), .B(n8256), .ZN(n8255)
         );
  NAND2_X1 U10130 ( .A1(n8260), .A2(n7572), .ZN(n8259) );
  NAND4_X1 U10131 ( .A1(n8259), .A2(n8258), .A3(n8257), .A4(n8255), .ZN(
        P2_U3192) );
  NAND3_X1 U10132 ( .A1(n8271), .A2(n8268), .A3(n8267), .ZN(n8276) );
  INV_X1 U10133 ( .A(n8276), .ZN(n14922) );
  AND2_X2 U10134 ( .A1(n8276), .A2(n8275), .ZN(n14925) );
  NAND2_X1 U10135 ( .A1(n8277), .A2(n14923), .ZN(n8275) );
  NOR2_X1 U10136 ( .A1(n7484), .A2(n8279), .ZN(n8278) );
  AND2_X1 U10137 ( .A1(n12702), .A2(n8281), .ZN(n8280) );
  OR2_X1 U10138 ( .A1(n11365), .A2(n7484), .ZN(n8281) );
  NAND2_X1 U10139 ( .A1(n11184), .A2(n8285), .ZN(n8284) );
  NAND2_X1 U10140 ( .A1(n8284), .A2(n8283), .ZN(n11101) );
  XNOR2_X2 U10141 ( .A(n10617), .B(SI_14_), .ZN(n10618) );
  INV_X1 U10142 ( .A(n8498), .ZN(n8501) );
  XNOR2_X1 U10143 ( .A(n13054), .B(n14936), .ZN(n10651) );
  NAND2_X2 U10144 ( .A1(n12814), .A2(n9874), .ZN(n10704) );
  NAND2_X2 U10145 ( .A1(n10019), .A2(n16240), .ZN(n12814) );
  NAND2_X1 U10146 ( .A1(n9724), .A2(n8312), .ZN(n9580) );
  AND2_X2 U10147 ( .A1(n7421), .A2(n11323), .ZN(n11642) );
  OR2_X1 U10148 ( .A1(n15198), .A2(n15468), .ZN(n8313) );
  AND2_X1 U10149 ( .A1(n15198), .A2(n8317), .ZN(n15139) );
  NAND2_X1 U10150 ( .A1(n15198), .A2(n15477), .ZN(n15183) );
  OAI21_X2 U10151 ( .B1(n16491), .B2(n8333), .A(n8330), .ZN(n11823) );
  NAND2_X1 U10152 ( .A1(n11920), .A2(n8335), .ZN(n8334) );
  NAND2_X1 U10153 ( .A1(n8334), .A2(n7577), .ZN(n11944) );
  CLKBUF_X1 U10154 ( .A(n14210), .Z(n8341) );
  AOI21_X2 U10155 ( .B1(n14210), .B2(n7508), .A(n8343), .ZN(n14171) );
  NAND4_X1 U10156 ( .A1(n8742), .A2(n8353), .A3(n8044), .A4(n9165), .ZN(n9227)
         );
  AOI21_X2 U10157 ( .B1(n8361), .B2(n8360), .A(n8357), .ZN(n13516) );
  INV_X2 U10158 ( .A(n10517), .ZN(n11817) );
  NAND2_X1 U10159 ( .A1(n12049), .A2(n8369), .ZN(n8368) );
  NAND2_X1 U10160 ( .A1(n8945), .A2(n8373), .ZN(n8887) );
  NAND2_X1 U10161 ( .A1(n8945), .A2(n7584), .ZN(n14903) );
  NAND3_X1 U10162 ( .A1(n16405), .A2(P3_ADDR_REG_19__SCAN_IN), .A3(n16441), 
        .ZN(n8377) );
  NAND3_X1 U10163 ( .A1(n8925), .A2(n8379), .A3(P2_ADDR_REG_19__SCAN_IN), .ZN(
        n8378) );
  NAND2_X1 U10164 ( .A1(n8384), .A2(n8381), .ZN(n11882) );
  NAND2_X1 U10165 ( .A1(n12511), .A2(n8401), .ZN(n8400) );
  INV_X1 U10166 ( .A(n12626), .ZN(n12855) );
  NAND3_X1 U10167 ( .A1(n13628), .A2(n15783), .A3(n8403), .ZN(n8402) );
  INV_X1 U10168 ( .A(n9669), .ZN(n8408) );
  NOR2_X1 U10169 ( .A1(n8408), .A2(n11411), .ZN(n8407) );
  NAND3_X1 U10170 ( .A1(n8411), .A2(n8410), .A3(n11310), .ZN(n8409) );
  OAI22_X1 U10171 ( .A1(n8962), .A2(n8413), .B1(P3_IR_REG_1__SCAN_IN), .B2(
        P3_IR_REG_31__SCAN_IN), .ZN(n8412) );
  INV_X1 U10172 ( .A(n8418), .ZN(n16421) );
  NAND2_X1 U10173 ( .A1(n8423), .A2(n8424), .ZN(n8422) );
  INV_X1 U10174 ( .A(n14014), .ZN(n8431) );
  NAND2_X1 U10175 ( .A1(n8431), .A2(n13999), .ZN(n14000) );
  NAND2_X1 U10176 ( .A1(n13999), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n8433) );
  AOI21_X1 U10177 ( .B1(n7500), .B2(n7459), .A(n8445), .ZN(n14623) );
  OAI22_X1 U10178 ( .A1(n10007), .A2(keyinput_117), .B1(n14614), .B2(
        P1_IR_REG_10__SCAN_IN), .ZN(n8454) );
  AND2_X1 U10179 ( .A1(n14611), .A2(n14612), .ZN(n8455) );
  NAND3_X1 U10180 ( .A1(n8484), .A2(n14488), .A3(n8483), .ZN(n8482) );
  AOI221_X1 U10181 ( .B1(n14581), .B2(n14580), .C1(keyinput_92), .C2(
        P3_DATAO_REG_4__SCAN_IN), .A(n14579), .ZN(n14589) );
  OAI21_X1 U10182 ( .B1(n14496), .B2(n14495), .A(n14494), .ZN(n14497) );
  NAND2_X1 U10183 ( .A1(n7468), .A2(n9701), .ZN(n8694) );
  NAND2_X1 U10184 ( .A1(n8496), .A2(n11047), .ZN(n8499) );
  AND2_X1 U10185 ( .A1(n10982), .A2(n9733), .ZN(n10566) );
  NOR2_X1 U10186 ( .A1(n14945), .A2(n14944), .ZN(n14958) );
  INV_X1 U10187 ( .A(n14944), .ZN(n8509) );
  NOR2_X1 U10188 ( .A1(n8517), .A2(P2_ADDR_REG_15__SCAN_IN), .ZN(n8512) );
  NAND3_X1 U10189 ( .A1(n16383), .A2(n16382), .A3(n8514), .ZN(n8513) );
  OAI21_X1 U10190 ( .B1(n16383), .B2(n11454), .A(n16382), .ZN(n16389) );
  NAND2_X1 U10191 ( .A1(n12709), .A2(n8523), .ZN(n12061) );
  NAND2_X1 U10192 ( .A1(n8541), .A2(n8540), .ZN(n11149) );
  AND2_X1 U10193 ( .A1(n8543), .A2(n13578), .ZN(n8540) );
  NAND2_X1 U10194 ( .A1(n11147), .A2(n8544), .ZN(n8541) );
  AND2_X1 U10195 ( .A1(n16554), .A2(n13678), .ZN(n8545) );
  NAND2_X1 U10196 ( .A1(n8551), .A2(n8550), .ZN(n11750) );
  OAI21_X1 U10197 ( .B1(n16468), .B2(n16461), .A(n13669), .ZN(n10933) );
  NAND2_X2 U10198 ( .A1(n13669), .A2(n10431), .ZN(n16468) );
  NAND2_X1 U10199 ( .A1(n8563), .A2(n8561), .ZN(n9189) );
  NAND2_X1 U10200 ( .A1(n9164), .A2(n8564), .ZN(n8563) );
  NAND2_X1 U10201 ( .A1(n8565), .A2(n8912), .ZN(n9177) );
  INV_X1 U10202 ( .A(n9176), .ZN(n8566) );
  OR2_X1 U10203 ( .A1(n9334), .A2(n9333), .ZN(n8593) );
  NAND2_X1 U10204 ( .A1(n8583), .A2(n8584), .ZN(n13499) );
  NAND2_X1 U10205 ( .A1(n9334), .A2(n8589), .ZN(n8583) );
  INV_X1 U10206 ( .A(n9333), .ZN(n8594) );
  INV_X1 U10207 ( .A(n16090), .ZN(n8605) );
  INV_X1 U10208 ( .A(n8611), .ZN(n15918) );
  INV_X1 U10209 ( .A(n15760), .ZN(n8610) );
  NAND2_X1 U10210 ( .A1(n11572), .A2(n8624), .ZN(n8621) );
  INV_X1 U10211 ( .A(n15686), .ZN(n8629) );
  NAND2_X1 U10212 ( .A1(n8630), .A2(n8631), .ZN(n15844) );
  NAND2_X1 U10213 ( .A1(n15876), .A2(n8843), .ZN(n15871) );
  NAND2_X1 U10214 ( .A1(n12324), .A2(n7449), .ZN(n12337) );
  XNOR2_X1 U10215 ( .A(n15690), .B(n16527), .ZN(n13671) );
  NAND2_X1 U10216 ( .A1(n9553), .A2(n8641), .ZN(n8636) );
  NAND2_X1 U10217 ( .A1(n13742), .A2(n13743), .ZN(n13741) );
  NAND2_X1 U10218 ( .A1(n13763), .A2(n13764), .ZN(n13762) );
  NAND2_X1 U10219 ( .A1(n13722), .A2(n13723), .ZN(n13721) );
  NAND2_X1 U10220 ( .A1(n13696), .A2(n13694), .ZN(n13688) );
  NAND2_X1 U10221 ( .A1(n8651), .A2(n13687), .ZN(n13694) );
  NAND2_X1 U10222 ( .A1(n8654), .A2(n13801), .ZN(n8652) );
  NAND2_X1 U10223 ( .A1(n8656), .A2(n13795), .ZN(n8655) );
  NAND3_X1 U10224 ( .A1(n13778), .A2(n13777), .A3(n7578), .ZN(n8657) );
  NAND4_X2 U10225 ( .A1(n9744), .A2(n9742), .A3(n9743), .A4(n8691), .ZN(n15043) );
  OR2_X1 U10226 ( .A1(n15239), .A2(n8700), .ZN(n8699) );
  AND2_X1 U10227 ( .A1(n8730), .A2(n11334), .ZN(n11419) );
  NAND2_X1 U10228 ( .A1(n8733), .A2(n11331), .ZN(n11334) );
  NAND2_X1 U10229 ( .A1(n9402), .A2(n7448), .ZN(n9447) );
  NAND2_X1 U10230 ( .A1(n8739), .A2(n9428), .ZN(n9418) );
  XNOR2_X1 U10231 ( .A(n11008), .B(n8739), .ZN(n9430) );
  NAND2_X1 U10232 ( .A1(n9390), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9391) );
  INV_X1 U10233 ( .A(n8755), .ZN(n8753) );
  AOI21_X2 U10234 ( .B1(n8757), .B2(n12498), .A(n7433), .ZN(n8755) );
  NAND2_X1 U10235 ( .A1(n8764), .A2(n8763), .ZN(n11237) );
  INV_X1 U10236 ( .A(n13142), .ZN(n8781) );
  INV_X1 U10237 ( .A(n13141), .ZN(n8782) );
  NAND2_X1 U10238 ( .A1(n8783), .A2(n7579), .ZN(n13116) );
  INV_X1 U10239 ( .A(n13110), .ZN(n8785) );
  NAND2_X1 U10240 ( .A1(n8786), .A2(n8787), .ZN(n13162) );
  NAND2_X1 U10241 ( .A1(n13154), .A2(n8789), .ZN(n8786) );
  INV_X1 U10242 ( .A(n13122), .ZN(n8793) );
  NAND2_X1 U10243 ( .A1(n8794), .A2(n8795), .ZN(n13192) );
  AOI21_X1 U10244 ( .B1(n13192), .B2(n13191), .A(n13190), .ZN(n13214) );
  AND2_X1 U10245 ( .A1(n13050), .A2(n13049), .ZN(n8799) );
  OR2_X1 U10246 ( .A1(n11688), .A2(n11689), .ZN(n8827) );
  NAND2_X1 U10247 ( .A1(n11019), .A2(n11020), .ZN(n8828) );
  NAND3_X1 U10248 ( .A1(n8830), .A2(n8829), .A3(n9543), .ZN(n9863) );
  INV_X1 U10249 ( .A(n8837), .ZN(n12401) );
  OR2_X1 U10250 ( .A1(n12378), .A2(n12379), .ZN(n8838) );
  NAND2_X1 U10251 ( .A1(n10247), .A2(n9994), .ZN(n9997) );
  INV_X1 U10252 ( .A(n15329), .ZN(n15504) );
  NAND2_X1 U10253 ( .A1(n10566), .A2(n10565), .ZN(n11128) );
  NAND2_X2 U10254 ( .A1(n12317), .A2(n12316), .ZN(n12345) );
  NOR2_X2 U10255 ( .A1(n15212), .A2(n15195), .ZN(n15198) );
  OR2_X2 U10256 ( .A1(n15227), .A2(n15211), .ZN(n15212) );
  XNOR2_X1 U10257 ( .A(n13216), .B(n13215), .ZN(n13599) );
  NAND2_X1 U10258 ( .A1(n11348), .A2(n11347), .ZN(n11572) );
  XNOR2_X1 U10259 ( .A(n12716), .B(n12714), .ZN(n15666) );
  NAND2_X1 U10260 ( .A1(n10362), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n10363) );
  INV_X1 U10261 ( .A(n13346), .ZN(n13337) );
  OR2_X1 U10262 ( .A1(n13808), .A2(n7411), .ZN(n11002) );
  XNOR2_X1 U10263 ( .A(n12892), .B(n7613), .ZN(n15532) );
  XNOR2_X1 U10264 ( .A(n13607), .B(n13606), .ZN(n13616) );
  NAND2_X2 U10265 ( .A1(n13368), .A2(n13364), .ZN(n16499) );
  OAI21_X1 U10266 ( .B1(n12577), .B2(n9465), .A(n12417), .ZN(n12576) );
  NOR2_X1 U10267 ( .A1(n8958), .A2(n8853), .ZN(n8961) );
  INV_X1 U10268 ( .A(n9389), .ZN(n9348) );
  INV_X1 U10269 ( .A(n10356), .ZN(n16120) );
  AND2_X2 U10270 ( .A1(n15526), .A2(n9704), .ZN(n9790) );
  INV_X2 U10271 ( .A(n16717), .ZN(n16718) );
  AND2_X1 U10272 ( .A1(n8842), .A2(n9426), .ZN(n8840) );
  INV_X1 U10273 ( .A(n14307), .ZN(n14319) );
  INV_X1 U10274 ( .A(n15675), .ZN(n15778) );
  XNOR2_X1 U10275 ( .A(n13606), .B(n13605), .ZN(n8841) );
  OR2_X1 U10276 ( .A1(n13810), .A2(n14896), .ZN(n8842) );
  OR2_X1 U10277 ( .A1(n15882), .A2(n15777), .ZN(n8843) );
  INV_X1 U10278 ( .A(n14937), .ZN(n14960) );
  INV_X1 U10279 ( .A(n11246), .ZN(n13223) );
  AND2_X1 U10280 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), 
        .ZN(n8845) );
  AND2_X1 U10281 ( .A1(n7600), .A2(n9443), .ZN(n8846) );
  AND2_X1 U10282 ( .A1(n12977), .A2(n12976), .ZN(n8847) );
  NAND2_X1 U10283 ( .A1(n16017), .A2(n16660), .ZN(n8848) );
  AND2_X1 U10284 ( .A1(n15000), .A2(n14960), .ZN(n8849) );
  AND2_X1 U10285 ( .A1(n16590), .A2(n13009), .ZN(n8850) );
  INV_X1 U10286 ( .A(n9704), .ZN(n12646) );
  NOR2_X1 U10287 ( .A1(n9491), .A2(n13854), .ZN(n8851) );
  INV_X1 U10288 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n16123) );
  INV_X1 U10289 ( .A(P3_D_REG_1__SCAN_IN), .ZN(n9403) );
  NAND2_X1 U10290 ( .A1(n13002), .A2(n13001), .ZN(n15266) );
  AND2_X1 U10291 ( .A1(n7416), .A2(P1_U3086), .ZN(n11168) );
  INV_X1 U10292 ( .A(n15308), .ZN(n15346) );
  AND2_X1 U10293 ( .A1(n8980), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n8853) );
  OR2_X1 U10294 ( .A1(n13798), .A2(n13797), .ZN(n8854) );
  AND2_X1 U10295 ( .A1(n10215), .A2(n10143), .ZN(n8856) );
  AND2_X1 U10296 ( .A1(n13280), .A2(n13212), .ZN(n8858) );
  NAND2_X1 U10297 ( .A1(n15819), .A2(n16606), .ZN(n8859) );
  INV_X1 U10298 ( .A(n15981), .ZN(n15754) );
  INV_X1 U10299 ( .A(n13680), .ZN(n13681) );
  NAND2_X1 U10300 ( .A1(n13682), .A2(n13681), .ZN(n13683) );
  NAND2_X1 U10301 ( .A1(n13698), .A2(n13697), .ZN(n13700) );
  OAI21_X1 U10302 ( .B1(n13058), .B2(n8104), .A(n13057), .ZN(n13060) );
  OAI21_X1 U10303 ( .B1(n13120), .B2(n8104), .A(n13119), .ZN(n13121) );
  NAND2_X1 U10304 ( .A1(n13147), .A2(n13146), .ZN(n13150) );
  AND2_X1 U10305 ( .A1(n13343), .A2(n13351), .ZN(n13224) );
  CLKBUF_X3 U10306 ( .A(n8104), .Z(n13299) );
  NOR2_X1 U10307 ( .A1(P3_IR_REG_16__SCAN_IN), .A2(P3_IR_REG_15__SCAN_IN), 
        .ZN(n8882) );
  INV_X1 U10308 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n9544) );
  AOI21_X1 U10309 ( .B1(n14308), .B2(n14307), .A(n9241), .ZN(n14294) );
  INV_X1 U10310 ( .A(P2_B_REG_SCAN_IN), .ZN(n15112) );
  INV_X1 U10311 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n9989) );
  INV_X1 U10312 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n9555) );
  INV_X1 U10313 ( .A(P3_REG3_REG_19__SCAN_IN), .ZN(n14703) );
  OR2_X1 U10314 ( .A1(n9323), .A2(n8871), .ZN(n9324) );
  INV_X1 U10315 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n14715) );
  NAND2_X1 U10316 ( .A1(n13525), .A2(n11403), .ZN(n11402) );
  INV_X1 U10317 ( .A(n12198), .ZN(n10842) );
  INV_X1 U10318 ( .A(n15167), .ZN(n15168) );
  INV_X1 U10319 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n12453) );
  INV_X1 U10320 ( .A(n15560), .ZN(n12847) );
  AND2_X1 U10321 ( .A1(n10693), .A2(n10692), .ZN(n10694) );
  INV_X1 U10322 ( .A(n15685), .ZN(n11686) );
  INV_X1 U10323 ( .A(n13607), .ZN(n10384) );
  OR2_X1 U10324 ( .A1(n9296), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n9305) );
  INV_X1 U10325 ( .A(P3_REG3_REG_18__SCAN_IN), .ZN(n14738) );
  OR2_X1 U10326 ( .A1(n9435), .A2(n9434), .ZN(n9431) );
  INV_X1 U10327 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n8883) );
  INV_X1 U10328 ( .A(n11068), .ZN(n14929) );
  OR2_X1 U10329 ( .A1(n13201), .A2(n13200), .ZN(n13260) );
  OR2_X1 U10330 ( .A1(n12996), .A2(n12995), .ZN(n13167) );
  NAND2_X1 U10331 ( .A1(n10842), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n12454) );
  OR2_X1 U10332 ( .A1(n10772), .A2(n10771), .ZN(n10799) );
  OAI22_X1 U10333 ( .A1(n15172), .A2(n15289), .B1(n15171), .B2(n15170), .ZN(
        n15173) );
  INV_X1 U10334 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n13256) );
  OAI21_X1 U10335 ( .B1(n9813), .B2(n9812), .A(n9811), .ZN(n10223) );
  INV_X1 U10336 ( .A(n12800), .ZN(n12817) );
  INV_X1 U10337 ( .A(n12816), .ZN(n12837) );
  NOR2_X1 U10338 ( .A1(n12764), .A2(n12763), .ZN(n12782) );
  OR2_X1 U10339 ( .A1(n12025), .A2(n12024), .ZN(n12308) );
  INV_X1 U10340 ( .A(n15762), .ZN(n15872) );
  INV_X1 U10341 ( .A(n15684), .ZN(n11696) );
  INV_X1 U10342 ( .A(P1_B_REG_SCAN_IN), .ZN(n15739) );
  NOR2_X1 U10343 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), 
        .ZN(n9558) );
  INV_X1 U10344 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n14712) );
  INV_X1 U10345 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n14634) );
  OR2_X1 U10346 ( .A1(n9285), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n9296) );
  AND2_X1 U10347 ( .A1(n9332), .A2(n9331), .ZN(n14184) );
  AND2_X1 U10348 ( .A1(n9644), .A2(n9667), .ZN(n9534) );
  INV_X1 U10349 ( .A(n13387), .ZN(n13534) );
  INV_X1 U10350 ( .A(n13557), .ZN(n9434) );
  OR2_X1 U10351 ( .A1(n9335), .A2(n14477), .ZN(n9321) );
  INV_X1 U10352 ( .A(n13877), .ZN(n14831) );
  INV_X1 U10353 ( .A(n16501), .ZN(n14310) );
  INV_X1 U10354 ( .A(n16647), .ZN(n16713) );
  AND2_X1 U10355 ( .A1(n9387), .A2(n9431), .ZN(n16521) );
  NAND2_X1 U10356 ( .A1(n7623), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9424) );
  NOR2_X1 U10357 ( .A1(n15157), .A2(n14960), .ZN(n14924) );
  INV_X1 U10358 ( .A(n15033), .ZN(n13089) );
  INV_X1 U10359 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n15002) );
  AND2_X1 U10360 ( .A1(n13260), .A2(n13202), .ZN(n15214) );
  OR2_X1 U10361 ( .A1(n12608), .A2(n15002), .ZN(n12962) );
  INV_X1 U10362 ( .A(n13338), .ZN(n13341) );
  INV_X1 U10363 ( .A(n15165), .ZN(n15179) );
  INV_X1 U10364 ( .A(n15145), .ZN(n15286) );
  INV_X1 U10365 ( .A(n15324), .ZN(n15317) );
  INV_X1 U10366 ( .A(n15031), .ZN(n12697) );
  INV_X1 U10367 ( .A(n15035), .ZN(n13079) );
  NAND2_X1 U10368 ( .A1(n15353), .A2(n11258), .ZN(n15330) );
  INV_X1 U10369 ( .A(n15034), .ZN(n12664) );
  AND2_X1 U10370 ( .A1(n10228), .A2(n10227), .ZN(n15308) );
  OR2_X1 U10371 ( .A1(n16147), .A2(P2_D_REG_0__SCAN_IN), .ZN(n9817) );
  OAI21_X1 U10372 ( .B1(n7460), .B2(P2_IR_REG_23__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9586) );
  OR2_X1 U10373 ( .A1(n10150), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n10449) );
  INV_X1 U10374 ( .A(n15658), .ZN(n15648) );
  AND2_X1 U10375 ( .A1(n12782), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n12799) );
  OR2_X1 U10376 ( .A1(n12745), .A2(n12744), .ZN(n12764) );
  INV_X1 U10377 ( .A(n12814), .ZN(n12759) );
  INV_X1 U10378 ( .A(n15860), .ZN(n15777) );
  INV_X1 U10379 ( .A(n15774), .ZN(n15910) );
  INV_X1 U10380 ( .A(n15678), .ZN(n12713) );
  OR2_X1 U10381 ( .A1(n10936), .A2(n13606), .ZN(n15993) );
  NOR2_X1 U10382 ( .A1(n9559), .A2(n9558), .ZN(n9560) );
  INV_X1 U10383 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n16316) );
  OAI21_X1 U10384 ( .B1(n14850), .B2(n13985), .A(n9539), .ZN(n9540) );
  AND2_X1 U10385 ( .A1(n11012), .A2(n16652), .ZN(n9523) );
  INV_X1 U10386 ( .A(n14311), .ZN(n14348) );
  INV_X1 U10387 ( .A(n11829), .ZN(n12250) );
  INV_X1 U10388 ( .A(n16418), .ZN(n14125) );
  NAND2_X1 U10389 ( .A1(n11010), .A2(n11009), .ZN(n11014) );
  AND2_X1 U10390 ( .A1(n9534), .A2(n13480), .ZN(n16498) );
  INV_X1 U10391 ( .A(n13533), .ZN(n13409) );
  AND2_X1 U10392 ( .A1(n14352), .A2(n16515), .ZN(n14240) );
  AND2_X1 U10393 ( .A1(n9430), .A2(n9429), .ZN(n11010) );
  NAND2_X1 U10394 ( .A1(n16521), .A2(n16615), .ZN(n16647) );
  INV_X1 U10395 ( .A(n16615), .ZN(n16596) );
  AND2_X1 U10396 ( .A1(n9405), .A2(n9404), .ZN(n11008) );
  INV_X1 U10397 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n9191) );
  OR2_X1 U10398 ( .A1(n9116), .A2(P3_IR_REG_10__SCAN_IN), .ZN(n9149) );
  NOR2_X1 U10399 ( .A1(n9831), .A2(n13351), .ZN(n14991) );
  NOR2_X1 U10400 ( .A1(n9831), .A2(n9821), .ZN(n15014) );
  OR2_X1 U10401 ( .A1(n15182), .A2(n13262), .ZN(n13268) );
  INV_X1 U10402 ( .A(n9790), .ZN(n13265) );
  OR3_X1 U10403 ( .A1(n15534), .A2(n15536), .A3(n15539), .ZN(n10076) );
  AND2_X1 U10404 ( .A1(n10095), .A2(n10081), .ZN(n16231) );
  INV_X1 U10405 ( .A(n15289), .ZN(n15341) );
  INV_X1 U10406 ( .A(n13319), .ZN(n11386) );
  OAI21_X1 U10407 ( .B1(n11245), .B2(n11244), .A(n15364), .ZN(n15327) );
  AND2_X1 U10408 ( .A1(n10226), .A2(n16590), .ZN(n16738) );
  INV_X1 U10409 ( .A(n16738), .ZN(n16641) );
  AND2_X1 U10410 ( .A1(n10151), .A2(n10449), .ZN(n16232) );
  XNOR2_X1 U10411 ( .A(n12943), .B(n12942), .ZN(n12944) );
  INV_X1 U10412 ( .A(n15673), .ZN(n16531) );
  AND2_X1 U10413 ( .A1(n16528), .A2(n16606), .ZN(n15671) );
  AND4_X1 U10414 ( .A1(n12939), .A2(n12938), .A3(n12937), .A4(n12936), .ZN(
        n15815) );
  INV_X1 U10415 ( .A(n10019), .ZN(n10401) );
  OR2_X1 U10416 ( .A1(n16249), .A2(n10025), .ZN(n15728) );
  INV_X1 U10417 ( .A(n15710), .ZN(n16259) );
  INV_X1 U10418 ( .A(n15727), .ZN(n16261) );
  INV_X1 U10419 ( .A(n16464), .ZN(n16079) );
  NAND4_X1 U10420 ( .A1(n10577), .A2(n10576), .A3(n10575), .A4(n10574), .ZN(
        n15838) );
  INV_X1 U10421 ( .A(n15847), .ZN(n15843) );
  INV_X1 U10422 ( .A(n15951), .ZN(n15971) );
  INV_X1 U10423 ( .A(n15983), .ZN(n15935) );
  INV_X1 U10424 ( .A(n15993), .ZN(n16472) );
  INV_X1 U10425 ( .A(n16561), .ZN(n16726) );
  INV_X1 U10426 ( .A(n16730), .ZN(n16540) );
  NAND2_X1 U10427 ( .A1(n15993), .A2(n16475), .ZN(n16730) );
  AND2_X1 U10428 ( .A1(n11137), .A2(n11136), .ZN(n11138) );
  OAI211_X1 U10429 ( .C1(n10379), .C2(n9968), .A(n10380), .B(n9967), .ZN(
        n10381) );
  AND2_X1 U10430 ( .A1(n10642), .A2(n11166), .ZN(n12339) );
  AND2_X1 U10431 ( .A1(n9689), .A2(n9688), .ZN(n16150) );
  INV_X1 U10432 ( .A(n9540), .ZN(n9541) );
  INV_X1 U10433 ( .A(n16451), .ZN(n13954) );
  INV_X1 U10434 ( .A(n13970), .ZN(n13979) );
  NAND2_X1 U10435 ( .A1(n9524), .A2(n9523), .ZN(n13985) );
  INV_X2 U10436 ( .A(n10989), .ZN(n11041) );
  OR2_X1 U10437 ( .A1(n11212), .A2(n9667), .ZN(n16423) );
  INV_X1 U10438 ( .A(n14146), .ZN(n16427) );
  INV_X1 U10439 ( .A(n14372), .ZN(n14358) );
  INV_X2 U10440 ( .A(n14352), .ZN(n16517) );
  NAND2_X1 U10441 ( .A1(n11010), .A2(n9441), .ZN(n16717) );
  OR2_X1 U10442 ( .A1(n16717), .A2(n16711), .ZN(n14455) );
  AND3_X1 U10443 ( .A1(n16600), .A2(n16599), .A3(n16598), .ZN(n16602) );
  NAND2_X1 U10444 ( .A1(n9398), .A2(n9397), .ZN(n12294) );
  INV_X1 U10445 ( .A(n9647), .ZN(n13997) );
  INV_X2 U10446 ( .A(n9852), .ZN(n14920) );
  INV_X1 U10447 ( .A(n15408), .ZN(n15228) );
  INV_X1 U10448 ( .A(n15014), .ZN(n15021) );
  INV_X1 U10449 ( .A(n15024), .ZN(n14994) );
  NAND2_X1 U10450 ( .A1(n13208), .A2(n13207), .ZN(n15162) );
  NAND2_X1 U10451 ( .A1(n12992), .A2(n12991), .ZN(n15145) );
  INV_X1 U10452 ( .A(n16231), .ZN(n16214) );
  INV_X1 U10453 ( .A(n15371), .ZN(n15233) );
  NAND2_X1 U10454 ( .A1(n16747), .A2(n16740), .ZN(n15464) );
  INV_X1 U10455 ( .A(n16747), .ZN(n16746) );
  AND2_X2 U10456 ( .A1(n10240), .A2(n11242), .ZN(n16747) );
  INV_X1 U10457 ( .A(n15291), .ZN(n15496) );
  NAND2_X1 U10458 ( .A1(n16751), .A2(n16740), .ZN(n15517) );
  INV_X1 U10459 ( .A(n16751), .ZN(n16748) );
  NAND2_X1 U10460 ( .A1(n16148), .A2(n16147), .ZN(n16149) );
  INV_X1 U10461 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n15525) );
  INV_X1 U10462 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n10632) );
  NAND2_X1 U10463 ( .A1(n10714), .A2(P1_STATE_REG_SCAN_IN), .ZN(n16535) );
  INV_X1 U10464 ( .A(n13719), .ZN(n16694) );
  INV_X1 U10465 ( .A(n15815), .ZN(n15791) );
  NAND4_X1 U10466 ( .A1(n12885), .A2(n12884), .A3(n12883), .A4(n12882), .ZN(
        n15859) );
  OR2_X1 U10467 ( .A1(n16249), .A2(n10401), .ZN(n15727) );
  OR2_X1 U10468 ( .A1(n16249), .A2(n10022), .ZN(n15710) );
  INV_X1 U10469 ( .A(n16246), .ZN(n16267) );
  OR2_X1 U10470 ( .A1(n15918), .A2(n15917), .ZN(n16064) );
  INV_X1 U10471 ( .A(n15855), .ZN(n15947) );
  OR2_X1 U10472 ( .A1(n7414), .A2(n10936), .ZN(n15983) );
  INV_X1 U10473 ( .A(n16734), .ZN(n16732) );
  INV_X1 U10474 ( .A(n16737), .ZN(n16735) );
  AND2_X1 U10475 ( .A1(n10392), .A2(n9969), .ZN(n10878) );
  INV_X1 U10476 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n12927) );
  INV_X1 U10477 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n16140) );
  INV_X1 U10478 ( .A(n12339), .ZN(n11898) );
  INV_X1 U10479 ( .A(n10989), .ZN(P3_U3897) );
  OR4_X1 U10480 ( .A1(n9695), .A2(n9694), .A3(n9693), .A4(n9692), .ZN(P3_U3194) );
  INV_X1 U10481 ( .A(n15044), .ZN(P2_U3947) );
  NAND2_X1 U10482 ( .A1(n14535), .A2(n14474), .ZN(n9022) );
  INV_X1 U10483 ( .A(n9022), .ZN(n8860) );
  NAND2_X1 U10484 ( .A1(n8860), .A2(n14716), .ZN(n9041) );
  INV_X1 U10485 ( .A(n9058), .ZN(n8862) );
  INV_X1 U10486 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n8861) );
  NAND2_X1 U10487 ( .A1(n8862), .A2(n8861), .ZN(n9087) );
  INV_X1 U10488 ( .A(n9089), .ZN(n8864) );
  INV_X1 U10489 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n8863) );
  NAND2_X1 U10490 ( .A1(n8864), .A2(n8863), .ZN(n9108) );
  INV_X1 U10491 ( .A(n9140), .ZN(n8866) );
  INV_X1 U10492 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n8865) );
  NAND2_X1 U10493 ( .A1(n8866), .A2(n8865), .ZN(n9158) );
  INV_X1 U10494 ( .A(n9158), .ZN(n8867) );
  NAND2_X1 U10495 ( .A1(n8867), .A2(n14632), .ZN(n9182) );
  NAND2_X1 U10496 ( .A1(n9217), .A2(n14715), .ZN(n9235) );
  NAND2_X1 U10497 ( .A1(n14703), .A2(n14738), .ZN(n8868) );
  INV_X1 U10498 ( .A(P3_REG3_REG_20__SCAN_IN), .ZN(n13926) );
  NAND2_X1 U10499 ( .A1(n9273), .A2(n14641), .ZN(n9285) );
  INV_X1 U10500 ( .A(n9305), .ZN(n8869) );
  NAND2_X1 U10501 ( .A1(n8869), .A2(n14634), .ZN(n9307) );
  INV_X1 U10502 ( .A(n9307), .ZN(n8870) );
  INV_X1 U10503 ( .A(P3_REG3_REG_26__SCAN_IN), .ZN(n14739) );
  INV_X1 U10504 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n14644) );
  NAND2_X1 U10505 ( .A1(n14739), .A2(n14644), .ZN(n8871) );
  INV_X1 U10506 ( .A(n9324), .ZN(n8873) );
  INV_X1 U10507 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n8872) );
  NAND2_X1 U10508 ( .A1(n8873), .A2(n8872), .ZN(n13808) );
  NAND2_X1 U10509 ( .A1(n9324), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n8874) );
  NAND2_X1 U10510 ( .A1(n13808), .A2(n8874), .ZN(n14165) );
  NOR2_X1 U10511 ( .A1(P3_IR_REG_9__SCAN_IN), .A2(P3_IR_REG_8__SCAN_IN), .ZN(
        n8881) );
  NOR2_X1 U10512 ( .A1(P3_IR_REG_7__SCAN_IN), .A2(P3_IR_REG_11__SCAN_IN), .ZN(
        n8880) );
  NOR2_X1 U10513 ( .A1(P3_IR_REG_10__SCAN_IN), .A2(P3_IR_REG_12__SCAN_IN), 
        .ZN(n8879) );
  NAND2_X1 U10514 ( .A1(n8887), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8889) );
  INV_X1 U10515 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n8895) );
  AND2_X2 U10516 ( .A1(n8890), .A2(n14915), .ZN(n8980) );
  NAND2_X1 U10517 ( .A1(n9308), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n8894) );
  INV_X2 U10518 ( .A(n8950), .ZN(n9314) );
  INV_X1 U10519 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n8892) );
  OR2_X1 U10520 ( .A1(n9314), .A2(n8892), .ZN(n8893) );
  OAI211_X1 U10521 ( .C1(n8895), .C2(n10998), .A(n8894), .B(n8893), .ZN(n8896)
         );
  AOI22_X1 U10522 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(n8582), .B1(
        P1_DATAO_REG_23__SCAN_IN), .B2(n16140), .ZN(n9292) );
  INV_X1 U10523 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8919) );
  AOI22_X1 U10524 ( .A1(P2_DATAO_REG_22__SCAN_IN), .A2(n7827), .B1(
        P1_DATAO_REG_22__SCAN_IN), .B2(n8919), .ZN(n9281) );
  INV_X1 U10525 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n12796) );
  INV_X1 U10526 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n12958) );
  AOI22_X1 U10527 ( .A1(P2_DATAO_REG_21__SCAN_IN), .A2(n12958), .B1(
        P1_DATAO_REG_21__SCAN_IN), .B2(n12796), .ZN(n9270) );
  INV_X1 U10528 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n12970) );
  AOI22_X1 U10529 ( .A1(P2_DATAO_REG_20__SCAN_IN), .A2(n12970), .B1(
        P1_DATAO_REG_20__SCAN_IN), .B2(n12779), .ZN(n9260) );
  NOR2_X1 U10530 ( .A1(P2_DATAO_REG_19__SCAN_IN), .A2(n11889), .ZN(n8918) );
  AOI22_X1 U10531 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(n11743), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n8120), .ZN(n8940) );
  XNOR2_X1 U10532 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(P2_DATAO_REG_17__SCAN_IN), 
        .ZN(n9225) );
  XNOR2_X1 U10533 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .ZN(n9146) );
  INV_X1 U10534 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n9894) );
  NAND2_X1 U10535 ( .A1(n9894), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n8897) );
  NAND2_X1 U10536 ( .A1(n8963), .A2(n8897), .ZN(n8983) );
  INV_X1 U10537 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n10407) );
  NAND2_X1 U10538 ( .A1(n10407), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n8898) );
  NAND2_X1 U10539 ( .A1(n8983), .A2(n8898), .ZN(n8900) );
  INV_X1 U10540 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n9882) );
  NAND2_X1 U10541 ( .A1(n9882), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n8899) );
  INV_X1 U10542 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n9895) );
  AND2_X1 U10543 ( .A1(n9895), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n8901) );
  NAND2_X1 U10544 ( .A1(n10684), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n8902) );
  INV_X1 U10545 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n10705) );
  NAND2_X1 U10546 ( .A1(n10705), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n8903) );
  NAND2_X1 U10547 ( .A1(n9914), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n8905) );
  INV_X1 U10548 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n9902) );
  NAND2_X1 U10549 ( .A1(n9902), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n8904) );
  NAND2_X1 U10550 ( .A1(n8905), .A2(n8904), .ZN(n9053) );
  XNOR2_X1 U10551 ( .A(n9923), .B(P1_DATAO_REG_7__SCAN_IN), .ZN(n9065) );
  NAND2_X1 U10552 ( .A1(n9096), .A2(n9095), .ZN(n8907) );
  NAND2_X1 U10553 ( .A1(n9943), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n8906) );
  NAND2_X1 U10554 ( .A1(n8907), .A2(n8906), .ZN(n9076) );
  NAND2_X1 U10555 ( .A1(n9959), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n8908) );
  NAND2_X1 U10556 ( .A1(n9978), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n8909) );
  XNOR2_X1 U10557 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .ZN(n9134) );
  NAND2_X1 U10558 ( .A1(n9146), .A2(n9148), .ZN(n8910) );
  NAND2_X1 U10559 ( .A1(n12005), .A2(n8911), .ZN(n8912) );
  XNOR2_X1 U10560 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .ZN(n9176) );
  NAND2_X1 U10561 ( .A1(n10457), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n8913) );
  XNOR2_X1 U10562 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .ZN(n9188) );
  NAND2_X1 U10563 ( .A1(n10644), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n8914) );
  XNOR2_X1 U10564 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(P2_DATAO_REG_16__SCAN_IN), 
        .ZN(n9207) );
  INV_X1 U10565 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n8915) );
  NAND2_X1 U10566 ( .A1(n9292), .A2(n9293), .ZN(n8920) );
  NOR2_X1 U10567 ( .A1(P2_DATAO_REG_24__SCAN_IN), .A2(n8921), .ZN(n8922) );
  INV_X1 U10568 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n15537) );
  AOI22_X1 U10569 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(
        P1_DATAO_REG_25__SCAN_IN), .B1(n15537), .B2(n16131), .ZN(n8929) );
  INV_X1 U10570 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n15533) );
  AOI22_X1 U10571 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(
        P1_DATAO_REG_26__SCAN_IN), .B1(n15533), .B2(n16125), .ZN(n9312) );
  INV_X1 U10572 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n10579) );
  AOI22_X1 U10573 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(
        P1_DATAO_REG_27__SCAN_IN), .B1(n10579), .B2(n16123), .ZN(n9318) );
  AOI22_X1 U10574 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(
        P1_DATAO_REG_28__SCAN_IN), .B1(n13256), .B2(n12927), .ZN(n9333) );
  XNOR2_X1 U10575 ( .A(n9334), .B(n8594), .ZN(n14916) );
  NAND2_X1 U10576 ( .A1(n14916), .A2(n13504), .ZN(n8928) );
  OR2_X1 U10577 ( .A1(n9335), .A2(n14919), .ZN(n8927) );
  INV_X1 U10578 ( .A(n14392), .ZN(n14167) );
  INV_X1 U10579 ( .A(n8929), .ZN(n8930) );
  XNOR2_X1 U10580 ( .A(n8931), .B(n8930), .ZN(n11934) );
  NAND2_X1 U10581 ( .A1(n11934), .A2(n13504), .ZN(n8933) );
  OR2_X1 U10582 ( .A1(n9335), .A2(n14656), .ZN(n8932) );
  NAND2_X1 U10583 ( .A1(n9307), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n8934) );
  NAND2_X1 U10584 ( .A1(n9323), .A2(n8934), .ZN(n14200) );
  NAND2_X1 U10585 ( .A1(n14200), .A2(n9326), .ZN(n8939) );
  INV_X1 U10586 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n14856) );
  NAND2_X1 U10587 ( .A1(n9308), .A2(P3_REG2_REG_25__SCAN_IN), .ZN(n8936) );
  INV_X1 U10588 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n14407) );
  OR2_X1 U10589 ( .A1(n9314), .A2(n14407), .ZN(n8935) );
  OAI211_X1 U10590 ( .C1(n14856), .C2(n10998), .A(n8936), .B(n8935), .ZN(n8937) );
  INV_X1 U10591 ( .A(n8937), .ZN(n8938) );
  INV_X1 U10592 ( .A(n8940), .ZN(n8941) );
  XNOR2_X1 U10593 ( .A(n8942), .B(n8941), .ZN(n10501) );
  NAND2_X1 U10594 ( .A1(n10501), .A2(n13504), .ZN(n8949) );
  NOR2_X1 U10595 ( .A1(n9229), .A2(n9077), .ZN(n8943) );
  MUX2_X1 U10596 ( .A(n9077), .B(n8943), .S(P3_IR_REG_18__SCAN_IN), .Z(n8944)
         );
  INV_X1 U10597 ( .A(n8944), .ZN(n8946) );
  INV_X1 U10598 ( .A(n8945), .ZN(n9245) );
  NAND2_X1 U10599 ( .A1(n8946), .A2(n9245), .ZN(n14137) );
  OAI22_X1 U10600 ( .A1(n9335), .A2(n14492), .B1(n9644), .B2(n14137), .ZN(
        n8947) );
  INV_X1 U10601 ( .A(n8947), .ZN(n8948) );
  NAND2_X1 U10602 ( .A1(n8949), .A2(n8948), .ZN(n14304) );
  INV_X1 U10603 ( .A(n14304), .ZN(n14433) );
  NAND2_X1 U10604 ( .A1(n8980), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n8955) );
  INV_X1 U10605 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n14113) );
  OR2_X1 U10606 ( .A1(n10995), .A2(n14113), .ZN(n8954) );
  XNOR2_X1 U10607 ( .A(n9249), .B(n14738), .ZN(n14301) );
  OR2_X1 U10608 ( .A1(n7411), .A2(n14301), .ZN(n8953) );
  INV_X1 U10609 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n8951) );
  OR2_X1 U10610 ( .A1(n10998), .A2(n8951), .ZN(n8952) );
  INV_X1 U10611 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n11531) );
  OR2_X1 U10612 ( .A1(n9253), .A2(n11531), .ZN(n8957) );
  INV_X1 U10613 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n9592) );
  OR2_X1 U10614 ( .A1(n8979), .A2(n9592), .ZN(n8956) );
  NAND2_X1 U10615 ( .A1(n8957), .A2(n8956), .ZN(n8958) );
  INV_X1 U10616 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n8959) );
  OR2_X1 U10617 ( .A1(n10998), .A2(n8959), .ZN(n8960) );
  NAND2_X1 U10618 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), 
        .ZN(n8962) );
  INV_X1 U10619 ( .A(SI_1_), .ZN(n9861) );
  OR2_X1 U10620 ( .A1(n9335), .A2(n9861), .ZN(n8967) );
  OAI21_X1 U10621 ( .B1(n8964), .B2(n8973), .A(n8963), .ZN(n8965) );
  INV_X1 U10622 ( .A(n8965), .ZN(n9862) );
  OR2_X1 U10623 ( .A1(n13494), .A2(n9862), .ZN(n8966) );
  OAI211_X1 U10624 ( .C1(n9644), .C2(n10898), .A(n8967), .B(n8966), .ZN(n11408) );
  NAND2_X1 U10625 ( .A1(n11333), .A2(n11408), .ZN(n13361) );
  NAND2_X1 U10626 ( .A1(n8980), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n8972) );
  INV_X1 U10627 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n11306) );
  OR2_X1 U10628 ( .A1(n7411), .A2(n11306), .ZN(n8971) );
  INV_X1 U10629 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n8968) );
  OR2_X1 U10630 ( .A1(n10998), .A2(n8968), .ZN(n8970) );
  INV_X1 U10631 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n9597) );
  INV_X1 U10632 ( .A(n8973), .ZN(n8975) );
  INV_X1 U10633 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n10266) );
  NAND2_X1 U10634 ( .A1(n10266), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n8974) );
  NAND2_X1 U10635 ( .A1(n8975), .A2(n8974), .ZN(n8977) );
  INV_X2 U10636 ( .A(n9874), .ZN(n8976) );
  MUX2_X1 U10637 ( .A(n8977), .B(SI_0_), .S(n7416), .Z(n9842) );
  MUX2_X1 U10638 ( .A(P3_IR_REG_0__SCAN_IN), .B(n9842), .S(n9644), .Z(n16450)
         );
  NAND2_X1 U10639 ( .A1(n11534), .A2(n16450), .ZN(n11403) );
  NAND2_X1 U10640 ( .A1(n11333), .A2(n11530), .ZN(n8978) );
  NAND2_X1 U10641 ( .A1(n11402), .A2(n8978), .ZN(n16500) );
  INV_X1 U10642 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n16509) );
  INV_X1 U10643 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n9598) );
  OR2_X1 U10644 ( .A1(n8979), .A2(n9598), .ZN(n8981) );
  INV_X1 U10645 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n9670) );
  OR2_X1 U10646 ( .A1(n9335), .A2(SI_2_), .ZN(n8988) );
  XNOR2_X1 U10647 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(P1_DATAO_REG_2__SCAN_IN), 
        .ZN(n8982) );
  XNOR2_X1 U10648 ( .A(n8983), .B(n8982), .ZN(n9856) );
  OR2_X1 U10649 ( .A1(n13494), .A2(n9856), .ZN(n8987) );
  INV_X1 U10650 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n9077) );
  OR2_X1 U10651 ( .A1(n9644), .A2(n9671), .ZN(n8986) );
  NAND2_X1 U10652 ( .A1(n11817), .A2(n9449), .ZN(n13368) );
  NAND2_X1 U10653 ( .A1(n16500), .A2(n16499), .ZN(n8990) );
  NAND2_X1 U10654 ( .A1(n11817), .A2(n16494), .ZN(n8989) );
  NAND2_X1 U10655 ( .A1(n9354), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n8994) );
  OR2_X1 U10656 ( .A1(n7411), .A2(P3_REG3_REG_3__SCAN_IN), .ZN(n8993) );
  INV_X1 U10657 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n9603) );
  OR2_X1 U10658 ( .A1(n9314), .A2(n9603), .ZN(n8992) );
  INV_X1 U10659 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n11820) );
  OR2_X1 U10660 ( .A1(n9157), .A2(n11820), .ZN(n8991) );
  AND4_X2 U10661 ( .A1(n8994), .A2(n8993), .A3(n8992), .A4(n8991), .ZN(n11828)
         );
  OR2_X1 U10662 ( .A1(n9335), .A2(SI_3_), .ZN(n9004) );
  XNOR2_X1 U10663 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .ZN(n8996) );
  XNOR2_X1 U10664 ( .A(n8997), .B(n8996), .ZN(n9859) );
  OR2_X1 U10665 ( .A1(n13494), .A2(n9859), .ZN(n9003) );
  NAND2_X1 U10666 ( .A1(n8998), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9000) );
  INV_X1 U10667 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n8999) );
  NAND2_X1 U10668 ( .A1(n9000), .A2(n8999), .ZN(n9015) );
  OR2_X1 U10669 ( .A1(n9000), .A2(n8999), .ZN(n9001) );
  OR2_X1 U10670 ( .A1(n9644), .A2(n9652), .ZN(n9002) );
  AND3_X2 U10671 ( .A1(n9004), .A2(n9003), .A3(n9002), .ZN(n16524) );
  NAND2_X1 U10672 ( .A1(n11828), .A2(n16524), .ZN(n13370) );
  INV_X1 U10673 ( .A(n16524), .ZN(n9005) );
  NAND2_X1 U10674 ( .A1(n16496), .A2(n9005), .ZN(n13363) );
  NAND2_X1 U10675 ( .A1(n16496), .A2(n16524), .ZN(n11824) );
  NAND2_X1 U10676 ( .A1(n8950), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n9011) );
  INV_X1 U10677 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n11833) );
  OR2_X1 U10678 ( .A1(n9157), .A2(n11833), .ZN(n9010) );
  NAND2_X1 U10679 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_REG3_REG_3__SCAN_IN), 
        .ZN(n9006) );
  AND2_X1 U10680 ( .A1(n9022), .A2(n9006), .ZN(n11834) );
  OR2_X1 U10681 ( .A1(n7411), .A2(n11834), .ZN(n9009) );
  INV_X1 U10682 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n9007) );
  OR2_X1 U10683 ( .A1(n10998), .A2(n9007), .ZN(n9008) );
  OR2_X1 U10684 ( .A1(n9335), .A2(SI_4_), .ZN(n9019) );
  INV_X1 U10685 ( .A(n9012), .ZN(n9013) );
  XNOR2_X1 U10686 ( .A(n9014), .B(n9013), .ZN(n9848) );
  OR2_X1 U10687 ( .A1(n13494), .A2(n9848), .ZN(n9018) );
  NAND2_X1 U10688 ( .A1(n9015), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9016) );
  XNOR2_X1 U10689 ( .A(n9016), .B(P3_IR_REG_4__SCAN_IN), .ZN(n9847) );
  OR2_X1 U10690 ( .A1(n9644), .A2(n9847), .ZN(n9017) );
  NAND2_X1 U10691 ( .A1(n11925), .A2(n11836), .ZN(n13374) );
  INV_X1 U10692 ( .A(n11836), .ZN(n16548) );
  NAND2_X1 U10693 ( .A1(n10554), .A2(n16548), .ZN(n13375) );
  NAND2_X1 U10694 ( .A1(n13374), .A2(n13375), .ZN(n13377) );
  NAND2_X1 U10695 ( .A1(n9020), .A2(n13377), .ZN(n11832) );
  NAND2_X1 U10696 ( .A1(n10554), .A2(n11836), .ZN(n9021) );
  NAND2_X1 U10697 ( .A1(n11832), .A2(n9021), .ZN(n11921) );
  INV_X1 U10698 ( .A(n11921), .ZN(n9039) );
  NAND2_X1 U10699 ( .A1(n9354), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n9028) );
  INV_X1 U10700 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n11928) );
  OR2_X1 U10701 ( .A1(n9157), .A2(n11928), .ZN(n9027) );
  NAND2_X1 U10702 ( .A1(n9022), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n9023) );
  AND2_X1 U10703 ( .A1(n9041), .A2(n9023), .ZN(n11929) );
  OR2_X1 U10704 ( .A1(n7411), .A2(n11929), .ZN(n9026) );
  INV_X1 U10705 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n9024) );
  OR2_X1 U10706 ( .A1(n10995), .A2(n9024), .ZN(n9025) );
  OR2_X1 U10707 ( .A1(n9335), .A2(SI_5_), .ZN(n9038) );
  INV_X1 U10708 ( .A(n9029), .ZN(n9030) );
  XNOR2_X1 U10709 ( .A(n9031), .B(n9030), .ZN(n9845) );
  OR2_X1 U10710 ( .A1(n13494), .A2(n9845), .ZN(n9037) );
  NAND2_X1 U10711 ( .A1(n9032), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9033) );
  MUX2_X1 U10712 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9033), .S(
        P3_IR_REG_5__SCAN_IN), .Z(n9034) );
  INV_X1 U10713 ( .A(n9034), .ZN(n9035) );
  NOR2_X1 U10714 ( .A1(n9035), .A2(n9048), .ZN(n10925) );
  OR2_X1 U10715 ( .A1(n9644), .A2(n10925), .ZN(n9036) );
  NAND2_X1 U10716 ( .A1(n11829), .A2(n11931), .ZN(n13379) );
  INV_X1 U10717 ( .A(n11931), .ZN(n16565) );
  NAND2_X1 U10718 ( .A1(n12250), .A2(n16565), .ZN(n13380) );
  NAND2_X1 U10719 ( .A1(n9039), .A2(n8336), .ZN(n11923) );
  NAND2_X1 U10720 ( .A1(n11829), .A2(n16565), .ZN(n9040) );
  NAND2_X1 U10721 ( .A1(n9308), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n9047) );
  INV_X1 U10722 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n9616) );
  OR2_X1 U10723 ( .A1(n9314), .A2(n9616), .ZN(n9046) );
  NAND2_X1 U10724 ( .A1(n9041), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n9042) );
  AND2_X1 U10725 ( .A1(n9058), .A2(n9042), .ZN(n12246) );
  OR2_X1 U10726 ( .A1(n7411), .A2(n12246), .ZN(n9045) );
  INV_X1 U10727 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n9043) );
  OR2_X1 U10728 ( .A1(n10998), .A2(n9043), .ZN(n9044) );
  NAND4_X1 U10729 ( .A1(n9047), .A2(n9046), .A3(n9045), .A4(n9044), .ZN(n13384) );
  NOR2_X1 U10730 ( .A1(n9048), .A2(n9077), .ZN(n9049) );
  MUX2_X1 U10731 ( .A(n9077), .B(n9049), .S(P3_IR_REG_6__SCAN_IN), .Z(n9050)
         );
  INV_X1 U10732 ( .A(n9050), .ZN(n9052) );
  NAND2_X1 U10733 ( .A1(n9052), .A2(n9051), .ZN(n9855) );
  INV_X1 U10734 ( .A(SI_6_), .ZN(n9853) );
  OR2_X1 U10735 ( .A1(n9335), .A2(n9853), .ZN(n9057) );
  INV_X1 U10736 ( .A(n9053), .ZN(n9054) );
  XNOR2_X1 U10737 ( .A(n9055), .B(n9054), .ZN(n9854) );
  OR2_X1 U10738 ( .A1(n13494), .A2(n9854), .ZN(n9056) );
  OAI211_X1 U10739 ( .C1(n9644), .C2(n9855), .A(n9057), .B(n9056), .ZN(n16580)
         );
  NAND2_X1 U10740 ( .A1(n9354), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n9063) );
  INV_X1 U10741 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n9621) );
  OR2_X1 U10742 ( .A1(n9157), .A2(n9621), .ZN(n9062) );
  INV_X1 U10743 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n9620) );
  OR2_X1 U10744 ( .A1(n9314), .A2(n9620), .ZN(n9061) );
  NAND2_X1 U10745 ( .A1(n9058), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n9059) );
  AND2_X1 U10746 ( .A1(n9087), .A2(n9059), .ZN(n11945) );
  OR2_X1 U10747 ( .A1(n7411), .A2(n11945), .ZN(n9060) );
  NAND4_X1 U10748 ( .A1(n9063), .A2(n9062), .A3(n9061), .A4(n9060), .ZN(n13391) );
  NAND2_X1 U10749 ( .A1(n9051), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9064) );
  INV_X1 U10750 ( .A(n9065), .ZN(n9066) );
  XNOR2_X1 U10751 ( .A(n9067), .B(n9066), .ZN(n9850) );
  OR2_X1 U10752 ( .A1(n13494), .A2(n9850), .ZN(n9069) );
  OR2_X1 U10753 ( .A1(n9335), .A2(SI_7_), .ZN(n9068) );
  OAI211_X1 U10754 ( .C1(n11524), .C2(n9644), .A(n9069), .B(n9068), .ZN(n13390) );
  XNOR2_X1 U10755 ( .A(n13391), .B(n13390), .ZN(n13387) );
  NAND2_X1 U10756 ( .A1(n9354), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n9074) );
  INV_X1 U10757 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n9628) );
  OR2_X1 U10758 ( .A1(n9314), .A2(n9628), .ZN(n9073) );
  INV_X1 U10759 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n12046) );
  OR2_X1 U10760 ( .A1(n9157), .A2(n12046), .ZN(n9072) );
  NAND2_X1 U10761 ( .A1(n9089), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n9070) );
  AND2_X1 U10762 ( .A1(n9108), .A2(n9070), .ZN(n12302) );
  OR2_X1 U10763 ( .A1(n7411), .A2(n12302), .ZN(n9071) );
  XNOR2_X1 U10764 ( .A(n9076), .B(n7833), .ZN(n9907) );
  OR2_X1 U10765 ( .A1(n13494), .A2(n9907), .ZN(n9085) );
  OR2_X1 U10766 ( .A1(n9335), .A2(SI_9_), .ZN(n9084) );
  NOR2_X1 U10767 ( .A1(n9097), .A2(P3_IR_REG_8__SCAN_IN), .ZN(n9080) );
  NOR2_X1 U10768 ( .A1(n9080), .A2(n9077), .ZN(n9078) );
  MUX2_X1 U10769 ( .A(n9077), .B(n9078), .S(P3_IR_REG_9__SCAN_IN), .Z(n9082)
         );
  INV_X1 U10770 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n9079) );
  NAND2_X1 U10771 ( .A1(n9080), .A2(n9079), .ZN(n9116) );
  INV_X1 U10772 ( .A(n9116), .ZN(n9081) );
  NOR2_X1 U10773 ( .A1(n9082), .A2(n9081), .ZN(n9630) );
  OR2_X1 U10774 ( .A1(n9644), .A2(n9630), .ZN(n9083) );
  NAND2_X1 U10775 ( .A1(n12420), .A2(n16651), .ZN(n13402) );
  INV_X1 U10776 ( .A(n16651), .ZN(n12045) );
  NAND2_X1 U10777 ( .A1(n12287), .A2(n12045), .ZN(n13403) );
  NAND2_X1 U10778 ( .A1(n13402), .A2(n13403), .ZN(n13395) );
  NAND2_X1 U10779 ( .A1(n8980), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n9094) );
  INV_X1 U10780 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n9086) );
  OR2_X1 U10781 ( .A1(n10998), .A2(n9086), .ZN(n9093) );
  NAND2_X1 U10782 ( .A1(n9087), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n9088) );
  AND2_X1 U10783 ( .A1(n9089), .A2(n9088), .ZN(n12241) );
  OR2_X1 U10784 ( .A1(n7411), .A2(n12241), .ZN(n9092) );
  INV_X1 U10785 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n9090) );
  OR2_X1 U10786 ( .A1(n10995), .A2(n9090), .ZN(n9091) );
  XNOR2_X1 U10787 ( .A(n9096), .B(n9095), .ZN(n9879) );
  OR2_X1 U10788 ( .A1(n13494), .A2(n9879), .ZN(n9102) );
  INV_X1 U10789 ( .A(SI_8_), .ZN(n9880) );
  OR2_X1 U10790 ( .A1(n9335), .A2(n9880), .ZN(n9101) );
  NAND2_X1 U10791 ( .A1(n9097), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9099) );
  INV_X1 U10792 ( .A(P3_IR_REG_8__SCAN_IN), .ZN(n9098) );
  XNOR2_X1 U10793 ( .A(n9099), .B(n9098), .ZN(n9881) );
  OR2_X1 U10794 ( .A1(n9644), .A2(n9881), .ZN(n9100) );
  NAND2_X1 U10795 ( .A1(n12300), .A2(n16614), .ZN(n12041) );
  NAND2_X1 U10796 ( .A1(n12287), .A2(n16651), .ZN(n12283) );
  INV_X1 U10797 ( .A(n16614), .ZN(n11972) );
  NAND2_X1 U10798 ( .A1(n13396), .A2(n11972), .ZN(n9104) );
  INV_X1 U10799 ( .A(n13390), .ZN(n16595) );
  NAND2_X1 U10800 ( .A1(n13391), .A2(n16595), .ZN(n9105) );
  NAND2_X1 U10801 ( .A1(n13384), .A2(n16580), .ZN(n11937) );
  OR2_X1 U10802 ( .A1(n13534), .A2(n11937), .ZN(n11939) );
  AND2_X1 U10803 ( .A1(n9105), .A2(n11939), .ZN(n12235) );
  AND2_X1 U10804 ( .A1(n12233), .A2(n12235), .ZN(n12040) );
  OR2_X1 U10805 ( .A1(n7467), .A2(n12040), .ZN(n12038) );
  AND2_X1 U10806 ( .A1(n12283), .A2(n12038), .ZN(n9106) );
  NAND2_X1 U10807 ( .A1(n8950), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n9114) );
  INV_X1 U10808 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n9107) );
  OR2_X1 U10809 ( .A1(n9157), .A2(n9107), .ZN(n9113) );
  NAND2_X1 U10810 ( .A1(n9108), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n9109) );
  AND2_X1 U10811 ( .A1(n9126), .A2(n9109), .ZN(n12426) );
  OR2_X1 U10812 ( .A1(n7411), .A2(n12426), .ZN(n9112) );
  INV_X1 U10813 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n9110) );
  OR2_X1 U10814 ( .A1(n10998), .A2(n9110), .ZN(n9111) );
  NAND4_X1 U10815 ( .A1(n9114), .A2(n9113), .A3(n9112), .A4(n9111), .ZN(n13406) );
  NAND2_X1 U10816 ( .A1(n9116), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9115) );
  MUX2_X1 U10817 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9115), .S(
        P3_IR_REG_10__SCAN_IN), .Z(n9117) );
  NAND2_X1 U10818 ( .A1(n9117), .A2(n9149), .ZN(n9935) );
  INV_X1 U10819 ( .A(n9935), .ZN(n11963) );
  OR2_X1 U10820 ( .A1(n9335), .A2(SI_10_), .ZN(n9122) );
  INV_X1 U10821 ( .A(n9118), .ZN(n9119) );
  XNOR2_X1 U10822 ( .A(n9120), .B(n9119), .ZN(n9933) );
  OR2_X1 U10823 ( .A1(n13494), .A2(n9933), .ZN(n9121) );
  OAI211_X1 U10824 ( .C1(n11963), .C2(n9644), .A(n9122), .B(n9121), .ZN(n16663) );
  XNOR2_X1 U10825 ( .A(n13406), .B(n16663), .ZN(n12282) );
  NAND2_X1 U10826 ( .A1(n9123), .A2(n12282), .ZN(n12286) );
  INV_X1 U10827 ( .A(n16663), .ZN(n12423) );
  NAND2_X1 U10828 ( .A1(n13406), .A2(n12423), .ZN(n9124) );
  NAND2_X1 U10829 ( .A1(n9354), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n9131) );
  INV_X1 U10830 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n9125) );
  OR2_X1 U10831 ( .A1(n9157), .A2(n9125), .ZN(n9130) );
  NAND2_X1 U10832 ( .A1(n9126), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n9127) );
  AND2_X1 U10833 ( .A1(n9140), .A2(n9127), .ZN(n12583) );
  OR2_X1 U10834 ( .A1(n7411), .A2(n12583), .ZN(n9129) );
  OR2_X1 U10835 ( .A1(n9314), .A2(n16690), .ZN(n9128) );
  NAND2_X1 U10836 ( .A1(n9149), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9132) );
  XNOR2_X1 U10837 ( .A(n9132), .B(P3_IR_REG_11__SCAN_IN), .ZN(n12166) );
  OR2_X1 U10838 ( .A1(n9335), .A2(SI_11_), .ZN(n9138) );
  INV_X1 U10839 ( .A(n9134), .ZN(n9135) );
  XNOR2_X1 U10840 ( .A(n9136), .B(n9135), .ZN(n9949) );
  OR2_X1 U10841 ( .A1(n13494), .A2(n9949), .ZN(n9137) );
  OAI211_X1 U10842 ( .C1(n12166), .C2(n9644), .A(n9138), .B(n9137), .ZN(n16686) );
  NAND2_X1 U10843 ( .A1(n12419), .A2(n16686), .ZN(n9139) );
  INV_X1 U10844 ( .A(n16686), .ZN(n12580) );
  NAND2_X1 U10845 ( .A1(n9354), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n9145) );
  INV_X1 U10846 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n9590) );
  OR2_X1 U10847 ( .A1(n9157), .A2(n9590), .ZN(n9144) );
  NAND2_X1 U10848 ( .A1(n9140), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n9141) );
  AND2_X1 U10849 ( .A1(n9158), .A2(n9141), .ZN(n14383) );
  OR2_X1 U10850 ( .A1(n7411), .A2(n14383), .ZN(n9143) );
  INV_X1 U10851 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n9591) );
  OR2_X1 U10852 ( .A1(n10995), .A2(n9591), .ZN(n9142) );
  INV_X1 U10853 ( .A(n9146), .ZN(n9147) );
  XNOR2_X1 U10854 ( .A(n9148), .B(n9147), .ZN(n9951) );
  OR2_X1 U10855 ( .A1(n9951), .A2(n13494), .ZN(n9153) );
  OR2_X1 U10856 ( .A1(n9335), .A2(SI_12_), .ZN(n9152) );
  OAI21_X1 U10857 ( .B1(n9149), .B2(P3_IR_REG_11__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9150) );
  XNOR2_X1 U10858 ( .A(n9150), .B(P3_IR_REG_12__SCAN_IN), .ZN(n9647) );
  OR2_X1 U10859 ( .A1(n9644), .A2(n9647), .ZN(n9151) );
  NAND2_X1 U10860 ( .A1(n13934), .A2(n13877), .ZN(n13417) );
  INV_X1 U10861 ( .A(n13934), .ZN(n10505) );
  NAND2_X1 U10862 ( .A1(n10505), .A2(n14831), .ZN(n13418) );
  NAND2_X1 U10863 ( .A1(n13417), .A2(n13418), .ZN(n14376) );
  INV_X1 U10864 ( .A(n14376), .ZN(n13537) );
  OR2_X1 U10865 ( .A1(n13934), .A2(n14831), .ZN(n9154) );
  NAND2_X1 U10866 ( .A1(n9354), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n9163) );
  INV_X1 U10867 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n9155) );
  OR2_X1 U10868 ( .A1(n9314), .A2(n9155), .ZN(n9162) );
  INV_X1 U10869 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n9156) );
  OR2_X1 U10870 ( .A1(n9157), .A2(n9156), .ZN(n9161) );
  NAND2_X1 U10871 ( .A1(n9158), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n9159) );
  AND2_X1 U10872 ( .A1(n9182), .A2(n9159), .ZN(n13937) );
  OR2_X1 U10873 ( .A1(n7411), .A2(n13937), .ZN(n9160) );
  NAND4_X1 U10874 ( .A1(n9163), .A2(n9162), .A3(n9161), .A4(n9160), .ZN(n14379) );
  XNOR2_X1 U10875 ( .A(n9164), .B(P1_DATAO_REG_13__SCAN_IN), .ZN(n9985) );
  NAND2_X1 U10876 ( .A1(n9985), .A2(n13504), .ZN(n9173) );
  INV_X1 U10877 ( .A(n9165), .ZN(n9166) );
  NOR2_X1 U10878 ( .A1(n9051), .A2(n9166), .ZN(n9169) );
  OR2_X1 U10879 ( .A1(n9169), .A2(n9077), .ZN(n9167) );
  MUX2_X1 U10880 ( .A(n9167), .B(P3_IR_REG_31__SCAN_IN), .S(n9168), .Z(n9170)
         );
  NAND2_X1 U10881 ( .A1(n9169), .A2(n9168), .ZN(n9190) );
  OAI22_X1 U10882 ( .A1(n9335), .A2(SI_13_), .B1(n14024), .B2(n9644), .ZN(
        n9171) );
  INV_X1 U10883 ( .A(n9171), .ZN(n9172) );
  NAND2_X1 U10884 ( .A1(n9173), .A2(n9172), .ZN(n16712) );
  NAND2_X1 U10885 ( .A1(n9174), .A2(n16712), .ZN(n9175) );
  XNOR2_X1 U10886 ( .A(n9177), .B(n9176), .ZN(n10016) );
  NAND2_X1 U10887 ( .A1(n10016), .A2(n13504), .ZN(n9181) );
  NAND2_X1 U10888 ( .A1(n9190), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9178) );
  XNOR2_X1 U10889 ( .A(n9178), .B(n9191), .ZN(n14046) );
  INV_X1 U10890 ( .A(n14046), .ZN(n14033) );
  OAI22_X1 U10891 ( .A1(n9335), .A2(SI_14_), .B1(n14033), .B2(n9644), .ZN(
        n9179) );
  INV_X1 U10892 ( .A(n9179), .ZN(n9180) );
  NAND2_X1 U10893 ( .A1(n9308), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n9187) );
  INV_X1 U10894 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n14453) );
  OR2_X1 U10895 ( .A1(n9314), .A2(n14453), .ZN(n9186) );
  NAND2_X1 U10896 ( .A1(n9182), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n9183) );
  AND2_X1 U10897 ( .A1(n9197), .A2(n9183), .ZN(n13837) );
  OR2_X1 U10898 ( .A1(n7411), .A2(n13837), .ZN(n9185) );
  INV_X1 U10899 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n14893) );
  OR2_X1 U10900 ( .A1(n10998), .A2(n14893), .ZN(n9184) );
  NAND4_X1 U10901 ( .A1(n9187), .A2(n9186), .A3(n9185), .A4(n9184), .ZN(n14347) );
  OR2_X1 U10902 ( .A1(n14895), .A2(n14347), .ZN(n13426) );
  NAND2_X1 U10903 ( .A1(n14895), .A2(n14347), .ZN(n13427) );
  XNOR2_X1 U10904 ( .A(n9189), .B(n9188), .ZN(n10123) );
  NAND2_X1 U10905 ( .A1(n10123), .A2(n13504), .ZN(n9196) );
  INV_X1 U10906 ( .A(n9190), .ZN(n9192) );
  NAND2_X1 U10907 ( .A1(n9192), .A2(n9191), .ZN(n9210) );
  NAND2_X1 U10908 ( .A1(n9210), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9193) );
  XNOR2_X1 U10909 ( .A(n9193), .B(P3_IR_REG_15__SCAN_IN), .ZN(n14063) );
  OAI22_X1 U10910 ( .A1(n9335), .A2(SI_15_), .B1(n14063), .B2(n9644), .ZN(
        n9194) );
  INV_X1 U10911 ( .A(n9194), .ZN(n9195) );
  NAND2_X1 U10912 ( .A1(n9196), .A2(n9195), .ZN(n14445) );
  NAND2_X1 U10913 ( .A1(n8980), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n9202) );
  INV_X1 U10914 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n14449) );
  OR2_X1 U10915 ( .A1(n9314), .A2(n14449), .ZN(n9201) );
  AND2_X1 U10916 ( .A1(n9197), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n9198) );
  NOR2_X1 U10917 ( .A1(n9217), .A2(n9198), .ZN(n14351) );
  OR2_X1 U10918 ( .A1(n7411), .A2(n14351), .ZN(n9200) );
  INV_X1 U10919 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n14889) );
  OR2_X1 U10920 ( .A1(n10998), .A2(n14889), .ZN(n9199) );
  NAND4_X1 U10921 ( .A1(n9202), .A2(n9201), .A3(n9200), .A4(n9199), .ZN(n14363) );
  INV_X1 U10922 ( .A(n14363), .ZN(n9469) );
  AND2_X1 U10923 ( .A1(n14445), .A2(n9469), .ZN(n9204) );
  OR2_X1 U10924 ( .A1(n14366), .A2(n9204), .ZN(n9203) );
  NOR2_X1 U10925 ( .A1(n14359), .A2(n9203), .ZN(n9206) );
  OR2_X1 U10926 ( .A1(n14445), .A2(n14363), .ZN(n14330) );
  NAND2_X1 U10927 ( .A1(n14445), .A2(n14363), .ZN(n13429) );
  NAND2_X1 U10928 ( .A1(n14330), .A2(n13429), .ZN(n14344) );
  INV_X1 U10929 ( .A(n14347), .ZN(n12570) );
  OR2_X1 U10930 ( .A1(n14895), .A2(n12570), .ZN(n14341) );
  AND2_X1 U10931 ( .A1(n14344), .A2(n14341), .ZN(n14342) );
  NOR2_X1 U10932 ( .A1(n9204), .A2(n14342), .ZN(n9205) );
  NOR2_X1 U10933 ( .A1(n9206), .A2(n9205), .ZN(n14327) );
  INV_X1 U10934 ( .A(n9207), .ZN(n9208) );
  XNOR2_X1 U10935 ( .A(n9209), .B(n9208), .ZN(n10237) );
  NAND2_X1 U10936 ( .A1(n10237), .A2(n13504), .ZN(n9215) );
  OAI21_X1 U10937 ( .B1(n9210), .B2(P3_IR_REG_15__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9212) );
  INV_X1 U10938 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n9211) );
  XNOR2_X1 U10939 ( .A(n9212), .B(n9211), .ZN(n14083) );
  OAI22_X1 U10940 ( .A1(n9335), .A2(n11160), .B1(n9644), .B2(n14083), .ZN(
        n9213) );
  INV_X1 U10941 ( .A(n9213), .ZN(n9214) );
  NAND2_X1 U10942 ( .A1(n9215), .A2(n9214), .ZN(n14441) );
  NAND2_X1 U10943 ( .A1(n9308), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n9223) );
  INV_X1 U10944 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n9216) );
  OR2_X1 U10945 ( .A1(n9314), .A2(n9216), .ZN(n9222) );
  OR2_X1 U10946 ( .A1(n9217), .A2(n14715), .ZN(n9218) );
  AND2_X1 U10947 ( .A1(n9235), .A2(n9218), .ZN(n14335) );
  OR2_X1 U10948 ( .A1(n7411), .A2(n14335), .ZN(n9221) );
  INV_X1 U10949 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n9219) );
  OR2_X1 U10950 ( .A1(n10998), .A2(n9219), .ZN(n9220) );
  XNOR2_X1 U10951 ( .A(n14441), .B(n14311), .ZN(n14326) );
  NOR2_X1 U10952 ( .A1(n14441), .A2(n14348), .ZN(n9224) );
  XNOR2_X1 U10953 ( .A(n9226), .B(n9225), .ZN(n10289) );
  NAND2_X1 U10954 ( .A1(n10289), .A2(n13504), .ZN(n9234) );
  NAND2_X1 U10955 ( .A1(n9227), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9228) );
  MUX2_X1 U10956 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9228), .S(
        P3_IR_REG_17__SCAN_IN), .Z(n9231) );
  INV_X1 U10957 ( .A(n9229), .ZN(n9230) );
  NAND2_X1 U10958 ( .A1(n9231), .A2(n9230), .ZN(n14108) );
  INV_X1 U10959 ( .A(n14108), .ZN(n14098) );
  OAI22_X1 U10960 ( .A1(n9335), .A2(SI_17_), .B1(n14098), .B2(n9644), .ZN(
        n9232) );
  INV_X1 U10961 ( .A(n9232), .ZN(n9233) );
  NAND2_X1 U10962 ( .A1(n9308), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n9240) );
  INV_X1 U10963 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n14884) );
  OR2_X1 U10964 ( .A1(n10998), .A2(n14884), .ZN(n9239) );
  NAND2_X1 U10965 ( .A1(n9235), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n9236) );
  AND2_X1 U10966 ( .A1(n9249), .A2(n9236), .ZN(n14321) );
  OR2_X1 U10967 ( .A1(n7411), .A2(n14321), .ZN(n9238) );
  INV_X1 U10968 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n14439) );
  OR2_X1 U10969 ( .A1(n10995), .A2(n14439), .ZN(n9237) );
  NAND4_X1 U10970 ( .A1(n9240), .A2(n9239), .A3(n9238), .A4(n9237), .ZN(n14328) );
  XNOR2_X1 U10971 ( .A(n14886), .B(n14328), .ZN(n14307) );
  INV_X1 U10972 ( .A(n14328), .ZN(n13905) );
  NOR2_X1 U10973 ( .A1(n14886), .A2(n13905), .ZN(n9241) );
  OR2_X1 U10974 ( .A1(n14304), .A2(n14313), .ZN(n13438) );
  NAND2_X1 U10975 ( .A1(n14304), .A2(n14313), .ZN(n14280) );
  NAND2_X1 U10976 ( .A1(n13438), .A2(n14280), .ZN(n14293) );
  AOI22_X1 U10977 ( .A1(P2_DATAO_REG_19__SCAN_IN), .A2(
        P1_DATAO_REG_19__SCAN_IN), .B1(n11889), .B2(n11887), .ZN(n9242) );
  XNOR2_X1 U10978 ( .A(n9243), .B(n9242), .ZN(n10675) );
  NAND2_X1 U10979 ( .A1(n9245), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9246) );
  MUX2_X1 U10980 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9246), .S(
        P3_IR_REG_19__SCAN_IN), .Z(n9247) );
  OAI22_X1 U10981 ( .A1(n9335), .A2(n14666), .B1(n9644), .B2(n14132), .ZN(
        n9248) );
  NAND2_X1 U10982 ( .A1(n8980), .A2(P3_REG2_REG_19__SCAN_IN), .ZN(n9257) );
  INV_X1 U10983 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n14431) );
  OR2_X1 U10984 ( .A1(n9314), .A2(n14431), .ZN(n9256) );
  OAI21_X1 U10985 ( .B1(n9249), .B2(P3_REG3_REG_18__SCAN_IN), .A(
        P3_REG3_REG_19__SCAN_IN), .ZN(n9250) );
  INV_X1 U10986 ( .A(n9250), .ZN(n9251) );
  OR2_X1 U10987 ( .A1(n9251), .A2(n9264), .ZN(n14287) );
  INV_X1 U10988 ( .A(n14287), .ZN(n9252) );
  OR2_X1 U10989 ( .A1(n7411), .A2(n9252), .ZN(n9255) );
  INV_X1 U10990 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n14879) );
  OR2_X1 U10991 ( .A1(n10998), .A2(n14879), .ZN(n9254) );
  NAND2_X1 U10992 ( .A1(n14881), .A2(n14264), .ZN(n9259) );
  NOR2_X1 U10993 ( .A1(n14881), .A2(n14264), .ZN(n9258) );
  XNOR2_X1 U10994 ( .A(n9261), .B(n9260), .ZN(n10785) );
  NAND2_X1 U10995 ( .A1(n10785), .A2(n13504), .ZN(n9263) );
  OR2_X1 U10996 ( .A1(n9335), .A2(n14664), .ZN(n9262) );
  NAND2_X1 U10997 ( .A1(n9308), .A2(P3_REG2_REG_20__SCAN_IN), .ZN(n9269) );
  NOR2_X1 U10998 ( .A1(n9264), .A2(n13926), .ZN(n9265) );
  OR2_X1 U10999 ( .A1(n9273), .A2(n9265), .ZN(n13929) );
  INV_X1 U11000 ( .A(n13929), .ZN(n14269) );
  OR2_X1 U11001 ( .A1(n14269), .A2(n7411), .ZN(n9268) );
  INV_X1 U11002 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n14427) );
  OR2_X1 U11003 ( .A1(n9314), .A2(n14427), .ZN(n9267) );
  INV_X1 U11004 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n14875) );
  OR2_X1 U11005 ( .A1(n10998), .A2(n14875), .ZN(n9266) );
  OR2_X1 U11006 ( .A1(n14272), .A2(n14278), .ZN(n13451) );
  NAND2_X1 U11007 ( .A1(n14272), .A2(n14278), .ZN(n13452) );
  XOR2_X1 U11008 ( .A(n9271), .B(n9270), .Z(n10834) );
  INV_X1 U11009 ( .A(SI_21_), .ZN(n14662) );
  OR2_X1 U11010 ( .A1(n9335), .A2(n14662), .ZN(n9272) );
  OAI21_X1 U11011 ( .B1(n10834), .B2(n13494), .A(n9272), .ZN(n14253) );
  INV_X1 U11012 ( .A(n14253), .ZN(n14873) );
  OR2_X1 U11013 ( .A1(n9273), .A2(n14641), .ZN(n9274) );
  AND2_X1 U11014 ( .A1(n9285), .A2(n9274), .ZN(n14250) );
  INV_X1 U11015 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n14423) );
  OR2_X1 U11016 ( .A1(n10995), .A2(n14423), .ZN(n9275) );
  OAI21_X1 U11017 ( .B1(n14250), .B2(n7411), .A(n9275), .ZN(n9276) );
  INV_X1 U11018 ( .A(n9276), .ZN(n9280) );
  NAND2_X1 U11019 ( .A1(n9308), .A2(P3_REG2_REG_21__SCAN_IN), .ZN(n9278) );
  INV_X1 U11020 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n14871) );
  OR2_X1 U11021 ( .A1(n10998), .A2(n14871), .ZN(n9277) );
  AND2_X1 U11022 ( .A1(n9278), .A2(n9277), .ZN(n9279) );
  NOR2_X1 U11023 ( .A1(n14873), .A2(n14265), .ZN(n9497) );
  INV_X1 U11024 ( .A(n14265), .ZN(n14233) );
  OR2_X1 U11025 ( .A1(n14253), .A2(n14233), .ZN(n9498) );
  XNOR2_X1 U11026 ( .A(n9282), .B(n9281), .ZN(n10960) );
  NAND2_X1 U11027 ( .A1(n10960), .A2(n13504), .ZN(n9284) );
  OR2_X1 U11028 ( .A1(n9335), .A2(n14655), .ZN(n9283) );
  NAND2_X1 U11029 ( .A1(n9285), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n9286) );
  NAND2_X1 U11030 ( .A1(n9296), .A2(n9286), .ZN(n14237) );
  NAND2_X1 U11031 ( .A1(n9287), .A2(n14237), .ZN(n9291) );
  INV_X1 U11032 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n14419) );
  OR2_X1 U11033 ( .A1(n10995), .A2(n14419), .ZN(n9290) );
  NAND2_X1 U11034 ( .A1(n9308), .A2(P3_REG2_REG_22__SCAN_IN), .ZN(n9289) );
  INV_X1 U11035 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n14867) );
  OR2_X1 U11036 ( .A1(n10998), .A2(n14867), .ZN(n9288) );
  NAND4_X1 U11037 ( .A1(n9291), .A2(n9290), .A3(n9289), .A4(n9288), .ZN(n14246) );
  NAND2_X1 U11038 ( .A1(n13942), .A2(n14246), .ZN(n13457) );
  NOR2_X1 U11039 ( .A1(n13942), .A2(n14246), .ZN(n13459) );
  XNOR2_X1 U11040 ( .A(n9293), .B(n9292), .ZN(n11356) );
  NAND2_X1 U11041 ( .A1(n11356), .A2(n13504), .ZN(n9295) );
  OR2_X1 U11042 ( .A1(n9335), .A2(n12618), .ZN(n9294) );
  INV_X1 U11043 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n14863) );
  NAND2_X1 U11044 ( .A1(n9296), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n9297) );
  NAND2_X1 U11045 ( .A1(n9305), .A2(n9297), .ZN(n14223) );
  NAND2_X1 U11046 ( .A1(n14223), .A2(n9326), .ZN(n9301) );
  NAND2_X1 U11047 ( .A1(n8980), .A2(P3_REG2_REG_23__SCAN_IN), .ZN(n9299) );
  INV_X1 U11048 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n14415) );
  OR2_X1 U11049 ( .A1(n9314), .A2(n14415), .ZN(n9298) );
  AND2_X1 U11050 ( .A1(n9299), .A2(n9298), .ZN(n9300) );
  OAI211_X1 U11051 ( .C1(n10998), .C2(n14863), .A(n9301), .B(n9300), .ZN(
        n14232) );
  XNOR2_X1 U11052 ( .A(n13847), .B(n14232), .ZN(n14221) );
  INV_X1 U11053 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n15541) );
  XNOR2_X1 U11054 ( .A(n15541), .B(n9302), .ZN(n13830) );
  NAND2_X1 U11055 ( .A1(n13830), .A2(n13504), .ZN(n9304) );
  INV_X1 U11056 ( .A(SI_24_), .ZN(n13832) );
  OR2_X1 U11057 ( .A1(n9335), .A2(n13832), .ZN(n9303) );
  INV_X1 U11058 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n14859) );
  NAND2_X1 U11059 ( .A1(n9305), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n9306) );
  NAND2_X1 U11060 ( .A1(n9307), .A2(n9306), .ZN(n14211) );
  NAND2_X1 U11061 ( .A1(n14211), .A2(n9326), .ZN(n9310) );
  AOI22_X1 U11062 ( .A1(n8950), .A2(P3_REG1_REG_24__SCAN_IN), .B1(n9308), .B2(
        P3_REG2_REG_24__SCAN_IN), .ZN(n9309) );
  OAI211_X1 U11063 ( .C1(n10998), .C2(n14859), .A(n9310), .B(n9309), .ZN(
        n14195) );
  NAND2_X1 U11064 ( .A1(n13470), .A2(n14195), .ZN(n9311) );
  INV_X1 U11065 ( .A(n14195), .ZN(n14220) );
  AOI22_X1 U11066 ( .A1(n14206), .A2(n9311), .B1(n14220), .B2(n14861), .ZN(
        n14194) );
  XNOR2_X1 U11067 ( .A(n9510), .B(n14209), .ZN(n14193) );
  XNOR2_X1 U11068 ( .A(n9313), .B(n8596), .ZN(n12292) );
  INV_X1 U11069 ( .A(SI_26_), .ZN(n14483) );
  XNOR2_X1 U11070 ( .A(n9323), .B(P3_REG3_REG_26__SCAN_IN), .ZN(n14187) );
  INV_X1 U11071 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n14852) );
  NAND2_X1 U11072 ( .A1(n8980), .A2(P3_REG2_REG_26__SCAN_IN), .ZN(n9316) );
  INV_X1 U11073 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n14403) );
  OR2_X1 U11074 ( .A1(n9314), .A2(n14403), .ZN(n9315) );
  OAI211_X1 U11075 ( .C1(n14852), .C2(n10998), .A(n9316), .B(n9315), .ZN(n9317) );
  INV_X1 U11076 ( .A(n9318), .ZN(n9319) );
  XNOR2_X1 U11077 ( .A(n9320), .B(n9319), .ZN(n13562) );
  NAND2_X1 U11078 ( .A1(n13562), .A2(n13504), .ZN(n9322) );
  INV_X1 U11079 ( .A(SI_27_), .ZN(n14477) );
  OAI21_X1 U11080 ( .B1(n9323), .B2(P3_REG3_REG_26__SCAN_IN), .A(
        P3_REG3_REG_27__SCAN_IN), .ZN(n9325) );
  NAND2_X1 U11081 ( .A1(n9325), .A2(n9324), .ZN(n14178) );
  NAND2_X1 U11082 ( .A1(n14178), .A2(n9326), .ZN(n9332) );
  INV_X1 U11083 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n9329) );
  NAND2_X1 U11084 ( .A1(n8980), .A2(P3_REG2_REG_27__SCAN_IN), .ZN(n9328) );
  INV_X1 U11085 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n14397) );
  OR2_X1 U11086 ( .A1(n10995), .A2(n14397), .ZN(n9327) );
  OAI211_X1 U11087 ( .C1(n9329), .C2(n10998), .A(n9328), .B(n9327), .ZN(n9330)
         );
  INV_X1 U11088 ( .A(n9330), .ZN(n9331) );
  NAND2_X1 U11089 ( .A1(n9448), .A2(n14184), .ZN(n13477) );
  NAND2_X1 U11090 ( .A1(n13478), .A2(n13477), .ZN(n14173) );
  OR2_X1 U11091 ( .A1(n14392), .A2(n11040), .ZN(n13356) );
  NAND2_X1 U11092 ( .A1(n14392), .A2(n11040), .ZN(n13355) );
  INV_X1 U11093 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n13600) );
  OAI22_X1 U11094 ( .A1(n13600), .A2(P1_DATAO_REG_29__SCAN_IN), .B1(n13493), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n13492) );
  NOR2_X1 U11095 ( .A1(n9335), .A2(n14914), .ZN(n9336) );
  INV_X1 U11096 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n9340) );
  NAND2_X1 U11097 ( .A1(n8980), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n9339) );
  INV_X1 U11098 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n9337) );
  OR2_X1 U11099 ( .A1(n10995), .A2(n9337), .ZN(n9338) );
  OAI211_X1 U11100 ( .C1(n10998), .C2(n9340), .A(n9339), .B(n9338), .ZN(n9341)
         );
  INV_X1 U11101 ( .A(n9341), .ZN(n9342) );
  NAND2_X1 U11102 ( .A1(n11002), .A2(n9342), .ZN(n10963) );
  NOR2_X1 U11103 ( .A1(n13810), .A2(n10963), .ZN(n13489) );
  INV_X1 U11104 ( .A(n13810), .ZN(n9343) );
  INV_X1 U11105 ( .A(n10963), .ZN(n14158) );
  INV_X1 U11106 ( .A(n9344), .ZN(n9346) );
  NAND2_X1 U11107 ( .A1(n13557), .A2(n14147), .ZN(n9417) );
  NAND2_X1 U11108 ( .A1(n9346), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9347) );
  MUX2_X1 U11109 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9347), .S(
        P3_IR_REG_21__SCAN_IN), .Z(n9349) );
  NAND2_X1 U11110 ( .A1(n9244), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9350) );
  INV_X1 U11111 ( .A(n10787), .ZN(n9416) );
  NAND2_X1 U11112 ( .A1(n13357), .A2(n9416), .ZN(n13517) );
  AOI22_X1 U11113 ( .A1(n8950), .A2(P3_REG1_REG_30__SCAN_IN), .B1(n8980), .B2(
        P3_REG2_REG_30__SCAN_IN), .ZN(n9351) );
  INV_X1 U11114 ( .A(n9351), .ZN(n9353) );
  INV_X1 U11115 ( .A(n11002), .ZN(n9352) );
  AOI211_X1 U11116 ( .C1(n9354), .C2(P3_REG0_REG_30__SCAN_IN), .A(n9353), .B(
        n9352), .ZN(n13507) );
  INV_X1 U11117 ( .A(n14921), .ZN(n9355) );
  NAND2_X1 U11118 ( .A1(n9355), .A2(n13555), .ZN(n9667) );
  INV_X1 U11119 ( .A(n9534), .ZN(n9535) );
  INV_X1 U11120 ( .A(P3_B_REG_SCAN_IN), .ZN(n9356) );
  OR2_X1 U11121 ( .A1(n14921), .A2(n9356), .ZN(n9357) );
  NAND2_X1 U11122 ( .A1(n16495), .A2(n9357), .ZN(n14149) );
  OAI22_X1 U11123 ( .A1(n13507), .A2(n14149), .B1(n11040), .B2(n14312), .ZN(
        n9358) );
  INV_X1 U11124 ( .A(n11534), .ZN(n11404) );
  NAND2_X1 U11125 ( .A1(n11404), .A2(n16450), .ZN(n11400) );
  NAND2_X1 U11126 ( .A1(n11400), .A2(n13361), .ZN(n9359) );
  INV_X1 U11127 ( .A(n13377), .ZN(n13522) );
  NAND2_X1 U11128 ( .A1(n11823), .A2(n13522), .ZN(n9360) );
  INV_X1 U11129 ( .A(n13384), .ZN(n11842) );
  NAND2_X1 U11130 ( .A1(n11842), .A2(n16580), .ZN(n13385) );
  NAND2_X1 U11131 ( .A1(n11944), .A2(n13534), .ZN(n9361) );
  INV_X1 U11132 ( .A(n13391), .ZN(n12240) );
  NAND2_X1 U11133 ( .A1(n12240), .A2(n16595), .ZN(n13392) );
  INV_X1 U11134 ( .A(n12233), .ZN(n13524) );
  NAND2_X1 U11135 ( .A1(n12234), .A2(n13524), .ZN(n9362) );
  NAND2_X1 U11136 ( .A1(n12300), .A2(n11972), .ZN(n13398) );
  NAND2_X1 U11137 ( .A1(n9362), .A2(n13398), .ZN(n12049) );
  NAND2_X1 U11138 ( .A1(n12577), .A2(n12423), .ZN(n13407) );
  NAND2_X1 U11139 ( .A1(n12419), .A2(n12580), .ZN(n13416) );
  NAND2_X1 U11140 ( .A1(n14380), .A2(n16686), .ZN(n13412) );
  NAND2_X1 U11141 ( .A1(n12391), .A2(n13533), .ZN(n9363) );
  NAND2_X1 U11142 ( .A1(n9363), .A2(n13416), .ZN(n14375) );
  NAND2_X1 U11143 ( .A1(n14375), .A2(n13418), .ZN(n9364) );
  NAND2_X1 U11144 ( .A1(n9364), .A2(n13417), .ZN(n12567) );
  NAND2_X1 U11145 ( .A1(n16712), .A2(n14379), .ZN(n9466) );
  NAND2_X1 U11146 ( .A1(n12567), .A2(n9466), .ZN(n9365) );
  OR2_X1 U11147 ( .A1(n16712), .A2(n14379), .ZN(n13425) );
  INV_X1 U11148 ( .A(n13426), .ZN(n9366) );
  INV_X1 U11149 ( .A(n14441), .ZN(n14334) );
  NAND2_X1 U11150 ( .A1(n14334), .A2(n14348), .ZN(n13434) );
  INV_X1 U11151 ( .A(n13434), .ZN(n9369) );
  OR2_X1 U11152 ( .A1(n14344), .A2(n9369), .ZN(n14316) );
  OR2_X1 U11153 ( .A1(n14316), .A2(n14307), .ZN(n9367) );
  NAND2_X1 U11154 ( .A1(n14441), .A2(n14311), .ZN(n13435) );
  AND2_X1 U11155 ( .A1(n14330), .A2(n13435), .ZN(n9368) );
  OR2_X1 U11156 ( .A1(n9369), .A2(n9368), .ZN(n14317) );
  OR2_X1 U11157 ( .A1(n14307), .A2(n14317), .ZN(n9370) );
  OR2_X1 U11158 ( .A1(n14886), .A2(n14328), .ZN(n14257) );
  INV_X1 U11159 ( .A(n14262), .ZN(n9373) );
  INV_X1 U11160 ( .A(n14881), .ZN(n9371) );
  NAND2_X1 U11161 ( .A1(n9371), .A2(n14264), .ZN(n13446) );
  INV_X1 U11162 ( .A(n14285), .ZN(n9372) );
  OR2_X1 U11163 ( .A1(n9372), .A2(n14280), .ZN(n14282) );
  AND2_X1 U11164 ( .A1(n13446), .A2(n14282), .ZN(n14260) );
  OR2_X1 U11165 ( .A1(n9373), .A2(n14260), .ZN(n9375) );
  AND2_X1 U11166 ( .A1(n14257), .A2(n9375), .ZN(n9374) );
  NAND2_X1 U11167 ( .A1(n14258), .A2(n9374), .ZN(n9379) );
  INV_X1 U11168 ( .A(n9375), .ZN(n9377) );
  INV_X1 U11169 ( .A(n14293), .ZN(n14279) );
  AND2_X1 U11170 ( .A1(n14279), .A2(n14285), .ZN(n14259) );
  AND2_X1 U11171 ( .A1(n14259), .A2(n14262), .ZN(n9376) );
  OR2_X1 U11172 ( .A1(n9377), .A2(n9376), .ZN(n9378) );
  NAND2_X1 U11173 ( .A1(n9379), .A2(n9378), .ZN(n9380) );
  NAND2_X1 U11174 ( .A1(n9380), .A2(n13452), .ZN(n14243) );
  OR2_X1 U11175 ( .A1(n14253), .A2(n14265), .ZN(n13456) );
  NAND2_X1 U11176 ( .A1(n14253), .A2(n14265), .ZN(n13455) );
  INV_X1 U11177 ( .A(n13455), .ZN(n9381) );
  AOI21_X1 U11178 ( .B1(n14243), .B2(n14245), .A(n9381), .ZN(n14228) );
  INV_X1 U11179 ( .A(n14246), .ZN(n14219) );
  NOR2_X1 U11180 ( .A1(n13942), .A2(n14219), .ZN(n13464) );
  NAND2_X1 U11181 ( .A1(n13942), .A2(n14219), .ZN(n13462) );
  OAI21_X2 U11182 ( .B1(n14228), .B2(n13464), .A(n13462), .ZN(n14222) );
  INV_X1 U11183 ( .A(n14232), .ZN(n14208) );
  NAND2_X1 U11184 ( .A1(n14861), .A2(n14195), .ZN(n9383) );
  NAND2_X1 U11185 ( .A1(n13470), .A2(n14220), .ZN(n9382) );
  INV_X1 U11186 ( .A(n9383), .ZN(n13484) );
  NAND2_X1 U11187 ( .A1(n9384), .A2(n14198), .ZN(n13473) );
  NAND2_X1 U11188 ( .A1(n14171), .A2(n7851), .ZN(n14170) );
  NAND2_X1 U11189 ( .A1(n14170), .A2(n13477), .ZN(n14164) );
  XNOR2_X1 U11190 ( .A(n13513), .B(n13520), .ZN(n13812) );
  NAND2_X1 U11191 ( .A1(n10835), .A2(n10787), .ZN(n9433) );
  XNOR2_X1 U11192 ( .A(n13557), .B(n9433), .ZN(n9386) );
  NAND2_X1 U11193 ( .A1(n10835), .A2(n14132), .ZN(n9385) );
  NAND2_X1 U11194 ( .A1(n9386), .A2(n9385), .ZN(n9528) );
  NAND2_X1 U11195 ( .A1(n10787), .A2(n14132), .ZN(n9432) );
  INV_X1 U11196 ( .A(n9432), .ZN(n13554) );
  NAND2_X1 U11197 ( .A1(n9434), .A2(n10835), .ZN(n16711) );
  NAND3_X1 U11198 ( .A1(n9528), .A2(n13554), .A3(n16711), .ZN(n9387) );
  NAND2_X1 U11199 ( .A1(n9417), .A2(n9432), .ZN(n9435) );
  XNOR2_X1 U11200 ( .A(n13831), .B(P3_B_REG_SCAN_IN), .ZN(n9399) );
  NAND2_X1 U11201 ( .A1(n9395), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9396) );
  MUX2_X1 U11202 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9396), .S(
        P3_IR_REG_26__SCAN_IN), .Z(n9398) );
  INV_X1 U11203 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n9400) );
  NAND2_X1 U11204 ( .A1(n10319), .A2(n9400), .ZN(n9402) );
  NAND2_X1 U11205 ( .A1(n13831), .A2(n12294), .ZN(n9401) );
  NAND2_X1 U11206 ( .A1(n10319), .A2(n9403), .ZN(n9405) );
  NAND2_X1 U11207 ( .A1(n11935), .A2(n12294), .ZN(n9404) );
  NOR2_X1 U11208 ( .A1(P3_D_REG_31__SCAN_IN), .A2(P3_D_REG_30__SCAN_IN), .ZN(
        n9409) );
  NOR4_X1 U11209 ( .A1(P3_D_REG_4__SCAN_IN), .A2(P3_D_REG_3__SCAN_IN), .A3(
        P3_D_REG_29__SCAN_IN), .A4(P3_D_REG_28__SCAN_IN), .ZN(n9408) );
  NOR4_X1 U11210 ( .A1(P3_D_REG_23__SCAN_IN), .A2(P3_D_REG_22__SCAN_IN), .A3(
        P3_D_REG_21__SCAN_IN), .A4(P3_D_REG_20__SCAN_IN), .ZN(n9407) );
  NOR4_X1 U11211 ( .A1(P3_D_REG_27__SCAN_IN), .A2(P3_D_REG_26__SCAN_IN), .A3(
        P3_D_REG_25__SCAN_IN), .A4(P3_D_REG_24__SCAN_IN), .ZN(n9406) );
  NAND4_X1 U11212 ( .A1(n9409), .A2(n9408), .A3(n9407), .A4(n9406), .ZN(n9415)
         );
  NOR4_X1 U11213 ( .A1(P3_D_REG_15__SCAN_IN), .A2(P3_D_REG_14__SCAN_IN), .A3(
        P3_D_REG_13__SCAN_IN), .A4(P3_D_REG_12__SCAN_IN), .ZN(n9413) );
  NOR4_X1 U11214 ( .A1(P3_D_REG_17__SCAN_IN), .A2(P3_D_REG_19__SCAN_IN), .A3(
        P3_D_REG_18__SCAN_IN), .A4(P3_D_REG_16__SCAN_IN), .ZN(n9412) );
  NOR4_X1 U11215 ( .A1(P3_D_REG_7__SCAN_IN), .A2(P3_D_REG_6__SCAN_IN), .A3(
        P3_D_REG_5__SCAN_IN), .A4(P3_D_REG_2__SCAN_IN), .ZN(n9411) );
  NOR4_X1 U11216 ( .A1(P3_D_REG_11__SCAN_IN), .A2(P3_D_REG_10__SCAN_IN), .A3(
        P3_D_REG_9__SCAN_IN), .A4(P3_D_REG_8__SCAN_IN), .ZN(n9410) );
  NAND4_X1 U11217 ( .A1(n9413), .A2(n9412), .A3(n9411), .A4(n9410), .ZN(n9414)
         );
  OAI21_X1 U11218 ( .B1(n9415), .B2(n9414), .A(n10319), .ZN(n9428) );
  NAND3_X1 U11219 ( .A1(n14900), .A2(n11008), .A3(n9428), .ZN(n9529) );
  OR2_X1 U11220 ( .A1(n13491), .A2(n9432), .ZN(n10789) );
  NAND2_X1 U11221 ( .A1(n10835), .A2(n9416), .ZN(n13549) );
  OR2_X1 U11222 ( .A1(n13549), .A2(n9417), .ZN(n9525) );
  AND2_X1 U11223 ( .A1(n10789), .A2(n9525), .ZN(n9420) );
  OR2_X1 U11224 ( .A1(n9418), .A2(n11008), .ZN(n9533) );
  INV_X1 U11225 ( .A(n9528), .ZN(n9419) );
  OAI22_X1 U11226 ( .A1(n9529), .A2(n9420), .B1(n9533), .B2(n9419), .ZN(n9425)
         );
  INV_X1 U11227 ( .A(n11935), .ZN(n9422) );
  NAND2_X1 U11228 ( .A1(n9442), .A2(n14891), .ZN(n9427) );
  NAND2_X1 U11229 ( .A1(n14891), .A2(n16652), .ZN(n14896) );
  NAND2_X1 U11230 ( .A1(n16719), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n9426) );
  NAND2_X1 U11231 ( .A1(n9427), .A2(n8840), .ZN(P3_U3456) );
  AND2_X1 U11232 ( .A1(n9428), .A2(n11012), .ZN(n9429) );
  INV_X1 U11233 ( .A(n11008), .ZN(n9439) );
  NAND2_X1 U11234 ( .A1(n9431), .A2(n13491), .ZN(n11006) );
  NAND2_X1 U11235 ( .A1(n13480), .A2(n9432), .ZN(n11004) );
  AND2_X1 U11236 ( .A1(n11006), .A2(n11004), .ZN(n9438) );
  AOI22_X1 U11237 ( .A1(n9435), .A2(n10835), .B1(n9434), .B2(n9433), .ZN(n9436) );
  NAND2_X1 U11238 ( .A1(n9439), .A2(n9436), .ZN(n9437) );
  OAI21_X1 U11239 ( .B1(n9439), .B2(n9438), .A(n9437), .ZN(n9440) );
  INV_X1 U11240 ( .A(n9440), .ZN(n9441) );
  NAND2_X1 U11241 ( .A1(n9442), .A2(n16718), .ZN(n9444) );
  NAND2_X1 U11242 ( .A1(n16717), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n9443) );
  NAND2_X1 U11243 ( .A1(n9444), .A2(n8846), .ZN(P3_U3488) );
  NAND2_X1 U11244 ( .A1(n10835), .A2(n14147), .ZN(n9445) );
  NAND2_X1 U11245 ( .A1(n9445), .A2(n10787), .ZN(n9446) );
  NAND2_X2 U11246 ( .A1(n9447), .A2(n9446), .ZN(n9450) );
  XNOR2_X1 U11247 ( .A(n9448), .B(n13815), .ZN(n13822) );
  NOR2_X1 U11248 ( .A1(n13822), .A2(n13821), .ZN(n13817) );
  AOI21_X1 U11249 ( .B1(n13822), .B2(n13821), .A(n13817), .ZN(n9520) );
  XNOR2_X1 U11250 ( .A(n9516), .B(n12423), .ZN(n9465) );
  XNOR2_X1 U11251 ( .A(n9516), .B(n16651), .ZN(n9464) );
  XNOR2_X1 U11252 ( .A(n9516), .B(n16614), .ZN(n9463) );
  XNOR2_X1 U11253 ( .A(n9516), .B(n16595), .ZN(n9462) );
  XNOR2_X1 U11254 ( .A(n9450), .B(n11836), .ZN(n9458) );
  INV_X1 U11255 ( .A(n9458), .ZN(n9459) );
  INV_X1 U11256 ( .A(n9456), .ZN(n9457) );
  AOI211_X1 U11257 ( .C1(n11400), .C2(n16497), .A(n11530), .B(n13815), .ZN(
        n9455) );
  OAI21_X1 U11258 ( .B1(n11403), .B2(n11333), .A(n11530), .ZN(n9452) );
  OAI211_X1 U11259 ( .C1(n13815), .C2(n16450), .A(n11333), .B(n11403), .ZN(
        n9451) );
  OAI21_X1 U11260 ( .B1(n9452), .B2(n9450), .A(n9451), .ZN(n9454) );
  XNOR2_X1 U11261 ( .A(n9456), .B(n11828), .ZN(n11421) );
  XNOR2_X1 U11262 ( .A(n9458), .B(n10554), .ZN(n11505) );
  NAND2_X1 U11263 ( .A1(n11504), .A2(n11505), .ZN(n11503) );
  XNOR2_X1 U11264 ( .A(n9460), .B(n12250), .ZN(n11660) );
  XNOR2_X1 U11265 ( .A(n9450), .B(n16580), .ZN(n9461) );
  XNOR2_X1 U11266 ( .A(n9461), .B(n13384), .ZN(n11680) );
  XNOR2_X1 U11267 ( .A(n9462), .B(n13391), .ZN(n11840) );
  XNOR2_X1 U11268 ( .A(n9463), .B(n12300), .ZN(n11968) );
  XNOR2_X1 U11269 ( .A(n9464), .B(n12420), .ZN(n12299) );
  XNOR2_X1 U11270 ( .A(n9465), .B(n12577), .ZN(n12415) );
  XNOR2_X1 U11271 ( .A(n13533), .B(n9516), .ZN(n12575) );
  XNOR2_X1 U11272 ( .A(n9516), .B(n14831), .ZN(n13874) );
  NAND2_X1 U11273 ( .A1(n13425), .A2(n9466), .ZN(n13414) );
  XOR2_X1 U11274 ( .A(n13414), .B(n9516), .Z(n13932) );
  NOR2_X1 U11275 ( .A1(n16712), .A2(n8160), .ZN(n9467) );
  INV_X1 U11276 ( .A(n9466), .ZN(n13421) );
  MUX2_X1 U11277 ( .A(n9467), .B(n13421), .S(n9516), .Z(n9468) );
  XNOR2_X1 U11278 ( .A(n14895), .B(n9516), .ZN(n9470) );
  XNOR2_X1 U11279 ( .A(n9470), .B(n12570), .ZN(n13835) );
  XNOR2_X1 U11280 ( .A(n14445), .B(n9516), .ZN(n9472) );
  XNOR2_X1 U11281 ( .A(n9472), .B(n9469), .ZN(n13976) );
  INV_X1 U11282 ( .A(n9470), .ZN(n9471) );
  NAND2_X1 U11283 ( .A1(n9471), .A2(n12570), .ZN(n13973) );
  NAND2_X1 U11284 ( .A1(n9472), .A2(n14363), .ZN(n13895) );
  XNOR2_X1 U11285 ( .A(n14886), .B(n13815), .ZN(n13906) );
  NAND2_X1 U11286 ( .A1(n13906), .A2(n13905), .ZN(n9484) );
  INV_X1 U11287 ( .A(n9484), .ZN(n9476) );
  XNOR2_X1 U11288 ( .A(n14441), .B(n9516), .ZN(n9483) );
  INV_X1 U11289 ( .A(n9483), .ZN(n9473) );
  NAND2_X1 U11290 ( .A1(n9473), .A2(n14348), .ZN(n13903) );
  OR2_X1 U11291 ( .A1(n13906), .A2(n13905), .ZN(n9474) );
  AND2_X1 U11292 ( .A1(n13903), .A2(n9474), .ZN(n9475) );
  OR2_X1 U11293 ( .A1(n9476), .A2(n9475), .ZN(n9482) );
  AND2_X1 U11294 ( .A1(n13895), .A2(n9482), .ZN(n13850) );
  XNOR2_X1 U11295 ( .A(n14881), .B(n9516), .ZN(n9479) );
  XNOR2_X1 U11296 ( .A(n9479), .B(n14264), .ZN(n13857) );
  INV_X1 U11297 ( .A(n13857), .ZN(n9478) );
  XNOR2_X1 U11298 ( .A(n14304), .B(n9516), .ZN(n9487) );
  INV_X1 U11299 ( .A(n9487), .ZN(n9477) );
  INV_X1 U11300 ( .A(n14313), .ZN(n13859) );
  NAND2_X1 U11301 ( .A1(n9477), .A2(n13859), .ZN(n13852) );
  OR2_X1 U11302 ( .A1(n9478), .A2(n13852), .ZN(n9481) );
  AND2_X1 U11303 ( .A1(n13850), .A2(n9481), .ZN(n13853) );
  INV_X1 U11304 ( .A(n14264), .ZN(n14298) );
  NAND2_X1 U11305 ( .A1(n9479), .A2(n14298), .ZN(n9480) );
  AND2_X1 U11306 ( .A1(n13853), .A2(n9480), .ZN(n9492) );
  INV_X1 U11307 ( .A(n9480), .ZN(n9491) );
  INV_X1 U11308 ( .A(n9481), .ZN(n9490) );
  INV_X1 U11309 ( .A(n9482), .ZN(n9486) );
  XNOR2_X1 U11310 ( .A(n9483), .B(n14348), .ZN(n13901) );
  AND2_X1 U11311 ( .A1(n13901), .A2(n9484), .ZN(n9485) );
  OR2_X1 U11312 ( .A1(n9486), .A2(n9485), .ZN(n13952) );
  XNOR2_X1 U11313 ( .A(n9487), .B(n14313), .ZN(n13955) );
  INV_X1 U11314 ( .A(n13955), .ZN(n9488) );
  AND2_X1 U11315 ( .A1(n13952), .A2(n9488), .ZN(n13851) );
  AND2_X1 U11316 ( .A1(n13851), .A2(n13857), .ZN(n9489) );
  OR2_X1 U11317 ( .A1(n9490), .A2(n9489), .ZN(n13854) );
  XNOR2_X1 U11318 ( .A(n14272), .B(n9516), .ZN(n9493) );
  XOR2_X1 U11319 ( .A(n14278), .B(n9493), .Z(n13924) );
  INV_X1 U11320 ( .A(n9493), .ZN(n9494) );
  NAND2_X1 U11321 ( .A1(n9494), .A2(n8153), .ZN(n9495) );
  INV_X1 U11322 ( .A(n13456), .ZN(n9496) );
  MUX2_X1 U11323 ( .A(n9497), .B(n9496), .S(n9516), .Z(n13866) );
  MUX2_X1 U11324 ( .A(n9498), .B(n13455), .S(n9516), .Z(n13864) );
  XNOR2_X1 U11325 ( .A(n13942), .B(n9516), .ZN(n9499) );
  XNOR2_X1 U11326 ( .A(n13847), .B(n9516), .ZN(n9505) );
  INV_X1 U11327 ( .A(n9505), .ZN(n9504) );
  OR2_X1 U11328 ( .A1(n14246), .A2(n9504), .ZN(n9502) );
  NAND2_X1 U11329 ( .A1(n13842), .A2(n13914), .ZN(n9509) );
  XNOR2_X1 U11330 ( .A(n13470), .B(n9516), .ZN(n9506) );
  NAND2_X1 U11331 ( .A1(n9506), .A2(n14220), .ZN(n13885) );
  INV_X1 U11332 ( .A(n9506), .ZN(n9507) );
  NAND2_X1 U11333 ( .A1(n9507), .A2(n14195), .ZN(n9508) );
  AND2_X1 U11334 ( .A1(n13885), .A2(n9508), .ZN(n13915) );
  NAND2_X1 U11335 ( .A1(n9509), .A2(n13915), .ZN(n13884) );
  NAND2_X1 U11336 ( .A1(n13884), .A2(n13885), .ZN(n9514) );
  XNOR2_X1 U11337 ( .A(n9510), .B(n9516), .ZN(n9511) );
  NAND2_X1 U11338 ( .A1(n9511), .A2(n14209), .ZN(n9515) );
  INV_X1 U11339 ( .A(n9511), .ZN(n9512) );
  NAND2_X1 U11340 ( .A1(n9512), .A2(n8350), .ZN(n9513) );
  NAND2_X1 U11341 ( .A1(n13888), .A2(n9515), .ZN(n13964) );
  XNOR2_X1 U11342 ( .A(n14854), .B(n9516), .ZN(n9517) );
  INV_X1 U11343 ( .A(n14198), .ZN(n14176) );
  NOR2_X1 U11344 ( .A1(n9517), .A2(n14176), .ZN(n9518) );
  AOI21_X1 U11345 ( .B1(n9517), .B2(n14176), .A(n9518), .ZN(n13965) );
  INV_X1 U11346 ( .A(n9518), .ZN(n9519) );
  NAND2_X1 U11347 ( .A1(n9528), .A2(n16711), .ZN(n9521) );
  OAI22_X1 U11348 ( .A1(n9529), .A2(n9521), .B1(n9533), .B2(n9525), .ZN(n9522)
         );
  NAND2_X1 U11349 ( .A1(n9529), .A2(n13550), .ZN(n9524) );
  NAND3_X1 U11350 ( .A1(n9589), .A2(n9642), .A3(n11004), .ZN(n9527) );
  INV_X1 U11351 ( .A(n9533), .ZN(n9531) );
  NOR2_X1 U11352 ( .A1(n9531), .A2(n9525), .ZN(n9526) );
  AOI211_X1 U11353 ( .C1(n9529), .C2(n9528), .A(n9527), .B(n9526), .ZN(n9532)
         );
  INV_X1 U11354 ( .A(n10789), .ZN(n9530) );
  NAND2_X1 U11355 ( .A1(n11012), .A2(n9530), .ZN(n13556) );
  OAI22_X2 U11356 ( .A1(n9532), .A2(P3_U3151), .B1(n9531), .B2(n13556), .ZN(
        n13970) );
  NOR2_X1 U11357 ( .A1(n9533), .A2(n13556), .ZN(n9536) );
  OAI22_X1 U11358 ( .A1(n14198), .A2(n13947), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n14644), .ZN(n9538) );
  NAND2_X2 U11359 ( .A1(n9536), .A2(n9535), .ZN(n13978) );
  NOR2_X1 U11360 ( .A1(n11040), .A2(n13978), .ZN(n9537) );
  AOI211_X1 U11361 ( .C1(n13970), .C2(n14178), .A(n9538), .B(n9537), .ZN(n9539) );
  NAND2_X1 U11362 ( .A1(n9542), .A2(n9541), .ZN(P3_U3154) );
  NAND4_X1 U11363 ( .A1(n10635), .A2(n9545), .A3(n14617), .A4(n9544), .ZN(
        n9551) );
  NOR2_X1 U11364 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n9549) );
  NOR2_X1 U11365 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), 
        .ZN(n9548) );
  NOR2_X1 U11366 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), 
        .ZN(n9547) );
  NOR2_X1 U11367 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n9546) );
  NAND4_X1 U11368 ( .A1(n9549), .A2(n9548), .A3(n9547), .A4(n9546), .ZN(n9550)
         );
  NAND2_X1 U11369 ( .A1(n9566), .A2(n9556), .ZN(n9569) );
  NOR2_X1 U11370 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), 
        .ZN(n9557) );
  NAND4_X1 U11371 ( .A1(n9557), .A2(n9552), .A3(n9556), .A4(n9555), .ZN(n9993)
         );
  NAND2_X1 U11372 ( .A1(n9563), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9564) );
  INV_X1 U11373 ( .A(n9566), .ZN(n9567) );
  NAND2_X1 U11374 ( .A1(n9567), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9568) );
  MUX2_X1 U11375 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9568), .S(
        P1_IR_REG_23__SCAN_IN), .Z(n9570) );
  INV_X1 U11376 ( .A(n9969), .ZN(n9571) );
  NOR2_X1 U11377 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), 
        .ZN(n9574) );
  NAND2_X1 U11378 ( .A1(n9586), .A2(n9696), .ZN(n9582) );
  NAND2_X1 U11379 ( .A1(n9585), .A2(n9697), .ZN(n9583) );
  XNOR2_X1 U11380 ( .A(n9586), .B(P2_IR_REG_24__SCAN_IN), .ZN(n9807) );
  NAND2_X1 U11381 ( .A1(n7460), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9587) );
  INV_X1 U11382 ( .A(n9818), .ZN(n9588) );
  XNOR2_X1 U11383 ( .A(n9647), .B(n9590), .ZN(n9687) );
  XNOR2_X1 U11384 ( .A(n9647), .B(n9591), .ZN(n9665) );
  MUX2_X1 U11385 ( .A(n9687), .B(n9665), .S(n14139), .Z(n9640) );
  INV_X1 U11386 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n11411) );
  MUX2_X1 U11387 ( .A(n11411), .B(n9592), .S(n14139), .Z(n9594) );
  INV_X1 U11388 ( .A(n10898), .ZN(n9593) );
  NAND2_X1 U11389 ( .A1(n9594), .A2(n9593), .ZN(n11224) );
  INV_X1 U11390 ( .A(n9594), .ZN(n9595) );
  NAND2_X1 U11391 ( .A1(n9595), .A2(n10898), .ZN(n9596) );
  AND2_X1 U11392 ( .A1(n11224), .A2(n9596), .ZN(n10893) );
  MUX2_X1 U11393 ( .A(n11017), .B(n9597), .S(n14139), .Z(n11302) );
  AND2_X1 U11394 ( .A1(n11302), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n11313) );
  NAND2_X1 U11395 ( .A1(n10893), .A2(n11313), .ZN(n11226) );
  NAND2_X1 U11396 ( .A1(n11226), .A2(n11224), .ZN(n9602) );
  MUX2_X1 U11397 ( .A(n9670), .B(n9598), .S(n14139), .Z(n9599) );
  NAND2_X1 U11398 ( .A1(n9599), .A2(n9671), .ZN(n10860) );
  INV_X1 U11399 ( .A(n9599), .ZN(n9600) );
  INV_X1 U11400 ( .A(n9671), .ZN(n11234) );
  NAND2_X1 U11401 ( .A1(n9600), .A2(n11234), .ZN(n9601) );
  AND2_X1 U11402 ( .A1(n10860), .A2(n9601), .ZN(n11223) );
  NAND2_X1 U11403 ( .A1(n9602), .A2(n11223), .ZN(n11228) );
  NAND2_X1 U11404 ( .A1(n11228), .A2(n10860), .ZN(n9607) );
  MUX2_X1 U11405 ( .A(n11820), .B(n9603), .S(n14139), .Z(n9604) );
  NAND2_X1 U11406 ( .A1(n9604), .A2(n9652), .ZN(n11206) );
  INV_X1 U11407 ( .A(n9604), .ZN(n9605) );
  INV_X1 U11408 ( .A(n9652), .ZN(n10868) );
  NAND2_X1 U11409 ( .A1(n9605), .A2(n10868), .ZN(n9606) );
  AND2_X1 U11410 ( .A1(n11206), .A2(n9606), .ZN(n10861) );
  NAND2_X1 U11411 ( .A1(n9607), .A2(n10861), .ZN(n11207) );
  NAND2_X1 U11412 ( .A1(n11207), .A2(n11206), .ZN(n9611) );
  INV_X1 U11413 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n9653) );
  MUX2_X1 U11414 ( .A(n11833), .B(n9653), .S(n14112), .Z(n9608) );
  NAND2_X1 U11415 ( .A1(n9608), .A2(n9847), .ZN(n9612) );
  INV_X1 U11416 ( .A(n9608), .ZN(n9609) );
  NAND2_X1 U11417 ( .A1(n9609), .A2(n7686), .ZN(n9610) );
  AND2_X1 U11418 ( .A1(n9612), .A2(n9610), .ZN(n11204) );
  NAND2_X1 U11419 ( .A1(n9611), .A2(n11204), .ZN(n11209) );
  NAND2_X1 U11420 ( .A1(n11209), .A2(n9612), .ZN(n10918) );
  MUX2_X1 U11421 ( .A(P3_REG2_REG_5__SCAN_IN), .B(P3_REG1_REG_5__SCAN_IN), .S(
        n14139), .Z(n9613) );
  XNOR2_X1 U11422 ( .A(n9613), .B(n10925), .ZN(n10917) );
  NAND2_X1 U11423 ( .A1(n10918), .A2(n10917), .ZN(n10916) );
  INV_X1 U11424 ( .A(n9613), .ZN(n9614) );
  NAND2_X1 U11425 ( .A1(n9614), .A2(n10925), .ZN(n9615) );
  NAND2_X1 U11426 ( .A1(n10916), .A2(n9615), .ZN(n10903) );
  INV_X1 U11427 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n9617) );
  MUX2_X1 U11428 ( .A(n9617), .B(n9616), .S(n14139), .Z(n9618) );
  AND2_X1 U11429 ( .A1(n9618), .A2(n7816), .ZN(n10899) );
  INV_X1 U11430 ( .A(n9618), .ZN(n9619) );
  NAND2_X1 U11431 ( .A1(n9619), .A2(n9855), .ZN(n10900) );
  MUX2_X1 U11432 ( .A(n9621), .B(n9620), .S(n14139), .Z(n9622) );
  XNOR2_X1 U11433 ( .A(n9622), .B(n11524), .ZN(n11514) );
  NAND2_X1 U11434 ( .A1(n9622), .A2(n11524), .ZN(n9623) );
  MUX2_X1 U11435 ( .A(P3_REG2_REG_8__SCAN_IN), .B(P3_REG1_REG_8__SCAN_IN), .S(
        n14139), .Z(n9624) );
  INV_X1 U11436 ( .A(n9881), .ZN(n11618) );
  XNOR2_X1 U11437 ( .A(n9624), .B(n11618), .ZN(n11607) );
  NAND2_X1 U11438 ( .A1(n11608), .A2(n11607), .ZN(n9627) );
  INV_X1 U11439 ( .A(n9624), .ZN(n9625) );
  NAND2_X1 U11440 ( .A1(n9625), .A2(n11618), .ZN(n9626) );
  NAND2_X1 U11441 ( .A1(n9627), .A2(n9626), .ZN(n16420) );
  MUX2_X1 U11442 ( .A(n12046), .B(n9628), .S(n14112), .Z(n9629) );
  XNOR2_X1 U11443 ( .A(n9629), .B(n9630), .ZN(n16419) );
  OR2_X1 U11444 ( .A1(n16420), .A2(n16419), .ZN(n16433) );
  INV_X1 U11445 ( .A(n9629), .ZN(n9631) );
  NAND2_X1 U11446 ( .A1(n9631), .A2(n16428), .ZN(n9632) );
  AND2_X1 U11447 ( .A1(n16433), .A2(n9632), .ZN(n11954) );
  MUX2_X1 U11448 ( .A(P3_REG2_REG_10__SCAN_IN), .B(P3_REG1_REG_10__SCAN_IN), 
        .S(n14139), .Z(n9633) );
  XNOR2_X1 U11449 ( .A(n9633), .B(n11963), .ZN(n11953) );
  NAND2_X1 U11450 ( .A1(n11954), .A2(n11953), .ZN(n11952) );
  INV_X1 U11451 ( .A(n9633), .ZN(n9634) );
  NAND2_X1 U11452 ( .A1(n9634), .A2(n11963), .ZN(n9635) );
  MUX2_X1 U11453 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n14139), .Z(n9636) );
  XNOR2_X1 U11454 ( .A(n9636), .B(n12166), .ZN(n12157) );
  INV_X1 U11455 ( .A(n9636), .ZN(n9637) );
  NAND2_X1 U11456 ( .A1(P3_U3897), .A2(n14921), .ZN(n16418) );
  INV_X1 U11457 ( .A(n13988), .ZN(n9638) );
  AOI211_X1 U11458 ( .C1(n9640), .C2(n9639), .A(n16418), .B(n9638), .ZN(n9695)
         );
  INV_X1 U11459 ( .A(n11012), .ZN(n9641) );
  OR2_X1 U11460 ( .A1(n9642), .A2(P3_U3151), .ZN(n13560) );
  NAND2_X1 U11461 ( .A1(n9641), .A2(n13560), .ZN(n9689) );
  NAND2_X1 U11462 ( .A1(n13480), .A2(n9642), .ZN(n9643) );
  NAND2_X1 U11463 ( .A1(n9644), .A2(n9643), .ZN(n9688) );
  INV_X1 U11464 ( .A(n9688), .ZN(n9645) );
  NAND2_X1 U11465 ( .A1(n9689), .A2(n9645), .ZN(n11212) );
  INV_X1 U11466 ( .A(n11212), .ZN(n9646) );
  MUX2_X1 U11467 ( .A(P3_U3897), .B(n9646), .S(n14921), .Z(n14146) );
  NOR2_X1 U11468 ( .A1(n16427), .A2(n13997), .ZN(n9694) );
  INV_X1 U11469 ( .A(n10925), .ZN(n9675) );
  NAND2_X1 U11470 ( .A1(n9668), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n9650) );
  INV_X1 U11471 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n11304) );
  NAND2_X1 U11472 ( .A1(P3_REG1_REG_0__SCAN_IN), .A2(n11304), .ZN(n9648) );
  OR2_X1 U11473 ( .A1(n9648), .A2(n9668), .ZN(n9649) );
  NAND2_X1 U11474 ( .A1(n10892), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n9651) );
  NAND2_X1 U11475 ( .A1(n9651), .A2(n9650), .ZN(n11221) );
  NOR2_X1 U11476 ( .A1(n9671), .A2(n9598), .ZN(n11222) );
  XNOR2_X1 U11477 ( .A(n9847), .B(n9653), .ZN(n11197) );
  AOI21_X1 U11478 ( .B1(P3_REG1_REG_4__SCAN_IN), .B2(n7686), .A(n11201), .ZN(
        n9654) );
  INV_X1 U11479 ( .A(n9654), .ZN(n9655) );
  XNOR2_X1 U11480 ( .A(n9654), .B(n10925), .ZN(n10920) );
  NAND2_X1 U11481 ( .A1(P3_REG1_REG_6__SCAN_IN), .A2(n9855), .ZN(n9656) );
  OAI21_X1 U11482 ( .B1(P3_REG1_REG_6__SCAN_IN), .B2(n9855), .A(n9656), .ZN(
        n10905) );
  NAND2_X1 U11483 ( .A1(P3_REG1_REG_8__SCAN_IN), .A2(n9881), .ZN(n9659) );
  OAI21_X1 U11484 ( .B1(P3_REG1_REG_8__SCAN_IN), .B2(n9881), .A(n9659), .ZN(
        n11613) );
  NAND2_X1 U11485 ( .A1(P3_REG1_REG_10__SCAN_IN), .A2(n9935), .ZN(n9660) );
  OAI21_X1 U11486 ( .B1(P3_REG1_REG_10__SCAN_IN), .B2(n9935), .A(n9660), .ZN(
        n11950) );
  AND2_X1 U11487 ( .A1(n9935), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n9661) );
  NAND2_X1 U11488 ( .A1(n9663), .A2(n9684), .ZN(n9662) );
  INV_X1 U11489 ( .A(n9662), .ZN(n9664) );
  INV_X1 U11490 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n16690) );
  AOI21_X1 U11491 ( .B1(n9665), .B2(n7456), .A(n13992), .ZN(n9666) );
  NOR2_X1 U11492 ( .A1(n16429), .A2(n9666), .ZN(n9693) );
  NAND2_X1 U11493 ( .A1(n9935), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n9683) );
  NAND2_X1 U11494 ( .A1(P3_REG2_REG_0__SCAN_IN), .A2(n11304), .ZN(n11310) );
  NAND2_X1 U11495 ( .A1(n9668), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n9669) );
  NAND2_X1 U11496 ( .A1(n9671), .A2(n9670), .ZN(n9672) );
  NAND2_X1 U11497 ( .A1(n11218), .A2(n9672), .ZN(n9673) );
  NAND2_X1 U11498 ( .A1(n11234), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n11215) );
  NAND2_X1 U11499 ( .A1(n11216), .A2(n10868), .ZN(n9674) );
  OAI21_X1 U11500 ( .B1(n11216), .B2(n10868), .A(n9674), .ZN(n10855) );
  INV_X1 U11501 ( .A(n9674), .ZN(n11192) );
  XNOR2_X1 U11502 ( .A(n9847), .B(P3_REG2_REG_4__SCAN_IN), .ZN(n11191) );
  NAND2_X1 U11503 ( .A1(P3_REG2_REG_6__SCAN_IN), .A2(n9855), .ZN(n9676) );
  OAI21_X1 U11504 ( .B1(P3_REG2_REG_6__SCAN_IN), .B2(n9855), .A(n9676), .ZN(
        n10908) );
  NAND2_X1 U11505 ( .A1(P3_REG2_REG_8__SCAN_IN), .A2(n9881), .ZN(n9679) );
  OAI21_X1 U11506 ( .B1(P3_REG2_REG_8__SCAN_IN), .B2(n9881), .A(n9679), .ZN(
        n11606) );
  AND2_X1 U11507 ( .A1(n9881), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n9680) );
  OAI21_X1 U11508 ( .B1(P3_REG2_REG_10__SCAN_IN), .B2(n9935), .A(n9683), .ZN(
        n11959) );
  NAND2_X1 U11509 ( .A1(n9683), .A2(n11956), .ZN(n9685) );
  INV_X1 U11510 ( .A(n12166), .ZN(n9684) );
  AOI21_X1 U11511 ( .B1(n9687), .B2(n9686), .A(n13996), .ZN(n9691) );
  NAND2_X1 U11512 ( .A1(P3_REG3_REG_12__SCAN_IN), .A2(P3_U3151), .ZN(n13878)
         );
  NAND2_X1 U11513 ( .A1(n16150), .A2(P3_ADDR_REG_12__SCAN_IN), .ZN(n9690) );
  OAI211_X1 U11514 ( .C1(n16423), .C2(n9691), .A(n13878), .B(n9690), .ZN(n9692) );
  INV_X4 U11515 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  INV_X4 U11516 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  NOR2_X1 U11517 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), 
        .ZN(n9700) );
  NAND2_X1 U11518 ( .A1(n9786), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n9709) );
  AND2_X2 U11519 ( .A1(n9705), .A2(n12646), .ZN(n9789) );
  NAND2_X1 U11520 ( .A1(n9789), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n9708) );
  AND2_X2 U11521 ( .A1(n15526), .A2(n12646), .ZN(n9788) );
  NAND2_X1 U11522 ( .A1(n9788), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n9707) );
  NAND2_X1 U11523 ( .A1(n9790), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n9706) );
  INV_X1 U11524 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n10130) );
  NAND2_X1 U11525 ( .A1(n7416), .A2(SI_0_), .ZN(n9711) );
  NAND2_X1 U11526 ( .A1(n9711), .A2(n9710), .ZN(n9712) );
  AND2_X1 U11527 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n9751) );
  NAND2_X1 U11528 ( .A1(n13247), .A2(n9751), .ZN(n9737) );
  NAND2_X1 U11529 ( .A1(n9712), .A2(n9737), .ZN(n15546) );
  INV_X1 U11530 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n9715) );
  INV_X1 U11531 ( .A(n13012), .ZN(n10984) );
  NAND2_X1 U11532 ( .A1(n9718), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9719) );
  MUX2_X1 U11533 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9719), .S(
        P2_IR_REG_22__SCAN_IN), .Z(n9720) );
  NAND2_X1 U11534 ( .A1(n9723), .A2(n9722), .ZN(n9729) );
  INV_X1 U11535 ( .A(n9724), .ZN(n9725) );
  NAND2_X1 U11536 ( .A1(n13345), .A2(n9730), .ZN(n13340) );
  XNOR2_X1 U11537 ( .A(n13340), .B(n8082), .ZN(n9732) );
  XNOR2_X1 U11538 ( .A(n9731), .B(P2_IR_REG_19__SCAN_IN), .ZN(n9824) );
  NAND2_X1 U11539 ( .A1(n9732), .A2(n13338), .ZN(n10226) );
  NAND2_X1 U11540 ( .A1(n10226), .A2(n13340), .ZN(n11068) );
  NAND2_X1 U11541 ( .A1(n14929), .A2(n13012), .ZN(n9733) );
  NAND2_X1 U11542 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n9734) );
  MUX2_X1 U11543 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9734), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n9736) );
  INV_X1 U11544 ( .A(n9758), .ZN(n9735) );
  NAND2_X1 U11545 ( .A1(n9736), .A2(n9735), .ZN(n10128) );
  AND2_X1 U11546 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(SI_0_), .ZN(n9748) );
  NAND2_X1 U11547 ( .A1(n9844), .A2(n9748), .ZN(n10269) );
  NAND2_X1 U11548 ( .A1(n10269), .A2(n9737), .ZN(n9738) );
  XNOR2_X1 U11549 ( .A(n11068), .B(n13024), .ZN(n11127) );
  NAND2_X1 U11550 ( .A1(n9789), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n9743) );
  NAND2_X1 U11551 ( .A1(n9790), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n9742) );
  XNOR2_X1 U11552 ( .A(n11127), .B(n9745), .ZN(n10565) );
  INV_X1 U11553 ( .A(n11127), .ZN(n9746) );
  NAND2_X1 U11554 ( .A1(n9746), .A2(n9745), .ZN(n9747) );
  NAND2_X1 U11555 ( .A1(n11128), .A2(n9747), .ZN(n9765) );
  OAI21_X1 U11556 ( .B1(P2_DATAO_REG_1__SCAN_IN), .B2(SI_1_), .A(n9748), .ZN(
        n9750) );
  NAND2_X1 U11557 ( .A1(P2_DATAO_REG_1__SCAN_IN), .A2(SI_1_), .ZN(n9749) );
  AND2_X1 U11558 ( .A1(n9750), .A2(n9749), .ZN(n9771) );
  OAI21_X1 U11559 ( .B1(SI_1_), .B2(P1_DATAO_REG_1__SCAN_IN), .A(n9751), .ZN(
        n9753) );
  NAND2_X1 U11560 ( .A1(SI_1_), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n9752) );
  NAND2_X1 U11561 ( .A1(n9753), .A2(n9752), .ZN(n9776) );
  NAND2_X1 U11562 ( .A1(n9874), .A2(n9776), .ZN(n9754) );
  OAI21_X1 U11563 ( .B1(n9771), .B2(n9874), .A(n9754), .ZN(n9755) );
  XNOR2_X1 U11564 ( .A(n9755), .B(SI_2_), .ZN(n9757) );
  MUX2_X1 U11565 ( .A(n10407), .B(n9882), .S(n9874), .Z(n9756) );
  OR2_X1 U11566 ( .A1(n9758), .A2(n9715), .ZN(n9760) );
  XNOR2_X1 U11567 ( .A(n9760), .B(n9759), .ZN(n15045) );
  XNOR2_X1 U11568 ( .A(n14936), .B(n13021), .ZN(n9766) );
  NAND2_X1 U11569 ( .A1(n9786), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n9764) );
  NAND2_X1 U11570 ( .A1(n9788), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n9763) );
  NAND2_X1 U11571 ( .A1(n9789), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n9762) );
  NAND2_X1 U11572 ( .A1(n9790), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n9761) );
  NAND2_X1 U11573 ( .A1(n15042), .A2(n14937), .ZN(n9767) );
  XNOR2_X1 U11574 ( .A(n9766), .B(n9767), .ZN(n11129) );
  NAND2_X1 U11575 ( .A1(n9765), .A2(n11129), .ZN(n11135) );
  INV_X1 U11576 ( .A(n9766), .ZN(n9768) );
  NAND2_X1 U11577 ( .A1(n9768), .A2(n9767), .ZN(n9769) );
  INV_X1 U11578 ( .A(n9771), .ZN(n9772) );
  OAI21_X1 U11579 ( .B1(P2_DATAO_REG_2__SCAN_IN), .B2(SI_2_), .A(n9772), .ZN(
        n9774) );
  NAND2_X1 U11580 ( .A1(P2_DATAO_REG_2__SCAN_IN), .A2(SI_2_), .ZN(n9773) );
  NAND2_X1 U11581 ( .A1(n9774), .A2(n9773), .ZN(n9775) );
  NAND2_X1 U11582 ( .A1(n8976), .A2(n9775), .ZN(n9781) );
  OAI21_X1 U11583 ( .B1(SI_2_), .B2(P1_DATAO_REG_2__SCAN_IN), .A(n9776), .ZN(
        n9778) );
  NAND2_X1 U11584 ( .A1(SI_2_), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n9777) );
  NAND2_X1 U11585 ( .A1(n9778), .A2(n9777), .ZN(n9779) );
  NAND2_X1 U11586 ( .A1(n9779), .A2(n13247), .ZN(n9780) );
  NAND2_X1 U11587 ( .A1(n9781), .A2(n9780), .ZN(n9868) );
  XNOR2_X1 U11588 ( .A(n9869), .B(n9868), .ZN(n10683) );
  OR2_X1 U11589 ( .A1(n9884), .A2(n9715), .ZN(n9782) );
  XNOR2_X1 U11590 ( .A(n9782), .B(n9883), .ZN(n10103) );
  OR2_X1 U11591 ( .A1(n11062), .A2(n10103), .ZN(n9785) );
  OR2_X1 U11592 ( .A1(n9783), .A2(n9895), .ZN(n9784) );
  XNOR2_X1 U11593 ( .A(n10581), .B(n14936), .ZN(n11170) );
  INV_X1 U11594 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n9787) );
  NAND2_X1 U11595 ( .A1(n9786), .A2(n9787), .ZN(n9794) );
  NAND2_X1 U11596 ( .A1(n10847), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n9793) );
  NAND2_X1 U11597 ( .A1(n9789), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n9792) );
  NAND2_X1 U11598 ( .A1(n9790), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n9791) );
  NAND4_X1 U11599 ( .A1(n9794), .A2(n9793), .A3(n9792), .A4(n9791), .ZN(n15041) );
  NAND2_X1 U11600 ( .A1(n15041), .A2(n14937), .ZN(n9795) );
  NAND2_X1 U11601 ( .A1(n11170), .A2(n9795), .ZN(n9798) );
  INV_X1 U11602 ( .A(n11170), .ZN(n9797) );
  INV_X1 U11603 ( .A(n9795), .ZN(n9796) );
  NAND2_X1 U11604 ( .A1(n9797), .A2(n9796), .ZN(n10645) );
  NAND2_X1 U11605 ( .A1(n9798), .A2(n10645), .ZN(n9822) );
  INV_X1 U11606 ( .A(n10647), .ZN(n11172) );
  NOR4_X1 U11607 ( .A1(P2_D_REG_19__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n9802) );
  NOR4_X1 U11608 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n9801) );
  NOR4_X1 U11609 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_6__SCAN_IN), .ZN(n9800) );
  NOR4_X1 U11610 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n9799) );
  NAND4_X1 U11611 ( .A1(n9802), .A2(n9801), .A3(n9800), .A4(n9799), .ZN(n9813)
         );
  NOR2_X1 U11612 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .ZN(
        n9806) );
  NOR4_X1 U11613 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n9805) );
  NOR4_X1 U11614 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n9804) );
  NOR4_X1 U11615 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n9803) );
  NAND4_X1 U11616 ( .A1(n9806), .A2(n9805), .A3(n9804), .A4(n9803), .ZN(n9812)
         );
  AOI22_X1 U11617 ( .A1(P2_B_REG_SCAN_IN), .A2(n15539), .B1(n9807), .B2(n15112), .ZN(n9808) );
  INV_X1 U11618 ( .A(n9808), .ZN(n9809) );
  AND2_X1 U11619 ( .A1(n15536), .A2(n9809), .ZN(n9810) );
  INV_X1 U11620 ( .A(n16147), .ZN(n9811) );
  OR2_X1 U11621 ( .A1(n16147), .A2(P2_D_REG_1__SCAN_IN), .ZN(n9815) );
  NAND2_X1 U11622 ( .A1(n15534), .A2(n15536), .ZN(n9814) );
  AND2_X1 U11623 ( .A1(n9815), .A2(n9814), .ZN(n11243) );
  NAND2_X1 U11624 ( .A1(n15534), .A2(n15539), .ZN(n9816) );
  AND3_X1 U11625 ( .A1(n11243), .A2(n11242), .A3(n16148), .ZN(n9819) );
  NAND2_X1 U11626 ( .A1(n10223), .A2(n9819), .ZN(n9831) );
  NAND2_X1 U11627 ( .A1(n10232), .A2(n13351), .ZN(n16678) );
  INV_X1 U11628 ( .A(n10077), .ZN(n9820) );
  NAND2_X1 U11629 ( .A1(n16678), .A2(n9820), .ZN(n9821) );
  AOI211_X1 U11630 ( .C1(n9823), .C2(n9822), .A(n11172), .B(n15021), .ZN(n9841) );
  INV_X1 U11631 ( .A(n11242), .ZN(n10239) );
  NAND2_X1 U11632 ( .A1(n11243), .A2(n10223), .ZN(n9825) );
  INV_X1 U11633 ( .A(n9829), .ZN(n10224) );
  OAI21_X1 U11634 ( .B1(n10239), .B2(n9825), .A(n10224), .ZN(n9827) );
  NAND2_X1 U11635 ( .A1(n10077), .A2(n13351), .ZN(n10222) );
  AND3_X1 U11636 ( .A1(n10076), .A2(n13350), .A3(n10222), .ZN(n9826) );
  NAND2_X1 U11637 ( .A1(n9827), .A2(n9826), .ZN(n10563) );
  NAND2_X1 U11638 ( .A1(n10563), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15003) );
  INV_X1 U11639 ( .A(n15003), .ZN(n15018) );
  MUX2_X1 U11640 ( .A(n15018), .B(P2_U3088), .S(P2_REG3_REG_3__SCAN_IN), .Z(
        n9840) );
  INV_X1 U11641 ( .A(n9831), .ZN(n9828) );
  AND2_X1 U11642 ( .A1(n10232), .A2(n13307), .ZN(n11258) );
  NAND2_X1 U11643 ( .A1(n9828), .A2(n11258), .ZN(n9830) );
  INV_X1 U11644 ( .A(n14991), .ZN(n15020) );
  INV_X1 U11645 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n9832) );
  XNOR2_X1 U11646 ( .A(n9832), .B(P2_REG3_REG_3__SCAN_IN), .ZN(n11282) );
  NAND2_X1 U11647 ( .A1(n9786), .A2(n11282), .ZN(n9836) );
  NAND2_X1 U11648 ( .A1(n10847), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n9835) );
  NAND2_X1 U11649 ( .A1(n9789), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n9834) );
  NAND2_X1 U11650 ( .A1(n9790), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n9833) );
  NAND4_X1 U11651 ( .A1(n9836), .A2(n9835), .A3(n9834), .A4(n9833), .ZN(n15040) );
  INV_X1 U11652 ( .A(n15040), .ZN(n10485) );
  INV_X1 U11653 ( .A(n15343), .ZN(n15287) );
  INV_X1 U11654 ( .A(n15042), .ZN(n10547) );
  INV_X1 U11655 ( .A(n10089), .ZN(n9837) );
  OAI22_X1 U11656 ( .A1(n10485), .A2(n15287), .B1(n10547), .B2(n15289), .ZN(
        n10541) );
  INV_X1 U11657 ( .A(n10541), .ZN(n9838) );
  OAI22_X1 U11658 ( .A1(n10581), .A2(n14994), .B1(n15020), .B2(n9838), .ZN(
        n9839) );
  OR3_X1 U11659 ( .A1(n9841), .A2(n9840), .A3(n9839), .ZN(P2_U3190) );
  NAND2_X1 U11660 ( .A1(n9842), .A2(P3_U3151), .ZN(n9843) );
  OAI21_X1 U11661 ( .B1(n11304), .B2(P3_U3151), .A(n9843), .ZN(P3_U3295) );
  AOI222_X1 U11662 ( .A1(n9845), .A2(n14901), .B1(SI_5_), .B2(n9852), .C1(
        n10925), .C2(P3_STATE_REG_SCAN_IN), .ZN(n9846) );
  INV_X1 U11663 ( .A(n9846), .ZN(P3_U3290) );
  AOI222_X1 U11664 ( .A1(n9848), .A2(n14901), .B1(n9847), .B2(
        P3_STATE_REG_SCAN_IN), .C1(SI_4_), .C2(n9852), .ZN(n9849) );
  INV_X1 U11665 ( .A(n9849), .ZN(P3_U3291) );
  AOI222_X1 U11666 ( .A1(n9850), .A2(n14901), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n11524), .C1(SI_7_), .C2(n9852), .ZN(n9851) );
  INV_X1 U11667 ( .A(n9851), .ZN(P3_U3288) );
  INV_X1 U11668 ( .A(n14901), .ZN(n14918) );
  OAI222_X1 U11669 ( .A1(P3_U3151), .A2(n9855), .B1(n14918), .B2(n9854), .C1(
        n9853), .C2(n14920), .ZN(P3_U3289) );
  INV_X1 U11670 ( .A(n9856), .ZN(n9858) );
  INV_X1 U11671 ( .A(SI_2_), .ZN(n9857) );
  OAI222_X1 U11672 ( .A1(n11234), .A2(P3_U3151), .B1(n14918), .B2(n9858), .C1(
        n9857), .C2(n14920), .ZN(P3_U3293) );
  INV_X1 U11673 ( .A(n9859), .ZN(n9860) );
  INV_X1 U11674 ( .A(SI_3_), .ZN(n9866) );
  OAI222_X1 U11675 ( .A1(n10868), .A2(P3_U3151), .B1(n14918), .B2(n9860), .C1(
        n9866), .C2(n14920), .ZN(P3_U3292) );
  OAI222_X1 U11676 ( .A1(P3_U3151), .A2(n10898), .B1(n14918), .B2(n9862), .C1(
        n9861), .C2(n14920), .ZN(P3_U3294) );
  INV_X2 U11677 ( .A(n11168), .ZN(n16139) );
  INV_X2 U11678 ( .A(n16135), .ZN(n11886) );
  NAND2_X1 U11679 ( .A1(n9863), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9865) );
  INV_X1 U11680 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n9864) );
  XNOR2_X1 U11681 ( .A(n9865), .B(n9864), .ZN(n10687) );
  OAI222_X1 U11682 ( .A1(n16139), .A2(n10684), .B1(n11886), .B2(n10683), .C1(
        P1_U3086), .C2(n10687), .ZN(P1_U3352) );
  INV_X1 U11683 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n10464) );
  INV_X1 U11684 ( .A(n9871), .ZN(n9872) );
  NAND2_X1 U11685 ( .A1(n9872), .A2(SI_4_), .ZN(n9873) );
  XNOR2_X1 U11686 ( .A(n9896), .B(n9897), .ZN(n10732) );
  INV_X1 U11687 ( .A(n10732), .ZN(n9886) );
  INV_X1 U11688 ( .A(n9875), .ZN(n9876) );
  NAND2_X1 U11689 ( .A1(n9876), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9877) );
  XNOR2_X1 U11690 ( .A(n9877), .B(P1_IR_REG_5__SCAN_IN), .ZN(n10731) );
  INV_X1 U11691 ( .A(n10731), .ZN(n10074) );
  OAI222_X1 U11692 ( .A1(n16139), .A2(n9878), .B1(n11886), .B2(n9886), .C1(
        P1_U3086), .C2(n10074), .ZN(P1_U3350) );
  OAI222_X1 U11693 ( .A1(P3_U3151), .A2(n9881), .B1(n14920), .B2(n9880), .C1(
        n14918), .C2(n9879), .ZN(P3_U3287) );
  INV_X2 U11694 ( .A(n15542), .ZN(n15540) );
  OAI222_X1 U11695 ( .A1(n15045), .A2(P2_U3088), .B1(n15540), .B2(n10408), 
        .C1(n9882), .C2(n15545), .ZN(P2_U3325) );
  INV_X1 U11696 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n9887) );
  NAND2_X1 U11697 ( .A1(n9884), .A2(n9883), .ZN(n9890) );
  NAND2_X1 U11698 ( .A1(n9910), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9885) );
  XNOR2_X1 U11699 ( .A(n9885), .B(P2_IR_REG_5__SCAN_IN), .ZN(n15083) );
  INV_X1 U11700 ( .A(n15083), .ZN(n15077) );
  OAI222_X1 U11701 ( .A1(n15545), .A2(n9887), .B1(n15540), .B2(n9886), .C1(
        P2_U3088), .C2(n15077), .ZN(P2_U3322) );
  XNOR2_X1 U11702 ( .A(n9889), .B(n9888), .ZN(n10703) );
  INV_X1 U11703 ( .A(n10703), .ZN(n9932) );
  NAND2_X1 U11704 ( .A1(n9890), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9891) );
  MUX2_X1 U11705 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9891), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n9892) );
  NAND2_X1 U11706 ( .A1(n9892), .A2(n9910), .ZN(n15069) );
  OAI222_X1 U11707 ( .A1(n15545), .A2(n10464), .B1(n15540), .B2(n9932), .C1(
        P2_U3088), .C2(n15069), .ZN(P2_U3323) );
  OAI222_X1 U11708 ( .A1(n10128), .A2(P2_U3088), .B1(n15540), .B2(n9893), .C1(
        n9894), .C2(n15545), .ZN(P2_U3326) );
  OAI222_X1 U11709 ( .A1(n15545), .A2(n9895), .B1(n15540), .B2(n10683), .C1(
        P2_U3088), .C2(n10103), .ZN(P2_U3324) );
  MUX2_X1 U11710 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n13247), .Z(n9918) );
  XNOR2_X1 U11711 ( .A(n9918), .B(SI_6_), .ZN(n9915) );
  XNOR2_X1 U11712 ( .A(n9917), .B(n9915), .ZN(n10811) );
  INV_X1 U11713 ( .A(n10811), .ZN(n9913) );
  INV_X1 U11714 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n9899) );
  AND2_X1 U11715 ( .A1(n9875), .A2(n9899), .ZN(n9921) );
  INV_X1 U11716 ( .A(n9921), .ZN(n9900) );
  NAND2_X1 U11717 ( .A1(n9900), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9901) );
  XNOR2_X1 U11718 ( .A(n9901), .B(P1_IR_REG_6__SCAN_IN), .ZN(n10812) );
  INV_X1 U11719 ( .A(n10812), .ZN(n10052) );
  OAI222_X1 U11720 ( .A1(n16139), .A2(n9902), .B1(n11886), .B2(n9913), .C1(
        P1_U3086), .C2(n10052), .ZN(P1_U3349) );
  NAND2_X1 U11721 ( .A1(n7469), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9903) );
  MUX2_X1 U11722 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9903), .S(
        P1_IR_REG_2__SCAN_IN), .Z(n9904) );
  NAND2_X1 U11723 ( .A1(n9904), .A2(n9863), .ZN(n10409) );
  OAI222_X1 U11724 ( .A1(n10409), .A2(P1_U3086), .B1(n11886), .B2(n10408), 
        .C1(n10407), .C2(n16139), .ZN(P1_U3353) );
  NAND2_X1 U11725 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n9905) );
  MUX2_X1 U11726 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9905), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n9906) );
  NAND2_X1 U11727 ( .A1(n9906), .A2(n7469), .ZN(n10364) );
  OAI222_X1 U11728 ( .A1(n10364), .A2(P1_U3086), .B1(n11886), .B2(n9893), .C1(
        n8094), .C2(n16139), .ZN(P1_U3354) );
  INV_X1 U11729 ( .A(SI_9_), .ZN(n9909) );
  INV_X1 U11730 ( .A(n9907), .ZN(n9908) );
  OAI222_X1 U11731 ( .A1(P3_U3151), .A2(n16428), .B1(n14920), .B2(n9909), .C1(
        n14918), .C2(n9908), .ZN(P3_U3286) );
  OR2_X1 U11732 ( .A1(n10148), .A2(n9715), .ZN(n9911) );
  XNOR2_X1 U11733 ( .A(n9911), .B(P2_IR_REG_6__SCAN_IN), .ZN(n15105) );
  INV_X1 U11734 ( .A(n15105), .ZN(n9912) );
  OAI222_X1 U11735 ( .A1(n15545), .A2(n9914), .B1(n15540), .B2(n9913), .C1(
        P2_U3088), .C2(n9912), .ZN(P2_U3321) );
  INV_X1 U11736 ( .A(n9915), .ZN(n9916) );
  NAND2_X1 U11737 ( .A1(n9918), .A2(SI_6_), .ZN(n9919) );
  XNOR2_X1 U11738 ( .A(n9939), .B(SI_7_), .ZN(n9936) );
  XNOR2_X1 U11739 ( .A(n9938), .B(n9936), .ZN(n11053) );
  INV_X1 U11740 ( .A(n11053), .ZN(n9927) );
  INV_X1 U11741 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n9920) );
  NAND2_X1 U11742 ( .A1(n9921), .A2(n9920), .ZN(n9941) );
  NAND2_X1 U11743 ( .A1(n9941), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9922) );
  XNOR2_X1 U11744 ( .A(n9922), .B(P1_IR_REG_7__SCAN_IN), .ZN(n11023) );
  INV_X1 U11745 ( .A(n11023), .ZN(n10202) );
  OAI222_X1 U11746 ( .A1(n16139), .A2(n9923), .B1(n11886), .B2(n9927), .C1(
        P1_U3086), .C2(n10202), .ZN(P1_U3348) );
  INV_X1 U11747 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n9924) );
  NAND2_X1 U11748 ( .A1(n10148), .A2(n9924), .ZN(n9944) );
  NAND2_X1 U11749 ( .A1(n9944), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9925) );
  XNOR2_X1 U11750 ( .A(n9925), .B(P2_IR_REG_7__SCAN_IN), .ZN(n16172) );
  INV_X1 U11751 ( .A(n16172), .ZN(n9926) );
  OAI222_X1 U11752 ( .A1(n15545), .A2(n9928), .B1(n15540), .B2(n9927), .C1(
        P2_U3088), .C2(n9926), .ZN(P2_U3320) );
  NAND2_X1 U11753 ( .A1(n9929), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9931) );
  INV_X1 U11754 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n9930) );
  XNOR2_X1 U11755 ( .A(n9931), .B(n9930), .ZN(n10708) );
  OAI222_X1 U11756 ( .A1(n16139), .A2(n10705), .B1(n11886), .B2(n9932), .C1(
        P1_U3086), .C2(n10708), .ZN(P1_U3351) );
  INV_X1 U11757 ( .A(SI_10_), .ZN(n14680) );
  INV_X1 U11758 ( .A(n9933), .ZN(n9934) );
  OAI222_X1 U11759 ( .A1(P3_U3151), .A2(n9935), .B1(n14920), .B2(n14680), .C1(
        n14918), .C2(n9934), .ZN(P3_U3285) );
  INV_X1 U11760 ( .A(n9936), .ZN(n9937) );
  NAND2_X1 U11761 ( .A1(n9939), .A2(SI_7_), .ZN(n9940) );
  MUX2_X1 U11762 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n13247), .Z(n9956) );
  XNOR2_X1 U11763 ( .A(n9955), .B(n9953), .ZN(n11539) );
  INV_X1 U11764 ( .A(n11539), .ZN(n9948) );
  NAND2_X1 U11765 ( .A1(n9957), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9942) );
  XNOR2_X1 U11766 ( .A(n9942), .B(P1_IR_REG_8__SCAN_IN), .ZN(n11540) );
  INV_X1 U11767 ( .A(n11540), .ZN(n10209) );
  OAI222_X1 U11768 ( .A1(n16139), .A2(n9943), .B1(n11886), .B2(n9948), .C1(
        P1_U3086), .C2(n10209), .ZN(P1_U3347) );
  INV_X1 U11769 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n11064) );
  NAND2_X1 U11770 ( .A1(n9946), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9945) );
  MUX2_X1 U11771 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9945), .S(
        P2_IR_REG_8__SCAN_IN), .Z(n9947) );
  NAND2_X1 U11772 ( .A1(n9947), .A2(n9979), .ZN(n11063) );
  OAI222_X1 U11773 ( .A1(n15545), .A2(n11064), .B1(n15540), .B2(n9948), .C1(
        P2_U3088), .C2(n11063), .ZN(P2_U3319) );
  INV_X1 U11774 ( .A(n9949), .ZN(n9950) );
  OAI222_X1 U11775 ( .A1(P3_U3151), .A2(n9684), .B1(n14920), .B2(n14679), .C1(
        n14918), .C2(n9950), .ZN(P3_U3284) );
  INV_X1 U11776 ( .A(n9951), .ZN(n9952) );
  OAI222_X1 U11777 ( .A1(P3_U3151), .A2(n13997), .B1(n14920), .B2(n14676), 
        .C1(n14918), .C2(n9952), .ZN(P3_U3283) );
  INV_X1 U11778 ( .A(n9953), .ZN(n9954) );
  MUX2_X1 U11779 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n7416), .Z(n9973) );
  XNOR2_X1 U11780 ( .A(n9972), .B(n9973), .ZN(n11545) );
  INV_X1 U11781 ( .A(n11545), .ZN(n9961) );
  INV_X1 U11782 ( .A(n10637), .ZN(n9958) );
  NAND2_X1 U11783 ( .A1(n9958), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9976) );
  XNOR2_X1 U11784 ( .A(n9976), .B(P1_IR_REG_9__SCAN_IN), .ZN(n11546) );
  INV_X1 U11785 ( .A(n11546), .ZN(n10605) );
  OAI222_X1 U11786 ( .A1(n16139), .A2(n9959), .B1(n11886), .B2(n9961), .C1(
        P1_U3086), .C2(n10605), .ZN(P1_U3346) );
  INV_X1 U11787 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n9962) );
  NAND2_X1 U11788 ( .A1(n9979), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9960) );
  XNOR2_X1 U11789 ( .A(n9960), .B(P2_IR_REG_9__SCAN_IN), .ZN(n11078) );
  INV_X1 U11790 ( .A(n11078), .ZN(n10187) );
  OAI222_X1 U11791 ( .A1(n15545), .A2(n9962), .B1(n15540), .B2(n9961), .C1(
        P2_U3088), .C2(n10187), .ZN(P2_U3318) );
  INV_X1 U11792 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n13501) );
  INV_X1 U11793 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n9965) );
  NAND2_X1 U11794 ( .A1(n9789), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n9964) );
  NAND2_X1 U11795 ( .A1(n10847), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n9963) );
  OAI211_X1 U11796 ( .C1(n13265), .C2(n9965), .A(n9964), .B(n9963), .ZN(n15114) );
  NAND2_X1 U11797 ( .A1(P2_U3947), .A2(n15114), .ZN(n9966) );
  OAI21_X1 U11798 ( .B1(P2_U3947), .B2(n13501), .A(n9966), .ZN(P2_U3562) );
  NAND2_X1 U11799 ( .A1(n10379), .A2(n15739), .ZN(n9967) );
  NAND2_X1 U11800 ( .A1(n10381), .A2(n10878), .ZN(n16144) );
  INV_X1 U11801 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n9971) );
  OR2_X1 U11802 ( .A1(n10380), .A2(n16128), .ZN(n10366) );
  INV_X1 U11803 ( .A(n10366), .ZN(n9970) );
  AOI22_X1 U11804 ( .A1(n16144), .A2(n9971), .B1(n9970), .B2(n10878), .ZN(
        P1_U3446) );
  NAND2_X1 U11805 ( .A1(n9974), .A2(SI_9_), .ZN(n9975) );
  MUX2_X1 U11806 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n9874), .Z(n10002) );
  XNOR2_X1 U11807 ( .A(n10002), .B(SI_10_), .ZN(n9999) );
  XNOR2_X1 U11808 ( .A(n10001), .B(n9999), .ZN(n11558) );
  INV_X1 U11809 ( .A(n11558), .ZN(n9983) );
  INV_X1 U11810 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n10633) );
  NAND2_X1 U11811 ( .A1(n9976), .A2(n10633), .ZN(n9977) );
  NAND2_X1 U11812 ( .A1(n9977), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10008) );
  XNOR2_X1 U11813 ( .A(n10008), .B(P1_IR_REG_10__SCAN_IN), .ZN(n11559) );
  INV_X1 U11814 ( .A(n11559), .ZN(n10613) );
  OAI222_X1 U11815 ( .A1(n16139), .A2(n9978), .B1(n11886), .B2(n9983), .C1(
        P1_U3086), .C2(n10613), .ZN(P1_U3345) );
  INV_X1 U11816 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n9984) );
  INV_X1 U11817 ( .A(n9979), .ZN(n9981) );
  INV_X1 U11818 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n9980) );
  NAND2_X1 U11819 ( .A1(n9981), .A2(n9980), .ZN(n10011) );
  NAND2_X1 U11820 ( .A1(n10011), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9982) );
  XNOR2_X1 U11821 ( .A(n9982), .B(P2_IR_REG_10__SCAN_IN), .ZN(n11091) );
  INV_X1 U11822 ( .A(n11091), .ZN(n10195) );
  OAI222_X1 U11823 ( .A1(n15545), .A2(n9984), .B1(n15540), .B2(n9983), .C1(
        P2_U3088), .C2(n10195), .ZN(P2_U3317) );
  INV_X1 U11824 ( .A(n14024), .ZN(n14008) );
  INV_X1 U11825 ( .A(SI_13_), .ZN(n14674) );
  OAI222_X1 U11826 ( .A1(n14008), .A2(P3_U3151), .B1(n14918), .B2(n9985), .C1(
        n14674), .C2(n14920), .ZN(P3_U3282) );
  INV_X1 U11827 ( .A(n10878), .ZN(n9986) );
  OR2_X1 U11828 ( .A1(n10389), .A2(P1_U3086), .ZN(n16137) );
  NAND2_X1 U11829 ( .A1(n9986), .A2(n16137), .ZN(n10018) );
  NAND2_X1 U11830 ( .A1(n10245), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9988) );
  NAND2_X1 U11831 ( .A1(n13607), .A2(n13608), .ZN(n13624) );
  INV_X1 U11832 ( .A(n13624), .ZN(n10402) );
  NAND3_X1 U11833 ( .A1(n9991), .A2(n9990), .A3(n9989), .ZN(n9992) );
  NOR2_X1 U11834 ( .A1(n9993), .A2(n9992), .ZN(n9994) );
  INV_X1 U11835 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n9995) );
  AOI21_X1 U11836 ( .B1(n10389), .B2(n10402), .A(n12759), .ZN(n10017) );
  INV_X1 U11837 ( .A(n10017), .ZN(n9998) );
  AND2_X1 U11838 ( .A1(n10018), .A2(n9998), .ZN(n16246) );
  NOR2_X1 U11839 ( .A1(n16246), .A2(P1_U4016), .ZN(P1_U3085) );
  INV_X1 U11840 ( .A(n9999), .ZN(n10000) );
  NAND2_X1 U11841 ( .A1(n10002), .A2(SI_10_), .ZN(n10003) );
  MUX2_X1 U11842 ( .A(n10010), .B(n10015), .S(n9874), .Z(n10004) );
  NAND2_X1 U11843 ( .A1(n10004), .A2(n14679), .ZN(n10139) );
  INV_X1 U11844 ( .A(n10004), .ZN(n10005) );
  NAND2_X1 U11845 ( .A1(n10005), .A2(SI_11_), .ZN(n10006) );
  NAND2_X1 U11846 ( .A1(n10139), .A2(n10006), .ZN(n10137) );
  XNOR2_X1 U11847 ( .A(n10136), .B(n10137), .ZN(n11851) );
  INV_X1 U11848 ( .A(n11851), .ZN(n10014) );
  INV_X1 U11849 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n10007) );
  NAND2_X1 U11850 ( .A1(n10008), .A2(n10007), .ZN(n10009) );
  NAND2_X1 U11851 ( .A1(n10009), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10145) );
  XNOR2_X1 U11852 ( .A(n10145), .B(P1_IR_REG_11__SCAN_IN), .ZN(n11852) );
  INV_X1 U11853 ( .A(n11852), .ZN(n10965) );
  OAI222_X1 U11854 ( .A1(n16139), .A2(n10010), .B1(n11886), .B2(n10014), .C1(
        P1_U3086), .C2(n10965), .ZN(P1_U3344) );
  OAI21_X1 U11855 ( .B1(n10011), .B2(P2_IR_REG_10__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n10012) );
  XNOR2_X1 U11856 ( .A(n10012), .B(P2_IR_REG_11__SCAN_IN), .ZN(n16184) );
  INV_X1 U11857 ( .A(n16184), .ZN(n10013) );
  OAI222_X1 U11858 ( .A1(n15545), .A2(n10015), .B1(n15540), .B2(n10014), .C1(
        P2_U3088), .C2(n10013), .ZN(P2_U3316) );
  OAI222_X1 U11859 ( .A1(P3_U3151), .A2(n14046), .B1(n14920), .B2(n14647), 
        .C1(n14918), .C2(n10016), .ZN(P3_U3281) );
  NAND2_X1 U11860 ( .A1(n10018), .A2(n10017), .ZN(n16249) );
  INV_X1 U11861 ( .A(n10409), .ZN(n10283) );
  INV_X1 U11862 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n16477) );
  AND2_X1 U11863 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n15696) );
  INV_X1 U11864 ( .A(n10364), .ZN(n15698) );
  NAND2_X1 U11865 ( .A1(n15698), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n10020) );
  NAND2_X1 U11866 ( .A1(n15695), .A2(n10020), .ZN(n10281) );
  XNOR2_X1 U11867 ( .A(n10409), .B(P1_REG1_REG_2__SCAN_IN), .ZN(n10282) );
  NAND2_X1 U11868 ( .A1(n10281), .A2(n10282), .ZN(n10280) );
  INV_X1 U11869 ( .A(n10280), .ZN(n10021) );
  XOR2_X1 U11870 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n10687), .Z(n10023) );
  NOR2_X1 U11871 ( .A1(n10024), .A2(n10023), .ZN(n10037) );
  INV_X1 U11872 ( .A(n7417), .ZN(n10022) );
  AOI211_X1 U11873 ( .C1(n10024), .C2(n10023), .A(n10037), .B(n15710), .ZN(
        n10033) );
  OR2_X1 U11874 ( .A1(n10019), .A2(n7417), .ZN(n10025) );
  INV_X1 U11875 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n10026) );
  MUX2_X1 U11876 ( .A(n10026), .B(P1_REG2_REG_1__SCAN_IN), .S(n10364), .Z(
        n15693) );
  AND2_X1 U11877 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n15694) );
  NAND2_X1 U11878 ( .A1(n15693), .A2(n15694), .ZN(n15692) );
  NAND2_X1 U11879 ( .A1(n15698), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n10027) );
  NAND2_X1 U11880 ( .A1(n15692), .A2(n10027), .ZN(n10278) );
  INV_X1 U11881 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n10885) );
  MUX2_X1 U11882 ( .A(n10885), .B(P1_REG2_REG_2__SCAN_IN), .S(n10409), .Z(
        n10279) );
  NAND2_X1 U11883 ( .A1(n10278), .A2(n10279), .ZN(n10277) );
  NAND2_X1 U11884 ( .A1(n10283), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n10030) );
  INV_X1 U11885 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n10028) );
  MUX2_X1 U11886 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n10028), .S(n10687), .Z(
        n10029) );
  AOI21_X1 U11887 ( .B1(n10277), .B2(n10030), .A(n10029), .ZN(n10296) );
  AND3_X1 U11888 ( .A1(n10277), .A2(n10030), .A3(n10029), .ZN(n10031) );
  NOR3_X1 U11889 ( .A1(n15728), .A2(n10296), .A3(n10031), .ZN(n10032) );
  NOR2_X1 U11890 ( .A1(n10033), .A2(n10032), .ZN(n10036) );
  AND2_X1 U11891 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n10034) );
  AOI21_X1 U11892 ( .B1(n16246), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n10034), .ZN(
        n10035) );
  OAI211_X1 U11893 ( .C1(n10687), .C2(n15727), .A(n10036), .B(n10035), .ZN(
        P1_U3246) );
  XNOR2_X1 U11894 ( .A(n10812), .B(P1_REG1_REG_6__SCAN_IN), .ZN(n10040) );
  INV_X1 U11895 ( .A(n10708), .ZN(n10041) );
  INV_X1 U11896 ( .A(n10687), .ZN(n10038) );
  AOI21_X1 U11897 ( .B1(P1_REG1_REG_3__SCAN_IN), .B2(n10038), .A(n10037), .ZN(
        n10292) );
  XOR2_X1 U11898 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n10708), .Z(n10291) );
  NOR2_X1 U11899 ( .A1(n10292), .A2(n10291), .ZN(n10290) );
  INV_X1 U11900 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n10715) );
  XNOR2_X1 U11901 ( .A(n10731), .B(n10715), .ZN(n10064) );
  NAND2_X1 U11902 ( .A1(n10063), .A2(n10064), .ZN(n10062) );
  OAI21_X1 U11903 ( .B1(n10731), .B2(P1_REG1_REG_5__SCAN_IN), .A(n10062), .ZN(
        n10039) );
  NOR2_X1 U11904 ( .A1(n10039), .A2(n10040), .ZN(n10155) );
  AOI211_X1 U11905 ( .C1(n10040), .C2(n10039), .A(n15710), .B(n10155), .ZN(
        n10048) );
  NOR2_X1 U11906 ( .A1(n10687), .A2(n10028), .ZN(n10295) );
  INV_X1 U11907 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n10695) );
  MUX2_X1 U11908 ( .A(n10695), .B(P1_REG2_REG_4__SCAN_IN), .S(n10708), .Z(
        n10294) );
  OAI21_X1 U11909 ( .B1(n10296), .B2(n10295), .A(n10294), .ZN(n10293) );
  NAND2_X1 U11910 ( .A1(n10041), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n10066) );
  INV_X1 U11911 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n10042) );
  MUX2_X1 U11912 ( .A(n10042), .B(P1_REG2_REG_5__SCAN_IN), .S(n10731), .Z(
        n10065) );
  AOI21_X1 U11913 ( .B1(n10293), .B2(n10066), .A(n10065), .ZN(n10068) );
  NOR2_X1 U11914 ( .A1(n10074), .A2(n10042), .ZN(n10044) );
  INV_X1 U11915 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n10739) );
  MUX2_X1 U11916 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n10739), .S(n10812), .Z(
        n10043) );
  OAI21_X1 U11917 ( .B1(n10068), .B2(n10044), .A(n10043), .ZN(n10161) );
  INV_X1 U11918 ( .A(n10161), .ZN(n10046) );
  NOR3_X1 U11919 ( .A1(n10068), .A2(n10044), .A3(n10043), .ZN(n10045) );
  NOR3_X1 U11920 ( .A1(n15728), .A2(n10046), .A3(n10045), .ZN(n10047) );
  NOR2_X1 U11921 ( .A1(n10048), .A2(n10047), .ZN(n10051) );
  NAND2_X1 U11922 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_U3086), .ZN(n10829) );
  INV_X1 U11923 ( .A(n10829), .ZN(n10049) );
  AOI21_X1 U11924 ( .B1(n16246), .B2(P1_ADDR_REG_6__SCAN_IN), .A(n10049), .ZN(
        n10050) );
  OAI211_X1 U11925 ( .C1(n10052), .C2(n15727), .A(n10051), .B(n10050), .ZN(
        P1_U3249) );
  INV_X1 U11926 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n13500) );
  XNOR2_X2 U11927 ( .A(n10250), .B(P1_IR_REG_30__SCAN_IN), .ZN(n10356) );
  INV_X1 U11928 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n10054) );
  NAND2_X1 U11929 ( .A1(n16120), .A2(n10355), .ZN(n10396) );
  INV_X1 U11930 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n10055) );
  OR2_X1 U11931 ( .A1(n12862), .A2(n10055), .ZN(n10060) );
  INV_X1 U11932 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n10056) );
  OR2_X1 U11933 ( .A1(n12929), .A2(n10056), .ZN(n10059) );
  NAND2_X2 U11934 ( .A1(n16120), .A2(n12655), .ZN(n10418) );
  INV_X1 U11935 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n10057) );
  OR2_X1 U11936 ( .A1(n7418), .A2(n10057), .ZN(n10058) );
  AND3_X1 U11937 ( .A1(n10060), .A2(n10059), .A3(n10058), .ZN(n15742) );
  INV_X1 U11938 ( .A(n15742), .ZN(n13615) );
  NAND2_X1 U11939 ( .A1(n13615), .A2(P1_U4016), .ZN(n10061) );
  OAI21_X1 U11940 ( .B1(P1_U4016), .B2(n13500), .A(n10061), .ZN(P1_U3591) );
  OAI21_X1 U11941 ( .B1(n10064), .B2(n10063), .A(n10062), .ZN(n10070) );
  AND3_X1 U11942 ( .A1(n10293), .A2(n10066), .A3(n10065), .ZN(n10067) );
  NOR3_X1 U11943 ( .A1(n15728), .A2(n10068), .A3(n10067), .ZN(n10069) );
  AOI21_X1 U11944 ( .B1(n16259), .B2(n10070), .A(n10069), .ZN(n10073) );
  AND2_X1 U11945 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n10071) );
  AOI21_X1 U11946 ( .B1(n16246), .B2(P1_ADDR_REG_5__SCAN_IN), .A(n10071), .ZN(
        n10072) );
  OAI211_X1 U11947 ( .C1(n10074), .C2(n15727), .A(n10073), .B(n10072), .ZN(
        P1_U3248) );
  INV_X1 U11948 ( .A(n13350), .ZN(n10075) );
  OR2_X1 U11949 ( .A1(n10076), .A2(n10075), .ZN(n10080) );
  NAND2_X1 U11950 ( .A1(n10077), .A2(n13350), .ZN(n10078) );
  NAND2_X1 U11951 ( .A1(n10078), .A2(n11062), .ZN(n10079) );
  NAND2_X1 U11952 ( .A1(n10080), .A2(n10079), .ZN(n10095) );
  AND2_X1 U11953 ( .A1(n10089), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10081) );
  INV_X1 U11954 ( .A(n15045), .ZN(n15057) );
  INV_X1 U11955 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10082) );
  MUX2_X1 U11956 ( .A(n10082), .B(P2_REG1_REG_1__SCAN_IN), .S(n10128), .Z(
        n10083) );
  NAND3_X1 U11957 ( .A1(n10083), .A2(P2_REG1_REG_0__SCAN_IN), .A3(
        P2_IR_REG_0__SCAN_IN), .ZN(n15054) );
  INV_X1 U11958 ( .A(n10128), .ZN(n10098) );
  NAND2_X1 U11959 ( .A1(n10098), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n15053) );
  INV_X1 U11960 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10084) );
  MUX2_X1 U11961 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n10084), .S(n15045), .Z(
        n15052) );
  AOI21_X1 U11962 ( .B1(n15054), .B2(n15053), .A(n15052), .ZN(n15051) );
  AOI21_X1 U11963 ( .B1(P2_REG1_REG_2__SCAN_IN), .B2(n15057), .A(n15051), .ZN(
        n16162) );
  INV_X1 U11964 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10085) );
  MUX2_X1 U11965 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n10085), .S(n10103), .Z(
        n16161) );
  OR2_X1 U11966 ( .A1(n16162), .A2(n16161), .ZN(n16164) );
  INV_X1 U11967 ( .A(n10103), .ZN(n16160) );
  NAND2_X1 U11968 ( .A1(n16160), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n15066) );
  INV_X1 U11969 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10086) );
  MUX2_X1 U11970 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n10086), .S(n15069), .Z(
        n15065) );
  AOI21_X1 U11971 ( .B1(n16164), .B2(n15066), .A(n15065), .ZN(n15088) );
  NOR2_X1 U11972 ( .A1(n15069), .A2(n10086), .ZN(n15084) );
  INV_X1 U11973 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n10087) );
  MUX2_X1 U11974 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n10087), .S(n15083), .Z(
        n10088) );
  OAI21_X1 U11975 ( .B1(n15088), .B2(n15084), .A(n10088), .ZN(n15100) );
  NAND2_X1 U11976 ( .A1(n15083), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n15099) );
  INV_X1 U11977 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n16592) );
  MUX2_X1 U11978 ( .A(n16592), .B(P2_REG1_REG_6__SCAN_IN), .S(n15105), .Z(
        n15098) );
  AOI21_X1 U11979 ( .B1(n15100), .B2(n15099), .A(n15098), .ZN(n15097) );
  AOI21_X1 U11980 ( .B1(P2_REG1_REG_6__SCAN_IN), .B2(n15105), .A(n15097), .ZN(
        n16174) );
  INV_X1 U11981 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n11322) );
  MUX2_X1 U11982 ( .A(n11322), .B(P2_REG1_REG_7__SCAN_IN), .S(n16172), .Z(
        n16173) );
  OR2_X1 U11983 ( .A1(n16174), .A2(n16173), .ZN(n16176) );
  NAND2_X1 U11984 ( .A1(n16172), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n10092) );
  INV_X1 U11985 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n16643) );
  MUX2_X1 U11986 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n16643), .S(n11063), .Z(
        n10091) );
  AOI21_X1 U11987 ( .B1(n16176), .B2(n10092), .A(n10091), .ZN(n10174) );
  INV_X1 U11988 ( .A(n10174), .ZN(n10094) );
  NOR2_X1 U11989 ( .A1(n10089), .A2(P2_U3088), .ZN(n15527) );
  AND2_X1 U11990 ( .A1(n10095), .A2(n15527), .ZN(n10116) );
  NAND2_X1 U11991 ( .A1(n10116), .A2(n10090), .ZN(n16190) );
  INV_X1 U11992 ( .A(n16190), .ZN(n16233) );
  NAND3_X1 U11993 ( .A1(n16176), .A2(n10092), .A3(n10091), .ZN(n10093) );
  NAND3_X1 U11994 ( .A1(n10094), .A2(n16233), .A3(n10093), .ZN(n10122) );
  NAND2_X1 U11995 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3088), .ZN(n12671) );
  INV_X1 U11996 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n11298) );
  MUX2_X1 U11997 ( .A(n11298), .B(P2_REG2_REG_1__SCAN_IN), .S(n10128), .Z(
        n10125) );
  AND2_X1 U11998 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n10097) );
  NAND2_X1 U11999 ( .A1(n10125), .A2(n10097), .ZN(n15048) );
  NAND2_X1 U12000 ( .A1(n10098), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n15047) );
  NAND2_X1 U12001 ( .A1(n15048), .A2(n15047), .ZN(n10101) );
  INV_X1 U12002 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n10099) );
  MUX2_X1 U12003 ( .A(n10099), .B(P2_REG2_REG_2__SCAN_IN), .S(n15045), .Z(
        n10100) );
  NAND2_X1 U12004 ( .A1(n10101), .A2(n10100), .ZN(n15050) );
  NAND2_X1 U12005 ( .A1(n15057), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n10102) );
  NAND2_X1 U12006 ( .A1(n15050), .A2(n10102), .ZN(n16167) );
  INV_X1 U12007 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n10104) );
  MUX2_X1 U12008 ( .A(n10104), .B(P2_REG2_REG_3__SCAN_IN), .S(n10103), .Z(
        n16166) );
  NAND2_X1 U12009 ( .A1(n16167), .A2(n16166), .ZN(n16165) );
  NAND2_X1 U12010 ( .A1(n16160), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n15071) );
  NAND2_X1 U12011 ( .A1(n16165), .A2(n15071), .ZN(n10106) );
  INV_X1 U12012 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n11289) );
  MUX2_X1 U12013 ( .A(n11289), .B(P2_REG2_REG_4__SCAN_IN), .S(n15069), .Z(
        n10105) );
  NAND2_X1 U12014 ( .A1(n10106), .A2(n10105), .ZN(n15081) );
  INV_X1 U12015 ( .A(n15069), .ZN(n10107) );
  NAND2_X1 U12016 ( .A1(n10107), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n15080) );
  NAND2_X1 U12017 ( .A1(n15081), .A2(n15080), .ZN(n10110) );
  INV_X1 U12018 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n10108) );
  MUX2_X1 U12019 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n10108), .S(n15083), .Z(
        n10109) );
  NAND2_X1 U12020 ( .A1(n10110), .A2(n10109), .ZN(n15094) );
  NAND2_X1 U12021 ( .A1(n15083), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n15093) );
  NAND2_X1 U12022 ( .A1(n15094), .A2(n15093), .ZN(n10112) );
  INV_X1 U12023 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n11273) );
  MUX2_X1 U12024 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n11273), .S(n15105), .Z(
        n10111) );
  NAND2_X1 U12025 ( .A1(n10112), .A2(n10111), .ZN(n15096) );
  NAND2_X1 U12026 ( .A1(n15105), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n10113) );
  NAND2_X1 U12027 ( .A1(n15096), .A2(n10113), .ZN(n16179) );
  INV_X1 U12028 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n11256) );
  MUX2_X1 U12029 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n11256), .S(n16172), .Z(
        n16178) );
  NAND2_X1 U12030 ( .A1(n16179), .A2(n16178), .ZN(n16177) );
  NAND2_X1 U12031 ( .A1(n16172), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n10114) );
  NAND2_X1 U12032 ( .A1(n16177), .A2(n10114), .ZN(n10118) );
  INV_X1 U12033 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n11647) );
  MUX2_X1 U12034 ( .A(n11647), .B(P2_REG2_REG_8__SCAN_IN), .S(n11063), .Z(
        n10117) );
  INV_X1 U12035 ( .A(n10090), .ZN(n10115) );
  AND2_X1 U12036 ( .A1(n10116), .A2(n10115), .ZN(n16229) );
  NAND2_X1 U12037 ( .A1(n10118), .A2(n10117), .ZN(n10170) );
  OAI211_X1 U12038 ( .C1(n10118), .C2(n10117), .A(n16229), .B(n10170), .ZN(
        n10119) );
  NAND2_X1 U12039 ( .A1(n12671), .A2(n10119), .ZN(n10120) );
  AOI21_X1 U12040 ( .B1(n10096), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n10120), .ZN(
        n10121) );
  OAI211_X1 U12041 ( .C1(n16214), .C2(n11063), .A(n10122), .B(n10121), .ZN(
        P2_U3222) );
  INV_X1 U12042 ( .A(n14063), .ZN(n14037) );
  OAI222_X1 U12043 ( .A1(P3_U3151), .A2(n14037), .B1(n14920), .B2(n10621), 
        .C1(n14918), .C2(n10123), .ZN(P3_U3280) );
  INV_X1 U12044 ( .A(n16229), .ZN(n16220) );
  INV_X1 U12045 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n10124) );
  NOR2_X1 U12046 ( .A1(n16220), .A2(n10124), .ZN(n16154) );
  AOI22_X1 U12047 ( .A1(n16154), .A2(P2_IR_REG_0__SCAN_IN), .B1(n16229), .B2(
        n10125), .ZN(n10135) );
  INV_X1 U12048 ( .A(n15048), .ZN(n10134) );
  NAND2_X1 U12049 ( .A1(P2_REG3_REG_1__SCAN_IN), .A2(P2_U3088), .ZN(n10126) );
  OAI21_X1 U12050 ( .B1(n16214), .B2(n10128), .A(n10126), .ZN(n10127) );
  AOI21_X1 U12051 ( .B1(n10096), .B2(P2_ADDR_REG_1__SCAN_IN), .A(n10127), .ZN(
        n10133) );
  INV_X1 U12052 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10236) );
  MUX2_X1 U12053 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n10082), .S(n10128), .Z(
        n10129) );
  OAI21_X1 U12054 ( .B1(n10236), .B2(n10130), .A(n10129), .ZN(n10131) );
  NAND3_X1 U12055 ( .A1(n16233), .A2(n15054), .A3(n10131), .ZN(n10132) );
  OAI211_X1 U12056 ( .C1(n10135), .C2(n10134), .A(n10133), .B(n10132), .ZN(
        P2_U3215) );
  INV_X1 U12057 ( .A(n10137), .ZN(n10138) );
  MUX2_X1 U12058 ( .A(n8078), .B(n10153), .S(n9874), .Z(n10141) );
  NAND2_X1 U12059 ( .A1(n10141), .A2(n14676), .ZN(n10215) );
  INV_X1 U12060 ( .A(n10141), .ZN(n10142) );
  NAND2_X1 U12061 ( .A1(n10142), .A2(SI_12_), .ZN(n10143) );
  XNOR2_X1 U12062 ( .A(n10214), .B(n8856), .ZN(n12000) );
  INV_X1 U12063 ( .A(n12000), .ZN(n10152) );
  INV_X1 U12064 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n10144) );
  NAND2_X1 U12065 ( .A1(n10145), .A2(n10144), .ZN(n10146) );
  NAND2_X1 U12066 ( .A1(n10146), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10217) );
  XNOR2_X1 U12067 ( .A(n10217), .B(P1_IR_REG_12__SCAN_IN), .ZN(n16262) );
  INV_X1 U12068 ( .A(n16262), .ZN(n10967) );
  OAI222_X1 U12069 ( .A1(n16139), .A2(n8078), .B1(n11886), .B2(n10152), .C1(
        n10967), .C2(P1_U3086), .ZN(P1_U3343) );
  NAND2_X1 U12070 ( .A1(n10148), .A2(n10147), .ZN(n10150) );
  NAND2_X1 U12071 ( .A1(n10150), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10149) );
  MUX2_X1 U12072 ( .A(P2_IR_REG_31__SCAN_IN), .B(n10149), .S(
        P2_IR_REG_12__SCAN_IN), .Z(n10151) );
  INV_X1 U12073 ( .A(n16232), .ZN(n10776) );
  OAI222_X1 U12074 ( .A1(n15545), .A2(n10153), .B1(n15540), .B2(n10152), .C1(
        n10776), .C2(P2_U3088), .ZN(P2_U3315) );
  NAND2_X1 U12075 ( .A1(n11008), .A2(n14899), .ZN(n10154) );
  OAI21_X1 U12076 ( .B1(n14899), .B2(n9403), .A(n10154), .ZN(P3_U3377) );
  INV_X1 U12077 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n10824) );
  MUX2_X1 U12078 ( .A(n10824), .B(P1_REG1_REG_7__SCAN_IN), .S(n11023), .Z(
        n10156) );
  NOR2_X1 U12079 ( .A1(n10157), .A2(n10156), .ZN(n10199) );
  AOI211_X1 U12080 ( .C1(n10157), .C2(n10156), .A(n15710), .B(n10199), .ZN(
        n10168) );
  INV_X1 U12081 ( .A(n15728), .ZN(n16263) );
  NAND2_X1 U12082 ( .A1(n10812), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n10160) );
  INV_X1 U12083 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n10158) );
  MUX2_X1 U12084 ( .A(n10158), .B(P1_REG2_REG_7__SCAN_IN), .S(n11023), .Z(
        n10159) );
  AOI21_X1 U12085 ( .B1(n10161), .B2(n10160), .A(n10159), .ZN(n10205) );
  INV_X1 U12086 ( .A(n10205), .ZN(n10163) );
  NAND3_X1 U12087 ( .A1(n10161), .A2(n10160), .A3(n10159), .ZN(n10162) );
  NAND3_X1 U12088 ( .A1(n16263), .A2(n10163), .A3(n10162), .ZN(n10166) );
  INV_X1 U12089 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n11035) );
  NOR2_X1 U12090 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n11035), .ZN(n10164) );
  AOI21_X1 U12091 ( .B1(n16246), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n10164), .ZN(
        n10165) );
  OAI211_X1 U12092 ( .C1(n15727), .C2(n10202), .A(n10166), .B(n10165), .ZN(
        n10167) );
  OR2_X1 U12093 ( .A1(n10168), .A2(n10167), .ZN(P1_U3250) );
  INV_X1 U12094 ( .A(n11063), .ZN(n10175) );
  NAND2_X1 U12095 ( .A1(n10175), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n10169) );
  NAND2_X1 U12096 ( .A1(n10170), .A2(n10169), .ZN(n10173) );
  INV_X1 U12097 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n10186) );
  MUX2_X1 U12098 ( .A(n10186), .B(P2_REG2_REG_9__SCAN_IN), .S(n11078), .Z(
        n10172) );
  OR2_X1 U12099 ( .A1(n10173), .A2(n10172), .ZN(n10189) );
  INV_X1 U12100 ( .A(n10189), .ZN(n10171) );
  AOI21_X1 U12101 ( .B1(n10173), .B2(n10172), .A(n10171), .ZN(n10182) );
  AOI21_X1 U12102 ( .B1(n10175), .B2(P2_REG1_REG_8__SCAN_IN), .A(n10174), .ZN(
        n10177) );
  INV_X1 U12103 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n11629) );
  MUX2_X1 U12104 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n11629), .S(n11078), .Z(
        n10176) );
  NAND2_X1 U12105 ( .A1(n10177), .A2(n10176), .ZN(n10183) );
  OAI21_X1 U12106 ( .B1(n10177), .B2(n10176), .A(n10183), .ZN(n10180) );
  NAND2_X1 U12107 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3088), .ZN(n12661) );
  NAND2_X1 U12108 ( .A1(n10096), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n10178) );
  OAI211_X1 U12109 ( .C1(n16214), .C2(n10187), .A(n12661), .B(n10178), .ZN(
        n10179) );
  AOI21_X1 U12110 ( .B1(n10180), .B2(n16233), .A(n10179), .ZN(n10181) );
  OAI21_X1 U12111 ( .B1(n10182), .B2(n16220), .A(n10181), .ZN(P2_U3223) );
  OAI21_X1 U12112 ( .B1(n11078), .B2(P2_REG1_REG_9__SCAN_IN), .A(n10183), .ZN(
        n10185) );
  INV_X1 U12113 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n16683) );
  MUX2_X1 U12114 ( .A(n16683), .B(P2_REG1_REG_10__SCAN_IN), .S(n11091), .Z(
        n10184) );
  NOR2_X1 U12115 ( .A1(n10185), .A2(n10184), .ZN(n10774) );
  AOI211_X1 U12116 ( .C1(n10185), .C2(n10184), .A(n16190), .B(n10774), .ZN(
        n10198) );
  NAND2_X1 U12117 ( .A1(n10187), .A2(n10186), .ZN(n10188) );
  NAND2_X1 U12118 ( .A1(n10189), .A2(n10188), .ZN(n10193) );
  INV_X1 U12119 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n10190) );
  MUX2_X1 U12120 ( .A(n10190), .B(P2_REG2_REG_10__SCAN_IN), .S(n11091), .Z(
        n10192) );
  OR2_X1 U12121 ( .A1(n10193), .A2(n10192), .ZN(n10766) );
  INV_X1 U12122 ( .A(n10766), .ZN(n10191) );
  AOI211_X1 U12123 ( .C1(n10193), .C2(n10192), .A(n16220), .B(n10191), .ZN(
        n10197) );
  NAND2_X1 U12124 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3088), .ZN(n11107)
         );
  NAND2_X1 U12125 ( .A1(n10096), .A2(P2_ADDR_REG_10__SCAN_IN), .ZN(n10194) );
  OAI211_X1 U12126 ( .C1(n16214), .C2(n10195), .A(n11107), .B(n10194), .ZN(
        n10196) );
  OR3_X1 U12127 ( .A1(n10198), .A2(n10197), .A3(n10196), .ZN(P2_U3224) );
  AOI21_X1 U12128 ( .B1(n11023), .B2(P1_REG1_REG_7__SCAN_IN), .A(n10199), .ZN(
        n10201) );
  INV_X1 U12129 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n11027) );
  MUX2_X1 U12130 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n11027), .S(n11540), .Z(
        n10200) );
  NAND2_X1 U12131 ( .A1(n10201), .A2(n10200), .ZN(n10309) );
  OAI21_X1 U12132 ( .B1(n10201), .B2(n10200), .A(n10309), .ZN(n10212) );
  NOR2_X1 U12133 ( .A1(n10202), .A2(n10158), .ZN(n10204) );
  INV_X1 U12134 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n16624) );
  MUX2_X1 U12135 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n16624), .S(n11540), .Z(
        n10203) );
  OAI21_X1 U12136 ( .B1(n10205), .B2(n10204), .A(n10203), .ZN(n10307) );
  INV_X1 U12137 ( .A(n10307), .ZN(n10207) );
  NOR3_X1 U12138 ( .A1(n10205), .A2(n10204), .A3(n10203), .ZN(n10206) );
  NOR3_X1 U12139 ( .A1(n15728), .A2(n10207), .A3(n10206), .ZN(n10211) );
  NAND2_X1 U12140 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n11711) );
  NAND2_X1 U12141 ( .A1(n16246), .A2(P1_ADDR_REG_8__SCAN_IN), .ZN(n10208) );
  OAI211_X1 U12142 ( .C1(n15727), .C2(n10209), .A(n11711), .B(n10208), .ZN(
        n10210) );
  AOI211_X1 U12143 ( .C1(n10212), .C2(n16259), .A(n10211), .B(n10210), .ZN(
        n10213) );
  INV_X1 U12144 ( .A(n10213), .ZN(P1_U3251) );
  MUX2_X1 U12145 ( .A(n12005), .B(n10221), .S(n13247), .Z(n10445) );
  XNOR2_X1 U12146 ( .A(n10445), .B(SI_13_), .ZN(n10444) );
  XNOR2_X1 U12147 ( .A(n10448), .B(n10444), .ZN(n12004) );
  INV_X1 U12148 ( .A(n12004), .ZN(n10220) );
  INV_X1 U12149 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n10216) );
  NAND2_X1 U12150 ( .A1(n10217), .A2(n10216), .ZN(n10218) );
  NAND2_X1 U12151 ( .A1(n10218), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10453) );
  XNOR2_X1 U12152 ( .A(n10453), .B(P1_IR_REG_13__SCAN_IN), .ZN(n12007) );
  INV_X1 U12153 ( .A(n12007), .ZN(n11473) );
  OAI222_X1 U12154 ( .A1(n16139), .A2(n12005), .B1(n11886), .B2(n10220), .C1(
        n11473), .C2(P1_U3086), .ZN(P1_U3342) );
  NAND2_X1 U12155 ( .A1(n10449), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10219) );
  XNOR2_X1 U12156 ( .A(n10219), .B(P2_IR_REG_13__SCAN_IN), .ZN(n11784) );
  INV_X1 U12157 ( .A(n11784), .ZN(n10800) );
  OAI222_X1 U12158 ( .A1(n15545), .A2(n10221), .B1(n15540), .B2(n10220), .C1(
        n10800), .C2(P2_U3088), .ZN(P2_U3314) );
  NAND2_X1 U12159 ( .A1(n10223), .A2(n10222), .ZN(n11245) );
  INV_X1 U12160 ( .A(n16148), .ZN(n16152) );
  NOR2_X1 U12161 ( .A1(n16152), .A2(n11243), .ZN(n16145) );
  NAND2_X1 U12162 ( .A1(n16145), .A2(n10224), .ZN(n10225) );
  OAI21_X1 U12163 ( .B1(n13013), .B2(n10984), .A(n10545), .ZN(n13308) );
  NAND2_X1 U12164 ( .A1(n13307), .A2(n13342), .ZN(n10228) );
  NAND2_X1 U12165 ( .A1(n8082), .A2(n13341), .ZN(n10227) );
  AND2_X1 U12166 ( .A1(n10226), .A2(n15308), .ZN(n10229) );
  OR2_X1 U12167 ( .A1(n13308), .A2(n10229), .ZN(n10231) );
  NAND2_X1 U12168 ( .A1(n15043), .A2(n15343), .ZN(n10230) );
  NAND2_X1 U12169 ( .A1(n10231), .A2(n10230), .ZN(n11413) );
  INV_X1 U12170 ( .A(n10232), .ZN(n10233) );
  NOR2_X1 U12171 ( .A1(n10233), .A2(n13012), .ZN(n10234) );
  NOR2_X1 U12172 ( .A1(n11413), .A2(n10234), .ZN(n11414) );
  OAI21_X1 U12173 ( .B1(n16590), .B2(n13308), .A(n11414), .ZN(n10241) );
  NAND2_X1 U12174 ( .A1(n16747), .A2(n10241), .ZN(n10235) );
  OAI21_X1 U12175 ( .B1(n16747), .B2(n10236), .A(n10235), .ZN(P2_U3499) );
  INV_X1 U12176 ( .A(n10237), .ZN(n10238) );
  OAI222_X1 U12177 ( .A1(P3_U3151), .A2(n14083), .B1(n14920), .B2(n11160), 
        .C1(n14918), .C2(n10238), .ZN(P3_U3279) );
  INV_X1 U12178 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n10243) );
  NAND2_X1 U12179 ( .A1(n16751), .A2(n10241), .ZN(n10242) );
  OAI21_X1 U12180 ( .B1(n16751), .B2(n10243), .A(n10242), .ZN(P2_U3430) );
  NAND2_X1 U12181 ( .A1(n9554), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10244) );
  MUX2_X1 U12182 ( .A(P1_IR_REG_31__SCAN_IN), .B(n10244), .S(
        P1_IR_REG_20__SCAN_IN), .Z(n10246) );
  NAND2_X1 U12183 ( .A1(n13608), .A2(n13610), .ZN(n13660) );
  NAND2_X1 U12184 ( .A1(n10384), .A2(n13610), .ZN(n13623) );
  INV_X1 U12185 ( .A(n13623), .ZN(n10429) );
  INV_X1 U12186 ( .A(n10247), .ZN(n10248) );
  NAND2_X1 U12187 ( .A1(n10248), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10249) );
  OR2_X1 U12188 ( .A1(n16464), .A2(n13606), .ZN(n12329) );
  INV_X1 U12189 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n16115) );
  AOI22_X1 U12190 ( .A1(n16115), .A2(P1_REG2_REG_0__SCAN_IN), .B1(
        P1_IR_REG_30__SCAN_IN), .B2(P1_REG0_REG_0__SCAN_IN), .ZN(n10255) );
  INV_X1 U12191 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n10252) );
  NAND2_X1 U12192 ( .A1(P1_REG2_REG_0__SCAN_IN), .A2(P1_IR_REG_30__SCAN_IN), 
        .ZN(n10251) );
  OAI21_X1 U12193 ( .B1(n10252), .B2(P1_IR_REG_30__SCAN_IN), .A(n10251), .ZN(
        n10253) );
  NAND2_X1 U12194 ( .A1(n10250), .A2(n10253), .ZN(n10254) );
  OAI21_X1 U12195 ( .B1(n10250), .B2(n10255), .A(n10254), .ZN(n10256) );
  NAND2_X1 U12196 ( .A1(n10256), .A2(n12655), .ZN(n10264) );
  AOI22_X1 U12197 ( .A1(n16115), .A2(P1_REG3_REG_0__SCAN_IN), .B1(
        P1_REG1_REG_0__SCAN_IN), .B2(P1_IR_REG_30__SCAN_IN), .ZN(n10261) );
  INV_X1 U12198 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n10258) );
  NAND2_X1 U12199 ( .A1(P1_IR_REG_30__SCAN_IN), .A2(P1_REG3_REG_0__SCAN_IN), 
        .ZN(n10257) );
  OAI21_X1 U12200 ( .B1(n10258), .B2(P1_IR_REG_30__SCAN_IN), .A(n10257), .ZN(
        n10259) );
  NAND2_X1 U12201 ( .A1(n10250), .A2(n10259), .ZN(n10260) );
  OAI21_X1 U12202 ( .B1(n10250), .B2(n10261), .A(n10260), .ZN(n10262) );
  NAND2_X1 U12203 ( .A1(n10262), .A2(n10355), .ZN(n10263) );
  NAND2_X1 U12204 ( .A1(n10264), .A2(n10263), .ZN(n15691) );
  INV_X1 U12205 ( .A(n15691), .ZN(n10265) );
  INV_X1 U12206 ( .A(n13660), .ZN(n10432) );
  INV_X1 U12207 ( .A(SI_0_), .ZN(n10267) );
  OAI21_X1 U12208 ( .B1(n7416), .B2(n10267), .A(n10266), .ZN(n10268) );
  NAND2_X1 U12209 ( .A1(n10269), .A2(n10268), .ZN(n16142) );
  MUX2_X1 U12210 ( .A(n8830), .B(n16142), .S(n12814), .Z(n15990) );
  OAI22_X1 U12211 ( .A1(n10271), .A2(n15990), .B1(n8830), .B2(n10392), .ZN(
        n10270) );
  NAND2_X1 U12212 ( .A1(n7413), .A2(n15691), .ZN(n10274) );
  INV_X1 U12213 ( .A(n10392), .ZN(n10272) );
  NAND2_X1 U12214 ( .A1(n10272), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n10273) );
  MUX2_X1 U12215 ( .A(n15694), .B(n12649), .S(n7417), .Z(n10276) );
  NOR2_X1 U12216 ( .A1(n7417), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n10275) );
  NOR2_X1 U12217 ( .A1(n10275), .A2(n10019), .ZN(n16241) );
  NOR2_X1 U12218 ( .A1(n16241), .A2(P1_IR_REG_0__SCAN_IN), .ZN(n16239) );
  AOI211_X1 U12219 ( .C1(n10276), .C2(n10401), .A(n16239), .B(n15677), .ZN(
        n10303) );
  OAI211_X1 U12220 ( .C1(n10279), .C2(n10278), .A(n16263), .B(n10277), .ZN(
        n10287) );
  OAI211_X1 U12221 ( .C1(n10282), .C2(n10281), .A(n16259), .B(n10280), .ZN(
        n10286) );
  AOI22_X1 U12222 ( .A1(n16246), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n10285) );
  NAND2_X1 U12223 ( .A1(n16261), .A2(n10283), .ZN(n10284) );
  NAND4_X1 U12224 ( .A1(n10287), .A2(n10286), .A3(n10285), .A4(n10284), .ZN(
        n10288) );
  OR2_X1 U12225 ( .A1(n10303), .A2(n10288), .ZN(P1_U3245) );
  OAI222_X1 U12226 ( .A1(P3_U3151), .A2(n14108), .B1(n14920), .B2(n11162), 
        .C1(n14918), .C2(n10289), .ZN(P3_U3278) );
  AOI211_X1 U12227 ( .C1(n10292), .C2(n10291), .A(n10290), .B(n15710), .ZN(
        n10302) );
  INV_X1 U12228 ( .A(n10293), .ZN(n10298) );
  NOR3_X1 U12229 ( .A1(n10296), .A2(n10295), .A3(n10294), .ZN(n10297) );
  NOR3_X1 U12230 ( .A1(n15728), .A2(n10298), .A3(n10297), .ZN(n10301) );
  NAND2_X1 U12231 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n10725) );
  NAND2_X1 U12232 ( .A1(n16246), .A2(P1_ADDR_REG_4__SCAN_IN), .ZN(n10299) );
  OAI211_X1 U12233 ( .C1(n15727), .C2(n10708), .A(n10725), .B(n10299), .ZN(
        n10300) );
  OR4_X1 U12234 ( .A1(n10303), .A2(n10302), .A3(n10301), .A4(n10300), .ZN(
        P1_U3247) );
  NAND2_X1 U12235 ( .A1(n11540), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n10306) );
  INV_X1 U12236 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n10304) );
  MUX2_X1 U12237 ( .A(n10304), .B(P1_REG2_REG_9__SCAN_IN), .S(n11546), .Z(
        n10305) );
  AOI21_X1 U12238 ( .B1(n10307), .B2(n10306), .A(n10305), .ZN(n10608) );
  NAND3_X1 U12239 ( .A1(n10307), .A2(n10306), .A3(n10305), .ZN(n10308) );
  NAND2_X1 U12240 ( .A1(n16263), .A2(n10308), .ZN(n10317) );
  INV_X1 U12241 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n11549) );
  MUX2_X1 U12242 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n11549), .S(n11546), .Z(
        n10311) );
  OAI21_X1 U12243 ( .B1(n11540), .B2(P1_REG1_REG_8__SCAN_IN), .A(n10309), .ZN(
        n10310) );
  NAND2_X1 U12244 ( .A1(n10310), .A2(n10311), .ZN(n10602) );
  OAI21_X1 U12245 ( .B1(n10311), .B2(n10310), .A(n10602), .ZN(n10312) );
  NAND2_X1 U12246 ( .A1(n10312), .A2(n16259), .ZN(n10316) );
  INV_X1 U12247 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n11704) );
  NOR2_X1 U12248 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n11704), .ZN(n10314) );
  NOR2_X1 U12249 ( .A1(n15727), .A2(n10605), .ZN(n10313) );
  AOI211_X1 U12250 ( .C1(n16246), .C2(P1_ADDR_REG_9__SCAN_IN), .A(n10314), .B(
        n10313), .ZN(n10315) );
  OAI211_X1 U12251 ( .C1(n10608), .C2(n10317), .A(n10316), .B(n10315), .ZN(
        P1_U3252) );
  NOR2_X1 U12252 ( .A1(n10319), .A2(n10318), .ZN(n10321) );
  INV_X1 U12253 ( .A(P3_D_REG_25__SCAN_IN), .ZN(n10320) );
  NOR2_X1 U12254 ( .A1(n10348), .A2(n10320), .ZN(P3_U3240) );
  CLKBUF_X1 U12255 ( .A(n10321), .Z(n10348) );
  INV_X1 U12256 ( .A(P3_D_REG_2__SCAN_IN), .ZN(n10322) );
  NOR2_X1 U12257 ( .A1(n10348), .A2(n10322), .ZN(P3_U3263) );
  INV_X1 U12258 ( .A(P3_D_REG_7__SCAN_IN), .ZN(n10323) );
  NOR2_X1 U12259 ( .A1(n10321), .A2(n10323), .ZN(P3_U3258) );
  INV_X1 U12260 ( .A(P3_D_REG_28__SCAN_IN), .ZN(n10324) );
  NOR2_X1 U12261 ( .A1(n10321), .A2(n10324), .ZN(P3_U3237) );
  INV_X1 U12262 ( .A(P3_D_REG_11__SCAN_IN), .ZN(n10325) );
  NOR2_X1 U12263 ( .A1(n10348), .A2(n10325), .ZN(P3_U3254) );
  INV_X1 U12264 ( .A(P3_D_REG_14__SCAN_IN), .ZN(n10326) );
  NOR2_X1 U12265 ( .A1(n10348), .A2(n10326), .ZN(P3_U3251) );
  INV_X1 U12266 ( .A(P3_D_REG_16__SCAN_IN), .ZN(n10327) );
  NOR2_X1 U12267 ( .A1(n10348), .A2(n10327), .ZN(P3_U3249) );
  INV_X1 U12268 ( .A(P3_D_REG_24__SCAN_IN), .ZN(n10328) );
  NOR2_X1 U12269 ( .A1(n10321), .A2(n10328), .ZN(P3_U3241) );
  INV_X1 U12270 ( .A(P3_D_REG_30__SCAN_IN), .ZN(n10329) );
  NOR2_X1 U12271 ( .A1(n10321), .A2(n10329), .ZN(P3_U3235) );
  INV_X1 U12272 ( .A(P3_D_REG_10__SCAN_IN), .ZN(n10330) );
  NOR2_X1 U12273 ( .A1(n10348), .A2(n10330), .ZN(P3_U3255) );
  INV_X1 U12274 ( .A(P3_D_REG_9__SCAN_IN), .ZN(n10331) );
  NOR2_X1 U12275 ( .A1(n10348), .A2(n10331), .ZN(P3_U3256) );
  INV_X1 U12276 ( .A(P3_D_REG_23__SCAN_IN), .ZN(n10332) );
  NOR2_X1 U12277 ( .A1(n10321), .A2(n10332), .ZN(P3_U3242) );
  INV_X1 U12278 ( .A(P3_D_REG_13__SCAN_IN), .ZN(n10333) );
  NOR2_X1 U12279 ( .A1(n10348), .A2(n10333), .ZN(P3_U3252) );
  INV_X1 U12280 ( .A(P3_D_REG_21__SCAN_IN), .ZN(n10334) );
  NOR2_X1 U12281 ( .A1(n10321), .A2(n10334), .ZN(P3_U3244) );
  INV_X1 U12282 ( .A(P3_D_REG_20__SCAN_IN), .ZN(n10335) );
  NOR2_X1 U12283 ( .A1(n10321), .A2(n10335), .ZN(P3_U3245) );
  INV_X1 U12284 ( .A(P3_D_REG_19__SCAN_IN), .ZN(n10336) );
  NOR2_X1 U12285 ( .A1(n10348), .A2(n10336), .ZN(P3_U3246) );
  INV_X1 U12286 ( .A(P3_D_REG_18__SCAN_IN), .ZN(n10337) );
  NOR2_X1 U12287 ( .A1(n10348), .A2(n10337), .ZN(P3_U3247) );
  INV_X1 U12288 ( .A(P3_D_REG_17__SCAN_IN), .ZN(n10338) );
  NOR2_X1 U12289 ( .A1(n10348), .A2(n10338), .ZN(P3_U3248) );
  INV_X1 U12290 ( .A(P3_D_REG_29__SCAN_IN), .ZN(n10339) );
  NOR2_X1 U12291 ( .A1(n10321), .A2(n10339), .ZN(P3_U3236) );
  INV_X1 U12292 ( .A(P3_D_REG_12__SCAN_IN), .ZN(n10340) );
  NOR2_X1 U12293 ( .A1(n10348), .A2(n10340), .ZN(P3_U3253) );
  INV_X1 U12294 ( .A(P3_D_REG_8__SCAN_IN), .ZN(n10341) );
  NOR2_X1 U12295 ( .A1(n10348), .A2(n10341), .ZN(P3_U3257) );
  INV_X1 U12296 ( .A(P3_D_REG_31__SCAN_IN), .ZN(n10342) );
  NOR2_X1 U12297 ( .A1(n10321), .A2(n10342), .ZN(P3_U3234) );
  INV_X1 U12298 ( .A(P3_D_REG_6__SCAN_IN), .ZN(n10343) );
  NOR2_X1 U12299 ( .A1(n10348), .A2(n10343), .ZN(P3_U3259) );
  INV_X1 U12300 ( .A(P3_D_REG_5__SCAN_IN), .ZN(n10344) );
  NOR2_X1 U12301 ( .A1(n10321), .A2(n10344), .ZN(P3_U3260) );
  INV_X1 U12302 ( .A(P3_D_REG_4__SCAN_IN), .ZN(n10345) );
  NOR2_X1 U12303 ( .A1(n10348), .A2(n10345), .ZN(P3_U3261) );
  INV_X1 U12304 ( .A(P3_D_REG_27__SCAN_IN), .ZN(n10346) );
  NOR2_X1 U12305 ( .A1(n10321), .A2(n10346), .ZN(P3_U3238) );
  INV_X1 U12306 ( .A(P3_D_REG_15__SCAN_IN), .ZN(n10347) );
  NOR2_X1 U12307 ( .A1(n10348), .A2(n10347), .ZN(P3_U3250) );
  INV_X1 U12308 ( .A(P3_D_REG_22__SCAN_IN), .ZN(n10349) );
  NOR2_X1 U12309 ( .A1(n10348), .A2(n10349), .ZN(P3_U3243) );
  INV_X1 U12310 ( .A(P3_D_REG_26__SCAN_IN), .ZN(n10350) );
  NOR2_X1 U12311 ( .A1(n10348), .A2(n10350), .ZN(P3_U3239) );
  INV_X1 U12312 ( .A(P3_D_REG_3__SCAN_IN), .ZN(n10351) );
  NOR2_X1 U12313 ( .A1(n10348), .A2(n10351), .ZN(P3_U3262) );
  NAND2_X1 U12314 ( .A1(n13607), .A2(n15733), .ZN(n10352) );
  OAI21_X1 U12315 ( .B1(n10354), .B2(n10817), .A(n10353), .ZN(n10416) );
  NAND2_X1 U12316 ( .A1(n7420), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n10361) );
  NAND2_X1 U12317 ( .A1(n12802), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n10360) );
  INV_X1 U12318 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n10357) );
  OR2_X1 U12319 ( .A1(n10418), .A2(n10357), .ZN(n10359) );
  OR2_X1 U12320 ( .A1(n10396), .A2(n16477), .ZN(n10358) );
  INV_X1 U12321 ( .A(n10704), .ZN(n10362) );
  OAI22_X1 U12322 ( .A1(n13667), .A2(n10271), .B1(n16480), .B2(n12940), .ZN(
        n10365) );
  XNOR2_X1 U12323 ( .A(n10365), .B(n10817), .ZN(n10414) );
  OAI22_X1 U12324 ( .A1(n12846), .A2(n13667), .B1(n16480), .B2(n10271), .ZN(
        n10415) );
  XNOR2_X1 U12325 ( .A(n10414), .B(n10415), .ZN(n10417) );
  XOR2_X1 U12326 ( .A(n10416), .B(n10417), .Z(n10406) );
  OAI21_X1 U12327 ( .B1(n10381), .B2(P1_D_REG_1__SCAN_IN), .A(n10366), .ZN(
        n10873) );
  NOR4_X1 U12328 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n10370) );
  NOR4_X1 U12329 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n10369) );
  NOR4_X1 U12330 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n10368) );
  NOR4_X1 U12331 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n10367) );
  NAND4_X1 U12332 ( .A1(n10370), .A2(n10369), .A3(n10368), .A4(n10367), .ZN(
        n10376) );
  NOR2_X1 U12333 ( .A1(P1_D_REG_31__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .ZN(
        n10374) );
  NOR4_X1 U12334 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_29__SCAN_IN), .A4(P1_D_REG_28__SCAN_IN), .ZN(n10373) );
  NOR4_X1 U12335 ( .A1(P1_D_REG_23__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_21__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n10372) );
  NOR4_X1 U12336 ( .A1(P1_D_REG_27__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_25__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n10371) );
  NAND4_X1 U12337 ( .A1(n10374), .A2(n10373), .A3(n10372), .A4(n10371), .ZN(
        n10375) );
  NOR2_X1 U12338 ( .A1(n10376), .A2(n10375), .ZN(n10377) );
  OR2_X1 U12339 ( .A1(n10381), .A2(n10377), .ZN(n10874) );
  INV_X1 U12340 ( .A(n10874), .ZN(n10378) );
  NOR2_X1 U12341 ( .A1(n10873), .A2(n10378), .ZN(n10383) );
  INV_X1 U12342 ( .A(n10379), .ZN(n16132) );
  INV_X1 U12343 ( .A(n10380), .ZN(n16127) );
  NAND2_X1 U12344 ( .A1(n16132), .A2(n16127), .ZN(n16114) );
  INV_X1 U12345 ( .A(n11137), .ZN(n10382) );
  NAND2_X1 U12346 ( .A1(n10383), .A2(n10382), .ZN(n10393) );
  INV_X1 U12347 ( .A(n13610), .ZN(n13614) );
  NAND2_X1 U12348 ( .A1(n15988), .A2(n13614), .ZN(n13803) );
  INV_X1 U12349 ( .A(n13803), .ZN(n10385) );
  NAND2_X1 U12350 ( .A1(n10384), .A2(n10385), .ZN(n10879) );
  NAND3_X1 U12351 ( .A1(n10878), .A2(n16725), .A3(n13624), .ZN(n10386) );
  NAND2_X1 U12352 ( .A1(n10393), .A2(n10876), .ZN(n10713) );
  NAND2_X1 U12353 ( .A1(n13607), .A2(n13606), .ZN(n10388) );
  NAND2_X1 U12354 ( .A1(n13608), .A2(n13614), .ZN(n10387) );
  NAND2_X1 U12355 ( .A1(n16561), .A2(n10402), .ZN(n10390) );
  AND2_X1 U12356 ( .A1(n10390), .A2(n10389), .ZN(n10391) );
  AND2_X1 U12357 ( .A1(n10392), .A2(n10391), .ZN(n10712) );
  NAND2_X1 U12358 ( .A1(n10712), .A2(P1_STATE_REG_SCAN_IN), .ZN(n13804) );
  INV_X1 U12359 ( .A(n13804), .ZN(n11136) );
  NAND2_X1 U12360 ( .A1(n10713), .A2(n11136), .ZN(n12647) );
  OR2_X1 U12361 ( .A1(n10393), .A2(n13804), .ZN(n15638) );
  INV_X1 U12362 ( .A(n16462), .ZN(n15953) );
  NOR2_X1 U12363 ( .A1(n15638), .A2(n15953), .ZN(n15658) );
  NAND2_X1 U12364 ( .A1(n7420), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n10400) );
  INV_X1 U12365 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n10880) );
  OR2_X1 U12366 ( .A1(n12946), .A2(n10880), .ZN(n10399) );
  INV_X1 U12367 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n10394) );
  OR2_X1 U12368 ( .A1(n7418), .A2(n10394), .ZN(n10398) );
  INV_X1 U12369 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10395) );
  OR2_X1 U12370 ( .A1(n10396), .A2(n10395), .ZN(n10397) );
  NAND2_X1 U12371 ( .A1(n15971), .A2(n15691), .ZN(n16469) );
  OAI22_X1 U12372 ( .A1(n15648), .A2(n8047), .B1(n16469), .B2(n15638), .ZN(
        n10404) );
  AND2_X1 U12373 ( .A1(n10713), .A2(n10878), .ZN(n16528) );
  INV_X1 U12374 ( .A(n15671), .ZN(n15653) );
  NOR2_X1 U12375 ( .A1(n15653), .A2(n16480), .ZN(n10403) );
  AOI211_X1 U12376 ( .C1(P1_REG3_REG_1__SCAN_IN), .C2(n12647), .A(n10404), .B(
        n10403), .ZN(n10405) );
  OAI21_X1 U12377 ( .B1(n10406), .B2(n15673), .A(n10405), .ZN(P1_U3222) );
  OR2_X1 U12378 ( .A1(n10704), .A2(n10407), .ZN(n10412) );
  OR2_X1 U12379 ( .A1(n10702), .A2(n10408), .ZN(n10411) );
  OR2_X1 U12380 ( .A1(n12814), .A2(n10409), .ZN(n10410) );
  AND3_X2 U12381 ( .A1(n10412), .A2(n10411), .A3(n10410), .ZN(n10934) );
  OAI22_X1 U12382 ( .A1(n12846), .A2(n8047), .B1(n10934), .B2(n10271), .ZN(
        n10678) );
  OAI22_X1 U12383 ( .A1(n8047), .A2(n10271), .B1(n10934), .B2(n12940), .ZN(
        n10413) );
  XNOR2_X1 U12384 ( .A(n10413), .B(n10817), .ZN(n10677) );
  XOR2_X1 U12385 ( .A(n10678), .B(n10677), .Z(n10681) );
  OAI22_X1 U12386 ( .A1(n10417), .A2(n10416), .B1(n10415), .B2(n10414), .ZN(
        n10682) );
  XOR2_X1 U12387 ( .A(n10682), .B(n10681), .Z(n10428) );
  NOR2_X1 U12388 ( .A1(n15653), .A2(n10934), .ZN(n10426) );
  NOR2_X2 U12389 ( .A1(n15638), .A2(n15951), .ZN(n15659) );
  INV_X1 U12390 ( .A(n15659), .ZN(n10424) );
  NAND2_X1 U12391 ( .A1(n13566), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n10423) );
  OR2_X1 U12392 ( .A1(n12946), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n10422) );
  INV_X1 U12393 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n10419) );
  OR2_X1 U12394 ( .A1(n10396), .A2(n10419), .ZN(n10420) );
  OAI22_X1 U12395 ( .A1(n13667), .A2(n10424), .B1(n15648), .B2(n13655), .ZN(
        n10425) );
  AOI211_X1 U12396 ( .C1(P1_REG3_REG_2__SCAN_IN), .C2(n12647), .A(n10426), .B(
        n10425), .ZN(n10427) );
  OAI21_X1 U12397 ( .B1(n15673), .B2(n10428), .A(n10427), .ZN(P1_U3237) );
  NAND2_X1 U12398 ( .A1(n10429), .A2(n13606), .ZN(n16475) );
  INV_X1 U12399 ( .A(n16475), .ZN(n16660) );
  NAND2_X1 U12400 ( .A1(n10430), .A2(n16466), .ZN(n10431) );
  INV_X1 U12401 ( .A(n15990), .ZN(n16465) );
  AND2_X1 U12402 ( .A1(n16465), .A2(n15691), .ZN(n16461) );
  NAND2_X1 U12403 ( .A1(n13665), .A2(n13668), .ZN(n10932) );
  XNOR2_X1 U12404 ( .A(n10933), .B(n13575), .ZN(n10888) );
  INV_X1 U12405 ( .A(n10888), .ZN(n10441) );
  OAI211_X1 U12406 ( .C1(n7458), .C2(n10934), .A(n16079), .B(n10940), .ZN(
        n10881) );
  OAI21_X1 U12407 ( .B1(n10934), .B2(n16725), .A(n10881), .ZN(n10440) );
  NAND2_X1 U12408 ( .A1(n10432), .A2(n13607), .ZN(n10433) );
  NAND2_X1 U12409 ( .A1(n10817), .A2(n10433), .ZN(n10936) );
  OR2_X1 U12410 ( .A1(n15990), .A2(n15691), .ZN(n16467) );
  INV_X1 U12411 ( .A(n16467), .ZN(n13663) );
  NAND2_X1 U12412 ( .A1(n16468), .A2(n13663), .ZN(n10435) );
  NAND2_X1 U12413 ( .A1(n13667), .A2(n16466), .ZN(n10434) );
  NAND2_X1 U12414 ( .A1(n10435), .A2(n10434), .ZN(n10436) );
  NAND2_X1 U12415 ( .A1(n10436), .A2(n13575), .ZN(n10944) );
  OAI21_X1 U12416 ( .B1(n13575), .B2(n10436), .A(n10944), .ZN(n10438) );
  OAI22_X1 U12417 ( .A1(n13667), .A2(n15951), .B1(n13655), .B2(n15953), .ZN(
        n10437) );
  AOI21_X1 U12418 ( .B1(n10438), .B2(n16561), .A(n10437), .ZN(n10439) );
  OAI21_X1 U12419 ( .B1(n10888), .B2(n15993), .A(n10439), .ZN(n10883) );
  AOI211_X1 U12420 ( .C1(n16660), .C2(n10441), .A(n10440), .B(n10883), .ZN(
        n16518) );
  AND3_X1 U12421 ( .A1(n10873), .A2(n10876), .A3(n10874), .ZN(n11139) );
  NOR2_X1 U12422 ( .A1(n11137), .A2(n13804), .ZN(n10442) );
  NAND2_X1 U12423 ( .A1(n16732), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n10443) );
  OAI21_X1 U12424 ( .B1(n16518), .B2(n16732), .A(n10443), .ZN(P1_U3530) );
  INV_X1 U12425 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n10451) );
  INV_X1 U12426 ( .A(n10444), .ZN(n10447) );
  INV_X1 U12427 ( .A(n10445), .ZN(n10446) );
  MUX2_X1 U12428 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(P1_DATAO_REG_14__SCAN_IN), 
        .S(n7416), .Z(n10619) );
  XNOR2_X1 U12429 ( .A(n10618), .B(n10619), .ZN(n12318) );
  INV_X1 U12430 ( .A(n12318), .ZN(n10456) );
  NAND2_X1 U12431 ( .A1(n10630), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10450) );
  XNOR2_X1 U12432 ( .A(n10450), .B(P2_IR_REG_14__SCAN_IN), .ZN(n12057) );
  INV_X1 U12433 ( .A(n12057), .ZN(n11456) );
  OAI222_X1 U12434 ( .A1(n15545), .A2(n10451), .B1(n15540), .B2(n10456), .C1(
        P2_U3088), .C2(n11456), .ZN(P2_U3313) );
  INV_X1 U12435 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n10452) );
  NAND2_X1 U12436 ( .A1(n10453), .A2(n10452), .ZN(n10454) );
  NAND2_X1 U12437 ( .A1(n10454), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10455) );
  XNOR2_X1 U12438 ( .A(n10455), .B(P1_IR_REG_14__SCAN_IN), .ZN(n12319) );
  INV_X1 U12439 ( .A(n12319), .ZN(n11894) );
  OAI222_X1 U12440 ( .A1(n16139), .A2(n10457), .B1(n11886), .B2(n10456), .C1(
        P1_U3086), .C2(n11894), .ZN(P1_U3341) );
  INV_X1 U12441 ( .A(P3_DATAO_REG_9__SCAN_IN), .ZN(n14459) );
  NAND2_X1 U12442 ( .A1(n12287), .A2(n11041), .ZN(n10458) );
  OAI21_X1 U12443 ( .B1(P3_U3897), .B2(n14459), .A(n10458), .ZN(P3_U3500) );
  INV_X1 U12444 ( .A(P3_DATAO_REG_11__SCAN_IN), .ZN(n14768) );
  NAND2_X1 U12445 ( .A1(n14380), .A2(n11041), .ZN(n10459) );
  OAI21_X1 U12446 ( .B1(n11041), .B2(n14768), .A(n10459), .ZN(P3_U3502) );
  OAI22_X1 U12447 ( .A1(n13309), .A2(n10460), .B1(n15043), .B2(n13024), .ZN(
        n10527) );
  XNOR2_X1 U12448 ( .A(n13021), .B(n15042), .ZN(n13310) );
  INV_X1 U12449 ( .A(n13310), .ZN(n10528) );
  NAND2_X1 U12450 ( .A1(n10527), .A2(n10528), .ZN(n10526) );
  NAND2_X1 U12451 ( .A1(n10547), .A2(n8321), .ZN(n10461) );
  NAND2_X1 U12452 ( .A1(n10526), .A2(n10461), .ZN(n10536) );
  NAND2_X1 U12453 ( .A1(n10536), .A2(n13311), .ZN(n10535) );
  NAND2_X1 U12454 ( .A1(n8111), .A2(n10581), .ZN(n10462) );
  NAND2_X1 U12455 ( .A1(n10535), .A2(n10462), .ZN(n10520) );
  NAND2_X1 U12456 ( .A1(n10703), .A2(n12053), .ZN(n10466) );
  OR2_X1 U12457 ( .A1(n9783), .A2(n10464), .ZN(n10465) );
  OAI211_X1 U12458 ( .C1(n11062), .C2(n15069), .A(n10466), .B(n10465), .ZN(
        n13048) );
  NAND2_X1 U12459 ( .A1(n10485), .A2(n11284), .ZN(n10467) );
  NAND2_X1 U12460 ( .A1(n10732), .A2(n12053), .ZN(n10469) );
  AOI22_X1 U12461 ( .A1(n12597), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n12596), 
        .B2(n15083), .ZN(n10468) );
  NAND2_X1 U12462 ( .A1(n9788), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n10478) );
  NAND2_X1 U12463 ( .A1(n9789), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n10477) );
  AND2_X1 U12464 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n10471) );
  NAND2_X1 U12465 ( .A1(n10471), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n10489) );
  INV_X1 U12466 ( .A(n10471), .ZN(n10473) );
  INV_X1 U12467 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n10472) );
  NAND2_X1 U12468 ( .A1(n10473), .A2(n10472), .ZN(n10474) );
  AND2_X1 U12469 ( .A1(n10489), .A2(n10474), .ZN(n11651) );
  NAND2_X1 U12470 ( .A1(n9786), .A2(n11651), .ZN(n10476) );
  NAND2_X1 U12471 ( .A1(n9790), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n10475) );
  NAND4_X1 U12472 ( .A1(n10478), .A2(n10477), .A3(n10476), .A4(n10475), .ZN(
        n15039) );
  XNOR2_X1 U12473 ( .A(n13054), .B(n15039), .ZN(n13314) );
  XNOR2_X1 U12474 ( .A(n11236), .B(n13314), .ZN(n11650) );
  INV_X1 U12475 ( .A(n15043), .ZN(n10987) );
  NAND2_X1 U12476 ( .A1(n10987), .A2(n13024), .ZN(n10479) );
  NAND2_X1 U12477 ( .A1(n10546), .A2(n10479), .ZN(n10529) );
  NAND2_X1 U12478 ( .A1(n10529), .A2(n13310), .ZN(n10481) );
  NAND2_X1 U12479 ( .A1(n10547), .A2(n13021), .ZN(n10480) );
  NAND2_X1 U12480 ( .A1(n10481), .A2(n10480), .ZN(n10540) );
  NAND2_X1 U12481 ( .A1(n8111), .A2(n13035), .ZN(n10482) );
  NAND2_X1 U12482 ( .A1(n10483), .A2(n10482), .ZN(n10523) );
  INV_X1 U12483 ( .A(n13312), .ZN(n10484) );
  NAND2_X1 U12484 ( .A1(n10485), .A2(n13048), .ZN(n10486) );
  XNOR2_X1 U12485 ( .A(n11249), .B(n13314), .ZN(n10497) );
  NAND2_X1 U12486 ( .A1(n15040), .A2(n15341), .ZN(n10496) );
  NAND2_X1 U12487 ( .A1(n10847), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n10494) );
  NAND2_X1 U12488 ( .A1(n9790), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n10493) );
  INV_X1 U12489 ( .A(n10489), .ZN(n10487) );
  NAND2_X1 U12490 ( .A1(n10487), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n10666) );
  INV_X1 U12491 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n10488) );
  NAND2_X1 U12492 ( .A1(n10489), .A2(n10488), .ZN(n10490) );
  AND2_X1 U12493 ( .A1(n10666), .A2(n10490), .ZN(n10662) );
  NAND2_X1 U12494 ( .A1(n9786), .A2(n10662), .ZN(n10492) );
  NAND2_X1 U12495 ( .A1(n9789), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n10491) );
  NAND4_X1 U12496 ( .A1(n10494), .A2(n10493), .A3(n10492), .A4(n10491), .ZN(
        n15038) );
  NAND2_X1 U12497 ( .A1(n15038), .A2(n15343), .ZN(n10495) );
  NAND2_X1 U12498 ( .A1(n10496), .A2(n10495), .ZN(n11043) );
  AOI21_X1 U12499 ( .B1(n10497), .B2(n15346), .A(n11043), .ZN(n11659) );
  AOI21_X1 U12500 ( .B1(n10522), .B2(n13054), .A(n14937), .ZN(n10498) );
  NAND2_X1 U12501 ( .A1(n10498), .A2(n11274), .ZN(n11655) );
  OAI211_X1 U12502 ( .C1(n11650), .C2(n16738), .A(n11659), .B(n11655), .ZN(
        n10599) );
  INV_X1 U12503 ( .A(n13054), .ZN(n11250) );
  OAI22_X1 U12504 ( .A1(n15464), .A2(n11250), .B1(n16747), .B2(n10087), .ZN(
        n10499) );
  AOI21_X1 U12505 ( .B1(n10599), .B2(n16747), .A(n10499), .ZN(n10500) );
  INV_X1 U12506 ( .A(n10500), .ZN(P2_U3504) );
  INV_X1 U12507 ( .A(n10501), .ZN(n10502) );
  OAI222_X1 U12508 ( .A1(P3_U3151), .A2(n14137), .B1(n14920), .B2(n14492), 
        .C1(n14918), .C2(n10502), .ZN(P3_U3277) );
  INV_X1 U12509 ( .A(P3_DATAO_REG_10__SCAN_IN), .ZN(n10504) );
  NAND2_X1 U12510 ( .A1(n13406), .A2(n11041), .ZN(n10503) );
  OAI21_X1 U12511 ( .B1(n11041), .B2(n10504), .A(n10503), .ZN(P3_U3501) );
  INV_X1 U12512 ( .A(P3_DATAO_REG_12__SCAN_IN), .ZN(n14763) );
  NAND2_X1 U12513 ( .A1(n10505), .A2(n11041), .ZN(n10506) );
  OAI21_X1 U12514 ( .B1(n11041), .B2(n14763), .A(n10506), .ZN(P3_U3503) );
  INV_X1 U12515 ( .A(P3_DATAO_REG_5__SCAN_IN), .ZN(n14578) );
  NAND2_X1 U12516 ( .A1(n12250), .A2(n11041), .ZN(n10507) );
  OAI21_X1 U12517 ( .B1(P3_U3897), .B2(n14578), .A(n10507), .ZN(P3_U3496) );
  INV_X1 U12518 ( .A(P3_DATAO_REG_14__SCAN_IN), .ZN(n14762) );
  NAND2_X1 U12519 ( .A1(n14347), .A2(n11041), .ZN(n10508) );
  OAI21_X1 U12520 ( .B1(n11041), .B2(n14762), .A(n10508), .ZN(P3_U3505) );
  INV_X1 U12521 ( .A(P3_DATAO_REG_13__SCAN_IN), .ZN(n14630) );
  NAND2_X1 U12522 ( .A1(n14379), .A2(n11041), .ZN(n10509) );
  OAI21_X1 U12523 ( .B1(n11041), .B2(n14630), .A(n10509), .ZN(P3_U3504) );
  INV_X1 U12524 ( .A(P3_DATAO_REG_15__SCAN_IN), .ZN(n14629) );
  NAND2_X1 U12525 ( .A1(n14363), .A2(n11041), .ZN(n10510) );
  OAI21_X1 U12526 ( .B1(n11041), .B2(n14629), .A(n10510), .ZN(P3_U3506) );
  INV_X1 U12527 ( .A(P3_DATAO_REG_17__SCAN_IN), .ZN(n14754) );
  NAND2_X1 U12528 ( .A1(n14328), .A2(n11041), .ZN(n10511) );
  OAI21_X1 U12529 ( .B1(n11041), .B2(n14754), .A(n10511), .ZN(P3_U3508) );
  INV_X1 U12530 ( .A(P3_DATAO_REG_16__SCAN_IN), .ZN(n14565) );
  NAND2_X1 U12531 ( .A1(n14348), .A2(n11041), .ZN(n10512) );
  OAI21_X1 U12532 ( .B1(n11041), .B2(n14565), .A(n10512), .ZN(P3_U3507) );
  INV_X1 U12533 ( .A(P3_DATAO_REG_20__SCAN_IN), .ZN(n14751) );
  NAND2_X1 U12534 ( .A1(n8153), .A2(n11041), .ZN(n10513) );
  OAI21_X1 U12535 ( .B1(P3_U3897), .B2(n14751), .A(n10513), .ZN(P3_U3511) );
  INV_X1 U12536 ( .A(P3_DATAO_REG_6__SCAN_IN), .ZN(n10515) );
  NAND2_X1 U12537 ( .A1(n13384), .A2(n11041), .ZN(n10514) );
  OAI21_X1 U12538 ( .B1(P3_U3897), .B2(n10515), .A(n10514), .ZN(P3_U3497) );
  INV_X1 U12539 ( .A(P3_DATAO_REG_8__SCAN_IN), .ZN(n14461) );
  NAND2_X1 U12540 ( .A1(n13396), .A2(n11041), .ZN(n10516) );
  OAI21_X1 U12541 ( .B1(P3_U3897), .B2(n14461), .A(n10516), .ZN(P3_U3499) );
  INV_X1 U12542 ( .A(P3_DATAO_REG_2__SCAN_IN), .ZN(n14778) );
  NAND2_X1 U12543 ( .A1(n10517), .A2(n11041), .ZN(n10518) );
  OAI21_X1 U12544 ( .B1(P3_U3897), .B2(n14778), .A(n10518), .ZN(P3_U3493) );
  OAI21_X1 U12545 ( .B1(n10520), .B2(n13312), .A(n10519), .ZN(n11281) );
  OR2_X1 U12546 ( .A1(n10537), .A2(n11284), .ZN(n10521) );
  AND3_X1 U12547 ( .A1(n10522), .A2(n14960), .A3(n10521), .ZN(n11286) );
  XNOR2_X1 U12548 ( .A(n10523), .B(n13312), .ZN(n10524) );
  AOI22_X1 U12549 ( .A1(n15341), .A2(n15041), .B1(n15039), .B2(n15343), .ZN(
        n11175) );
  OAI21_X1 U12550 ( .B1(n10524), .B2(n15308), .A(n11175), .ZN(n11287) );
  AOI211_X1 U12551 ( .C1(n16641), .C2(n11281), .A(n11286), .B(n11287), .ZN(
        n10592) );
  INV_X1 U12552 ( .A(n15464), .ZN(n15457) );
  AOI22_X1 U12553 ( .A1(n15457), .A2(n13048), .B1(n16746), .B2(
        P2_REG1_REG_4__SCAN_IN), .ZN(n10525) );
  OAI21_X1 U12554 ( .B1(n10592), .B2(n16746), .A(n10525), .ZN(P2_U3503) );
  OAI21_X1 U12555 ( .B1(n10527), .B2(n10528), .A(n10526), .ZN(n11675) );
  OAI211_X1 U12556 ( .C1(n7627), .C2(n8321), .A(n14960), .B(n10538), .ZN(
        n11678) );
  INV_X1 U12557 ( .A(n11678), .ZN(n10533) );
  XNOR2_X1 U12558 ( .A(n10529), .B(n10528), .ZN(n10532) );
  NAND2_X1 U12559 ( .A1(n15043), .A2(n15341), .ZN(n10531) );
  NAND2_X1 U12560 ( .A1(n15041), .A2(n15343), .ZN(n10530) );
  AND2_X1 U12561 ( .A1(n10531), .A2(n10530), .ZN(n11126) );
  OAI21_X1 U12562 ( .B1(n10532), .B2(n15308), .A(n11126), .ZN(n11674) );
  AOI211_X1 U12563 ( .C1(n16641), .C2(n11675), .A(n10533), .B(n11674), .ZN(
        n10588) );
  AOI22_X1 U12564 ( .A1(n15457), .A2(n13021), .B1(n16746), .B2(
        P2_REG1_REG_2__SCAN_IN), .ZN(n10534) );
  OAI21_X1 U12565 ( .B1(n10588), .B2(n16746), .A(n10534), .ZN(P2_U3501) );
  OAI21_X1 U12566 ( .B1(n10536), .B2(n13311), .A(n10535), .ZN(n11669) );
  AOI211_X1 U12567 ( .C1(n13035), .C2(n10538), .A(n14937), .B(n10537), .ZN(
        n11668) );
  XNOR2_X1 U12568 ( .A(n10540), .B(n10539), .ZN(n10542) );
  AOI21_X1 U12569 ( .B1(n10542), .B2(n15346), .A(n10541), .ZN(n11672) );
  INV_X1 U12570 ( .A(n11672), .ZN(n10543) );
  AOI211_X1 U12571 ( .C1(n16641), .C2(n11669), .A(n11668), .B(n10543), .ZN(
        n10584) );
  AOI22_X1 U12572 ( .A1(n15457), .A2(n13035), .B1(n16746), .B2(
        P2_REG1_REG_3__SCAN_IN), .ZN(n10544) );
  OAI21_X1 U12573 ( .B1(n10584), .B2(n16746), .A(n10544), .ZN(P2_U3502) );
  XNOR2_X1 U12574 ( .A(n13309), .B(n10545), .ZN(n11301) );
  INV_X1 U12575 ( .A(n11301), .ZN(n10550) );
  AOI211_X1 U12576 ( .C1(n10984), .C2(n13024), .A(n14937), .B(n7627), .ZN(
        n11296) );
  OAI21_X1 U12577 ( .B1(n13015), .B2(n13309), .A(n10546), .ZN(n10548) );
  INV_X1 U12578 ( .A(n13013), .ZN(n10981) );
  OAI22_X1 U12579 ( .A1(n10981), .A2(n15289), .B1(n10547), .B2(n15287), .ZN(
        n10564) );
  AOI21_X1 U12580 ( .B1(n10548), .B2(n15346), .A(n10564), .ZN(n11297) );
  INV_X1 U12581 ( .A(n11297), .ZN(n10549) );
  AOI211_X1 U12582 ( .C1(n10550), .C2(n16641), .A(n11296), .B(n10549), .ZN(
        n10596) );
  AOI22_X1 U12583 ( .A1(n15457), .A2(n13024), .B1(n16746), .B2(
        P2_REG1_REG_1__SCAN_IN), .ZN(n10551) );
  OAI21_X1 U12584 ( .B1(n10596), .B2(n16746), .A(n10551), .ZN(P2_U3500) );
  INV_X1 U12585 ( .A(P3_DATAO_REG_23__SCAN_IN), .ZN(n10553) );
  NAND2_X1 U12586 ( .A1(n14232), .A2(n11041), .ZN(n10552) );
  OAI21_X1 U12587 ( .B1(n11041), .B2(n10553), .A(n10552), .ZN(P3_U3514) );
  INV_X1 U12588 ( .A(P3_DATAO_REG_4__SCAN_IN), .ZN(n14775) );
  NAND2_X1 U12589 ( .A1(n10554), .A2(n11041), .ZN(n10555) );
  OAI21_X1 U12590 ( .B1(P3_U3897), .B2(n14775), .A(n10555), .ZN(P3_U3495) );
  INV_X1 U12591 ( .A(P3_DATAO_REG_7__SCAN_IN), .ZN(n14766) );
  NAND2_X1 U12592 ( .A1(n13391), .A2(n11041), .ZN(n10556) );
  OAI21_X1 U12593 ( .B1(n11041), .B2(n14766), .A(n10556), .ZN(P3_U3498) );
  INV_X1 U12594 ( .A(P3_DATAO_REG_19__SCAN_IN), .ZN(n14562) );
  NAND2_X1 U12595 ( .A1(n14298), .A2(n11041), .ZN(n10557) );
  OAI21_X1 U12596 ( .B1(n11041), .B2(n14562), .A(n10557), .ZN(P3_U3510) );
  INV_X1 U12597 ( .A(P3_DATAO_REG_3__SCAN_IN), .ZN(n14777) );
  NAND2_X1 U12598 ( .A1(n16496), .A2(n11041), .ZN(n10558) );
  OAI21_X1 U12599 ( .B1(P3_U3897), .B2(n14777), .A(n10558), .ZN(P3_U3494) );
  INV_X1 U12600 ( .A(P3_DATAO_REG_0__SCAN_IN), .ZN(n14584) );
  NAND2_X1 U12601 ( .A1(n11534), .A2(n11041), .ZN(n10559) );
  OAI21_X1 U12602 ( .B1(P3_U3897), .B2(n14584), .A(n10559), .ZN(P3_U3491) );
  INV_X1 U12603 ( .A(P3_DATAO_REG_18__SCAN_IN), .ZN(n14563) );
  NAND2_X1 U12604 ( .A1(n13859), .A2(n11041), .ZN(n10560) );
  OAI21_X1 U12605 ( .B1(n11041), .B2(n14563), .A(n10560), .ZN(P3_U3509) );
  INV_X1 U12606 ( .A(P3_DATAO_REG_21__SCAN_IN), .ZN(n14752) );
  NAND2_X1 U12607 ( .A1(n14233), .A2(n11041), .ZN(n10561) );
  OAI21_X1 U12608 ( .B1(n11041), .B2(n14752), .A(n10561), .ZN(P3_U3512) );
  INV_X1 U12609 ( .A(P3_DATAO_REG_1__SCAN_IN), .ZN(n14780) );
  NAND2_X1 U12610 ( .A1(n16497), .A2(n11041), .ZN(n10562) );
  OAI21_X1 U12611 ( .B1(n11041), .B2(n14780), .A(n10562), .ZN(P3_U3492) );
  OR2_X1 U12612 ( .A1(n10563), .A2(P2_U3088), .ZN(n11123) );
  AOI22_X1 U12613 ( .A1(n14991), .A2(n10564), .B1(P2_REG3_REG_1__SCAN_IN), 
        .B2(n11123), .ZN(n10569) );
  OAI21_X1 U12614 ( .B1(n10566), .B2(n10565), .A(n11128), .ZN(n10567) );
  NAND2_X1 U12615 ( .A1(n15000), .A2(n10567), .ZN(n10568) );
  OAI211_X1 U12616 ( .C1(n14994), .C2(n11294), .A(n10569), .B(n10568), .ZN(
        P2_U3194) );
  INV_X2 U12617 ( .A(n12862), .ZN(n12945) );
  NAND2_X1 U12618 ( .A1(n12945), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n10577) );
  INV_X1 U12619 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n15821) );
  OR2_X1 U12620 ( .A1(n12929), .A2(n15821), .ZN(n10576) );
  AND2_X1 U12621 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n10696) );
  NAND2_X1 U12622 ( .A1(n10696), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n10821) );
  NAND2_X1 U12623 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_REG3_REG_7__SCAN_IN), 
        .ZN(n10570) );
  NOR2_X1 U12624 ( .A1(n10821), .A2(n10570), .ZN(n10822) );
  NAND2_X1 U12625 ( .A1(n10822), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n11550) );
  INV_X1 U12626 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n11564) );
  NOR2_X1 U12627 ( .A1(n11565), .A2(n11564), .ZN(n11563) );
  AND2_X1 U12628 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_REG3_REG_12__SCAN_IN), 
        .ZN(n10571) );
  NAND2_X1 U12629 ( .A1(n11859), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n12025) );
  INV_X1 U12630 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n12024) );
  INV_X1 U12631 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n12307) );
  INV_X1 U12632 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n12350) );
  NAND2_X1 U12633 ( .A1(n12349), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n12745) );
  INV_X1 U12634 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n12744) );
  INV_X1 U12635 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n12763) );
  NAND2_X1 U12636 ( .A1(n12799), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n12800) );
  NAND2_X1 U12637 ( .A1(n12817), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n12816) );
  NAND2_X1 U12638 ( .A1(n12837), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n12836) );
  INV_X1 U12639 ( .A(n12836), .ZN(n12860) );
  NAND2_X1 U12640 ( .A1(n12860), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n12859) );
  INV_X1 U12641 ( .A(n12859), .ZN(n12880) );
  NAND2_X1 U12642 ( .A1(P1_REG3_REG_25__SCAN_IN), .A2(n12880), .ZN(n12897) );
  INV_X1 U12643 ( .A(n12897), .ZN(n10572) );
  NAND2_X1 U12644 ( .A1(n10572), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n12931) );
  INV_X1 U12645 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n15552) );
  XNOR2_X1 U12646 ( .A(n12931), .B(n15552), .ZN(n15820) );
  OR2_X1 U12647 ( .A1(n12946), .A2(n15820), .ZN(n10575) );
  INV_X1 U12648 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n10573) );
  OR2_X1 U12649 ( .A1(n7418), .A2(n10573), .ZN(n10574) );
  NAND2_X1 U12650 ( .A1(P1_U4016), .A2(n15838), .ZN(n10578) );
  OAI21_X1 U12651 ( .B1(P1_U4016), .B2(n10579), .A(n10578), .ZN(P1_U3587) );
  INV_X1 U12652 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10580) );
  OAI22_X1 U12653 ( .A1(n15517), .A2(n10581), .B1(n16751), .B2(n10580), .ZN(
        n10582) );
  INV_X1 U12654 ( .A(n10582), .ZN(n10583) );
  OAI21_X1 U12655 ( .B1(n10584), .B2(n16748), .A(n10583), .ZN(P2_U3439) );
  INV_X1 U12656 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10585) );
  OAI22_X1 U12657 ( .A1(n15517), .A2(n8321), .B1(n16751), .B2(n10585), .ZN(
        n10586) );
  INV_X1 U12658 ( .A(n10586), .ZN(n10587) );
  OAI21_X1 U12659 ( .B1(n10588), .B2(n16748), .A(n10587), .ZN(P2_U3436) );
  INV_X1 U12660 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10589) );
  OAI22_X1 U12661 ( .A1(n15517), .A2(n11284), .B1(n16751), .B2(n10589), .ZN(
        n10590) );
  INV_X1 U12662 ( .A(n10590), .ZN(n10591) );
  OAI21_X1 U12663 ( .B1(n10592), .B2(n16748), .A(n10591), .ZN(P2_U3442) );
  INV_X1 U12664 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10593) );
  OAI22_X1 U12665 ( .A1(n15517), .A2(n11294), .B1(n16751), .B2(n10593), .ZN(
        n10594) );
  INV_X1 U12666 ( .A(n10594), .ZN(n10595) );
  OAI21_X1 U12667 ( .B1(n10596), .B2(n16748), .A(n10595), .ZN(P2_U3433) );
  INV_X1 U12668 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10597) );
  OAI22_X1 U12669 ( .A1(n15517), .A2(n11250), .B1(n16751), .B2(n10597), .ZN(
        n10598) );
  AOI21_X1 U12670 ( .B1(n10599), .B2(n16751), .A(n10598), .ZN(n10600) );
  INV_X1 U12671 ( .A(n10600), .ZN(P2_U3445) );
  INV_X1 U12672 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n10601) );
  MUX2_X1 U12673 ( .A(n10601), .B(P1_REG1_REG_10__SCAN_IN), .S(n11559), .Z(
        n10604) );
  OAI21_X1 U12674 ( .B1(P1_REG1_REG_9__SCAN_IN), .B2(n11546), .A(n10602), .ZN(
        n10603) );
  NOR2_X1 U12675 ( .A1(n10603), .A2(n10604), .ZN(n10755) );
  AOI211_X1 U12676 ( .C1(n10604), .C2(n10603), .A(n15710), .B(n10755), .ZN(
        n10616) );
  NOR2_X1 U12677 ( .A1(n10605), .A2(n10304), .ZN(n10607) );
  INV_X1 U12678 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n11562) );
  MUX2_X1 U12679 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n11562), .S(n11559), .Z(
        n10606) );
  OAI21_X1 U12680 ( .B1(n10608), .B2(n10607), .A(n10606), .ZN(n10753) );
  INV_X1 U12681 ( .A(n10753), .ZN(n10610) );
  NOR3_X1 U12682 ( .A1(n10608), .A2(n10607), .A3(n10606), .ZN(n10609) );
  NOR3_X1 U12683 ( .A1(n10610), .A2(n10609), .A3(n15728), .ZN(n10615) );
  NAND2_X1 U12684 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_U3086), .ZN(n12124)
         );
  INV_X1 U12685 ( .A(n12124), .ZN(n10611) );
  AOI21_X1 U12686 ( .B1(n16246), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n10611), 
        .ZN(n10612) );
  OAI21_X1 U12687 ( .B1(n15727), .B2(n10613), .A(n10612), .ZN(n10614) );
  OR3_X1 U12688 ( .A1(n10616), .A2(n10615), .A3(n10614), .ZN(P1_U3253) );
  INV_X1 U12689 ( .A(n10617), .ZN(n10620) );
  MUX2_X1 U12690 ( .A(n10644), .B(n10632), .S(n7416), .Z(n10622) );
  NAND2_X1 U12691 ( .A1(n10622), .A2(n10621), .ZN(n10869) );
  INV_X1 U12692 ( .A(n10622), .ZN(n10623) );
  NAND2_X1 U12693 ( .A1(n10623), .A2(SI_15_), .ZN(n10624) );
  NAND2_X1 U12694 ( .A1(n10869), .A2(n10624), .ZN(n10627) );
  NAND2_X1 U12695 ( .A1(n10628), .A2(n10627), .ZN(n10629) );
  NAND2_X1 U12696 ( .A1(n10870), .A2(n10629), .ZN(n12338) );
  INV_X1 U12697 ( .A(n12338), .ZN(n10643) );
  OAI21_X1 U12698 ( .B1(n10630), .B2(P2_IR_REG_14__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n10631) );
  XNOR2_X1 U12699 ( .A(n10631), .B(P2_IR_REG_15__SCAN_IN), .ZN(n12054) );
  INV_X1 U12700 ( .A(n12054), .ZN(n11457) );
  OAI222_X1 U12701 ( .A1(n15545), .A2(n10632), .B1(n15540), .B2(n10643), .C1(
        P2_U3088), .C2(n11457), .ZN(P2_U3312) );
  NOR2_X1 U12702 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), 
        .ZN(n10634) );
  AND4_X1 U12703 ( .A1(n10635), .A2(n10634), .A3(n10633), .A4(n14617), .ZN(
        n10636) );
  NAND2_X1 U12704 ( .A1(n10637), .A2(n10636), .ZN(n10639) );
  NAND2_X1 U12705 ( .A1(n10639), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10638) );
  MUX2_X1 U12706 ( .A(P1_IR_REG_31__SCAN_IN), .B(n10638), .S(
        P1_IR_REG_15__SCAN_IN), .Z(n10642) );
  INV_X1 U12707 ( .A(n10639), .ZN(n10641) );
  INV_X1 U12708 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n10640) );
  NAND2_X1 U12709 ( .A1(n10641), .A2(n10640), .ZN(n11166) );
  OAI222_X1 U12710 ( .A1(n16139), .A2(n10644), .B1(n11886), .B2(n10643), .C1(
        P1_U3086), .C2(n11898), .ZN(P1_U3340) );
  XNOR2_X1 U12711 ( .A(n14936), .B(n13048), .ZN(n11046) );
  NAND2_X1 U12712 ( .A1(n15040), .A2(n14937), .ZN(n10648) );
  XNOR2_X1 U12713 ( .A(n11046), .B(n10648), .ZN(n11179) );
  AND2_X1 U12714 ( .A1(n11179), .A2(n10645), .ZN(n10646) );
  INV_X1 U12715 ( .A(n11046), .ZN(n10649) );
  NAND2_X1 U12716 ( .A1(n10649), .A2(n10648), .ZN(n10650) );
  NAND2_X1 U12717 ( .A1(n15039), .A2(n14937), .ZN(n10652) );
  INV_X1 U12718 ( .A(n10651), .ZN(n10653) );
  NAND2_X1 U12719 ( .A1(n10811), .A2(n12053), .ZN(n10655) );
  AOI22_X1 U12720 ( .A1(n12597), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n12596), 
        .B2(n15105), .ZN(n10654) );
  XNOR2_X1 U12721 ( .A(n16586), .B(n14936), .ZN(n10656) );
  AND2_X1 U12722 ( .A1(n15038), .A2(n14937), .ZN(n10657) );
  NAND2_X1 U12723 ( .A1(n10656), .A2(n10657), .ZN(n11056) );
  INV_X1 U12724 ( .A(n10656), .ZN(n11181) );
  INV_X1 U12725 ( .A(n10657), .ZN(n10658) );
  NAND2_X1 U12726 ( .A1(n11181), .A2(n10658), .ZN(n10659) );
  NAND2_X1 U12727 ( .A1(n11056), .A2(n10659), .ZN(n10660) );
  INV_X1 U12728 ( .A(n11058), .ZN(n11183) );
  AOI211_X1 U12729 ( .C1(n10661), .C2(n10660), .A(n15021), .B(n11183), .ZN(
        n10674) );
  INV_X1 U12730 ( .A(n10662), .ZN(n11275) );
  NAND2_X1 U12731 ( .A1(n15024), .A2(n16586), .ZN(n10663) );
  NAND2_X1 U12732 ( .A1(P2_U3088), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n15103) );
  OAI211_X1 U12733 ( .C1(n15003), .C2(n11275), .A(n10663), .B(n15103), .ZN(
        n10673) );
  NAND2_X1 U12734 ( .A1(n10847), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n10671) );
  NAND2_X1 U12735 ( .A1(n9790), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n10670) );
  INV_X1 U12736 ( .A(n10666), .ZN(n10664) );
  NAND2_X1 U12737 ( .A1(n10664), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n11070) );
  INV_X1 U12738 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n10665) );
  NAND2_X1 U12739 ( .A1(n10666), .A2(n10665), .ZN(n10667) );
  AND2_X1 U12740 ( .A1(n11070), .A2(n10667), .ZN(n11259) );
  NAND2_X1 U12741 ( .A1(n9786), .A2(n11259), .ZN(n10669) );
  NAND2_X1 U12742 ( .A1(n9789), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n10668) );
  NAND4_X1 U12743 ( .A1(n10671), .A2(n10670), .A3(n10669), .A4(n10668), .ZN(
        n15037) );
  NAND2_X1 U12744 ( .A1(n14991), .A2(n15343), .ZN(n14972) );
  NAND2_X1 U12745 ( .A1(n14991), .A2(n15341), .ZN(n12994) );
  INV_X1 U12746 ( .A(n15039), .ZN(n11265) );
  OAI22_X1 U12747 ( .A1(n13064), .A2(n14972), .B1(n12994), .B2(n11265), .ZN(
        n10672) );
  OR3_X1 U12748 ( .A1(n10674), .A2(n10673), .A3(n10672), .ZN(P2_U3211) );
  INV_X1 U12749 ( .A(n10675), .ZN(n10676) );
  OAI222_X1 U12750 ( .A1(P3_U3151), .A2(n14132), .B1(n14918), .B2(n10676), 
        .C1(n14666), .C2(n14920), .ZN(P3_U3276) );
  INV_X1 U12751 ( .A(n10677), .ZN(n10680) );
  INV_X1 U12752 ( .A(n10678), .ZN(n10679) );
  NAND2_X1 U12753 ( .A1(n7413), .A2(n15690), .ZN(n10689) );
  OR2_X1 U12754 ( .A1(n10702), .A2(n10683), .ZN(n10686) );
  OR2_X1 U12755 ( .A1(n10704), .A2(n10684), .ZN(n10685) );
  NAND2_X1 U12756 ( .A1(n7412), .A2(n16527), .ZN(n10688) );
  NAND2_X1 U12757 ( .A1(n10689), .A2(n10688), .ZN(n10690) );
  XNOR2_X1 U12758 ( .A(n10690), .B(n12720), .ZN(n10691) );
  INV_X1 U12759 ( .A(n16527), .ZN(n13653) );
  OAI22_X1 U12760 ( .A1(n12846), .A2(n13655), .B1(n13653), .B2(n10271), .ZN(
        n10692) );
  XNOR2_X1 U12761 ( .A(n10691), .B(n10692), .ZN(n16529) );
  INV_X1 U12762 ( .A(n10691), .ZN(n10693) );
  OR2_X1 U12763 ( .A1(n12929), .A2(n10695), .ZN(n10700) );
  INV_X1 U12764 ( .A(n10696), .ZN(n10716) );
  OAI21_X1 U12765 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(n10716), .ZN(n10951) );
  OR2_X1 U12766 ( .A1(n12946), .A2(n10951), .ZN(n10699) );
  INV_X1 U12767 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10697) );
  OR2_X1 U12768 ( .A1(n10418), .A2(n10697), .ZN(n10698) );
  NAND2_X1 U12769 ( .A1(n11544), .A2(n10703), .ZN(n10707) );
  OR2_X1 U12770 ( .A1(n10704), .A2(n10705), .ZN(n10706) );
  OAI211_X1 U12771 ( .C1(n12814), .C2(n10708), .A(n10707), .B(n10706), .ZN(
        n16554) );
  AOI22_X1 U12772 ( .A1(n12921), .A2(n15689), .B1(n7413), .B2(n16554), .ZN(
        n10709) );
  NOR2_X1 U12773 ( .A1(n10729), .A2(n7631), .ZN(n10711) );
  INV_X1 U12774 ( .A(n15689), .ZN(n13678) );
  OAI22_X1 U12775 ( .A1(n13678), .A2(n10271), .B1(n13677), .B2(n12940), .ZN(
        n10710) );
  XNOR2_X1 U12776 ( .A(n10710), .B(n10817), .ZN(n10730) );
  XNOR2_X1 U12777 ( .A(n10711), .B(n10730), .ZN(n10728) );
  NAND2_X1 U12778 ( .A1(n10713), .A2(n10712), .ZN(n10714) );
  INV_X1 U12779 ( .A(n15638), .ZN(n16530) );
  NAND2_X1 U12780 ( .A1(n13566), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n10721) );
  OR2_X1 U12781 ( .A1(n12862), .A2(n10715), .ZN(n10720) );
  OR2_X1 U12782 ( .A1(n12929), .A2(n10042), .ZN(n10719) );
  INV_X1 U12783 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n10745) );
  NAND2_X1 U12784 ( .A1(n10716), .A2(n10745), .ZN(n10717) );
  NAND2_X1 U12785 ( .A1(n10821), .A2(n10717), .ZN(n11442) );
  OR2_X1 U12786 ( .A1(n12946), .A2(n11442), .ZN(n10718) );
  OR2_X1 U12787 ( .A1(n13684), .A2(n15953), .ZN(n10723) );
  NAND2_X1 U12788 ( .A1(n15690), .A2(n15971), .ZN(n10722) );
  NAND2_X1 U12789 ( .A1(n10723), .A2(n10722), .ZN(n16553) );
  NAND2_X1 U12790 ( .A1(n16530), .A2(n16553), .ZN(n10724) );
  OAI211_X1 U12791 ( .C1(n16535), .C2(n10951), .A(n10725), .B(n10724), .ZN(
        n10726) );
  AOI21_X1 U12792 ( .B1(n15671), .B2(n16554), .A(n10726), .ZN(n10727) );
  OAI21_X1 U12793 ( .B1(n10728), .B2(n15673), .A(n10727), .ZN(P1_U3230) );
  NAND2_X1 U12794 ( .A1(n10732), .A2(n11544), .ZN(n10733) );
  OAI22_X1 U12795 ( .A1(n13684), .A2(n10271), .B1(n16572), .B2(n12940), .ZN(
        n10734) );
  XNOR2_X1 U12796 ( .A(n10734), .B(n10817), .ZN(n10736) );
  OAI22_X1 U12797 ( .A1(n12846), .A2(n13684), .B1(n16572), .B2(n10271), .ZN(
        n10735) );
  NOR2_X1 U12798 ( .A1(n10736), .A2(n10735), .ZN(n10808) );
  INV_X1 U12799 ( .A(n10808), .ZN(n10737) );
  NAND2_X1 U12800 ( .A1(n10736), .A2(n10735), .ZN(n10809) );
  NAND2_X1 U12801 ( .A1(n10737), .A2(n10809), .ZN(n10738) );
  XNOR2_X1 U12802 ( .A(n10810), .B(n10738), .ZN(n10749) );
  NAND2_X1 U12803 ( .A1(n12945), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n10744) );
  OR2_X1 U12804 ( .A1(n12929), .A2(n10739), .ZN(n10743) );
  INV_X1 U12805 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n10820) );
  XNOR2_X1 U12806 ( .A(n10821), .B(n10820), .ZN(n11427) );
  OR2_X1 U12807 ( .A1(n12946), .A2(n11427), .ZN(n10742) );
  INV_X1 U12808 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10740) );
  OR2_X1 U12809 ( .A1(n10418), .A2(n10740), .ZN(n10741) );
  NAND4_X1 U12810 ( .A1(n10744), .A2(n10743), .A3(n10742), .A4(n10741), .ZN(
        n15687) );
  INV_X1 U12811 ( .A(n15687), .ZN(n10819) );
  OAI22_X1 U12812 ( .A1(n15648), .A2(n10819), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10745), .ZN(n10747) );
  OAI22_X1 U12813 ( .A1(n15653), .A2(n16572), .B1(n16535), .B2(n11442), .ZN(
        n10746) );
  AOI211_X1 U12814 ( .C1(n15659), .C2(n15689), .A(n10747), .B(n10746), .ZN(
        n10748) );
  OAI21_X1 U12815 ( .B1(n10749), .B2(n15673), .A(n10748), .ZN(P1_U3227) );
  NAND2_X1 U12816 ( .A1(n11559), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n10752) );
  INV_X1 U12817 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n10750) );
  MUX2_X1 U12818 ( .A(n10750), .B(P1_REG2_REG_11__SCAN_IN), .S(n11852), .Z(
        n10751) );
  AOI21_X1 U12819 ( .B1(n10753), .B2(n10752), .A(n10751), .ZN(n10970) );
  NAND3_X1 U12820 ( .A1(n10753), .A2(n10752), .A3(n10751), .ZN(n10754) );
  NAND2_X1 U12821 ( .A1(n10754), .A2(n16263), .ZN(n10763) );
  INV_X1 U12822 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n11575) );
  MUX2_X1 U12823 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n11575), .S(n11852), .Z(
        n10756) );
  NAND2_X1 U12824 ( .A1(n10757), .A2(n10756), .ZN(n16256) );
  OAI21_X1 U12825 ( .B1(n10757), .B2(n10756), .A(n16256), .ZN(n10758) );
  NAND2_X1 U12826 ( .A1(n10758), .A2(n16259), .ZN(n10762) );
  NAND2_X1 U12827 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n11990)
         );
  INV_X1 U12828 ( .A(n11990), .ZN(n10760) );
  NOR2_X1 U12829 ( .A1(n15727), .A2(n10965), .ZN(n10759) );
  AOI211_X1 U12830 ( .C1(n16246), .C2(P1_ADDR_REG_11__SCAN_IN), .A(n10760), 
        .B(n10759), .ZN(n10761) );
  OAI211_X1 U12831 ( .C1(n10970), .C2(n10763), .A(n10762), .B(n10761), .ZN(
        P1_U3254) );
  INV_X1 U12832 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n10764) );
  MUX2_X1 U12833 ( .A(n10764), .B(P2_REG2_REG_13__SCAN_IN), .S(n11784), .Z(
        n10771) );
  NAND2_X1 U12834 ( .A1(n11091), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n10765) );
  AND2_X1 U12835 ( .A1(n10766), .A2(n10765), .ZN(n16186) );
  INV_X1 U12836 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n10767) );
  MUX2_X1 U12837 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n10767), .S(n16184), .Z(
        n16187) );
  NAND2_X1 U12838 ( .A1(n16186), .A2(n16187), .ZN(n16185) );
  OR2_X1 U12839 ( .A1(n16184), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n10768) );
  NAND2_X1 U12840 ( .A1(n16185), .A2(n10768), .ZN(n10769) );
  NAND2_X1 U12841 ( .A1(n10769), .A2(n10776), .ZN(n10770) );
  OAI21_X1 U12842 ( .B1(n10769), .B2(n10776), .A(n10770), .ZN(n16226) );
  OR2_X1 U12843 ( .A1(n16226), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n16228) );
  NAND2_X1 U12844 ( .A1(n16228), .A2(n10770), .ZN(n10772) );
  AOI21_X1 U12845 ( .B1(n10771), .B2(n10772), .A(n16220), .ZN(n10773) );
  NAND2_X1 U12846 ( .A1(n10773), .A2(n10799), .ZN(n10781) );
  INV_X1 U12847 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n16708) );
  AOI21_X1 U12848 ( .B1(n11091), .B2(P2_REG1_REG_10__SCAN_IN), .A(n10774), 
        .ZN(n16192) );
  INV_X1 U12849 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n10775) );
  MUX2_X1 U12850 ( .A(n10775), .B(P2_REG1_REG_11__SCAN_IN), .S(n16184), .Z(
        n16191) );
  NOR2_X1 U12851 ( .A1(n16192), .A2(n16191), .ZN(n16189) );
  AOI21_X1 U12852 ( .B1(n16184), .B2(P2_REG1_REG_11__SCAN_IN), .A(n16189), 
        .ZN(n16225) );
  MUX2_X1 U12853 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n16708), .S(n16232), .Z(
        n16224) );
  AND2_X1 U12854 ( .A1(n16225), .A2(n16224), .ZN(n16222) );
  AOI21_X1 U12855 ( .B1(n16708), .B2(n10776), .A(n16222), .ZN(n10779) );
  INV_X1 U12856 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n10777) );
  MUX2_X1 U12857 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n10777), .S(n11784), .Z(
        n10778) );
  NAND2_X1 U12858 ( .A1(n10779), .A2(n10778), .ZN(n10794) );
  OAI211_X1 U12859 ( .C1(n10779), .C2(n10778), .A(n16233), .B(n10794), .ZN(
        n10780) );
  NAND2_X1 U12860 ( .A1(n10781), .A2(n10780), .ZN(n10783) );
  NAND2_X1 U12861 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_U3088), .ZN(n11809)
         );
  INV_X1 U12862 ( .A(n11809), .ZN(n10782) );
  AOI211_X1 U12863 ( .C1(n10096), .C2(P2_ADDR_REG_13__SCAN_IN), .A(n10783), 
        .B(n10782), .ZN(n10784) );
  OAI21_X1 U12864 ( .B1(n10800), .B2(n16214), .A(n10784), .ZN(P2_U3227) );
  INV_X1 U12865 ( .A(n10785), .ZN(n10786) );
  OAI222_X1 U12866 ( .A1(P3_U3151), .A2(n10787), .B1(n14918), .B2(n10786), 
        .C1(n14664), .C2(n14920), .ZN(P3_U3275) );
  INV_X1 U12867 ( .A(P3_DATAO_REG_25__SCAN_IN), .ZN(n14468) );
  NAND2_X1 U12868 ( .A1(n8350), .A2(n11041), .ZN(n10788) );
  OAI21_X1 U12869 ( .B1(n11041), .B2(n14468), .A(n10788), .ZN(P3_U3516) );
  INV_X1 U12870 ( .A(n16450), .ZN(n11637) );
  AND2_X1 U12871 ( .A1(n11534), .A2(n11637), .ZN(n13362) );
  INV_X1 U12872 ( .A(n13362), .ZN(n13358) );
  AND2_X1 U12873 ( .A1(n13358), .A2(n11400), .ZN(n16447) );
  NAND2_X1 U12874 ( .A1(n10789), .A2(n16711), .ZN(n10790) );
  OAI22_X1 U12875 ( .A1(n16447), .A2(n10790), .B1(n11333), .B2(n14314), .ZN(
        n11635) );
  NOR2_X1 U12876 ( .A1(n16718), .A2(n9597), .ZN(n10791) );
  AOI21_X1 U12877 ( .B1(n16718), .B2(n11635), .A(n10791), .ZN(n10792) );
  OAI21_X1 U12878 ( .B1(n11637), .B2(n14455), .A(n10792), .ZN(P3_U3459) );
  INV_X1 U12879 ( .A(n10096), .ZN(n16237) );
  INV_X1 U12880 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n10793) );
  NAND2_X1 U12881 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3088), .ZN(n12683)
         );
  OAI21_X1 U12882 ( .B1(n16237), .B2(n10793), .A(n12683), .ZN(n10806) );
  OAI21_X1 U12883 ( .B1(n10777), .B2(n10800), .A(n10794), .ZN(n10796) );
  INV_X1 U12884 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n11807) );
  MUX2_X1 U12885 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n11807), .S(n12057), .Z(
        n10795) );
  NAND2_X1 U12886 ( .A1(n10796), .A2(n10795), .ZN(n11455) );
  OAI211_X1 U12887 ( .C1(n10796), .C2(n10795), .A(n11455), .B(n16233), .ZN(
        n10804) );
  INV_X1 U12888 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n10797) );
  MUX2_X1 U12889 ( .A(n10797), .B(P2_REG2_REG_14__SCAN_IN), .S(n12057), .Z(
        n10798) );
  INV_X1 U12890 ( .A(n10798), .ZN(n10802) );
  OAI21_X1 U12891 ( .B1(n10764), .B2(n10800), .A(n10799), .ZN(n10801) );
  NAND2_X1 U12892 ( .A1(n10802), .A2(n10801), .ZN(n11459) );
  OAI211_X1 U12893 ( .C1(n10802), .C2(n10801), .A(n16229), .B(n11459), .ZN(
        n10803) );
  NAND2_X1 U12894 ( .A1(n10804), .A2(n10803), .ZN(n10805) );
  AOI211_X1 U12895 ( .C1(n16231), .C2(n12057), .A(n10806), .B(n10805), .ZN(
        n10807) );
  INV_X1 U12896 ( .A(n10807), .ZN(P2_U3228) );
  NAND2_X1 U12897 ( .A1(n10811), .A2(n11544), .ZN(n10814) );
  AOI22_X1 U12898 ( .A1(n12760), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n12759), 
        .B2(n10812), .ZN(n10813) );
  NAND2_X1 U12899 ( .A1(n10814), .A2(n10813), .ZN(n13689) );
  NAND2_X1 U12900 ( .A1(n7412), .A2(n13689), .ZN(n10816) );
  NAND2_X1 U12901 ( .A1(n7413), .A2(n15687), .ZN(n10815) );
  NAND2_X1 U12902 ( .A1(n10816), .A2(n10815), .ZN(n10818) );
  XNOR2_X1 U12903 ( .A(n10818), .B(n12720), .ZN(n11018) );
  INV_X1 U12904 ( .A(n13689), .ZN(n11341) );
  OAI22_X1 U12905 ( .A1(n12846), .A2(n10819), .B1(n11341), .B2(n10271), .ZN(
        n11020) );
  XNOR2_X1 U12906 ( .A(n11018), .B(n11020), .ZN(n11021) );
  XNOR2_X1 U12907 ( .A(n11022), .B(n11021), .ZN(n10833) );
  NAND2_X1 U12908 ( .A1(n13566), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n10828) );
  OR2_X1 U12909 ( .A1(n12929), .A2(n10158), .ZN(n10827) );
  OAI21_X1 U12910 ( .B1(n10821), .B2(n10820), .A(n11035), .ZN(n10823) );
  INV_X1 U12911 ( .A(n10822), .ZN(n11029) );
  NAND2_X1 U12912 ( .A1(n10823), .A2(n11029), .ZN(n11352) );
  OR2_X1 U12913 ( .A1(n12946), .A2(n11352), .ZN(n10826) );
  OR2_X1 U12914 ( .A1(n12862), .A2(n10824), .ZN(n10825) );
  NAND4_X1 U12915 ( .A1(n10828), .A2(n10827), .A3(n10826), .A4(n10825), .ZN(
        n15686) );
  OAI21_X1 U12916 ( .B1(n15648), .B2(n8629), .A(n10829), .ZN(n10831) );
  OAI22_X1 U12917 ( .A1(n15653), .A2(n11341), .B1(n11427), .B2(n16535), .ZN(
        n10830) );
  AOI211_X1 U12918 ( .C1(n15659), .C2(n15688), .A(n10831), .B(n10830), .ZN(
        n10832) );
  OAI21_X1 U12919 ( .B1(n10833), .B2(n15673), .A(n10832), .ZN(P1_U3239) );
  OAI222_X1 U12920 ( .A1(P3_U3151), .A2(n10835), .B1(n14918), .B2(n10834), 
        .C1(n14662), .C2(n14920), .ZN(P3_U3274) );
  INV_X1 U12921 ( .A(P3_DATAO_REG_26__SCAN_IN), .ZN(n14465) );
  NAND2_X1 U12922 ( .A1(n14176), .A2(n11041), .ZN(n10836) );
  OAI21_X1 U12923 ( .B1(n11041), .B2(n14465), .A(n10836), .ZN(P3_U3517) );
  INV_X1 U12924 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n11069) );
  INV_X1 U12925 ( .A(n11095), .ZN(n10837) );
  NAND2_X1 U12926 ( .A1(n10837), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n11111) );
  INV_X1 U12927 ( .A(n11111), .ZN(n10838) );
  NAND2_X1 U12928 ( .A1(n10838), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n11369) );
  INV_X1 U12929 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n11368) );
  INV_X1 U12930 ( .A(n11768), .ZN(n10839) );
  NAND2_X1 U12931 ( .A1(n10839), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n11803) );
  INV_X1 U12932 ( .A(n11803), .ZN(n10840) );
  NAND2_X1 U12933 ( .A1(n10840), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n12067) );
  INV_X1 U12934 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n12066) );
  INV_X1 U12935 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n12178) );
  INV_X1 U12936 ( .A(n12962), .ZN(n10843) );
  NAND2_X1 U12937 ( .A1(n10843), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n12985) );
  INV_X1 U12938 ( .A(n12985), .ZN(n10844) );
  NAND2_X1 U12939 ( .A1(n10844), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n12996) );
  INV_X1 U12940 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n12995) );
  INV_X1 U12941 ( .A(n13167), .ZN(n10845) );
  NAND2_X1 U12942 ( .A1(n10845), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n13180) );
  INV_X1 U12943 ( .A(n13180), .ZN(n10846) );
  NAND2_X1 U12944 ( .A1(n10846), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n13201) );
  INV_X1 U12945 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n13200) );
  XNOR2_X1 U12946 ( .A(n13260), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n15199) );
  NAND2_X1 U12947 ( .A1(n15199), .A2(n9786), .ZN(n10852) );
  INV_X1 U12948 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n15398) );
  NAND2_X1 U12949 ( .A1(n9789), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n10849) );
  NAND2_X1 U12950 ( .A1(n10847), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n10848) );
  OAI211_X1 U12951 ( .C1(n13265), .C2(n15398), .A(n10849), .B(n10848), .ZN(
        n10850) );
  INV_X1 U12952 ( .A(n10850), .ZN(n10851) );
  NAND2_X1 U12953 ( .A1(n10852), .A2(n10851), .ZN(n15017) );
  NAND2_X1 U12954 ( .A1(n15017), .A2(P2_U3947), .ZN(n10853) );
  OAI21_X1 U12955 ( .B1(n16123), .B2(P2_U3947), .A(n10853), .ZN(P2_U3558) );
  INV_X1 U12956 ( .A(n16429), .ZN(n11199) );
  OAI21_X1 U12957 ( .B1(n10854), .B2(P3_REG1_REG_3__SCAN_IN), .A(n11198), .ZN(
        n10859) );
  AOI21_X1 U12958 ( .B1(n11820), .B2(n10855), .A(n11193), .ZN(n10857) );
  NOR2_X1 U12959 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n14474), .ZN(n11424) );
  AOI21_X1 U12960 ( .B1(n16150), .B2(P3_ADDR_REG_3__SCAN_IN), .A(n11424), .ZN(
        n10856) );
  OAI21_X1 U12961 ( .B1(n10857), .B2(n16423), .A(n10856), .ZN(n10858) );
  AOI21_X1 U12962 ( .B1(n11199), .B2(n10859), .A(n10858), .ZN(n10867) );
  INV_X1 U12963 ( .A(n11228), .ZN(n10863) );
  INV_X1 U12964 ( .A(n10860), .ZN(n10862) );
  NOR3_X1 U12965 ( .A1(n10863), .A2(n10862), .A3(n10861), .ZN(n10865) );
  INV_X1 U12966 ( .A(n11207), .ZN(n10864) );
  OAI21_X1 U12967 ( .B1(n10865), .B2(n10864), .A(n14125), .ZN(n10866) );
  OAI211_X1 U12968 ( .C1(n16427), .C2(n10868), .A(n10867), .B(n10866), .ZN(
        P3_U3185) );
  MUX2_X1 U12969 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(P1_DATAO_REG_16__SCAN_IN), 
        .S(n7416), .Z(n11159) );
  INV_X1 U12970 ( .A(n12539), .ZN(n10992) );
  NAND2_X1 U12971 ( .A1(n11166), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10871) );
  XNOR2_X1 U12972 ( .A(n10871), .B(P1_IR_REG_16__SCAN_IN), .ZN(n12540) );
  AOI22_X1 U12973 ( .A1(n12540), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n11168), .ZN(n10872) );
  OAI21_X1 U12974 ( .B1(n10992), .B2(n11886), .A(n10872), .ZN(P1_U3339) );
  INV_X1 U12975 ( .A(n10873), .ZN(n10875) );
  NAND4_X1 U12976 ( .A1(n10875), .A2(n11136), .A3(n10874), .A4(n11137), .ZN(
        n15790) );
  INV_X1 U12977 ( .A(n10876), .ZN(n10877) );
  OR2_X1 U12978 ( .A1(n13660), .A2(n15733), .ZN(n13625) );
  OR2_X1 U12979 ( .A1(n7414), .A2(n13625), .ZN(n15826) );
  OAI22_X1 U12980 ( .A1(n16631), .A2(n10881), .B1(n10880), .B2(n16622), .ZN(
        n10882) );
  AOI21_X1 U12981 ( .B1(n16628), .B2(n8046), .A(n10882), .ZN(n10887) );
  INV_X1 U12982 ( .A(n10883), .ZN(n10884) );
  MUX2_X1 U12983 ( .A(n10885), .B(n10884), .S(n16625), .Z(n10886) );
  OAI211_X1 U12984 ( .C1(n10888), .C2(n15826), .A(n10887), .B(n10886), .ZN(
        P1_U3291) );
  INV_X1 U12985 ( .A(n16423), .ZN(n14120) );
  OAI21_X1 U12986 ( .B1(n7635), .B2(P3_REG2_REG_1__SCAN_IN), .A(n10889), .ZN(
        n10891) );
  OAI22_X1 U12987 ( .A1(n16438), .A2(n16272), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n11531), .ZN(n10890) );
  AOI21_X1 U12988 ( .B1(n14120), .B2(n10891), .A(n10890), .ZN(n10897) );
  XNOR2_X1 U12989 ( .A(n10892), .B(P3_REG1_REG_1__SCAN_IN), .ZN(n10895) );
  OAI21_X1 U12990 ( .B1(n11313), .B2(n10893), .A(n11226), .ZN(n10894) );
  AOI22_X1 U12991 ( .A1(n11199), .A2(n10895), .B1(n14125), .B2(n10894), .ZN(
        n10896) );
  OAI211_X1 U12992 ( .C1(n10898), .C2(n16427), .A(n10897), .B(n10896), .ZN(
        P3_U3183) );
  INV_X1 U12993 ( .A(n10899), .ZN(n10901) );
  NAND2_X1 U12994 ( .A1(n10901), .A2(n10900), .ZN(n10902) );
  XNOR2_X1 U12995 ( .A(n10903), .B(n10902), .ZN(n10915) );
  AOI21_X1 U12996 ( .B1(n10906), .B2(n10905), .A(n10904), .ZN(n10912) );
  INV_X1 U12997 ( .A(P3_REG3_REG_6__SCAN_IN), .ZN(n14741) );
  NOR2_X1 U12998 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n14741), .ZN(n11683) );
  AOI21_X1 U12999 ( .B1(n7628), .B2(n10908), .A(n10907), .ZN(n10909) );
  NOR2_X1 U13000 ( .A1(n16423), .A2(n10909), .ZN(n10910) );
  AOI211_X1 U13001 ( .C1(n16150), .C2(P3_ADDR_REG_6__SCAN_IN), .A(n11683), .B(
        n10910), .ZN(n10911) );
  OAI21_X1 U13002 ( .B1(n10912), .B2(n16429), .A(n10911), .ZN(n10913) );
  AOI21_X1 U13003 ( .B1(n7816), .B2(n14146), .A(n10913), .ZN(n10914) );
  OAI21_X1 U13004 ( .B1(n16418), .B2(n10915), .A(n10914), .ZN(P3_U3188) );
  OAI21_X1 U13005 ( .B1(n10918), .B2(n10917), .A(n10916), .ZN(n10930) );
  AOI21_X1 U13006 ( .B1(n9024), .B2(n10920), .A(n10919), .ZN(n10928) );
  INV_X1 U13007 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n14716) );
  NOR2_X1 U13008 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n14716), .ZN(n11664) );
  AOI21_X1 U13009 ( .B1(n11928), .B2(n10922), .A(n10921), .ZN(n10923) );
  NOR2_X1 U13010 ( .A1(n16423), .A2(n10923), .ZN(n10924) );
  AOI211_X1 U13011 ( .C1(n16150), .C2(P3_ADDR_REG_5__SCAN_IN), .A(n11664), .B(
        n10924), .ZN(n10927) );
  NAND2_X1 U13012 ( .A1(n14146), .A2(n10925), .ZN(n10926) );
  OAI211_X1 U13013 ( .C1(n10928), .C2(n16429), .A(n10927), .B(n10926), .ZN(
        n10929) );
  AOI21_X1 U13014 ( .B1(n14125), .B2(n10930), .A(n10929), .ZN(n10931) );
  INV_X1 U13015 ( .A(n10931), .ZN(P3_U3187) );
  NAND2_X1 U13016 ( .A1(n8047), .A2(n10934), .ZN(n10935) );
  XNOR2_X1 U13017 ( .A(n10948), .B(n13671), .ZN(n16541) );
  NAND2_X1 U13018 ( .A1(n15689), .A2(n16462), .ZN(n10938) );
  NAND2_X1 U13019 ( .A1(n16463), .A2(n15971), .ZN(n10937) );
  NAND2_X1 U13020 ( .A1(n10938), .A2(n10937), .ZN(n16537) );
  MUX2_X1 U13021 ( .A(n16537), .B(P1_REG2_REG_3__SCAN_IN), .S(n7414), .Z(
        n10943) );
  NAND2_X1 U13022 ( .A1(n10940), .A2(n16527), .ZN(n10939) );
  NAND2_X1 U13023 ( .A1(n10939), .A2(n16079), .ZN(n10941) );
  OR2_X1 U13024 ( .A1(n10941), .A2(n10950), .ZN(n16538) );
  OAI22_X1 U13025 ( .A1(n16631), .A2(n16538), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(n16622), .ZN(n10942) );
  AOI211_X1 U13026 ( .C1(n16628), .C2(n16527), .A(n10943), .B(n10942), .ZN(
        n10946) );
  NAND2_X1 U13027 ( .A1(n10944), .A2(n13665), .ZN(n10954) );
  XNOR2_X1 U13028 ( .A(n10954), .B(n13671), .ZN(n16543) );
  NAND2_X1 U13029 ( .A1(n15855), .A2(n16543), .ZN(n10945) );
  OAI211_X1 U13030 ( .C1(n16541), .C2(n15983), .A(n10946), .B(n10945), .ZN(
        P1_U3290) );
  INV_X1 U13031 ( .A(n13671), .ZN(n10947) );
  NAND2_X1 U13032 ( .A1(n13655), .A2(n13653), .ZN(n10949) );
  INV_X1 U13033 ( .A(n13675), .ZN(n13576) );
  XNOR2_X1 U13034 ( .A(n11142), .B(n13576), .ZN(n16552) );
  INV_X1 U13035 ( .A(n16552), .ZN(n10959) );
  MUX2_X1 U13036 ( .A(n16553), .B(P1_REG2_REG_4__SCAN_IN), .S(n7414), .Z(
        n10953) );
  OAI211_X1 U13037 ( .C1(n10950), .C2(n13677), .A(n16079), .B(n11439), .ZN(
        n16556) );
  OAI22_X1 U13038 ( .A1(n16631), .A2(n16556), .B1(n10951), .B2(n16622), .ZN(
        n10952) );
  AOI211_X1 U13039 ( .C1(n16628), .C2(n16554), .A(n10953), .B(n10952), .ZN(
        n10958) );
  NAND2_X1 U13040 ( .A1(n10954), .A2(n13671), .ZN(n10956) );
  NAND2_X1 U13041 ( .A1(n13655), .A2(n16527), .ZN(n10955) );
  NAND2_X1 U13042 ( .A1(n10956), .A2(n10955), .ZN(n11147) );
  XNOR2_X1 U13043 ( .A(n11147), .B(n13675), .ZN(n16560) );
  NAND2_X1 U13044 ( .A1(n16560), .A2(n15855), .ZN(n10957) );
  OAI211_X1 U13045 ( .C1(n10959), .C2(n15983), .A(n10958), .B(n10957), .ZN(
        P1_U3289) );
  INV_X1 U13046 ( .A(n10960), .ZN(n10962) );
  OAI22_X1 U13047 ( .A1(n13557), .A2(P3_U3151), .B1(SI_22_), .B2(n14920), .ZN(
        n10961) );
  AOI21_X1 U13048 ( .B1(n10962), .B2(n14901), .A(n10961), .ZN(P3_U3273) );
  INV_X1 U13049 ( .A(P3_DATAO_REG_29__SCAN_IN), .ZN(n14729) );
  NAND2_X1 U13050 ( .A1(n10963), .A2(n11041), .ZN(n10964) );
  OAI21_X1 U13051 ( .B1(P3_U3897), .B2(n14729), .A(n10964), .ZN(P3_U3520) );
  INV_X1 U13052 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n10966) );
  NAND2_X1 U13053 ( .A1(n10965), .A2(n11575), .ZN(n16255) );
  MUX2_X1 U13054 ( .A(n10966), .B(P1_REG1_REG_12__SCAN_IN), .S(n16262), .Z(
        n16254) );
  AOI21_X1 U13055 ( .B1(n16256), .B2(n16255), .A(n16254), .ZN(n16253) );
  AOI21_X1 U13056 ( .B1(n10967), .B2(n10966), .A(n16253), .ZN(n10969) );
  INV_X1 U13057 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n16733) );
  MUX2_X1 U13058 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n16733), .S(n12007), .Z(
        n10968) );
  NAND2_X1 U13059 ( .A1(n10969), .A2(n10968), .ZN(n11467) );
  OAI211_X1 U13060 ( .C1(n10969), .C2(n10968), .A(n11467), .B(n16259), .ZN(
        n10979) );
  AOI21_X1 U13061 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n11852), .A(n10970), 
        .ZN(n16251) );
  INV_X1 U13062 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n10971) );
  MUX2_X1 U13063 ( .A(P1_REG2_REG_12__SCAN_IN), .B(n10971), .S(n16262), .Z(
        n16252) );
  NAND2_X1 U13064 ( .A1(n16251), .A2(n16252), .ZN(n16250) );
  OAI21_X1 U13065 ( .B1(n16262), .B2(P1_REG2_REG_12__SCAN_IN), .A(n16250), 
        .ZN(n10973) );
  INV_X1 U13066 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n12023) );
  MUX2_X1 U13067 ( .A(n12023), .B(P1_REG2_REG_13__SCAN_IN), .S(n12007), .Z(
        n10972) );
  NOR2_X1 U13068 ( .A1(n10973), .A2(n10972), .ZN(n11479) );
  AOI211_X1 U13069 ( .C1(n10973), .C2(n10972), .A(n15728), .B(n11479), .ZN(
        n10977) );
  INV_X1 U13070 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n12010) );
  NOR2_X1 U13071 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n12010), .ZN(n10974) );
  AOI21_X1 U13072 ( .B1(n16246), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n10974), 
        .ZN(n10975) );
  OAI21_X1 U13073 ( .B1(n15727), .B2(n11473), .A(n10975), .ZN(n10976) );
  NOR2_X1 U13074 ( .A1(n10977), .A2(n10976), .ZN(n10978) );
  NAND2_X1 U13075 ( .A1(n10979), .A2(n10978), .ZN(P1_U3256) );
  INV_X1 U13076 ( .A(P3_DATAO_REG_27__SCAN_IN), .ZN(n14726) );
  NAND2_X1 U13077 ( .A1(n13821), .A2(n11041), .ZN(n10980) );
  OAI21_X1 U13078 ( .B1(n11041), .B2(n14726), .A(n10980), .ZN(P3_U3518) );
  INV_X1 U13079 ( .A(n14961), .ZN(n15011) );
  OAI22_X1 U13080 ( .A1(n15011), .A2(n10981), .B1(n13012), .B2(n15021), .ZN(
        n10983) );
  NAND2_X1 U13081 ( .A1(n10983), .A2(n10982), .ZN(n10986) );
  AOI22_X1 U13082 ( .A1(n15024), .A2(n10984), .B1(P2_REG3_REG_0__SCAN_IN), 
        .B2(n11123), .ZN(n10985) );
  OAI211_X1 U13083 ( .C1(n10987), .C2(n14972), .A(n10986), .B(n10985), .ZN(
        P2_U3204) );
  NAND2_X1 U13084 ( .A1(n10989), .A2(P3_DATAO_REG_30__SCAN_IN), .ZN(n10988) );
  OAI21_X1 U13085 ( .B1(n13507), .B2(n10989), .A(n10988), .ZN(P3_U3521) );
  INV_X1 U13086 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n10993) );
  NAND2_X1 U13087 ( .A1(n10990), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10991) );
  XNOR2_X1 U13088 ( .A(n10991), .B(P2_IR_REG_16__SCAN_IN), .ZN(n12170) );
  INV_X1 U13089 ( .A(n12170), .ZN(n16199) );
  OAI222_X1 U13090 ( .A1(n15545), .A2(n10993), .B1(n15540), .B2(n10992), .C1(
        n16199), .C2(P2_U3088), .ZN(P2_U3311) );
  INV_X1 U13091 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n14728) );
  INV_X1 U13092 ( .A(P3_REG0_REG_31__SCAN_IN), .ZN(n10999) );
  NAND2_X1 U13093 ( .A1(n8980), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n10997) );
  INV_X1 U13094 ( .A(P3_REG1_REG_31__SCAN_IN), .ZN(n10994) );
  OR2_X1 U13095 ( .A1(n10995), .A2(n10994), .ZN(n10996) );
  OAI211_X1 U13096 ( .C1(n10999), .C2(n10998), .A(n10997), .B(n10996), .ZN(
        n11000) );
  INV_X1 U13097 ( .A(n11000), .ZN(n11001) );
  NAND2_X1 U13098 ( .A1(n11002), .A2(n11001), .ZN(n14151) );
  NAND2_X1 U13099 ( .A1(n14151), .A2(n11041), .ZN(n11003) );
  OAI21_X1 U13100 ( .B1(P3_U3897), .B2(n14728), .A(n11003), .ZN(P3_U3522) );
  INV_X1 U13101 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n11017) );
  INV_X1 U13102 ( .A(n11004), .ZN(n11005) );
  NOR2_X1 U13103 ( .A1(n11008), .A2(n11005), .ZN(n11007) );
  MUX2_X1 U13104 ( .A(n11008), .B(n11007), .S(n11006), .Z(n11009) );
  NOR2_X1 U13105 ( .A1(n16711), .A2(n13550), .ZN(n11011) );
  INV_X1 U13106 ( .A(n13550), .ZN(n16510) );
  OR2_X1 U13107 ( .A1(n16711), .A2(n16510), .ZN(n11013) );
  INV_X1 U13108 ( .A(n14384), .ZN(n14354) );
  AOI22_X1 U13109 ( .A1(n14354), .A2(n16450), .B1(P3_REG3_REG_0__SCAN_IN), 
        .B2(n14369), .ZN(n11016) );
  NAND2_X1 U13110 ( .A1(n11635), .A2(n14352), .ZN(n11015) );
  OAI211_X1 U13111 ( .C1(n11017), .C2(n14352), .A(n11016), .B(n11015), .ZN(
        P3_U3233) );
  INV_X1 U13112 ( .A(n11018), .ZN(n11019) );
  NAND2_X1 U13113 ( .A1(n11053), .A2(n11544), .ZN(n11025) );
  AOI22_X1 U13114 ( .A1(n12760), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n12759), 
        .B2(n11023), .ZN(n11024) );
  NAND2_X1 U13115 ( .A1(n11025), .A2(n11024), .ZN(n16607) );
  AOI22_X1 U13116 ( .A1(n16607), .A2(n7412), .B1(n7413), .B2(n15686), .ZN(
        n11026) );
  XNOR2_X1 U13117 ( .A(n11026), .B(n10817), .ZN(n11688) );
  AOI22_X1 U13118 ( .A1(n12921), .A2(n15686), .B1(n16607), .B2(n7413), .ZN(
        n11689) );
  XNOR2_X1 U13119 ( .A(n11688), .B(n11689), .ZN(n11690) );
  XNOR2_X1 U13120 ( .A(n11691), .B(n11690), .ZN(n11039) );
  NAND2_X1 U13121 ( .A1(n13566), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n11034) );
  OR2_X1 U13122 ( .A1(n12929), .A2(n16624), .ZN(n11033) );
  OR2_X1 U13123 ( .A1(n12862), .A2(n11027), .ZN(n11032) );
  INV_X1 U13124 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n11028) );
  NAND2_X1 U13125 ( .A1(n11029), .A2(n11028), .ZN(n11030) );
  NAND2_X1 U13126 ( .A1(n11550), .A2(n11030), .ZN(n16623) );
  OR2_X1 U13127 ( .A1(n12946), .A2(n16623), .ZN(n11031) );
  NAND4_X1 U13128 ( .A1(n11034), .A2(n11033), .A3(n11032), .A4(n11031), .ZN(
        n15685) );
  AOI22_X1 U13129 ( .A1(n15971), .A2(n15687), .B1(n15685), .B2(n16462), .ZN(
        n16603) );
  OAI22_X1 U13130 ( .A1(n15638), .A2(n16603), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n11035), .ZN(n11037) );
  NOR2_X1 U13131 ( .A1(n16535), .A2(n11352), .ZN(n11036) );
  AOI211_X1 U13132 ( .C1(n15671), .C2(n16607), .A(n11037), .B(n11036), .ZN(
        n11038) );
  OAI21_X1 U13133 ( .B1(n11039), .B2(n15673), .A(n11038), .ZN(P1_U3213) );
  INV_X1 U13134 ( .A(P3_DATAO_REG_28__SCAN_IN), .ZN(n14732) );
  INV_X1 U13135 ( .A(n11040), .ZN(n14175) );
  NAND2_X1 U13136 ( .A1(n14175), .A2(n11041), .ZN(n11042) );
  OAI21_X1 U13137 ( .B1(n11041), .B2(n14732), .A(n11042), .ZN(P3_U3519) );
  INV_X1 U13138 ( .A(n11043), .ZN(n11045) );
  AOI22_X1 U13139 ( .A1(n15018), .A2(n11651), .B1(P2_REG3_REG_5__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11044) );
  OAI21_X1 U13140 ( .B1(n15020), .B2(n11045), .A(n11044), .ZN(n11050) );
  AOI22_X1 U13141 ( .A1(n14961), .A2(n15040), .B1(n15000), .B2(n11046), .ZN(
        n11048) );
  NOR3_X1 U13142 ( .A1(n11048), .A2(n8496), .A3(n11047), .ZN(n11049) );
  AOI211_X1 U13143 ( .C1(n13054), .C2(n15024), .A(n11050), .B(n11049), .ZN(
        n11051) );
  OAI21_X1 U13144 ( .B1(n11052), .B2(n15021), .A(n11051), .ZN(P2_U3199) );
  NAND2_X1 U13145 ( .A1(n11053), .A2(n12053), .ZN(n11055) );
  AOI22_X1 U13146 ( .A1(n12597), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n12596), 
        .B2(n16172), .ZN(n11054) );
  NAND2_X1 U13147 ( .A1(n11055), .A2(n11054), .ZN(n13062) );
  XNOR2_X1 U13148 ( .A(n13062), .B(n14936), .ZN(n12675) );
  NAND2_X1 U13149 ( .A1(n15037), .A2(n14937), .ZN(n11059) );
  XNOR2_X1 U13150 ( .A(n12675), .B(n11059), .ZN(n11189) );
  AND2_X1 U13151 ( .A1(n11189), .A2(n11056), .ZN(n11057) );
  NAND2_X1 U13152 ( .A1(n11058), .A2(n11057), .ZN(n11184) );
  INV_X1 U13153 ( .A(n12675), .ZN(n11060) );
  NAND2_X1 U13154 ( .A1(n11060), .A2(n11059), .ZN(n11061) );
  NAND2_X1 U13155 ( .A1(n11539), .A2(n12053), .ZN(n11067) );
  OAI22_X1 U13156 ( .A1(n9783), .A2(n11064), .B1(n11063), .B2(n11062), .ZN(
        n11065) );
  INV_X1 U13157 ( .A(n11065), .ZN(n11066) );
  NAND2_X1 U13158 ( .A1(n11067), .A2(n11066), .ZN(n13071) );
  XNOR2_X1 U13159 ( .A(n13071), .B(n14959), .ZN(n11076) );
  NAND2_X1 U13160 ( .A1(n9788), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n11075) );
  NAND2_X1 U13161 ( .A1(n9790), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n11074) );
  NAND2_X1 U13162 ( .A1(n11070), .A2(n11069), .ZN(n11071) );
  AND2_X1 U13163 ( .A1(n11082), .A2(n11071), .ZN(n12670) );
  NAND2_X1 U13164 ( .A1(n9786), .A2(n12670), .ZN(n11073) );
  NAND2_X1 U13165 ( .A1(n9789), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n11072) );
  NAND4_X1 U13166 ( .A1(n11075), .A2(n11074), .A3(n11073), .A4(n11072), .ZN(
        n15036) );
  NAND2_X1 U13167 ( .A1(n15036), .A2(n14937), .ZN(n11077) );
  XNOR2_X1 U13168 ( .A(n11076), .B(n11077), .ZN(n12676) );
  INV_X1 U13169 ( .A(n11076), .ZN(n12658) );
  NAND2_X1 U13170 ( .A1(n11545), .A2(n12053), .ZN(n11080) );
  AOI22_X1 U13171 ( .A1(n12596), .A2(n11078), .B1(n12597), .B2(
        P1_DATAO_REG_9__SCAN_IN), .ZN(n11079) );
  NAND2_X1 U13172 ( .A1(n11080), .A2(n11079), .ZN(n13077) );
  XNOR2_X1 U13173 ( .A(n13077), .B(n14959), .ZN(n11103) );
  NAND2_X1 U13174 ( .A1(n9788), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n11087) );
  NAND2_X1 U13175 ( .A1(n9790), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n11086) );
  NAND2_X1 U13176 ( .A1(n11082), .A2(n11081), .ZN(n11083) );
  NAND2_X1 U13177 ( .A1(n11095), .A2(n11083), .ZN(n12662) );
  INV_X1 U13178 ( .A(n12662), .ZN(n11395) );
  NAND2_X1 U13179 ( .A1(n9786), .A2(n11395), .ZN(n11085) );
  NAND2_X1 U13180 ( .A1(n9789), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n11084) );
  NAND4_X1 U13181 ( .A1(n11087), .A2(n11086), .A3(n11085), .A4(n11084), .ZN(
        n15035) );
  NAND2_X1 U13182 ( .A1(n15035), .A2(n14937), .ZN(n11088) );
  XNOR2_X1 U13183 ( .A(n11103), .B(n11088), .ZN(n12656) );
  INV_X1 U13184 ( .A(n11103), .ZN(n11089) );
  NAND2_X1 U13185 ( .A1(n11089), .A2(n11088), .ZN(n11090) );
  NAND2_X1 U13186 ( .A1(n11558), .A2(n12053), .ZN(n11093) );
  AOI22_X1 U13187 ( .A1(n11091), .A2(n12596), .B1(n12597), .B2(
        P1_DATAO_REG_10__SCAN_IN), .ZN(n11092) );
  XNOR2_X1 U13188 ( .A(n13083), .B(n14959), .ZN(n11364) );
  NAND2_X1 U13189 ( .A1(n9790), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n11100) );
  NAND2_X1 U13190 ( .A1(n10847), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n11099) );
  INV_X1 U13191 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n11094) );
  NAND2_X1 U13192 ( .A1(n11095), .A2(n11094), .ZN(n11096) );
  AND2_X1 U13193 ( .A1(n11111), .A2(n11096), .ZN(n11599) );
  NAND2_X1 U13194 ( .A1(n9786), .A2(n11599), .ZN(n11098) );
  NAND2_X1 U13195 ( .A1(n9789), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n11097) );
  NAND4_X1 U13196 ( .A1(n11100), .A2(n11099), .A3(n11098), .A4(n11097), .ZN(
        n15034) );
  NAND2_X1 U13197 ( .A1(n15034), .A2(n14937), .ZN(n11358) );
  XNOR2_X1 U13198 ( .A(n11364), .B(n11358), .ZN(n11102) );
  INV_X1 U13199 ( .A(n11361), .ZN(n11367) );
  NAND2_X1 U13200 ( .A1(n11103), .A2(n15000), .ZN(n11105) );
  NAND2_X1 U13201 ( .A1(n14961), .A2(n15035), .ZN(n11104) );
  NAND2_X1 U13202 ( .A1(n11105), .A2(n11104), .ZN(n11106) );
  NAND3_X1 U13203 ( .A1(n11101), .A2(n7920), .A3(n11106), .ZN(n11120) );
  INV_X1 U13204 ( .A(n12994), .ZN(n14974) );
  INV_X1 U13205 ( .A(n11599), .ZN(n11108) );
  OAI21_X1 U13206 ( .B1(n15003), .B2(n11108), .A(n11107), .ZN(n11109) );
  AOI21_X1 U13207 ( .B1(n14974), .B2(n15035), .A(n11109), .ZN(n11119) );
  NAND2_X1 U13208 ( .A1(n13083), .A2(n15024), .ZN(n11118) );
  NAND2_X1 U13209 ( .A1(n9790), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n11116) );
  NAND2_X1 U13210 ( .A1(n10847), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n11115) );
  INV_X1 U13211 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n11110) );
  NAND2_X1 U13212 ( .A1(n11111), .A2(n11110), .ZN(n11112) );
  AND2_X1 U13213 ( .A1(n11369), .A2(n11112), .ZN(n11375) );
  NAND2_X1 U13214 ( .A1(n9786), .A2(n11375), .ZN(n11114) );
  NAND2_X1 U13215 ( .A1(n9789), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n11113) );
  NAND4_X1 U13216 ( .A1(n11116), .A2(n11115), .A3(n11114), .A4(n11113), .ZN(
        n15033) );
  OR2_X1 U13217 ( .A1(n14972), .A2(n13089), .ZN(n11117) );
  NAND4_X1 U13218 ( .A1(n11120), .A2(n11119), .A3(n11118), .A4(n11117), .ZN(
        n11121) );
  AOI21_X1 U13219 ( .B1(n11367), .B2(n15000), .A(n11121), .ZN(n11122) );
  INV_X1 U13220 ( .A(n11122), .ZN(P2_U3189) );
  INV_X1 U13221 ( .A(n11123), .ZN(n11125) );
  INV_X1 U13222 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n11124) );
  OAI22_X1 U13223 ( .A1(n15020), .A2(n11126), .B1(n11125), .B2(n11124), .ZN(
        n11133) );
  AOI22_X1 U13224 ( .A1(n14961), .A2(n15043), .B1(n15000), .B2(n11127), .ZN(
        n11131) );
  INV_X1 U13225 ( .A(n11128), .ZN(n11130) );
  NOR3_X1 U13226 ( .A1(n11131), .A2(n11130), .A3(n11129), .ZN(n11132) );
  AOI211_X1 U13227 ( .C1(n13021), .C2(n15024), .A(n11133), .B(n11132), .ZN(
        n11134) );
  OAI21_X1 U13228 ( .B1(n11135), .B2(n15021), .A(n11134), .ZN(P2_U3209) );
  NOR2_X1 U13229 ( .A1(n15689), .A2(n16554), .ZN(n11141) );
  NAND2_X1 U13230 ( .A1(n15689), .A2(n16554), .ZN(n11140) );
  OAI21_X1 U13231 ( .B1(n11142), .B2(n11141), .A(n11140), .ZN(n11436) );
  INV_X1 U13232 ( .A(n11436), .ZN(n11143) );
  XNOR2_X1 U13233 ( .A(n15688), .B(n13685), .ZN(n13578) );
  INV_X1 U13234 ( .A(n13578), .ZN(n11445) );
  NAND2_X1 U13235 ( .A1(n11143), .A2(n11445), .ZN(n11438) );
  NAND2_X1 U13236 ( .A1(n13684), .A2(n16572), .ZN(n11144) );
  XNOR2_X1 U13237 ( .A(n15687), .B(n13689), .ZN(n13579) );
  INV_X1 U13238 ( .A(n13579), .ZN(n11145) );
  NAND2_X1 U13239 ( .A1(n11345), .A2(n11145), .ZN(n11344) );
  OAI21_X1 U13240 ( .B1(n11345), .B2(n11145), .A(n11344), .ZN(n11434) );
  INV_X1 U13241 ( .A(n11440), .ZN(n11146) );
  OAI211_X1 U13242 ( .C1(n11341), .C2(n11146), .A(n11349), .B(n16079), .ZN(
        n11430) );
  OAI21_X1 U13243 ( .B1(n11341), .B2(n16725), .A(n11430), .ZN(n11153) );
  OR2_X1 U13244 ( .A1(n13684), .A2(n13685), .ZN(n11148) );
  NAND2_X1 U13245 ( .A1(n11149), .A2(n11148), .ZN(n11340) );
  XNOR2_X1 U13246 ( .A(n11340), .B(n13579), .ZN(n11152) );
  NAND2_X1 U13247 ( .A1(n11434), .A2(n16472), .ZN(n11151) );
  AOI22_X1 U13248 ( .A1(n15688), .A2(n15971), .B1(n16462), .B2(n15686), .ZN(
        n11150) );
  OAI211_X1 U13249 ( .C1(n16726), .C2(n11152), .A(n11151), .B(n11150), .ZN(
        n11431) );
  AOI211_X1 U13250 ( .C1(n16660), .C2(n11434), .A(n11153), .B(n11431), .ZN(
        n11155) );
  OR2_X1 U13251 ( .A1(n11155), .A2(n16735), .ZN(n11154) );
  OAI21_X1 U13252 ( .B1(n16737), .B2(n10740), .A(n11154), .ZN(P1_U3477) );
  INV_X1 U13253 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n11157) );
  OR2_X1 U13254 ( .A1(n11155), .A2(n16732), .ZN(n11156) );
  OAI21_X1 U13255 ( .B1(n16734), .B2(n11157), .A(n11156), .ZN(P1_U3534) );
  MUX2_X1 U13256 ( .A(n8040), .B(n11329), .S(n7416), .Z(n11163) );
  NAND2_X1 U13257 ( .A1(n11163), .A2(n11162), .ZN(n11741) );
  INV_X1 U13258 ( .A(n11163), .ZN(n11164) );
  NAND2_X1 U13259 ( .A1(n11164), .A2(SI_17_), .ZN(n11165) );
  NAND2_X1 U13260 ( .A1(n11741), .A2(n11165), .ZN(n11742) );
  INV_X1 U13261 ( .A(n12728), .ZN(n11328) );
  NAND2_X1 U13262 ( .A1(n11744), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n11167) );
  XNOR2_X1 U13263 ( .A(n11167), .B(P1_IR_REG_17__SCAN_IN), .ZN(n15709) );
  AOI22_X1 U13264 ( .A1(n15709), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n11168), .ZN(n11169) );
  OAI21_X1 U13265 ( .B1(n11328), .B2(n11886), .A(n11169), .ZN(P1_U3338) );
  NOR3_X1 U13266 ( .A1(n15011), .A2(n11170), .A3(n8111), .ZN(n11171) );
  AOI21_X1 U13267 ( .B1(n15000), .B2(n11172), .A(n11171), .ZN(n11180) );
  NOR2_X1 U13268 ( .A1(n15021), .A2(n11173), .ZN(n11177) );
  NAND2_X1 U13269 ( .A1(P2_U3088), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n15062) );
  NAND2_X1 U13270 ( .A1(n15018), .A2(n11282), .ZN(n11174) );
  OAI211_X1 U13271 ( .C1(n15020), .C2(n11175), .A(n15062), .B(n11174), .ZN(
        n11176) );
  AOI211_X1 U13272 ( .C1(n13048), .C2(n15024), .A(n11177), .B(n11176), .ZN(
        n11178) );
  OAI21_X1 U13273 ( .B1(n11180), .B2(n11179), .A(n11178), .ZN(P2_U3202) );
  INV_X1 U13274 ( .A(n15038), .ZN(n13058) );
  NOR3_X1 U13275 ( .A1(n15011), .A2(n11181), .A3(n13058), .ZN(n11182) );
  AOI21_X1 U13276 ( .B1(n15014), .B2(n11183), .A(n11182), .ZN(n11190) );
  INV_X1 U13277 ( .A(n11184), .ZN(n12678) );
  NAND2_X1 U13278 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(P2_U3088), .ZN(n16182) );
  NAND2_X1 U13279 ( .A1(n15018), .A2(n11259), .ZN(n11185) );
  OAI211_X1 U13280 ( .C1(n12994), .C2(n13058), .A(n16182), .B(n11185), .ZN(
        n11187) );
  INV_X1 U13281 ( .A(n13062), .ZN(n11323) );
  INV_X1 U13282 ( .A(n15036), .ZN(n11391) );
  OAI22_X1 U13283 ( .A1(n11323), .A2(n14994), .B1(n14972), .B2(n11391), .ZN(
        n11186) );
  AOI211_X1 U13284 ( .C1(n12678), .C2(n15014), .A(n11187), .B(n11186), .ZN(
        n11188) );
  OAI21_X1 U13285 ( .B1(n11190), .B2(n11189), .A(n11188), .ZN(P2_U3185) );
  NOR2_X1 U13286 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n14535), .ZN(n11508) );
  OR3_X1 U13287 ( .A1(n11193), .A2(n11192), .A3(n11191), .ZN(n11194) );
  AOI21_X1 U13288 ( .B1(n11195), .B2(n11194), .A(n16423), .ZN(n11196) );
  AOI211_X1 U13289 ( .C1(n16150), .C2(P3_ADDR_REG_4__SCAN_IN), .A(n11508), .B(
        n11196), .ZN(n11203) );
  AND3_X1 U13290 ( .A1(n11198), .A2(n11197), .A3(n7480), .ZN(n11200) );
  OAI21_X1 U13291 ( .B1(n11201), .B2(n11200), .A(n11199), .ZN(n11202) );
  OAI211_X1 U13292 ( .C1(n16427), .C2(n7686), .A(n11203), .B(n11202), .ZN(
        n11211) );
  INV_X1 U13293 ( .A(n11204), .ZN(n11205) );
  NAND3_X1 U13294 ( .A1(n11207), .A2(n11206), .A3(n11205), .ZN(n11208) );
  AOI21_X1 U13295 ( .B1(n11209), .B2(n11208), .A(n16418), .ZN(n11210) );
  OR2_X1 U13296 ( .A1(n11211), .A2(n11210), .ZN(P3_U3186) );
  NOR3_X1 U13297 ( .A1(n16429), .A2(P3_REG1_REG_2__SCAN_IN), .A3(n11221), .ZN(
        n11214) );
  NOR4_X1 U13298 ( .A1(n11212), .A2(P3_REG2_REG_2__SCAN_IN), .A3(n14139), .A4(
        n11218), .ZN(n11213) );
  NOR3_X1 U13299 ( .A1(n11214), .A2(n14146), .A3(n11213), .ZN(n11235) );
  INV_X1 U13300 ( .A(n11215), .ZN(n11219) );
  INV_X1 U13301 ( .A(n11216), .ZN(n11217) );
  AOI211_X1 U13302 ( .C1(n11219), .C2(n11218), .A(n11217), .B(n16423), .ZN(
        n11232) );
  AOI211_X1 U13303 ( .C1(n11222), .C2(n11221), .A(n11220), .B(n16429), .ZN(
        n11231) );
  INV_X1 U13304 ( .A(n11223), .ZN(n11225) );
  NAND3_X1 U13305 ( .A1(n11226), .A2(n11225), .A3(n11224), .ZN(n11227) );
  AOI21_X1 U13306 ( .B1(n11228), .B2(n11227), .A(n16418), .ZN(n11230) );
  OAI22_X1 U13307 ( .A1(n16438), .A2(n16281), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n16509), .ZN(n11229) );
  NOR4_X1 U13308 ( .A1(n11232), .A2(n11231), .A3(n11230), .A4(n11229), .ZN(
        n11233) );
  OAI21_X1 U13309 ( .B1(n11235), .B2(n11234), .A(n11233), .ZN(P3_U3184) );
  XNOR2_X1 U13310 ( .A(n13062), .B(n13064), .ZN(n13319) );
  NAND2_X1 U13311 ( .A1(n11237), .A2(n15038), .ZN(n11239) );
  INV_X1 U13312 ( .A(n11383), .ZN(n11240) );
  AOI21_X1 U13313 ( .B1(n11386), .B2(n11241), .A(n11240), .ZN(n11315) );
  NOR2_X1 U13314 ( .A1(n16152), .A2(n11242), .ZN(n16151) );
  NAND2_X1 U13315 ( .A1(n16151), .A2(n11243), .ZN(n11244) );
  NAND2_X1 U13316 ( .A1(n13223), .A2(n13342), .ZN(n11279) );
  INV_X1 U13317 ( .A(n11279), .ZN(n11247) );
  NAND2_X1 U13318 ( .A1(n15353), .A2(n11247), .ZN(n15336) );
  AND2_X1 U13319 ( .A1(n11265), .A2(n13054), .ZN(n11248) );
  XNOR2_X1 U13320 ( .A(n16586), .B(n15038), .ZN(n13315) );
  INV_X1 U13321 ( .A(n13315), .ZN(n11266) );
  NAND2_X1 U13322 ( .A1(n16586), .A2(n13058), .ZN(n11251) );
  NAND2_X1 U13323 ( .A1(n11269), .A2(n11251), .ZN(n11387) );
  XNOR2_X1 U13324 ( .A(n11387), .B(n11386), .ZN(n11253) );
  OAI22_X1 U13325 ( .A1(n11391), .A2(n15287), .B1(n13058), .B2(n15289), .ZN(
        n11252) );
  AOI21_X1 U13326 ( .B1(n11253), .B2(n15346), .A(n11252), .ZN(n11254) );
  OAI21_X1 U13327 ( .B1(n11315), .B2(n10226), .A(n11254), .ZN(n11316) );
  INV_X1 U13328 ( .A(n11316), .ZN(n11255) );
  MUX2_X1 U13329 ( .A(n11256), .B(n11255), .S(n15327), .Z(n11263) );
  OAI21_X1 U13330 ( .B1(n7421), .B2(n11323), .A(n14960), .ZN(n11257) );
  NOR2_X1 U13331 ( .A1(n11257), .A2(n11642), .ZN(n11317) );
  INV_X1 U13332 ( .A(n11259), .ZN(n11260) );
  OAI22_X1 U13333 ( .A1(n15330), .A2(n11323), .B1(n11260), .B2(n15364), .ZN(
        n11261) );
  AOI21_X1 U13334 ( .B1(n15371), .B2(n11317), .A(n11261), .ZN(n11262) );
  OAI211_X1 U13335 ( .C1(n11315), .C2(n15336), .A(n11263), .B(n11262), .ZN(
        P2_U3258) );
  XNOR2_X1 U13336 ( .A(n11264), .B(n11266), .ZN(n11272) );
  INV_X1 U13337 ( .A(n11272), .ZN(n16589) );
  INV_X1 U13338 ( .A(n10226), .ZN(n12139) );
  OAI22_X1 U13339 ( .A1(n13064), .A2(n15287), .B1(n11265), .B2(n15289), .ZN(
        n11271) );
  NAND2_X1 U13340 ( .A1(n11267), .A2(n11266), .ZN(n11268) );
  AOI21_X1 U13341 ( .B1(n11269), .B2(n11268), .A(n15308), .ZN(n11270) );
  AOI211_X1 U13342 ( .C1(n11272), .C2(n12139), .A(n11271), .B(n11270), .ZN(
        n16588) );
  MUX2_X1 U13343 ( .A(n11273), .B(n16588), .S(n15353), .Z(n11278) );
  AOI211_X1 U13344 ( .C1(n16586), .C2(n11274), .A(n14937), .B(n7421), .ZN(
        n16585) );
  OAI22_X1 U13345 ( .A1(n15330), .A2(n7669), .B1(n15364), .B2(n11275), .ZN(
        n11276) );
  AOI21_X1 U13346 ( .B1(n15371), .B2(n16585), .A(n11276), .ZN(n11277) );
  OAI211_X1 U13347 ( .C1(n16589), .C2(n15336), .A(n11278), .B(n11277), .ZN(
        P2_U3259) );
  NAND2_X1 U13348 ( .A1(n10226), .A2(n11279), .ZN(n11280) );
  INV_X1 U13349 ( .A(n11281), .ZN(n11292) );
  INV_X1 U13350 ( .A(n11282), .ZN(n11283) );
  OAI22_X1 U13351 ( .A1(n15330), .A2(n11284), .B1(n11283), .B2(n15364), .ZN(
        n11285) );
  AOI21_X1 U13352 ( .B1(n15371), .B2(n11286), .A(n11285), .ZN(n11291) );
  INV_X1 U13353 ( .A(n11287), .ZN(n11288) );
  MUX2_X1 U13354 ( .A(n11289), .B(n11288), .S(n15353), .Z(n11290) );
  OAI211_X1 U13355 ( .C1(n15359), .C2(n11292), .A(n11291), .B(n11290), .ZN(
        P2_U3261) );
  INV_X1 U13356 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n11293) );
  OAI22_X1 U13357 ( .A1(n15330), .A2(n11294), .B1(n11293), .B2(n15364), .ZN(
        n11295) );
  AOI21_X1 U13358 ( .B1(n15371), .B2(n11296), .A(n11295), .ZN(n11300) );
  MUX2_X1 U13359 ( .A(n11298), .B(n11297), .S(n15353), .Z(n11299) );
  OAI211_X1 U13360 ( .C1(n15359), .C2(n11301), .A(n11300), .B(n11299), .ZN(
        P2_U3264) );
  NAND3_X1 U13361 ( .A1(n16429), .A2(n16423), .A3(n16418), .ZN(n11312) );
  NAND2_X1 U13362 ( .A1(n16429), .A2(n16418), .ZN(n11305) );
  INV_X1 U13363 ( .A(n11302), .ZN(n11303) );
  NAND3_X1 U13364 ( .A1(n11305), .A2(n11304), .A3(n11303), .ZN(n11309) );
  NOR2_X1 U13365 ( .A1(n11306), .A2(P3_STATE_REG_SCAN_IN), .ZN(n11307) );
  AOI21_X1 U13366 ( .B1(n16150), .B2(P3_ADDR_REG_0__SCAN_IN), .A(n11307), .ZN(
        n11308) );
  OAI211_X1 U13367 ( .C1(n11310), .C2(n16423), .A(n11309), .B(n11308), .ZN(
        n11311) );
  AOI21_X1 U13368 ( .B1(n11313), .B2(n11312), .A(n11311), .ZN(n11314) );
  OAI21_X1 U13369 ( .B1(n11304), .B2(n16427), .A(n11314), .ZN(P3_U3182) );
  INV_X1 U13370 ( .A(n11315), .ZN(n11318) );
  AOI211_X1 U13371 ( .C1(n16704), .C2(n11318), .A(n11317), .B(n11316), .ZN(
        n11326) );
  INV_X1 U13372 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n11319) );
  OAI22_X1 U13373 ( .A1(n15517), .A2(n11323), .B1(n16751), .B2(n11319), .ZN(
        n11320) );
  INV_X1 U13374 ( .A(n11320), .ZN(n11321) );
  OAI21_X1 U13375 ( .B1(n11326), .B2(n16748), .A(n11321), .ZN(P2_U3451) );
  OAI22_X1 U13376 ( .A1(n15464), .A2(n11323), .B1(n16747), .B2(n11322), .ZN(
        n11324) );
  INV_X1 U13377 ( .A(n11324), .ZN(n11325) );
  OAI21_X1 U13378 ( .B1(n11326), .B2(n16746), .A(n11325), .ZN(P2_U3506) );
  NAND2_X1 U13379 ( .A1(n11327), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n11738) );
  XNOR2_X1 U13380 ( .A(n11738), .B(P2_IR_REG_17__SCAN_IN), .ZN(n12194) );
  INV_X1 U13381 ( .A(n12194), .ZN(n12109) );
  OAI222_X1 U13382 ( .A1(n15545), .A2(n11329), .B1(n15540), .B2(n11328), .C1(
        P2_U3088), .C2(n12109), .ZN(P2_U3310) );
  NOR2_X1 U13383 ( .A1(n13970), .A2(P3_U3151), .ZN(n16454) );
  XNOR2_X1 U13384 ( .A(n9516), .B(n11530), .ZN(n11330) );
  INV_X1 U13385 ( .A(n11330), .ZN(n11332) );
  XNOR2_X1 U13386 ( .A(n11330), .B(n16497), .ZN(n11529) );
  MUX2_X1 U13387 ( .A(n9516), .B(n11534), .S(n16450), .Z(n11528) );
  NOR2_X1 U13388 ( .A1(n11529), .A2(n11528), .ZN(n11527) );
  AOI211_X1 U13389 ( .C1(n11333), .C2(n11332), .A(n11331), .B(n11527), .ZN(
        n11336) );
  INV_X1 U13390 ( .A(n11334), .ZN(n11335) );
  OAI21_X1 U13391 ( .B1(n11336), .B2(n11335), .A(n16451), .ZN(n11339) );
  INV_X1 U13392 ( .A(n13947), .ZN(n13982) );
  OAI22_X1 U13393 ( .A1(n13978), .A2(n11828), .B1(n13985), .B2(n16494), .ZN(
        n11337) );
  AOI21_X1 U13394 ( .B1(n13982), .B2(n16497), .A(n11337), .ZN(n11338) );
  OAI211_X1 U13395 ( .C1(n16454), .C2(n16509), .A(n11339), .B(n11338), .ZN(
        P3_U3177) );
  NAND2_X1 U13396 ( .A1(n11340), .A2(n13579), .ZN(n11343) );
  NAND2_X1 U13397 ( .A1(n11341), .A2(n15687), .ZN(n11342) );
  XNOR2_X1 U13398 ( .A(n11537), .B(n13580), .ZN(n16609) );
  NAND2_X1 U13399 ( .A1(n11344), .A2(n15687), .ZN(n11348) );
  INV_X1 U13400 ( .A(n11345), .ZN(n11346) );
  NAND2_X1 U13401 ( .A1(n11346), .A2(n13689), .ZN(n11347) );
  XNOR2_X1 U13402 ( .A(n11572), .B(n13580), .ZN(n16611) );
  NAND2_X1 U13403 ( .A1(n16611), .A2(n15935), .ZN(n11355) );
  AOI211_X1 U13404 ( .C1(n16607), .C2(n11349), .A(n16464), .B(n11748), .ZN(
        n16604) );
  NAND2_X1 U13405 ( .A1(n16628), .A2(n16607), .ZN(n11351) );
  MUX2_X1 U13406 ( .A(n16603), .B(n10158), .S(n7414), .Z(n11350) );
  OAI211_X1 U13407 ( .C1(n16622), .C2(n11352), .A(n11351), .B(n11350), .ZN(
        n11353) );
  AOI21_X1 U13408 ( .B1(n16604), .B2(n16486), .A(n11353), .ZN(n11354) );
  OAI211_X1 U13409 ( .C1(n16609), .C2(n15947), .A(n11355), .B(n11354), .ZN(
        P1_U3286) );
  NAND2_X1 U13410 ( .A1(n11356), .A2(n14901), .ZN(n11357) );
  OAI211_X1 U13411 ( .C1(n12618), .C2(n14920), .A(n11357), .B(n13560), .ZN(
        P3_U3272) );
  INV_X1 U13412 ( .A(n11364), .ZN(n11359) );
  NAND2_X1 U13413 ( .A1(n11359), .A2(n11358), .ZN(n11360) );
  NAND2_X1 U13414 ( .A1(n11851), .A2(n12053), .ZN(n11363) );
  AOI22_X1 U13415 ( .A1(n16184), .A2(n12596), .B1(n12597), .B2(
        P1_DATAO_REG_11__SCAN_IN), .ZN(n11362) );
  XNOR2_X1 U13416 ( .A(n15368), .B(n14959), .ZN(n11791) );
  NAND2_X1 U13417 ( .A1(n15033), .A2(n14937), .ZN(n11792) );
  XNOR2_X1 U13418 ( .A(n11791), .B(n11792), .ZN(n11365) );
  AOI22_X1 U13419 ( .A1(n11364), .A2(n15014), .B1(n14961), .B2(n15034), .ZN(
        n11366) );
  NOR3_X1 U13420 ( .A1(n11367), .A2(n11366), .A3(n11365), .ZN(n11380) );
  NAND2_X1 U13421 ( .A1(n10847), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n11374) );
  NAND2_X1 U13422 ( .A1(n9790), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n11373) );
  NAND2_X1 U13423 ( .A1(n11369), .A2(n11368), .ZN(n11370) );
  AND2_X1 U13424 ( .A1(n11768), .A2(n11370), .ZN(n12698) );
  NAND2_X1 U13425 ( .A1(n9786), .A2(n12698), .ZN(n11372) );
  NAND2_X1 U13426 ( .A1(n9789), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n11371) );
  NAND4_X1 U13427 ( .A1(n11374), .A2(n11373), .A3(n11372), .A4(n11371), .ZN(
        n15032) );
  INV_X1 U13428 ( .A(n11375), .ZN(n15365) );
  NAND2_X1 U13429 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(P2_U3088), .ZN(n16196)
         );
  OAI21_X1 U13430 ( .B1(n15003), .B2(n15365), .A(n16196), .ZN(n11376) );
  AOI21_X1 U13431 ( .B1(n14974), .B2(n15034), .A(n11376), .ZN(n11378) );
  NAND2_X1 U13432 ( .A1(n15368), .A2(n15024), .ZN(n11377) );
  OAI211_X1 U13433 ( .C1(n12137), .C2(n14972), .A(n11378), .B(n11377), .ZN(
        n11379) );
  NOR2_X1 U13434 ( .A1(n11380), .A2(n11379), .ZN(n11381) );
  OAI21_X1 U13435 ( .B1(n12706), .B2(n15021), .A(n11381), .ZN(P2_U3208) );
  OR2_X1 U13436 ( .A1(n13062), .A2(n15037), .ZN(n11382) );
  NAND2_X1 U13437 ( .A1(n13071), .A2(n15036), .ZN(n11385) );
  OR2_X1 U13438 ( .A1(n13071), .A2(n15036), .ZN(n11384) );
  NAND2_X1 U13439 ( .A1(n11385), .A2(n11384), .ZN(n13317) );
  XNOR2_X1 U13440 ( .A(n13077), .B(n13079), .ZN(n13320) );
  XNOR2_X1 U13441 ( .A(n11590), .B(n13320), .ZN(n11622) );
  NAND2_X1 U13442 ( .A1(n11387), .A2(n11386), .ZN(n11389) );
  NAND2_X1 U13443 ( .A1(n13062), .A2(n13064), .ZN(n11388) );
  AND2_X1 U13444 ( .A1(n13071), .A2(n11391), .ZN(n11390) );
  XNOR2_X1 U13445 ( .A(n11587), .B(n13320), .ZN(n11393) );
  OAI22_X1 U13446 ( .A1(n12664), .A2(n15287), .B1(n11391), .B2(n15289), .ZN(
        n11392) );
  AOI21_X1 U13447 ( .B1(n11393), .B2(n15346), .A(n11392), .ZN(n11394) );
  OAI21_X1 U13448 ( .B1(n11622), .B2(n10226), .A(n11394), .ZN(n11623) );
  NAND2_X1 U13449 ( .A1(n11623), .A2(n15327), .ZN(n11399) );
  INV_X1 U13450 ( .A(n13071), .ZN(n16639) );
  INV_X1 U13451 ( .A(n11596), .ZN(n11598) );
  AOI211_X1 U13452 ( .C1(n13077), .C2(n11641), .A(n14937), .B(n11598), .ZN(
        n11624) );
  INV_X1 U13453 ( .A(n13077), .ZN(n11630) );
  INV_X1 U13454 ( .A(n15364), .ZN(n15292) );
  AOI22_X1 U13455 ( .A1(n15362), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n11395), 
        .B2(n15292), .ZN(n11396) );
  OAI21_X1 U13456 ( .B1(n11630), .B2(n15330), .A(n11396), .ZN(n11397) );
  AOI21_X1 U13457 ( .B1(n11624), .B2(n15371), .A(n11397), .ZN(n11398) );
  OAI211_X1 U13458 ( .C1(n11622), .C2(n15336), .A(n11399), .B(n11398), .ZN(
        P2_U3256) );
  INV_X1 U13459 ( .A(n11400), .ZN(n11401) );
  XNOR2_X1 U13460 ( .A(n13525), .B(n11401), .ZN(n16455) );
  NAND2_X1 U13461 ( .A1(n13357), .A2(n16510), .ZN(n11813) );
  INV_X1 U13462 ( .A(n11813), .ZN(n16515) );
  INV_X1 U13463 ( .A(n14240), .ZN(n14388) );
  OAI21_X1 U13464 ( .B1(n13525), .B2(n11403), .A(n11402), .ZN(n11406) );
  OAI22_X1 U13465 ( .A1(n11404), .A2(n14312), .B1(n11817), .B2(n14314), .ZN(
        n11405) );
  AOI21_X1 U13466 ( .B1(n11406), .B2(n16501), .A(n11405), .ZN(n11407) );
  OAI21_X1 U13467 ( .B1(n16455), .B2(n16521), .A(n11407), .ZN(n16457) );
  NAND2_X1 U13468 ( .A1(n11408), .A2(n16652), .ZN(n16456) );
  OAI22_X1 U13469 ( .A1(n11531), .A2(n16508), .B1(n16456), .B2(n16510), .ZN(
        n11409) );
  NOR2_X1 U13470 ( .A1(n16457), .A2(n11409), .ZN(n11410) );
  MUX2_X1 U13471 ( .A(n11411), .B(n11410), .S(n14352), .Z(n11412) );
  OAI21_X1 U13472 ( .B1(n16455), .B2(n14388), .A(n11412), .ZN(P3_U3232) );
  INV_X1 U13473 ( .A(n11413), .ZN(n11415) );
  AOI211_X1 U13474 ( .C1(n13223), .C2(n11415), .A(n11414), .B(n15362), .ZN(
        n11416) );
  AOI21_X1 U13475 ( .B1(n15292), .B2(P2_REG3_REG_0__SCAN_IN), .A(n11416), .ZN(
        n11418) );
  NAND2_X1 U13476 ( .A1(n15362), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n11417) );
  OAI211_X1 U13477 ( .C1(n15336), .C2(n13308), .A(n11418), .B(n11417), .ZN(
        P2_U3265) );
  AOI211_X1 U13478 ( .C1(n11421), .C2(n11420), .A(n13954), .B(n11419), .ZN(
        n11422) );
  INV_X1 U13479 ( .A(n11422), .ZN(n11426) );
  INV_X1 U13480 ( .A(n13985), .ZN(n16449) );
  OAI22_X1 U13481 ( .A1(n11817), .A2(n13947), .B1(n13978), .B2(n11925), .ZN(
        n11423) );
  AOI211_X1 U13482 ( .C1(n16449), .C2(n16524), .A(n11424), .B(n11423), .ZN(
        n11425) );
  OAI211_X1 U13483 ( .C1(P3_REG3_REG_3__SCAN_IN), .C2(n13979), .A(n11426), .B(
        n11425), .ZN(P3_U3158) );
  INV_X1 U13484 ( .A(n15826), .ZN(n16633) );
  INV_X1 U13485 ( .A(n11427), .ZN(n11428) );
  INV_X1 U13486 ( .A(n16622), .ZN(n15991) );
  AOI22_X1 U13487 ( .A1(n16628), .A2(n13689), .B1(n11428), .B2(n15991), .ZN(
        n11429) );
  OAI21_X1 U13488 ( .B1(n16631), .B2(n11430), .A(n11429), .ZN(n11433) );
  MUX2_X1 U13489 ( .A(n11431), .B(P1_REG2_REG_6__SCAN_IN), .S(n7414), .Z(
        n11432) );
  AOI211_X1 U13490 ( .C1(n16633), .C2(n11434), .A(n11433), .B(n11432), .ZN(
        n11435) );
  INV_X1 U13491 ( .A(n11435), .ZN(P1_U3287) );
  NAND2_X1 U13492 ( .A1(n11436), .A2(n13578), .ZN(n11437) );
  NAND2_X1 U13493 ( .A1(n11438), .A2(n11437), .ZN(n16575) );
  AOI21_X1 U13494 ( .B1(n11439), .B2(n13685), .A(n16464), .ZN(n11441) );
  NAND2_X1 U13495 ( .A1(n11441), .A2(n11440), .ZN(n16571) );
  INV_X1 U13496 ( .A(n11442), .ZN(n11443) );
  AOI22_X1 U13497 ( .A1(n16628), .A2(n13685), .B1(n15991), .B2(n11443), .ZN(
        n11444) );
  OAI21_X1 U13498 ( .B1(n16631), .B2(n16571), .A(n11444), .ZN(n11452) );
  NAND2_X1 U13499 ( .A1(n16575), .A2(n16472), .ZN(n11450) );
  XNOR2_X1 U13500 ( .A(n11446), .B(n11445), .ZN(n11447) );
  NAND2_X1 U13501 ( .A1(n11447), .A2(n16561), .ZN(n11449) );
  AOI22_X1 U13502 ( .A1(n15971), .A2(n15689), .B1(n15687), .B2(n16462), .ZN(
        n11448) );
  NAND3_X1 U13503 ( .A1(n11450), .A2(n11449), .A3(n11448), .ZN(n16573) );
  MUX2_X1 U13504 ( .A(n16573), .B(P1_REG2_REG_5__SCAN_IN), .S(n7414), .Z(
        n11451) );
  AOI211_X1 U13505 ( .C1(n16633), .C2(n16575), .A(n11452), .B(n11451), .ZN(
        n11453) );
  INV_X1 U13506 ( .A(n11453), .ZN(P1_U3288) );
  INV_X1 U13507 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n11454) );
  NAND2_X1 U13508 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(P2_U3088), .ZN(n12077)
         );
  OAI21_X1 U13509 ( .B1(n16237), .B2(n11454), .A(n12077), .ZN(n11465) );
  OAI21_X1 U13510 ( .B1(n11807), .B2(n11456), .A(n11455), .ZN(n11483) );
  XNOR2_X1 U13511 ( .A(n11483), .B(n11457), .ZN(n11458) );
  NAND2_X1 U13512 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n11458), .ZN(n11484) );
  OAI211_X1 U13513 ( .C1(n11458), .C2(P2_REG1_REG_15__SCAN_IN), .A(n16233), 
        .B(n11484), .ZN(n11463) );
  NAND2_X1 U13514 ( .A1(n12057), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n11460) );
  NAND2_X1 U13515 ( .A1(n11460), .A2(n11459), .ZN(n11493) );
  XOR2_X1 U13516 ( .A(n12054), .B(n11493), .Z(n11461) );
  NAND2_X1 U13517 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n11461), .ZN(n11494) );
  OAI211_X1 U13518 ( .C1(P2_REG2_REG_15__SCAN_IN), .C2(n11461), .A(n16229), 
        .B(n11494), .ZN(n11462) );
  NAND2_X1 U13519 ( .A1(n11463), .A2(n11462), .ZN(n11464) );
  AOI211_X1 U13520 ( .C1(n16231), .C2(n12054), .A(n11465), .B(n11464), .ZN(
        n11466) );
  INV_X1 U13521 ( .A(n11466), .ZN(P2_U3229) );
  INV_X1 U13522 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n12490) );
  MUX2_X1 U13523 ( .A(n12490), .B(P1_REG1_REG_14__SCAN_IN), .S(n12319), .Z(
        n11469) );
  OAI21_X1 U13524 ( .B1(n11473), .B2(n16733), .A(n11467), .ZN(n11468) );
  AOI21_X1 U13525 ( .B1(n11469), .B2(n11468), .A(n11890), .ZN(n11482) );
  NAND2_X1 U13526 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n12531)
         );
  INV_X1 U13527 ( .A(n12531), .ZN(n11471) );
  NOR2_X1 U13528 ( .A1(n15727), .A2(n11894), .ZN(n11470) );
  AOI211_X1 U13529 ( .C1(n16246), .C2(P1_ADDR_REG_14__SCAN_IN), .A(n11471), 
        .B(n11470), .ZN(n11481) );
  INV_X1 U13530 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n11472) );
  MUX2_X1 U13531 ( .A(n11472), .B(P1_REG2_REG_14__SCAN_IN), .S(n12319), .Z(
        n11475) );
  NOR2_X1 U13532 ( .A1(n11473), .A2(n12023), .ZN(n11477) );
  INV_X1 U13533 ( .A(n11477), .ZN(n11474) );
  NAND2_X1 U13534 ( .A1(n11475), .A2(n11474), .ZN(n11478) );
  MUX2_X1 U13535 ( .A(P1_REG2_REG_14__SCAN_IN), .B(n11472), .S(n12319), .Z(
        n11476) );
  OAI21_X1 U13536 ( .B1(n11479), .B2(n11477), .A(n11476), .ZN(n11893) );
  OAI211_X1 U13537 ( .C1(n11479), .C2(n11478), .A(n11893), .B(n16263), .ZN(
        n11480) );
  OAI211_X1 U13538 ( .C1(n11482), .C2(n15710), .A(n11481), .B(n11480), .ZN(
        P1_U3257) );
  NAND2_X1 U13539 ( .A1(n12054), .A2(n11483), .ZN(n11485) );
  NAND2_X1 U13540 ( .A1(n11485), .A2(n11484), .ZN(n16201) );
  INV_X1 U13541 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n11486) );
  XNOR2_X1 U13542 ( .A(n12170), .B(n11486), .ZN(n16202) );
  NAND2_X1 U13543 ( .A1(n16201), .A2(n16202), .ZN(n11488) );
  NAND2_X1 U13544 ( .A1(n12170), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n11487) );
  NAND2_X1 U13545 ( .A1(n11488), .A2(n11487), .ZN(n12103) );
  INV_X1 U13546 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n15451) );
  XNOR2_X1 U13547 ( .A(n12194), .B(n15451), .ZN(n12102) );
  XNOR2_X1 U13548 ( .A(n12103), .B(n12102), .ZN(n11502) );
  NAND2_X1 U13549 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(P2_U3088), .ZN(n12206)
         );
  INV_X1 U13550 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n11490) );
  NOR2_X1 U13551 ( .A1(n12109), .A2(n11490), .ZN(n11489) );
  AOI21_X1 U13552 ( .B1(n11490), .B2(n12109), .A(n11489), .ZN(n11498) );
  NAND2_X1 U13553 ( .A1(n12170), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n11496) );
  INV_X1 U13554 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n11492) );
  INV_X1 U13555 ( .A(n11496), .ZN(n11491) );
  AOI21_X1 U13556 ( .B1(n11492), .B2(n16199), .A(n11491), .ZN(n16206) );
  NAND2_X1 U13557 ( .A1(n12054), .A2(n11493), .ZN(n11495) );
  NAND2_X1 U13558 ( .A1(n11495), .A2(n11494), .ZN(n16205) );
  NAND2_X1 U13559 ( .A1(n16206), .A2(n16205), .ZN(n16204) );
  NAND2_X1 U13560 ( .A1(n11496), .A2(n16204), .ZN(n11497) );
  NAND2_X1 U13561 ( .A1(n11498), .A2(n11497), .ZN(n12108) );
  OAI211_X1 U13562 ( .C1(n11498), .C2(n11497), .A(n16229), .B(n12108), .ZN(
        n11499) );
  AND2_X1 U13563 ( .A1(n12206), .A2(n11499), .ZN(n11501) );
  AOI22_X1 U13564 ( .A1(n10096), .A2(P2_ADDR_REG_17__SCAN_IN), .B1(n16231), 
        .B2(n12194), .ZN(n11500) );
  OAI211_X1 U13565 ( .C1(n11502), .C2(n16190), .A(n11501), .B(n11500), .ZN(
        P2_U3231) );
  OAI21_X1 U13566 ( .B1(n11505), .B2(n11504), .A(n11503), .ZN(n11506) );
  NAND2_X1 U13567 ( .A1(n11506), .A2(n16451), .ZN(n11510) );
  OAI22_X1 U13568 ( .A1(n11829), .A2(n13978), .B1(n13947), .B2(n11828), .ZN(
        n11507) );
  AOI211_X1 U13569 ( .C1(n16449), .C2(n11836), .A(n11508), .B(n11507), .ZN(
        n11509) );
  OAI211_X1 U13570 ( .C1(n11834), .C2(n13979), .A(n11510), .B(n11509), .ZN(
        P3_U3170) );
  INV_X1 U13571 ( .A(n11511), .ZN(n11512) );
  AOI21_X1 U13572 ( .B1(n11514), .B2(n11513), .A(n11512), .ZN(n11526) );
  AOI21_X1 U13573 ( .B1(n11516), .B2(n9620), .A(n11515), .ZN(n11522) );
  NOR2_X1 U13574 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n8861), .ZN(n11844) );
  AOI21_X1 U13575 ( .B1(n11518), .B2(n9621), .A(n11517), .ZN(n11519) );
  NOR2_X1 U13576 ( .A1(n16423), .A2(n11519), .ZN(n11520) );
  AOI211_X1 U13577 ( .C1(n16150), .C2(P3_ADDR_REG_7__SCAN_IN), .A(n11844), .B(
        n11520), .ZN(n11521) );
  OAI21_X1 U13578 ( .B1(n11522), .B2(n16429), .A(n11521), .ZN(n11523) );
  AOI21_X1 U13579 ( .B1(n11524), .B2(n14146), .A(n11523), .ZN(n11525) );
  OAI21_X1 U13580 ( .B1(n11526), .B2(n16418), .A(n11525), .ZN(P3_U3189) );
  AOI21_X1 U13581 ( .B1(n11529), .B2(n11528), .A(n11527), .ZN(n11536) );
  OAI22_X1 U13582 ( .A1(n13978), .A2(n11817), .B1(n13985), .B2(n11530), .ZN(
        n11533) );
  NOR2_X1 U13583 ( .A1(n16454), .A2(n11531), .ZN(n11532) );
  AOI211_X1 U13584 ( .C1(n13982), .C2(n11534), .A(n11533), .B(n11532), .ZN(
        n11535) );
  OAI21_X1 U13585 ( .B1(n11536), .B2(n13954), .A(n11535), .ZN(P3_U3162) );
  NAND2_X1 U13586 ( .A1(n16607), .A2(n8629), .ZN(n11538) );
  NAND2_X1 U13587 ( .A1(n11539), .A2(n11544), .ZN(n11542) );
  AOI22_X1 U13588 ( .A1(n12760), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n12759), 
        .B2(n11540), .ZN(n11541) );
  NAND2_X1 U13589 ( .A1(n11542), .A2(n11541), .ZN(n16627) );
  XNOR2_X1 U13590 ( .A(n16627), .B(n11686), .ZN(n13582) );
  OR2_X1 U13591 ( .A1(n16627), .A2(n11686), .ZN(n11543) );
  NAND2_X1 U13592 ( .A1(n11545), .A2(n11544), .ZN(n11548) );
  AOI22_X1 U13593 ( .A1(n12760), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n12759), 
        .B2(n11546), .ZN(n11547) );
  NAND2_X1 U13594 ( .A1(n11548), .A2(n11547), .ZN(n13711) );
  NAND2_X1 U13595 ( .A1(n13566), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n11555) );
  OR2_X1 U13596 ( .A1(n12862), .A2(n11549), .ZN(n11554) );
  OR2_X1 U13597 ( .A1(n12929), .A2(n10304), .ZN(n11553) );
  NAND2_X1 U13598 ( .A1(n11550), .A2(n11704), .ZN(n11551) );
  NAND2_X1 U13599 ( .A1(n11565), .A2(n11551), .ZN(n11701) );
  OR2_X1 U13600 ( .A1(n12946), .A2(n11701), .ZN(n11552) );
  NAND4_X1 U13601 ( .A1(n11555), .A2(n11554), .A3(n11553), .A4(n11552), .ZN(
        n15684) );
  NAND2_X1 U13602 ( .A1(n13711), .A2(n11696), .ZN(n11556) );
  OR2_X1 U13603 ( .A1(n13711), .A2(n11696), .ZN(n11557) );
  NAND2_X1 U13604 ( .A1(n11558), .A2(n11544), .ZN(n11561) );
  AOI22_X1 U13605 ( .A1(n11559), .A2(n12759), .B1(n12760), .B2(
        P2_DATAO_REG_10__SCAN_IN), .ZN(n11560) );
  NAND2_X1 U13606 ( .A1(n11561), .A2(n11560), .ZN(n13715) );
  NAND2_X1 U13607 ( .A1(n12945), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n11571) );
  OR2_X1 U13608 ( .A1(n12929), .A2(n11562), .ZN(n11570) );
  INV_X1 U13609 ( .A(n11563), .ZN(n11858) );
  NAND2_X1 U13610 ( .A1(n11565), .A2(n11564), .ZN(n11566) );
  NAND2_X1 U13611 ( .A1(n11858), .A2(n11566), .ZN(n12122) );
  OR2_X1 U13612 ( .A1(n12946), .A2(n12122), .ZN(n11569) );
  INV_X1 U13613 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n11567) );
  OR2_X1 U13614 ( .A1(n10418), .A2(n11567), .ZN(n11568) );
  NAND4_X1 U13615 ( .A1(n11571), .A2(n11570), .A3(n11569), .A4(n11568), .ZN(
        n15683) );
  INV_X1 U13616 ( .A(n15683), .ZN(n11979) );
  XNOR2_X1 U13617 ( .A(n13715), .B(n11979), .ZN(n13585) );
  INV_X1 U13618 ( .A(n13585), .ZN(n11847) );
  XNOR2_X1 U13619 ( .A(n11848), .B(n11847), .ZN(n16672) );
  XNOR2_X1 U13620 ( .A(n13711), .B(n11696), .ZN(n13583) );
  OR2_X1 U13621 ( .A1(n13711), .A2(n15684), .ZN(n11573) );
  NAND2_X1 U13622 ( .A1(n11906), .A2(n11573), .ZN(n11574) );
  OAI21_X1 U13623 ( .B1(n11574), .B2(n13585), .A(n11869), .ZN(n16675) );
  NAND2_X1 U13624 ( .A1(n13566), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n11579) );
  OR2_X1 U13625 ( .A1(n12862), .A2(n11575), .ZN(n11578) );
  OR2_X1 U13626 ( .A1(n12929), .A2(n10750), .ZN(n11577) );
  INV_X1 U13627 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n11857) );
  XNOR2_X1 U13628 ( .A(n11858), .B(n11857), .ZN(n11989) );
  OR2_X1 U13629 ( .A1(n12946), .A2(n11989), .ZN(n11576) );
  NAND4_X1 U13630 ( .A1(n11579), .A2(n11578), .A3(n11577), .A4(n11576), .ZN(
        n15682) );
  INV_X1 U13631 ( .A(n16627), .ZN(n11749) );
  NAND2_X1 U13632 ( .A1(n11748), .A2(n11749), .ZN(n11908) );
  OR2_X1 U13633 ( .A1(n11908), .A2(n13711), .ZN(n11909) );
  AOI211_X1 U13634 ( .C1(n13715), .C2(n11909), .A(n16464), .B(n11872), .ZN(
        n11580) );
  AOI21_X1 U13635 ( .B1(n16462), .B2(n15682), .A(n11580), .ZN(n16670) );
  NAND2_X1 U13636 ( .A1(n15684), .A2(n15971), .ZN(n16669) );
  OAI22_X1 U13637 ( .A1(n7414), .A2(n16669), .B1(n12122), .B2(n16622), .ZN(
        n11582) );
  INV_X1 U13638 ( .A(n13715), .ZN(n16671) );
  NOR2_X1 U13639 ( .A1(n16671), .A2(n16481), .ZN(n11581) );
  AOI211_X1 U13640 ( .C1(n7414), .C2(P1_REG2_REG_10__SCAN_IN), .A(n11582), .B(
        n11581), .ZN(n11583) );
  OAI21_X1 U13641 ( .B1(n16670), .B2(n16631), .A(n11583), .ZN(n11584) );
  AOI21_X1 U13642 ( .B1(n16675), .B2(n15935), .A(n11584), .ZN(n11585) );
  OAI21_X1 U13643 ( .B1(n15947), .B2(n16672), .A(n11585), .ZN(P1_U3283) );
  INV_X1 U13644 ( .A(n13320), .ZN(n11586) );
  NAND2_X1 U13645 ( .A1(n11587), .A2(n11586), .ZN(n11589) );
  OR2_X1 U13646 ( .A1(n13077), .A2(n13079), .ZN(n11588) );
  NAND2_X1 U13647 ( .A1(n11589), .A2(n11588), .ZN(n11726) );
  XNOR2_X1 U13648 ( .A(n13083), .B(n12664), .ZN(n13321) );
  INV_X1 U13649 ( .A(n13321), .ZN(n11725) );
  XNOR2_X1 U13650 ( .A(n11726), .B(n11725), .ZN(n11595) );
  NAND2_X1 U13651 ( .A1(n13077), .A2(n15035), .ZN(n11591) );
  OAI21_X1 U13652 ( .B1(n7606), .B2(n13321), .A(n11719), .ZN(n16682) );
  OAI22_X1 U13653 ( .A1(n13089), .A2(n15287), .B1(n13079), .B2(n15289), .ZN(
        n11593) );
  AOI21_X1 U13654 ( .B1(n16682), .B2(n12139), .A(n11593), .ZN(n11594) );
  OAI21_X1 U13655 ( .B1(n15308), .B2(n11595), .A(n11594), .ZN(n16680) );
  INV_X1 U13656 ( .A(n16680), .ZN(n11604) );
  INV_X1 U13657 ( .A(n15336), .ZN(n11782) );
  INV_X1 U13658 ( .A(n13083), .ZN(n16679) );
  INV_X1 U13659 ( .A(n11723), .ZN(n11597) );
  OAI211_X1 U13660 ( .C1(n16679), .C2(n11598), .A(n11597), .B(n14960), .ZN(
        n16677) );
  AOI22_X1 U13661 ( .A1(n15362), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n11599), 
        .B2(n15292), .ZN(n11601) );
  NAND2_X1 U13662 ( .A1(n15367), .A2(n13083), .ZN(n11600) );
  OAI211_X1 U13663 ( .C1(n16677), .C2(n15233), .A(n11601), .B(n11600), .ZN(
        n11602) );
  AOI21_X1 U13664 ( .B1(n16682), .B2(n11782), .A(n11602), .ZN(n11603) );
  OAI21_X1 U13665 ( .B1(n11604), .B2(n15362), .A(n11603), .ZN(P2_U3255) );
  AOI21_X1 U13666 ( .B1(n7629), .B2(n11606), .A(n11605), .ZN(n11621) );
  XNOR2_X1 U13667 ( .A(n11608), .B(n11607), .ZN(n11609) );
  NAND2_X1 U13668 ( .A1(n11609), .A2(n14125), .ZN(n11620) );
  INV_X1 U13669 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n11611) );
  INV_X1 U13670 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n14525) );
  NOR2_X1 U13671 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n14525), .ZN(n11971) );
  INV_X1 U13672 ( .A(n11971), .ZN(n11610) );
  OAI21_X1 U13673 ( .B1(n16438), .B2(n11611), .A(n11610), .ZN(n11617) );
  AOI21_X1 U13674 ( .B1(n11614), .B2(n11613), .A(n11612), .ZN(n11615) );
  NOR2_X1 U13675 ( .A1(n11615), .A2(n16429), .ZN(n11616) );
  AOI211_X1 U13676 ( .C1(n14146), .C2(n11618), .A(n11617), .B(n11616), .ZN(
        n11619) );
  OAI211_X1 U13677 ( .C1(n11621), .C2(n16423), .A(n11620), .B(n11619), .ZN(
        P3_U3190) );
  INV_X1 U13678 ( .A(n11622), .ZN(n11625) );
  AOI211_X1 U13679 ( .C1(n16704), .C2(n11625), .A(n11624), .B(n11623), .ZN(
        n11633) );
  INV_X1 U13680 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n11626) );
  OAI22_X1 U13681 ( .A1(n15517), .A2(n11630), .B1(n16751), .B2(n11626), .ZN(
        n11627) );
  INV_X1 U13682 ( .A(n11627), .ZN(n11628) );
  OAI21_X1 U13683 ( .B1(n11633), .B2(n16748), .A(n11628), .ZN(P2_U3457) );
  OAI22_X1 U13684 ( .A1(n15464), .A2(n11630), .B1(n16747), .B2(n11629), .ZN(
        n11631) );
  INV_X1 U13685 ( .A(n11631), .ZN(n11632) );
  OAI21_X1 U13686 ( .B1(n11633), .B2(n16746), .A(n11632), .ZN(P2_U3508) );
  NOR2_X1 U13687 ( .A1(n14891), .A2(n8968), .ZN(n11634) );
  AOI21_X1 U13688 ( .B1(n14891), .B2(n11635), .A(n11634), .ZN(n11636) );
  OAI21_X1 U13689 ( .B1(n11637), .B2(n14896), .A(n11636), .ZN(P3_U3390) );
  INV_X1 U13690 ( .A(n11638), .ZN(n11639) );
  AOI21_X1 U13691 ( .B1(n13317), .B2(n11640), .A(n11639), .ZN(n16642) );
  OAI211_X1 U13692 ( .C1(n11642), .C2(n16639), .A(n14960), .B(n11641), .ZN(
        n16637) );
  AOI22_X1 U13693 ( .A1(n15367), .A2(n13071), .B1(n12670), .B2(n15292), .ZN(
        n11643) );
  OAI21_X1 U13694 ( .B1(n15233), .B2(n16637), .A(n11643), .ZN(n11644) );
  AOI21_X1 U13695 ( .B1(n16642), .B2(n15369), .A(n11644), .ZN(n11649) );
  XNOR2_X1 U13696 ( .A(n11645), .B(n13317), .ZN(n11646) );
  AOI222_X1 U13697 ( .A1(n15346), .A2(n11646), .B1(n15037), .B2(n15341), .C1(
        n15035), .C2(n15343), .ZN(n16638) );
  MUX2_X1 U13698 ( .A(n11647), .B(n16638), .S(n15327), .Z(n11648) );
  NAND2_X1 U13699 ( .A1(n11649), .A2(n11648), .ZN(P2_U3257) );
  INV_X1 U13700 ( .A(n11650), .ZN(n11657) );
  INV_X1 U13701 ( .A(n11651), .ZN(n11652) );
  OAI22_X1 U13702 ( .A1(n15327), .A2(n10108), .B1(n11652), .B2(n15364), .ZN(
        n11653) );
  AOI21_X1 U13703 ( .B1(n15367), .B2(n13054), .A(n11653), .ZN(n11654) );
  OAI21_X1 U13704 ( .B1(n15233), .B2(n11655), .A(n11654), .ZN(n11656) );
  AOI21_X1 U13705 ( .B1(n11657), .B2(n15369), .A(n11656), .ZN(n11658) );
  OAI21_X1 U13706 ( .B1(n15362), .B2(n11659), .A(n11658), .ZN(P2_U3260) );
  XNOR2_X1 U13707 ( .A(n11661), .B(n11660), .ZN(n11662) );
  NAND2_X1 U13708 ( .A1(n11662), .A2(n16451), .ZN(n11666) );
  OAI22_X1 U13709 ( .A1(n11925), .A2(n13947), .B1(n13978), .B2(n11842), .ZN(
        n11663) );
  AOI211_X1 U13710 ( .C1(n16449), .C2(n11931), .A(n11664), .B(n11663), .ZN(
        n11665) );
  OAI211_X1 U13711 ( .C1(n11929), .C2(n13979), .A(n11666), .B(n11665), .ZN(
        P3_U3167) );
  OAI22_X1 U13712 ( .A1(n15353), .A2(n10104), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(n15364), .ZN(n11667) );
  AOI21_X1 U13713 ( .B1(n15367), .B2(n13035), .A(n11667), .ZN(n11671) );
  AOI22_X1 U13714 ( .A1(n15369), .A2(n11669), .B1(n15371), .B2(n11668), .ZN(
        n11670) );
  OAI211_X1 U13715 ( .C1(n15362), .C2(n11672), .A(n11671), .B(n11670), .ZN(
        P2_U3262) );
  OAI22_X1 U13716 ( .A1(n15353), .A2(n10099), .B1(n11124), .B2(n15364), .ZN(
        n11673) );
  AOI21_X1 U13717 ( .B1(n15367), .B2(n13021), .A(n11673), .ZN(n11677) );
  AOI22_X1 U13718 ( .A1(n15369), .A2(n11675), .B1(n15327), .B2(n11674), .ZN(
        n11676) );
  OAI211_X1 U13719 ( .C1(n15233), .C2(n11678), .A(n11677), .B(n11676), .ZN(
        P2_U3263) );
  OAI211_X1 U13720 ( .C1(n11681), .C2(n11680), .A(n11679), .B(n16451), .ZN(
        n11685) );
  OAI22_X1 U13721 ( .A1(n12240), .A2(n13978), .B1(n13947), .B2(n11829), .ZN(
        n11682) );
  AOI211_X1 U13722 ( .C1(n16449), .C2(n16580), .A(n11683), .B(n11682), .ZN(
        n11684) );
  OAI211_X1 U13723 ( .C1(n12246), .C2(n13979), .A(n11685), .B(n11684), .ZN(
        P3_U3179) );
  INV_X1 U13724 ( .A(n13711), .ZN(n16656) );
  OAI22_X1 U13725 ( .A1(n11749), .A2(n10271), .B1(n11686), .B2(n12846), .ZN(
        n11692) );
  INV_X1 U13726 ( .A(n11692), .ZN(n11695) );
  OAI22_X1 U13727 ( .A1(n11749), .A2(n12940), .B1(n11686), .B2(n10271), .ZN(
        n11687) );
  XNOR2_X1 U13728 ( .A(n11687), .B(n10817), .ZN(n11693) );
  INV_X1 U13729 ( .A(n11693), .ZN(n11694) );
  XNOR2_X1 U13730 ( .A(n11693), .B(n11692), .ZN(n11713) );
  NOR2_X1 U13731 ( .A1(n12846), .A2(n11696), .ZN(n11697) );
  AOI21_X1 U13732 ( .B1(n13711), .B2(n7413), .A(n11697), .ZN(n11978) );
  AOI22_X1 U13733 ( .A1(n13711), .A2(n7412), .B1(n7413), .B2(n15684), .ZN(
        n11698) );
  XNOR2_X1 U13734 ( .A(n11698), .B(n10817), .ZN(n11977) );
  XOR2_X1 U13735 ( .A(n11978), .B(n11977), .Z(n11699) );
  OAI211_X1 U13736 ( .C1(n11700), .C2(n11699), .A(n11976), .B(n16531), .ZN(
        n11707) );
  INV_X1 U13737 ( .A(n11701), .ZN(n11911) );
  INV_X1 U13738 ( .A(n16535), .ZN(n15640) );
  NAND2_X1 U13739 ( .A1(n15658), .A2(n15683), .ZN(n11703) );
  NAND2_X1 U13740 ( .A1(n15659), .A2(n15685), .ZN(n11702) );
  OAI211_X1 U13741 ( .C1(P1_STATE_REG_SCAN_IN), .C2(n11704), .A(n11703), .B(
        n11702), .ZN(n11705) );
  AOI21_X1 U13742 ( .B1(n11911), .B2(n15640), .A(n11705), .ZN(n11706) );
  OAI211_X1 U13743 ( .C1(n16656), .C2(n15653), .A(n11707), .B(n11706), .ZN(
        P1_U3231) );
  NAND2_X1 U13744 ( .A1(n15684), .A2(n16462), .ZN(n11709) );
  NAND2_X1 U13745 ( .A1(n15686), .A2(n15971), .ZN(n11708) );
  NAND2_X1 U13746 ( .A1(n11709), .A2(n11708), .ZN(n11754) );
  NAND2_X1 U13747 ( .A1(n16530), .A2(n11754), .ZN(n11710) );
  OAI211_X1 U13748 ( .C1(n16535), .C2(n16623), .A(n11711), .B(n11710), .ZN(
        n11716) );
  AOI21_X1 U13749 ( .B1(n11713), .B2(n11712), .A(n7621), .ZN(n11714) );
  NOR2_X1 U13750 ( .A1(n11714), .A2(n15673), .ZN(n11715) );
  AOI211_X1 U13751 ( .C1(n15671), .C2(n16627), .A(n11716), .B(n11715), .ZN(
        n11717) );
  INV_X1 U13752 ( .A(n11717), .ZN(P1_U3221) );
  XNOR2_X1 U13753 ( .A(n15368), .B(n13089), .ZN(n13322) );
  INV_X1 U13754 ( .A(n13322), .ZN(n11722) );
  OR2_X1 U13755 ( .A1(n13083), .A2(n15034), .ZN(n11718) );
  INV_X1 U13756 ( .A(n11760), .ZN(n11720) );
  AOI21_X1 U13757 ( .B1(n11722), .B2(n11721), .A(n11720), .ZN(n15370) );
  INV_X1 U13758 ( .A(n15368), .ZN(n11732) );
  OR2_X1 U13759 ( .A1(n11732), .A2(n11723), .ZN(n11724) );
  AND3_X1 U13760 ( .A1(n11777), .A2(n14960), .A3(n11724), .ZN(n15372) );
  OR2_X1 U13761 ( .A1(n13083), .A2(n12664), .ZN(n11727) );
  INV_X1 U13762 ( .A(n11764), .ZN(n11728) );
  AOI21_X1 U13763 ( .B1(n13322), .B2(n11729), .A(n11728), .ZN(n11730) );
  OAI222_X1 U13764 ( .A1(n15287), .A2(n12137), .B1(n15289), .B2(n12664), .C1(
        n15308), .C2(n11730), .ZN(n15363) );
  AOI211_X1 U13765 ( .C1(n15370), .C2(n16641), .A(n15372), .B(n15363), .ZN(
        n11736) );
  INV_X1 U13766 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n11731) );
  OAI22_X1 U13767 ( .A1(n11732), .A2(n15517), .B1(n16751), .B2(n11731), .ZN(
        n11733) );
  INV_X1 U13768 ( .A(n11733), .ZN(n11734) );
  OAI21_X1 U13769 ( .B1(n11736), .B2(n16748), .A(n11734), .ZN(P2_U3463) );
  AOI22_X1 U13770 ( .A1(n15457), .A2(n15368), .B1(n16746), .B2(
        P2_REG1_REG_11__SCAN_IN), .ZN(n11735) );
  OAI21_X1 U13771 ( .B1(n11736), .B2(n16746), .A(n11735), .ZN(P2_U3510) );
  INV_X1 U13772 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n11737) );
  NAND2_X1 U13773 ( .A1(n11738), .A2(n11737), .ZN(n11739) );
  NAND2_X1 U13774 ( .A1(n11739), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n11740) );
  XNOR2_X1 U13775 ( .A(n11740), .B(P2_IR_REG_18__SCAN_IN), .ZN(n12438) );
  INV_X1 U13776 ( .A(n12438), .ZN(n16213) );
  MUX2_X1 U13777 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(P1_DATAO_REG_18__SCAN_IN), 
        .S(n7416), .Z(n11880) );
  XNOR2_X1 U13778 ( .A(n11881), .B(n11880), .ZN(n12740) );
  INV_X1 U13779 ( .A(n12740), .ZN(n11746) );
  OAI222_X1 U13780 ( .A1(P2_U3088), .A2(n16213), .B1(n15540), .B2(n11746), 
        .C1(n11743), .C2(n15545), .ZN(P2_U3309) );
  OAI21_X1 U13781 ( .B1(n11744), .B2(P1_IR_REG_17__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n11745) );
  XNOR2_X1 U13782 ( .A(n11745), .B(P1_IR_REG_18__SCAN_IN), .ZN(n15723) );
  INV_X1 U13783 ( .A(n15723), .ZN(n15717) );
  OAI222_X1 U13784 ( .A1(P1_U3086), .A2(n15717), .B1(n11886), .B2(n11746), 
        .C1(n8120), .C2(n16139), .ZN(P1_U3337) );
  AOI21_X1 U13785 ( .B1(n11751), .B2(n11747), .A(n7619), .ZN(n16634) );
  OAI211_X1 U13786 ( .C1(n11748), .C2(n11749), .A(n11908), .B(n16079), .ZN(
        n16630) );
  OAI21_X1 U13787 ( .B1(n11749), .B2(n16725), .A(n16630), .ZN(n11757) );
  OAI211_X1 U13788 ( .C1(n11752), .C2(n11751), .A(n11750), .B(n16561), .ZN(
        n11753) );
  INV_X1 U13789 ( .A(n11753), .ZN(n11755) );
  AOI211_X1 U13790 ( .C1(n16634), .C2(n16472), .A(n11755), .B(n11754), .ZN(
        n16636) );
  INV_X1 U13791 ( .A(n16636), .ZN(n11756) );
  AOI211_X1 U13792 ( .C1(n16660), .C2(n16634), .A(n11757), .B(n11756), .ZN(
        n11903) );
  NAND2_X1 U13793 ( .A1(n16732), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n11758) );
  OAI21_X1 U13794 ( .B1(n11903), .B2(n16732), .A(n11758), .ZN(P1_U3536) );
  NAND2_X1 U13795 ( .A1(n15368), .A2(n15033), .ZN(n11759) );
  NAND2_X1 U13796 ( .A1(n11760), .A2(n11759), .ZN(n12133) );
  NAND2_X1 U13797 ( .A1(n12000), .A2(n12053), .ZN(n11762) );
  AOI22_X1 U13798 ( .A1(n12597), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n12596), 
        .B2(n16232), .ZN(n11761) );
  XNOR2_X1 U13799 ( .A(n16700), .B(n12137), .ZN(n13324) );
  XNOR2_X1 U13800 ( .A(n12133), .B(n8706), .ZN(n16705) );
  NAND2_X1 U13801 ( .A1(n15368), .A2(n13089), .ZN(n11763) );
  NAND2_X1 U13802 ( .A1(n11765), .A2(n13324), .ZN(n11766) );
  NAND3_X1 U13803 ( .A1(n12136), .A2(n15346), .A3(n11766), .ZN(n11775) );
  INV_X1 U13804 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n11767) );
  NAND2_X1 U13805 ( .A1(n11768), .A2(n11767), .ZN(n11769) );
  AND2_X1 U13806 ( .A1(n11803), .A2(n11769), .ZN(n12144) );
  NAND2_X1 U13807 ( .A1(n12144), .A2(n9786), .ZN(n11773) );
  NAND2_X1 U13808 ( .A1(n9790), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n11772) );
  NAND2_X1 U13809 ( .A1(n10847), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n11771) );
  NAND2_X1 U13810 ( .A1(n9789), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n11770) );
  NAND4_X1 U13811 ( .A1(n11773), .A2(n11772), .A3(n11771), .A4(n11770), .ZN(
        n15031) );
  AOI22_X1 U13812 ( .A1(n15341), .A2(n15033), .B1(n15031), .B2(n15343), .ZN(
        n11774) );
  NAND2_X1 U13813 ( .A1(n11775), .A2(n11774), .ZN(n11776) );
  AOI21_X1 U13814 ( .B1(n16705), .B2(n12139), .A(n11776), .ZN(n16707) );
  NAND2_X1 U13815 ( .A1(n11777), .A2(n16700), .ZN(n11778) );
  NAND3_X1 U13816 ( .A1(n12143), .A2(n14960), .A3(n11778), .ZN(n16702) );
  AOI22_X1 U13817 ( .A1(n15362), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n12698), 
        .B2(n15292), .ZN(n11780) );
  NAND2_X1 U13818 ( .A1(n16700), .A2(n15367), .ZN(n11779) );
  OAI211_X1 U13819 ( .C1(n16702), .C2(n15233), .A(n11780), .B(n11779), .ZN(
        n11781) );
  AOI21_X1 U13820 ( .B1(n16705), .B2(n11782), .A(n11781), .ZN(n11783) );
  OAI21_X1 U13821 ( .B1(n16707), .B2(n15362), .A(n11783), .ZN(P2_U3253) );
  NAND2_X1 U13822 ( .A1(n12004), .A2(n12053), .ZN(n11786) );
  AOI22_X1 U13823 ( .A1(n12597), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n12596), 
        .B2(n11784), .ZN(n11785) );
  XNOR2_X1 U13824 ( .A(n13102), .B(n14959), .ZN(n11787) );
  AND2_X1 U13825 ( .A1(n15031), .A2(n14937), .ZN(n11788) );
  NAND2_X1 U13826 ( .A1(n11787), .A2(n11788), .ZN(n12060) );
  INV_X1 U13827 ( .A(n11787), .ZN(n12688) );
  INV_X1 U13828 ( .A(n11788), .ZN(n11789) );
  NAND2_X1 U13829 ( .A1(n12688), .A2(n11789), .ZN(n11790) );
  NAND2_X1 U13830 ( .A1(n12060), .A2(n11790), .ZN(n11798) );
  INV_X1 U13831 ( .A(n11791), .ZN(n12703) );
  XNOR2_X1 U13832 ( .A(n16700), .B(n14959), .ZN(n11793) );
  NAND2_X1 U13833 ( .A1(n15032), .A2(n14937), .ZN(n11794) );
  XNOR2_X1 U13834 ( .A(n11793), .B(n11794), .ZN(n12702) );
  INV_X1 U13835 ( .A(n11793), .ZN(n11795) );
  NAND2_X1 U13836 ( .A1(n11795), .A2(n11794), .ZN(n11796) );
  INV_X1 U13837 ( .A(n12061), .ZN(n12690) );
  AOI211_X1 U13838 ( .C1(n11798), .C2(n11797), .A(n15021), .B(n12690), .ZN(
        n11799) );
  INV_X1 U13839 ( .A(n11799), .ZN(n11812) );
  NAND2_X1 U13840 ( .A1(n10847), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n11801) );
  NAND2_X1 U13841 ( .A1(n9789), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n11800) );
  AND2_X1 U13842 ( .A1(n11801), .A2(n11800), .ZN(n11806) );
  INV_X1 U13843 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n11802) );
  NAND2_X1 U13844 ( .A1(n11803), .A2(n11802), .ZN(n11804) );
  NAND2_X1 U13845 ( .A1(n12067), .A2(n11804), .ZN(n12684) );
  OR2_X1 U13846 ( .A1(n12684), .A2(n13262), .ZN(n11805) );
  OAI211_X1 U13847 ( .C1(n13265), .C2(n11807), .A(n11806), .B(n11805), .ZN(
        n15030) );
  INV_X1 U13848 ( .A(n15030), .ZN(n12468) );
  NAND2_X1 U13849 ( .A1(n15018), .A2(n12144), .ZN(n11808) );
  OAI211_X1 U13850 ( .C1(n14972), .C2(n12468), .A(n11809), .B(n11808), .ZN(
        n11810) );
  AOI21_X1 U13851 ( .B1(n14974), .B2(n15032), .A(n11810), .ZN(n11811) );
  OAI211_X1 U13852 ( .C1(n8319), .C2(n14994), .A(n11812), .B(n11811), .ZN(
        P2_U3206) );
  NAND2_X1 U13853 ( .A1(n16521), .A2(n11813), .ZN(n11814) );
  XOR2_X1 U13854 ( .A(n13527), .B(n11815), .Z(n16520) );
  AOI21_X1 U13855 ( .B1(n11816), .B2(n13527), .A(n14310), .ZN(n11819) );
  OAI22_X1 U13856 ( .A1(n11817), .A2(n14312), .B1(n11925), .B2(n14314), .ZN(
        n11818) );
  AOI21_X1 U13857 ( .B1(n11819), .B2(n11827), .A(n11818), .ZN(n16519) );
  MUX2_X1 U13858 ( .A(n11820), .B(n16519), .S(n14352), .Z(n11822) );
  AOI22_X1 U13859 ( .A1(n14354), .A2(n16524), .B1(n14369), .B2(n14474), .ZN(
        n11821) );
  OAI211_X1 U13860 ( .C1(n14358), .C2(n16520), .A(n11822), .B(n11821), .ZN(
        P3_U3230) );
  XNOR2_X1 U13861 ( .A(n11823), .B(n13377), .ZN(n16546) );
  INV_X1 U13862 ( .A(n11824), .ZN(n11825) );
  NOR2_X1 U13863 ( .A1(n13377), .A2(n11825), .ZN(n11826) );
  AOI21_X1 U13864 ( .B1(n11827), .B2(n11826), .A(n14310), .ZN(n11831) );
  OAI22_X1 U13865 ( .A1(n11829), .A2(n14314), .B1(n11828), .B2(n14312), .ZN(
        n11830) );
  AOI21_X1 U13866 ( .B1(n11832), .B2(n11831), .A(n11830), .ZN(n16547) );
  MUX2_X1 U13867 ( .A(n11833), .B(n16547), .S(n14352), .Z(n11838) );
  INV_X1 U13868 ( .A(n11834), .ZN(n11835) );
  AOI22_X1 U13869 ( .A1(n14354), .A2(n11836), .B1(n14369), .B2(n11835), .ZN(
        n11837) );
  OAI211_X1 U13870 ( .C1(n14358), .C2(n16546), .A(n11838), .B(n11837), .ZN(
        P3_U3229) );
  OAI211_X1 U13871 ( .C1(n11841), .C2(n11840), .A(n11839), .B(n16451), .ZN(
        n11846) );
  OAI22_X1 U13872 ( .A1(n11842), .A2(n13947), .B1(n13978), .B2(n12300), .ZN(
        n11843) );
  AOI211_X1 U13873 ( .C1(n16449), .C2(n16595), .A(n11844), .B(n11843), .ZN(
        n11845) );
  OAI211_X1 U13874 ( .C1(n11945), .C2(n13979), .A(n11846), .B(n11845), .ZN(
        P3_U3153) );
  OR2_X1 U13875 ( .A1(n13715), .A2(n11979), .ZN(n11849) );
  NAND2_X1 U13876 ( .A1(n11850), .A2(n11849), .ZN(n11996) );
  NAND2_X1 U13877 ( .A1(n11851), .A2(n11544), .ZN(n11854) );
  AOI22_X1 U13878 ( .A1(n11852), .A2(n12759), .B1(n12760), .B2(
        P2_DATAO_REG_11__SCAN_IN), .ZN(n11853) );
  NAND2_X1 U13879 ( .A1(n11854), .A2(n11853), .ZN(n13719) );
  XNOR2_X1 U13880 ( .A(n13719), .B(n11997), .ZN(n13587) );
  XNOR2_X1 U13881 ( .A(n11996), .B(n13587), .ZN(n11855) );
  NAND2_X1 U13882 ( .A1(n11855), .A2(n16561), .ZN(n11867) );
  NAND2_X1 U13883 ( .A1(n12945), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n11865) );
  OR2_X1 U13884 ( .A1(n12929), .A2(n10971), .ZN(n11864) );
  INV_X1 U13885 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n11856) );
  OAI21_X1 U13886 ( .B1(n11858), .B2(n11857), .A(n11856), .ZN(n11860) );
  INV_X1 U13887 ( .A(n11859), .ZN(n12011) );
  NAND2_X1 U13888 ( .A1(n11860), .A2(n12011), .ZN(n12400) );
  OR2_X1 U13889 ( .A1(n12946), .A2(n12400), .ZN(n11863) );
  INV_X1 U13890 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n11861) );
  OR2_X1 U13891 ( .A1(n10418), .A2(n11861), .ZN(n11862) );
  NAND4_X1 U13892 ( .A1(n11865), .A2(n11864), .A3(n11863), .A4(n11862), .ZN(
        n15681) );
  AOI22_X1 U13893 ( .A1(n15971), .A2(n15683), .B1(n15681), .B2(n16462), .ZN(
        n11866) );
  NAND2_X1 U13894 ( .A1(n11867), .A2(n11866), .ZN(n16696) );
  INV_X1 U13895 ( .A(n16696), .ZN(n11879) );
  INV_X1 U13896 ( .A(n13587), .ZN(n11995) );
  OR2_X1 U13897 ( .A1(n13715), .A2(n15683), .ZN(n11868) );
  INV_X1 U13898 ( .A(n12019), .ZN(n11870) );
  AOI21_X1 U13899 ( .B1(n11995), .B2(n11871), .A(n11870), .ZN(n16697) );
  OAI21_X1 U13900 ( .B1(n11872), .B2(n16694), .A(n16079), .ZN(n11873) );
  OR2_X1 U13901 ( .A1(n12095), .A2(n11873), .ZN(n16693) );
  NAND2_X1 U13902 ( .A1(n7414), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n11874) );
  OAI21_X1 U13903 ( .B1(n16622), .B2(n11989), .A(n11874), .ZN(n11875) );
  AOI21_X1 U13904 ( .B1(n13719), .B2(n16628), .A(n11875), .ZN(n11876) );
  OAI21_X1 U13905 ( .B1(n16693), .B2(n16631), .A(n11876), .ZN(n11877) );
  AOI21_X1 U13906 ( .B1(n16697), .B2(n15935), .A(n11877), .ZN(n11878) );
  OAI21_X1 U13907 ( .B1(n7414), .B2(n11879), .A(n11878), .ZN(P1_U3282) );
  MUX2_X1 U13908 ( .A(n11887), .B(n11889), .S(n7416), .Z(n11883) );
  INV_X1 U13909 ( .A(n11883), .ZN(n11884) );
  NAND2_X1 U13910 ( .A1(n11884), .A2(SI_19_), .ZN(n11885) );
  NAND2_X1 U13911 ( .A1(n12150), .A2(n11885), .ZN(n12151) );
  INV_X1 U13912 ( .A(n12758), .ZN(n11888) );
  OAI222_X1 U13913 ( .A1(n16139), .A2(n11887), .B1(n11886), .B2(n11888), .C1(
        P1_U3086), .C2(n15733), .ZN(P1_U3336) );
  OAI222_X1 U13914 ( .A1(n15545), .A2(n11889), .B1(n15540), .B2(n11888), .C1(
        n13338), .C2(P2_U3088), .ZN(P2_U3308) );
  AOI21_X1 U13915 ( .B1(n12490), .B2(n11894), .A(n11890), .ZN(n12258) );
  XNOR2_X1 U13916 ( .A(n12258), .B(n11898), .ZN(n11892) );
  INV_X1 U13917 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n11891) );
  NAND2_X1 U13918 ( .A1(n11892), .A2(n11891), .ZN(n12257) );
  OAI21_X1 U13919 ( .B1(n11892), .B2(n11891), .A(n12257), .ZN(n11901) );
  OAI21_X1 U13920 ( .B1(n11894), .B2(n11472), .A(n11893), .ZN(n12263) );
  XOR2_X1 U13921 ( .A(n11898), .B(n12263), .Z(n11895) );
  NOR2_X1 U13922 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n11895), .ZN(n12264) );
  AOI21_X1 U13923 ( .B1(P1_REG2_REG_15__SCAN_IN), .B2(n11895), .A(n12264), 
        .ZN(n11896) );
  NOR2_X1 U13924 ( .A1(n11896), .A2(n15728), .ZN(n11900) );
  NAND2_X1 U13925 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n15668)
         );
  NAND2_X1 U13926 ( .A1(n16246), .A2(P1_ADDR_REG_15__SCAN_IN), .ZN(n11897) );
  OAI211_X1 U13927 ( .C1(n15727), .C2(n11898), .A(n15668), .B(n11897), .ZN(
        n11899) );
  AOI211_X1 U13928 ( .C1(n11901), .C2(n16259), .A(n11900), .B(n11899), .ZN(
        n11902) );
  INV_X1 U13929 ( .A(n11902), .ZN(P1_U3258) );
  INV_X1 U13930 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n11905) );
  OR2_X1 U13931 ( .A1(n11903), .A2(n16735), .ZN(n11904) );
  OAI21_X1 U13932 ( .B1(n16737), .B2(n11905), .A(n11904), .ZN(P1_U3483) );
  OAI21_X1 U13933 ( .B1(n11907), .B2(n13583), .A(n11906), .ZN(n16659) );
  AOI21_X1 U13934 ( .B1(n11908), .B2(n13711), .A(n16464), .ZN(n11910) );
  NAND2_X1 U13935 ( .A1(n11910), .A2(n11909), .ZN(n16655) );
  AOI22_X1 U13936 ( .A1(n16628), .A2(n13711), .B1(n11911), .B2(n15991), .ZN(
        n11912) );
  OAI21_X1 U13937 ( .B1(n16655), .B2(n16631), .A(n11912), .ZN(n11918) );
  XNOR2_X1 U13938 ( .A(n11913), .B(n8620), .ZN(n11916) );
  NAND2_X1 U13939 ( .A1(n16659), .A2(n16472), .ZN(n11915) );
  AOI22_X1 U13940 ( .A1(n15971), .A2(n15685), .B1(n15683), .B2(n16462), .ZN(
        n11914) );
  OAI211_X1 U13941 ( .C1(n16726), .C2(n11916), .A(n11915), .B(n11914), .ZN(
        n16657) );
  MUX2_X1 U13942 ( .A(n16657), .B(P1_REG2_REG_9__SCAN_IN), .S(n7414), .Z(
        n11917) );
  AOI211_X1 U13943 ( .C1(n16633), .C2(n16659), .A(n11918), .B(n11917), .ZN(
        n11919) );
  INV_X1 U13944 ( .A(n11919), .ZN(P1_U3284) );
  XOR2_X1 U13945 ( .A(n13526), .B(n11920), .Z(n16566) );
  NAND2_X1 U13946 ( .A1(n11921), .A2(n13526), .ZN(n11922) );
  NAND2_X1 U13947 ( .A1(n11923), .A2(n11922), .ZN(n11927) );
  NAND2_X1 U13948 ( .A1(n13384), .A2(n16495), .ZN(n11924) );
  OAI21_X1 U13949 ( .B1(n11925), .B2(n14312), .A(n11924), .ZN(n11926) );
  AOI21_X1 U13950 ( .B1(n11927), .B2(n16501), .A(n11926), .ZN(n16564) );
  MUX2_X1 U13951 ( .A(n11928), .B(n16564), .S(n14352), .Z(n11933) );
  INV_X1 U13952 ( .A(n11929), .ZN(n11930) );
  AOI22_X1 U13953 ( .A1(n14354), .A2(n11931), .B1(n14369), .B2(n11930), .ZN(
        n11932) );
  OAI211_X1 U13954 ( .C1(n14358), .C2(n16566), .A(n11933), .B(n11932), .ZN(
        P3_U3228) );
  INV_X1 U13955 ( .A(n11934), .ZN(n11936) );
  OAI222_X1 U13956 ( .A1(n14918), .A2(n11936), .B1(n14920), .B2(n14656), .C1(
        P3_U3151), .C2(n11935), .ZN(P3_U3270) );
  OR2_X1 U13957 ( .A1(n12247), .A2(n13532), .ZN(n12249) );
  NAND2_X1 U13958 ( .A1(n12249), .A2(n11937), .ZN(n11941) );
  OR2_X1 U13959 ( .A1(n12247), .A2(n11938), .ZN(n12236) );
  AND2_X1 U13960 ( .A1(n12236), .A2(n11939), .ZN(n11940) );
  OAI211_X1 U13961 ( .C1(n11941), .C2(n13387), .A(n11940), .B(n16501), .ZN(
        n11943) );
  AOI22_X1 U13962 ( .A1(n13396), .A2(n16495), .B1(n16498), .B2(n13384), .ZN(
        n11942) );
  AND2_X1 U13963 ( .A1(n11943), .A2(n11942), .ZN(n16600) );
  XNOR2_X1 U13964 ( .A(n11944), .B(n13534), .ZN(n16597) );
  NOR2_X1 U13965 ( .A1(n14352), .A2(n9621), .ZN(n11947) );
  OAI22_X1 U13966 ( .A1(n14384), .A2(n13390), .B1(n11945), .B2(n16508), .ZN(
        n11946) );
  AOI211_X1 U13967 ( .C1(n16597), .C2(n14372), .A(n11947), .B(n11946), .ZN(
        n11948) );
  OAI21_X1 U13968 ( .B1(n16600), .B2(n16517), .A(n11948), .ZN(P3_U3226) );
  AOI21_X1 U13969 ( .B1(n11951), .B2(n11950), .A(n11949), .ZN(n11966) );
  OAI21_X1 U13970 ( .B1(n11954), .B2(n11953), .A(n11952), .ZN(n11955) );
  NAND2_X1 U13971 ( .A1(n11955), .A2(n14125), .ZN(n11965) );
  INV_X1 U13972 ( .A(n11956), .ZN(n11957) );
  AOI21_X1 U13973 ( .B1(n11959), .B2(n11958), .A(n11957), .ZN(n11961) );
  INV_X1 U13974 ( .A(P3_REG3_REG_10__SCAN_IN), .ZN(n14699) );
  NOR2_X1 U13975 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n14699), .ZN(n12422) );
  AOI21_X1 U13976 ( .B1(n16150), .B2(P3_ADDR_REG_10__SCAN_IN), .A(n12422), 
        .ZN(n11960) );
  OAI21_X1 U13977 ( .B1(n11961), .B2(n16423), .A(n11960), .ZN(n11962) );
  AOI21_X1 U13978 ( .B1(n11963), .B2(n14146), .A(n11962), .ZN(n11964) );
  OAI211_X1 U13979 ( .C1(n11966), .C2(n16429), .A(n11965), .B(n11964), .ZN(
        P3_U3192) );
  OAI211_X1 U13980 ( .C1(n11969), .C2(n11968), .A(n11967), .B(n16451), .ZN(
        n11974) );
  OAI22_X1 U13981 ( .A1(n12240), .A2(n13947), .B1(n13978), .B2(n12420), .ZN(
        n11970) );
  AOI211_X1 U13982 ( .C1(n16449), .C2(n11972), .A(n11971), .B(n11970), .ZN(
        n11973) );
  OAI211_X1 U13983 ( .C1(n12241), .C2(n13979), .A(n11974), .B(n11973), .ZN(
        P3_U3161) );
  OAI22_X1 U13984 ( .A1(n16694), .A2(n10271), .B1(n11997), .B2(n12846), .ZN(
        n12379) );
  OAI22_X1 U13985 ( .A1(n16694), .A2(n12940), .B1(n11997), .B2(n10271), .ZN(
        n11975) );
  XNOR2_X1 U13986 ( .A(n11975), .B(n10817), .ZN(n12378) );
  XOR2_X1 U13987 ( .A(n12379), .B(n12378), .Z(n11987) );
  NOR2_X1 U13988 ( .A1(n12846), .A2(n11979), .ZN(n11980) );
  AOI21_X1 U13989 ( .B1(n13715), .B2(n7413), .A(n11980), .ZN(n11982) );
  AOI22_X1 U13990 ( .A1(n13715), .A2(n7412), .B1(n7413), .B2(n15683), .ZN(
        n11981) );
  XNOR2_X1 U13991 ( .A(n11981), .B(n10817), .ZN(n11983) );
  XOR2_X1 U13992 ( .A(n11982), .B(n11983), .Z(n12127) );
  INV_X1 U13993 ( .A(n11982), .ZN(n11985) );
  INV_X1 U13994 ( .A(n11983), .ZN(n11984) );
  OAI21_X1 U13995 ( .B1(n11987), .B2(n11986), .A(n12377), .ZN(n11988) );
  NAND2_X1 U13996 ( .A1(n11988), .A2(n16531), .ZN(n11994) );
  NOR2_X1 U13997 ( .A1(n16535), .A2(n11989), .ZN(n11992) );
  INV_X1 U13998 ( .A(n15681), .ZN(n12374) );
  OAI21_X1 U13999 ( .B1(n15648), .B2(n12374), .A(n11990), .ZN(n11991) );
  AOI211_X1 U14000 ( .C1(n15659), .C2(n15683), .A(n11992), .B(n11991), .ZN(
        n11993) );
  OAI211_X1 U14001 ( .C1(n16694), .C2(n15653), .A(n11994), .B(n11993), .ZN(
        P1_U3236) );
  NAND2_X1 U14002 ( .A1(n11996), .A2(n11995), .ZN(n11999) );
  OR2_X1 U14003 ( .A1(n13719), .A2(n11997), .ZN(n11998) );
  NAND2_X1 U14004 ( .A1(n12000), .A2(n11544), .ZN(n12002) );
  AOI22_X1 U14005 ( .A1(n16262), .A2(n12759), .B1(n12760), .B2(
        P2_DATAO_REG_12__SCAN_IN), .ZN(n12001) );
  NAND2_X1 U14006 ( .A1(n12002), .A2(n12001), .ZN(n13728) );
  XNOR2_X1 U14007 ( .A(n13728), .B(n15681), .ZN(n13588) );
  OR2_X1 U14008 ( .A1(n13728), .A2(n12374), .ZN(n12003) );
  NAND2_X1 U14009 ( .A1(n12004), .A2(n11544), .ZN(n12009) );
  NOR2_X1 U14010 ( .A1(n10704), .A2(n12005), .ZN(n12006) );
  AOI21_X1 U14011 ( .B1(n12007), .B2(n12759), .A(n12006), .ZN(n12008) );
  NAND2_X1 U14012 ( .A1(n7420), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n12017) );
  OR2_X1 U14013 ( .A1(n12862), .A2(n16733), .ZN(n12016) );
  NAND2_X1 U14014 ( .A1(n12011), .A2(n12010), .ZN(n12012) );
  NAND2_X1 U14015 ( .A1(n12025), .A2(n12012), .ZN(n12387) );
  OR2_X1 U14016 ( .A1(n12946), .A2(n12387), .ZN(n12015) );
  INV_X1 U14017 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n12013) );
  OR2_X1 U14018 ( .A1(n10418), .A2(n12013), .ZN(n12014) );
  NAND4_X1 U14019 ( .A1(n12017), .A2(n12016), .A3(n12015), .A4(n12014), .ZN(
        n15680) );
  XNOR2_X1 U14020 ( .A(n16722), .B(n15680), .ZN(n13590) );
  XNOR2_X1 U14021 ( .A(n12315), .B(n13590), .ZN(n16727) );
  NAND2_X1 U14022 ( .A1(n13719), .A2(n15682), .ZN(n12018) );
  INV_X1 U14023 ( .A(n13588), .ZN(n12088) );
  INV_X1 U14024 ( .A(n13590), .ZN(n12020) );
  OAI21_X1 U14025 ( .B1(n12021), .B2(n12020), .A(n12324), .ZN(n16731) );
  INV_X1 U14026 ( .A(n13728), .ZN(n12375) );
  AOI21_X1 U14027 ( .B1(n12094), .B2(n16722), .A(n16464), .ZN(n12022) );
  NAND2_X1 U14028 ( .A1(n12022), .A2(n12327), .ZN(n16724) );
  NOR2_X1 U14029 ( .A1(n16625), .A2(n12023), .ZN(n12034) );
  NAND2_X1 U14030 ( .A1(n13566), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n12030) );
  OR2_X1 U14031 ( .A1(n12929), .A2(n11472), .ZN(n12029) );
  NAND2_X1 U14032 ( .A1(n12025), .A2(n12024), .ZN(n12026) );
  NAND2_X1 U14033 ( .A1(n12308), .A2(n12026), .ZN(n12534) );
  OR2_X1 U14034 ( .A1(n12946), .A2(n12534), .ZN(n12028) );
  OR2_X1 U14035 ( .A1(n12862), .A2(n12490), .ZN(n12027) );
  NAND4_X1 U14036 ( .A1(n12030), .A2(n12029), .A3(n12028), .A4(n12027), .ZN(
        n15679) );
  NAND2_X1 U14037 ( .A1(n15679), .A2(n16462), .ZN(n12032) );
  NAND2_X1 U14038 ( .A1(n15681), .A2(n15971), .ZN(n12031) );
  NAND2_X1 U14039 ( .A1(n12032), .A2(n12031), .ZN(n12385) );
  INV_X1 U14040 ( .A(n12385), .ZN(n16723) );
  OAI22_X1 U14041 ( .A1(n7414), .A2(n16723), .B1(n12387), .B2(n16622), .ZN(
        n12033) );
  AOI211_X1 U14042 ( .C1(n16722), .C2(n16628), .A(n12034), .B(n12033), .ZN(
        n12035) );
  OAI21_X1 U14043 ( .B1(n16724), .B2(n16631), .A(n12035), .ZN(n12036) );
  AOI21_X1 U14044 ( .B1(n16731), .B2(n15935), .A(n12036), .ZN(n12037) );
  OAI21_X1 U14045 ( .B1(n15947), .B2(n16727), .A(n12037), .ZN(P1_U3280) );
  AND2_X1 U14046 ( .A1(n12039), .A2(n12038), .ZN(n12284) );
  NAND2_X1 U14047 ( .A1(n12284), .A2(n16501), .ZN(n12044) );
  NAND2_X1 U14048 ( .A1(n12236), .A2(n12040), .ZN(n12237) );
  AOI21_X1 U14049 ( .B1(n12237), .B2(n12041), .A(n13395), .ZN(n12043) );
  AOI22_X1 U14050 ( .A1(n13396), .A2(n16498), .B1(n16495), .B2(n13406), .ZN(
        n12042) );
  OAI21_X1 U14051 ( .B1(n12044), .B2(n12043), .A(n12042), .ZN(n16649) );
  INV_X1 U14052 ( .A(n16649), .ZN(n12052) );
  OAI22_X1 U14053 ( .A1(n14384), .A2(n12045), .B1(n12302), .B2(n16508), .ZN(
        n12048) );
  NOR2_X1 U14054 ( .A1(n14352), .A2(n12046), .ZN(n12047) );
  NOR2_X1 U14055 ( .A1(n12048), .A2(n12047), .ZN(n12051) );
  NAND2_X1 U14056 ( .A1(n12049), .A2(n13395), .ZN(n16646) );
  NAND3_X1 U14057 ( .A1(n16648), .A2(n16646), .A3(n14372), .ZN(n12050) );
  OAI211_X1 U14058 ( .C1(n12052), .C2(n16517), .A(n12051), .B(n12050), .ZN(
        P3_U3224) );
  NAND2_X1 U14059 ( .A1(n12338), .A2(n12053), .ZN(n12056) );
  AOI22_X1 U14060 ( .A1(n12054), .A2(n12596), .B1(n12597), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n12055) );
  NAND2_X1 U14061 ( .A1(n12318), .A2(n12053), .ZN(n12059) );
  AOI22_X1 U14062 ( .A1(n12596), .A2(n12057), .B1(n12597), .B2(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n12058) );
  XNOR2_X1 U14063 ( .A(n16741), .B(n14959), .ZN(n12062) );
  NAND2_X1 U14064 ( .A1(n15030), .A2(n14937), .ZN(n12063) );
  XNOR2_X1 U14065 ( .A(n12062), .B(n12063), .ZN(n12691) );
  NAND3_X1 U14066 ( .A1(n12061), .A2(n12691), .A3(n12060), .ZN(n12696) );
  INV_X1 U14067 ( .A(n12062), .ZN(n12064) );
  NAND2_X1 U14068 ( .A1(n12064), .A2(n12063), .ZN(n12065) );
  XNOR2_X1 U14069 ( .A(n13113), .B(n14936), .ZN(n12173) );
  NAND2_X1 U14070 ( .A1(n12067), .A2(n12066), .ZN(n12068) );
  NAND2_X1 U14071 ( .A1(n12079), .A2(n12068), .ZN(n12475) );
  AOI22_X1 U14072 ( .A1(n9790), .A2(P2_REG1_REG_15__SCAN_IN), .B1(n10847), 
        .B2(P2_REG0_REG_15__SCAN_IN), .ZN(n12070) );
  NAND2_X1 U14073 ( .A1(n9789), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n12069) );
  OAI211_X1 U14074 ( .C1(n12475), .C2(n13262), .A(n12070), .B(n12069), .ZN(
        n15029) );
  AND2_X1 U14075 ( .A1(n15029), .A2(n14937), .ZN(n12071) );
  NAND2_X1 U14076 ( .A1(n12173), .A2(n12071), .ZN(n12172) );
  INV_X1 U14077 ( .A(n12173), .ZN(n12073) );
  INV_X1 U14078 ( .A(n12071), .ZN(n12072) );
  NAND2_X1 U14079 ( .A1(n12073), .A2(n12072), .ZN(n12074) );
  AND2_X1 U14080 ( .A1(n12172), .A2(n12074), .ZN(n12075) );
  OAI211_X1 U14081 ( .C1(n12076), .C2(n12075), .A(n12175), .B(n15000), .ZN(
        n12086) );
  OAI21_X1 U14082 ( .B1(n15003), .B2(n12475), .A(n12077), .ZN(n12084) );
  INV_X1 U14083 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n12078) );
  NAND2_X1 U14084 ( .A1(n12079), .A2(n12078), .ZN(n12080) );
  NAND2_X1 U14085 ( .A1(n12179), .A2(n12080), .ZN(n12503) );
  OR2_X1 U14086 ( .A1(n12503), .A2(n13262), .ZN(n12082) );
  AOI22_X1 U14087 ( .A1(n9790), .A2(P2_REG1_REG_16__SCAN_IN), .B1(n10847), 
        .B2(P2_REG0_REG_16__SCAN_IN), .ZN(n12081) );
  OAI211_X1 U14088 ( .C1(n10470), .C2(n11492), .A(n12082), .B(n12081), .ZN(
        n15028) );
  INV_X1 U14089 ( .A(n15028), .ZN(n13120) );
  NOR2_X1 U14090 ( .A1(n14972), .A2(n13120), .ZN(n12083) );
  AOI211_X1 U14091 ( .C1(n14974), .C2(n15030), .A(n12084), .B(n12083), .ZN(
        n12085) );
  OAI211_X1 U14092 ( .C1(n15518), .C2(n14994), .A(n12086), .B(n12085), .ZN(
        P2_U3213) );
  OAI21_X1 U14093 ( .B1(n12089), .B2(n12088), .A(n12087), .ZN(n12272) );
  INV_X1 U14094 ( .A(n12272), .ZN(n12100) );
  XNOR2_X1 U14095 ( .A(n12090), .B(n13588), .ZN(n12093) );
  NAND2_X1 U14096 ( .A1(n12272), .A2(n16472), .ZN(n12092) );
  AOI22_X1 U14097 ( .A1(n15971), .A2(n15682), .B1(n15680), .B2(n16462), .ZN(
        n12091) );
  OAI211_X1 U14098 ( .C1(n16726), .C2(n12093), .A(n12092), .B(n12091), .ZN(
        n12276) );
  NAND2_X1 U14099 ( .A1(n12276), .A2(n16625), .ZN(n12099) );
  OAI22_X1 U14100 ( .A1(n16625), .A2(n10971), .B1(n12400), .B2(n16622), .ZN(
        n12097) );
  OAI211_X1 U14101 ( .C1(n12095), .C2(n12375), .A(n16079), .B(n12094), .ZN(
        n12273) );
  NOR2_X1 U14102 ( .A1(n12273), .A2(n16631), .ZN(n12096) );
  AOI211_X1 U14103 ( .C1(n16628), .C2(n13728), .A(n12097), .B(n12096), .ZN(
        n12098) );
  OAI211_X1 U14104 ( .C1(n12100), .C2(n15826), .A(n12099), .B(n12098), .ZN(
        P1_U3281) );
  AND2_X1 U14105 ( .A1(n12194), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n12101) );
  AOI21_X1 U14106 ( .B1(n12103), .B2(n12102), .A(n12101), .ZN(n12104) );
  XNOR2_X1 U14107 ( .A(n12104), .B(n12438), .ZN(n16216) );
  INV_X1 U14108 ( .A(n12104), .ZN(n12105) );
  AOI22_X1 U14109 ( .A1(n16216), .A2(P2_REG1_REG_18__SCAN_IN), .B1(n12438), 
        .B2(n12105), .ZN(n12107) );
  XNOR2_X1 U14110 ( .A(n13341), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n12106) );
  XNOR2_X1 U14111 ( .A(n12107), .B(n12106), .ZN(n12121) );
  OAI21_X1 U14112 ( .B1(n12109), .B2(n11490), .A(n12108), .ZN(n12110) );
  NOR2_X1 U14113 ( .A1(n12110), .A2(n12438), .ZN(n12112) );
  AOI21_X1 U14114 ( .B1(n12438), .B2(n12110), .A(n12112), .ZN(n12111) );
  INV_X1 U14115 ( .A(n12111), .ZN(n16211) );
  NOR2_X1 U14116 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n16211), .ZN(n16210) );
  NOR2_X1 U14117 ( .A1(n12112), .A2(n16210), .ZN(n12115) );
  INV_X1 U14118 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n12113) );
  MUX2_X1 U14119 ( .A(n12113), .B(P2_REG2_REG_19__SCAN_IN), .S(n13341), .Z(
        n12114) );
  XNOR2_X1 U14120 ( .A(n12115), .B(n12114), .ZN(n12119) );
  NAND2_X1 U14121 ( .A1(n10096), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n12117) );
  NAND2_X1 U14122 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n12607)
         );
  NAND2_X1 U14123 ( .A1(n16231), .A2(n13341), .ZN(n12116) );
  NAND3_X1 U14124 ( .A1(n12117), .A2(n12607), .A3(n12116), .ZN(n12118) );
  AOI21_X1 U14125 ( .B1(n12119), .B2(n16229), .A(n12118), .ZN(n12120) );
  OAI21_X1 U14126 ( .B1(n12121), .B2(n16190), .A(n12120), .ZN(P2_U3233) );
  NAND2_X1 U14127 ( .A1(n15659), .A2(n15684), .ZN(n12126) );
  NAND2_X1 U14128 ( .A1(n15658), .A2(n15682), .ZN(n12125) );
  OR2_X1 U14129 ( .A1(n16535), .A2(n12122), .ZN(n12123) );
  NAND4_X1 U14130 ( .A1(n12126), .A2(n12125), .A3(n12124), .A4(n12123), .ZN(
        n12131) );
  XNOR2_X1 U14131 ( .A(n12128), .B(n12127), .ZN(n12129) );
  NOR2_X1 U14132 ( .A1(n12129), .A2(n15673), .ZN(n12130) );
  AOI211_X1 U14133 ( .C1(n15671), .C2(n13715), .A(n12131), .B(n12130), .ZN(
        n12132) );
  INV_X1 U14134 ( .A(n12132), .ZN(P1_U3217) );
  NAND2_X1 U14135 ( .A1(n16700), .A2(n15032), .ZN(n12134) );
  XNOR2_X1 U14136 ( .A(n13102), .B(n12697), .ZN(n13325) );
  INV_X1 U14137 ( .A(n13325), .ZN(n12216) );
  OAI21_X1 U14138 ( .B1(n7602), .B2(n13325), .A(n12224), .ZN(n12409) );
  INV_X1 U14139 ( .A(n12409), .ZN(n12149) );
  OR2_X1 U14140 ( .A1(n16700), .A2(n12137), .ZN(n12135) );
  XNOR2_X1 U14141 ( .A(n12217), .B(n12216), .ZN(n12141) );
  OAI22_X1 U14142 ( .A1(n12468), .A2(n15287), .B1(n12137), .B2(n15289), .ZN(
        n12138) );
  AOI21_X1 U14143 ( .B1(n12409), .B2(n12139), .A(n12138), .ZN(n12140) );
  OAI21_X1 U14144 ( .B1(n15308), .B2(n12141), .A(n12140), .ZN(n12407) );
  NAND2_X1 U14145 ( .A1(n12407), .A2(n15353), .ZN(n12148) );
  INV_X1 U14146 ( .A(n12226), .ZN(n12142) );
  AOI211_X1 U14147 ( .C1(n13102), .C2(n12143), .A(n14937), .B(n12142), .ZN(
        n12408) );
  AOI22_X1 U14148 ( .A1(n15362), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n12144), 
        .B2(n15292), .ZN(n12145) );
  OAI21_X1 U14149 ( .B1(n8319), .B2(n15330), .A(n12145), .ZN(n12146) );
  AOI21_X1 U14150 ( .B1(n12408), .B2(n15371), .A(n12146), .ZN(n12147) );
  OAI211_X1 U14151 ( .C1(n12149), .C2(n15336), .A(n12148), .B(n12147), .ZN(
        P2_U3252) );
  MUX2_X1 U14152 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(P1_DATAO_REG_20__SCAN_IN), 
        .S(n7416), .Z(n12367) );
  XNOR2_X1 U14153 ( .A(n12367), .B(n14664), .ZN(n12153) );
  INV_X1 U14154 ( .A(n12969), .ZN(n12295) );
  OAI222_X1 U14155 ( .A1(n16139), .A2(n12779), .B1(n11886), .B2(n12295), .C1(
        n13610), .C2(P1_U3086), .ZN(P1_U3335) );
  AOI21_X1 U14156 ( .B1(n12155), .B2(n16690), .A(n12154), .ZN(n12169) );
  OAI21_X1 U14157 ( .B1(n12158), .B2(n12157), .A(n12156), .ZN(n12159) );
  NAND2_X1 U14158 ( .A1(n12159), .A2(n14125), .ZN(n12168) );
  AOI21_X1 U14159 ( .B1(n12161), .B2(n9125), .A(n12160), .ZN(n12164) );
  INV_X1 U14160 ( .A(P3_REG3_REG_11__SCAN_IN), .ZN(n14719) );
  NOR2_X1 U14161 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n14719), .ZN(n12579) );
  INV_X1 U14162 ( .A(n12579), .ZN(n12163) );
  NAND2_X1 U14163 ( .A1(n16150), .A2(P3_ADDR_REG_11__SCAN_IN), .ZN(n12162) );
  OAI211_X1 U14164 ( .C1(n16423), .C2(n12164), .A(n12163), .B(n12162), .ZN(
        n12165) );
  AOI21_X1 U14165 ( .B1(n12166), .B2(n14146), .A(n12165), .ZN(n12167) );
  OAI211_X1 U14166 ( .C1(n12169), .C2(n16429), .A(n12168), .B(n12167), .ZN(
        P3_U3193) );
  AOI22_X1 U14167 ( .A1(n12597), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n12596), 
        .B2(n12170), .ZN(n12171) );
  XNOR2_X1 U14168 ( .A(n15511), .B(n14929), .ZN(n12210) );
  NAND2_X1 U14169 ( .A1(n15028), .A2(n14937), .ZN(n12192) );
  XNOR2_X1 U14170 ( .A(n12210), .B(n12192), .ZN(n12176) );
  NAND3_X1 U14171 ( .A1(n12173), .A2(n14961), .A3(n15029), .ZN(n12174) );
  OAI21_X1 U14172 ( .B1(n12175), .B2(n15021), .A(n12174), .ZN(n12177) );
  NAND2_X1 U14173 ( .A1(n12177), .A2(n12176), .ZN(n12191) );
  NAND2_X1 U14174 ( .A1(n12179), .A2(n12178), .ZN(n12180) );
  AND2_X1 U14175 ( .A1(n12198), .A2(n12180), .ZN(n12590) );
  NAND2_X1 U14176 ( .A1(n12590), .A2(n9786), .ZN(n12185) );
  NAND2_X1 U14177 ( .A1(n9789), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n12182) );
  NAND2_X1 U14178 ( .A1(n9788), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n12181) );
  OAI211_X1 U14179 ( .C1(n13265), .C2(n15451), .A(n12182), .B(n12181), .ZN(
        n12183) );
  INV_X1 U14180 ( .A(n12183), .ZN(n12184) );
  NAND2_X1 U14181 ( .A1(n12185), .A2(n12184), .ZN(n15342) );
  NAND2_X1 U14182 ( .A1(n15342), .A2(n15343), .ZN(n12187) );
  NAND2_X1 U14183 ( .A1(n15029), .A2(n15341), .ZN(n12186) );
  NAND2_X1 U14184 ( .A1(n12187), .A2(n12186), .ZN(n12494) );
  NAND2_X1 U14185 ( .A1(n14991), .A2(n12494), .ZN(n12188) );
  NAND2_X1 U14186 ( .A1(P2_U3088), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n16198)
         );
  OAI211_X1 U14187 ( .C1(n15003), .C2(n12503), .A(n12188), .B(n16198), .ZN(
        n12189) );
  AOI21_X1 U14188 ( .B1(n15511), .B2(n15024), .A(n12189), .ZN(n12190) );
  OAI211_X1 U14189 ( .C1(n12212), .C2(n15021), .A(n12191), .B(n12190), .ZN(
        P2_U3198) );
  NAND2_X1 U14190 ( .A1(n12210), .A2(n12192), .ZN(n12193) );
  NAND2_X1 U14191 ( .A1(n12212), .A2(n12193), .ZN(n12196) );
  AOI22_X1 U14192 ( .A1(n12597), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n12596), 
        .B2(n12194), .ZN(n12195) );
  XNOR2_X1 U14193 ( .A(n15146), .B(n14959), .ZN(n12445) );
  NAND2_X1 U14194 ( .A1(n15342), .A2(n14937), .ZN(n12446) );
  XNOR2_X1 U14195 ( .A(n12445), .B(n12446), .ZN(n12209) );
  INV_X1 U14196 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n12197) );
  NAND2_X1 U14197 ( .A1(n12198), .A2(n12197), .ZN(n12199) );
  NAND2_X1 U14198 ( .A1(n12454), .A2(n12199), .ZN(n15351) );
  OR2_X1 U14199 ( .A1(n15351), .A2(n13262), .ZN(n12204) );
  INV_X1 U14200 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n15352) );
  NAND2_X1 U14201 ( .A1(n9790), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n12201) );
  NAND2_X1 U14202 ( .A1(n10847), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n12200) );
  OAI211_X1 U14203 ( .C1(n15352), .C2(n10470), .A(n12201), .B(n12200), .ZN(
        n12202) );
  INV_X1 U14204 ( .A(n12202), .ZN(n12203) );
  NAND2_X1 U14205 ( .A1(n12204), .A2(n12203), .ZN(n15319) );
  INV_X1 U14206 ( .A(n15319), .ZN(n15150) );
  NOR2_X1 U14207 ( .A1(n14972), .A2(n15150), .ZN(n12208) );
  NAND2_X1 U14208 ( .A1(n15018), .A2(n12590), .ZN(n12205) );
  OAI211_X1 U14209 ( .C1(n12994), .C2(n13120), .A(n12206), .B(n12205), .ZN(
        n12207) );
  AOI211_X1 U14210 ( .C1(n8008), .C2(n15024), .A(n12208), .B(n12207), .ZN(
        n12215) );
  INV_X1 U14211 ( .A(n12209), .ZN(n12213) );
  OAI22_X1 U14212 ( .A1(n12210), .A2(n15021), .B1(n13120), .B2(n15011), .ZN(
        n12211) );
  NAND3_X1 U14213 ( .A1(n12213), .A2(n12212), .A3(n12211), .ZN(n12214) );
  OAI211_X1 U14214 ( .C1(n12449), .C2(n15021), .A(n12215), .B(n12214), .ZN(
        P2_U3200) );
  XNOR2_X1 U14215 ( .A(n16741), .B(n12468), .ZN(n13327) );
  NAND2_X1 U14216 ( .A1(n12218), .A2(n13327), .ZN(n12219) );
  NAND2_X1 U14217 ( .A1(n12470), .A2(n12219), .ZN(n12222) );
  NAND2_X1 U14218 ( .A1(n15029), .A2(n15343), .ZN(n12220) );
  OAI21_X1 U14219 ( .B1(n12697), .B2(n15289), .A(n12220), .ZN(n12221) );
  AOI21_X1 U14220 ( .B1(n12222), .B2(n15346), .A(n12221), .ZN(n16744) );
  OR2_X1 U14221 ( .A1(n13102), .A2(n15031), .ZN(n12223) );
  OAI21_X1 U14222 ( .B1(n12225), .B2(n13327), .A(n12466), .ZN(n16739) );
  INV_X1 U14223 ( .A(n16739), .ZN(n12231) );
  AOI21_X1 U14224 ( .B1(n16741), .B2(n12226), .A(n14937), .ZN(n12227) );
  NAND2_X1 U14225 ( .A1(n12227), .A2(n12474), .ZN(n16743) );
  OAI22_X1 U14226 ( .A1(n15327), .A2(n10797), .B1(n12684), .B2(n15364), .ZN(
        n12228) );
  AOI21_X1 U14227 ( .B1(n16741), .B2(n15367), .A(n12228), .ZN(n12229) );
  OAI21_X1 U14228 ( .B1(n16743), .B2(n15233), .A(n12229), .ZN(n12230) );
  AOI21_X1 U14229 ( .B1(n12231), .B2(n15369), .A(n12230), .ZN(n12232) );
  OAI21_X1 U14230 ( .B1(n15362), .B2(n16744), .A(n12232), .ZN(P2_U3251) );
  XNOR2_X1 U14231 ( .A(n12234), .B(n12233), .ZN(n16616) );
  INV_X1 U14232 ( .A(n12237), .ZN(n12238) );
  AOI21_X1 U14233 ( .B1(n13524), .B2(n7604), .A(n12238), .ZN(n12239) );
  OAI222_X1 U14234 ( .A1(n14314), .A2(n12420), .B1(n14312), .B2(n12240), .C1(
        n14310), .C2(n12239), .ZN(n16617) );
  NAND2_X1 U14235 ( .A1(n16617), .A2(n14352), .ZN(n12244) );
  OAI22_X1 U14236 ( .A1(n14384), .A2(n16614), .B1(n12241), .B2(n16508), .ZN(
        n12242) );
  AOI21_X1 U14237 ( .B1(P3_REG2_REG_8__SCAN_IN), .B2(n16517), .A(n12242), .ZN(
        n12243) );
  OAI211_X1 U14238 ( .C1(n14358), .C2(n16616), .A(n12244), .B(n12243), .ZN(
        P3_U3225) );
  XNOR2_X1 U14239 ( .A(n12245), .B(n13532), .ZN(n16579) );
  INV_X1 U14240 ( .A(n16580), .ZN(n13383) );
  OAI22_X1 U14241 ( .A1(n14384), .A2(n13383), .B1(n12246), .B2(n16508), .ZN(
        n12254) );
  NAND2_X1 U14242 ( .A1(n12247), .A2(n13532), .ZN(n12248) );
  NAND3_X1 U14243 ( .A1(n12249), .A2(n16501), .A3(n12248), .ZN(n12252) );
  AOI22_X1 U14244 ( .A1(n12250), .A2(n16498), .B1(n16495), .B2(n13391), .ZN(
        n12251) );
  NAND2_X1 U14245 ( .A1(n12252), .A2(n12251), .ZN(n16578) );
  MUX2_X1 U14246 ( .A(n16578), .B(P3_REG2_REG_6__SCAN_IN), .S(n16517), .Z(
        n12253) );
  AOI211_X1 U14247 ( .C1(n14372), .C2(n16579), .A(n12254), .B(n12253), .ZN(
        n12255) );
  INV_X1 U14248 ( .A(n12255), .ZN(P3_U3227) );
  INV_X1 U14249 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n12256) );
  NAND2_X1 U14250 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n15596)
         );
  OAI21_X1 U14251 ( .B1(n16267), .B2(n12256), .A(n15596), .ZN(n12262) );
  OAI21_X1 U14252 ( .B1(n12258), .B2(n12339), .A(n12257), .ZN(n12260) );
  XNOR2_X1 U14253 ( .A(n12540), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n12259) );
  NOR2_X1 U14254 ( .A1(n12259), .A2(n12260), .ZN(n12431) );
  AOI211_X1 U14255 ( .C1(n12260), .C2(n12259), .A(n12431), .B(n15710), .ZN(
        n12261) );
  AOI211_X1 U14256 ( .C1(n16261), .C2(n12540), .A(n12262), .B(n12261), .ZN(
        n12271) );
  NOR2_X1 U14257 ( .A1(n12339), .A2(n12263), .ZN(n12265) );
  NOR2_X1 U14258 ( .A1(n12265), .A2(n12264), .ZN(n12269) );
  INV_X1 U14259 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n12266) );
  MUX2_X1 U14260 ( .A(n12266), .B(P1_REG2_REG_16__SCAN_IN), .S(n12540), .Z(
        n12267) );
  INV_X1 U14261 ( .A(n12267), .ZN(n12268) );
  NAND2_X1 U14262 ( .A1(n12268), .A2(n12269), .ZN(n12427) );
  OAI211_X1 U14263 ( .C1(n12269), .C2(n12268), .A(n16263), .B(n12427), .ZN(
        n12270) );
  NAND2_X1 U14264 ( .A1(n12271), .A2(n12270), .ZN(P1_U3259) );
  NAND2_X1 U14265 ( .A1(n12272), .A2(n16660), .ZN(n12274) );
  OAI211_X1 U14266 ( .C1(n12375), .C2(n16725), .A(n12274), .B(n12273), .ZN(
        n12275) );
  NOR2_X1 U14267 ( .A1(n12276), .A2(n12275), .ZN(n12278) );
  MUX2_X1 U14268 ( .A(n10966), .B(n12278), .S(n16734), .Z(n12277) );
  INV_X1 U14269 ( .A(n12277), .ZN(P1_U3540) );
  MUX2_X1 U14270 ( .A(n11861), .B(n12278), .S(n16737), .Z(n12279) );
  INV_X1 U14271 ( .A(n12279), .ZN(P1_U3495) );
  AOI21_X1 U14272 ( .B1(n12282), .B2(n12280), .A(n7618), .ZN(n16664) );
  OAI22_X1 U14273 ( .A1(n14384), .A2(n16663), .B1(n12426), .B2(n16508), .ZN(
        n12281) );
  AOI21_X1 U14274 ( .B1(P3_REG2_REG_10__SCAN_IN), .B2(n16517), .A(n12281), 
        .ZN(n12291) );
  INV_X1 U14275 ( .A(n12282), .ZN(n13538) );
  NAND3_X1 U14276 ( .A1(n12284), .A2(n13538), .A3(n12283), .ZN(n12285) );
  NAND3_X1 U14277 ( .A1(n12286), .A2(n16501), .A3(n12285), .ZN(n12289) );
  AOI22_X1 U14278 ( .A1(n16498), .A2(n12287), .B1(n14380), .B2(n16495), .ZN(
        n12288) );
  NAND2_X1 U14279 ( .A1(n12289), .A2(n12288), .ZN(n16665) );
  NAND2_X1 U14280 ( .A1(n16665), .A2(n14352), .ZN(n12290) );
  OAI211_X1 U14281 ( .C1(n16664), .C2(n14358), .A(n12291), .B(n12290), .ZN(
        P3_U3223) );
  INV_X1 U14282 ( .A(n12292), .ZN(n12293) );
  OAI222_X1 U14283 ( .A1(P3_U3151), .A2(n12294), .B1(n14920), .B2(n14483), 
        .C1(n14918), .C2(n12293), .ZN(P3_U3269) );
  OAI222_X1 U14284 ( .A1(n15545), .A2(n12970), .B1(P2_U3088), .B2(n13345), 
        .C1(n15540), .C2(n12295), .ZN(P2_U3307) );
  INV_X1 U14285 ( .A(n12296), .ZN(n12297) );
  AOI21_X1 U14286 ( .B1(n12299), .B2(n12298), .A(n12297), .ZN(n12306) );
  NOR2_X1 U14287 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n8863), .ZN(n16435) );
  OAI22_X1 U14288 ( .A1(n12300), .A2(n13947), .B1(n13978), .B2(n12577), .ZN(
        n12301) );
  AOI211_X1 U14289 ( .C1(n16449), .C2(n16651), .A(n16435), .B(n12301), .ZN(
        n12305) );
  INV_X1 U14290 ( .A(n12302), .ZN(n12303) );
  NAND2_X1 U14291 ( .A1(n13970), .A2(n12303), .ZN(n12304) );
  OAI211_X1 U14292 ( .C1(n12306), .C2(n13954), .A(n12305), .B(n12304), .ZN(
        P3_U3171) );
  NAND2_X1 U14293 ( .A1(n12945), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n12314) );
  INV_X1 U14294 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n12361) );
  OR2_X1 U14295 ( .A1(n12929), .A2(n12361), .ZN(n12313) );
  NAND2_X1 U14296 ( .A1(n12308), .A2(n12307), .ZN(n12309) );
  NAND2_X1 U14297 ( .A1(n12351), .A2(n12309), .ZN(n15669) );
  OR2_X1 U14298 ( .A1(n12946), .A2(n15669), .ZN(n12312) );
  INV_X1 U14299 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n12310) );
  OR2_X1 U14300 ( .A1(n10418), .A2(n12310), .ZN(n12311) );
  NAND4_X1 U14301 ( .A1(n12314), .A2(n12313), .A3(n12312), .A4(n12311), .ZN(
        n15678) );
  INV_X1 U14302 ( .A(n15680), .ZN(n12397) );
  OR2_X1 U14303 ( .A1(n16722), .A2(n12397), .ZN(n12316) );
  NAND2_X1 U14304 ( .A1(n12318), .A2(n11544), .ZN(n12321) );
  AOI22_X1 U14305 ( .A1(n12319), .A2(n12759), .B1(n12760), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n12320) );
  XNOR2_X1 U14306 ( .A(n13736), .B(n15679), .ZN(n13593) );
  XNOR2_X1 U14307 ( .A(n12345), .B(n13593), .ZN(n12322) );
  OAI222_X1 U14308 ( .A1(n15953), .A2(n12713), .B1(n15951), .B2(n12397), .C1(
        n12322), .C2(n16726), .ZN(n12485) );
  INV_X1 U14309 ( .A(n12485), .ZN(n12335) );
  OR2_X1 U14310 ( .A1(n16722), .A2(n15680), .ZN(n12323) );
  INV_X1 U14311 ( .A(n12337), .ZN(n12325) );
  AOI21_X1 U14312 ( .B1(n13593), .B2(n12326), .A(n12325), .ZN(n12486) );
  AND2_X1 U14313 ( .A1(n13736), .A2(n12327), .ZN(n12328) );
  OR2_X1 U14314 ( .A1(n12347), .A2(n12328), .ZN(n12483) );
  NOR2_X1 U14315 ( .A1(n7414), .A2(n12329), .ZN(n15986) );
  INV_X1 U14316 ( .A(n15986), .ZN(n12364) );
  NAND2_X1 U14317 ( .A1(n7414), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n12330) );
  OAI21_X1 U14318 ( .B1(n16622), .B2(n12534), .A(n12330), .ZN(n12331) );
  AOI21_X1 U14319 ( .B1(n13736), .B2(n16628), .A(n12331), .ZN(n12332) );
  OAI21_X1 U14320 ( .B1(n12483), .B2(n12364), .A(n12332), .ZN(n12333) );
  AOI21_X1 U14321 ( .B1(n12486), .B2(n15935), .A(n12333), .ZN(n12334) );
  OAI21_X1 U14322 ( .B1(n7414), .B2(n12335), .A(n12334), .ZN(P1_U3279) );
  NAND2_X1 U14323 ( .A1(n13736), .A2(n15679), .ZN(n12336) );
  NAND2_X1 U14324 ( .A1(n12338), .A2(n11544), .ZN(n12341) );
  AOI22_X1 U14325 ( .A1(n12339), .A2(n12759), .B1(n12760), .B2(
        P2_DATAO_REG_15__SCAN_IN), .ZN(n12340) );
  NAND2_X1 U14326 ( .A1(n16090), .A2(n12713), .ZN(n12342) );
  NAND2_X1 U14327 ( .A1(n12538), .A2(n12342), .ZN(n13592) );
  XNOR2_X1 U14328 ( .A(n12555), .B(n13592), .ZN(n16096) );
  INV_X1 U14329 ( .A(n13593), .ZN(n12344) );
  INV_X1 U14330 ( .A(n15679), .ZN(n12520) );
  NAND2_X1 U14331 ( .A1(n13736), .A2(n12520), .ZN(n12343) );
  AOI21_X1 U14332 ( .B1(n13592), .B2(n12346), .A(n7607), .ZN(n16094) );
  NAND2_X1 U14333 ( .A1(n8605), .A2(n12347), .ZN(n12561) );
  OR2_X1 U14334 ( .A1(n8605), .A2(n12347), .ZN(n12348) );
  NAND2_X1 U14335 ( .A1(n12561), .A2(n12348), .ZN(n16092) );
  INV_X1 U14336 ( .A(n12349), .ZN(n12545) );
  NAND2_X1 U14337 ( .A1(n12351), .A2(n12350), .ZN(n12352) );
  NAND2_X1 U14338 ( .A1(n12545), .A2(n12352), .ZN(n15599) );
  OR2_X1 U14339 ( .A1(n12946), .A2(n15599), .ZN(n12358) );
  INV_X1 U14340 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n12353) );
  OR2_X1 U14341 ( .A1(n12862), .A2(n12353), .ZN(n12357) );
  OR2_X1 U14342 ( .A1(n12929), .A2(n12266), .ZN(n12356) );
  INV_X1 U14343 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n12354) );
  OR2_X1 U14344 ( .A1(n10418), .A2(n12354), .ZN(n12355) );
  NAND4_X1 U14345 ( .A1(n12358), .A2(n12357), .A3(n12356), .A4(n12355), .ZN(
        n15972) );
  INV_X1 U14346 ( .A(n15972), .ZN(n12722) );
  OAI22_X1 U14347 ( .A1(n12520), .A2(n15951), .B1(n12722), .B2(n15953), .ZN(
        n16089) );
  NOR2_X1 U14348 ( .A1(n15669), .A2(n16622), .ZN(n12359) );
  AOI21_X1 U14349 ( .B1(n16625), .B2(n16089), .A(n12359), .ZN(n12360) );
  OAI21_X1 U14350 ( .B1(n12361), .B2(n16625), .A(n12360), .ZN(n12362) );
  AOI21_X1 U14351 ( .B1(n16090), .B2(n16628), .A(n12362), .ZN(n12363) );
  OAI21_X1 U14352 ( .B1(n16092), .B2(n12364), .A(n12363), .ZN(n12365) );
  AOI21_X1 U14353 ( .B1(n16094), .B2(n15855), .A(n12365), .ZN(n12366) );
  OAI21_X1 U14354 ( .B1(n16096), .B2(n15983), .A(n12366), .ZN(P1_U3278) );
  NAND2_X1 U14355 ( .A1(n12368), .A2(n12367), .ZN(n12370) );
  MUX2_X1 U14356 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n7416), .Z(n12512) );
  XNOR2_X1 U14357 ( .A(n12512), .B(SI_21_), .ZN(n12509) );
  XNOR2_X1 U14358 ( .A(n12511), .B(n12509), .ZN(n12957) );
  INV_X1 U14359 ( .A(n12957), .ZN(n12372) );
  OAI222_X1 U14360 ( .A1(n16139), .A2(n12796), .B1(n11886), .B2(n12372), .C1(
        P1_U3086), .C2(n15988), .ZN(P1_U3334) );
  OAI222_X1 U14361 ( .A1(n15545), .A2(n12958), .B1(n15540), .B2(n12372), .C1(
        n12371), .C2(P2_U3088), .ZN(P2_U3306) );
  NOR2_X1 U14362 ( .A1(n12846), .A2(n12374), .ZN(n12373) );
  AOI21_X1 U14363 ( .B1(n13728), .B2(n7413), .A(n12373), .ZN(n12380) );
  INV_X1 U14364 ( .A(n12380), .ZN(n12382) );
  OAI22_X1 U14365 ( .A1(n12375), .A2(n12940), .B1(n12374), .B2(n10271), .ZN(
        n12376) );
  XNOR2_X1 U14366 ( .A(n12376), .B(n10817), .ZN(n12381) );
  XOR2_X1 U14367 ( .A(n12380), .B(n12381), .Z(n12403) );
  AOI22_X1 U14368 ( .A1(n16722), .A2(n7412), .B1(n7413), .B2(n15680), .ZN(
        n12383) );
  XNOR2_X1 U14369 ( .A(n12383), .B(n10817), .ZN(n12524) );
  NOR2_X1 U14370 ( .A1(n12846), .A2(n12397), .ZN(n12384) );
  AOI21_X1 U14371 ( .B1(n16722), .B2(n7413), .A(n12384), .ZN(n12525) );
  XNOR2_X1 U14372 ( .A(n12524), .B(n12525), .ZN(n12526) );
  XNOR2_X1 U14373 ( .A(n12527), .B(n12526), .ZN(n12390) );
  AOI22_X1 U14374 ( .A1(n16530), .A2(n12385), .B1(P1_REG3_REG_13__SCAN_IN), 
        .B2(P1_U3086), .ZN(n12386) );
  OAI21_X1 U14375 ( .B1(n12387), .B2(n16535), .A(n12386), .ZN(n12388) );
  AOI21_X1 U14376 ( .B1(n16722), .B2(n15671), .A(n12388), .ZN(n12389) );
  OAI21_X1 U14377 ( .B1(n12390), .B2(n15673), .A(n12389), .ZN(P1_U3234) );
  XNOR2_X1 U14378 ( .A(n12391), .B(n13409), .ZN(n16687) );
  XNOR2_X1 U14379 ( .A(n12392), .B(n13409), .ZN(n12393) );
  OAI222_X1 U14380 ( .A1(n14314), .A2(n13934), .B1(n14312), .B2(n12577), .C1(
        n12393), .C2(n14310), .ZN(n16689) );
  NAND2_X1 U14381 ( .A1(n16689), .A2(n14352), .ZN(n12396) );
  OAI22_X1 U14382 ( .A1(n14384), .A2(n16686), .B1(n12583), .B2(n16508), .ZN(
        n12394) );
  AOI21_X1 U14383 ( .B1(P3_REG2_REG_11__SCAN_IN), .B2(n16517), .A(n12394), 
        .ZN(n12395) );
  OAI211_X1 U14384 ( .C1(n14358), .C2(n16687), .A(n12396), .B(n12395), .ZN(
        P3_U3222) );
  NAND2_X1 U14385 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_U3086), .ZN(n16265)
         );
  OAI21_X1 U14386 ( .B1(n15648), .B2(n12397), .A(n16265), .ZN(n12398) );
  AOI21_X1 U14387 ( .B1(n15659), .B2(n15682), .A(n12398), .ZN(n12399) );
  OAI21_X1 U14388 ( .B1(n12400), .B2(n16535), .A(n12399), .ZN(n12405) );
  AOI211_X1 U14389 ( .C1(n12403), .C2(n12402), .A(n15673), .B(n12401), .ZN(
        n12404) );
  AOI211_X1 U14390 ( .C1(n15671), .C2(n13728), .A(n12405), .B(n12404), .ZN(
        n12406) );
  INV_X1 U14391 ( .A(n12406), .ZN(P1_U3224) );
  AOI211_X1 U14392 ( .C1(n16704), .C2(n12409), .A(n12408), .B(n12407), .ZN(
        n12414) );
  INV_X1 U14393 ( .A(n15517), .ZN(n15512) );
  INV_X1 U14394 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n12410) );
  NOR2_X1 U14395 ( .A1(n16751), .A2(n12410), .ZN(n12411) );
  AOI21_X1 U14396 ( .B1(n13102), .B2(n15512), .A(n12411), .ZN(n12412) );
  OAI21_X1 U14397 ( .B1(n12414), .B2(n16748), .A(n12412), .ZN(P2_U3469) );
  AOI22_X1 U14398 ( .A1(n13102), .A2(n15457), .B1(n16746), .B2(
        P2_REG1_REG_13__SCAN_IN), .ZN(n12413) );
  OAI21_X1 U14399 ( .B1(n12414), .B2(n16746), .A(n12413), .ZN(P2_U3512) );
  AOI21_X1 U14400 ( .B1(n12416), .B2(n12415), .A(n13954), .ZN(n12418) );
  NAND2_X1 U14401 ( .A1(n12418), .A2(n12417), .ZN(n12425) );
  OAI22_X1 U14402 ( .A1(n12420), .A2(n13947), .B1(n13978), .B2(n12419), .ZN(
        n12421) );
  AOI211_X1 U14403 ( .C1(n16449), .C2(n12423), .A(n12422), .B(n12421), .ZN(
        n12424) );
  OAI211_X1 U14404 ( .C1(n12426), .C2(n13979), .A(n12425), .B(n12424), .ZN(
        P3_U3157) );
  NAND2_X1 U14405 ( .A1(n12540), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n12428) );
  NAND2_X1 U14406 ( .A1(n12428), .A2(n12427), .ZN(n12430) );
  INV_X1 U14407 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n12547) );
  XNOR2_X1 U14408 ( .A(n15709), .B(n12547), .ZN(n12429) );
  NAND2_X1 U14409 ( .A1(n12429), .A2(n12430), .ZN(n15703) );
  OAI211_X1 U14410 ( .C1(n12430), .C2(n12429), .A(n16263), .B(n15703), .ZN(
        n12437) );
  NAND2_X1 U14411 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n15607)
         );
  OAI21_X1 U14412 ( .B1(n16267), .B2(n7644), .A(n15607), .ZN(n12435) );
  AOI21_X1 U14413 ( .B1(n12540), .B2(P1_REG1_REG_16__SCAN_IN), .A(n12431), 
        .ZN(n12433) );
  XNOR2_X1 U14414 ( .A(n15709), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n12432) );
  NOR2_X1 U14415 ( .A1(n12433), .A2(n12432), .ZN(n15708) );
  AOI211_X1 U14416 ( .C1(n12433), .C2(n12432), .A(n15708), .B(n15710), .ZN(
        n12434) );
  AOI211_X1 U14417 ( .C1(n16261), .C2(n15709), .A(n12435), .B(n12434), .ZN(
        n12436) );
  NAND2_X1 U14418 ( .A1(n12437), .A2(n12436), .ZN(P1_U3260) );
  NAND2_X1 U14419 ( .A1(n12740), .A2(n12053), .ZN(n12440) );
  AOI22_X1 U14420 ( .A1(n12597), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n12596), 
        .B2(n12438), .ZN(n12439) );
  XNOR2_X1 U14421 ( .A(n15444), .B(n14936), .ZN(n12441) );
  AND2_X1 U14422 ( .A1(n15319), .A2(n14937), .ZN(n12442) );
  NAND2_X1 U14423 ( .A1(n12441), .A2(n12442), .ZN(n12604) );
  INV_X1 U14424 ( .A(n12441), .ZN(n12600) );
  INV_X1 U14425 ( .A(n12442), .ZN(n12443) );
  NAND2_X1 U14426 ( .A1(n12600), .A2(n12443), .ZN(n12444) );
  NAND2_X1 U14427 ( .A1(n12604), .A2(n12444), .ZN(n12451) );
  INV_X1 U14428 ( .A(n12445), .ZN(n12447) );
  NAND2_X1 U14429 ( .A1(n12447), .A2(n12446), .ZN(n12448) );
  AOI21_X1 U14430 ( .B1(n12451), .B2(n12450), .A(n15021), .ZN(n12452) );
  NAND2_X1 U14431 ( .A1(n12452), .A2(n12603), .ZN(n12464) );
  NAND2_X1 U14432 ( .A1(P2_U3088), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n16212)
         );
  OAI21_X1 U14433 ( .B1(n15003), .B2(n15351), .A(n16212), .ZN(n12462) );
  NAND2_X1 U14434 ( .A1(n12454), .A2(n12453), .ZN(n12455) );
  NAND2_X1 U14435 ( .A1(n12608), .A2(n12455), .ZN(n15331) );
  OR2_X1 U14436 ( .A1(n15331), .A2(n13262), .ZN(n12460) );
  NAND2_X1 U14437 ( .A1(n9790), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n12457) );
  NAND2_X1 U14438 ( .A1(n9788), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n12456) );
  OAI211_X1 U14439 ( .C1(n12113), .C2(n10470), .A(n12457), .B(n12456), .ZN(
        n12458) );
  INV_X1 U14440 ( .A(n12458), .ZN(n12459) );
  NAND2_X1 U14441 ( .A1(n12460), .A2(n12459), .ZN(n15344) );
  INV_X1 U14442 ( .A(n15344), .ZN(n14995) );
  NOR2_X1 U14443 ( .A1(n14972), .A2(n14995), .ZN(n12461) );
  AOI211_X1 U14444 ( .C1(n14974), .C2(n15342), .A(n12462), .B(n12461), .ZN(
        n12463) );
  OAI211_X1 U14445 ( .C1(n8329), .C2(n14994), .A(n12464), .B(n12463), .ZN(
        P2_U3210) );
  NAND2_X1 U14446 ( .A1(n16741), .A2(n15030), .ZN(n12465) );
  INV_X1 U14447 ( .A(n15029), .ZN(n12687) );
  XNOR2_X1 U14448 ( .A(n13113), .B(n12687), .ZN(n13328) );
  OAI21_X1 U14449 ( .B1(n12467), .B2(n13328), .A(n12497), .ZN(n15461) );
  INV_X1 U14450 ( .A(n15461), .ZN(n12481) );
  AOI22_X1 U14451 ( .A1(n15028), .A2(n15343), .B1(n15341), .B2(n15030), .ZN(
        n12473) );
  NAND2_X1 U14452 ( .A1(n16741), .A2(n12468), .ZN(n12469) );
  OAI211_X1 U14453 ( .C1(n8713), .C2(n8712), .A(n15346), .B(n12493), .ZN(
        n12472) );
  OAI211_X1 U14454 ( .C1(n12481), .C2(n10226), .A(n12473), .B(n12472), .ZN(
        n15459) );
  NAND2_X1 U14455 ( .A1(n15459), .A2(n15327), .ZN(n12480) );
  AOI211_X1 U14456 ( .C1(n13113), .C2(n12474), .A(n14937), .B(n8328), .ZN(
        n15460) );
  NOR2_X1 U14457 ( .A1(n15518), .A2(n15330), .ZN(n12478) );
  INV_X1 U14458 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n12476) );
  OAI22_X1 U14459 ( .A1(n15353), .A2(n12476), .B1(n12475), .B2(n15364), .ZN(
        n12477) );
  AOI211_X1 U14460 ( .C1(n15460), .C2(n15371), .A(n12478), .B(n12477), .ZN(
        n12479) );
  OAI211_X1 U14461 ( .C1(n12481), .C2(n15336), .A(n12480), .B(n12479), .ZN(
        P2_U3250) );
  INV_X1 U14462 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n12487) );
  INV_X1 U14463 ( .A(n13736), .ZN(n12482) );
  OAI22_X1 U14464 ( .A1(n12483), .A2(n16464), .B1(n12482), .B2(n16725), .ZN(
        n12484) );
  AOI211_X1 U14465 ( .C1(n12486), .C2(n16730), .A(n12485), .B(n12484), .ZN(
        n12489) );
  MUX2_X1 U14466 ( .A(n12487), .B(n12489), .S(n16737), .Z(n12488) );
  INV_X1 U14467 ( .A(n12488), .ZN(P1_U3501) );
  MUX2_X1 U14468 ( .A(n12490), .B(n12489), .S(n16734), .Z(n12491) );
  INV_X1 U14469 ( .A(n12491), .ZN(P1_U3542) );
  OR2_X1 U14470 ( .A1(n13113), .A2(n12687), .ZN(n12492) );
  XNOR2_X1 U14471 ( .A(n15511), .B(n13120), .ZN(n13329) );
  XNOR2_X1 U14472 ( .A(n12585), .B(n13329), .ZN(n12495) );
  AOI21_X1 U14473 ( .B1(n12495), .B2(n15346), .A(n12494), .ZN(n15454) );
  OR2_X1 U14474 ( .A1(n13113), .A2(n15029), .ZN(n12496) );
  INV_X1 U14475 ( .A(n13329), .ZN(n12498) );
  NAND2_X1 U14476 ( .A1(n12499), .A2(n12498), .ZN(n12500) );
  NAND2_X1 U14477 ( .A1(n12588), .A2(n12500), .ZN(n15455) );
  INV_X1 U14478 ( .A(n15455), .ZN(n12507) );
  AOI21_X1 U14479 ( .B1(n15511), .B2(n12501), .A(n14937), .ZN(n12502) );
  NAND2_X1 U14480 ( .A1(n12502), .A2(n12589), .ZN(n15453) );
  OAI22_X1 U14481 ( .A1(n15353), .A2(n11492), .B1(n12503), .B2(n15364), .ZN(
        n12504) );
  AOI21_X1 U14482 ( .B1(n15511), .B2(n15367), .A(n12504), .ZN(n12505) );
  OAI21_X1 U14483 ( .B1(n15453), .B2(n15233), .A(n12505), .ZN(n12506) );
  AOI21_X1 U14484 ( .B1(n12507), .B2(n15369), .A(n12506), .ZN(n12508) );
  OAI21_X1 U14485 ( .B1(n15362), .B2(n15454), .A(n12508), .ZN(P2_U3249) );
  INV_X1 U14486 ( .A(n12509), .ZN(n12510) );
  MUX2_X1 U14487 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(P1_DATAO_REG_22__SCAN_IN), 
        .S(n7416), .Z(n12622) );
  XNOR2_X1 U14488 ( .A(n12829), .B(n12622), .ZN(n12981) );
  INV_X1 U14489 ( .A(n12981), .ZN(n12516) );
  INV_X1 U14490 ( .A(n8082), .ZN(n12515) );
  OAI222_X1 U14491 ( .A1(n15545), .A2(n7827), .B1(n15540), .B2(n12516), .C1(
        n12515), .C2(P2_U3088), .ZN(P2_U3305) );
  NAND2_X1 U14492 ( .A1(n13736), .A2(n7412), .ZN(n12518) );
  NAND2_X1 U14493 ( .A1(n7413), .A2(n15679), .ZN(n12517) );
  NAND2_X1 U14494 ( .A1(n12518), .A2(n12517), .ZN(n12519) );
  XNOR2_X1 U14495 ( .A(n12519), .B(n12720), .ZN(n12523) );
  NOR2_X1 U14496 ( .A1(n12846), .A2(n12520), .ZN(n12521) );
  AOI21_X1 U14497 ( .B1(n13736), .B2(n7413), .A(n12521), .ZN(n12522) );
  NAND2_X1 U14498 ( .A1(n12523), .A2(n12522), .ZN(n12710) );
  OAI21_X1 U14499 ( .B1(n12523), .B2(n12522), .A(n12710), .ZN(n12530) );
  INV_X1 U14500 ( .A(n12711), .ZN(n12528) );
  AOI21_X1 U14501 ( .B1(n12530), .B2(n12529), .A(n12528), .ZN(n12537) );
  OAI21_X1 U14502 ( .B1(n15648), .B2(n12713), .A(n12531), .ZN(n12532) );
  AOI21_X1 U14503 ( .B1(n15659), .B2(n15680), .A(n12532), .ZN(n12533) );
  OAI21_X1 U14504 ( .B1(n12534), .B2(n16535), .A(n12533), .ZN(n12535) );
  AOI21_X1 U14505 ( .B1(n13736), .B2(n15671), .A(n12535), .ZN(n12536) );
  OAI21_X1 U14506 ( .B1(n12537), .B2(n15673), .A(n12536), .ZN(P1_U3215) );
  NAND2_X1 U14507 ( .A1(n12539), .A2(n11544), .ZN(n12542) );
  AOI22_X1 U14508 ( .A1(n12540), .A2(n12759), .B1(n12760), .B2(
        P2_DATAO_REG_16__SCAN_IN), .ZN(n12541) );
  NAND2_X1 U14509 ( .A1(n16085), .A2(n12722), .ZN(n15766) );
  OR2_X1 U14510 ( .A1(n16085), .A2(n12722), .ZN(n12543) );
  OAI21_X1 U14511 ( .B1(n7603), .B2(n13595), .A(n15767), .ZN(n12553) );
  INV_X1 U14512 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n12544) );
  NAND2_X1 U14513 ( .A1(n12545), .A2(n12544), .ZN(n12546) );
  NAND2_X1 U14514 ( .A1(n12745), .A2(n12546), .ZN(n15978) );
  OR2_X1 U14515 ( .A1(n15978), .A2(n12946), .ZN(n12552) );
  NAND2_X1 U14516 ( .A1(n13566), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n12551) );
  OR2_X1 U14517 ( .A1(n12929), .A2(n12547), .ZN(n12550) );
  INV_X1 U14518 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n12548) );
  OR2_X1 U14519 ( .A1(n12862), .A2(n12548), .ZN(n12549) );
  NAND4_X1 U14520 ( .A1(n12552), .A2(n12551), .A3(n12550), .A4(n12549), .ZN(
        n15755) );
  AOI222_X1 U14521 ( .A1(n16561), .A2(n12553), .B1(n15755), .B2(n16462), .C1(
        n15678), .C2(n15971), .ZN(n16087) );
  INV_X1 U14522 ( .A(n13592), .ZN(n12554) );
  OAI21_X1 U14523 ( .B1(n12557), .B2(n12556), .A(n15753), .ZN(n12558) );
  INV_X1 U14524 ( .A(n12558), .ZN(n16088) );
  NAND2_X1 U14525 ( .A1(n7414), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n12559) );
  OAI21_X1 U14526 ( .B1(n16622), .B2(n15599), .A(n12559), .ZN(n12560) );
  AOI21_X1 U14527 ( .B1(n16085), .B2(n16628), .A(n12560), .ZN(n12564) );
  AOI21_X1 U14528 ( .B1(n16085), .B2(n12561), .A(n16464), .ZN(n12562) );
  AND2_X1 U14529 ( .A1(n12562), .A2(n15977), .ZN(n16084) );
  NAND2_X1 U14530 ( .A1(n16084), .A2(n16486), .ZN(n12563) );
  OAI211_X1 U14531 ( .C1(n16088), .C2(n15983), .A(n12564), .B(n12563), .ZN(
        n12565) );
  INV_X1 U14532 ( .A(n12565), .ZN(n12566) );
  OAI21_X1 U14533 ( .B1(n7414), .B2(n16087), .A(n12566), .ZN(P1_U3277) );
  XNOR2_X1 U14534 ( .A(n12567), .B(n13414), .ZN(n16714) );
  XNOR2_X1 U14535 ( .A(n12568), .B(n13414), .ZN(n12569) );
  OAI222_X1 U14536 ( .A1(n14314), .A2(n12570), .B1(n14312), .B2(n13934), .C1(
        n12569), .C2(n14310), .ZN(n16716) );
  NAND2_X1 U14537 ( .A1(n16716), .A2(n14352), .ZN(n12573) );
  INV_X1 U14538 ( .A(n16712), .ZN(n13939) );
  OAI22_X1 U14539 ( .A1(n14352), .A2(n9156), .B1(n13937), .B2(n16508), .ZN(
        n12571) );
  AOI21_X1 U14540 ( .B1(n13939), .B2(n14354), .A(n12571), .ZN(n12572) );
  OAI211_X1 U14541 ( .C1(n14358), .C2(n16714), .A(n12573), .B(n12572), .ZN(
        P3_U3220) );
  OAI211_X1 U14542 ( .C1(n12576), .C2(n12575), .A(n12574), .B(n16451), .ZN(
        n12582) );
  OAI22_X1 U14543 ( .A1(n12577), .A2(n13947), .B1(n13978), .B2(n13934), .ZN(
        n12578) );
  AOI211_X1 U14544 ( .C1(n16449), .C2(n12580), .A(n12579), .B(n12578), .ZN(
        n12581) );
  OAI211_X1 U14545 ( .C1(n12583), .C2(n13979), .A(n12582), .B(n12581), .ZN(
        P3_U3176) );
  NAND2_X1 U14546 ( .A1(n15511), .A2(n13120), .ZN(n12584) );
  XNOR2_X1 U14547 ( .A(n15149), .B(n15148), .ZN(n12586) );
  OAI222_X1 U14548 ( .A1(n15287), .A2(n15150), .B1(n15289), .B2(n13120), .C1(
        n12586), .C2(n15308), .ZN(n15448) );
  INV_X1 U14549 ( .A(n15448), .ZN(n12595) );
  NAND2_X1 U14550 ( .A1(n15511), .A2(n15028), .ZN(n12587) );
  XNOR2_X1 U14551 ( .A(n15122), .B(n15148), .ZN(n15450) );
  AOI211_X1 U14552 ( .C1(n8008), .C2(n12589), .A(n14937), .B(n8326), .ZN(
        n15449) );
  NAND2_X1 U14553 ( .A1(n15449), .A2(n15371), .ZN(n12592) );
  AOI22_X1 U14554 ( .A1(n15362), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n12590), 
        .B2(n15292), .ZN(n12591) );
  OAI211_X1 U14555 ( .C1(n8761), .C2(n15330), .A(n12592), .B(n12591), .ZN(
        n12593) );
  AOI21_X1 U14556 ( .B1(n15450), .B2(n15369), .A(n12593), .ZN(n12594) );
  OAI21_X1 U14557 ( .B1(n15362), .B2(n12595), .A(n12594), .ZN(P2_U3248) );
  NAND2_X1 U14558 ( .A1(n12758), .A2(n12053), .ZN(n12599) );
  AOI22_X1 U14559 ( .A1(n12597), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n12596), 
        .B2(n13341), .ZN(n12598) );
  NOR3_X1 U14560 ( .A1(n12600), .A2(n15150), .A3(n15011), .ZN(n12606) );
  XNOR2_X1 U14561 ( .A(n15329), .B(n14959), .ZN(n14996) );
  AND2_X1 U14562 ( .A1(n15344), .A2(n14937), .ZN(n12601) );
  NAND2_X1 U14563 ( .A1(n14996), .A2(n12601), .ZN(n12973) );
  OAI21_X1 U14564 ( .B1(n14996), .B2(n12601), .A(n12973), .ZN(n12602) );
  AOI21_X1 U14565 ( .B1(n12602), .B2(n12603), .A(n15021), .ZN(n12605) );
  OAI21_X1 U14566 ( .B1(n12606), .B2(n12605), .A(n8292), .ZN(n12617) );
  OAI21_X1 U14567 ( .B1(n15003), .B2(n15331), .A(n12607), .ZN(n12615) );
  NAND2_X1 U14568 ( .A1(n12608), .A2(n15002), .ZN(n12609) );
  NAND2_X1 U14569 ( .A1(n12962), .A2(n12609), .ZN(n15301) );
  INV_X1 U14570 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n15436) );
  NAND2_X1 U14571 ( .A1(n9789), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n12611) );
  NAND2_X1 U14572 ( .A1(n9788), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n12610) );
  OAI211_X1 U14573 ( .C1(n13265), .C2(n15436), .A(n12611), .B(n12610), .ZN(
        n12612) );
  INV_X1 U14574 ( .A(n12612), .ZN(n12613) );
  OAI21_X1 U14575 ( .B1(n15301), .B2(n13262), .A(n12613), .ZN(n15320) );
  INV_X1 U14576 ( .A(n15320), .ZN(n15288) );
  NOR2_X1 U14577 ( .A1(n14972), .A2(n15288), .ZN(n12614) );
  AOI211_X1 U14578 ( .C1(n14974), .C2(n15319), .A(n12615), .B(n12614), .ZN(
        n12616) );
  OAI211_X1 U14579 ( .C1(n15504), .C2(n14994), .A(n12617), .B(n12616), .ZN(
        P2_U3191) );
  MUX2_X1 U14580 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n7416), .Z(n12832) );
  INV_X1 U14581 ( .A(n12832), .ZN(n12619) );
  NAND2_X1 U14582 ( .A1(n12619), .A2(n12618), .ZN(n12623) );
  OAI21_X1 U14583 ( .B1(SI_22_), .B2(n12622), .A(n12623), .ZN(n12620) );
  INV_X1 U14584 ( .A(n12620), .ZN(n12621) );
  INV_X1 U14585 ( .A(n12622), .ZN(n12831) );
  NOR2_X1 U14586 ( .A1(n12831), .A2(n14655), .ZN(n12624) );
  AOI22_X1 U14587 ( .A1(n12624), .A2(n12623), .B1(n12832), .B2(SI_23_), .ZN(
        n12625) );
  MUX2_X1 U14588 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n7416), .Z(n12854) );
  NAND2_X1 U14589 ( .A1(n12626), .A2(n12854), .ZN(n12629) );
  MUX2_X1 U14590 ( .A(n16131), .B(n15537), .S(n7416), .Z(n12630) );
  NAND2_X1 U14591 ( .A1(n12630), .A2(n14656), .ZN(n12633) );
  INV_X1 U14592 ( .A(n12630), .ZN(n12631) );
  NAND2_X1 U14593 ( .A1(n12631), .A2(SI_25_), .ZN(n12632) );
  NAND2_X1 U14594 ( .A1(n12633), .A2(n12632), .ZN(n12875) );
  MUX2_X1 U14595 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(P1_DATAO_REG_26__SCAN_IN), 
        .S(n7416), .Z(n12634) );
  MUX2_X1 U14596 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(P1_DATAO_REG_27__SCAN_IN), 
        .S(n7416), .Z(n12636) );
  XNOR2_X1 U14597 ( .A(n12636), .B(SI_27_), .ZN(n12914) );
  INV_X1 U14598 ( .A(n12914), .ZN(n12635) );
  NAND2_X1 U14599 ( .A1(n12636), .A2(SI_27_), .ZN(n12637) );
  MUX2_X1 U14600 ( .A(n12927), .B(n13256), .S(n7416), .Z(n12639) );
  NAND2_X1 U14601 ( .A1(n12639), .A2(n14919), .ZN(n12642) );
  INV_X1 U14602 ( .A(n12639), .ZN(n12640) );
  NAND2_X1 U14603 ( .A1(n12640), .A2(SI_28_), .ZN(n12641) );
  NAND2_X1 U14604 ( .A1(n12642), .A2(n12641), .ZN(n12652) );
  MUX2_X1 U14605 ( .A(n13600), .B(n13493), .S(n7416), .Z(n12643) );
  NAND2_X1 U14606 ( .A1(n12643), .A2(n14914), .ZN(n13217) );
  INV_X1 U14607 ( .A(n12643), .ZN(n12644) );
  NAND2_X1 U14608 ( .A1(n12644), .A2(SI_29_), .ZN(n12645) );
  INV_X1 U14609 ( .A(n13599), .ZN(n12654) );
  OAI222_X1 U14610 ( .A1(n15540), .A2(n12654), .B1(P2_U3088), .B2(n12646), 
        .C1(n13493), .C2(n15545), .ZN(P2_U3298) );
  NAND2_X1 U14611 ( .A1(P1_REG3_REG_0__SCAN_IN), .A2(n12647), .ZN(n12648) );
  OAI21_X1 U14612 ( .B1(n12649), .B2(n15673), .A(n12648), .ZN(n12650) );
  AOI21_X1 U14613 ( .B1(n15658), .B2(n10430), .A(n12650), .ZN(n12651) );
  OAI21_X1 U14614 ( .B1(n15653), .B2(n15990), .A(n12651), .ZN(P1_U3232) );
  INV_X1 U14615 ( .A(n13255), .ZN(n15530) );
  OAI222_X1 U14616 ( .A1(n16139), .A2(n12927), .B1(n11886), .B2(n15530), .C1(
        P1_U3086), .C2(n10019), .ZN(P1_U3327) );
  OAI222_X1 U14617 ( .A1(n16139), .A2(n13600), .B1(P1_U3086), .B2(n12655), 
        .C1(n11886), .C2(n12654), .ZN(P1_U3326) );
  INV_X1 U14618 ( .A(n12656), .ZN(n12660) );
  NAND2_X1 U14619 ( .A1(n14961), .A2(n15036), .ZN(n12657) );
  OAI21_X1 U14620 ( .B1(n12658), .B2(n15021), .A(n12657), .ZN(n12659) );
  NAND3_X1 U14621 ( .A1(n12682), .A2(n12660), .A3(n12659), .ZN(n12668) );
  OAI21_X1 U14622 ( .B1(n15003), .B2(n12662), .A(n12661), .ZN(n12663) );
  AOI21_X1 U14623 ( .B1(n14974), .B2(n15036), .A(n12663), .ZN(n12667) );
  NAND2_X1 U14624 ( .A1(n15024), .A2(n13077), .ZN(n12666) );
  OR2_X1 U14625 ( .A1(n14972), .A2(n12664), .ZN(n12665) );
  AND4_X1 U14626 ( .A1(n12668), .A2(n12667), .A3(n12666), .A4(n12665), .ZN(
        n12669) );
  OAI21_X1 U14627 ( .B1(n11101), .B2(n15021), .A(n12669), .ZN(P2_U3203) );
  INV_X1 U14628 ( .A(n12670), .ZN(n12672) );
  OAI21_X1 U14629 ( .B1(n15003), .B2(n12672), .A(n12671), .ZN(n12673) );
  AOI21_X1 U14630 ( .B1(n14974), .B2(n15037), .A(n12673), .ZN(n12674) );
  OAI21_X1 U14631 ( .B1(n13079), .B2(n14972), .A(n12674), .ZN(n12680) );
  AOI22_X1 U14632 ( .A1(n14961), .A2(n15037), .B1(n15000), .B2(n12675), .ZN(
        n12677) );
  NOR3_X1 U14633 ( .A1(n12678), .A2(n12677), .A3(n12676), .ZN(n12679) );
  AOI211_X1 U14634 ( .C1(n13071), .C2(n15024), .A(n12680), .B(n12679), .ZN(
        n12681) );
  OAI21_X1 U14635 ( .B1(n12682), .B2(n15021), .A(n12681), .ZN(P2_U3193) );
  OAI21_X1 U14636 ( .B1(n15003), .B2(n12684), .A(n12683), .ZN(n12685) );
  AOI21_X1 U14637 ( .B1(n14974), .B2(n15031), .A(n12685), .ZN(n12686) );
  OAI21_X1 U14638 ( .B1(n12687), .B2(n14972), .A(n12686), .ZN(n12694) );
  NOR3_X1 U14639 ( .A1(n12688), .A2(n12697), .A3(n15011), .ZN(n12689) );
  AOI21_X1 U14640 ( .B1(n12690), .B2(n15014), .A(n12689), .ZN(n12692) );
  NOR2_X1 U14641 ( .A1(n12692), .A2(n12691), .ZN(n12693) );
  AOI211_X1 U14642 ( .C1(n16741), .C2(n15024), .A(n12694), .B(n12693), .ZN(
        n12695) );
  OAI21_X1 U14643 ( .B1(n12696), .B2(n15021), .A(n12695), .ZN(P2_U3187) );
  NOR2_X1 U14644 ( .A1(n14972), .A2(n12697), .ZN(n12701) );
  NAND2_X1 U14645 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3088), .ZN(n16235)
         );
  NAND2_X1 U14646 ( .A1(n15018), .A2(n12698), .ZN(n12699) );
  OAI211_X1 U14647 ( .C1(n12994), .C2(n13089), .A(n16235), .B(n12699), .ZN(
        n12700) );
  AOI211_X1 U14648 ( .C1(n16700), .C2(n15024), .A(n12701), .B(n12700), .ZN(
        n12708) );
  INV_X1 U14649 ( .A(n12702), .ZN(n12705) );
  OAI22_X1 U14650 ( .A1(n12703), .A2(n15021), .B1(n13089), .B2(n15011), .ZN(
        n12704) );
  NAND3_X1 U14651 ( .A1(n12706), .A2(n12705), .A3(n12704), .ZN(n12707) );
  OAI211_X1 U14652 ( .C1(n12709), .C2(n15021), .A(n12708), .B(n12707), .ZN(
        P2_U3196) );
  NAND2_X1 U14653 ( .A1(n12711), .A2(n12710), .ZN(n12716) );
  OAI22_X1 U14654 ( .A1(n8605), .A2(n12940), .B1(n12713), .B2(n10271), .ZN(
        n12712) );
  XNOR2_X1 U14655 ( .A(n12712), .B(n10817), .ZN(n12714) );
  OAI22_X1 U14656 ( .A1(n8605), .A2(n10271), .B1(n12713), .B2(n12846), .ZN(
        n15665) );
  NAND2_X1 U14657 ( .A1(n15666), .A2(n15665), .ZN(n12717) );
  INV_X1 U14658 ( .A(n12714), .ZN(n12715) );
  NAND2_X1 U14659 ( .A1(n16085), .A2(n7412), .ZN(n12719) );
  NAND2_X1 U14660 ( .A1(n7413), .A2(n15972), .ZN(n12718) );
  NAND2_X1 U14661 ( .A1(n12719), .A2(n12718), .ZN(n12721) );
  XNOR2_X1 U14662 ( .A(n12721), .B(n12720), .ZN(n12725) );
  NOR2_X1 U14663 ( .A1(n12846), .A2(n12722), .ZN(n12723) );
  AOI21_X1 U14664 ( .B1(n16085), .B2(n7413), .A(n12723), .ZN(n12724) );
  NAND2_X1 U14665 ( .A1(n12725), .A2(n12724), .ZN(n12727) );
  OAI21_X1 U14666 ( .B1(n12725), .B2(n12724), .A(n12727), .ZN(n15595) );
  INV_X1 U14667 ( .A(n15595), .ZN(n12726) );
  AOI22_X1 U14668 ( .A1(n15709), .A2(n12759), .B1(n12760), .B2(
        P2_DATAO_REG_17__SCAN_IN), .ZN(n12729) );
  NAND2_X1 U14669 ( .A1(n16078), .A2(n7412), .ZN(n12732) );
  NAND2_X1 U14670 ( .A1(n7413), .A2(n15755), .ZN(n12731) );
  NAND2_X1 U14671 ( .A1(n12732), .A2(n12731), .ZN(n12733) );
  XNOR2_X1 U14672 ( .A(n12733), .B(n10817), .ZN(n12737) );
  NAND2_X1 U14673 ( .A1(n16078), .A2(n7413), .ZN(n12735) );
  NAND2_X1 U14674 ( .A1(n12921), .A2(n15755), .ZN(n12734) );
  NAND2_X1 U14675 ( .A1(n12735), .A2(n12734), .ZN(n12736) );
  NOR2_X1 U14676 ( .A1(n12737), .A2(n12736), .ZN(n12738) );
  AOI21_X1 U14677 ( .B1(n12737), .B2(n12736), .A(n12738), .ZN(n15605) );
  INV_X1 U14678 ( .A(n12738), .ZN(n12739) );
  NAND2_X1 U14679 ( .A1(n15603), .A2(n12739), .ZN(n15645) );
  NAND2_X1 U14680 ( .A1(n12740), .A2(n11544), .ZN(n12743) );
  NOR2_X1 U14681 ( .A1(n10704), .A2(n8120), .ZN(n12741) );
  AOI21_X1 U14682 ( .B1(n15723), .B2(n12759), .A(n12741), .ZN(n12742) );
  NAND2_X1 U14683 ( .A1(n16074), .A2(n7412), .ZN(n12752) );
  NAND2_X1 U14684 ( .A1(n12745), .A2(n12744), .ZN(n12746) );
  NAND2_X1 U14685 ( .A1(n12764), .A2(n12746), .ZN(n15963) );
  INV_X1 U14686 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n15711) );
  OR2_X1 U14687 ( .A1(n12862), .A2(n15711), .ZN(n12748) );
  INV_X1 U14688 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n15964) );
  OR2_X1 U14689 ( .A1(n12929), .A2(n15964), .ZN(n12747) );
  AND2_X1 U14690 ( .A1(n12748), .A2(n12747), .ZN(n12750) );
  NAND2_X1 U14691 ( .A1(n13566), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n12749) );
  OAI211_X1 U14692 ( .C1(n15963), .C2(n12946), .A(n12750), .B(n12749), .ZN(
        n15973) );
  NAND2_X1 U14693 ( .A1(n15973), .A2(n7413), .ZN(n12751) );
  NAND2_X1 U14694 ( .A1(n12752), .A2(n12751), .ZN(n12753) );
  XNOR2_X1 U14695 ( .A(n12753), .B(n10817), .ZN(n12754) );
  AOI22_X1 U14696 ( .A1(n16074), .A2(n7413), .B1(n12921), .B2(n15973), .ZN(
        n12755) );
  XNOR2_X1 U14697 ( .A(n12754), .B(n12755), .ZN(n15646) );
  INV_X1 U14698 ( .A(n12754), .ZN(n12756) );
  NAND2_X1 U14699 ( .A1(n12756), .A2(n12755), .ZN(n12757) );
  NAND2_X1 U14700 ( .A1(n12758), .A2(n11544), .ZN(n12762) );
  AOI22_X1 U14701 ( .A1(n12760), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n13606), 
        .B2(n12759), .ZN(n12761) );
  NAND2_X1 U14702 ( .A1(n16068), .A2(n7412), .ZN(n12771) );
  INV_X1 U14703 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n12769) );
  INV_X1 U14704 ( .A(n12782), .ZN(n12766) );
  NAND2_X1 U14705 ( .A1(n12764), .A2(n12763), .ZN(n12765) );
  NAND2_X1 U14706 ( .A1(n12766), .A2(n12765), .ZN(n15940) );
  OR2_X1 U14707 ( .A1(n15940), .A2(n12946), .ZN(n12768) );
  AOI22_X1 U14708 ( .A1(n7420), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n13566), 
        .B2(P1_REG0_REG_19__SCAN_IN), .ZN(n12767) );
  OAI211_X1 U14709 ( .C1(n12862), .C2(n12769), .A(n12768), .B(n12767), .ZN(
        n15756) );
  NAND2_X1 U14710 ( .A1(n15756), .A2(n7413), .ZN(n12770) );
  NAND2_X1 U14711 ( .A1(n12771), .A2(n12770), .ZN(n12772) );
  XNOR2_X1 U14712 ( .A(n12772), .B(n10817), .ZN(n12775) );
  NAND2_X1 U14713 ( .A1(n16068), .A2(n7413), .ZN(n12774) );
  NAND2_X1 U14714 ( .A1(n15756), .A2(n12921), .ZN(n12773) );
  NAND2_X1 U14715 ( .A1(n12774), .A2(n12773), .ZN(n12776) );
  NAND2_X1 U14716 ( .A1(n12775), .A2(n12776), .ZN(n15566) );
  INV_X1 U14717 ( .A(n12775), .ZN(n12778) );
  INV_X1 U14718 ( .A(n12776), .ZN(n12777) );
  NAND2_X1 U14719 ( .A1(n12778), .A2(n12777), .ZN(n15565) );
  OR2_X1 U14720 ( .A1(n10704), .A2(n12779), .ZN(n12780) );
  NOR2_X1 U14721 ( .A1(n12782), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n12783) );
  OR2_X1 U14722 ( .A1(n12799), .A2(n12783), .ZN(n15919) );
  INV_X1 U14723 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n12786) );
  NAND2_X1 U14724 ( .A1(n13566), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n12785) );
  NAND2_X1 U14725 ( .A1(n7420), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n12784) );
  OAI211_X1 U14726 ( .C1(n12862), .C2(n12786), .A(n12785), .B(n12784), .ZN(
        n12787) );
  INV_X1 U14727 ( .A(n12787), .ZN(n12788) );
  OAI21_X1 U14728 ( .B1(n15919), .B2(n12946), .A(n12788), .ZN(n15759) );
  AOI22_X1 U14729 ( .A1(n16059), .A2(n7412), .B1(n7413), .B2(n15759), .ZN(
        n12789) );
  XNOR2_X1 U14730 ( .A(n12789), .B(n10817), .ZN(n12791) );
  AOI22_X1 U14731 ( .A1(n16059), .A2(n7413), .B1(n12921), .B2(n15759), .ZN(
        n12792) );
  XNOR2_X1 U14732 ( .A(n12791), .B(n12792), .ZN(n15628) );
  INV_X1 U14733 ( .A(n15628), .ZN(n12790) );
  INV_X1 U14734 ( .A(n12791), .ZN(n12794) );
  INV_X1 U14735 ( .A(n12792), .ZN(n12793) );
  NAND2_X1 U14736 ( .A1(n12794), .A2(n12793), .ZN(n12795) );
  NAND2_X1 U14737 ( .A1(n12957), .A2(n11544), .ZN(n12798) );
  OR2_X1 U14738 ( .A1(n10704), .A2(n12796), .ZN(n12797) );
  OR2_X1 U14739 ( .A1(n12799), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n12801) );
  AND2_X1 U14740 ( .A1(n12801), .A2(n12800), .ZN(n15905) );
  NAND2_X1 U14741 ( .A1(n15905), .A2(n12802), .ZN(n12808) );
  INV_X1 U14742 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n12805) );
  NAND2_X1 U14743 ( .A1(n7420), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n12804) );
  NAND2_X1 U14744 ( .A1(n13566), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n12803) );
  OAI211_X1 U14745 ( .C1(n12805), .C2(n12862), .A(n12804), .B(n12803), .ZN(
        n12806) );
  INV_X1 U14746 ( .A(n12806), .ZN(n12807) );
  NAND2_X1 U14747 ( .A1(n12808), .A2(n12807), .ZN(n15676) );
  INV_X1 U14748 ( .A(n15676), .ZN(n15772) );
  OAI22_X1 U14749 ( .A1(n16053), .A2(n12940), .B1(n15772), .B2(n10271), .ZN(
        n12809) );
  XNOR2_X1 U14750 ( .A(n12809), .B(n10817), .ZN(n12811) );
  OAI22_X1 U14751 ( .A1(n16053), .A2(n10271), .B1(n15772), .B2(n12846), .ZN(
        n12810) );
  XNOR2_X1 U14752 ( .A(n12811), .B(n12810), .ZN(n15577) );
  OR2_X1 U14753 ( .A1(n12811), .A2(n12810), .ZN(n12812) );
  NAND2_X1 U14754 ( .A1(n12945), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n12822) );
  INV_X1 U14755 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n12815) );
  OR2_X1 U14756 ( .A1(n12929), .A2(n12815), .ZN(n12821) );
  OAI21_X1 U14757 ( .B1(P1_REG3_REG_22__SCAN_IN), .B2(n12817), .A(n12816), 
        .ZN(n15895) );
  OR2_X1 U14758 ( .A1(n12946), .A2(n15895), .ZN(n12820) );
  INV_X1 U14759 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n12818) );
  OR2_X1 U14760 ( .A1(n10418), .A2(n12818), .ZN(n12819) );
  OAI22_X1 U14761 ( .A1(n16046), .A2(n12940), .B1(n15761), .B2(n10271), .ZN(
        n12823) );
  XNOR2_X1 U14762 ( .A(n12823), .B(n10817), .ZN(n12825) );
  OAI22_X1 U14763 ( .A1(n16046), .A2(n10271), .B1(n15761), .B2(n12846), .ZN(
        n12826) );
  XNOR2_X1 U14764 ( .A(n12825), .B(n12826), .ZN(n15632) );
  INV_X1 U14765 ( .A(n15632), .ZN(n12824) );
  INV_X1 U14766 ( .A(n12825), .ZN(n12828) );
  INV_X1 U14767 ( .A(n12826), .ZN(n12827) );
  INV_X1 U14768 ( .A(n15559), .ZN(n12848) );
  NAND2_X1 U14769 ( .A1(n16136), .A2(n11544), .ZN(n12834) );
  OR2_X1 U14770 ( .A1(n10704), .A2(n16140), .ZN(n12833) );
  NAND2_X1 U14771 ( .A1(n16040), .A2(n7412), .ZN(n12844) );
  NAND2_X1 U14772 ( .A1(n12945), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n12842) );
  INV_X1 U14773 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n12835) );
  OR2_X1 U14774 ( .A1(n12929), .A2(n12835), .ZN(n12841) );
  OAI21_X1 U14775 ( .B1(P1_REG3_REG_23__SCAN_IN), .B2(n12837), .A(n12836), 
        .ZN(n15878) );
  OR2_X1 U14776 ( .A1(n12946), .A2(n15878), .ZN(n12840) );
  INV_X1 U14777 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n12838) );
  OR2_X1 U14778 ( .A1(n10418), .A2(n12838), .ZN(n12839) );
  NAND4_X1 U14779 ( .A1(n12842), .A2(n12841), .A3(n12840), .A4(n12839), .ZN(
        n15860) );
  NAND2_X1 U14780 ( .A1(n7413), .A2(n15860), .ZN(n12843) );
  NAND2_X1 U14781 ( .A1(n12844), .A2(n12843), .ZN(n12845) );
  XNOR2_X1 U14782 ( .A(n12845), .B(n10817), .ZN(n12849) );
  INV_X1 U14783 ( .A(n16040), .ZN(n15882) );
  OAI22_X1 U14784 ( .A1(n15882), .A2(n10271), .B1(n15777), .B2(n12846), .ZN(
        n12850) );
  XNOR2_X1 U14785 ( .A(n12849), .B(n12850), .ZN(n15560) );
  INV_X1 U14786 ( .A(n12849), .ZN(n12852) );
  INV_X1 U14787 ( .A(n12850), .ZN(n12851) );
  NAND2_X1 U14788 ( .A1(n12852), .A2(n12851), .ZN(n12853) );
  NAND2_X1 U14789 ( .A1(n15538), .A2(n11544), .ZN(n12857) );
  INV_X1 U14790 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n16134) );
  OR2_X1 U14791 ( .A1(n10704), .A2(n16134), .ZN(n12856) );
  INV_X1 U14792 ( .A(n15869), .ZN(n15763) );
  NAND2_X1 U14793 ( .A1(n7420), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n12866) );
  INV_X1 U14794 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n12858) );
  OR2_X1 U14795 ( .A1(n7418), .A2(n12858), .ZN(n12865) );
  OAI21_X1 U14796 ( .B1(P1_REG3_REG_24__SCAN_IN), .B2(n12860), .A(n12859), 
        .ZN(n15867) );
  OR2_X1 U14797 ( .A1(n12946), .A2(n15867), .ZN(n12864) );
  INV_X1 U14798 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n12861) );
  OR2_X1 U14799 ( .A1(n12862), .A2(n12861), .ZN(n12863) );
  NAND4_X1 U14800 ( .A1(n12866), .A2(n12865), .A3(n12864), .A4(n12863), .ZN(
        n15675) );
  OAI22_X1 U14801 ( .A1(n15763), .A2(n10271), .B1(n15778), .B2(n12846), .ZN(
        n12871) );
  NAND2_X1 U14802 ( .A1(n15869), .A2(n7412), .ZN(n12868) );
  NAND2_X1 U14803 ( .A1(n7413), .A2(n15675), .ZN(n12867) );
  NAND2_X1 U14804 ( .A1(n12868), .A2(n12867), .ZN(n12869) );
  XNOR2_X1 U14805 ( .A(n12869), .B(n10817), .ZN(n12870) );
  XOR2_X1 U14806 ( .A(n12871), .B(n12870), .Z(n15614) );
  INV_X1 U14807 ( .A(n12870), .ZN(n12873) );
  INV_X1 U14808 ( .A(n12871), .ZN(n12872) );
  NAND2_X1 U14809 ( .A1(n12873), .A2(n12872), .ZN(n12874) );
  NAND2_X1 U14810 ( .A1(n15535), .A2(n11544), .ZN(n12878) );
  OR2_X1 U14811 ( .A1(n10704), .A2(n16131), .ZN(n12877) );
  NAND2_X1 U14812 ( .A1(n15738), .A2(n7412), .ZN(n12887) );
  NAND2_X1 U14813 ( .A1(n12945), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n12885) );
  INV_X1 U14814 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n12879) );
  OR2_X1 U14815 ( .A1(n12929), .A2(n12879), .ZN(n12884) );
  OAI21_X1 U14816 ( .B1(P1_REG3_REG_25__SCAN_IN), .B2(n12880), .A(n12897), 
        .ZN(n15850) );
  OR2_X1 U14817 ( .A1(n12946), .A2(n15850), .ZN(n12883) );
  INV_X1 U14818 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n12881) );
  OR2_X1 U14819 ( .A1(n10418), .A2(n12881), .ZN(n12882) );
  NAND2_X1 U14820 ( .A1(n7413), .A2(n15859), .ZN(n12886) );
  NAND2_X1 U14821 ( .A1(n12887), .A2(n12886), .ZN(n12888) );
  XNOR2_X1 U14822 ( .A(n12888), .B(n10817), .ZN(n12889) );
  AOI22_X1 U14823 ( .A1(n15738), .A2(n7413), .B1(n12921), .B2(n15859), .ZN(
        n12890) );
  XNOR2_X1 U14824 ( .A(n12889), .B(n12890), .ZN(n15585) );
  INV_X1 U14825 ( .A(n12889), .ZN(n12891) );
  NAND2_X1 U14826 ( .A1(n15532), .A2(n11544), .ZN(n12894) );
  OR2_X1 U14827 ( .A1(n10704), .A2(n16125), .ZN(n12893) );
  NAND2_X1 U14828 ( .A1(n16021), .A2(n7412), .ZN(n12905) );
  NAND2_X1 U14829 ( .A1(n12945), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n12903) );
  INV_X1 U14830 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n12895) );
  OR2_X1 U14831 ( .A1(n12929), .A2(n12895), .ZN(n12902) );
  INV_X1 U14832 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n12896) );
  NAND2_X1 U14833 ( .A1(n12897), .A2(n12896), .ZN(n12898) );
  NAND2_X1 U14834 ( .A1(n12931), .A2(n12898), .ZN(n15831) );
  OR2_X1 U14835 ( .A1(n12946), .A2(n15831), .ZN(n12901) );
  INV_X1 U14836 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n12899) );
  OR2_X1 U14837 ( .A1(n7418), .A2(n12899), .ZN(n12900) );
  NAND4_X1 U14838 ( .A1(n12903), .A2(n12902), .A3(n12901), .A4(n12900), .ZN(
        n15765) );
  NAND2_X1 U14839 ( .A1(n7413), .A2(n15765), .ZN(n12904) );
  NAND2_X1 U14840 ( .A1(n12905), .A2(n12904), .ZN(n12906) );
  XNOR2_X1 U14841 ( .A(n12906), .B(n10817), .ZN(n12909) );
  NAND2_X1 U14842 ( .A1(n16021), .A2(n7413), .ZN(n12908) );
  NAND2_X1 U14843 ( .A1(n12921), .A2(n15765), .ZN(n12907) );
  NAND2_X1 U14844 ( .A1(n12908), .A2(n12907), .ZN(n12910) );
  NAND2_X1 U14845 ( .A1(n12909), .A2(n12910), .ZN(n15655) );
  NAND2_X1 U14846 ( .A1(n15654), .A2(n15655), .ZN(n12913) );
  INV_X1 U14847 ( .A(n12909), .ZN(n12912) );
  INV_X1 U14848 ( .A(n12910), .ZN(n12911) );
  NAND2_X1 U14849 ( .A1(n12912), .A2(n12911), .ZN(n15656) );
  NAND2_X1 U14850 ( .A1(n15531), .A2(n11544), .ZN(n12917) );
  OR2_X1 U14851 ( .A1(n10704), .A2(n16123), .ZN(n12916) );
  NAND2_X1 U14852 ( .A1(n15819), .A2(n7412), .ZN(n12919) );
  NAND2_X1 U14853 ( .A1(n7413), .A2(n15838), .ZN(n12918) );
  NAND2_X1 U14854 ( .A1(n12919), .A2(n12918), .ZN(n12920) );
  XNOR2_X1 U14855 ( .A(n12920), .B(n10817), .ZN(n12925) );
  NAND2_X1 U14856 ( .A1(n15819), .A2(n7413), .ZN(n12923) );
  NAND2_X1 U14857 ( .A1(n12921), .A2(n15838), .ZN(n12922) );
  NAND2_X1 U14858 ( .A1(n12923), .A2(n12922), .ZN(n12924) );
  NOR2_X1 U14859 ( .A1(n12925), .A2(n12924), .ZN(n12926) );
  AOI21_X1 U14860 ( .B1(n12925), .B2(n12924), .A(n12926), .ZN(n15550) );
  NAND2_X1 U14861 ( .A1(n12945), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n12939) );
  INV_X1 U14862 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n12928) );
  OR2_X1 U14863 ( .A1(n12929), .A2(n12928), .ZN(n12938) );
  INV_X1 U14864 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n12930) );
  OAI21_X1 U14865 ( .B1(n12931), .B2(n15552), .A(n12930), .ZN(n12934) );
  INV_X1 U14866 ( .A(n12931), .ZN(n12933) );
  AND2_X1 U14867 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n12932) );
  NAND2_X1 U14868 ( .A1(n12933), .A2(n12932), .ZN(n15789) );
  NAND2_X1 U14869 ( .A1(n12934), .A2(n15789), .ZN(n15805) );
  OR2_X1 U14870 ( .A1(n12946), .A2(n15805), .ZN(n12937) );
  INV_X1 U14871 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n12935) );
  OR2_X1 U14872 ( .A1(n10418), .A2(n12935), .ZN(n12936) );
  OAI22_X1 U14873 ( .A1(n15808), .A2(n12940), .B1(n15815), .B2(n10271), .ZN(
        n12941) );
  XNOR2_X1 U14874 ( .A(n12941), .B(n10817), .ZN(n12943) );
  OAI22_X1 U14875 ( .A1(n15808), .A2(n10271), .B1(n15815), .B2(n12846), .ZN(
        n12942) );
  INV_X1 U14876 ( .A(n15808), .ZN(n16011) );
  AOI22_X1 U14877 ( .A1(n15659), .A2(n15838), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n12953) );
  NAND2_X1 U14878 ( .A1(n12945), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n12951) );
  NAND2_X1 U14879 ( .A1(n7420), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n12950) );
  OR2_X1 U14880 ( .A1(n12946), .A2(n15789), .ZN(n12949) );
  INV_X1 U14881 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n12947) );
  OR2_X1 U14882 ( .A1(n10418), .A2(n12947), .ZN(n12948) );
  NAND4_X1 U14883 ( .A1(n12951), .A2(n12950), .A3(n12949), .A4(n12948), .ZN(
        n15800) );
  NAND2_X1 U14884 ( .A1(n15658), .A2(n15800), .ZN(n12952) );
  OAI211_X1 U14885 ( .C1(n16535), .C2(n15805), .A(n12953), .B(n12952), .ZN(
        n12954) );
  AOI21_X1 U14886 ( .B1(n16011), .B2(n15671), .A(n12954), .ZN(n12955) );
  OAI21_X1 U14887 ( .B1(n12956), .B2(n15673), .A(n12955), .ZN(P1_U3220) );
  NAND2_X1 U14888 ( .A1(n12957), .A2(n12053), .ZN(n12960) );
  OR2_X1 U14889 ( .A1(n9783), .A2(n12958), .ZN(n12959) );
  XNOR2_X1 U14890 ( .A(n15291), .B(n14936), .ZN(n12978) );
  INV_X1 U14891 ( .A(n12978), .ZN(n12980) );
  INV_X1 U14892 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n12961) );
  NAND2_X1 U14893 ( .A1(n12962), .A2(n12961), .ZN(n12963) );
  AND2_X1 U14894 ( .A1(n12985), .A2(n12963), .ZN(n15293) );
  NAND2_X1 U14895 ( .A1(n15293), .A2(n9786), .ZN(n12968) );
  INV_X1 U14896 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n15431) );
  NAND2_X1 U14897 ( .A1(n10847), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n12965) );
  NAND2_X1 U14898 ( .A1(n9789), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n12964) );
  OAI211_X1 U14899 ( .C1(n15431), .C2(n13265), .A(n12965), .B(n12964), .ZN(
        n12966) );
  INV_X1 U14900 ( .A(n12966), .ZN(n12967) );
  NAND2_X1 U14901 ( .A1(n12968), .A2(n12967), .ZN(n15267) );
  NAND2_X1 U14902 ( .A1(n15267), .A2(n14937), .ZN(n12979) );
  NAND2_X1 U14903 ( .A1(n15320), .A2(n14937), .ZN(n12976) );
  NAND2_X1 U14904 ( .A1(n12969), .A2(n12053), .ZN(n12972) );
  OR2_X1 U14905 ( .A1(n9783), .A2(n12970), .ZN(n12971) );
  XOR2_X1 U14906 ( .A(n12976), .B(n12975), .Z(n14999) );
  INV_X1 U14907 ( .A(n12973), .ZN(n12974) );
  INV_X1 U14908 ( .A(n12975), .ZN(n12977) );
  XNOR2_X1 U14909 ( .A(n12978), .B(n12979), .ZN(n14969) );
  NAND2_X1 U14910 ( .A1(n12981), .A2(n12053), .ZN(n12983) );
  OR2_X1 U14911 ( .A1(n9783), .A2(n7827), .ZN(n12982) );
  NAND2_X2 U14912 ( .A1(n12983), .A2(n12982), .ZN(n15424) );
  INV_X1 U14913 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n12984) );
  NAND2_X1 U14914 ( .A1(n12985), .A2(n12984), .ZN(n12986) );
  NAND2_X1 U14915 ( .A1(n12996), .A2(n12986), .ZN(n15271) );
  OR2_X1 U14916 ( .A1(n15271), .A2(n13262), .ZN(n12992) );
  INV_X1 U14917 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n12989) );
  NAND2_X1 U14918 ( .A1(n9789), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n12988) );
  NAND2_X1 U14919 ( .A1(n10847), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n12987) );
  OAI211_X1 U14920 ( .C1(n13265), .C2(n12989), .A(n12988), .B(n12987), .ZN(
        n12990) );
  INV_X1 U14921 ( .A(n12990), .ZN(n12991) );
  NAND2_X1 U14922 ( .A1(n15145), .A2(n14937), .ZN(n12993) );
  AOI22_X1 U14923 ( .A1(n7507), .A2(n15014), .B1(n14961), .B2(n15145), .ZN(
        n13008) );
  INV_X1 U14924 ( .A(n15267), .ZN(n15153) );
  NOR2_X1 U14925 ( .A1(n15153), .A2(n12994), .ZN(n13006) );
  NAND2_X1 U14926 ( .A1(n12996), .A2(n12995), .ZN(n12997) );
  AND2_X1 U14927 ( .A1(n13167), .A2(n12997), .ZN(n15259) );
  NAND2_X1 U14928 ( .A1(n15259), .A2(n9786), .ZN(n13002) );
  INV_X1 U14929 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n15421) );
  NAND2_X1 U14930 ( .A1(n9789), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n12999) );
  NAND2_X1 U14931 ( .A1(n9788), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n12998) );
  OAI211_X1 U14932 ( .C1(n13265), .C2(n15421), .A(n12999), .B(n12998), .ZN(
        n13000) );
  INV_X1 U14933 ( .A(n13000), .ZN(n13001) );
  INV_X1 U14934 ( .A(n15266), .ZN(n15157) );
  INV_X1 U14935 ( .A(n15271), .ZN(n13003) );
  AOI22_X1 U14936 ( .A1(n13003), .A2(n15018), .B1(P2_REG3_REG_22__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13004) );
  OAI21_X1 U14937 ( .B1(n15157), .B2(n14972), .A(n13004), .ZN(n13005) );
  AOI211_X1 U14938 ( .C1(n15424), .C2(n15024), .A(n13006), .B(n13005), .ZN(
        n13007) );
  OAI21_X1 U14939 ( .B1(n14922), .B2(n13008), .A(n13007), .ZN(P2_U3207) );
  NAND2_X1 U14940 ( .A1(n13013), .A2(n13012), .ZN(n13010) );
  INV_X1 U14941 ( .A(n13340), .ZN(n13009) );
  NAND2_X1 U14942 ( .A1(n13010), .A2(n8850), .ZN(n13014) );
  NAND2_X1 U14943 ( .A1(n13015), .A2(n8104), .ZN(n13016) );
  INV_X2 U14944 ( .A(n13302), .ZN(n13239) );
  NAND2_X1 U14945 ( .A1(n15043), .A2(n13239), .ZN(n13018) );
  NAND2_X1 U14946 ( .A1(n8104), .A2(n13024), .ZN(n13017) );
  NAND2_X1 U14947 ( .A1(n13018), .A2(n13017), .ZN(n13026) );
  NAND2_X1 U14948 ( .A1(n13239), .A2(n13021), .ZN(n13020) );
  NAND2_X1 U14949 ( .A1(n15042), .A2(n8104), .ZN(n13019) );
  NAND2_X1 U14950 ( .A1(n15042), .A2(n13239), .ZN(n13023) );
  NAND2_X1 U14951 ( .A1(n8104), .A2(n13021), .ZN(n13022) );
  NAND2_X1 U14952 ( .A1(n13023), .A2(n13022), .ZN(n13028) );
  OAI22_X1 U14953 ( .A1(n13027), .A2(n13026), .B1(n13029), .B2(n13028), .ZN(
        n13032) );
  AOI22_X1 U14954 ( .A1(n15043), .A2(n8104), .B1(n13239), .B2(n13024), .ZN(
        n13025) );
  AOI21_X1 U14955 ( .B1(n13027), .B2(n13026), .A(n13025), .ZN(n13031) );
  NAND2_X1 U14956 ( .A1(n13029), .A2(n13028), .ZN(n13030) );
  NAND2_X1 U14957 ( .A1(n15041), .A2(n13160), .ZN(n13034) );
  NAND2_X1 U14958 ( .A1(n8104), .A2(n13035), .ZN(n13033) );
  NAND2_X1 U14959 ( .A1(n13034), .A2(n13033), .ZN(n13041) );
  NAND2_X1 U14960 ( .A1(n13040), .A2(n13041), .ZN(n13039) );
  NAND2_X1 U14961 ( .A1(n15041), .A2(n8104), .ZN(n13037) );
  NAND2_X1 U14962 ( .A1(n13160), .A2(n13035), .ZN(n13036) );
  NAND2_X1 U14963 ( .A1(n13037), .A2(n13036), .ZN(n13038) );
  NAND2_X1 U14964 ( .A1(n13039), .A2(n13038), .ZN(n13045) );
  INV_X1 U14965 ( .A(n13040), .ZN(n13043) );
  INV_X1 U14966 ( .A(n13041), .ZN(n13042) );
  NAND2_X1 U14967 ( .A1(n13043), .A2(n13042), .ZN(n13044) );
  NAND2_X1 U14968 ( .A1(n13045), .A2(n13044), .ZN(n13051) );
  NAND2_X1 U14969 ( .A1(n15040), .A2(n8104), .ZN(n13047) );
  NAND2_X1 U14970 ( .A1(n13160), .A2(n13048), .ZN(n13046) );
  NAND2_X1 U14971 ( .A1(n13047), .A2(n13046), .ZN(n13050) );
  AOI22_X1 U14972 ( .A1(n13160), .A2(n15040), .B1(n8104), .B2(n13048), .ZN(
        n13049) );
  NAND2_X1 U14973 ( .A1(n13054), .A2(n13299), .ZN(n13053) );
  NAND2_X1 U14974 ( .A1(n15039), .A2(n13160), .ZN(n13052) );
  NAND2_X1 U14975 ( .A1(n13053), .A2(n13052), .ZN(n13056) );
  AOI22_X1 U14976 ( .A1(n13160), .A2(n13054), .B1(n15039), .B2(n13299), .ZN(
        n13055) );
  AOI22_X1 U14977 ( .A1(n16586), .A2(n13239), .B1(n15038), .B2(n13299), .ZN(
        n13059) );
  NAND2_X1 U14978 ( .A1(n16586), .A2(n13299), .ZN(n13057) );
  AND2_X1 U14979 ( .A1(n15037), .A2(n13239), .ZN(n13061) );
  AOI21_X1 U14980 ( .B1(n13062), .B2(n13299), .A(n13061), .ZN(n13066) );
  NAND2_X1 U14981 ( .A1(n13067), .A2(n13066), .ZN(n13068) );
  NAND2_X1 U14982 ( .A1(n13062), .A2(n13160), .ZN(n13063) );
  OAI21_X1 U14983 ( .B1(n13064), .B2(n13160), .A(n13063), .ZN(n13065) );
  NAND2_X1 U14984 ( .A1(n13071), .A2(n13239), .ZN(n13070) );
  NAND2_X1 U14985 ( .A1(n15036), .A2(n13299), .ZN(n13069) );
  NAND2_X1 U14986 ( .A1(n13070), .A2(n13069), .ZN(n13073) );
  AOI22_X1 U14987 ( .A1(n13071), .A2(n13299), .B1(n13239), .B2(n15036), .ZN(
        n13072) );
  NAND2_X1 U14988 ( .A1(n13077), .A2(n13299), .ZN(n13076) );
  NAND2_X1 U14989 ( .A1(n15035), .A2(n13239), .ZN(n13075) );
  NAND2_X1 U14990 ( .A1(n13077), .A2(n13160), .ZN(n13078) );
  OAI21_X1 U14991 ( .B1(n13079), .B2(n13160), .A(n13078), .ZN(n13080) );
  NAND2_X1 U14992 ( .A1(n13083), .A2(n13160), .ZN(n13082) );
  NAND2_X1 U14993 ( .A1(n15034), .A2(n13299), .ZN(n13081) );
  AOI22_X1 U14994 ( .A1(n13083), .A2(n13299), .B1(n13239), .B2(n15034), .ZN(
        n13084) );
  NAND2_X1 U14995 ( .A1(n15368), .A2(n13299), .ZN(n13087) );
  NAND2_X1 U14996 ( .A1(n15033), .A2(n13239), .ZN(n13086) );
  NAND2_X1 U14997 ( .A1(n13087), .A2(n13086), .ZN(n13093) );
  NAND2_X1 U14998 ( .A1(n13092), .A2(n13093), .ZN(n13091) );
  NAND2_X1 U14999 ( .A1(n15368), .A2(n13160), .ZN(n13088) );
  OAI21_X1 U15000 ( .B1(n13089), .B2(n13160), .A(n13088), .ZN(n13090) );
  INV_X1 U15001 ( .A(n13093), .ZN(n13094) );
  NAND2_X1 U15002 ( .A1(n13095), .A2(n13094), .ZN(n13096) );
  NAND2_X1 U15003 ( .A1(n16700), .A2(n13239), .ZN(n13098) );
  NAND2_X1 U15004 ( .A1(n15032), .A2(n13299), .ZN(n13097) );
  AOI22_X1 U15005 ( .A1(n16700), .A2(n13299), .B1(n13239), .B2(n15032), .ZN(
        n13099) );
  NAND2_X1 U15006 ( .A1(n13102), .A2(n13299), .ZN(n13101) );
  NAND2_X1 U15007 ( .A1(n15031), .A2(n13239), .ZN(n13100) );
  NAND2_X1 U15008 ( .A1(n13101), .A2(n13100), .ZN(n13104) );
  AOI22_X1 U15009 ( .A1(n13102), .A2(n13160), .B1(n15031), .B2(n13299), .ZN(
        n13103) );
  NAND2_X1 U15010 ( .A1(n16741), .A2(n13160), .ZN(n13106) );
  NAND2_X1 U15011 ( .A1(n15030), .A2(n13299), .ZN(n13105) );
  NAND2_X1 U15012 ( .A1(n13106), .A2(n13105), .ZN(n13110) );
  NAND2_X1 U15013 ( .A1(n16741), .A2(n13299), .ZN(n13108) );
  NAND2_X1 U15014 ( .A1(n15030), .A2(n13239), .ZN(n13107) );
  NAND2_X1 U15015 ( .A1(n13108), .A2(n13107), .ZN(n13109) );
  NAND2_X1 U15016 ( .A1(n13113), .A2(n13299), .ZN(n13112) );
  NAND2_X1 U15017 ( .A1(n15029), .A2(n13160), .ZN(n13111) );
  NAND2_X1 U15018 ( .A1(n13112), .A2(n13111), .ZN(n13115) );
  AOI22_X1 U15019 ( .A1(n13113), .A2(n13160), .B1(n15029), .B2(n13299), .ZN(
        n13114) );
  NAND2_X1 U15020 ( .A1(n15511), .A2(n13239), .ZN(n13118) );
  NAND2_X1 U15021 ( .A1(n15028), .A2(n13299), .ZN(n13117) );
  NAND2_X1 U15022 ( .A1(n13118), .A2(n13117), .ZN(n13122) );
  NAND2_X1 U15023 ( .A1(n15511), .A2(n13299), .ZN(n13119) );
  NAND2_X1 U15024 ( .A1(n8008), .A2(n13299), .ZN(n13124) );
  NAND2_X1 U15025 ( .A1(n15342), .A2(n13239), .ZN(n13123) );
  NAND2_X1 U15026 ( .A1(n13124), .A2(n13123), .ZN(n13126) );
  AOI22_X1 U15027 ( .A1(n8008), .A2(n13239), .B1(n15342), .B2(n13299), .ZN(
        n13125) );
  AOI21_X1 U15028 ( .B1(n13127), .B2(n13126), .A(n13125), .ZN(n13128) );
  NAND2_X1 U15029 ( .A1(n15444), .A2(n13239), .ZN(n13130) );
  NAND2_X1 U15030 ( .A1(n15319), .A2(n13299), .ZN(n13129) );
  NAND2_X1 U15031 ( .A1(n13130), .A2(n13129), .ZN(n13131) );
  NAND2_X1 U15032 ( .A1(n15444), .A2(n13299), .ZN(n13133) );
  NAND2_X1 U15033 ( .A1(n15319), .A2(n13160), .ZN(n13132) );
  NAND2_X1 U15034 ( .A1(n13133), .A2(n13132), .ZN(n13134) );
  NAND2_X1 U15035 ( .A1(n15329), .A2(n13299), .ZN(n13136) );
  NAND2_X1 U15036 ( .A1(n15344), .A2(n13160), .ZN(n13135) );
  NAND2_X1 U15037 ( .A1(n13136), .A2(n13135), .ZN(n13138) );
  AOI22_X1 U15038 ( .A1(n15329), .A2(n13239), .B1(n15344), .B2(n13299), .ZN(
        n13137) );
  NAND2_X1 U15039 ( .A1(n15304), .A2(n13239), .ZN(n13140) );
  NAND2_X1 U15040 ( .A1(n15320), .A2(n13299), .ZN(n13139) );
  NAND2_X1 U15041 ( .A1(n13140), .A2(n13139), .ZN(n13142) );
  AOI22_X1 U15042 ( .A1(n15304), .A2(n13299), .B1(n13160), .B2(n15320), .ZN(
        n13141) );
  NAND2_X1 U15043 ( .A1(n15291), .A2(n13299), .ZN(n13144) );
  NAND2_X1 U15044 ( .A1(n15267), .A2(n13160), .ZN(n13143) );
  NAND2_X1 U15045 ( .A1(n13144), .A2(n13143), .ZN(n13148) );
  NAND2_X1 U15046 ( .A1(n15291), .A2(n13239), .ZN(n13145) );
  OAI21_X1 U15047 ( .B1(n15153), .B2(n13160), .A(n13145), .ZN(n13146) );
  NAND2_X1 U15048 ( .A1(n15424), .A2(n13160), .ZN(n13152) );
  NAND2_X1 U15049 ( .A1(n15145), .A2(n13299), .ZN(n13151) );
  AOI22_X1 U15050 ( .A1(n15424), .A2(n13299), .B1(n13239), .B2(n15145), .ZN(
        n13153) );
  NAND2_X1 U15051 ( .A1(n16136), .A2(n12053), .ZN(n13156) );
  OR2_X1 U15052 ( .A1(n9783), .A2(n8582), .ZN(n13155) );
  NAND2_X1 U15053 ( .A1(n15256), .A2(n13299), .ZN(n13158) );
  NAND2_X1 U15054 ( .A1(n15266), .A2(n13160), .ZN(n13157) );
  NAND2_X1 U15055 ( .A1(n13158), .A2(n13157), .ZN(n13163) );
  NAND2_X1 U15056 ( .A1(n15256), .A2(n13239), .ZN(n13159) );
  OAI21_X1 U15057 ( .B1(n15157), .B2(n13160), .A(n13159), .ZN(n13161) );
  NAND2_X1 U15058 ( .A1(n13162), .A2(n13161), .ZN(n13164) );
  NAND2_X1 U15059 ( .A1(n15538), .A2(n12053), .ZN(n13166) );
  OR2_X1 U15060 ( .A1(n9783), .A2(n15541), .ZN(n13165) );
  NAND2_X2 U15061 ( .A1(n13166), .A2(n13165), .ZN(n15414) );
  NAND2_X1 U15062 ( .A1(n15414), .A2(n13239), .ZN(n13176) );
  INV_X1 U15063 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n14989) );
  NAND2_X1 U15064 ( .A1(n13167), .A2(n14989), .ZN(n13168) );
  NAND2_X1 U15065 ( .A1(n13180), .A2(n13168), .ZN(n15242) );
  INV_X1 U15066 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n13171) );
  NAND2_X1 U15067 ( .A1(n9788), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n13170) );
  NAND2_X1 U15068 ( .A1(n9789), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n13169) );
  OAI211_X1 U15069 ( .C1(n13265), .C2(n13171), .A(n13170), .B(n13169), .ZN(
        n13172) );
  INV_X1 U15070 ( .A(n13172), .ZN(n13173) );
  NAND2_X1 U15071 ( .A1(n15132), .A2(n13299), .ZN(n13175) );
  AOI22_X1 U15072 ( .A1(n15414), .A2(n13299), .B1(n13239), .B2(n15132), .ZN(
        n13177) );
  NAND2_X1 U15073 ( .A1(n15535), .A2(n12053), .ZN(n13179) );
  OR2_X1 U15074 ( .A1(n9783), .A2(n15537), .ZN(n13178) );
  NAND2_X2 U15075 ( .A1(n13179), .A2(n13178), .ZN(n15408) );
  NAND2_X1 U15076 ( .A1(n15408), .A2(n13299), .ZN(n13189) );
  INV_X1 U15077 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n14982) );
  NAND2_X1 U15078 ( .A1(n13180), .A2(n14982), .ZN(n13181) );
  NAND2_X1 U15079 ( .A1(n13201), .A2(n13181), .ZN(n15230) );
  OR2_X1 U15080 ( .A1(n15230), .A2(n13262), .ZN(n13187) );
  INV_X1 U15081 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n13184) );
  NAND2_X1 U15082 ( .A1(n9789), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n13183) );
  NAND2_X1 U15083 ( .A1(n10847), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n13182) );
  OAI211_X1 U15084 ( .C1(n13265), .C2(n13184), .A(n13183), .B(n13182), .ZN(
        n13185) );
  INV_X1 U15085 ( .A(n13185), .ZN(n13186) );
  NAND2_X1 U15086 ( .A1(n13187), .A2(n13186), .ZN(n15134) );
  NAND2_X1 U15087 ( .A1(n15134), .A2(n13239), .ZN(n13188) );
  NAND2_X1 U15088 ( .A1(n13189), .A2(n13188), .ZN(n13191) );
  AOI22_X1 U15089 ( .A1(n15408), .A2(n13160), .B1(n15134), .B2(n13299), .ZN(
        n13190) );
  NOR2_X1 U15090 ( .A1(n13192), .A2(n13191), .ZN(n13213) );
  NAND2_X1 U15091 ( .A1(n15531), .A2(n12053), .ZN(n13194) );
  OR2_X1 U15092 ( .A1(n9783), .A2(n10579), .ZN(n13193) );
  AND2_X1 U15093 ( .A1(n15017), .A2(n13299), .ZN(n13195) );
  AOI21_X1 U15094 ( .B1(n15195), .B2(n13160), .A(n13195), .ZN(n13273) );
  NAND2_X1 U15095 ( .A1(n15195), .A2(n13299), .ZN(n13197) );
  NAND2_X1 U15096 ( .A1(n15017), .A2(n13239), .ZN(n13196) );
  NAND2_X1 U15097 ( .A1(n13197), .A2(n13196), .ZN(n13272) );
  NAND2_X1 U15098 ( .A1(n13273), .A2(n13272), .ZN(n13280) );
  NAND2_X1 U15099 ( .A1(n15532), .A2(n12053), .ZN(n13199) );
  OR2_X1 U15100 ( .A1(n9783), .A2(n15533), .ZN(n13198) );
  NAND2_X1 U15101 ( .A1(n13201), .A2(n13200), .ZN(n13202) );
  NAND2_X1 U15102 ( .A1(n15214), .A2(n9786), .ZN(n13208) );
  INV_X1 U15103 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n13205) );
  NAND2_X1 U15104 ( .A1(n10847), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n13204) );
  NAND2_X1 U15105 ( .A1(n9789), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n13203) );
  OAI211_X1 U15106 ( .C1(n13205), .C2(n13265), .A(n13204), .B(n13203), .ZN(
        n13206) );
  INV_X1 U15107 ( .A(n13206), .ZN(n13207) );
  AND2_X1 U15108 ( .A1(n15162), .A2(n13299), .ZN(n13209) );
  AOI21_X1 U15109 ( .B1(n15211), .B2(n13239), .A(n13209), .ZN(n13277) );
  NAND2_X1 U15110 ( .A1(n15211), .A2(n13299), .ZN(n13211) );
  NAND2_X1 U15111 ( .A1(n15162), .A2(n13160), .ZN(n13210) );
  NAND2_X1 U15112 ( .A1(n13211), .A2(n13210), .ZN(n13276) );
  NAND2_X1 U15113 ( .A1(n13277), .A2(n13276), .ZN(n13212) );
  INV_X1 U15114 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n16121) );
  MUX2_X1 U15115 ( .A(n16121), .B(n15525), .S(n7416), .Z(n13244) );
  XNOR2_X1 U15116 ( .A(n13244), .B(SI_30_), .ZN(n13243) );
  NAND2_X1 U15117 ( .A1(n15524), .A2(n12053), .ZN(n13219) );
  OR2_X1 U15118 ( .A1(n9783), .A2(n15525), .ZN(n13218) );
  INV_X1 U15119 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n15382) );
  NAND2_X1 U15120 ( .A1(n9789), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n13221) );
  NAND2_X1 U15121 ( .A1(n10847), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n13220) );
  OAI211_X1 U15122 ( .C1(n13265), .C2(n15382), .A(n13221), .B(n13220), .ZN(
        n15169) );
  AND2_X1 U15123 ( .A1(n15169), .A2(n13239), .ZN(n13222) );
  AOI21_X1 U15124 ( .B1(n15110), .B2(n13299), .A(n13222), .ZN(n13294) );
  NAND2_X1 U15125 ( .A1(n15110), .A2(n13160), .ZN(n13228) );
  NAND2_X1 U15126 ( .A1(n13299), .A2(n15114), .ZN(n13225) );
  NAND2_X1 U15127 ( .A1(n13223), .A2(n8082), .ZN(n13343) );
  NAND3_X1 U15128 ( .A1(n13225), .A2(n13224), .A3(n13342), .ZN(n13226) );
  NAND2_X1 U15129 ( .A1(n13226), .A2(n15169), .ZN(n13227) );
  NAND2_X1 U15130 ( .A1(n13228), .A2(n13227), .ZN(n13293) );
  NAND2_X1 U15131 ( .A1(n13599), .A2(n12053), .ZN(n13230) );
  OR2_X1 U15132 ( .A1(n9783), .A2(n13493), .ZN(n13229) );
  INV_X1 U15133 ( .A(n13260), .ZN(n13232) );
  AND2_X1 U15134 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(P2_REG3_REG_28__SCAN_IN), 
        .ZN(n13231) );
  NAND2_X1 U15135 ( .A1(n13232), .A2(n13231), .ZN(n15140) );
  OR2_X1 U15136 ( .A1(n15140), .A2(n13262), .ZN(n13238) );
  INV_X1 U15137 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n13235) );
  NAND2_X1 U15138 ( .A1(n9789), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n13234) );
  NAND2_X1 U15139 ( .A1(n9788), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n13233) );
  OAI211_X1 U15140 ( .C1(n13265), .C2(n13235), .A(n13234), .B(n13233), .ZN(
        n13236) );
  INV_X1 U15141 ( .A(n13236), .ZN(n13237) );
  NAND2_X1 U15142 ( .A1(n13238), .A2(n13237), .ZN(n15027) );
  AND2_X1 U15143 ( .A1(n15027), .A2(n13239), .ZN(n13240) );
  AOI21_X1 U15144 ( .B1(n15386), .B2(n13299), .A(n13240), .ZN(n13291) );
  NAND2_X1 U15145 ( .A1(n15386), .A2(n13239), .ZN(n13242) );
  NAND2_X1 U15146 ( .A1(n15027), .A2(n13299), .ZN(n13241) );
  NAND2_X1 U15147 ( .A1(n13242), .A2(n13241), .ZN(n13290) );
  AOI22_X1 U15148 ( .A1(n13294), .A2(n13293), .B1(n13291), .B2(n13290), .ZN(
        n13254) );
  INV_X1 U15149 ( .A(n13243), .ZN(n13245) );
  MUX2_X1 U15150 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n7416), .Z(n13248) );
  XNOR2_X1 U15151 ( .A(n13248), .B(SI_31_), .ZN(n13249) );
  NAND2_X1 U15152 ( .A1(n15519), .A2(n12053), .ZN(n13252) );
  OR2_X1 U15153 ( .A1(n9783), .A2(n13500), .ZN(n13251) );
  INV_X1 U15154 ( .A(n15114), .ZN(n13300) );
  NAND2_X1 U15155 ( .A1(n15111), .A2(n13300), .ZN(n13298) );
  OR2_X1 U15156 ( .A1(n15111), .A2(n13300), .ZN(n13253) );
  OR2_X1 U15157 ( .A1(n9783), .A2(n13256), .ZN(n13257) );
  INV_X1 U15158 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n13259) );
  INV_X1 U15159 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n14964) );
  OAI21_X1 U15160 ( .B1(n13260), .B2(n13259), .A(n14964), .ZN(n13261) );
  NAND2_X1 U15161 ( .A1(n15140), .A2(n13261), .ZN(n15182) );
  INV_X1 U15162 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n15393) );
  NAND2_X1 U15163 ( .A1(n10847), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n13264) );
  NAND2_X1 U15164 ( .A1(n9789), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n13263) );
  OAI211_X1 U15165 ( .C1(n15393), .C2(n13265), .A(n13264), .B(n13263), .ZN(
        n13266) );
  INV_X1 U15166 ( .A(n13266), .ZN(n13267) );
  NAND2_X1 U15167 ( .A1(n13268), .A2(n13267), .ZN(n15137) );
  AND2_X1 U15168 ( .A1(n15137), .A2(n13299), .ZN(n13269) );
  AOI21_X1 U15169 ( .B1(n15184), .B2(n13239), .A(n13269), .ZN(n13287) );
  NAND2_X1 U15170 ( .A1(n15184), .A2(n13299), .ZN(n13271) );
  NAND2_X1 U15171 ( .A1(n15137), .A2(n13160), .ZN(n13270) );
  NAND2_X1 U15172 ( .A1(n13271), .A2(n13270), .ZN(n13286) );
  INV_X1 U15173 ( .A(n13272), .ZN(n13275) );
  INV_X1 U15174 ( .A(n13273), .ZN(n13274) );
  NAND2_X1 U15175 ( .A1(n13275), .A2(n13274), .ZN(n13282) );
  INV_X1 U15176 ( .A(n13276), .ZN(n13279) );
  INV_X1 U15177 ( .A(n13277), .ZN(n13278) );
  NAND3_X1 U15178 ( .A1(n13280), .A2(n13279), .A3(n13278), .ZN(n13281) );
  OAI211_X1 U15179 ( .C1(n13287), .C2(n13286), .A(n13282), .B(n13281), .ZN(
        n13283) );
  INV_X1 U15180 ( .A(n13283), .ZN(n13284) );
  INV_X1 U15181 ( .A(n13286), .ZN(n13289) );
  INV_X1 U15182 ( .A(n13287), .ZN(n13288) );
  OAI22_X1 U15183 ( .A1(n13291), .A2(n13290), .B1(n13289), .B2(n13288), .ZN(
        n13292) );
  INV_X1 U15184 ( .A(n13293), .ZN(n13296) );
  INV_X1 U15185 ( .A(n13294), .ZN(n13295) );
  NAND2_X1 U15186 ( .A1(n13296), .A2(n13295), .ZN(n13297) );
  INV_X1 U15187 ( .A(n13298), .ZN(n13303) );
  NOR2_X1 U15188 ( .A1(n13300), .A2(n13299), .ZN(n13301) );
  AOI22_X1 U15189 ( .A1(n13303), .A2(n8104), .B1(n13301), .B2(n15468), .ZN(
        n13304) );
  INV_X1 U15190 ( .A(n15137), .ZN(n15172) );
  NAND2_X1 U15191 ( .A1(n15184), .A2(n15172), .ZN(n13305) );
  NAND2_X1 U15192 ( .A1(n15166), .A2(n13305), .ZN(n15165) );
  INV_X1 U15193 ( .A(n15017), .ZN(n15163) );
  XNOR2_X1 U15194 ( .A(n15195), .B(n15163), .ZN(n15193) );
  INV_X1 U15195 ( .A(n15162), .ZN(n15136) );
  XNOR2_X1 U15196 ( .A(n15211), .B(n15136), .ZN(n15209) );
  XNOR2_X1 U15197 ( .A(n15408), .B(n15134), .ZN(n15220) );
  XNOR2_X1 U15198 ( .A(n15304), .B(n15288), .ZN(n15299) );
  XNOR2_X1 U15199 ( .A(n15291), .B(n15153), .ZN(n15284) );
  OR2_X1 U15200 ( .A1(n15329), .A2(n14995), .ZN(n15151) );
  NAND2_X1 U15201 ( .A1(n15329), .A2(n14995), .ZN(n13306) );
  AND2_X2 U15202 ( .A1(n15151), .A2(n13306), .ZN(n15324) );
  NAND4_X1 U15203 ( .A1(n13310), .A2(n13309), .A3(n13308), .A4(n13307), .ZN(
        n13313) );
  NOR3_X1 U15204 ( .A1(n13313), .A2(n13312), .A3(n13311), .ZN(n13316) );
  NAND4_X1 U15205 ( .A1(n13317), .A2(n13316), .A3(n13315), .A4(n13314), .ZN(
        n13318) );
  OR4_X1 U15206 ( .A1(n13321), .A2(n13320), .A3(n13319), .A4(n13318), .ZN(
        n13323) );
  OR4_X1 U15207 ( .A1(n13325), .A2(n13324), .A3(n13323), .A4(n13322), .ZN(
        n13326) );
  NOR4_X1 U15208 ( .A1(n13329), .A2(n13328), .A3(n13327), .A4(n13326), .ZN(
        n13330) );
  XNOR2_X1 U15209 ( .A(n15444), .B(n15319), .ZN(n15339) );
  NAND4_X1 U15210 ( .A1(n15324), .A2(n13330), .A3(n15148), .A4(n15339), .ZN(
        n13331) );
  NOR4_X1 U15211 ( .A1(n15269), .A2(n15299), .A3(n15284), .A4(n13331), .ZN(
        n13332) );
  XNOR2_X1 U15212 ( .A(n15256), .B(n15266), .ZN(n15254) );
  NAND4_X1 U15213 ( .A1(n15220), .A2(n13332), .A3(n15239), .A4(n15254), .ZN(
        n13333) );
  XNOR2_X1 U15214 ( .A(n15386), .B(n15027), .ZN(n15167) );
  XNOR2_X1 U15215 ( .A(n15110), .B(n15169), .ZN(n13334) );
  NAND2_X1 U15216 ( .A1(n13342), .A2(n13338), .ZN(n13339) );
  OAI211_X1 U15217 ( .C1(n13340), .C2(n8082), .A(n13351), .B(n13339), .ZN(
        n13348) );
  NAND2_X1 U15218 ( .A1(n13342), .A2(n13341), .ZN(n13344) );
  OAI21_X1 U15219 ( .B1(n13345), .B2(n13344), .A(n13343), .ZN(n13347) );
  OR2_X1 U15220 ( .A1(n13350), .A2(P2_U3088), .ZN(n15543) );
  NOR4_X1 U15221 ( .A1(n16152), .A2(n10090), .A3(n13351), .A4(n15289), .ZN(
        n13353) );
  OAI21_X1 U15222 ( .B1(n15543), .B2(n8082), .A(P2_B_REG_SCAN_IN), .ZN(n13352)
         );
  OAI22_X1 U15223 ( .A1(n13354), .A2(n15543), .B1(n13353), .B2(n13352), .ZN(
        P2_U3328) );
  MUX2_X1 U15224 ( .A(n13356), .B(n13355), .S(n13491), .Z(n13488) );
  INV_X1 U15225 ( .A(n13363), .ZN(n13373) );
  OAI21_X1 U15226 ( .B1(n16499), .B2(n13359), .A(n16491), .ZN(n13367) );
  AOI21_X1 U15227 ( .B1(n13362), .B2(n13361), .A(n13360), .ZN(n13365) );
  OAI211_X1 U15228 ( .C1(n13365), .C2(n16499), .A(n13364), .B(n13363), .ZN(
        n13366) );
  MUX2_X1 U15229 ( .A(n13367), .B(n13366), .S(n13480), .Z(n13371) );
  AOI21_X1 U15230 ( .B1(n13370), .B2(n13368), .A(n13480), .ZN(n13369) );
  AOI21_X1 U15231 ( .B1(n13371), .B2(n13370), .A(n13369), .ZN(n13372) );
  AOI21_X1 U15232 ( .B1(n13373), .B2(n13491), .A(n13372), .ZN(n13378) );
  MUX2_X1 U15233 ( .A(n13375), .B(n13374), .S(n13480), .Z(n13376) );
  OAI211_X1 U15234 ( .C1(n13378), .C2(n13377), .A(n13526), .B(n13376), .ZN(
        n13382) );
  MUX2_X1 U15235 ( .A(n13380), .B(n13379), .S(n13491), .Z(n13381) );
  NAND3_X1 U15236 ( .A1(n13382), .A2(n13532), .A3(n13381), .ZN(n13389) );
  NAND2_X1 U15237 ( .A1(n13384), .A2(n13383), .ZN(n13386) );
  MUX2_X1 U15238 ( .A(n13386), .B(n13385), .S(n13480), .Z(n13388) );
  AOI21_X1 U15239 ( .B1(n13389), .B2(n13388), .A(n13387), .ZN(n13401) );
  NAND2_X1 U15240 ( .A1(n13391), .A2(n13390), .ZN(n13393) );
  MUX2_X1 U15241 ( .A(n13393), .B(n13392), .S(n13480), .Z(n13394) );
  NAND2_X1 U15242 ( .A1(n13524), .A2(n13394), .ZN(n13400) );
  INV_X1 U15243 ( .A(n13395), .ZN(n13528) );
  NAND2_X1 U15244 ( .A1(n13396), .A2(n16614), .ZN(n13397) );
  MUX2_X1 U15245 ( .A(n13398), .B(n13397), .S(n13480), .Z(n13399) );
  OAI211_X1 U15246 ( .C1(n13401), .C2(n13400), .A(n13528), .B(n13399), .ZN(
        n13405) );
  MUX2_X1 U15247 ( .A(n13403), .B(n13402), .S(n13480), .Z(n13404) );
  NAND3_X1 U15248 ( .A1(n13405), .A2(n13538), .A3(n13404), .ZN(n13411) );
  NAND2_X1 U15249 ( .A1(n13406), .A2(n16663), .ZN(n13408) );
  MUX2_X1 U15250 ( .A(n13408), .B(n13407), .S(n13491), .Z(n13410) );
  AOI21_X1 U15251 ( .B1(n13411), .B2(n13410), .A(n13409), .ZN(n13420) );
  NAND2_X1 U15252 ( .A1(n13418), .A2(n13412), .ZN(n13413) );
  OAI21_X1 U15253 ( .B1(n13420), .B2(n13413), .A(n13417), .ZN(n13415) );
  INV_X1 U15254 ( .A(n13414), .ZN(n13539) );
  NAND2_X1 U15255 ( .A1(n13415), .A2(n13539), .ZN(n13424) );
  NAND2_X1 U15256 ( .A1(n13417), .A2(n13416), .ZN(n13419) );
  OAI21_X1 U15257 ( .B1(n13420), .B2(n13419), .A(n13418), .ZN(n13422) );
  AOI21_X1 U15258 ( .B1(n13422), .B2(n13539), .A(n13421), .ZN(n13423) );
  MUX2_X1 U15259 ( .A(n13424), .B(n13423), .S(n13491), .Z(n13433) );
  INV_X1 U15260 ( .A(n14366), .ZN(n14361) );
  OR2_X1 U15261 ( .A1(n14361), .A2(n14344), .ZN(n13541) );
  INV_X1 U15262 ( .A(n14326), .ZN(n14332) );
  AOI21_X1 U15263 ( .B1(n13426), .B2(n13425), .A(n13491), .ZN(n13428) );
  MUX2_X1 U15264 ( .A(n13491), .B(n13428), .S(n13427), .Z(n13431) );
  MUX2_X1 U15265 ( .A(n13429), .B(n14330), .S(n13491), .Z(n13430) );
  OAI21_X1 U15266 ( .B1(n13431), .B2(n14344), .A(n13430), .ZN(n13432) );
  OAI211_X1 U15267 ( .C1(n13433), .C2(n13541), .A(n14332), .B(n13432), .ZN(
        n13437) );
  MUX2_X1 U15268 ( .A(n13435), .B(n13434), .S(n13480), .Z(n13436) );
  NAND2_X1 U15269 ( .A1(n14279), .A2(n14319), .ZN(n13441) );
  AOI21_X1 U15270 ( .B1(n13437), .B2(n13436), .A(n13441), .ZN(n13450) );
  INV_X1 U15271 ( .A(n13438), .ZN(n13439) );
  OAI21_X1 U15272 ( .B1(n13439), .B2(n14257), .A(n14280), .ZN(n13443) );
  INV_X1 U15273 ( .A(n13443), .ZN(n13440) );
  NAND2_X1 U15274 ( .A1(n13440), .A2(n13446), .ZN(n13445) );
  INV_X1 U15275 ( .A(n13441), .ZN(n13442) );
  OAI21_X1 U15276 ( .B1(n13443), .B2(n13442), .A(n13447), .ZN(n13444) );
  MUX2_X1 U15277 ( .A(n13445), .B(n13444), .S(n13480), .Z(n13449) );
  MUX2_X1 U15278 ( .A(n13447), .B(n13446), .S(n13480), .Z(n13448) );
  OAI211_X1 U15279 ( .C1(n13450), .C2(n13449), .A(n14262), .B(n13448), .ZN(
        n13454) );
  MUX2_X1 U15280 ( .A(n13452), .B(n13451), .S(n13480), .Z(n13453) );
  NAND3_X1 U15281 ( .A1(n13454), .A2(n14245), .A3(n13453), .ZN(n13461) );
  MUX2_X1 U15282 ( .A(n13456), .B(n13455), .S(n13480), .Z(n13460) );
  INV_X1 U15283 ( .A(n13457), .ZN(n13458) );
  NAND3_X1 U15284 ( .A1(n13461), .A2(n13460), .A3(n14230), .ZN(n13469) );
  INV_X1 U15285 ( .A(n13462), .ZN(n13463) );
  MUX2_X1 U15286 ( .A(n13464), .B(n13463), .S(n13491), .Z(n13465) );
  NOR2_X1 U15287 ( .A1(n13465), .A2(n14216), .ZN(n13468) );
  NOR3_X1 U15288 ( .A1(n14865), .A2(n14232), .A3(n13491), .ZN(n13467) );
  NOR3_X1 U15289 ( .A1(n13847), .A2(n14208), .A3(n13480), .ZN(n13466) );
  AOI211_X1 U15290 ( .C1(n13469), .C2(n13468), .A(n13467), .B(n13466), .ZN(
        n13472) );
  NAND3_X1 U15291 ( .A1(n13470), .A2(n14220), .A3(n13480), .ZN(n13471) );
  OAI21_X1 U15292 ( .B1(n8349), .B2(n13472), .A(n13471), .ZN(n13481) );
  OAI21_X1 U15293 ( .B1(n8351), .B2(n8350), .A(n13473), .ZN(n13475) );
  NAND2_X1 U15294 ( .A1(n13475), .A2(n13474), .ZN(n13476) );
  NAND2_X1 U15295 ( .A1(n13477), .A2(n13476), .ZN(n13479) );
  AOI22_X1 U15296 ( .A1(n13545), .A2(n13481), .B1(n13480), .B2(n13482), .ZN(
        n13486) );
  INV_X1 U15297 ( .A(n13482), .ZN(n13483) );
  AND3_X1 U15298 ( .A1(n13487), .A2(n13488), .A3(n13520), .ZN(n13490) );
  INV_X1 U15299 ( .A(n13489), .ZN(n13511) );
  AOI22_X1 U15300 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(n16121), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n15525), .ZN(n13498) );
  XNOR2_X1 U15301 ( .A(n13497), .B(n13498), .ZN(n14909) );
  OR2_X1 U15302 ( .A1(n13494), .A2(n14909), .ZN(n13496) );
  OR2_X1 U15303 ( .A1(n9335), .A2(n14910), .ZN(n13495) );
  OAI21_X1 U15304 ( .B1(n15525), .B2(P2_DATAO_REG_30__SCAN_IN), .A(n13499), 
        .ZN(n13503) );
  AOI22_X1 U15305 ( .A1(P1_DATAO_REG_31__SCAN_IN), .A2(
        P2_DATAO_REG_31__SCAN_IN), .B1(n13501), .B2(n13500), .ZN(n13502) );
  XNOR2_X1 U15306 ( .A(n13503), .B(n13502), .ZN(n14902) );
  NAND2_X1 U15307 ( .A1(n14902), .A2(n13504), .ZN(n13506) );
  INV_X1 U15308 ( .A(SI_31_), .ZN(n14908) );
  OR2_X1 U15309 ( .A1(n9335), .A2(n14908), .ZN(n13505) );
  NOR2_X1 U15310 ( .A1(n14840), .A2(n14151), .ZN(n13546) );
  AOI21_X1 U15311 ( .B1(n13508), .B2(n13521), .A(n13546), .ZN(n13553) );
  INV_X1 U15312 ( .A(n14840), .ZN(n13515) );
  INV_X1 U15313 ( .A(n13509), .ZN(n13514) );
  OAI211_X1 U15314 ( .C1(n14843), .C2(n14151), .A(n13521), .B(n13511), .ZN(
        n13512) );
  XNOR2_X1 U15315 ( .A(n13516), .B(n14132), .ZN(n13519) );
  INV_X1 U15316 ( .A(n13517), .ZN(n13518) );
  INV_X1 U15317 ( .A(n13520), .ZN(n13547) );
  INV_X1 U15318 ( .A(n16499), .ZN(n13523) );
  NAND4_X1 U15319 ( .A1(n13524), .A2(n13523), .A3(n13522), .A4(n16447), .ZN(
        n13531) );
  INV_X1 U15320 ( .A(n13525), .ZN(n13529) );
  NAND4_X1 U15321 ( .A1(n13529), .A2(n13528), .A3(n13527), .A4(n13526), .ZN(
        n13530) );
  NOR2_X1 U15322 ( .A1(n13531), .A2(n13530), .ZN(n13535) );
  AND4_X1 U15323 ( .A1(n13535), .A2(n13534), .A3(n13533), .A4(n13532), .ZN(
        n13536) );
  NAND4_X1 U15324 ( .A1(n13539), .A2(n13538), .A3(n13537), .A4(n13536), .ZN(
        n13540) );
  NOR4_X1 U15325 ( .A1(n14293), .A2(n14326), .A3(n13541), .A4(n13540), .ZN(
        n13542) );
  AND4_X1 U15326 ( .A1(n14319), .A2(n14285), .A3(n14262), .A4(n13542), .ZN(
        n13543) );
  XNOR2_X1 U15327 ( .A(n13548), .B(n14132), .ZN(n13551) );
  NOR3_X1 U15328 ( .A1(n13556), .A2(n13555), .A3(n14921), .ZN(n13559) );
  OAI21_X1 U15329 ( .B1(n13560), .B2(n13557), .A(P3_B_REG_SCAN_IN), .ZN(n13558) );
  OAI22_X1 U15330 ( .A1(n13561), .A2(n13560), .B1(n13559), .B2(n13558), .ZN(
        P3_U3296) );
  INV_X1 U15331 ( .A(n13562), .ZN(n13563) );
  OAI222_X1 U15332 ( .A1(n14918), .A2(n13563), .B1(n14920), .B2(n14477), .C1(
        P3_U3151), .C2(n14139), .ZN(P3_U3268) );
  NAND2_X1 U15333 ( .A1(n15519), .A2(n11544), .ZN(n13565) );
  OR2_X1 U15334 ( .A1(n10704), .A2(n13501), .ZN(n13564) );
  XNOR2_X1 U15335 ( .A(n15743), .B(n13615), .ZN(n13628) );
  INV_X1 U15336 ( .A(n13628), .ZN(n13645) );
  INV_X1 U15337 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n13569) );
  NAND2_X1 U15338 ( .A1(n7420), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n13568) );
  NAND2_X1 U15339 ( .A1(n13566), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n13567) );
  OAI211_X1 U15340 ( .C1(n12862), .C2(n13569), .A(n13568), .B(n13567), .ZN(
        n15788) );
  INV_X1 U15341 ( .A(n16002), .ZN(n13613) );
  XOR2_X1 U15342 ( .A(n15788), .B(n13613), .Z(n13604) );
  OR2_X1 U15343 ( .A1(n15819), .A2(n13570), .ZN(n13571) );
  INV_X1 U15344 ( .A(n15765), .ZN(n15816) );
  NAND2_X1 U15345 ( .A1(n16021), .A2(n15816), .ZN(n15779) );
  OR2_X1 U15346 ( .A1(n16021), .A2(n15816), .ZN(n13572) );
  NAND2_X1 U15347 ( .A1(n15779), .A2(n13572), .ZN(n15828) );
  NAND2_X1 U15348 ( .A1(n15738), .A2(n15859), .ZN(n15764) );
  OR2_X1 U15349 ( .A1(n15738), .A2(n15859), .ZN(n13573) );
  NAND2_X1 U15350 ( .A1(n15764), .A2(n13573), .ZN(n15847) );
  INV_X1 U15351 ( .A(n15759), .ZN(n15939) );
  NAND2_X1 U15352 ( .A1(n16059), .A2(n15939), .ZN(n13574) );
  NAND2_X1 U15353 ( .A1(n15771), .A2(n13574), .ZN(n15925) );
  INV_X1 U15354 ( .A(n15756), .ZN(n15954) );
  INV_X1 U15355 ( .A(n15973), .ZN(n15938) );
  XNOR2_X1 U15356 ( .A(n16074), .B(n15938), .ZN(n15958) );
  NAND2_X1 U15357 ( .A1(n15990), .A2(n15691), .ZN(n13661) );
  AND2_X1 U15358 ( .A1(n16467), .A2(n13661), .ZN(n15992) );
  NAND4_X1 U15359 ( .A1(n13575), .A2(n15992), .A3(n13671), .A4(n16468), .ZN(
        n13577) );
  NOR2_X1 U15360 ( .A1(n13577), .A2(n13576), .ZN(n13581) );
  NAND4_X1 U15361 ( .A1(n13581), .A2(n13580), .A3(n13579), .A4(n13578), .ZN(
        n13584) );
  OR4_X1 U15362 ( .A1(n13585), .A2(n13584), .A3(n13583), .A4(n13582), .ZN(
        n13586) );
  NOR2_X1 U15363 ( .A1(n13587), .A2(n13586), .ZN(n13589) );
  NAND3_X1 U15364 ( .A1(n13590), .A2(n13589), .A3(n13588), .ZN(n13591) );
  NOR2_X1 U15365 ( .A1(n13592), .A2(n13591), .ZN(n13594) );
  NAND4_X1 U15366 ( .A1(n15981), .A2(n13595), .A3(n13594), .A4(n13593), .ZN(
        n13596) );
  NOR4_X1 U15367 ( .A1(n15925), .A2(n15933), .A3(n15958), .A4(n13596), .ZN(
        n13597) );
  XNOR2_X1 U15368 ( .A(n15906), .B(n15676), .ZN(n15774) );
  NAND4_X1 U15369 ( .A1(n15891), .A2(n15847), .A3(n13597), .A4(n15774), .ZN(
        n13598) );
  NOR4_X1 U15370 ( .A1(n15828), .A2(n13598), .A3(n15884), .A4(n15762), .ZN(
        n13603) );
  NAND2_X1 U15371 ( .A1(n13599), .A2(n11544), .ZN(n13602) );
  OR2_X1 U15372 ( .A1(n10704), .A2(n13600), .ZN(n13601) );
  XNOR2_X1 U15373 ( .A(n15786), .B(n15800), .ZN(n15783) );
  MUX2_X1 U15374 ( .A(n13608), .B(n13610), .S(n13616), .Z(n13652) );
  MUX2_X1 U15375 ( .A(n15800), .B(n15786), .S(n13782), .Z(n13630) );
  INV_X1 U15376 ( .A(n13630), .ZN(n13609) );
  MUX2_X1 U15377 ( .A(n15786), .B(n15800), .S(n13779), .Z(n13629) );
  NOR2_X1 U15378 ( .A1(n13609), .A2(n13629), .ZN(n13797) );
  OAI21_X1 U15379 ( .B1(n13615), .B2(n13610), .A(n15788), .ZN(n13611) );
  MUX2_X1 U15380 ( .A(n16002), .B(n13611), .S(n13779), .Z(n13635) );
  INV_X1 U15381 ( .A(n13635), .ZN(n13622) );
  NAND2_X1 U15382 ( .A1(n13613), .A2(n13782), .ZN(n13620) );
  AND2_X1 U15383 ( .A1(n13615), .A2(n13614), .ZN(n13617) );
  MUX2_X1 U15384 ( .A(n15988), .B(n13617), .S(n13616), .Z(n13618) );
  NAND2_X1 U15385 ( .A1(n13618), .A2(n15788), .ZN(n13619) );
  NAND2_X1 U15386 ( .A1(n13620), .A2(n13619), .ZN(n13634) );
  INV_X1 U15387 ( .A(n13634), .ZN(n13621) );
  AND2_X1 U15388 ( .A1(n13622), .A2(n13621), .ZN(n13637) );
  NAND2_X1 U15389 ( .A1(n13624), .A2(n13623), .ZN(n13626) );
  NAND2_X1 U15390 ( .A1(n13626), .A2(n13625), .ZN(n13648) );
  INV_X1 U15391 ( .A(n13648), .ZN(n13627) );
  NAND2_X1 U15392 ( .A1(n13628), .A2(n13627), .ZN(n13639) );
  INV_X1 U15393 ( .A(n13629), .ZN(n13631) );
  NOR2_X1 U15394 ( .A1(n13631), .A2(n13630), .ZN(n13799) );
  NAND2_X1 U15395 ( .A1(n15743), .A2(n15742), .ZN(n13633) );
  MUX2_X1 U15396 ( .A(n13633), .B(n13632), .S(n13782), .Z(n13646) );
  AND2_X1 U15397 ( .A1(n13648), .A2(n13803), .ZN(n13644) );
  NAND2_X1 U15398 ( .A1(n13635), .A2(n13634), .ZN(n13638) );
  NAND2_X1 U15399 ( .A1(n13636), .A2(n13638), .ZN(n13798) );
  INV_X1 U15400 ( .A(n13798), .ZN(n13643) );
  INV_X1 U15401 ( .A(n13636), .ZN(n13641) );
  INV_X1 U15402 ( .A(n13637), .ZN(n13640) );
  OAI22_X1 U15403 ( .A1(n13641), .A2(n13640), .B1(n13639), .B2(n13638), .ZN(
        n13642) );
  AOI21_X1 U15404 ( .B1(n13799), .B2(n13643), .A(n13642), .ZN(n13651) );
  NAND2_X1 U15405 ( .A1(n13645), .A2(n13644), .ZN(n13649) );
  INV_X1 U15406 ( .A(n13646), .ZN(n13647) );
  MUX2_X1 U15407 ( .A(n13649), .B(n13648), .S(n13647), .Z(n13650) );
  MUX2_X1 U15408 ( .A(n15815), .B(n15808), .S(n13735), .Z(n13795) );
  AOI21_X1 U15409 ( .B1(n13655), .B2(n13782), .A(n13653), .ZN(n13658) );
  AOI21_X1 U15410 ( .B1(n15690), .B2(n13612), .A(n16527), .ZN(n13657) );
  OAI211_X1 U15411 ( .C1(n13655), .C2(n16527), .A(n13654), .B(n13779), .ZN(
        n13656) );
  OAI21_X1 U15412 ( .B1(n13658), .B2(n13657), .A(n13656), .ZN(n13659) );
  INV_X1 U15413 ( .A(n13659), .ZN(n13676) );
  NAND2_X1 U15414 ( .A1(n16467), .A2(n13660), .ZN(n13662) );
  NAND3_X1 U15415 ( .A1(n13664), .A2(n13668), .A3(n16468), .ZN(n13673) );
  OAI21_X1 U15416 ( .B1(n13668), .B2(n13612), .A(n13665), .ZN(n13666) );
  INV_X1 U15417 ( .A(n13666), .ZN(n13672) );
  NAND4_X1 U15418 ( .A1(n13673), .A2(n13672), .A3(n13671), .A4(n13670), .ZN(
        n13674) );
  AOI21_X1 U15419 ( .B1(n13678), .B2(n13612), .A(n13677), .ZN(n13679) );
  AOI21_X1 U15420 ( .B1(n15689), .B2(n13779), .A(n16554), .ZN(n13680) );
  MUX2_X1 U15421 ( .A(n13684), .B(n16572), .S(n13652), .Z(n13687) );
  MUX2_X1 U15422 ( .A(n13685), .B(n15688), .S(n13782), .Z(n13686) );
  MUX2_X1 U15423 ( .A(n13689), .B(n15687), .S(n13652), .Z(n13692) );
  NAND2_X1 U15424 ( .A1(n13688), .A2(n13692), .ZN(n13691) );
  MUX2_X1 U15425 ( .A(n15687), .B(n13689), .S(n13779), .Z(n13690) );
  NAND2_X1 U15426 ( .A1(n13691), .A2(n13690), .ZN(n13698) );
  INV_X1 U15427 ( .A(n13692), .ZN(n13693) );
  AND2_X1 U15428 ( .A1(n13694), .A2(n13693), .ZN(n13695) );
  NAND2_X1 U15429 ( .A1(n13696), .A2(n13695), .ZN(n13697) );
  MUX2_X1 U15430 ( .A(n15686), .B(n16607), .S(n13782), .Z(n13701) );
  MUX2_X1 U15431 ( .A(n16607), .B(n15686), .S(n13782), .Z(n13699) );
  INV_X1 U15432 ( .A(n13701), .ZN(n13702) );
  MUX2_X1 U15433 ( .A(n15685), .B(n16627), .S(n13735), .Z(n13706) );
  MUX2_X1 U15434 ( .A(n15685), .B(n16627), .S(n13779), .Z(n13703) );
  NAND2_X1 U15435 ( .A1(n13704), .A2(n13703), .ZN(n13710) );
  INV_X1 U15436 ( .A(n13705), .ZN(n13708) );
  INV_X1 U15437 ( .A(n13706), .ZN(n13707) );
  NAND2_X1 U15438 ( .A1(n13708), .A2(n13707), .ZN(n13709) );
  MUX2_X1 U15439 ( .A(n15684), .B(n13711), .S(n13782), .Z(n13713) );
  MUX2_X1 U15440 ( .A(n15684), .B(n13711), .S(n13735), .Z(n13712) );
  INV_X1 U15441 ( .A(n13713), .ZN(n13714) );
  MUX2_X1 U15442 ( .A(n15683), .B(n13715), .S(n13735), .Z(n13717) );
  MUX2_X1 U15443 ( .A(n15683), .B(n13715), .S(n13782), .Z(n13716) );
  INV_X1 U15444 ( .A(n13717), .ZN(n13718) );
  MUX2_X1 U15445 ( .A(n15682), .B(n13719), .S(n13779), .Z(n13723) );
  MUX2_X1 U15446 ( .A(n15682), .B(n13719), .S(n13735), .Z(n13720) );
  NAND2_X1 U15447 ( .A1(n13721), .A2(n13720), .ZN(n13727) );
  INV_X1 U15448 ( .A(n13722), .ZN(n13725) );
  INV_X1 U15449 ( .A(n13723), .ZN(n13724) );
  NAND2_X1 U15450 ( .A1(n13725), .A2(n13724), .ZN(n13726) );
  MUX2_X1 U15451 ( .A(n15681), .B(n13728), .S(n13735), .Z(n13730) );
  MUX2_X1 U15452 ( .A(n15681), .B(n13728), .S(n13782), .Z(n13729) );
  INV_X1 U15453 ( .A(n13730), .ZN(n13731) );
  MUX2_X1 U15454 ( .A(n15680), .B(n16722), .S(n13652), .Z(n13734) );
  MUX2_X1 U15455 ( .A(n15680), .B(n16722), .S(n13735), .Z(n13732) );
  MUX2_X1 U15456 ( .A(n15679), .B(n13736), .S(n13735), .Z(n13738) );
  MUX2_X1 U15457 ( .A(n15679), .B(n13736), .S(n13779), .Z(n13737) );
  INV_X1 U15458 ( .A(n13738), .ZN(n13739) );
  MUX2_X1 U15459 ( .A(n15678), .B(n16090), .S(n13782), .Z(n13743) );
  MUX2_X1 U15460 ( .A(n15678), .B(n16090), .S(n13735), .Z(n13740) );
  NAND2_X1 U15461 ( .A1(n13741), .A2(n13740), .ZN(n13747) );
  INV_X1 U15462 ( .A(n13742), .ZN(n13745) );
  INV_X1 U15463 ( .A(n13743), .ZN(n13744) );
  NAND2_X1 U15464 ( .A1(n13745), .A2(n13744), .ZN(n13746) );
  MUX2_X1 U15465 ( .A(n15972), .B(n16085), .S(n13735), .Z(n13749) );
  MUX2_X1 U15466 ( .A(n15972), .B(n16085), .S(n13782), .Z(n13748) );
  MUX2_X1 U15467 ( .A(n15755), .B(n16078), .S(n13779), .Z(n13751) );
  MUX2_X1 U15468 ( .A(n15755), .B(n16078), .S(n13735), .Z(n13750) );
  MUX2_X1 U15469 ( .A(n15973), .B(n16074), .S(n13735), .Z(n13753) );
  MUX2_X1 U15470 ( .A(n15973), .B(n16074), .S(n13782), .Z(n13752) );
  INV_X1 U15471 ( .A(n13753), .ZN(n13754) );
  MUX2_X1 U15472 ( .A(n15756), .B(n16068), .S(n13652), .Z(n13757) );
  MUX2_X1 U15473 ( .A(n15756), .B(n16068), .S(n13735), .Z(n13755) );
  MUX2_X1 U15474 ( .A(n15759), .B(n16059), .S(n13735), .Z(n13759) );
  MUX2_X1 U15475 ( .A(n15759), .B(n16059), .S(n13779), .Z(n13758) );
  INV_X1 U15476 ( .A(n13759), .ZN(n13760) );
  MUX2_X1 U15477 ( .A(n15676), .B(n15906), .S(n13782), .Z(n13764) );
  MUX2_X1 U15478 ( .A(n15676), .B(n15906), .S(n13735), .Z(n13761) );
  INV_X1 U15479 ( .A(n13763), .ZN(n13766) );
  INV_X1 U15480 ( .A(n13764), .ZN(n13765) );
  MUX2_X1 U15481 ( .A(n16046), .B(n15761), .S(n13782), .Z(n13768) );
  MUX2_X1 U15482 ( .A(n15761), .B(n16046), .S(n13779), .Z(n13767) );
  MUX2_X1 U15483 ( .A(n15860), .B(n16040), .S(n13782), .Z(n13770) );
  MUX2_X1 U15484 ( .A(n15675), .B(n15869), .S(n13735), .Z(n13774) );
  NAND2_X1 U15485 ( .A1(n13773), .A2(n13774), .ZN(n13772) );
  MUX2_X1 U15486 ( .A(n15675), .B(n15869), .S(n13782), .Z(n13771) );
  NAND2_X1 U15487 ( .A1(n13772), .A2(n13771), .ZN(n13778) );
  INV_X1 U15488 ( .A(n13773), .ZN(n13776) );
  INV_X1 U15489 ( .A(n13774), .ZN(n13775) );
  NAND2_X1 U15490 ( .A1(n13776), .A2(n13775), .ZN(n13777) );
  MUX2_X1 U15491 ( .A(n15859), .B(n15738), .S(n13779), .Z(n13781) );
  MUX2_X1 U15492 ( .A(n15859), .B(n15738), .S(n13735), .Z(n13780) );
  MUX2_X1 U15493 ( .A(n15765), .B(n16021), .S(n13735), .Z(n13785) );
  MUX2_X1 U15494 ( .A(n15765), .B(n16021), .S(n13782), .Z(n13783) );
  MUX2_X1 U15495 ( .A(n15838), .B(n15819), .S(n13652), .Z(n13789) );
  MUX2_X1 U15496 ( .A(n15838), .B(n15819), .S(n13735), .Z(n13786) );
  NAND2_X1 U15497 ( .A1(n13787), .A2(n13786), .ZN(n13793) );
  INV_X1 U15498 ( .A(n13788), .ZN(n13791) );
  INV_X1 U15499 ( .A(n13789), .ZN(n13790) );
  NAND2_X1 U15500 ( .A1(n13791), .A2(n13790), .ZN(n13792) );
  MUX2_X1 U15501 ( .A(n15791), .B(n16011), .S(n13652), .Z(n13794) );
  NOR2_X1 U15502 ( .A1(n13800), .A2(n13799), .ZN(n13801) );
  NOR3_X1 U15503 ( .A1(n13804), .A2(n7417), .A3(n15951), .ZN(n13806) );
  OAI21_X1 U15504 ( .B1(n16137), .B2(n13607), .A(P1_B_REG_SCAN_IN), .ZN(n13805) );
  OAI22_X1 U15505 ( .A1(n13807), .A2(n16137), .B1(n13806), .B2(n13805), .ZN(
        P1_U3242) );
  NOR2_X1 U15506 ( .A1(n13808), .A2(n16508), .ZN(n14152) );
  AOI21_X1 U15507 ( .B1(n16517), .B2(P3_REG2_REG_29__SCAN_IN), .A(n14152), 
        .ZN(n13809) );
  OAI21_X1 U15508 ( .B1(n13810), .B2(n14384), .A(n13809), .ZN(n13811) );
  AOI21_X1 U15509 ( .B1(n13812), .B2(n14372), .A(n13811), .ZN(n13813) );
  OAI21_X1 U15510 ( .B1(n13814), .B2(n16517), .A(n13813), .ZN(P3_U3204) );
  XNOR2_X1 U15511 ( .A(n14163), .B(n13815), .ZN(n13823) );
  INV_X1 U15512 ( .A(n13823), .ZN(n13816) );
  NAND2_X1 U15513 ( .A1(n13816), .A2(n16451), .ZN(n13829) );
  INV_X1 U15514 ( .A(n13817), .ZN(n13818) );
  NAND4_X1 U15515 ( .A1(n13828), .A2(n16451), .A3(n13818), .A4(n13823), .ZN(
        n13827) );
  NAND2_X1 U15516 ( .A1(n13970), .A2(n14165), .ZN(n13820) );
  AOI22_X1 U15517 ( .A1(n13821), .A2(n13982), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13819) );
  OAI211_X1 U15518 ( .C1(n14158), .C2(n13978), .A(n13820), .B(n13819), .ZN(
        n13825) );
  NOR4_X1 U15519 ( .A1(n13823), .A2(n13822), .A3(n13821), .A4(n13954), .ZN(
        n13824) );
  AOI211_X1 U15520 ( .C1(n16449), .C2(n14392), .A(n13825), .B(n13824), .ZN(
        n13826) );
  OAI211_X1 U15521 ( .C1(n13829), .C2(n13828), .A(n13827), .B(n13826), .ZN(
        P3_U3160) );
  INV_X1 U15522 ( .A(n13830), .ZN(n13833) );
  OAI222_X1 U15523 ( .A1(n14918), .A2(n13833), .B1(n14920), .B2(n13832), .C1(
        P3_U3151), .C2(n13831), .ZN(P3_U3271) );
  OAI21_X1 U15524 ( .B1(n13835), .B2(n13834), .A(n13974), .ZN(n13836) );
  NAND2_X1 U15525 ( .A1(n13836), .A2(n16451), .ZN(n13841) );
  INV_X1 U15526 ( .A(n13837), .ZN(n14368) );
  INV_X1 U15527 ( .A(n13978), .ZN(n16448) );
  INV_X1 U15528 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n14643) );
  NOR2_X1 U15529 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n14643), .ZN(n14019) );
  AOI21_X1 U15530 ( .B1(n16448), .B2(n14363), .A(n14019), .ZN(n13838) );
  OAI21_X1 U15531 ( .B1(n8160), .B2(n13947), .A(n13838), .ZN(n13839) );
  AOI21_X1 U15532 ( .B1(n13970), .B2(n14368), .A(n13839), .ZN(n13840) );
  OAI211_X1 U15533 ( .C1(n13985), .C2(n14895), .A(n13841), .B(n13840), .ZN(
        P3_U3155) );
  INV_X1 U15534 ( .A(n13842), .ZN(n13916) );
  AOI21_X1 U15535 ( .B1(n13843), .B2(n14232), .A(n13916), .ZN(n13849) );
  NAND2_X1 U15536 ( .A1(n13970), .A2(n14223), .ZN(n13845) );
  AOI22_X1 U15537 ( .A1(n13982), .A2(n14246), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13844) );
  OAI211_X1 U15538 ( .C1(n14220), .C2(n13978), .A(n13845), .B(n13844), .ZN(
        n13846) );
  AOI21_X1 U15539 ( .B1(n13847), .B2(n16449), .A(n13846), .ZN(n13848) );
  OAI21_X1 U15540 ( .B1(n13849), .B2(n13954), .A(n13848), .ZN(P3_U3156) );
  NAND2_X1 U15541 ( .A1(n13975), .A2(n13850), .ZN(n13953) );
  NAND2_X1 U15542 ( .A1(n13953), .A2(n13851), .ZN(n13957) );
  NAND2_X1 U15543 ( .A1(n13957), .A2(n13852), .ZN(n13858) );
  NAND2_X1 U15544 ( .A1(n13975), .A2(n13853), .ZN(n13855) );
  NAND2_X1 U15545 ( .A1(n13855), .A2(n13854), .ZN(n13856) );
  OAI211_X1 U15546 ( .C1(n13858), .C2(n13857), .A(n13856), .B(n16451), .ZN(
        n13863) );
  NAND2_X1 U15547 ( .A1(n13982), .A2(n13859), .ZN(n13860) );
  NAND2_X1 U15548 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n14135)
         );
  OAI211_X1 U15549 ( .C1(n14278), .C2(n13978), .A(n13860), .B(n14135), .ZN(
        n13861) );
  AOI21_X1 U15550 ( .B1(n13970), .B2(n14287), .A(n13861), .ZN(n13862) );
  OAI211_X1 U15551 ( .C1(n14881), .C2(n13985), .A(n13863), .B(n13862), .ZN(
        P3_U3159) );
  INV_X1 U15552 ( .A(n13864), .ZN(n13865) );
  NOR2_X1 U15553 ( .A1(n13866), .A2(n13865), .ZN(n13867) );
  XNOR2_X1 U15554 ( .A(n13868), .B(n13867), .ZN(n13873) );
  OAI22_X1 U15555 ( .A1(n13978), .A2(n14219), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n14641), .ZN(n13869) );
  AOI21_X1 U15556 ( .B1(n13982), .B2(n8153), .A(n13869), .ZN(n13870) );
  OAI21_X1 U15557 ( .B1(n13979), .B2(n14250), .A(n13870), .ZN(n13871) );
  AOI21_X1 U15558 ( .B1(n14253), .B2(n16449), .A(n13871), .ZN(n13872) );
  OAI21_X1 U15559 ( .B1(n13873), .B2(n13954), .A(n13872), .ZN(P3_U3163) );
  XNOR2_X1 U15560 ( .A(n13874), .B(n13934), .ZN(n13875) );
  XNOR2_X1 U15561 ( .A(n13876), .B(n13875), .ZN(n13883) );
  INV_X1 U15562 ( .A(n14383), .ZN(n13881) );
  AOI22_X1 U15563 ( .A1(n13982), .A2(n14380), .B1(n16449), .B2(n13877), .ZN(
        n13879) );
  OAI211_X1 U15564 ( .C1(n8160), .C2(n13978), .A(n13879), .B(n13878), .ZN(
        n13880) );
  AOI21_X1 U15565 ( .B1(n13970), .B2(n13881), .A(n13880), .ZN(n13882) );
  OAI21_X1 U15566 ( .B1(n13883), .B2(n13954), .A(n13882), .ZN(P3_U3164) );
  INV_X1 U15567 ( .A(n13884), .ZN(n13917) );
  INV_X1 U15568 ( .A(n13885), .ZN(n13887) );
  NOR3_X1 U15569 ( .A1(n13917), .A2(n13887), .A3(n13886), .ZN(n13890) );
  INV_X1 U15570 ( .A(n13888), .ZN(n13889) );
  OAI21_X1 U15571 ( .B1(n13890), .B2(n13889), .A(n16451), .ZN(n13894) );
  NOR2_X1 U15572 ( .A1(n13947), .A2(n14220), .ZN(n13892) );
  OAI22_X1 U15573 ( .A1(n14198), .A2(n13978), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n14712), .ZN(n13891) );
  AOI211_X1 U15574 ( .C1(n13970), .C2(n14200), .A(n13892), .B(n13891), .ZN(
        n13893) );
  OAI211_X1 U15575 ( .C1(n8351), .C2(n13985), .A(n13894), .B(n13893), .ZN(
        P3_U3165) );
  NAND2_X1 U15576 ( .A1(n13975), .A2(n13895), .ZN(n13902) );
  XNOR2_X1 U15577 ( .A(n13902), .B(n13901), .ZN(n13900) );
  NAND2_X1 U15578 ( .A1(P3_REG3_REG_16__SCAN_IN), .A2(P3_U3151), .ZN(n14073)
         );
  OAI21_X1 U15579 ( .B1(n13978), .B2(n13905), .A(n14073), .ZN(n13896) );
  AOI21_X1 U15580 ( .B1(n13982), .B2(n14363), .A(n13896), .ZN(n13897) );
  OAI21_X1 U15581 ( .B1(n13979), .B2(n14335), .A(n13897), .ZN(n13898) );
  AOI21_X1 U15582 ( .B1(n16449), .B2(n14441), .A(n13898), .ZN(n13899) );
  OAI21_X1 U15583 ( .B1(n13900), .B2(n13954), .A(n13899), .ZN(P3_U3166) );
  NAND2_X1 U15584 ( .A1(n13902), .A2(n13901), .ZN(n13904) );
  NAND2_X1 U15585 ( .A1(n13904), .A2(n13903), .ZN(n13908) );
  XNOR2_X1 U15586 ( .A(n13906), .B(n13905), .ZN(n13907) );
  XNOR2_X1 U15587 ( .A(n13908), .B(n13907), .ZN(n13909) );
  NAND2_X1 U15588 ( .A1(n13909), .A2(n16451), .ZN(n13913) );
  NAND2_X1 U15589 ( .A1(P3_U3151), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n14085)
         );
  OAI21_X1 U15590 ( .B1(n13978), .B2(n14313), .A(n14085), .ZN(n13911) );
  NOR2_X1 U15591 ( .A1(n13979), .A2(n14321), .ZN(n13910) );
  AOI211_X1 U15592 ( .C1(n13982), .C2(n14348), .A(n13911), .B(n13910), .ZN(
        n13912) );
  OAI211_X1 U15593 ( .C1(n13985), .C2(n14886), .A(n13913), .B(n13912), .ZN(
        P3_U3168) );
  NOR3_X1 U15594 ( .A1(n13916), .A2(n8735), .A3(n13915), .ZN(n13918) );
  OAI21_X1 U15595 ( .B1(n13918), .B2(n13917), .A(n16451), .ZN(n13922) );
  NOR2_X1 U15596 ( .A1(n13947), .A2(n14208), .ZN(n13920) );
  OAI22_X1 U15597 ( .A1(n14209), .A2(n13978), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n14634), .ZN(n13919) );
  AOI211_X1 U15598 ( .C1(n13970), .C2(n14211), .A(n13920), .B(n13919), .ZN(
        n13921) );
  OAI211_X1 U15599 ( .C1(n14861), .C2(n13985), .A(n13922), .B(n13921), .ZN(
        P3_U3169) );
  OAI211_X1 U15600 ( .C1(n13925), .C2(n13924), .A(n13923), .B(n16451), .ZN(
        n13931) );
  NOR2_X1 U15601 ( .A1(n13947), .A2(n14264), .ZN(n13928) );
  OAI22_X1 U15602 ( .A1(n13978), .A2(n14265), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n13926), .ZN(n13927) );
  AOI211_X1 U15603 ( .C1(n13970), .C2(n13929), .A(n13928), .B(n13927), .ZN(
        n13930) );
  OAI211_X1 U15604 ( .C1(n14877), .C2(n13985), .A(n13931), .B(n13930), .ZN(
        P3_U3173) );
  XNOR2_X1 U15605 ( .A(n13933), .B(n13932), .ZN(n13941) );
  INV_X1 U15606 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n14632) );
  NOR2_X1 U15607 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n14632), .ZN(n14002) );
  NOR2_X1 U15608 ( .A1(n13947), .A2(n13934), .ZN(n13935) );
  AOI211_X1 U15609 ( .C1(n16448), .C2(n14347), .A(n14002), .B(n13935), .ZN(
        n13936) );
  OAI21_X1 U15610 ( .B1(n13979), .B2(n13937), .A(n13936), .ZN(n13938) );
  AOI21_X1 U15611 ( .B1(n13939), .B2(n16449), .A(n13938), .ZN(n13940) );
  OAI21_X1 U15612 ( .B1(n13941), .B2(n13954), .A(n13940), .ZN(P3_U3174) );
  INV_X1 U15613 ( .A(n13943), .ZN(n13945) );
  OAI21_X1 U15614 ( .B1(n13945), .B2(n14219), .A(n13944), .ZN(n13946) );
  NAND2_X1 U15615 ( .A1(n13946), .A2(n16451), .ZN(n13951) );
  NOR2_X1 U15616 ( .A1(n13947), .A2(n14265), .ZN(n13949) );
  INV_X1 U15617 ( .A(P3_REG3_REG_22__SCAN_IN), .ZN(n14720) );
  OAI22_X1 U15618 ( .A1(n13978), .A2(n14208), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n14720), .ZN(n13948) );
  AOI211_X1 U15619 ( .C1(n13970), .C2(n14237), .A(n13949), .B(n13948), .ZN(
        n13950) );
  OAI211_X1 U15620 ( .C1(n14869), .C2(n13985), .A(n13951), .B(n13950), .ZN(
        P3_U3175) );
  NAND2_X1 U15621 ( .A1(n13953), .A2(n13952), .ZN(n13956) );
  AOI21_X1 U15622 ( .B1(n13956), .B2(n13955), .A(n13954), .ZN(n13958) );
  NAND2_X1 U15623 ( .A1(n13958), .A2(n13957), .ZN(n13962) );
  NAND2_X1 U15624 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n14123)
         );
  OAI21_X1 U15625 ( .B1(n13978), .B2(n14264), .A(n14123), .ZN(n13960) );
  NOR2_X1 U15626 ( .A1(n13979), .A2(n14301), .ZN(n13959) );
  AOI211_X1 U15627 ( .C1(n13982), .C2(n14328), .A(n13960), .B(n13959), .ZN(
        n13961) );
  OAI211_X1 U15628 ( .C1(n14433), .C2(n13985), .A(n13962), .B(n13961), .ZN(
        P3_U3178) );
  OAI21_X1 U15629 ( .B1(n13965), .B2(n13964), .A(n13963), .ZN(n13966) );
  NAND2_X1 U15630 ( .A1(n13966), .A2(n16451), .ZN(n13972) );
  AOI22_X1 U15631 ( .A1(n8350), .A2(n13982), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13968) );
  OAI21_X1 U15632 ( .B1(n14184), .B2(n13978), .A(n13968), .ZN(n13969) );
  AOI21_X1 U15633 ( .B1(n13970), .B2(n14187), .A(n13969), .ZN(n13971) );
  OAI211_X1 U15634 ( .C1(n14854), .C2(n13985), .A(n13972), .B(n13971), .ZN(
        P3_U3180) );
  AND2_X1 U15635 ( .A1(n13974), .A2(n13973), .ZN(n13977) );
  OAI211_X1 U15636 ( .C1(n13977), .C2(n13976), .A(n16451), .B(n13975), .ZN(
        n13984) );
  INV_X1 U15637 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n14470) );
  OR2_X1 U15638 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n14470), .ZN(n14042) );
  OAI21_X1 U15639 ( .B1(n13978), .B2(n14311), .A(n14042), .ZN(n13981) );
  NOR2_X1 U15640 ( .A1(n13979), .A2(n14351), .ZN(n13980) );
  AOI211_X1 U15641 ( .C1(n13982), .C2(n14347), .A(n13981), .B(n13980), .ZN(
        n13983) );
  OAI211_X1 U15642 ( .C1(n13985), .C2(n14445), .A(n13984), .B(n13983), .ZN(
        P3_U3181) );
  MUX2_X1 U15643 ( .A(P3_DATAO_REG_24__SCAN_IN), .B(n14195), .S(P3_U3897), .Z(
        P3_U3515) );
  MUX2_X1 U15644 ( .A(P3_DATAO_REG_22__SCAN_IN), .B(n14246), .S(P3_U3897), .Z(
        P3_U3513) );
  MUX2_X1 U15645 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n14112), .Z(n13986) );
  NAND2_X1 U15646 ( .A1(n13986), .A2(n13997), .ZN(n13987) );
  MUX2_X1 U15647 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n14139), .Z(n14023) );
  XNOR2_X1 U15648 ( .A(n14023), .B(n14024), .ZN(n13989) );
  NAND2_X1 U15649 ( .A1(n13990), .A2(n13989), .ZN(n14027) );
  OAI21_X1 U15650 ( .B1(n13990), .B2(n13989), .A(n14027), .ZN(n13991) );
  NAND2_X1 U15651 ( .A1(n13991), .A2(n14125), .ZN(n14007) );
  AOI21_X1 U15652 ( .B1(n13994), .B2(n9155), .A(n14009), .ZN(n13995) );
  NOR2_X1 U15653 ( .A1(n16429), .A2(n13995), .ZN(n14005) );
  INV_X1 U15654 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n16365) );
  NOR2_X1 U15655 ( .A1(n16438), .A2(n16365), .ZN(n14004) );
  AOI21_X1 U15656 ( .B1(n13997), .B2(P3_REG2_REG_12__SCAN_IN), .A(n13996), 
        .ZN(n13998) );
  NOR2_X1 U15657 ( .A1(n13998), .A2(n14024), .ZN(n14014) );
  NAND2_X1 U15658 ( .A1(n13998), .A2(n14024), .ZN(n13999) );
  AOI21_X1 U15659 ( .B1(n14000), .B2(n9156), .A(n14015), .ZN(n14001) );
  NOR2_X1 U15660 ( .A1(n16423), .A2(n14001), .ZN(n14003) );
  NOR4_X1 U15661 ( .A1(n14005), .A2(n14004), .A3(n14003), .A4(n14002), .ZN(
        n14006) );
  OAI211_X1 U15662 ( .C1(n16427), .C2(n14008), .A(n14007), .B(n14006), .ZN(
        P3_U3195) );
  AOI22_X1 U15663 ( .A1(P3_REG1_REG_14__SCAN_IN), .A2(n14033), .B1(n14046), 
        .B2(n14453), .ZN(n14011) );
  AOI21_X1 U15664 ( .B1(n14012), .B2(n14011), .A(n14036), .ZN(n14035) );
  INV_X1 U15665 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n14022) );
  INV_X1 U15666 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n14013) );
  AOI22_X1 U15667 ( .A1(P3_REG2_REG_14__SCAN_IN), .A2(n14033), .B1(n14046), 
        .B2(n14013), .ZN(n14017) );
  AOI21_X1 U15668 ( .B1(n14017), .B2(n14016), .A(n14039), .ZN(n14018) );
  OR2_X1 U15669 ( .A1(n16423), .A2(n14018), .ZN(n14021) );
  INV_X1 U15670 ( .A(n14019), .ZN(n14020) );
  OAI211_X1 U15671 ( .C1(n16438), .C2(n14022), .A(n14021), .B(n14020), .ZN(
        n14032) );
  MUX2_X1 U15672 ( .A(P3_REG2_REG_14__SCAN_IN), .B(P3_REG1_REG_14__SCAN_IN), 
        .S(n14139), .Z(n14047) );
  XNOR2_X1 U15673 ( .A(n14047), .B(n14046), .ZN(n14030) );
  INV_X1 U15674 ( .A(n14023), .ZN(n14025) );
  NAND2_X1 U15675 ( .A1(n14025), .A2(n14024), .ZN(n14026) );
  INV_X1 U15676 ( .A(n14049), .ZN(n14028) );
  AOI211_X1 U15677 ( .C1(n14030), .C2(n14029), .A(n16418), .B(n14028), .ZN(
        n14031) );
  AOI211_X1 U15678 ( .C1(n14146), .C2(n14033), .A(n14032), .B(n14031), .ZN(
        n14034) );
  OAI21_X1 U15679 ( .B1(n14035), .B2(n16429), .A(n14034), .ZN(P3_U3196) );
  AOI21_X1 U15680 ( .B1(n14038), .B2(n14449), .A(n14057), .ZN(n14055) );
  AOI21_X1 U15681 ( .B1(n8857), .B2(n8435), .A(n7440), .ZN(n14041) );
  NOR2_X1 U15682 ( .A1(n16423), .A2(n14041), .ZN(n14045) );
  INV_X1 U15683 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n14043) );
  OAI21_X1 U15684 ( .B1(n16438), .B2(n14043), .A(n14042), .ZN(n14044) );
  AOI211_X1 U15685 ( .C1(n14146), .C2(n14063), .A(n14045), .B(n14044), .ZN(
        n14054) );
  NAND2_X1 U15686 ( .A1(n14047), .A2(n14046), .ZN(n14048) );
  MUX2_X1 U15687 ( .A(n8435), .B(n14449), .S(n14139), .Z(n14050) );
  NAND2_X1 U15688 ( .A1(n14051), .A2(n14050), .ZN(n14066) );
  OAI21_X1 U15689 ( .B1(n14051), .B2(n14050), .A(n14066), .ZN(n14052) );
  NAND2_X1 U15690 ( .A1(n14052), .A2(n14125), .ZN(n14053) );
  OAI211_X1 U15691 ( .C1(n14055), .C2(n16429), .A(n14054), .B(n14053), .ZN(
        P3_U3197) );
  INV_X1 U15692 ( .A(n14056), .ZN(n14058) );
  NAND2_X1 U15693 ( .A1(P3_REG1_REG_16__SCAN_IN), .A2(n14083), .ZN(n14059) );
  OAI21_X1 U15694 ( .B1(P3_REG1_REG_16__SCAN_IN), .B2(n14083), .A(n14059), 
        .ZN(n14060) );
  AOI21_X1 U15695 ( .B1(n14061), .B2(n14060), .A(n14080), .ZN(n14079) );
  INV_X1 U15696 ( .A(n14062), .ZN(n14064) );
  NAND2_X1 U15697 ( .A1(n14064), .A2(n14063), .ZN(n14065) );
  NAND2_X1 U15698 ( .A1(n14066), .A2(n14065), .ZN(n14068) );
  MUX2_X1 U15699 ( .A(P3_REG2_REG_16__SCAN_IN), .B(P3_REG1_REG_16__SCAN_IN), 
        .S(n14139), .Z(n14088) );
  INV_X1 U15700 ( .A(n14083), .ZN(n14089) );
  XNOR2_X1 U15701 ( .A(n14088), .B(n14089), .ZN(n14067) );
  NAND2_X1 U15702 ( .A1(n14068), .A2(n14067), .ZN(n14092) );
  OAI21_X1 U15703 ( .B1(n14068), .B2(n14067), .A(n14092), .ZN(n14077) );
  NOR2_X1 U15704 ( .A1(n16427), .A2(n14083), .ZN(n14076) );
  NAND2_X1 U15705 ( .A1(P3_REG2_REG_16__SCAN_IN), .A2(n14083), .ZN(n14069) );
  OAI21_X1 U15706 ( .B1(P3_REG2_REG_16__SCAN_IN), .B2(n14083), .A(n14069), 
        .ZN(n14071) );
  NOR2_X1 U15707 ( .A1(n14070), .A2(n14071), .ZN(n14082) );
  AOI21_X1 U15708 ( .B1(n14071), .B2(n14070), .A(n14082), .ZN(n14074) );
  NAND2_X1 U15709 ( .A1(n16150), .A2(P3_ADDR_REG_16__SCAN_IN), .ZN(n14072) );
  OAI211_X1 U15710 ( .C1(n16423), .C2(n14074), .A(n14073), .B(n14072), .ZN(
        n14075) );
  AOI211_X1 U15711 ( .C1(n14077), .C2(n14125), .A(n14076), .B(n14075), .ZN(
        n14078) );
  OAI21_X1 U15712 ( .B1(n14079), .B2(n16429), .A(n14078), .ZN(P3_U3198) );
  AOI21_X1 U15713 ( .B1(n14439), .B2(n14081), .A(n14105), .ZN(n14100) );
  INV_X1 U15714 ( .A(P3_ADDR_REG_17__SCAN_IN), .ZN(n14087) );
  NOR2_X1 U15715 ( .A1(n7502), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n14084) );
  OAI21_X1 U15716 ( .B1(n14119), .B2(n14084), .A(n14120), .ZN(n14086) );
  OAI211_X1 U15717 ( .C1(n16438), .C2(n14087), .A(n14086), .B(n14085), .ZN(
        n14097) );
  MUX2_X1 U15718 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n14139), .Z(n14109) );
  XNOR2_X1 U15719 ( .A(n14109), .B(n14108), .ZN(n14095) );
  INV_X1 U15720 ( .A(n14088), .ZN(n14090) );
  NAND2_X1 U15721 ( .A1(n14090), .A2(n14089), .ZN(n14091) );
  NAND2_X1 U15722 ( .A1(n14092), .A2(n14091), .ZN(n14094) );
  INV_X1 U15723 ( .A(n14111), .ZN(n14093) );
  AOI211_X1 U15724 ( .C1(n14095), .C2(n14094), .A(n16418), .B(n14093), .ZN(
        n14096) );
  AOI211_X1 U15725 ( .C1(n14146), .C2(n14098), .A(n14097), .B(n14096), .ZN(
        n14099) );
  OAI21_X1 U15726 ( .B1(n14100), .B2(n16429), .A(n14099), .ZN(P3_U3199) );
  INV_X1 U15727 ( .A(n14101), .ZN(n14104) );
  OR2_X1 U15728 ( .A1(n14137), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n14102) );
  NAND2_X1 U15729 ( .A1(n14137), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n14128) );
  AND2_X1 U15730 ( .A1(n14102), .A2(n14128), .ZN(n14103) );
  INV_X1 U15731 ( .A(n14129), .ZN(n14107) );
  NOR3_X1 U15732 ( .A1(n14105), .A2(n14104), .A3(n14103), .ZN(n14106) );
  NOR2_X1 U15733 ( .A1(n14107), .A2(n14106), .ZN(n14127) );
  NAND2_X1 U15734 ( .A1(n14109), .A2(n14108), .ZN(n14110) );
  INV_X1 U15735 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n14302) );
  MUX2_X1 U15736 ( .A(n14302), .B(n14113), .S(n14112), .Z(n14114) );
  OAI21_X1 U15737 ( .B1(n14115), .B2(n14114), .A(n14136), .ZN(n14126) );
  NOR2_X1 U15738 ( .A1(n16427), .A2(n14137), .ZN(n14124) );
  INV_X1 U15739 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n16404) );
  OR2_X1 U15740 ( .A1(n14137), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n14116) );
  NAND2_X1 U15741 ( .A1(n14137), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n14130) );
  AND2_X1 U15742 ( .A1(n14116), .A2(n14130), .ZN(n14117) );
  INV_X1 U15743 ( .A(n14131), .ZN(n14122) );
  NOR3_X1 U15744 ( .A1(n14119), .A2(n14118), .A3(n14117), .ZN(n14121) );
  XNOR2_X1 U15745 ( .A(n14132), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n14140) );
  NAND2_X1 U15746 ( .A1(n14131), .A2(n14130), .ZN(n14133) );
  XNOR2_X1 U15747 ( .A(n14132), .B(P3_REG2_REG_19__SCAN_IN), .ZN(n14141) );
  NAND2_X1 U15748 ( .A1(n16150), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n14134) );
  OAI21_X1 U15749 ( .B1(n14138), .B2(n14137), .A(n14136), .ZN(n14143) );
  MUX2_X1 U15750 ( .A(n14141), .B(n14140), .S(n14139), .Z(n14142) );
  XNOR2_X1 U15751 ( .A(n14143), .B(n14142), .ZN(n14144) );
  NOR2_X1 U15752 ( .A1(n14144), .A2(n16418), .ZN(n14145) );
  INV_X1 U15753 ( .A(n14149), .ZN(n14150) );
  NAND2_X1 U15754 ( .A1(n14151), .A2(n14150), .ZN(n14838) );
  INV_X1 U15755 ( .A(n14838), .ZN(n14153) );
  NOR3_X1 U15756 ( .A1(n14153), .A2(n16517), .A3(n14152), .ZN(n14156) );
  NOR2_X1 U15757 ( .A1(n14352), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n14154) );
  OAI22_X1 U15758 ( .A1(n14840), .A2(n14384), .B1(n14156), .B2(n14154), .ZN(
        P3_U3202) );
  NOR2_X1 U15759 ( .A1(n14352), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n14155) );
  OAI22_X1 U15760 ( .A1(n14156), .A2(n14155), .B1(n14843), .B2(n14384), .ZN(
        P3_U3203) );
  AOI21_X1 U15761 ( .B1(n14157), .B2(n14163), .A(n14310), .ZN(n14161) );
  OAI22_X1 U15762 ( .A1(n14158), .A2(n14314), .B1(n14184), .B2(n14312), .ZN(
        n14159) );
  AOI21_X1 U15763 ( .B1(n14161), .B2(n14160), .A(n14159), .ZN(n14395) );
  OAI21_X1 U15764 ( .B1(n14164), .B2(n14163), .A(n14162), .ZN(n14393) );
  AOI22_X1 U15765 ( .A1(n16517), .A2(P3_REG2_REG_28__SCAN_IN), .B1(n14369), 
        .B2(n14165), .ZN(n14166) );
  OAI21_X1 U15766 ( .B1(n14167), .B2(n14384), .A(n14166), .ZN(n14168) );
  AOI21_X1 U15767 ( .B1(n14393), .B2(n14372), .A(n14168), .ZN(n14169) );
  OAI21_X1 U15768 ( .B1(n14395), .B2(n16517), .A(n14169), .ZN(P3_U3205) );
  OAI21_X1 U15769 ( .B1(n14171), .B2(n7851), .A(n14170), .ZN(n14181) );
  INV_X1 U15770 ( .A(n14181), .ZN(n14845) );
  OAI21_X1 U15771 ( .B1(n14174), .B2(n14173), .A(n14172), .ZN(n14177) );
  AOI222_X1 U15772 ( .A1(n16501), .A2(n14177), .B1(n14176), .B2(n16498), .C1(
        n14175), .C2(n16495), .ZN(n14396) );
  OAI21_X1 U15773 ( .B1(n16521), .B2(n14845), .A(n14396), .ZN(n14847) );
  INV_X1 U15774 ( .A(n14847), .ZN(n14183) );
  AOI22_X1 U15775 ( .A1(n16517), .A2(P3_REG2_REG_27__SCAN_IN), .B1(n14369), 
        .B2(n14178), .ZN(n14179) );
  OAI21_X1 U15776 ( .B1(n14850), .B2(n14384), .A(n14179), .ZN(n14180) );
  AOI21_X1 U15777 ( .B1(n14181), .B2(n14240), .A(n14180), .ZN(n14182) );
  OAI21_X1 U15778 ( .B1(n14183), .B2(n16517), .A(n14182), .ZN(P3_U3206) );
  INV_X1 U15779 ( .A(n14401), .ZN(n14191) );
  XOR2_X1 U15780 ( .A(n14186), .B(n14185), .Z(n14402) );
  AOI22_X1 U15781 ( .A1(n16517), .A2(P3_REG2_REG_26__SCAN_IN), .B1(n14187), 
        .B2(n14369), .ZN(n14188) );
  OAI21_X1 U15782 ( .B1(n14854), .B2(n14384), .A(n14188), .ZN(n14189) );
  AOI21_X1 U15783 ( .B1(n14402), .B2(n14372), .A(n14189), .ZN(n14190) );
  OAI21_X1 U15784 ( .B1(n14191), .B2(n16517), .A(n14190), .ZN(P3_U3207) );
  OAI211_X1 U15785 ( .C1(n14194), .C2(n14193), .A(n14192), .B(n16501), .ZN(
        n14197) );
  NAND2_X1 U15786 ( .A1(n14195), .A2(n16498), .ZN(n14196) );
  OAI211_X1 U15787 ( .C1(n14198), .C2(n14314), .A(n14197), .B(n14196), .ZN(
        n14405) );
  INV_X1 U15788 ( .A(n14405), .ZN(n14204) );
  XNOR2_X1 U15789 ( .A(n14199), .B(n8347), .ZN(n14406) );
  AOI22_X1 U15790 ( .A1(n16517), .A2(P3_REG2_REG_25__SCAN_IN), .B1(n14369), 
        .B2(n14200), .ZN(n14201) );
  OAI21_X1 U15791 ( .B1(n8351), .B2(n14384), .A(n14201), .ZN(n14202) );
  AOI21_X1 U15792 ( .B1(n14406), .B2(n14372), .A(n14202), .ZN(n14203) );
  OAI21_X1 U15793 ( .B1(n14204), .B2(n16517), .A(n14203), .ZN(P3_U3208) );
  XNOR2_X1 U15794 ( .A(n14206), .B(n14205), .ZN(n14207) );
  OAI222_X1 U15795 ( .A1(n14314), .A2(n14209), .B1(n14312), .B2(n14208), .C1(
        n14207), .C2(n14310), .ZN(n14409) );
  INV_X1 U15796 ( .A(n14409), .ZN(n14215) );
  XNOR2_X1 U15797 ( .A(n14210), .B(n8349), .ZN(n14410) );
  AOI22_X1 U15798 ( .A1(n16517), .A2(P3_REG2_REG_24__SCAN_IN), .B1(n14369), 
        .B2(n14211), .ZN(n14212) );
  OAI21_X1 U15799 ( .B1(n14861), .B2(n14384), .A(n14212), .ZN(n14213) );
  AOI21_X1 U15800 ( .B1(n14410), .B2(n14372), .A(n14213), .ZN(n14214) );
  OAI21_X1 U15801 ( .B1(n14215), .B2(n16517), .A(n14214), .ZN(P3_U3209) );
  XNOR2_X1 U15802 ( .A(n14217), .B(n14216), .ZN(n14218) );
  OAI222_X1 U15803 ( .A1(n14314), .A2(n14220), .B1(n14312), .B2(n14219), .C1(
        n14218), .C2(n14310), .ZN(n14413) );
  INV_X1 U15804 ( .A(n14413), .ZN(n14227) );
  XNOR2_X1 U15805 ( .A(n14222), .B(n14221), .ZN(n14414) );
  AOI22_X1 U15806 ( .A1(n16517), .A2(P3_REG2_REG_23__SCAN_IN), .B1(n14369), 
        .B2(n14223), .ZN(n14224) );
  OAI21_X1 U15807 ( .B1(n14865), .B2(n14384), .A(n14224), .ZN(n14225) );
  AOI21_X1 U15808 ( .B1(n14414), .B2(n14372), .A(n14225), .ZN(n14226) );
  OAI21_X1 U15809 ( .B1(n14227), .B2(n16517), .A(n14226), .ZN(P3_U3210) );
  XNOR2_X1 U15810 ( .A(n14228), .B(n14230), .ZN(n14236) );
  XOR2_X1 U15811 ( .A(n14230), .B(n14229), .Z(n14231) );
  NAND2_X1 U15812 ( .A1(n14231), .A2(n16501), .ZN(n14235) );
  AOI22_X1 U15813 ( .A1(n14233), .A2(n16498), .B1(n14232), .B2(n16495), .ZN(
        n14234) );
  OAI211_X1 U15814 ( .C1(n16521), .C2(n14236), .A(n14235), .B(n14234), .ZN(
        n14417) );
  INV_X1 U15815 ( .A(n14417), .ZN(n14242) );
  INV_X1 U15816 ( .A(n14236), .ZN(n14418) );
  AOI22_X1 U15817 ( .A1(n16517), .A2(P3_REG2_REG_22__SCAN_IN), .B1(n14369), 
        .B2(n14237), .ZN(n14238) );
  OAI21_X1 U15818 ( .B1(n14869), .B2(n14384), .A(n14238), .ZN(n14239) );
  AOI21_X1 U15819 ( .B1(n14418), .B2(n14240), .A(n14239), .ZN(n14241) );
  OAI21_X1 U15820 ( .B1(n14242), .B2(n16517), .A(n14241), .ZN(P3_U3211) );
  XNOR2_X1 U15821 ( .A(n14243), .B(n14245), .ZN(n14422) );
  INV_X1 U15822 ( .A(n14422), .ZN(n14256) );
  XOR2_X1 U15823 ( .A(n14245), .B(n14244), .Z(n14249) );
  AOI22_X1 U15824 ( .A1(n8153), .A2(n16498), .B1(n16495), .B2(n14246), .ZN(
        n14248) );
  INV_X1 U15825 ( .A(n16521), .ZN(n16620) );
  NAND2_X1 U15826 ( .A1(n14422), .A2(n16620), .ZN(n14247) );
  OAI211_X1 U15827 ( .C1(n14249), .C2(n14310), .A(n14248), .B(n14247), .ZN(
        n14421) );
  NAND2_X1 U15828 ( .A1(n14421), .A2(n14352), .ZN(n14255) );
  INV_X1 U15829 ( .A(P3_REG2_REG_21__SCAN_IN), .ZN(n14251) );
  OAI22_X1 U15830 ( .A1(n14352), .A2(n14251), .B1(n14250), .B2(n16508), .ZN(
        n14252) );
  AOI21_X1 U15831 ( .B1(n14253), .B2(n14354), .A(n14252), .ZN(n14254) );
  OAI211_X1 U15832 ( .C1(n14256), .C2(n14388), .A(n14255), .B(n14254), .ZN(
        P3_U3212) );
  NAND2_X1 U15833 ( .A1(n14258), .A2(n14257), .ZN(n14292) );
  NAND2_X1 U15834 ( .A1(n14292), .A2(n14259), .ZN(n14283) );
  NAND2_X1 U15835 ( .A1(n14283), .A2(n14260), .ZN(n14261) );
  XNOR2_X1 U15836 ( .A(n14261), .B(n14262), .ZN(n14426) );
  INV_X1 U15837 ( .A(n14426), .ZN(n14275) );
  XNOR2_X1 U15838 ( .A(n14263), .B(n14262), .ZN(n14268) );
  OAI22_X1 U15839 ( .A1(n14265), .A2(n14314), .B1(n14264), .B2(n14312), .ZN(
        n14266) );
  AOI21_X1 U15840 ( .B1(n14426), .B2(n16620), .A(n14266), .ZN(n14267) );
  OAI21_X1 U15841 ( .B1(n14268), .B2(n14310), .A(n14267), .ZN(n14425) );
  NAND2_X1 U15842 ( .A1(n14425), .A2(n14352), .ZN(n14274) );
  INV_X1 U15843 ( .A(P3_REG2_REG_20__SCAN_IN), .ZN(n14270) );
  OAI22_X1 U15844 ( .A1(n14352), .A2(n14270), .B1(n14269), .B2(n16508), .ZN(
        n14271) );
  AOI21_X1 U15845 ( .B1(n14272), .B2(n14354), .A(n14271), .ZN(n14273) );
  OAI211_X1 U15846 ( .C1(n14275), .C2(n14388), .A(n14274), .B(n14273), .ZN(
        P3_U3213) );
  XOR2_X1 U15847 ( .A(n14285), .B(n14276), .Z(n14277) );
  OAI222_X1 U15848 ( .A1(n14312), .A2(n14313), .B1(n14314), .B2(n14278), .C1(
        n14310), .C2(n14277), .ZN(n14429) );
  INV_X1 U15849 ( .A(n14429), .ZN(n14291) );
  NAND2_X1 U15850 ( .A1(n14292), .A2(n14279), .ZN(n14281) );
  NAND2_X1 U15851 ( .A1(n14281), .A2(n14280), .ZN(n14286) );
  AND2_X1 U15852 ( .A1(n14283), .A2(n14282), .ZN(n14284) );
  OAI21_X1 U15853 ( .B1(n14286), .B2(n14285), .A(n14284), .ZN(n14430) );
  AOI22_X1 U15854 ( .A1(n16517), .A2(P3_REG2_REG_19__SCAN_IN), .B1(n14369), 
        .B2(n14287), .ZN(n14288) );
  OAI21_X1 U15855 ( .B1(n14881), .B2(n14384), .A(n14288), .ZN(n14289) );
  AOI21_X1 U15856 ( .B1(n14430), .B2(n14372), .A(n14289), .ZN(n14290) );
  OAI21_X1 U15857 ( .B1(n14291), .B2(n16517), .A(n14290), .ZN(P3_U3214) );
  XNOR2_X1 U15858 ( .A(n14292), .B(n14293), .ZN(n14434) );
  NOR2_X1 U15859 ( .A1(n14294), .A2(n14293), .ZN(n14295) );
  OR2_X1 U15860 ( .A1(n14296), .A2(n14295), .ZN(n14297) );
  NAND2_X1 U15861 ( .A1(n14297), .A2(n16501), .ZN(n14300) );
  AOI22_X1 U15862 ( .A1(n14298), .A2(n16495), .B1(n16498), .B2(n14328), .ZN(
        n14299) );
  NAND2_X1 U15863 ( .A1(n14300), .A2(n14299), .ZN(n14436) );
  NAND2_X1 U15864 ( .A1(n14436), .A2(n14352), .ZN(n14306) );
  OAI22_X1 U15865 ( .A1(n14352), .A2(n14302), .B1(n14301), .B2(n16508), .ZN(
        n14303) );
  AOI21_X1 U15866 ( .B1(n14304), .B2(n14354), .A(n14303), .ZN(n14305) );
  OAI211_X1 U15867 ( .C1(n14434), .C2(n14358), .A(n14306), .B(n14305), .ZN(
        P3_U3215) );
  XNOR2_X1 U15868 ( .A(n14308), .B(n14307), .ZN(n14309) );
  OAI222_X1 U15869 ( .A1(n14314), .A2(n14313), .B1(n14312), .B2(n14311), .C1(
        n14310), .C2(n14309), .ZN(n14437) );
  INV_X1 U15870 ( .A(n14437), .ZN(n14325) );
  OR2_X1 U15871 ( .A1(n14315), .A2(n14316), .ZN(n14318) );
  NAND2_X1 U15872 ( .A1(n14318), .A2(n14317), .ZN(n14320) );
  XNOR2_X1 U15873 ( .A(n14320), .B(n14319), .ZN(n14438) );
  NOR2_X1 U15874 ( .A1(n14886), .A2(n14384), .ZN(n14323) );
  OAI22_X1 U15875 ( .A1(n14352), .A2(n8426), .B1(n14321), .B2(n16508), .ZN(
        n14322) );
  AOI211_X1 U15876 ( .C1(n14438), .C2(n14372), .A(n14323), .B(n14322), .ZN(
        n14324) );
  OAI21_X1 U15877 ( .B1(n14325), .B2(n16517), .A(n14324), .ZN(P3_U3216) );
  XNOR2_X1 U15878 ( .A(n14327), .B(n14326), .ZN(n14329) );
  AOI222_X1 U15879 ( .A1(n16501), .A2(n14329), .B1(n14328), .B2(n16495), .C1(
        n14363), .C2(n16498), .ZN(n14444) );
  OR2_X1 U15880 ( .A1(n14315), .A2(n14344), .ZN(n14331) );
  NAND2_X1 U15881 ( .A1(n14331), .A2(n14330), .ZN(n14333) );
  XNOR2_X1 U15882 ( .A(n14333), .B(n14332), .ZN(n14442) );
  NOR2_X1 U15883 ( .A1(n14334), .A2(n14384), .ZN(n14338) );
  INV_X1 U15884 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n14336) );
  OAI22_X1 U15885 ( .A1(n14352), .A2(n14336), .B1(n14335), .B2(n16508), .ZN(
        n14337) );
  AOI211_X1 U15886 ( .C1(n14442), .C2(n14372), .A(n14338), .B(n14337), .ZN(
        n14339) );
  OAI21_X1 U15887 ( .B1(n14444), .B2(n16517), .A(n14339), .ZN(P3_U3217) );
  INV_X1 U15888 ( .A(n14344), .ZN(n14340) );
  XNOR2_X1 U15889 ( .A(n14315), .B(n14340), .ZN(n14446) );
  AND2_X1 U15890 ( .A1(n14360), .A2(n14341), .ZN(n14345) );
  NAND2_X1 U15891 ( .A1(n14360), .A2(n14342), .ZN(n14343) );
  OAI21_X1 U15892 ( .B1(n14345), .B2(n14344), .A(n14343), .ZN(n14346) );
  NAND2_X1 U15893 ( .A1(n14346), .A2(n16501), .ZN(n14350) );
  AOI22_X1 U15894 ( .A1(n14348), .A2(n16495), .B1(n16498), .B2(n14347), .ZN(
        n14349) );
  NAND2_X1 U15895 ( .A1(n14350), .A2(n14349), .ZN(n14448) );
  NAND2_X1 U15896 ( .A1(n14448), .A2(n14352), .ZN(n14357) );
  INV_X1 U15897 ( .A(n14445), .ZN(n14355) );
  OAI22_X1 U15898 ( .A1(n14352), .A2(n8435), .B1(n14351), .B2(n16508), .ZN(
        n14353) );
  AOI21_X1 U15899 ( .B1(n14355), .B2(n14354), .A(n14353), .ZN(n14356) );
  OAI211_X1 U15900 ( .C1(n14446), .C2(n14358), .A(n14357), .B(n14356), .ZN(
        P3_U3218) );
  INV_X1 U15901 ( .A(n14359), .ZN(n14362) );
  OAI211_X1 U15902 ( .C1(n14362), .C2(n14361), .A(n14360), .B(n16501), .ZN(
        n14365) );
  AOI22_X1 U15903 ( .A1(n16495), .A2(n14363), .B1(n14379), .B2(n16498), .ZN(
        n14364) );
  NAND2_X1 U15904 ( .A1(n14365), .A2(n14364), .ZN(n14451) );
  INV_X1 U15905 ( .A(n14451), .ZN(n14374) );
  XNOR2_X1 U15906 ( .A(n14367), .B(n14366), .ZN(n14452) );
  AOI22_X1 U15907 ( .A1(n16517), .A2(P3_REG2_REG_14__SCAN_IN), .B1(n14369), 
        .B2(n14368), .ZN(n14370) );
  OAI21_X1 U15908 ( .B1(n14895), .B2(n14384), .A(n14370), .ZN(n14371) );
  AOI21_X1 U15909 ( .B1(n14452), .B2(n14372), .A(n14371), .ZN(n14373) );
  OAI21_X1 U15910 ( .B1(n14374), .B2(n16517), .A(n14373), .ZN(P3_U3219) );
  XNOR2_X1 U15911 ( .A(n14375), .B(n14376), .ZN(n14832) );
  XNOR2_X1 U15912 ( .A(n14377), .B(n14376), .ZN(n14378) );
  NAND2_X1 U15913 ( .A1(n14378), .A2(n16501), .ZN(n14382) );
  AOI22_X1 U15914 ( .A1(n16498), .A2(n14380), .B1(n14379), .B2(n16495), .ZN(
        n14381) );
  OAI211_X1 U15915 ( .C1(n16521), .C2(n14832), .A(n14382), .B(n14381), .ZN(
        n14834) );
  NAND2_X1 U15916 ( .A1(n14834), .A2(n14352), .ZN(n14387) );
  OAI22_X1 U15917 ( .A1(n14384), .A2(n14831), .B1(n14383), .B2(n16508), .ZN(
        n14385) );
  AOI21_X1 U15918 ( .B1(P3_REG2_REG_12__SCAN_IN), .B2(n16517), .A(n14385), 
        .ZN(n14386) );
  OAI211_X1 U15919 ( .C1(n14388), .C2(n14832), .A(n14387), .B(n14386), .ZN(
        P3_U3221) );
  NOR2_X1 U15920 ( .A1(n16717), .A2(n14838), .ZN(n14390) );
  AOI21_X1 U15921 ( .B1(n16717), .B2(P3_REG1_REG_31__SCAN_IN), .A(n14390), 
        .ZN(n14389) );
  OAI21_X1 U15922 ( .B1(n14840), .B2(n14455), .A(n14389), .ZN(P3_U3490) );
  AOI21_X1 U15923 ( .B1(n16717), .B2(P3_REG1_REG_30__SCAN_IN), .A(n14390), 
        .ZN(n14391) );
  OAI21_X1 U15924 ( .B1(n14455), .B2(n14843), .A(n14391), .ZN(P3_U3489) );
  AOI22_X1 U15925 ( .A1(n14393), .A2(n16647), .B1(n16652), .B2(n14392), .ZN(
        n14394) );
  NAND2_X1 U15926 ( .A1(n14395), .A2(n14394), .ZN(n14844) );
  MUX2_X1 U15927 ( .A(P3_REG1_REG_28__SCAN_IN), .B(n14844), .S(n16718), .Z(
        P3_U3487) );
  OAI21_X1 U15928 ( .B1(n16713), .B2(n14845), .A(n14396), .ZN(n14399) );
  OAI22_X1 U15929 ( .A1(n14850), .A2(n14455), .B1(n16718), .B2(n14397), .ZN(
        n14398) );
  AOI21_X1 U15930 ( .B1(n14399), .B2(n16718), .A(n14398), .ZN(n14400) );
  INV_X1 U15931 ( .A(n14400), .ZN(P3_U3486) );
  AOI21_X1 U15932 ( .B1(n16647), .B2(n14402), .A(n14401), .ZN(n14851) );
  MUX2_X1 U15933 ( .A(n14403), .B(n14851), .S(n16718), .Z(n14404) );
  OAI21_X1 U15934 ( .B1(n14854), .B2(n14455), .A(n14404), .ZN(P3_U3485) );
  AOI21_X1 U15935 ( .B1(n14406), .B2(n16647), .A(n14405), .ZN(n14855) );
  MUX2_X1 U15936 ( .A(n14407), .B(n14855), .S(n16718), .Z(n14408) );
  OAI21_X1 U15937 ( .B1(n8351), .B2(n14455), .A(n14408), .ZN(P3_U3484) );
  INV_X1 U15938 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n14411) );
  AOI21_X1 U15939 ( .B1(n16647), .B2(n14410), .A(n14409), .ZN(n14858) );
  MUX2_X1 U15940 ( .A(n14411), .B(n14858), .S(n16718), .Z(n14412) );
  OAI21_X1 U15941 ( .B1(n14861), .B2(n14455), .A(n14412), .ZN(P3_U3483) );
  AOI21_X1 U15942 ( .B1(n16647), .B2(n14414), .A(n14413), .ZN(n14862) );
  MUX2_X1 U15943 ( .A(n14415), .B(n14862), .S(n16718), .Z(n14416) );
  OAI21_X1 U15944 ( .B1(n14865), .B2(n14455), .A(n14416), .ZN(P3_U3482) );
  AOI21_X1 U15945 ( .B1(n16596), .B2(n14418), .A(n14417), .ZN(n14866) );
  MUX2_X1 U15946 ( .A(n14419), .B(n14866), .S(n16718), .Z(n14420) );
  OAI21_X1 U15947 ( .B1(n14869), .B2(n14455), .A(n14420), .ZN(P3_U3481) );
  AOI21_X1 U15948 ( .B1(n16596), .B2(n14422), .A(n14421), .ZN(n14870) );
  MUX2_X1 U15949 ( .A(n14423), .B(n14870), .S(n16718), .Z(n14424) );
  OAI21_X1 U15950 ( .B1(n14873), .B2(n14455), .A(n14424), .ZN(P3_U3480) );
  AOI21_X1 U15951 ( .B1(n16596), .B2(n14426), .A(n14425), .ZN(n14874) );
  MUX2_X1 U15952 ( .A(n14427), .B(n14874), .S(n16718), .Z(n14428) );
  OAI21_X1 U15953 ( .B1(n14877), .B2(n14455), .A(n14428), .ZN(P3_U3479) );
  AOI21_X1 U15954 ( .B1(n16647), .B2(n14430), .A(n14429), .ZN(n14878) );
  MUX2_X1 U15955 ( .A(n14431), .B(n14878), .S(n16718), .Z(n14432) );
  OAI21_X1 U15956 ( .B1(n14881), .B2(n14455), .A(n14432), .ZN(P3_U3478) );
  OAI22_X1 U15957 ( .A1(n14434), .A2(n16713), .B1(n14433), .B2(n16711), .ZN(
        n14435) );
  MUX2_X1 U15958 ( .A(n14882), .B(P3_REG1_REG_18__SCAN_IN), .S(n16717), .Z(
        P3_U3477) );
  AOI21_X1 U15959 ( .B1(n14438), .B2(n16647), .A(n14437), .ZN(n14883) );
  MUX2_X1 U15960 ( .A(n14439), .B(n14883), .S(n16718), .Z(n14440) );
  OAI21_X1 U15961 ( .B1(n14455), .B2(n14886), .A(n14440), .ZN(P3_U3476) );
  AOI22_X1 U15962 ( .A1(n14442), .A2(n16647), .B1(n16652), .B2(n14441), .ZN(
        n14443) );
  NAND2_X1 U15963 ( .A1(n14444), .A2(n14443), .ZN(n14887) );
  MUX2_X1 U15964 ( .A(P3_REG1_REG_16__SCAN_IN), .B(n14887), .S(n16718), .Z(
        P3_U3475) );
  OAI22_X1 U15965 ( .A1(n14446), .A2(n16713), .B1(n14445), .B2(n16711), .ZN(
        n14447) );
  NOR2_X1 U15966 ( .A1(n14448), .A2(n14447), .ZN(n14888) );
  MUX2_X1 U15967 ( .A(n14449), .B(n14888), .S(n16718), .Z(n14450) );
  INV_X1 U15968 ( .A(n14450), .ZN(P3_U3474) );
  AOI21_X1 U15969 ( .B1(n14452), .B2(n16647), .A(n14451), .ZN(n14892) );
  MUX2_X1 U15970 ( .A(n14453), .B(n14892), .S(n16718), .Z(n14454) );
  OAI21_X1 U15971 ( .B1(n14455), .B2(n14895), .A(n14454), .ZN(P3_U3473) );
  OAI22_X1 U15972 ( .A1(n10452), .A2(keyinput_120), .B1(keyinput_119), .B2(
        P1_IR_REG_12__SCAN_IN), .ZN(n14456) );
  AOI221_X1 U15973 ( .B1(n10452), .B2(keyinput_120), .C1(P1_IR_REG_12__SCAN_IN), .C2(keyinput_119), .A(n14456), .ZN(n14619) );
  INV_X1 U15974 ( .A(keyinput_118), .ZN(n14615) );
  INV_X1 U15975 ( .A(keyinput_117), .ZN(n14614) );
  INV_X1 U15976 ( .A(keyinput_110), .ZN(n14605) );
  INV_X1 U15977 ( .A(keyinput_106), .ZN(n14598) );
  INV_X1 U15978 ( .A(keyinput_105), .ZN(n14597) );
  INV_X1 U15979 ( .A(keyinput_104), .ZN(n14596) );
  INV_X1 U15980 ( .A(keyinput_103), .ZN(n14595) );
  OAI22_X1 U15981 ( .A1(n16281), .A2(keyinput_99), .B1(keyinput_100), .B2(
        P3_ADDR_REG_3__SCAN_IN), .ZN(n14457) );
  AOI221_X1 U15982 ( .B1(n16281), .B2(keyinput_99), .C1(P3_ADDR_REG_3__SCAN_IN), .C2(keyinput_100), .A(n14457), .ZN(n14593) );
  XOR2_X1 U15983 ( .A(P3_DATAO_REG_11__SCAN_IN), .B(keyinput_85), .Z(n14576)
         );
  OAI22_X1 U15984 ( .A1(n14459), .A2(keyinput_87), .B1(keyinput_86), .B2(
        P3_DATAO_REG_10__SCAN_IN), .ZN(n14458) );
  AOI221_X1 U15985 ( .B1(n14459), .B2(keyinput_87), .C1(
        P3_DATAO_REG_10__SCAN_IN), .C2(keyinput_86), .A(n14458), .ZN(n14575)
         );
  OAI22_X1 U15986 ( .A1(n14461), .A2(keyinput_88), .B1(P3_DATAO_REG_7__SCAN_IN), .B2(keyinput_89), .ZN(n14460) );
  AOI221_X1 U15987 ( .B1(n14461), .B2(keyinput_88), .C1(keyinput_89), .C2(
        P3_DATAO_REG_7__SCAN_IN), .A(n14460), .ZN(n14574) );
  INV_X1 U15988 ( .A(keyinput_84), .ZN(n14572) );
  OAI22_X1 U15989 ( .A1(P3_DATAO_REG_21__SCAN_IN), .A2(keyinput_75), .B1(
        P3_DATAO_REG_20__SCAN_IN), .B2(keyinput_76), .ZN(n14462) );
  AOI221_X1 U15990 ( .B1(P3_DATAO_REG_21__SCAN_IN), .B2(keyinput_75), .C1(
        keyinput_76), .C2(P3_DATAO_REG_20__SCAN_IN), .A(n14462), .ZN(n14569)
         );
  AOI22_X1 U15991 ( .A1(n14732), .A2(keyinput_68), .B1(n14728), .B2(
        keyinput_65), .ZN(n14463) );
  OAI221_X1 U15992 ( .B1(n14732), .B2(keyinput_68), .C1(n14728), .C2(
        keyinput_65), .A(n14463), .ZN(n14560) );
  INV_X1 U15993 ( .A(P3_DATAO_REG_30__SCAN_IN), .ZN(n14725) );
  OAI22_X1 U15994 ( .A1(n14725), .A2(keyinput_66), .B1(n14465), .B2(
        keyinput_70), .ZN(n14464) );
  AOI221_X1 U15995 ( .B1(n14725), .B2(keyinput_66), .C1(keyinput_70), .C2(
        n14465), .A(n14464), .ZN(n14556) );
  OAI22_X1 U15996 ( .A1(P3_DATAO_REG_27__SCAN_IN), .A2(keyinput_69), .B1(
        keyinput_67), .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n14466) );
  AOI221_X1 U15997 ( .B1(P3_DATAO_REG_27__SCAN_IN), .B2(keyinput_69), .C1(
        P3_DATAO_REG_29__SCAN_IN), .C2(keyinput_67), .A(n14466), .ZN(n14555)
         );
  OAI22_X1 U15998 ( .A1(n14468), .A2(keyinput_71), .B1(keyinput_72), .B2(
        P3_DATAO_REG_24__SCAN_IN), .ZN(n14467) );
  AOI221_X1 U15999 ( .B1(n14468), .B2(keyinput_71), .C1(
        P3_DATAO_REG_24__SCAN_IN), .C2(keyinput_72), .A(n14467), .ZN(n14554)
         );
  XNOR2_X1 U16000 ( .A(keyinput_60), .B(n14738), .ZN(n14552) );
  OAI22_X1 U16001 ( .A1(n14470), .A2(keyinput_63), .B1(keyinput_62), .B2(
        P3_REG3_REG_26__SCAN_IN), .ZN(n14469) );
  AOI221_X1 U16002 ( .B1(n14470), .B2(keyinput_63), .C1(
        P3_REG3_REG_26__SCAN_IN), .C2(keyinput_62), .A(n14469), .ZN(n14551) );
  OAI22_X1 U16003 ( .A1(n14741), .A2(keyinput_61), .B1(P3_B_REG_SCAN_IN), .B2(
        keyinput_64), .ZN(n14471) );
  AOI221_X1 U16004 ( .B1(n14741), .B2(keyinput_61), .C1(keyinput_64), .C2(
        P3_B_REG_SCAN_IN), .A(n14471), .ZN(n14550) );
  INV_X1 U16005 ( .A(keyinput_59), .ZN(n14548) );
  INV_X1 U16006 ( .A(keyinput_49), .ZN(n14533) );
  INV_X1 U16007 ( .A(keyinput_48), .ZN(n14532) );
  AOI22_X1 U16008 ( .A1(P3_REG3_REG_12__SCAN_IN), .A2(keyinput_46), .B1(n14641), .B2(keyinput_45), .ZN(n14472) );
  OAI221_X1 U16009 ( .B1(P3_REG3_REG_12__SCAN_IN), .B2(keyinput_46), .C1(
        n14641), .C2(keyinput_45), .A(n14472), .ZN(n14531) );
  OAI22_X1 U16010 ( .A1(n14474), .A2(keyinput_40), .B1(P3_REG3_REG_19__SCAN_IN), .B2(keyinput_41), .ZN(n14473) );
  AOI221_X1 U16011 ( .B1(n14474), .B2(keyinput_40), .C1(keyinput_41), .C2(
        P3_REG3_REG_19__SCAN_IN), .A(n14473), .ZN(n14529) );
  INV_X1 U16012 ( .A(keyinput_35), .ZN(n14518) );
  INV_X1 U16013 ( .A(keyinput_21), .ZN(n14503) );
  INV_X1 U16014 ( .A(keyinput_20), .ZN(n14501) );
  OAI22_X1 U16015 ( .A1(n14647), .A2(keyinput_18), .B1(SI_15_), .B2(
        keyinput_17), .ZN(n14475) );
  AOI221_X1 U16016 ( .B1(n14647), .B2(keyinput_18), .C1(keyinput_17), .C2(
        SI_15_), .A(n14475), .ZN(n14498) );
  INV_X1 U16017 ( .A(keyinput_12), .ZN(n14490) );
  INV_X1 U16018 ( .A(keyinput_11), .ZN(n14489) );
  OAI22_X1 U16019 ( .A1(n14919), .A2(keyinput_4), .B1(n14477), .B2(keyinput_5), 
        .ZN(n14476) );
  AOI221_X1 U16020 ( .B1(n14919), .B2(keyinput_4), .C1(keyinput_5), .C2(n14477), .A(n14476), .ZN(n14488) );
  OAI221_X1 U16021 ( .B1(SI_29_), .B2(keyinput_3), .C1(n14910), .C2(keyinput_2), .A(n14478), .ZN(n14481) );
  OAI22_X1 U16022 ( .A1(SI_31_), .A2(keyinput_1), .B1(P3_WR_REG_SCAN_IN), .B2(
        keyinput_0), .ZN(n14479) );
  OAI22_X1 U16023 ( .A1(n14481), .A2(n14480), .B1(n14483), .B2(keyinput_6), 
        .ZN(n14482) );
  AOI22_X1 U16024 ( .A1(SI_24_), .A2(keyinput_8), .B1(SI_25_), .B2(keyinput_7), 
        .ZN(n14484) );
  OAI221_X1 U16025 ( .B1(SI_24_), .B2(keyinput_8), .C1(SI_25_), .C2(keyinput_7), .A(n14484), .ZN(n14487) );
  AOI22_X1 U16026 ( .A1(SI_22_), .A2(keyinput_10), .B1(SI_23_), .B2(keyinput_9), .ZN(n14485) );
  OAI221_X1 U16027 ( .B1(SI_22_), .B2(keyinput_10), .C1(SI_23_), .C2(
        keyinput_9), .A(n14485), .ZN(n14486) );
  AOI22_X1 U16028 ( .A1(n14492), .A2(keyinput_14), .B1(n14666), .B2(
        keyinput_13), .ZN(n14491) );
  OAI221_X1 U16029 ( .B1(n14492), .B2(keyinput_14), .C1(n14666), .C2(
        keyinput_13), .A(n14491), .ZN(n14495) );
  OAI22_X1 U16030 ( .A1(SI_17_), .A2(keyinput_15), .B1(SI_16_), .B2(
        keyinput_16), .ZN(n14493) );
  AOI221_X1 U16031 ( .B1(SI_17_), .B2(keyinput_15), .C1(keyinput_16), .C2(
        SI_16_), .A(n14493), .ZN(n14494) );
  AOI22_X1 U16032 ( .A1(keyinput_19), .A2(n14674), .B1(n14498), .B2(n14497), 
        .ZN(n14499) );
  OAI21_X1 U16033 ( .B1(n14674), .B2(keyinput_19), .A(n14499), .ZN(n14500) );
  OAI221_X1 U16034 ( .B1(SI_12_), .B2(keyinput_20), .C1(n14676), .C2(n14501), 
        .A(n14500), .ZN(n14502) );
  OAI221_X1 U16035 ( .B1(SI_11_), .B2(n14503), .C1(n14679), .C2(keyinput_21), 
        .A(n14502), .ZN(n14510) );
  XNOR2_X1 U16036 ( .A(keyinput_22), .B(n14680), .ZN(n14509) );
  XOR2_X1 U16037 ( .A(SI_8_), .B(keyinput_24), .Z(n14507) );
  XNOR2_X1 U16038 ( .A(SI_7_), .B(keyinput_25), .ZN(n14506) );
  XNOR2_X1 U16039 ( .A(SI_6_), .B(keyinput_26), .ZN(n14505) );
  XNOR2_X1 U16040 ( .A(SI_9_), .B(keyinput_23), .ZN(n14504) );
  NAND4_X1 U16041 ( .A1(n14507), .A2(n14506), .A3(n14505), .A4(n14504), .ZN(
        n14508) );
  AOI21_X1 U16042 ( .B1(n14510), .B2(n14509), .A(n14508), .ZN(n14511) );
  XOR2_X1 U16043 ( .A(SI_1_), .B(keyinput_31), .Z(n14514) );
  XOR2_X1 U16044 ( .A(SI_2_), .B(keyinput_30), .Z(n14513) );
  XNOR2_X1 U16045 ( .A(SI_3_), .B(keyinput_29), .ZN(n14512) );
  XOR2_X1 U16046 ( .A(P3_RD_REG_SCAN_IN), .B(keyinput_33), .Z(n14516) );
  XNOR2_X1 U16047 ( .A(SI_0_), .B(keyinput_32), .ZN(n14515) );
  AOI221_X1 U16048 ( .B1(P3_REG3_REG_7__SCAN_IN), .B2(n14518), .C1(n8861), 
        .C2(keyinput_35), .A(n14517), .ZN(n14523) );
  AOI22_X1 U16049 ( .A1(P3_REG3_REG_14__SCAN_IN), .A2(keyinput_37), .B1(
        P3_REG3_REG_27__SCAN_IN), .B2(keyinput_36), .ZN(n14519) );
  OAI221_X1 U16050 ( .B1(P3_REG3_REG_14__SCAN_IN), .B2(keyinput_37), .C1(
        P3_REG3_REG_27__SCAN_IN), .C2(keyinput_36), .A(n14519), .ZN(n14522) );
  OAI22_X1 U16051 ( .A1(P3_REG3_REG_23__SCAN_IN), .A2(keyinput_38), .B1(
        keyinput_39), .B2(P3_REG3_REG_10__SCAN_IN), .ZN(n14520) );
  AOI221_X1 U16052 ( .B1(P3_REG3_REG_23__SCAN_IN), .B2(keyinput_38), .C1(
        P3_REG3_REG_10__SCAN_IN), .C2(keyinput_39), .A(n14520), .ZN(n14521) );
  OAI21_X1 U16053 ( .B1(n14523), .B2(n14522), .A(n14521), .ZN(n14528) );
  XOR2_X1 U16054 ( .A(P3_REG3_REG_28__SCAN_IN), .B(keyinput_42), .Z(n14527) );
  AOI22_X1 U16055 ( .A1(P3_REG3_REG_1__SCAN_IN), .A2(keyinput_44), .B1(n14525), 
        .B2(keyinput_43), .ZN(n14524) );
  OAI221_X1 U16056 ( .B1(P3_REG3_REG_1__SCAN_IN), .B2(keyinput_44), .C1(n14525), .C2(keyinput_43), .A(n14524), .ZN(n14526) );
  AOI211_X1 U16057 ( .C1(n14529), .C2(n14528), .A(n14527), .B(n14526), .ZN(
        n14530) );
  OAI22_X1 U16058 ( .A1(n14632), .A2(keyinput_56), .B1(n14535), .B2(
        keyinput_52), .ZN(n14534) );
  AOI221_X1 U16059 ( .B1(n14632), .B2(keyinput_56), .C1(keyinput_52), .C2(
        n14535), .A(n14534), .ZN(n14542) );
  INV_X1 U16060 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n14537) );
  OAI22_X1 U16061 ( .A1(n14537), .A2(keyinput_50), .B1(keyinput_53), .B2(
        P3_REG3_REG_9__SCAN_IN), .ZN(n14536) );
  AOI221_X1 U16062 ( .B1(n14537), .B2(keyinput_50), .C1(P3_REG3_REG_9__SCAN_IN), .C2(keyinput_53), .A(n14536), .ZN(n14541) );
  OAI22_X1 U16063 ( .A1(P3_REG3_REG_24__SCAN_IN), .A2(keyinput_51), .B1(
        keyinput_55), .B2(P3_REG3_REG_20__SCAN_IN), .ZN(n14538) );
  AOI221_X1 U16064 ( .B1(P3_REG3_REG_24__SCAN_IN), .B2(keyinput_51), .C1(
        P3_REG3_REG_20__SCAN_IN), .C2(keyinput_55), .A(n14538), .ZN(n14540) );
  XNOR2_X1 U16065 ( .A(P3_REG3_REG_0__SCAN_IN), .B(keyinput_54), .ZN(n14539)
         );
  NAND4_X1 U16066 ( .A1(n14542), .A2(n14541), .A3(n14540), .A4(n14539), .ZN(
        n14545) );
  OAI22_X1 U16067 ( .A1(P3_REG3_REG_22__SCAN_IN), .A2(keyinput_57), .B1(
        keyinput_58), .B2(P3_REG3_REG_11__SCAN_IN), .ZN(n14543) );
  AOI221_X1 U16068 ( .B1(P3_REG3_REG_22__SCAN_IN), .B2(keyinput_57), .C1(
        P3_REG3_REG_11__SCAN_IN), .C2(keyinput_58), .A(n14543), .ZN(n14544) );
  OAI21_X1 U16069 ( .B1(n14546), .B2(n14545), .A(n14544), .ZN(n14547) );
  OAI221_X1 U16070 ( .B1(P3_REG3_REG_2__SCAN_IN), .B2(n14548), .C1(n16509), 
        .C2(keyinput_59), .A(n14547), .ZN(n14549) );
  NAND4_X1 U16071 ( .A1(n14552), .A2(n14551), .A3(n14550), .A4(n14549), .ZN(
        n14553) );
  NAND4_X1 U16072 ( .A1(n14556), .A2(n14555), .A3(n14554), .A4(n14553), .ZN(
        n14559) );
  OAI22_X1 U16073 ( .A1(P3_DATAO_REG_22__SCAN_IN), .A2(keyinput_74), .B1(
        keyinput_73), .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n14557) );
  AOI221_X1 U16074 ( .B1(P3_DATAO_REG_22__SCAN_IN), .B2(keyinput_74), .C1(
        P3_DATAO_REG_23__SCAN_IN), .C2(keyinput_73), .A(n14557), .ZN(n14558)
         );
  OAI21_X1 U16075 ( .B1(n14560), .B2(n14559), .A(n14558), .ZN(n14568) );
  AOI22_X1 U16076 ( .A1(n14563), .A2(keyinput_78), .B1(n14562), .B2(
        keyinput_77), .ZN(n14561) );
  OAI221_X1 U16077 ( .B1(n14563), .B2(keyinput_78), .C1(n14562), .C2(
        keyinput_77), .A(n14561), .ZN(n14567) );
  AOI22_X1 U16078 ( .A1(P3_DATAO_REG_17__SCAN_IN), .A2(keyinput_79), .B1(
        n14565), .B2(keyinput_80), .ZN(n14564) );
  OAI221_X1 U16079 ( .B1(P3_DATAO_REG_17__SCAN_IN), .B2(keyinput_79), .C1(
        n14565), .C2(keyinput_80), .A(n14564), .ZN(n14566) );
  AOI22_X1 U16080 ( .A1(P3_DATAO_REG_15__SCAN_IN), .A2(keyinput_81), .B1(
        n14630), .B2(keyinput_83), .ZN(n14570) );
  OAI221_X1 U16081 ( .B1(P3_DATAO_REG_15__SCAN_IN), .B2(keyinput_81), .C1(
        n14630), .C2(keyinput_83), .A(n14570), .ZN(n14571) );
  NAND4_X1 U16082 ( .A1(n14576), .A2(n14575), .A3(n14574), .A4(n14573), .ZN(
        n14581) );
  OAI22_X1 U16083 ( .A1(n14578), .A2(keyinput_91), .B1(P3_DATAO_REG_6__SCAN_IN), .B2(keyinput_90), .ZN(n14577) );
  AOI221_X1 U16084 ( .B1(n14578), .B2(keyinput_91), .C1(keyinput_90), .C2(
        P3_DATAO_REG_6__SCAN_IN), .A(n14577), .ZN(n14580) );
  NOR2_X1 U16085 ( .A1(P3_DATAO_REG_4__SCAN_IN), .A2(keyinput_92), .ZN(n14579)
         );
  AOI22_X1 U16086 ( .A1(P3_DATAO_REG_2__SCAN_IN), .A2(keyinput_94), .B1(n14777), .B2(keyinput_93), .ZN(n14582) );
  OAI221_X1 U16087 ( .B1(P3_DATAO_REG_2__SCAN_IN), .B2(keyinput_94), .C1(
        n14777), .C2(keyinput_93), .A(n14582), .ZN(n14588) );
  OAI22_X1 U16088 ( .A1(n14584), .A2(keyinput_96), .B1(n16274), .B2(
        keyinput_97), .ZN(n14583) );
  AOI221_X1 U16089 ( .B1(n14584), .B2(keyinput_96), .C1(keyinput_97), .C2(
        n16274), .A(n14583), .ZN(n14587) );
  OAI22_X1 U16090 ( .A1(n16272), .A2(keyinput_98), .B1(n14780), .B2(
        keyinput_95), .ZN(n14585) );
  AOI221_X1 U16091 ( .B1(n16272), .B2(keyinput_98), .C1(keyinput_95), .C2(
        n14780), .A(n14585), .ZN(n14586) );
  OAI211_X1 U16092 ( .C1(n14589), .C2(n14588), .A(n14587), .B(n14586), .ZN(
        n14592) );
  AOI22_X1 U16093 ( .A1(P3_ADDR_REG_4__SCAN_IN), .A2(keyinput_101), .B1(n16306), .B2(keyinput_102), .ZN(n14590) );
  OAI221_X1 U16094 ( .B1(P3_ADDR_REG_4__SCAN_IN), .B2(keyinput_101), .C1(
        n16306), .C2(keyinput_102), .A(n14590), .ZN(n14591) );
  AOI21_X1 U16095 ( .B1(n14593), .B2(n14592), .A(n14591), .ZN(n14594) );
  XOR2_X1 U16096 ( .A(keyinput_108), .B(n8829), .Z(n14600) );
  XNOR2_X1 U16097 ( .A(P1_IR_REG_0__SCAN_IN), .B(keyinput_107), .ZN(n14599) );
  NAND2_X1 U16098 ( .A1(n14600), .A2(n14599), .ZN(n14601) );
  OAI22_X1 U16099 ( .A1(n14602), .A2(n14601), .B1(keyinput_109), .B2(n9543), 
        .ZN(n14603) );
  AOI21_X1 U16100 ( .B1(keyinput_109), .B2(n9543), .A(n14603), .ZN(n14604) );
  AOI221_X1 U16101 ( .B1(P1_IR_REG_3__SCAN_IN), .B2(n14605), .C1(n9864), .C2(
        keyinput_110), .A(n14604), .ZN(n14608) );
  INV_X1 U16102 ( .A(keyinput_111), .ZN(n14606) );
  MUX2_X1 U16103 ( .A(keyinput_111), .B(n14606), .S(P1_IR_REG_4__SCAN_IN), .Z(
        n14607) );
  AOI22_X1 U16104 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(keyinput_113), .B1(n9899), 
        .B2(keyinput_112), .ZN(n14609) );
  OAI221_X1 U16105 ( .B1(P1_IR_REG_6__SCAN_IN), .B2(keyinput_113), .C1(n9899), 
        .C2(keyinput_112), .A(n14609), .ZN(n14613) );
  XNOR2_X1 U16106 ( .A(P1_IR_REG_8__SCAN_IN), .B(keyinput_115), .ZN(n14612) );
  OAI22_X1 U16107 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(keyinput_114), .B1(
        keyinput_116), .B2(P1_IR_REG_9__SCAN_IN), .ZN(n14610) );
  AOI221_X1 U16108 ( .B1(P1_IR_REG_7__SCAN_IN), .B2(keyinput_114), .C1(
        P1_IR_REG_9__SCAN_IN), .C2(keyinput_116), .A(n14610), .ZN(n14611) );
  AOI22_X1 U16109 ( .A1(n10640), .A2(keyinput_122), .B1(keyinput_121), .B2(
        n14617), .ZN(n14616) );
  OAI221_X1 U16110 ( .B1(n10640), .B2(keyinput_122), .C1(n14617), .C2(
        keyinput_121), .A(n14616), .ZN(n14618) );
  XOR2_X1 U16111 ( .A(P1_IR_REG_16__SCAN_IN), .B(keyinput_123), .Z(n14622) );
  XNOR2_X1 U16112 ( .A(P1_IR_REG_18__SCAN_IN), .B(keyinput_125), .ZN(n14621)
         );
  XNOR2_X1 U16113 ( .A(P1_IR_REG_17__SCAN_IN), .B(keyinput_124), .ZN(n14620)
         );
  NOR4_X1 U16114 ( .A1(n14623), .A2(n14622), .A3(n14621), .A4(n14620), .ZN(
        n14830) );
  XOR2_X1 U16115 ( .A(P1_IR_REG_19__SCAN_IN), .B(keyinput_126), .Z(n14829) );
  OAI22_X1 U16116 ( .A1(n10452), .A2(keyinput_248), .B1(n10216), .B2(
        keyinput_247), .ZN(n14624) );
  AOI221_X1 U16117 ( .B1(n10452), .B2(keyinput_248), .C1(keyinput_247), .C2(
        n10216), .A(n14624), .ZN(n14816) );
  INV_X1 U16118 ( .A(keyinput_246), .ZN(n14812) );
  INV_X1 U16119 ( .A(keyinput_245), .ZN(n14810) );
  INV_X1 U16120 ( .A(keyinput_238), .ZN(n14799) );
  AOI22_X1 U16121 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(keyinput_235), .B1(n8829), 
        .B2(keyinput_236), .ZN(n14625) );
  OAI221_X1 U16122 ( .B1(P1_IR_REG_0__SCAN_IN), .B2(keyinput_235), .C1(n8829), 
        .C2(keyinput_236), .A(n14625), .ZN(n14796) );
  INV_X1 U16123 ( .A(keyinput_234), .ZN(n14794) );
  INV_X1 U16124 ( .A(keyinput_233), .ZN(n14793) );
  INV_X1 U16125 ( .A(keyinput_232), .ZN(n14792) );
  INV_X1 U16126 ( .A(keyinput_231), .ZN(n14791) );
  OAI22_X1 U16127 ( .A1(P3_ADDR_REG_2__SCAN_IN), .A2(keyinput_227), .B1(
        P3_ADDR_REG_3__SCAN_IN), .B2(keyinput_228), .ZN(n14626) );
  AOI221_X1 U16128 ( .B1(P3_ADDR_REG_2__SCAN_IN), .B2(keyinput_227), .C1(
        keyinput_228), .C2(P3_ADDR_REG_3__SCAN_IN), .A(n14626), .ZN(n14789) );
  AOI22_X1 U16129 ( .A1(P3_DATAO_REG_5__SCAN_IN), .A2(keyinput_219), .B1(
        P3_DATAO_REG_6__SCAN_IN), .B2(keyinput_218), .ZN(n14627) );
  OAI221_X1 U16130 ( .B1(P3_DATAO_REG_5__SCAN_IN), .B2(keyinput_219), .C1(
        P3_DATAO_REG_6__SCAN_IN), .C2(keyinput_218), .A(n14627), .ZN(n14773)
         );
  INV_X1 U16131 ( .A(keyinput_212), .ZN(n14764) );
  OAI22_X1 U16132 ( .A1(n14630), .A2(keyinput_211), .B1(n14629), .B2(
        keyinput_209), .ZN(n14628) );
  AOI221_X1 U16133 ( .B1(n14630), .B2(keyinput_211), .C1(keyinput_209), .C2(
        n14629), .A(n14628), .ZN(n14761) );
  INV_X1 U16134 ( .A(keyinput_187), .ZN(n14723) );
  XOR2_X1 U16135 ( .A(P3_REG3_REG_0__SCAN_IN), .B(keyinput_182), .Z(n14639) );
  AOI22_X1 U16136 ( .A1(n8863), .A2(keyinput_181), .B1(n14632), .B2(
        keyinput_184), .ZN(n14631) );
  OAI221_X1 U16137 ( .B1(n8863), .B2(keyinput_181), .C1(n14632), .C2(
        keyinput_184), .A(n14631), .ZN(n14638) );
  AOI22_X1 U16138 ( .A1(P3_REG3_REG_17__SCAN_IN), .A2(keyinput_178), .B1(
        n14634), .B2(keyinput_179), .ZN(n14633) );
  OAI221_X1 U16139 ( .B1(P3_REG3_REG_17__SCAN_IN), .B2(keyinput_178), .C1(
        n14634), .C2(keyinput_179), .A(n14633), .ZN(n14637) );
  AOI22_X1 U16140 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(keyinput_180), .B1(
        P3_REG3_REG_20__SCAN_IN), .B2(keyinput_183), .ZN(n14635) );
  OAI221_X1 U16141 ( .B1(P3_REG3_REG_4__SCAN_IN), .B2(keyinput_180), .C1(
        P3_REG3_REG_20__SCAN_IN), .C2(keyinput_183), .A(n14635), .ZN(n14636)
         );
  NOR4_X1 U16142 ( .A1(n14639), .A2(n14638), .A3(n14637), .A4(n14636), .ZN(
        n14722) );
  INV_X1 U16143 ( .A(keyinput_177), .ZN(n14717) );
  INV_X1 U16144 ( .A(keyinput_176), .ZN(n14714) );
  OAI22_X1 U16145 ( .A1(n14641), .A2(keyinput_173), .B1(
        P3_REG3_REG_12__SCAN_IN), .B2(keyinput_174), .ZN(n14640) );
  AOI221_X1 U16146 ( .B1(n14641), .B2(keyinput_173), .C1(keyinput_174), .C2(
        P3_REG3_REG_12__SCAN_IN), .A(n14640), .ZN(n14710) );
  OAI22_X1 U16147 ( .A1(n14644), .A2(keyinput_164), .B1(n14643), .B2(
        keyinput_165), .ZN(n14642) );
  AOI221_X1 U16148 ( .B1(n14644), .B2(keyinput_164), .C1(keyinput_165), .C2(
        n14643), .A(n14642), .ZN(n14701) );
  INV_X1 U16149 ( .A(keyinput_163), .ZN(n14696) );
  OAI22_X1 U16150 ( .A1(SI_0_), .A2(keyinput_160), .B1(P3_RD_REG_SCAN_IN), 
        .B2(keyinput_161), .ZN(n14645) );
  AOI221_X1 U16151 ( .B1(SI_0_), .B2(keyinput_160), .C1(keyinput_161), .C2(
        P3_RD_REG_SCAN_IN), .A(n14645), .ZN(n14695) );
  INV_X1 U16152 ( .A(keyinput_149), .ZN(n14678) );
  INV_X1 U16153 ( .A(keyinput_148), .ZN(n14677) );
  OAI22_X1 U16154 ( .A1(n14647), .A2(keyinput_146), .B1(keyinput_145), .B2(
        SI_15_), .ZN(n14646) );
  AOI221_X1 U16155 ( .B1(n14647), .B2(keyinput_146), .C1(SI_15_), .C2(
        keyinput_145), .A(n14646), .ZN(n14672) );
  INV_X1 U16156 ( .A(keyinput_140), .ZN(n14663) );
  INV_X1 U16157 ( .A(keyinput_139), .ZN(n14661) );
  OAI221_X1 U16158 ( .B1(SI_30_), .B2(keyinput_130), .C1(n14914), .C2(
        keyinput_131), .A(n14648), .ZN(n14651) );
  OAI22_X1 U16159 ( .A1(SI_31_), .A2(keyinput_129), .B1(P3_WR_REG_SCAN_IN), 
        .B2(keyinput_128), .ZN(n14649) );
  AOI221_X1 U16160 ( .B1(SI_31_), .B2(keyinput_129), .C1(keyinput_128), .C2(
        P3_WR_REG_SCAN_IN), .A(n14649), .ZN(n14650) );
  OAI22_X1 U16161 ( .A1(n14651), .A2(n14650), .B1(SI_26_), .B2(keyinput_134), 
        .ZN(n14652) );
  OAI22_X1 U16162 ( .A1(SI_28_), .A2(keyinput_132), .B1(keyinput_133), .B2(
        SI_27_), .ZN(n14653) );
  AOI221_X1 U16163 ( .B1(SI_28_), .B2(keyinput_132), .C1(SI_27_), .C2(
        keyinput_133), .A(n14653), .ZN(n14660) );
  INV_X1 U16164 ( .A(SI_22_), .ZN(n14655) );
  AOI22_X1 U16165 ( .A1(n14656), .A2(keyinput_135), .B1(keyinput_138), .B2(
        n14655), .ZN(n14654) );
  OAI221_X1 U16166 ( .B1(n14656), .B2(keyinput_135), .C1(n14655), .C2(
        keyinput_138), .A(n14654), .ZN(n14659) );
  AOI22_X1 U16167 ( .A1(SI_23_), .A2(keyinput_137), .B1(SI_24_), .B2(
        keyinput_136), .ZN(n14657) );
  OAI221_X1 U16168 ( .B1(SI_23_), .B2(keyinput_137), .C1(SI_24_), .C2(
        keyinput_136), .A(n14657), .ZN(n14658) );
  AOI22_X1 U16169 ( .A1(SI_18_), .A2(keyinput_142), .B1(n14666), .B2(
        keyinput_141), .ZN(n14665) );
  OAI221_X1 U16170 ( .B1(SI_18_), .B2(keyinput_142), .C1(n14666), .C2(
        keyinput_141), .A(n14665), .ZN(n14669) );
  OAI22_X1 U16171 ( .A1(SI_17_), .A2(keyinput_143), .B1(keyinput_144), .B2(
        SI_16_), .ZN(n14667) );
  AOI221_X1 U16172 ( .B1(SI_17_), .B2(keyinput_143), .C1(SI_16_), .C2(
        keyinput_144), .A(n14667), .ZN(n14668) );
  OAI21_X1 U16173 ( .B1(n14670), .B2(n14669), .A(n14668), .ZN(n14671) );
  AOI22_X1 U16174 ( .A1(keyinput_147), .A2(n14674), .B1(n14672), .B2(n14671), 
        .ZN(n14673) );
  OAI21_X1 U16175 ( .B1(n14674), .B2(keyinput_147), .A(n14673), .ZN(n14675) );
  XNOR2_X1 U16176 ( .A(keyinput_150), .B(n14680), .ZN(n14686) );
  AOI22_X1 U16177 ( .A1(SI_8_), .A2(keyinput_152), .B1(SI_9_), .B2(
        keyinput_151), .ZN(n14681) );
  OAI221_X1 U16178 ( .B1(SI_8_), .B2(keyinput_152), .C1(SI_9_), .C2(
        keyinput_151), .A(n14681), .ZN(n14685) );
  XNOR2_X1 U16179 ( .A(SI_6_), .B(keyinput_154), .ZN(n14683) );
  XNOR2_X1 U16180 ( .A(SI_7_), .B(keyinput_153), .ZN(n14682) );
  NAND2_X1 U16181 ( .A1(n14683), .A2(n14682), .ZN(n14684) );
  AOI22_X1 U16182 ( .A1(SI_4_), .A2(keyinput_156), .B1(SI_5_), .B2(
        keyinput_155), .ZN(n14687) );
  OAI221_X1 U16183 ( .B1(SI_4_), .B2(keyinput_156), .C1(SI_5_), .C2(
        keyinput_155), .A(n14687), .ZN(n14688) );
  XNOR2_X1 U16184 ( .A(SI_1_), .B(keyinput_159), .ZN(n14692) );
  INV_X1 U16185 ( .A(keyinput_158), .ZN(n14689) );
  XNOR2_X1 U16186 ( .A(n14689), .B(SI_2_), .ZN(n14691) );
  XNOR2_X1 U16187 ( .A(SI_3_), .B(keyinput_157), .ZN(n14690) );
  NAND4_X1 U16188 ( .A1(n14693), .A2(n14692), .A3(n14691), .A4(n14690), .ZN(
        n14694) );
  INV_X1 U16189 ( .A(P3_REG3_REG_23__SCAN_IN), .ZN(n14698) );
  AOI22_X1 U16190 ( .A1(n14699), .A2(keyinput_167), .B1(n14698), .B2(
        keyinput_166), .ZN(n14697) );
  OAI221_X1 U16191 ( .B1(n14699), .B2(keyinput_167), .C1(n14698), .C2(
        keyinput_166), .A(n14697), .ZN(n14700) );
  AOI22_X1 U16192 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(keyinput_168), .B1(n14703), .B2(keyinput_169), .ZN(n14702) );
  OAI221_X1 U16193 ( .B1(P3_REG3_REG_3__SCAN_IN), .B2(keyinput_168), .C1(
        n14703), .C2(keyinput_169), .A(n14702), .ZN(n14707) );
  OAI22_X1 U16194 ( .A1(P3_REG3_REG_28__SCAN_IN), .A2(keyinput_170), .B1(
        P3_REG3_REG_1__SCAN_IN), .B2(keyinput_172), .ZN(n14704) );
  AOI221_X1 U16195 ( .B1(P3_REG3_REG_28__SCAN_IN), .B2(keyinput_170), .C1(
        keyinput_172), .C2(P3_REG3_REG_1__SCAN_IN), .A(n14704), .ZN(n14706) );
  XNOR2_X1 U16196 ( .A(P3_REG3_REG_8__SCAN_IN), .B(keyinput_171), .ZN(n14705)
         );
  OAI211_X1 U16197 ( .C1(n14708), .C2(n14707), .A(n14706), .B(n14705), .ZN(
        n14709) );
  AOI22_X1 U16198 ( .A1(keyinput_175), .A2(n14712), .B1(n14710), .B2(n14709), 
        .ZN(n14711) );
  OAI21_X1 U16199 ( .B1(n14712), .B2(keyinput_175), .A(n14711), .ZN(n14713) );
  AOI22_X1 U16200 ( .A1(n14720), .A2(keyinput_185), .B1(keyinput_186), .B2(
        n14719), .ZN(n14718) );
  OAI221_X1 U16201 ( .B1(n14720), .B2(keyinput_185), .C1(n14719), .C2(
        keyinput_186), .A(n14718), .ZN(n14721) );
  AOI22_X1 U16202 ( .A1(n14726), .A2(keyinput_197), .B1(keyinput_194), .B2(
        n14725), .ZN(n14724) );
  OAI221_X1 U16203 ( .B1(n14726), .B2(keyinput_197), .C1(n14725), .C2(
        keyinput_194), .A(n14724), .ZN(n14736) );
  AOI22_X1 U16204 ( .A1(n14729), .A2(keyinput_195), .B1(keyinput_193), .B2(
        n14728), .ZN(n14727) );
  OAI221_X1 U16205 ( .B1(n14729), .B2(keyinput_195), .C1(n14728), .C2(
        keyinput_193), .A(n14727), .ZN(n14735) );
  AOI22_X1 U16206 ( .A1(P3_DATAO_REG_24__SCAN_IN), .A2(keyinput_200), .B1(
        P3_DATAO_REG_26__SCAN_IN), .B2(keyinput_198), .ZN(n14730) );
  OAI221_X1 U16207 ( .B1(P3_DATAO_REG_24__SCAN_IN), .B2(keyinput_200), .C1(
        P3_DATAO_REG_26__SCAN_IN), .C2(keyinput_198), .A(n14730), .ZN(n14734)
         );
  AOI22_X1 U16208 ( .A1(keyinput_199), .A2(P3_DATAO_REG_25__SCAN_IN), .B1(
        n14732), .B2(keyinput_196), .ZN(n14731) );
  OAI221_X1 U16209 ( .B1(keyinput_199), .B2(P3_DATAO_REG_25__SCAN_IN), .C1(
        n14732), .C2(keyinput_196), .A(n14731), .ZN(n14733) );
  NOR4_X1 U16210 ( .A1(n14736), .A2(n14735), .A3(n14734), .A4(n14733), .ZN(
        n14748) );
  AOI22_X1 U16211 ( .A1(n14739), .A2(keyinput_190), .B1(keyinput_188), .B2(
        n14738), .ZN(n14737) );
  OAI221_X1 U16212 ( .B1(n14739), .B2(keyinput_190), .C1(n14738), .C2(
        keyinput_188), .A(n14737), .ZN(n14743) );
  AOI22_X1 U16213 ( .A1(P3_B_REG_SCAN_IN), .A2(keyinput_192), .B1(n14741), 
        .B2(keyinput_189), .ZN(n14740) );
  OAI221_X1 U16214 ( .B1(P3_B_REG_SCAN_IN), .B2(keyinput_192), .C1(n14741), 
        .C2(keyinput_189), .A(n14740), .ZN(n14742) );
  AOI211_X1 U16215 ( .C1(keyinput_191), .C2(P3_REG3_REG_15__SCAN_IN), .A(
        n14743), .B(n14742), .ZN(n14744) );
  OAI21_X1 U16216 ( .B1(keyinput_191), .B2(P3_REG3_REG_15__SCAN_IN), .A(n14744), .ZN(n14747) );
  AOI22_X1 U16217 ( .A1(P3_DATAO_REG_23__SCAN_IN), .A2(keyinput_201), .B1(
        P3_DATAO_REG_22__SCAN_IN), .B2(keyinput_202), .ZN(n14745) );
  OAI221_X1 U16218 ( .B1(P3_DATAO_REG_23__SCAN_IN), .B2(keyinput_201), .C1(
        P3_DATAO_REG_22__SCAN_IN), .C2(keyinput_202), .A(n14745), .ZN(n14746)
         );
  AOI221_X1 U16219 ( .B1(n14749), .B2(n14748), .C1(n14747), .C2(n14748), .A(
        n14746), .ZN(n14759) );
  AOI22_X1 U16220 ( .A1(n14752), .A2(keyinput_203), .B1(keyinput_204), .B2(
        n14751), .ZN(n14750) );
  OAI221_X1 U16221 ( .B1(n14752), .B2(keyinput_203), .C1(n14751), .C2(
        keyinput_204), .A(n14750), .ZN(n14758) );
  OAI22_X1 U16222 ( .A1(n14754), .A2(keyinput_207), .B1(
        P3_DATAO_REG_18__SCAN_IN), .B2(keyinput_206), .ZN(n14753) );
  AOI221_X1 U16223 ( .B1(n14754), .B2(keyinput_207), .C1(keyinput_206), .C2(
        P3_DATAO_REG_18__SCAN_IN), .A(n14753), .ZN(n14757) );
  OAI22_X1 U16224 ( .A1(P3_DATAO_REG_19__SCAN_IN), .A2(keyinput_205), .B1(
        P3_DATAO_REG_16__SCAN_IN), .B2(keyinput_208), .ZN(n14755) );
  AOI221_X1 U16225 ( .B1(P3_DATAO_REG_19__SCAN_IN), .B2(keyinput_205), .C1(
        keyinput_208), .C2(P3_DATAO_REG_16__SCAN_IN), .A(n14755), .ZN(n14756)
         );
  OAI211_X1 U16226 ( .C1(n14759), .C2(n14758), .A(n14757), .B(n14756), .ZN(
        n14760) );
  XNOR2_X1 U16227 ( .A(P3_DATAO_REG_10__SCAN_IN), .B(keyinput_214), .ZN(n14771) );
  AOI22_X1 U16228 ( .A1(keyinput_215), .A2(P3_DATAO_REG_9__SCAN_IN), .B1(
        n14766), .B2(keyinput_217), .ZN(n14765) );
  OAI221_X1 U16229 ( .B1(keyinput_215), .B2(P3_DATAO_REG_9__SCAN_IN), .C1(
        n14766), .C2(keyinput_217), .A(n14765), .ZN(n14770) );
  AOI22_X1 U16230 ( .A1(P3_DATAO_REG_8__SCAN_IN), .A2(keyinput_216), .B1(
        n14768), .B2(keyinput_213), .ZN(n14767) );
  OAI221_X1 U16231 ( .B1(P3_DATAO_REG_8__SCAN_IN), .B2(keyinput_216), .C1(
        n14768), .C2(keyinput_213), .A(n14767), .ZN(n14769) );
  OAI22_X1 U16232 ( .A1(keyinput_220), .A2(n14775), .B1(n14773), .B2(n14772), 
        .ZN(n14774) );
  AOI21_X1 U16233 ( .B1(keyinput_220), .B2(n14775), .A(n14774), .ZN(n14785) );
  AOI22_X1 U16234 ( .A1(n14778), .A2(keyinput_222), .B1(keyinput_221), .B2(
        n14777), .ZN(n14776) );
  OAI221_X1 U16235 ( .B1(n14778), .B2(keyinput_222), .C1(n14777), .C2(
        keyinput_221), .A(n14776), .ZN(n14784) );
  OAI22_X1 U16236 ( .A1(n16274), .A2(keyinput_225), .B1(n14780), .B2(
        keyinput_223), .ZN(n14779) );
  AOI221_X1 U16237 ( .B1(n16274), .B2(keyinput_225), .C1(keyinput_223), .C2(
        n14780), .A(n14779), .ZN(n14783) );
  OAI22_X1 U16238 ( .A1(P3_ADDR_REG_1__SCAN_IN), .A2(keyinput_226), .B1(
        P3_DATAO_REG_0__SCAN_IN), .B2(keyinput_224), .ZN(n14781) );
  AOI221_X1 U16239 ( .B1(P3_ADDR_REG_1__SCAN_IN), .B2(keyinput_226), .C1(
        keyinput_224), .C2(P3_DATAO_REG_0__SCAN_IN), .A(n14781), .ZN(n14782)
         );
  OAI211_X1 U16240 ( .C1(n14785), .C2(n14784), .A(n14783), .B(n14782), .ZN(
        n14788) );
  AOI22_X1 U16241 ( .A1(P3_ADDR_REG_5__SCAN_IN), .A2(keyinput_230), .B1(
        P3_ADDR_REG_4__SCAN_IN), .B2(keyinput_229), .ZN(n14786) );
  OAI221_X1 U16242 ( .B1(P3_ADDR_REG_5__SCAN_IN), .B2(keyinput_230), .C1(
        P3_ADDR_REG_4__SCAN_IN), .C2(keyinput_229), .A(n14786), .ZN(n14787) );
  AOI21_X1 U16243 ( .B1(n14789), .B2(n14788), .A(n14787), .ZN(n14790) );
  OAI22_X1 U16244 ( .A1(keyinput_237), .A2(n9543), .B1(n14796), .B2(n14795), 
        .ZN(n14797) );
  AOI21_X1 U16245 ( .B1(keyinput_237), .B2(n9543), .A(n14797), .ZN(n14798) );
  AOI221_X1 U16246 ( .B1(P1_IR_REG_3__SCAN_IN), .B2(n14799), .C1(n9864), .C2(
        keyinput_238), .A(n14798), .ZN(n14804) );
  INV_X1 U16247 ( .A(keyinput_239), .ZN(n14800) );
  MUX2_X1 U16248 ( .A(n14800), .B(keyinput_239), .S(P1_IR_REG_4__SCAN_IN), .Z(
        n14803) );
  XOR2_X1 U16249 ( .A(n9899), .B(keyinput_240), .Z(n14802) );
  XNOR2_X1 U16250 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput_241), .ZN(n14801) );
  OAI211_X1 U16251 ( .C1(n14804), .C2(n14803), .A(n14802), .B(n14801), .ZN(
        n14808) );
  XNOR2_X1 U16252 ( .A(P1_IR_REG_9__SCAN_IN), .B(keyinput_244), .ZN(n14807) );
  OAI22_X1 U16253 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(keyinput_242), .B1(
        keyinput_243), .B2(P1_IR_REG_8__SCAN_IN), .ZN(n14805) );
  AOI221_X1 U16254 ( .B1(P1_IR_REG_7__SCAN_IN), .B2(keyinput_242), .C1(
        P1_IR_REG_8__SCAN_IN), .C2(keyinput_243), .A(n14805), .ZN(n14806) );
  NAND3_X1 U16255 ( .A1(n14808), .A2(n14807), .A3(n14806), .ZN(n14809) );
  OAI221_X1 U16256 ( .B1(P1_IR_REG_10__SCAN_IN), .B2(keyinput_245), .C1(n10007), .C2(n14810), .A(n14809), .ZN(n14811) );
  OAI221_X1 U16257 ( .B1(P1_IR_REG_11__SCAN_IN), .B2(keyinput_246), .C1(n10144), .C2(n14812), .A(n14811), .ZN(n14815) );
  AOI22_X1 U16258 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(keyinput_249), .B1(n10640), 
        .B2(keyinput_250), .ZN(n14813) );
  OAI221_X1 U16259 ( .B1(P1_IR_REG_14__SCAN_IN), .B2(keyinput_249), .C1(n10640), .C2(keyinput_250), .A(n14813), .ZN(n14814) );
  AOI21_X1 U16260 ( .B1(n14816), .B2(n14815), .A(n14814), .ZN(n14823) );
  XOR2_X1 U16261 ( .A(P1_IR_REG_17__SCAN_IN), .B(keyinput_252), .Z(n14819) );
  XOR2_X1 U16262 ( .A(P1_IR_REG_16__SCAN_IN), .B(keyinput_251), .Z(n14818) );
  XNOR2_X1 U16263 ( .A(P1_IR_REG_18__SCAN_IN), .B(keyinput_253), .ZN(n14817)
         );
  NAND3_X1 U16264 ( .A1(n14819), .A2(n14818), .A3(n14817), .ZN(n14822) );
  INV_X1 U16265 ( .A(keyinput_254), .ZN(n14820) );
  MUX2_X1 U16266 ( .A(keyinput_254), .B(n14820), .S(P1_IR_REG_19__SCAN_IN), 
        .Z(n14821) );
  OAI21_X1 U16267 ( .B1(n14823), .B2(n14822), .A(n14821), .ZN(n14827) );
  INV_X1 U16268 ( .A(keyinput_255), .ZN(n14824) );
  MUX2_X1 U16269 ( .A(keyinput_255), .B(n14824), .S(P1_IR_REG_20__SCAN_IN), 
        .Z(n14826) );
  XNOR2_X1 U16270 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput_127), .ZN(n14825)
         );
  AOI21_X1 U16271 ( .B1(n14827), .B2(n14826), .A(n14825), .ZN(n14828) );
  OAI22_X1 U16272 ( .A1(n14832), .A2(n16615), .B1(n14831), .B2(n16711), .ZN(
        n14833) );
  NOR2_X1 U16273 ( .A1(n14834), .A2(n14833), .ZN(n14898) );
  NOR2_X1 U16274 ( .A1(n16718), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n14835) );
  AOI21_X1 U16275 ( .B1(n14898), .B2(n16718), .A(n14835), .ZN(n14836) );
  XNOR2_X1 U16276 ( .A(n14837), .B(n14836), .ZN(P3_U3471) );
  NOR2_X1 U16277 ( .A1(n16719), .A2(n14838), .ZN(n14841) );
  AOI21_X1 U16278 ( .B1(n16719), .B2(P3_REG0_REG_31__SCAN_IN), .A(n14841), 
        .ZN(n14839) );
  OAI21_X1 U16279 ( .B1(n14840), .B2(n14896), .A(n14839), .ZN(P3_U3458) );
  AOI21_X1 U16280 ( .B1(n16719), .B2(P3_REG0_REG_30__SCAN_IN), .A(n14841), 
        .ZN(n14842) );
  OAI21_X1 U16281 ( .B1(n14843), .B2(n14896), .A(n14842), .ZN(P3_U3457) );
  MUX2_X1 U16282 ( .A(P3_REG0_REG_28__SCAN_IN), .B(n14844), .S(n14891), .Z(
        P3_U3455) );
  NOR2_X1 U16283 ( .A1(n14845), .A2(n16615), .ZN(n14846) );
  OAI21_X1 U16284 ( .B1(n14847), .B2(n14846), .A(n14891), .ZN(n14849) );
  NAND2_X1 U16285 ( .A1(n16719), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n14848) );
  OAI211_X1 U16286 ( .C1(n14850), .C2(n14896), .A(n14849), .B(n14848), .ZN(
        P3_U3454) );
  MUX2_X1 U16287 ( .A(n14852), .B(n14851), .S(n14891), .Z(n14853) );
  OAI21_X1 U16288 ( .B1(n14854), .B2(n14896), .A(n14853), .ZN(P3_U3453) );
  MUX2_X1 U16289 ( .A(n14856), .B(n14855), .S(n14891), .Z(n14857) );
  OAI21_X1 U16290 ( .B1(n8351), .B2(n14896), .A(n14857), .ZN(P3_U3452) );
  MUX2_X1 U16291 ( .A(n14859), .B(n14858), .S(n14891), .Z(n14860) );
  OAI21_X1 U16292 ( .B1(n14861), .B2(n14896), .A(n14860), .ZN(P3_U3451) );
  MUX2_X1 U16293 ( .A(n14863), .B(n14862), .S(n14891), .Z(n14864) );
  OAI21_X1 U16294 ( .B1(n14865), .B2(n14896), .A(n14864), .ZN(P3_U3450) );
  MUX2_X1 U16295 ( .A(n14867), .B(n14866), .S(n14891), .Z(n14868) );
  OAI21_X1 U16296 ( .B1(n14869), .B2(n14896), .A(n14868), .ZN(P3_U3449) );
  MUX2_X1 U16297 ( .A(n14871), .B(n14870), .S(n14891), .Z(n14872) );
  OAI21_X1 U16298 ( .B1(n14873), .B2(n14896), .A(n14872), .ZN(P3_U3448) );
  MUX2_X1 U16299 ( .A(n14875), .B(n14874), .S(n14891), .Z(n14876) );
  OAI21_X1 U16300 ( .B1(n14877), .B2(n14896), .A(n14876), .ZN(P3_U3447) );
  MUX2_X1 U16301 ( .A(n14879), .B(n14878), .S(n14891), .Z(n14880) );
  OAI21_X1 U16302 ( .B1(n14881), .B2(n14896), .A(n14880), .ZN(P3_U3446) );
  MUX2_X1 U16303 ( .A(n14882), .B(P3_REG0_REG_18__SCAN_IN), .S(n16719), .Z(
        P3_U3444) );
  MUX2_X1 U16304 ( .A(n14884), .B(n14883), .S(n14891), .Z(n14885) );
  OAI21_X1 U16305 ( .B1(n14896), .B2(n14886), .A(n14885), .ZN(P3_U3441) );
  MUX2_X1 U16306 ( .A(P3_REG0_REG_16__SCAN_IN), .B(n14887), .S(n14891), .Z(
        P3_U3438) );
  MUX2_X1 U16307 ( .A(n14889), .B(n14888), .S(n14891), .Z(n14890) );
  INV_X1 U16308 ( .A(n14890), .ZN(P3_U3435) );
  MUX2_X1 U16309 ( .A(n14893), .B(n14892), .S(n14891), .Z(n14894) );
  OAI21_X1 U16310 ( .B1(n14896), .B2(n14895), .A(n14894), .ZN(P3_U3432) );
  NAND2_X1 U16311 ( .A1(n16719), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n14897) );
  OAI21_X1 U16312 ( .B1(n14898), .B2(n16719), .A(n14897), .ZN(P3_U3426) );
  MUX2_X1 U16313 ( .A(P3_D_REG_0__SCAN_IN), .B(n14900), .S(n14899), .Z(
        P3_U3376) );
  NAND2_X1 U16314 ( .A1(n14902), .A2(n14901), .ZN(n14907) );
  INV_X1 U16315 ( .A(n14903), .ZN(n14905) );
  INV_X1 U16316 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n14904) );
  NAND4_X1 U16317 ( .A1(n14905), .A2(P3_IR_REG_31__SCAN_IN), .A3(
        P3_STATE_REG_SCAN_IN), .A4(n14904), .ZN(n14906) );
  OAI211_X1 U16318 ( .C1(n14920), .C2(n14908), .A(n14907), .B(n14906), .ZN(
        P3_U3264) );
  OAI222_X1 U16319 ( .A1(n14911), .A2(P3_U3151), .B1(n14920), .B2(n14910), 
        .C1(n14918), .C2(n14909), .ZN(P3_U3265) );
  INV_X1 U16320 ( .A(n14912), .ZN(n14913) );
  OAI222_X1 U16321 ( .A1(n14915), .A2(P3_U3151), .B1(n14920), .B2(n14914), 
        .C1(n14918), .C2(n14913), .ZN(P3_U3266) );
  INV_X1 U16322 ( .A(n14916), .ZN(n14917) );
  OAI222_X1 U16323 ( .A1(n14921), .A2(P3_U3151), .B1(n14920), .B2(n14919), 
        .C1(n14918), .C2(n14917), .ZN(P3_U3267) );
  XNOR2_X1 U16324 ( .A(n15256), .B(n14959), .ZN(n14926) );
  XNOR2_X1 U16325 ( .A(n14925), .B(n14926), .ZN(n14950) );
  NAND2_X1 U16326 ( .A1(n14950), .A2(n14924), .ZN(n14949) );
  INV_X1 U16327 ( .A(n14925), .ZN(n14927) );
  NAND2_X1 U16328 ( .A1(n14949), .A2(n14928), .ZN(n14987) );
  XNOR2_X1 U16329 ( .A(n15414), .B(n14929), .ZN(n14979) );
  NAND2_X1 U16330 ( .A1(n15132), .A2(n14937), .ZN(n14930) );
  NOR2_X1 U16331 ( .A1(n14979), .A2(n14930), .ZN(n14935) );
  AOI21_X1 U16332 ( .B1(n14979), .B2(n14930), .A(n14935), .ZN(n14988) );
  AND2_X2 U16333 ( .A1(n14987), .A2(n14988), .ZN(n14977) );
  XNOR2_X1 U16334 ( .A(n15408), .B(n14959), .ZN(n14931) );
  AND2_X1 U16335 ( .A1(n15134), .A2(n14937), .ZN(n14932) );
  NAND2_X1 U16336 ( .A1(n14931), .A2(n14932), .ZN(n14938) );
  INV_X1 U16337 ( .A(n14931), .ZN(n15012) );
  INV_X1 U16338 ( .A(n14932), .ZN(n14933) );
  NAND2_X1 U16339 ( .A1(n15012), .A2(n14933), .ZN(n14934) );
  AND2_X1 U16340 ( .A1(n14938), .A2(n14934), .ZN(n14978) );
  XNOR2_X1 U16341 ( .A(n15211), .B(n14936), .ZN(n14941) );
  NAND2_X1 U16342 ( .A1(n15162), .A2(n14937), .ZN(n14939) );
  XNOR2_X1 U16343 ( .A(n14941), .B(n14939), .ZN(n15025) );
  INV_X1 U16344 ( .A(n14939), .ZN(n14940) );
  XNOR2_X1 U16345 ( .A(n15195), .B(n14959), .ZN(n14943) );
  AND2_X1 U16346 ( .A1(n15017), .A2(n14937), .ZN(n14942) );
  NAND2_X1 U16347 ( .A1(n14943), .A2(n14942), .ZN(n14956) );
  OAI21_X1 U16348 ( .B1(n14943), .B2(n14942), .A(n14956), .ZN(n14944) );
  AOI22_X1 U16349 ( .A1(n15137), .A2(n15343), .B1(n15341), .B2(n15162), .ZN(
        n15191) );
  NAND2_X1 U16350 ( .A1(n15195), .A2(n15024), .ZN(n14947) );
  AOI22_X1 U16351 ( .A1(n15199), .A2(n15018), .B1(P2_REG3_REG_27__SCAN_IN), 
        .B2(P2_U3088), .ZN(n14946) );
  OAI211_X1 U16352 ( .C1(n15191), .C2(n15020), .A(n14947), .B(n14946), .ZN(
        n14948) );
  INV_X1 U16353 ( .A(n14949), .ZN(n14955) );
  AOI22_X1 U16354 ( .A1(n14950), .A2(n15014), .B1(n14961), .B2(n15266), .ZN(
        n14954) );
  AOI22_X1 U16355 ( .A1(n15132), .A2(n15343), .B1(n15341), .B2(n15145), .ZN(
        n15252) );
  AOI22_X1 U16356 ( .A1(n15259), .A2(n15018), .B1(P2_REG3_REG_23__SCAN_IN), 
        .B2(P2_U3088), .ZN(n14951) );
  OAI21_X1 U16357 ( .B1(n15252), .B2(n15020), .A(n14951), .ZN(n14952) );
  AOI21_X1 U16358 ( .B1(n15256), .B2(n15024), .A(n14952), .ZN(n14953) );
  OAI21_X1 U16359 ( .B1(n14955), .B2(n14954), .A(n14953), .ZN(P2_U3188) );
  INV_X1 U16360 ( .A(n14956), .ZN(n14957) );
  NAND2_X1 U16361 ( .A1(n15017), .A2(n15341), .ZN(n14963) );
  NAND2_X1 U16362 ( .A1(n15027), .A2(n15343), .ZN(n14962) );
  NAND2_X1 U16363 ( .A1(n14963), .A2(n14962), .ZN(n15181) );
  OAI22_X1 U16364 ( .A1(n15182), .A2(n15003), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14964), .ZN(n14965) );
  AOI21_X1 U16365 ( .B1(n15181), .B2(n14991), .A(n14965), .ZN(n14967) );
  NAND2_X1 U16366 ( .A1(n15184), .A2(n15024), .ZN(n14966) );
  OAI211_X1 U16367 ( .C1(n14970), .C2(n14969), .A(n14968), .B(n15000), .ZN(
        n14976) );
  AOI22_X1 U16368 ( .A1(n15293), .A2(n15018), .B1(P2_REG3_REG_21__SCAN_IN), 
        .B2(P2_U3088), .ZN(n14971) );
  OAI21_X1 U16369 ( .B1(n15286), .B2(n14972), .A(n14971), .ZN(n14973) );
  AOI21_X1 U16370 ( .B1(n14974), .B2(n15320), .A(n14973), .ZN(n14975) );
  OAI211_X1 U16371 ( .C1(n15496), .C2(n14994), .A(n14976), .B(n14975), .ZN(
        P2_U3195) );
  INV_X1 U16372 ( .A(n14977), .ZN(n14986) );
  AOI21_X1 U16373 ( .B1(n14986), .B2(n7925), .A(n15021), .ZN(n14981) );
  INV_X1 U16374 ( .A(n15132), .ZN(n15159) );
  NOR3_X1 U16375 ( .A1(n14979), .A2(n15159), .A3(n15011), .ZN(n14980) );
  OAI21_X1 U16376 ( .B1(n14981), .B2(n14980), .A(n15010), .ZN(n14985) );
  OAI22_X1 U16377 ( .A1(n15136), .A2(n15287), .B1(n15159), .B2(n15289), .ZN(
        n15222) );
  OAI22_X1 U16378 ( .A1(n15230), .A2(n15003), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14982), .ZN(n14983) );
  AOI21_X1 U16379 ( .B1(n15222), .B2(n14991), .A(n14983), .ZN(n14984) );
  OAI211_X1 U16380 ( .C1(n15228), .C2(n14994), .A(n14985), .B(n14984), .ZN(
        P2_U3197) );
  OAI211_X1 U16381 ( .C1(n14988), .C2(n14987), .A(n14986), .B(n15000), .ZN(
        n14993) );
  INV_X1 U16382 ( .A(n15134), .ZN(n15161) );
  OAI22_X1 U16383 ( .A1(n15161), .A2(n15287), .B1(n15157), .B2(n15289), .ZN(
        n15237) );
  OAI22_X1 U16384 ( .A1(n15242), .A2(n15003), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14989), .ZN(n14990) );
  AOI21_X1 U16385 ( .B1(n15237), .B2(n14991), .A(n14990), .ZN(n14992) );
  OAI211_X1 U16386 ( .C1(n8322), .C2(n14994), .A(n14993), .B(n14992), .ZN(
        P2_U3201) );
  NOR2_X1 U16387 ( .A1(n15011), .A2(n14995), .ZN(n14997) );
  AOI22_X1 U16388 ( .A1(n14998), .A2(n15000), .B1(n14997), .B2(n14996), .ZN(
        n15009) );
  INV_X1 U16389 ( .A(n14999), .ZN(n15008) );
  NAND2_X1 U16390 ( .A1(n15001), .A2(n15000), .ZN(n15007) );
  AOI22_X1 U16391 ( .A1(n15267), .A2(n15343), .B1(n15341), .B2(n15344), .ZN(
        n15307) );
  NOR2_X1 U16392 ( .A1(n15307), .A2(n15020), .ZN(n15005) );
  OAI22_X1 U16393 ( .A1(n15003), .A2(n15301), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n15002), .ZN(n15004) );
  AOI211_X1 U16394 ( .C1(n15304), .C2(n15024), .A(n15005), .B(n15004), .ZN(
        n15006) );
  OAI211_X1 U16395 ( .C1(n15009), .C2(n15008), .A(n15007), .B(n15006), .ZN(
        P2_U3205) );
  INV_X1 U16396 ( .A(n15010), .ZN(n15015) );
  NOR3_X1 U16397 ( .A1(n15012), .A2(n15161), .A3(n15011), .ZN(n15013) );
  AOI21_X1 U16398 ( .B1(n15015), .B2(n15014), .A(n15013), .ZN(n15026) );
  AND2_X1 U16399 ( .A1(n15134), .A2(n15341), .ZN(n15016) );
  AOI21_X1 U16400 ( .B1(n15017), .B2(n15343), .A(n15016), .ZN(n15207) );
  AOI22_X1 U16401 ( .A1(n15214), .A2(n15018), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3088), .ZN(n15019) );
  OAI21_X1 U16402 ( .B1(n15207), .B2(n15020), .A(n15019), .ZN(n15023) );
  MUX2_X1 U16403 ( .A(n15169), .B(P2_DATAO_REG_30__SCAN_IN), .S(n15044), .Z(
        P2_U3561) );
  MUX2_X1 U16404 ( .A(n15027), .B(P2_DATAO_REG_29__SCAN_IN), .S(n15044), .Z(
        P2_U3560) );
  MUX2_X1 U16405 ( .A(n15137), .B(P2_DATAO_REG_28__SCAN_IN), .S(n15044), .Z(
        P2_U3559) );
  MUX2_X1 U16406 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n15162), .S(P2_U3947), .Z(
        P2_U3557) );
  MUX2_X1 U16407 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n15134), .S(P2_U3947), .Z(
        P2_U3556) );
  MUX2_X1 U16408 ( .A(n15132), .B(P2_DATAO_REG_24__SCAN_IN), .S(n15044), .Z(
        P2_U3555) );
  MUX2_X1 U16409 ( .A(n15266), .B(P2_DATAO_REG_23__SCAN_IN), .S(n15044), .Z(
        P2_U3554) );
  MUX2_X1 U16410 ( .A(n15145), .B(P2_DATAO_REG_22__SCAN_IN), .S(n15044), .Z(
        P2_U3553) );
  MUX2_X1 U16411 ( .A(n15267), .B(P2_DATAO_REG_21__SCAN_IN), .S(n15044), .Z(
        P2_U3552) );
  MUX2_X1 U16412 ( .A(n15320), .B(P2_DATAO_REG_20__SCAN_IN), .S(n15044), .Z(
        P2_U3551) );
  MUX2_X1 U16413 ( .A(n15344), .B(P2_DATAO_REG_19__SCAN_IN), .S(n15044), .Z(
        P2_U3550) );
  MUX2_X1 U16414 ( .A(n15319), .B(P2_DATAO_REG_18__SCAN_IN), .S(n15044), .Z(
        P2_U3549) );
  MUX2_X1 U16415 ( .A(n15342), .B(P2_DATAO_REG_17__SCAN_IN), .S(n15044), .Z(
        P2_U3548) );
  MUX2_X1 U16416 ( .A(n15028), .B(P2_DATAO_REG_16__SCAN_IN), .S(n15044), .Z(
        P2_U3547) );
  MUX2_X1 U16417 ( .A(n15029), .B(P2_DATAO_REG_15__SCAN_IN), .S(n15044), .Z(
        P2_U3546) );
  MUX2_X1 U16418 ( .A(n15030), .B(P2_DATAO_REG_14__SCAN_IN), .S(n15044), .Z(
        P2_U3545) );
  MUX2_X1 U16419 ( .A(n15031), .B(P2_DATAO_REG_13__SCAN_IN), .S(n15044), .Z(
        P2_U3544) );
  MUX2_X1 U16420 ( .A(n15032), .B(P2_DATAO_REG_12__SCAN_IN), .S(n15044), .Z(
        P2_U3543) );
  MUX2_X1 U16421 ( .A(n15033), .B(P2_DATAO_REG_11__SCAN_IN), .S(n15044), .Z(
        P2_U3542) );
  MUX2_X1 U16422 ( .A(n15034), .B(P2_DATAO_REG_10__SCAN_IN), .S(n15044), .Z(
        P2_U3541) );
  MUX2_X1 U16423 ( .A(n15035), .B(P2_DATAO_REG_9__SCAN_IN), .S(n15044), .Z(
        P2_U3540) );
  MUX2_X1 U16424 ( .A(n15036), .B(P2_DATAO_REG_8__SCAN_IN), .S(n15044), .Z(
        P2_U3539) );
  MUX2_X1 U16425 ( .A(n15037), .B(P2_DATAO_REG_7__SCAN_IN), .S(n15044), .Z(
        P2_U3538) );
  MUX2_X1 U16426 ( .A(n15038), .B(P2_DATAO_REG_6__SCAN_IN), .S(n15044), .Z(
        P2_U3537) );
  MUX2_X1 U16427 ( .A(n15039), .B(P2_DATAO_REG_5__SCAN_IN), .S(n15044), .Z(
        P2_U3536) );
  MUX2_X1 U16428 ( .A(n15040), .B(P2_DATAO_REG_4__SCAN_IN), .S(n15044), .Z(
        P2_U3535) );
  MUX2_X1 U16429 ( .A(n15041), .B(P2_DATAO_REG_3__SCAN_IN), .S(n15044), .Z(
        P2_U3534) );
  MUX2_X1 U16430 ( .A(n15042), .B(P2_DATAO_REG_2__SCAN_IN), .S(n15044), .Z(
        P2_U3533) );
  MUX2_X1 U16431 ( .A(n15043), .B(P2_DATAO_REG_1__SCAN_IN), .S(n15044), .Z(
        P2_U3532) );
  MUX2_X1 U16432 ( .A(n13013), .B(P2_DATAO_REG_0__SCAN_IN), .S(n15044), .Z(
        P2_U3531) );
  MUX2_X1 U16433 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n10099), .S(n15045), .Z(
        n15046) );
  NAND3_X1 U16434 ( .A1(n15048), .A2(n15047), .A3(n15046), .ZN(n15049) );
  NAND3_X1 U16435 ( .A1(n16229), .A2(n15050), .A3(n15049), .ZN(n15061) );
  INV_X1 U16436 ( .A(n15051), .ZN(n15056) );
  NAND3_X1 U16437 ( .A1(n15054), .A2(n15053), .A3(n15052), .ZN(n15055) );
  NAND3_X1 U16438 ( .A1(n16233), .A2(n15056), .A3(n15055), .ZN(n15060) );
  AOI22_X1 U16439 ( .A1(n10096), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3088), .ZN(n15059) );
  NAND2_X1 U16440 ( .A1(n16231), .A2(n15057), .ZN(n15058) );
  NAND4_X1 U16441 ( .A1(n15061), .A2(n15060), .A3(n15059), .A4(n15058), .ZN(
        P2_U3216) );
  INV_X1 U16442 ( .A(n15062), .ZN(n15064) );
  NOR2_X1 U16443 ( .A1(n16214), .A2(n15069), .ZN(n15063) );
  AOI211_X1 U16444 ( .C1(n10096), .C2(P2_ADDR_REG_4__SCAN_IN), .A(n15064), .B(
        n15063), .ZN(n15075) );
  INV_X1 U16445 ( .A(n15088), .ZN(n15068) );
  NAND3_X1 U16446 ( .A1(n16164), .A2(n15066), .A3(n15065), .ZN(n15067) );
  NAND3_X1 U16447 ( .A1(n16233), .A2(n15068), .A3(n15067), .ZN(n15074) );
  MUX2_X1 U16448 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n11289), .S(n15069), .Z(
        n15070) );
  NAND3_X1 U16449 ( .A1(n16165), .A2(n15071), .A3(n15070), .ZN(n15072) );
  NAND3_X1 U16450 ( .A1(n16229), .A2(n15081), .A3(n15072), .ZN(n15073) );
  NAND3_X1 U16451 ( .A1(n15075), .A2(n15074), .A3(n15073), .ZN(P2_U3218) );
  NAND2_X1 U16452 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3088), .ZN(n15076) );
  OAI21_X1 U16453 ( .B1(n16214), .B2(n15077), .A(n15076), .ZN(n15078) );
  AOI21_X1 U16454 ( .B1(n10096), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n15078), .ZN(
        n15091) );
  MUX2_X1 U16455 ( .A(n10108), .B(P2_REG2_REG_5__SCAN_IN), .S(n15083), .Z(
        n15079) );
  NAND3_X1 U16456 ( .A1(n15081), .A2(n15080), .A3(n15079), .ZN(n15082) );
  NAND3_X1 U16457 ( .A1(n16229), .A2(n15094), .A3(n15082), .ZN(n15090) );
  MUX2_X1 U16458 ( .A(n10087), .B(P2_REG1_REG_5__SCAN_IN), .S(n15083), .Z(
        n15086) );
  INV_X1 U16459 ( .A(n15084), .ZN(n15085) );
  NAND2_X1 U16460 ( .A1(n15086), .A2(n15085), .ZN(n15087) );
  OAI211_X1 U16461 ( .C1(n15088), .C2(n15087), .A(n16233), .B(n15100), .ZN(
        n15089) );
  NAND3_X1 U16462 ( .A1(n15091), .A2(n15090), .A3(n15089), .ZN(P2_U3219) );
  MUX2_X1 U16463 ( .A(n11273), .B(P2_REG2_REG_6__SCAN_IN), .S(n15105), .Z(
        n15092) );
  NAND3_X1 U16464 ( .A1(n15094), .A2(n15093), .A3(n15092), .ZN(n15095) );
  NAND3_X1 U16465 ( .A1(n16229), .A2(n15096), .A3(n15095), .ZN(n15109) );
  INV_X1 U16466 ( .A(n15097), .ZN(n15102) );
  NAND3_X1 U16467 ( .A1(n15100), .A2(n15099), .A3(n15098), .ZN(n15101) );
  NAND3_X1 U16468 ( .A1(n16233), .A2(n15102), .A3(n15101), .ZN(n15108) );
  INV_X1 U16469 ( .A(n15103), .ZN(n15104) );
  AOI21_X1 U16470 ( .B1(n10096), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n15104), .ZN(
        n15107) );
  NAND2_X1 U16471 ( .A1(n16231), .A2(n15105), .ZN(n15106) );
  NAND4_X1 U16472 ( .A1(n15109), .A2(n15108), .A3(n15107), .A4(n15106), .ZN(
        P2_U3220) );
  NAND2_X1 U16473 ( .A1(n15500), .A2(n15328), .ZN(n15311) );
  OR2_X1 U16474 ( .A1(n10090), .A2(n15112), .ZN(n15113) );
  NAND2_X1 U16475 ( .A1(n15343), .A2(n15113), .ZN(n15171) );
  INV_X1 U16476 ( .A(n15171), .ZN(n15115) );
  NAND2_X1 U16477 ( .A1(n15115), .A2(n15114), .ZN(n15380) );
  NOR2_X1 U16478 ( .A1(n15362), .A2(n15380), .ZN(n15120) );
  NOR2_X1 U16479 ( .A1(n15468), .A2(n15330), .ZN(n15116) );
  AOI211_X1 U16480 ( .C1(n15362), .C2(P2_REG2_REG_31__SCAN_IN), .A(n15120), 
        .B(n15116), .ZN(n15117) );
  OAI21_X1 U16481 ( .B1(n15377), .B2(n15233), .A(n15117), .ZN(P2_U3234) );
  OAI211_X1 U16482 ( .C1(n15472), .C2(n15139), .A(n14960), .B(n15118), .ZN(
        n15381) );
  NOR2_X1 U16483 ( .A1(n15472), .A2(n15330), .ZN(n15119) );
  AOI211_X1 U16484 ( .C1(n15362), .C2(P2_REG2_REG_30__SCAN_IN), .A(n15120), 
        .B(n15119), .ZN(n15121) );
  OAI21_X1 U16485 ( .B1(n15233), .B2(n15381), .A(n15121), .ZN(P2_U3235) );
  INV_X1 U16486 ( .A(n15339), .ZN(n15348) );
  OR2_X1 U16487 ( .A1(n15329), .A2(n15344), .ZN(n15123) );
  NAND2_X1 U16488 ( .A1(n15300), .A2(n15299), .ZN(n15125) );
  OR2_X1 U16489 ( .A1(n15304), .A2(n15320), .ZN(n15124) );
  NOR2_X1 U16490 ( .A1(n15291), .A2(n15267), .ZN(n15126) );
  NAND2_X1 U16491 ( .A1(n15291), .A2(n15267), .ZN(n15127) );
  NAND2_X1 U16492 ( .A1(n15424), .A2(n15145), .ZN(n15128) );
  AND2_X1 U16493 ( .A1(n15256), .A2(n15266), .ZN(n15129) );
  OR2_X1 U16494 ( .A1(n15256), .A2(n15266), .ZN(n15130) );
  NAND2_X1 U16495 ( .A1(n15414), .A2(n15132), .ZN(n15133) );
  INV_X1 U16496 ( .A(n15220), .ZN(n15225) );
  OR2_X1 U16497 ( .A1(n15408), .A2(n15134), .ZN(n15135) );
  INV_X1 U16498 ( .A(n15193), .ZN(n15164) );
  AOI211_X1 U16499 ( .C1(n15386), .C2(n15183), .A(n14937), .B(n15139), .ZN(
        n15385) );
  INV_X1 U16500 ( .A(n15386), .ZN(n15143) );
  INV_X1 U16501 ( .A(n15140), .ZN(n15141) );
  AOI22_X1 U16502 ( .A1(n15141), .A2(n15292), .B1(P2_REG2_REG_29__SCAN_IN), 
        .B2(n15362), .ZN(n15142) );
  OAI21_X1 U16503 ( .B1(n15143), .B2(n15330), .A(n15142), .ZN(n15144) );
  AOI21_X1 U16504 ( .B1(n15385), .B2(n15371), .A(n15144), .ZN(n15176) );
  NAND2_X1 U16505 ( .A1(n15269), .A2(n15145), .ZN(n15156) );
  INV_X1 U16506 ( .A(n15299), .ZN(n15306) );
  NOR2_X1 U16507 ( .A1(n8008), .A2(n8760), .ZN(n15147) );
  NAND2_X1 U16508 ( .A1(n15444), .A2(n15150), .ZN(n15321) );
  OR2_X1 U16509 ( .A1(n15304), .A2(n15288), .ZN(n15152) );
  NAND2_X1 U16510 ( .A1(n15291), .A2(n15153), .ZN(n15154) );
  NAND2_X1 U16511 ( .A1(n15424), .A2(n15286), .ZN(n15155) );
  NAND2_X1 U16512 ( .A1(n15256), .A2(n15157), .ZN(n15158) );
  NAND2_X1 U16513 ( .A1(n15414), .A2(n15159), .ZN(n15160) );
  NAND2_X1 U16514 ( .A1(n15180), .A2(n15179), .ZN(n15178) );
  INV_X1 U16515 ( .A(n15169), .ZN(n15170) );
  INV_X1 U16516 ( .A(n15173), .ZN(n15174) );
  NAND2_X1 U16517 ( .A1(n15384), .A2(n15353), .ZN(n15175) );
  OAI211_X1 U16518 ( .C1(n15387), .C2(n15359), .A(n15176), .B(n15175), .ZN(
        P2_U3236) );
  XNOR2_X1 U16519 ( .A(n15177), .B(n15179), .ZN(n15392) );
  INV_X1 U16520 ( .A(n15392), .ZN(n15189) );
  OAI211_X1 U16521 ( .C1(n15180), .C2(n15179), .A(n15178), .B(n15346), .ZN(
        n15390) );
  INV_X1 U16522 ( .A(n15181), .ZN(n15389) );
  OAI211_X1 U16523 ( .C1(n15364), .C2(n15182), .A(n15390), .B(n15389), .ZN(
        n15187) );
  OAI211_X1 U16524 ( .C1(n15477), .C2(n15198), .A(n14960), .B(n15183), .ZN(
        n15388) );
  AOI22_X1 U16525 ( .A1(n15184), .A2(n15367), .B1(P2_REG2_REG_28__SCAN_IN), 
        .B2(n15362), .ZN(n15185) );
  OAI21_X1 U16526 ( .B1(n15388), .B2(n15233), .A(n15185), .ZN(n15186) );
  AOI21_X1 U16527 ( .B1(n15187), .B2(n15353), .A(n15186), .ZN(n15188) );
  OAI21_X1 U16528 ( .B1(n15189), .B2(n15359), .A(n15188), .ZN(P2_U3237) );
  XNOR2_X1 U16529 ( .A(n15190), .B(n15193), .ZN(n15192) );
  OAI21_X1 U16530 ( .B1(n15192), .B2(n15308), .A(n15191), .ZN(n15395) );
  INV_X1 U16531 ( .A(n15395), .ZN(n15204) );
  XNOR2_X1 U16532 ( .A(n15194), .B(n15193), .ZN(n15397) );
  NAND2_X1 U16533 ( .A1(n15212), .A2(n15195), .ZN(n15196) );
  NAND2_X1 U16534 ( .A1(n15196), .A2(n14960), .ZN(n15197) );
  NOR2_X1 U16535 ( .A1(n15198), .A2(n15197), .ZN(n15396) );
  NAND2_X1 U16536 ( .A1(n15396), .A2(n15371), .ZN(n15201) );
  AOI22_X1 U16537 ( .A1(n15199), .A2(n15292), .B1(P2_REG2_REG_27__SCAN_IN), 
        .B2(n15362), .ZN(n15200) );
  OAI211_X1 U16538 ( .C1(n15481), .C2(n15330), .A(n15201), .B(n15200), .ZN(
        n15202) );
  AOI21_X1 U16539 ( .B1(n15397), .B2(n15369), .A(n15202), .ZN(n15203) );
  OAI21_X1 U16540 ( .B1(n15204), .B2(n15362), .A(n15203), .ZN(P2_U3238) );
  XNOR2_X1 U16541 ( .A(n15205), .B(n15209), .ZN(n15206) );
  NAND2_X1 U16542 ( .A1(n15206), .A2(n15346), .ZN(n15208) );
  NAND2_X1 U16543 ( .A1(n15208), .A2(n15207), .ZN(n15402) );
  INV_X1 U16544 ( .A(n15402), .ZN(n15219) );
  XNOR2_X1 U16545 ( .A(n15210), .B(n15209), .ZN(n15400) );
  AOI21_X1 U16546 ( .B1(n15227), .B2(n15211), .A(n14937), .ZN(n15213) );
  AND2_X1 U16547 ( .A1(n15213), .A2(n15212), .ZN(n15401) );
  NAND2_X1 U16548 ( .A1(n15401), .A2(n15371), .ZN(n15216) );
  AOI22_X1 U16549 ( .A1(n15214), .A2(n15292), .B1(P2_REG2_REG_26__SCAN_IN), 
        .B2(n15362), .ZN(n15215) );
  OAI211_X1 U16550 ( .C1(n15485), .C2(n15330), .A(n15216), .B(n15215), .ZN(
        n15217) );
  AOI21_X1 U16551 ( .B1(n15400), .B2(n15369), .A(n15217), .ZN(n15218) );
  OAI21_X1 U16552 ( .B1(n15362), .B2(n15219), .A(n15218), .ZN(P2_U3239) );
  XNOR2_X1 U16553 ( .A(n15221), .B(n15220), .ZN(n15223) );
  AOI21_X1 U16554 ( .B1(n15223), .B2(n15346), .A(n15222), .ZN(n15411) );
  OAI21_X1 U16555 ( .B1(n15226), .B2(n15225), .A(n15224), .ZN(n15407) );
  OAI211_X1 U16556 ( .C1(n15246), .C2(n15228), .A(n14960), .B(n15227), .ZN(
        n15410) );
  INV_X1 U16557 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n15229) );
  OAI22_X1 U16558 ( .A1(n15230), .A2(n15364), .B1(n15229), .B2(n15353), .ZN(
        n15231) );
  AOI21_X1 U16559 ( .B1(n15408), .B2(n15367), .A(n15231), .ZN(n15232) );
  OAI21_X1 U16560 ( .B1(n15410), .B2(n15233), .A(n15232), .ZN(n15234) );
  AOI21_X1 U16561 ( .B1(n15407), .B2(n15369), .A(n15234), .ZN(n15235) );
  OAI21_X1 U16562 ( .B1(n15362), .B2(n15411), .A(n15235), .ZN(P2_U3240) );
  XNOR2_X1 U16563 ( .A(n15236), .B(n15239), .ZN(n15238) );
  AOI21_X1 U16564 ( .B1(n15238), .B2(n15346), .A(n15237), .ZN(n15416) );
  OAI21_X1 U16565 ( .B1(n7520), .B2(n8770), .A(n15240), .ZN(n15417) );
  INV_X1 U16566 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n15241) );
  OAI22_X1 U16567 ( .A1(n15242), .A2(n15364), .B1(n15241), .B2(n15327), .ZN(
        n15243) );
  AOI21_X1 U16568 ( .B1(n15414), .B2(n15367), .A(n15243), .ZN(n15248) );
  NAND2_X1 U16569 ( .A1(n15257), .A2(n15414), .ZN(n15244) );
  NAND2_X1 U16570 ( .A1(n15244), .A2(n14960), .ZN(n15245) );
  NOR2_X1 U16571 ( .A1(n15246), .A2(n15245), .ZN(n15413) );
  NAND2_X1 U16572 ( .A1(n15413), .A2(n15371), .ZN(n15247) );
  OAI211_X1 U16573 ( .C1(n15417), .C2(n15359), .A(n15248), .B(n15247), .ZN(
        n15249) );
  INV_X1 U16574 ( .A(n15249), .ZN(n15250) );
  OAI21_X1 U16575 ( .B1(n15362), .B2(n15416), .A(n15250), .ZN(P2_U3241) );
  XNOR2_X1 U16576 ( .A(n15251), .B(n15254), .ZN(n15253) );
  OAI21_X1 U16577 ( .B1(n15253), .B2(n15308), .A(n15252), .ZN(n15418) );
  INV_X1 U16578 ( .A(n15418), .ZN(n15264) );
  XNOR2_X1 U16579 ( .A(n15255), .B(n15254), .ZN(n15420) );
  INV_X1 U16580 ( .A(n15256), .ZN(n15491) );
  AOI21_X1 U16581 ( .B1(n15256), .B2(n15274), .A(n14937), .ZN(n15258) );
  AND2_X1 U16582 ( .A1(n15258), .A2(n15257), .ZN(n15419) );
  NAND2_X1 U16583 ( .A1(n15419), .A2(n15371), .ZN(n15261) );
  AOI22_X1 U16584 ( .A1(n15259), .A2(n15292), .B1(n15362), .B2(
        P2_REG2_REG_23__SCAN_IN), .ZN(n15260) );
  OAI211_X1 U16585 ( .C1(n15491), .C2(n15330), .A(n15261), .B(n15260), .ZN(
        n15262) );
  AOI21_X1 U16586 ( .B1(n15420), .B2(n15369), .A(n15262), .ZN(n15263) );
  OAI21_X1 U16587 ( .B1(n15264), .B2(n15362), .A(n15263), .ZN(P2_U3242) );
  XNOR2_X1 U16588 ( .A(n15265), .B(n15269), .ZN(n15268) );
  AOI222_X1 U16589 ( .A1(n15346), .A2(n15268), .B1(n15267), .B2(n15341), .C1(
        n15266), .C2(n15343), .ZN(n15426) );
  XNOR2_X1 U16590 ( .A(n15270), .B(n15269), .ZN(n15427) );
  INV_X1 U16591 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n15272) );
  OAI22_X1 U16592 ( .A1(n15353), .A2(n15272), .B1(n15271), .B2(n15364), .ZN(
        n15273) );
  AOI21_X1 U16593 ( .B1(n15424), .B2(n15367), .A(n15273), .ZN(n15277) );
  AOI21_X1 U16594 ( .B1(n15424), .B2(n15290), .A(n14937), .ZN(n15275) );
  AND2_X1 U16595 ( .A1(n15275), .A2(n15274), .ZN(n15423) );
  NAND2_X1 U16596 ( .A1(n15423), .A2(n15371), .ZN(n15276) );
  OAI211_X1 U16597 ( .C1(n15427), .C2(n15359), .A(n15277), .B(n15276), .ZN(
        n15278) );
  INV_X1 U16598 ( .A(n15278), .ZN(n15279) );
  OAI21_X1 U16599 ( .B1(n15426), .B2(n15362), .A(n15279), .ZN(P2_U3243) );
  XNOR2_X1 U16600 ( .A(n15280), .B(n15284), .ZN(n15430) );
  INV_X1 U16601 ( .A(n15430), .ZN(n15298) );
  INV_X1 U16602 ( .A(n15281), .ZN(n15282) );
  AOI21_X1 U16603 ( .B1(n15284), .B2(n15283), .A(n15282), .ZN(n15285) );
  OAI222_X1 U16604 ( .A1(n15289), .A2(n15288), .B1(n15287), .B2(n15286), .C1(
        n15308), .C2(n15285), .ZN(n15428) );
  AOI211_X1 U16605 ( .C1(n15291), .C2(n15311), .A(n14937), .B(n8325), .ZN(
        n15429) );
  NAND2_X1 U16606 ( .A1(n15429), .A2(n15371), .ZN(n15295) );
  AOI22_X1 U16607 ( .A1(n15362), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n15293), 
        .B2(n15292), .ZN(n15294) );
  OAI211_X1 U16608 ( .C1(n15496), .C2(n15330), .A(n15295), .B(n15294), .ZN(
        n15296) );
  AOI21_X1 U16609 ( .B1(n15428), .B2(n15353), .A(n15296), .ZN(n15297) );
  OAI21_X1 U16610 ( .B1(n15359), .B2(n15298), .A(n15297), .ZN(P2_U3244) );
  XNOR2_X1 U16611 ( .A(n15300), .B(n15299), .ZN(n15435) );
  NAND2_X1 U16612 ( .A1(n15435), .A2(n15369), .ZN(n15315) );
  INV_X1 U16613 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n15302) );
  OAI22_X1 U16614 ( .A1(n15353), .A2(n15302), .B1(n15301), .B2(n15364), .ZN(
        n15303) );
  AOI21_X1 U16615 ( .B1(n15304), .B2(n15367), .A(n15303), .ZN(n15314) );
  XNOR2_X1 U16616 ( .A(n15305), .B(n15306), .ZN(n15309) );
  OAI21_X1 U16617 ( .B1(n15309), .B2(n15308), .A(n15307), .ZN(n15433) );
  NAND2_X1 U16618 ( .A1(n15433), .A2(n15353), .ZN(n15313) );
  OR2_X1 U16619 ( .A1(n15500), .A2(n15328), .ZN(n15310) );
  AND3_X1 U16620 ( .A1(n15311), .A2(n15310), .A3(n14960), .ZN(n15434) );
  NAND2_X1 U16621 ( .A1(n15434), .A2(n15371), .ZN(n15312) );
  NAND4_X1 U16622 ( .A1(n15315), .A2(n15314), .A3(n15313), .A4(n15312), .ZN(
        P2_U3245) );
  OAI21_X1 U16623 ( .B1(n15318), .B2(n15317), .A(n15316), .ZN(n15440) );
  INV_X1 U16624 ( .A(n15440), .ZN(n15337) );
  AOI22_X1 U16625 ( .A1(n15320), .A2(n15343), .B1(n15341), .B2(n15319), .ZN(
        n15326) );
  AND2_X1 U16626 ( .A1(n15338), .A2(n15321), .ZN(n15323) );
  OAI211_X1 U16627 ( .C1(n15324), .C2(n15323), .A(n15322), .B(n15346), .ZN(
        n15325) );
  OAI211_X1 U16628 ( .C1(n15337), .C2(n10226), .A(n15326), .B(n15325), .ZN(
        n15438) );
  NAND2_X1 U16629 ( .A1(n15438), .A2(n15327), .ZN(n15335) );
  AOI211_X1 U16630 ( .C1(n15329), .C2(n15355), .A(n14937), .B(n15328), .ZN(
        n15439) );
  NOR2_X1 U16631 ( .A1(n15504), .A2(n15330), .ZN(n15333) );
  OAI22_X1 U16632 ( .A1(n15353), .A2(n12113), .B1(n15331), .B2(n15364), .ZN(
        n15332) );
  AOI211_X1 U16633 ( .C1(n15439), .C2(n15371), .A(n15333), .B(n15332), .ZN(
        n15334) );
  OAI211_X1 U16634 ( .C1(n15337), .C2(n15336), .A(n15335), .B(n15334), .ZN(
        P2_U3246) );
  OAI21_X1 U16635 ( .B1(n15340), .B2(n15339), .A(n15338), .ZN(n15345) );
  AOI222_X1 U16636 ( .A1(n15346), .A2(n15345), .B1(n15344), .B2(n15343), .C1(
        n15342), .C2(n15341), .ZN(n15446) );
  OAI21_X1 U16637 ( .B1(n15349), .B2(n15348), .A(n15347), .ZN(n15350) );
  INV_X1 U16638 ( .A(n15350), .ZN(n15447) );
  OAI22_X1 U16639 ( .A1(n15353), .A2(n15352), .B1(n15351), .B2(n15364), .ZN(
        n15354) );
  AOI21_X1 U16640 ( .B1(n15444), .B2(n15367), .A(n15354), .ZN(n15358) );
  AOI21_X1 U16641 ( .B1(n15444), .B2(n7668), .A(n14937), .ZN(n15356) );
  AND2_X1 U16642 ( .A1(n15356), .A2(n15355), .ZN(n15443) );
  NAND2_X1 U16643 ( .A1(n15443), .A2(n15371), .ZN(n15357) );
  OAI211_X1 U16644 ( .C1(n15447), .C2(n15359), .A(n15358), .B(n15357), .ZN(
        n15360) );
  INV_X1 U16645 ( .A(n15360), .ZN(n15361) );
  OAI21_X1 U16646 ( .B1(n15362), .B2(n15446), .A(n15361), .ZN(P2_U3247) );
  NAND2_X1 U16647 ( .A1(n15363), .A2(n15353), .ZN(n15376) );
  OAI22_X1 U16648 ( .A1(n15353), .A2(n10767), .B1(n15365), .B2(n15364), .ZN(
        n15366) );
  AOI21_X1 U16649 ( .B1(n15368), .B2(n15367), .A(n15366), .ZN(n15375) );
  NAND2_X1 U16650 ( .A1(n15370), .A2(n15369), .ZN(n15374) );
  NAND2_X1 U16651 ( .A1(n15372), .A2(n15371), .ZN(n15373) );
  NAND4_X1 U16652 ( .A1(n15376), .A2(n15375), .A3(n15374), .A4(n15373), .ZN(
        P2_U3254) );
  NAND2_X1 U16653 ( .A1(n15377), .A2(n15380), .ZN(n15465) );
  MUX2_X1 U16654 ( .A(n15465), .B(P2_REG1_REG_31__SCAN_IN), .S(n16746), .Z(
        n15378) );
  INV_X1 U16655 ( .A(n15378), .ZN(n15379) );
  OAI21_X1 U16656 ( .B1(n15468), .B2(n15464), .A(n15379), .ZN(P2_U3530) );
  AND2_X1 U16657 ( .A1(n15381), .A2(n15380), .ZN(n15469) );
  MUX2_X1 U16658 ( .A(n15382), .B(n15469), .S(n16747), .Z(n15383) );
  OAI21_X1 U16659 ( .B1(n15472), .B2(n15464), .A(n15383), .ZN(P2_U3529) );
  MUX2_X1 U16660 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n15473), .S(n16747), .Z(
        P2_U3528) );
  NAND3_X1 U16661 ( .A1(n15390), .A2(n15389), .A3(n15388), .ZN(n15391) );
  AOI21_X1 U16662 ( .B1(n15392), .B2(n16641), .A(n15391), .ZN(n15474) );
  MUX2_X1 U16663 ( .A(n15393), .B(n15474), .S(n16747), .Z(n15394) );
  AOI211_X1 U16664 ( .C1(n15397), .C2(n16641), .A(n15396), .B(n15395), .ZN(
        n15478) );
  MUX2_X1 U16665 ( .A(n15398), .B(n15478), .S(n16747), .Z(n15399) );
  OAI21_X1 U16666 ( .B1(n15481), .B2(n15464), .A(n15399), .ZN(P2_U3526) );
  NAND2_X1 U16667 ( .A1(n15400), .A2(n16641), .ZN(n15404) );
  NOR2_X1 U16668 ( .A1(n15402), .A2(n15401), .ZN(n15403) );
  NAND2_X1 U16669 ( .A1(n15404), .A2(n15403), .ZN(n15482) );
  MUX2_X1 U16670 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n15482), .S(n16747), .Z(
        n15405) );
  INV_X1 U16671 ( .A(n15405), .ZN(n15406) );
  OAI21_X1 U16672 ( .B1(n15485), .B2(n15464), .A(n15406), .ZN(P2_U3525) );
  NAND2_X1 U16673 ( .A1(n15407), .A2(n16641), .ZN(n15412) );
  NAND2_X1 U16674 ( .A1(n15408), .A2(n16740), .ZN(n15409) );
  NAND4_X1 U16675 ( .A1(n15412), .A2(n15411), .A3(n15410), .A4(n15409), .ZN(
        n15486) );
  MUX2_X1 U16676 ( .A(n15486), .B(P2_REG1_REG_25__SCAN_IN), .S(n16746), .Z(
        P2_U3524) );
  AOI21_X1 U16677 ( .B1(n16740), .B2(n15414), .A(n15413), .ZN(n15415) );
  OAI211_X1 U16678 ( .C1(n15417), .C2(n16738), .A(n15416), .B(n15415), .ZN(
        n15487) );
  MUX2_X1 U16679 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n15487), .S(n16747), .Z(
        P2_U3523) );
  AOI211_X1 U16680 ( .C1(n16641), .C2(n15420), .A(n15419), .B(n15418), .ZN(
        n15488) );
  MUX2_X1 U16681 ( .A(n15421), .B(n15488), .S(n16747), .Z(n15422) );
  OAI21_X1 U16682 ( .B1(n15491), .B2(n15464), .A(n15422), .ZN(P2_U3522) );
  AOI21_X1 U16683 ( .B1(n16740), .B2(n15424), .A(n15423), .ZN(n15425) );
  OAI211_X1 U16684 ( .C1(n16738), .C2(n15427), .A(n15426), .B(n15425), .ZN(
        n15492) );
  MUX2_X1 U16685 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n15492), .S(n16747), .Z(
        P2_U3521) );
  AOI211_X1 U16686 ( .C1(n15430), .C2(n16641), .A(n15429), .B(n15428), .ZN(
        n15493) );
  MUX2_X1 U16687 ( .A(n15431), .B(n15493), .S(n16747), .Z(n15432) );
  OAI21_X1 U16688 ( .B1(n15496), .B2(n15464), .A(n15432), .ZN(P2_U3520) );
  AOI211_X1 U16689 ( .C1(n15435), .C2(n16641), .A(n15434), .B(n15433), .ZN(
        n15497) );
  MUX2_X1 U16690 ( .A(n15436), .B(n15497), .S(n16747), .Z(n15437) );
  OAI21_X1 U16691 ( .B1(n15500), .B2(n15464), .A(n15437), .ZN(P2_U3519) );
  INV_X1 U16692 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n15441) );
  AOI211_X1 U16693 ( .C1(n16704), .C2(n15440), .A(n15439), .B(n15438), .ZN(
        n15501) );
  MUX2_X1 U16694 ( .A(n15441), .B(n15501), .S(n16747), .Z(n15442) );
  OAI21_X1 U16695 ( .B1(n15504), .B2(n15464), .A(n15442), .ZN(P2_U3518) );
  AOI21_X1 U16696 ( .B1(n16740), .B2(n15444), .A(n15443), .ZN(n15445) );
  OAI211_X1 U16697 ( .C1(n15447), .C2(n16738), .A(n15446), .B(n15445), .ZN(
        n15505) );
  MUX2_X1 U16698 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n15505), .S(n16747), .Z(
        P2_U3517) );
  AOI211_X1 U16699 ( .C1(n16641), .C2(n15450), .A(n15449), .B(n15448), .ZN(
        n15506) );
  MUX2_X1 U16700 ( .A(n15451), .B(n15506), .S(n16747), .Z(n15452) );
  OAI21_X1 U16701 ( .B1(n8761), .B2(n15464), .A(n15452), .ZN(P2_U3516) );
  OAI211_X1 U16702 ( .C1(n15455), .C2(n16738), .A(n15454), .B(n15453), .ZN(
        n15509) );
  MUX2_X1 U16703 ( .A(n15509), .B(P2_REG1_REG_16__SCAN_IN), .S(n16746), .Z(
        n15456) );
  AOI21_X1 U16704 ( .B1(n15457), .B2(n15511), .A(n15456), .ZN(n15458) );
  INV_X1 U16705 ( .A(n15458), .ZN(P2_U3515) );
  INV_X1 U16706 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n15462) );
  AOI211_X1 U16707 ( .C1(n16704), .C2(n15461), .A(n15460), .B(n15459), .ZN(
        n15514) );
  MUX2_X1 U16708 ( .A(n15462), .B(n15514), .S(n16747), .Z(n15463) );
  OAI21_X1 U16709 ( .B1(n15518), .B2(n15464), .A(n15463), .ZN(P2_U3514) );
  MUX2_X1 U16710 ( .A(n15465), .B(P2_REG0_REG_31__SCAN_IN), .S(n16748), .Z(
        n15466) );
  INV_X1 U16711 ( .A(n15466), .ZN(n15467) );
  OAI21_X1 U16712 ( .B1(n15468), .B2(n15517), .A(n15467), .ZN(P2_U3498) );
  INV_X1 U16713 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n15470) );
  MUX2_X1 U16714 ( .A(n15470), .B(n15469), .S(n16751), .Z(n15471) );
  OAI21_X1 U16715 ( .B1(n15472), .B2(n15517), .A(n15471), .ZN(P2_U3497) );
  MUX2_X1 U16716 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n15473), .S(n16751), .Z(
        P2_U3496) );
  INV_X1 U16717 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n15475) );
  MUX2_X1 U16718 ( .A(n15475), .B(n15474), .S(n16751), .Z(n15476) );
  INV_X1 U16719 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n15479) );
  MUX2_X1 U16720 ( .A(n15479), .B(n15478), .S(n16751), .Z(n15480) );
  OAI21_X1 U16721 ( .B1(n15481), .B2(n15517), .A(n15480), .ZN(P2_U3494) );
  MUX2_X1 U16722 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n15482), .S(n16751), .Z(
        n15483) );
  INV_X1 U16723 ( .A(n15483), .ZN(n15484) );
  OAI21_X1 U16724 ( .B1(n15485), .B2(n15517), .A(n15484), .ZN(P2_U3493) );
  MUX2_X1 U16725 ( .A(n15486), .B(P2_REG0_REG_25__SCAN_IN), .S(n16748), .Z(
        P2_U3492) );
  MUX2_X1 U16726 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n15487), .S(n16751), .Z(
        P2_U3491) );
  INV_X1 U16727 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n15489) );
  MUX2_X1 U16728 ( .A(n15489), .B(n15488), .S(n16751), .Z(n15490) );
  OAI21_X1 U16729 ( .B1(n15491), .B2(n15517), .A(n15490), .ZN(P2_U3490) );
  MUX2_X1 U16730 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n15492), .S(n16751), .Z(
        P2_U3489) );
  INV_X1 U16731 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n15494) );
  MUX2_X1 U16732 ( .A(n15494), .B(n15493), .S(n16751), .Z(n15495) );
  OAI21_X1 U16733 ( .B1(n15496), .B2(n15517), .A(n15495), .ZN(P2_U3488) );
  INV_X1 U16734 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n15498) );
  MUX2_X1 U16735 ( .A(n15498), .B(n15497), .S(n16751), .Z(n15499) );
  OAI21_X1 U16736 ( .B1(n15500), .B2(n15517), .A(n15499), .ZN(P2_U3487) );
  INV_X1 U16737 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n15502) );
  MUX2_X1 U16738 ( .A(n15502), .B(n15501), .S(n16751), .Z(n15503) );
  OAI21_X1 U16739 ( .B1(n15504), .B2(n15517), .A(n15503), .ZN(P2_U3486) );
  MUX2_X1 U16740 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n15505), .S(n16751), .Z(
        P2_U3484) );
  INV_X1 U16741 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n15507) );
  MUX2_X1 U16742 ( .A(n15507), .B(n15506), .S(n16751), .Z(n15508) );
  OAI21_X1 U16743 ( .B1(n8761), .B2(n15517), .A(n15508), .ZN(P2_U3481) );
  MUX2_X1 U16744 ( .A(n15509), .B(P2_REG0_REG_16__SCAN_IN), .S(n16748), .Z(
        n15510) );
  AOI21_X1 U16745 ( .B1(n15512), .B2(n15511), .A(n15510), .ZN(n15513) );
  INV_X1 U16746 ( .A(n15513), .ZN(P2_U3478) );
  INV_X1 U16747 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n15515) );
  MUX2_X1 U16748 ( .A(n15515), .B(n15514), .S(n16751), .Z(n15516) );
  OAI21_X1 U16749 ( .B1(n15518), .B2(n15517), .A(n15516), .ZN(P2_U3475) );
  INV_X1 U16750 ( .A(n15519), .ZN(n15523) );
  NOR4_X1 U16751 ( .A1(n15520), .A2(P2_IR_REG_30__SCAN_IN), .A3(n9715), .A4(
        P2_U3088), .ZN(n15521) );
  AOI21_X1 U16752 ( .B1(n15528), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n15521), 
        .ZN(n15522) );
  OAI21_X1 U16753 ( .B1(n15523), .B2(n15540), .A(n15522), .ZN(P2_U3296) );
  INV_X1 U16754 ( .A(n15524), .ZN(n16122) );
  OAI222_X1 U16755 ( .A1(n15540), .A2(n16122), .B1(P2_U3088), .B2(n15526), 
        .C1(n15525), .C2(n15545), .ZN(P2_U3297) );
  AOI21_X1 U16756 ( .B1(n15528), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n15527), 
        .ZN(n15529) );
  OAI21_X1 U16757 ( .B1(n15530), .B2(n15540), .A(n15529), .ZN(P2_U3299) );
  INV_X1 U16758 ( .A(n15531), .ZN(n16124) );
  OAI222_X1 U16759 ( .A1(n15545), .A2(n10579), .B1(n15540), .B2(n16124), .C1(
        n10090), .C2(P2_U3088), .ZN(P2_U3300) );
  INV_X1 U16760 ( .A(n15532), .ZN(n16126) );
  OAI222_X1 U16761 ( .A1(P2_U3088), .A2(n15534), .B1(n15540), .B2(n16126), 
        .C1(n15533), .C2(n15545), .ZN(P2_U3301) );
  INV_X1 U16762 ( .A(n15535), .ZN(n16130) );
  OAI222_X1 U16763 ( .A1(n15545), .A2(n15537), .B1(n15540), .B2(n16130), .C1(
        P2_U3088), .C2(n15536), .ZN(P2_U3302) );
  INV_X1 U16764 ( .A(n15538), .ZN(n16133) );
  OAI222_X1 U16765 ( .A1(n15545), .A2(n15541), .B1(n15540), .B2(n16133), .C1(
        P2_U3088), .C2(n15539), .ZN(P2_U3303) );
  NAND2_X1 U16766 ( .A1(n16136), .A2(n15542), .ZN(n15544) );
  OAI211_X1 U16767 ( .C1(n8582), .C2(n15545), .A(n15544), .B(n15543), .ZN(
        P2_U3304) );
  INV_X1 U16768 ( .A(n15546), .ZN(n15547) );
  MUX2_X1 U16769 ( .A(n15547), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  INV_X1 U16770 ( .A(n16528), .ZN(n15622) );
  OAI21_X1 U16771 ( .B1(n15550), .B2(n15549), .A(n15548), .ZN(n15551) );
  NAND2_X1 U16772 ( .A1(n15551), .A2(n16531), .ZN(n15556) );
  NOR2_X1 U16773 ( .A1(n16535), .A2(n15820), .ZN(n15554) );
  OAI22_X1 U16774 ( .A1(n15648), .A2(n15815), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15552), .ZN(n15553) );
  AOI211_X1 U16775 ( .C1(n15659), .C2(n15765), .A(n15554), .B(n15553), .ZN(
        n15555) );
  OAI211_X1 U16776 ( .C1(n8859), .C2(n15622), .A(n15556), .B(n15555), .ZN(
        P1_U3214) );
  INV_X1 U16777 ( .A(n15557), .ZN(n15558) );
  AOI21_X1 U16778 ( .B1(n15560), .B2(n15559), .A(n15558), .ZN(n15564) );
  OAI22_X1 U16779 ( .A1(n15778), .A2(n15953), .B1(n15761), .B2(n15951), .ZN(
        n16039) );
  AOI22_X1 U16780 ( .A1(n16530), .A2(n16039), .B1(P1_REG3_REG_23__SCAN_IN), 
        .B2(P1_U3086), .ZN(n15561) );
  OAI21_X1 U16781 ( .B1(n15878), .B2(n16535), .A(n15561), .ZN(n15562) );
  AOI21_X1 U16782 ( .B1(n16040), .B2(n15671), .A(n15562), .ZN(n15563) );
  OAI21_X1 U16783 ( .B1(n15564), .B2(n15673), .A(n15563), .ZN(P1_U3216) );
  NAND2_X1 U16784 ( .A1(n15566), .A2(n15565), .ZN(n15567) );
  XNOR2_X1 U16785 ( .A(n15568), .B(n15567), .ZN(n15573) );
  NAND2_X1 U16786 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n15736)
         );
  OAI21_X1 U16787 ( .B1(n15648), .B2(n15939), .A(n15736), .ZN(n15569) );
  AOI21_X1 U16788 ( .B1(n15659), .B2(n15973), .A(n15569), .ZN(n15570) );
  OAI21_X1 U16789 ( .B1(n15940), .B2(n16535), .A(n15570), .ZN(n15571) );
  AOI21_X1 U16790 ( .B1(n16068), .B2(n15671), .A(n15571), .ZN(n15572) );
  OAI21_X1 U16791 ( .B1(n15573), .B2(n15673), .A(n15572), .ZN(P1_U3219) );
  INV_X1 U16792 ( .A(n15574), .ZN(n15575) );
  AOI21_X1 U16793 ( .B1(n15577), .B2(n15576), .A(n15575), .ZN(n15583) );
  NOR2_X1 U16794 ( .A1(n15761), .A2(n15953), .ZN(n15578) );
  AOI21_X1 U16795 ( .B1(n15759), .B2(n15971), .A(n15578), .ZN(n16051) );
  INV_X1 U16796 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n15579) );
  OAI22_X1 U16797 ( .A1(n16051), .A2(n15638), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15579), .ZN(n15581) );
  NOR2_X1 U16798 ( .A1(n16053), .A2(n15653), .ZN(n15580) );
  AOI211_X1 U16799 ( .C1(n15640), .C2(n15905), .A(n15581), .B(n15580), .ZN(
        n15582) );
  OAI21_X1 U16800 ( .B1(n15583), .B2(n15673), .A(n15582), .ZN(P1_U3223) );
  XOR2_X1 U16801 ( .A(n15585), .B(n15584), .Z(n15591) );
  NAND2_X1 U16802 ( .A1(n15675), .A2(n15971), .ZN(n15587) );
  NAND2_X1 U16803 ( .A1(n15765), .A2(n16462), .ZN(n15586) );
  NAND2_X1 U16804 ( .A1(n15587), .A2(n15586), .ZN(n15849) );
  AOI22_X1 U16805 ( .A1(n16530), .A2(n15849), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3086), .ZN(n15588) );
  OAI21_X1 U16806 ( .B1(n15850), .B2(n16535), .A(n15588), .ZN(n15589) );
  AOI21_X1 U16807 ( .B1(n15738), .B2(n15671), .A(n15589), .ZN(n15590) );
  OAI21_X1 U16808 ( .B1(n15591), .B2(n15673), .A(n15590), .ZN(P1_U3225) );
  INV_X1 U16809 ( .A(n15593), .ZN(n15594) );
  AOI21_X1 U16810 ( .B1(n15595), .B2(n15592), .A(n15594), .ZN(n15602) );
  INV_X1 U16811 ( .A(n15755), .ZN(n15952) );
  OAI21_X1 U16812 ( .B1(n15648), .B2(n15952), .A(n15596), .ZN(n15597) );
  AOI21_X1 U16813 ( .B1(n15659), .B2(n15678), .A(n15597), .ZN(n15598) );
  OAI21_X1 U16814 ( .B1(n15599), .B2(n16535), .A(n15598), .ZN(n15600) );
  AOI21_X1 U16815 ( .B1(n16085), .B2(n15671), .A(n15600), .ZN(n15601) );
  OAI21_X1 U16816 ( .B1(n15602), .B2(n15673), .A(n15601), .ZN(P1_U3226) );
  OAI21_X1 U16817 ( .B1(n15605), .B2(n15604), .A(n15603), .ZN(n15606) );
  NAND2_X1 U16818 ( .A1(n15606), .A2(n16531), .ZN(n15611) );
  NOR2_X1 U16819 ( .A1(n16535), .A2(n15978), .ZN(n15609) );
  OAI21_X1 U16820 ( .B1(n15648), .B2(n15938), .A(n15607), .ZN(n15608) );
  AOI211_X1 U16821 ( .C1(n15659), .C2(n15972), .A(n15609), .B(n15608), .ZN(
        n15610) );
  OAI211_X1 U16822 ( .C1(n8309), .C2(n15653), .A(n15611), .B(n15610), .ZN(
        P1_U3228) );
  NAND2_X1 U16823 ( .A1(n15869), .A2(n16606), .ZN(n16032) );
  OAI21_X1 U16824 ( .B1(n15614), .B2(n15613), .A(n15612), .ZN(n15615) );
  NAND2_X1 U16825 ( .A1(n15615), .A2(n16531), .ZN(n15621) );
  NOR2_X1 U16826 ( .A1(n16535), .A2(n15867), .ZN(n15619) );
  INV_X1 U16827 ( .A(n15859), .ZN(n15617) );
  INV_X1 U16828 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n15616) );
  OAI22_X1 U16829 ( .A1(n15648), .A2(n15617), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15616), .ZN(n15618) );
  AOI211_X1 U16830 ( .C1(n15659), .C2(n15860), .A(n15619), .B(n15618), .ZN(
        n15620) );
  OAI211_X1 U16831 ( .C1(n15622), .C2(n16032), .A(n15621), .B(n15620), .ZN(
        P1_U3229) );
  NAND2_X1 U16832 ( .A1(n15676), .A2(n16462), .ZN(n15624) );
  NAND2_X1 U16833 ( .A1(n15756), .A2(n15971), .ZN(n15623) );
  NAND2_X1 U16834 ( .A1(n15624), .A2(n15623), .ZN(n16058) );
  AOI22_X1 U16835 ( .A1(n16530), .A2(n16058), .B1(P1_REG3_REG_20__SCAN_IN), 
        .B2(P1_U3086), .ZN(n15625) );
  OAI21_X1 U16836 ( .B1(n15919), .B2(n16535), .A(n15625), .ZN(n15630) );
  AOI211_X1 U16837 ( .C1(n15628), .C2(n15627), .A(n15673), .B(n7786), .ZN(
        n15629) );
  AOI211_X1 U16838 ( .C1(n15671), .C2(n16059), .A(n15630), .B(n15629), .ZN(
        n15631) );
  INV_X1 U16839 ( .A(n15631), .ZN(P1_U3233) );
  AOI21_X1 U16840 ( .B1(n15633), .B2(n15632), .A(n15673), .ZN(n15635) );
  NAND2_X1 U16841 ( .A1(n15635), .A2(n15634), .ZN(n15643) );
  INV_X1 U16842 ( .A(n15895), .ZN(n15641) );
  AND2_X1 U16843 ( .A1(n15860), .A2(n16462), .ZN(n15636) );
  AOI21_X1 U16844 ( .B1(n15676), .B2(n15971), .A(n15636), .ZN(n16044) );
  INV_X1 U16845 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n15637) );
  OAI22_X1 U16846 ( .A1(n16044), .A2(n15638), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15637), .ZN(n15639) );
  AOI21_X1 U16847 ( .B1(n15641), .B2(n15640), .A(n15639), .ZN(n15642) );
  OAI211_X1 U16848 ( .C1(n15653), .C2(n16046), .A(n15643), .B(n15642), .ZN(
        P1_U3235) );
  INV_X1 U16849 ( .A(n16074), .ZN(n15962) );
  OAI21_X1 U16850 ( .B1(n15646), .B2(n15645), .A(n15644), .ZN(n15647) );
  NAND2_X1 U16851 ( .A1(n15647), .A2(n16531), .ZN(n15652) );
  NOR2_X1 U16852 ( .A1(n16535), .A2(n15963), .ZN(n15650) );
  NAND2_X1 U16853 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n15706)
         );
  OAI21_X1 U16854 ( .B1(n15648), .B2(n15954), .A(n15706), .ZN(n15649) );
  AOI211_X1 U16855 ( .C1(n15659), .C2(n15755), .A(n15650), .B(n15649), .ZN(
        n15651) );
  OAI211_X1 U16856 ( .C1(n15962), .C2(n15653), .A(n15652), .B(n15651), .ZN(
        P1_U3238) );
  NAND2_X1 U16857 ( .A1(n15656), .A2(n15655), .ZN(n15657) );
  XNOR2_X1 U16858 ( .A(n15654), .B(n15657), .ZN(n15664) );
  AOI22_X1 U16859 ( .A1(n15658), .A2(n15838), .B1(P1_REG3_REG_26__SCAN_IN), 
        .B2(P1_U3086), .ZN(n15661) );
  NAND2_X1 U16860 ( .A1(n15659), .A2(n15859), .ZN(n15660) );
  OAI211_X1 U16861 ( .C1(n16535), .C2(n15831), .A(n15661), .B(n15660), .ZN(
        n15662) );
  AOI21_X1 U16862 ( .B1(n16021), .B2(n15671), .A(n15662), .ZN(n15663) );
  OAI21_X1 U16863 ( .B1(n15664), .B2(n15673), .A(n15663), .ZN(P1_U3240) );
  XNOR2_X1 U16864 ( .A(n15666), .B(n15665), .ZN(n15674) );
  NAND2_X1 U16865 ( .A1(n16530), .A2(n16089), .ZN(n15667) );
  OAI211_X1 U16866 ( .C1(n16535), .C2(n15669), .A(n15668), .B(n15667), .ZN(
        n15670) );
  AOI21_X1 U16867 ( .B1(n16090), .B2(n15671), .A(n15670), .ZN(n15672) );
  OAI21_X1 U16868 ( .B1(n15674), .B2(n15673), .A(n15672), .ZN(P1_U3241) );
  MUX2_X1 U16869 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n15788), .S(P1_U4016), .Z(
        P1_U3590) );
  MUX2_X1 U16870 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n15800), .S(P1_U4016), .Z(
        P1_U3589) );
  MUX2_X1 U16871 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n15791), .S(P1_U4016), .Z(
        P1_U3588) );
  MUX2_X1 U16872 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n15765), .S(P1_U4016), .Z(
        P1_U3586) );
  MUX2_X1 U16873 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n15859), .S(P1_U4016), .Z(
        P1_U3585) );
  MUX2_X1 U16874 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n15675), .S(P1_U4016), .Z(
        P1_U3584) );
  MUX2_X1 U16875 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n15860), .S(P1_U4016), .Z(
        P1_U3583) );
  INV_X1 U16876 ( .A(n15761), .ZN(n15775) );
  MUX2_X1 U16877 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n15775), .S(P1_U4016), .Z(
        P1_U3582) );
  MUX2_X1 U16878 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n15676), .S(P1_U4016), .Z(
        P1_U3581) );
  MUX2_X1 U16879 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n15759), .S(P1_U4016), .Z(
        P1_U3580) );
  MUX2_X1 U16880 ( .A(n15756), .B(P1_DATAO_REG_19__SCAN_IN), .S(n15677), .Z(
        P1_U3579) );
  MUX2_X1 U16881 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n15973), .S(P1_U4016), .Z(
        P1_U3578) );
  MUX2_X1 U16882 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n15755), .S(P1_U4016), .Z(
        P1_U3577) );
  MUX2_X1 U16883 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n15972), .S(P1_U4016), .Z(
        P1_U3576) );
  MUX2_X1 U16884 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n15678), .S(P1_U4016), .Z(
        P1_U3575) );
  MUX2_X1 U16885 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n15679), .S(P1_U4016), .Z(
        P1_U3574) );
  MUX2_X1 U16886 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n15680), .S(P1_U4016), .Z(
        P1_U3573) );
  MUX2_X1 U16887 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n15681), .S(P1_U4016), .Z(
        P1_U3572) );
  MUX2_X1 U16888 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n15682), .S(P1_U4016), .Z(
        P1_U3571) );
  MUX2_X1 U16889 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n15683), .S(P1_U4016), .Z(
        P1_U3570) );
  MUX2_X1 U16890 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n15684), .S(P1_U4016), .Z(
        P1_U3569) );
  MUX2_X1 U16891 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n15685), .S(P1_U4016), .Z(
        P1_U3568) );
  MUX2_X1 U16892 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n15686), .S(P1_U4016), .Z(
        P1_U3567) );
  MUX2_X1 U16893 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n15687), .S(P1_U4016), .Z(
        P1_U3566) );
  MUX2_X1 U16894 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n15688), .S(P1_U4016), .Z(
        P1_U3565) );
  MUX2_X1 U16895 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n15689), .S(P1_U4016), .Z(
        P1_U3564) );
  MUX2_X1 U16896 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n15690), .S(P1_U4016), .Z(
        P1_U3563) );
  MUX2_X1 U16897 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n16463), .S(P1_U4016), .Z(
        P1_U3562) );
  MUX2_X1 U16898 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n10430), .S(P1_U4016), .Z(
        P1_U3561) );
  MUX2_X1 U16899 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n15691), .S(P1_U4016), .Z(
        P1_U3560) );
  OAI211_X1 U16900 ( .C1(n15694), .C2(n15693), .A(n16263), .B(n15692), .ZN(
        n15702) );
  OAI211_X1 U16901 ( .C1(n15697), .C2(n15696), .A(n16259), .B(n15695), .ZN(
        n15701) );
  AOI22_X1 U16902 ( .A1(n16246), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n15700) );
  NAND2_X1 U16903 ( .A1(n16261), .A2(n15698), .ZN(n15699) );
  NAND4_X1 U16904 ( .A1(n15702), .A2(n15701), .A3(n15700), .A4(n15699), .ZN(
        P1_U3244) );
  NAND2_X1 U16905 ( .A1(n15709), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n15704) );
  NAND2_X1 U16906 ( .A1(n15704), .A2(n15703), .ZN(n15722) );
  XNOR2_X1 U16907 ( .A(n15722), .B(n15717), .ZN(n15705) );
  NAND2_X1 U16908 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n15705), .ZN(n15724) );
  OAI211_X1 U16909 ( .C1(n15705), .C2(P1_REG2_REG_18__SCAN_IN), .A(n16263), 
        .B(n15724), .ZN(n15716) );
  INV_X1 U16910 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n15707) );
  OAI21_X1 U16911 ( .B1(n16267), .B2(n15707), .A(n15706), .ZN(n15714) );
  NOR2_X1 U16912 ( .A1(n15711), .A2(n15712), .ZN(n15720) );
  AOI211_X1 U16913 ( .C1(n15712), .C2(n15711), .A(n15720), .B(n15710), .ZN(
        n15713) );
  AOI211_X1 U16914 ( .C1(n16261), .C2(n15723), .A(n15714), .B(n15713), .ZN(
        n15715) );
  NAND2_X1 U16915 ( .A1(n15716), .A2(n15715), .ZN(P1_U3261) );
  NOR2_X1 U16916 ( .A1(n15718), .A2(n15717), .ZN(n15719) );
  NOR2_X1 U16917 ( .A1(n15720), .A2(n15719), .ZN(n15721) );
  XNOR2_X1 U16918 ( .A(n15721), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n15732) );
  INV_X1 U16919 ( .A(n15732), .ZN(n15730) );
  NAND2_X1 U16920 ( .A1(n15723), .A2(n15722), .ZN(n15725) );
  NAND2_X1 U16921 ( .A1(n15725), .A2(n15724), .ZN(n15726) );
  XOR2_X1 U16922 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n15726), .Z(n15731) );
  OAI21_X1 U16923 ( .B1(n15731), .B2(n15728), .A(n15727), .ZN(n15729) );
  AOI21_X1 U16924 ( .B1(n15730), .B2(n16259), .A(n15729), .ZN(n15735) );
  AOI22_X1 U16925 ( .A1(n15732), .A2(n16259), .B1(n16263), .B2(n15731), .ZN(
        n15734) );
  OAI211_X1 U16926 ( .C1(n8926), .C2(n16267), .A(n15737), .B(n15736), .ZN(
        P1_U3262) );
  NAND2_X1 U16927 ( .A1(n16002), .A2(n15785), .ZN(n15746) );
  OR2_X1 U16928 ( .A1(n7417), .A2(n15739), .ZN(n15740) );
  AND2_X1 U16929 ( .A1(n16462), .A2(n15740), .ZN(n15787) );
  INV_X1 U16930 ( .A(n15787), .ZN(n15741) );
  OR2_X1 U16931 ( .A1(n15742), .A2(n15741), .ZN(n16000) );
  NOR2_X1 U16932 ( .A1(n7414), .A2(n16000), .ZN(n15747) );
  NOR2_X1 U16933 ( .A1(n8074), .A2(n16481), .ZN(n15744) );
  AOI211_X1 U16934 ( .C1(n7414), .C2(P1_REG2_REG_31__SCAN_IN), .A(n15747), .B(
        n15744), .ZN(n15745) );
  OAI21_X1 U16935 ( .B1(n16631), .B2(n15999), .A(n15745), .ZN(P1_U3263) );
  OAI211_X1 U16936 ( .C1(n15785), .C2(n16002), .A(n15746), .B(n16079), .ZN(
        n16001) );
  NAND2_X1 U16937 ( .A1(n7414), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n15749) );
  INV_X1 U16938 ( .A(n15747), .ZN(n15748) );
  OAI211_X1 U16939 ( .C1(n16002), .C2(n16481), .A(n15749), .B(n15748), .ZN(
        n15750) );
  INV_X1 U16940 ( .A(n15750), .ZN(n15751) );
  OAI21_X1 U16941 ( .B1(n16001), .B2(n16631), .A(n15751), .ZN(P1_U3264) );
  OR2_X1 U16942 ( .A1(n16085), .A2(n15972), .ZN(n15752) );
  INV_X1 U16943 ( .A(n16003), .ZN(n15798) );
  NAND2_X1 U16944 ( .A1(n15970), .A2(n15981), .ZN(n15969) );
  NAND2_X1 U16945 ( .A1(n16078), .A2(n15952), .ZN(n15768) );
  NAND2_X1 U16946 ( .A1(n15969), .A2(n15768), .ZN(n15957) );
  OR2_X1 U16947 ( .A1(n16074), .A2(n15938), .ZN(n15769) );
  NAND2_X1 U16948 ( .A1(n16068), .A2(n15954), .ZN(n15770) );
  NOR2_X1 U16949 ( .A1(n15906), .A2(n15772), .ZN(n15773) );
  NOR2_X1 U16950 ( .A1(n16046), .A2(n15775), .ZN(n15776) );
  NOR2_X1 U16951 ( .A1(n16027), .A2(n15859), .ZN(n15835) );
  INV_X1 U16952 ( .A(n15781), .ZN(n15782) );
  XNOR2_X1 U16953 ( .A(n15784), .B(n15783), .ZN(n16009) );
  INV_X1 U16954 ( .A(n15786), .ZN(n16006) );
  AOI211_X1 U16955 ( .C1(n15786), .C2(n7497), .A(n16464), .B(n15785), .ZN(
        n16008) );
  NAND2_X1 U16956 ( .A1(n16008), .A2(n16486), .ZN(n15795) );
  NAND2_X1 U16957 ( .A1(n15788), .A2(n15787), .ZN(n16004) );
  OAI22_X1 U16958 ( .A1(n15790), .A2(n16004), .B1(n15789), .B2(n16622), .ZN(
        n15793) );
  NAND2_X1 U16959 ( .A1(n15791), .A2(n15971), .ZN(n16005) );
  NOR2_X1 U16960 ( .A1(n7414), .A2(n16005), .ZN(n15792) );
  AOI211_X1 U16961 ( .C1(n7414), .C2(P1_REG2_REG_29__SCAN_IN), .A(n15793), .B(
        n15792), .ZN(n15794) );
  OAI211_X1 U16962 ( .C1(n16006), .C2(n16481), .A(n15795), .B(n15794), .ZN(
        n15796) );
  AOI21_X1 U16963 ( .B1(n16009), .B2(n15855), .A(n15796), .ZN(n15797) );
  OAI21_X1 U16964 ( .B1(n15798), .B2(n15983), .A(n15797), .ZN(P1_U3356) );
  AOI21_X1 U16965 ( .B1(n15804), .B2(n15803), .A(n15802), .ZN(n16010) );
  OAI211_X1 U16966 ( .C1(n15818), .C2(n15808), .A(n16079), .B(n7497), .ZN(
        n16013) );
  NOR2_X1 U16967 ( .A1(n16013), .A2(n16631), .ZN(n15810) );
  NOR2_X1 U16968 ( .A1(n16622), .A2(n15805), .ZN(n15806) );
  AOI21_X1 U16969 ( .B1(n7414), .B2(P1_REG2_REG_28__SCAN_IN), .A(n15806), .ZN(
        n15807) );
  OAI21_X1 U16970 ( .B1(n15808), .B2(n16481), .A(n15807), .ZN(n15809) );
  AOI211_X1 U16971 ( .C1(n16010), .C2(n15935), .A(n15810), .B(n15809), .ZN(
        n15811) );
  OAI21_X1 U16972 ( .B1(n16014), .B2(n7414), .A(n15811), .ZN(P1_U3265) );
  OAI22_X1 U16973 ( .A1(n15816), .A2(n15951), .B1(n15815), .B2(n15953), .ZN(
        n15817) );
  NAND2_X1 U16974 ( .A1(n16015), .A2(n16625), .ZN(n15825) );
  AOI211_X1 U16975 ( .C1(n15819), .C2(n15830), .A(n16464), .B(n15818), .ZN(
        n16016) );
  NOR2_X1 U16976 ( .A1(n8618), .A2(n16481), .ZN(n15823) );
  OAI22_X1 U16977 ( .A1(n16625), .A2(n15821), .B1(n15820), .B2(n16622), .ZN(
        n15822) );
  AOI211_X1 U16978 ( .C1(n16016), .C2(n16486), .A(n15823), .B(n15822), .ZN(
        n15824) );
  OAI211_X1 U16979 ( .C1(n15827), .C2(n15826), .A(n15825), .B(n15824), .ZN(
        P1_U3266) );
  XNOR2_X1 U16980 ( .A(n15829), .B(n15828), .ZN(n16024) );
  AOI211_X1 U16981 ( .C1(n16021), .C2(n15848), .A(n16464), .B(n8307), .ZN(
        n16020) );
  INV_X1 U16982 ( .A(n16021), .ZN(n15834) );
  INV_X1 U16983 ( .A(n15831), .ZN(n15832) );
  AOI22_X1 U16984 ( .A1(n7414), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n15832), 
        .B2(n15991), .ZN(n15833) );
  OAI21_X1 U16985 ( .B1(n15834), .B2(n16481), .A(n15833), .ZN(n15840) );
  OR3_X1 U16986 ( .A1(n15845), .A2(n8615), .A3(n15835), .ZN(n15836) );
  NOR2_X1 U16987 ( .A1(n16023), .A2(n7414), .ZN(n15839) );
  AOI211_X1 U16988 ( .C1(n16020), .C2(n16486), .A(n15840), .B(n15839), .ZN(
        n15841) );
  OAI21_X1 U16989 ( .B1(n16024), .B2(n15983), .A(n15841), .ZN(P1_U3267) );
  OAI21_X1 U16990 ( .B1(n15844), .B2(n15843), .A(n15842), .ZN(n16031) );
  INV_X1 U16991 ( .A(n15845), .ZN(n15846) );
  OAI21_X1 U16992 ( .B1(n7518), .B2(n15847), .A(n15846), .ZN(n16029) );
  OAI211_X1 U16993 ( .C1(n15864), .C2(n16027), .A(n15848), .B(n16079), .ZN(
        n16026) );
  INV_X1 U16994 ( .A(n15849), .ZN(n16025) );
  OAI22_X1 U16995 ( .A1(n7414), .A2(n16025), .B1(n15850), .B2(n16622), .ZN(
        n15852) );
  NOR2_X1 U16996 ( .A1(n16027), .A2(n16481), .ZN(n15851) );
  AOI211_X1 U16997 ( .C1(n7414), .C2(P1_REG2_REG_25__SCAN_IN), .A(n15852), .B(
        n15851), .ZN(n15853) );
  OAI21_X1 U16998 ( .B1(n16631), .B2(n16026), .A(n15853), .ZN(n15854) );
  AOI21_X1 U16999 ( .B1(n16029), .B2(n15855), .A(n15854), .ZN(n15856) );
  OAI21_X1 U17000 ( .B1(n16031), .B2(n15983), .A(n15856), .ZN(P1_U3268) );
  OAI211_X1 U17001 ( .C1(n15858), .C2(n15872), .A(n15857), .B(n16561), .ZN(
        n15862) );
  AOI22_X1 U17002 ( .A1(n15971), .A2(n15860), .B1(n15859), .B2(n16462), .ZN(
        n15861) );
  NAND2_X1 U17003 ( .A1(n15862), .A2(n15861), .ZN(n16035) );
  NAND2_X1 U17004 ( .A1(n15877), .A2(n15869), .ZN(n15863) );
  NAND2_X1 U17005 ( .A1(n15863), .A2(n16079), .ZN(n15865) );
  OR2_X1 U17006 ( .A1(n15865), .A2(n15864), .ZN(n16033) );
  NAND2_X1 U17007 ( .A1(n7414), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n15866) );
  OAI21_X1 U17008 ( .B1(n16622), .B2(n15867), .A(n15866), .ZN(n15868) );
  AOI21_X1 U17009 ( .B1(n15869), .B2(n16628), .A(n15868), .ZN(n15870) );
  OAI21_X1 U17010 ( .B1(n16033), .B2(n16631), .A(n15870), .ZN(n15874) );
  AOI21_X1 U17011 ( .B1(n15872), .B2(n15871), .A(n7534), .ZN(n16034) );
  NOR2_X1 U17012 ( .A1(n16034), .A2(n15983), .ZN(n15873) );
  AOI211_X1 U17013 ( .C1(n16625), .C2(n16035), .A(n15874), .B(n15873), .ZN(
        n15875) );
  INV_X1 U17014 ( .A(n15875), .ZN(P1_U3269) );
  OAI21_X1 U17015 ( .B1(n7466), .B2(n15884), .A(n15876), .ZN(n16037) );
  INV_X1 U17016 ( .A(n16039), .ZN(n15879) );
  OAI22_X1 U17017 ( .A1(n7414), .A2(n15879), .B1(n15878), .B2(n16622), .ZN(
        n15880) );
  AOI21_X1 U17018 ( .B1(P1_REG2_REG_23__SCAN_IN), .B2(n7414), .A(n15880), .ZN(
        n15881) );
  OAI21_X1 U17019 ( .B1(n15882), .B2(n16481), .A(n15881), .ZN(n15887) );
  AOI21_X1 U17020 ( .B1(n15885), .B2(n15884), .A(n15883), .ZN(n16043) );
  NOR2_X1 U17021 ( .A1(n16043), .A2(n15947), .ZN(n15886) );
  AOI211_X1 U17022 ( .C1(n16038), .C2(n16486), .A(n15887), .B(n15886), .ZN(
        n15888) );
  OAI21_X1 U17023 ( .B1(n16037), .B2(n15983), .A(n15888), .ZN(P1_U3270) );
  XOR2_X1 U17024 ( .A(n15891), .B(n15889), .Z(n16050) );
  AOI21_X1 U17025 ( .B1(n15892), .B2(n15891), .A(n15890), .ZN(n15893) );
  INV_X1 U17026 ( .A(n15893), .ZN(n16048) );
  OAI211_X1 U17027 ( .C1(n16046), .C2(n15904), .A(n16079), .B(n15894), .ZN(
        n16045) );
  OAI21_X1 U17028 ( .B1(n15895), .B2(n16622), .A(n16044), .ZN(n15896) );
  MUX2_X1 U17029 ( .A(n15896), .B(P1_REG2_REG_22__SCAN_IN), .S(n7414), .Z(
        n15897) );
  AOI21_X1 U17030 ( .B1(n7726), .B2(n16628), .A(n15897), .ZN(n15898) );
  OAI21_X1 U17031 ( .B1(n16045), .B2(n16631), .A(n15898), .ZN(n15899) );
  AOI21_X1 U17032 ( .B1(n16048), .B2(n15935), .A(n15899), .ZN(n15900) );
  OAI21_X1 U17033 ( .B1(n16050), .B2(n15947), .A(n15900), .ZN(P1_U3271) );
  XNOR2_X1 U17034 ( .A(n15901), .B(n15910), .ZN(n16056) );
  NAND2_X1 U17035 ( .A1(n15906), .A2(n15921), .ZN(n15902) );
  NAND2_X1 U17036 ( .A1(n15902), .A2(n16079), .ZN(n15903) );
  OR2_X1 U17037 ( .A1(n15904), .A2(n15903), .ZN(n16052) );
  AOI22_X1 U17038 ( .A1(n7414), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n15905), 
        .B2(n15991), .ZN(n15908) );
  NAND2_X1 U17039 ( .A1(n15906), .A2(n16628), .ZN(n15907) );
  OAI211_X1 U17040 ( .C1(n16052), .C2(n16631), .A(n15908), .B(n15907), .ZN(
        n15909) );
  AOI21_X1 U17041 ( .B1(n16056), .B2(n15935), .A(n15909), .ZN(n15915) );
  XNOR2_X1 U17042 ( .A(n15911), .B(n15910), .ZN(n15912) );
  AND2_X1 U17043 ( .A1(n15912), .A2(n16561), .ZN(n16055) );
  INV_X1 U17044 ( .A(n16051), .ZN(n15913) );
  OAI21_X1 U17045 ( .B1(n16055), .B2(n15913), .A(n16625), .ZN(n15914) );
  NAND2_X1 U17046 ( .A1(n15915), .A2(n15914), .ZN(P1_U3272) );
  NOR2_X1 U17047 ( .A1(n15916), .A2(n15925), .ZN(n15917) );
  INV_X1 U17048 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n15920) );
  OAI22_X1 U17049 ( .A1(n16625), .A2(n15920), .B1(n15919), .B2(n16622), .ZN(
        n15924) );
  AOI21_X1 U17050 ( .B1(n16059), .B2(n15936), .A(n16464), .ZN(n15922) );
  NAND2_X1 U17051 ( .A1(n15922), .A2(n15921), .ZN(n16060) );
  NOR2_X1 U17052 ( .A1(n16060), .A2(n16631), .ZN(n15923) );
  AOI211_X1 U17053 ( .C1(n16628), .C2(n16059), .A(n15924), .B(n15923), .ZN(
        n15931) );
  NAND2_X1 U17054 ( .A1(n15926), .A2(n15925), .ZN(n15927) );
  NAND3_X1 U17055 ( .A1(n15928), .A2(n16561), .A3(n15927), .ZN(n16062) );
  INV_X1 U17056 ( .A(n16062), .ZN(n15929) );
  OAI21_X1 U17057 ( .B1(n15929), .B2(n16058), .A(n16625), .ZN(n15930) );
  OAI211_X1 U17058 ( .C1(n16064), .C2(n15983), .A(n15931), .B(n15930), .ZN(
        P1_U3273) );
  XOR2_X1 U17059 ( .A(n15933), .B(n15932), .Z(n16071) );
  XNOR2_X1 U17060 ( .A(n15934), .B(n15933), .ZN(n16065) );
  NAND2_X1 U17061 ( .A1(n16065), .A2(n15935), .ZN(n15946) );
  INV_X1 U17062 ( .A(n15936), .ZN(n15937) );
  AOI211_X1 U17063 ( .C1(n16068), .C2(n15961), .A(n16464), .B(n15937), .ZN(
        n16066) );
  OAI22_X1 U17064 ( .A1(n15939), .A2(n15953), .B1(n15938), .B2(n15951), .ZN(
        n16067) );
  INV_X1 U17065 ( .A(n15940), .ZN(n15941) );
  AOI22_X1 U17066 ( .A1(n16067), .A2(n16625), .B1(n15941), .B2(n15991), .ZN(
        n15943) );
  NAND2_X1 U17067 ( .A1(n7414), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n15942) );
  OAI211_X1 U17068 ( .C1(n8311), .C2(n16481), .A(n15943), .B(n15942), .ZN(
        n15944) );
  AOI21_X1 U17069 ( .B1(n16066), .B2(n16486), .A(n15944), .ZN(n15945) );
  OAI211_X1 U17070 ( .C1(n16071), .C2(n15947), .A(n15946), .B(n15945), .ZN(
        P1_U3274) );
  INV_X1 U17071 ( .A(n15948), .ZN(n15950) );
  OAI21_X1 U17072 ( .B1(n15950), .B2(n15958), .A(n15949), .ZN(n16072) );
  OAI22_X1 U17073 ( .A1(n15954), .A2(n15953), .B1(n15952), .B2(n15951), .ZN(
        n15960) );
  AOI211_X1 U17074 ( .C1(n15958), .C2(n15957), .A(n16726), .B(n15956), .ZN(
        n15959) );
  AOI211_X1 U17075 ( .C1(n16072), .C2(n16472), .A(n15960), .B(n15959), .ZN(
        n16076) );
  AOI211_X1 U17076 ( .C1(n16074), .C2(n15975), .A(n16464), .B(n8308), .ZN(
        n16073) );
  NOR2_X1 U17077 ( .A1(n15962), .A2(n16481), .ZN(n15966) );
  OAI22_X1 U17078 ( .A1(n16625), .A2(n15964), .B1(n15963), .B2(n16622), .ZN(
        n15965) );
  AOI211_X1 U17079 ( .C1(n16073), .C2(n16486), .A(n15966), .B(n15965), .ZN(
        n15968) );
  NAND2_X1 U17080 ( .A1(n16072), .A2(n16633), .ZN(n15967) );
  OAI211_X1 U17081 ( .C1(n16076), .C2(n7414), .A(n15968), .B(n15967), .ZN(
        P1_U3275) );
  OAI21_X1 U17082 ( .B1(n15970), .B2(n15981), .A(n15969), .ZN(n15974) );
  AOI222_X1 U17083 ( .A1(n16561), .A2(n15974), .B1(n15973), .B2(n16462), .C1(
        n15972), .C2(n15971), .ZN(n16082) );
  INV_X1 U17084 ( .A(n15975), .ZN(n15976) );
  AOI21_X1 U17085 ( .B1(n16078), .B2(n15977), .A(n15976), .ZN(n16080) );
  INV_X1 U17086 ( .A(n15978), .ZN(n15979) );
  AOI22_X1 U17087 ( .A1(n7414), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n15979), 
        .B2(n15991), .ZN(n15980) );
  OAI21_X1 U17088 ( .B1(n8309), .B2(n16481), .A(n15980), .ZN(n15985) );
  OAI21_X1 U17089 ( .B1(n7611), .B2(n15754), .A(n15982), .ZN(n16083) );
  NOR2_X1 U17090 ( .A1(n16083), .A2(n15983), .ZN(n15984) );
  AOI211_X1 U17091 ( .C1(n16080), .C2(n15986), .A(n15985), .B(n15984), .ZN(
        n15987) );
  OAI21_X1 U17092 ( .B1(n7414), .B2(n16082), .A(n15987), .ZN(P1_U3276) );
  INV_X1 U17093 ( .A(n15992), .ZN(n16445) );
  AOI22_X1 U17094 ( .A1(n16465), .A2(n16628), .B1(n16633), .B2(n16445), .ZN(
        n15998) );
  NAND2_X1 U17095 ( .A1(n10384), .A2(n15988), .ZN(n15989) );
  NOR2_X1 U17096 ( .A1(n15990), .A2(n15989), .ZN(n16444) );
  AOI22_X1 U17097 ( .A1(n16486), .A2(n16444), .B1(P1_REG3_REG_0__SCAN_IN), 
        .B2(n15991), .ZN(n15997) );
  AOI21_X1 U17098 ( .B1(n16726), .B2(n15993), .A(n15992), .ZN(n15994) );
  AOI21_X1 U17099 ( .B1(n16462), .B2(n10430), .A(n15994), .ZN(n16442) );
  NOR2_X1 U17100 ( .A1(n7414), .A2(n16442), .ZN(n15995) );
  AOI21_X1 U17101 ( .B1(n7414), .B2(P1_REG2_REG_0__SCAN_IN), .A(n15995), .ZN(
        n15996) );
  NAND3_X1 U17102 ( .A1(n15998), .A2(n15997), .A3(n15996), .ZN(P1_U3293) );
  MUX2_X1 U17103 ( .A(n16097), .B(P1_REG1_REG_31__SCAN_IN), .S(n16732), .Z(
        P1_U3559) );
  OAI211_X1 U17104 ( .C1(n16725), .C2(n16002), .A(n16001), .B(n16000), .ZN(
        n16098) );
  MUX2_X1 U17105 ( .A(n16098), .B(P1_REG1_REG_30__SCAN_IN), .S(n16732), .Z(
        P1_U3558) );
  OAI211_X1 U17106 ( .C1(n16006), .C2(n16725), .A(n16005), .B(n16004), .ZN(
        n16007) );
  MUX2_X1 U17107 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n16099), .S(n16734), .Z(
        P1_U3557) );
  NAND2_X1 U17108 ( .A1(n16011), .A2(n16606), .ZN(n16012) );
  MUX2_X1 U17109 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n16100), .S(n16734), .Z(
        P1_U3556) );
  INV_X1 U17110 ( .A(n16015), .ZN(n16019) );
  INV_X1 U17111 ( .A(n16016), .ZN(n16018) );
  MUX2_X1 U17112 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n16101), .S(n16734), .Z(
        P1_U3555) );
  AOI21_X1 U17113 ( .B1(n16021), .B2(n16606), .A(n16020), .ZN(n16022) );
  OAI211_X1 U17114 ( .C1(n16024), .C2(n16540), .A(n16023), .B(n16022), .ZN(
        n16102) );
  MUX2_X1 U17115 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n16102), .S(n16734), .Z(
        P1_U3554) );
  OAI211_X1 U17116 ( .C1(n16027), .C2(n16725), .A(n16026), .B(n16025), .ZN(
        n16028) );
  AOI21_X1 U17117 ( .B1(n16029), .B2(n16561), .A(n16028), .ZN(n16030) );
  OAI21_X1 U17118 ( .B1(n16031), .B2(n16540), .A(n16030), .ZN(n16103) );
  MUX2_X1 U17119 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n16103), .S(n16734), .Z(
        P1_U3553) );
  OAI211_X1 U17120 ( .C1(n16034), .C2(n16540), .A(n16033), .B(n16032), .ZN(
        n16036) );
  MUX2_X1 U17121 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n16104), .S(n16734), .Z(
        P1_U3552) );
  OR2_X1 U17122 ( .A1(n16037), .A2(n16540), .ZN(n16042) );
  OAI211_X1 U17123 ( .C1(n16726), .C2(n16043), .A(n16042), .B(n16041), .ZN(
        n16105) );
  MUX2_X1 U17124 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n16105), .S(n16734), .Z(
        P1_U3551) );
  OAI211_X1 U17125 ( .C1(n16725), .C2(n16046), .A(n16045), .B(n16044), .ZN(
        n16047) );
  AOI21_X1 U17126 ( .B1(n16048), .B2(n16730), .A(n16047), .ZN(n16049) );
  OAI21_X1 U17127 ( .B1(n16726), .B2(n16050), .A(n16049), .ZN(n16106) );
  MUX2_X1 U17128 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n16106), .S(n16734), .Z(
        P1_U3550) );
  OAI211_X1 U17129 ( .C1(n16053), .C2(n16725), .A(n16052), .B(n16051), .ZN(
        n16054) );
  AOI211_X1 U17130 ( .C1(n16056), .C2(n16730), .A(n16055), .B(n16054), .ZN(
        n16057) );
  INV_X1 U17131 ( .A(n16057), .ZN(n16107) );
  MUX2_X1 U17132 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n16107), .S(n16734), .Z(
        P1_U3549) );
  AOI21_X1 U17133 ( .B1(n16059), .B2(n16606), .A(n16058), .ZN(n16061) );
  AND3_X1 U17134 ( .A1(n16062), .A2(n16061), .A3(n16060), .ZN(n16063) );
  OAI21_X1 U17135 ( .B1(n16064), .B2(n16540), .A(n16063), .ZN(n16108) );
  MUX2_X1 U17136 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n16108), .S(n16734), .Z(
        P1_U3548) );
  NAND2_X1 U17137 ( .A1(n16065), .A2(n16730), .ZN(n16070) );
  AOI211_X1 U17138 ( .C1(n16068), .C2(n16606), .A(n16067), .B(n16066), .ZN(
        n16069) );
  OAI211_X1 U17139 ( .C1(n16726), .C2(n16071), .A(n16070), .B(n16069), .ZN(
        n16109) );
  MUX2_X1 U17140 ( .A(n16109), .B(P1_REG1_REG_19__SCAN_IN), .S(n16732), .Z(
        P1_U3547) );
  INV_X1 U17141 ( .A(n16072), .ZN(n16077) );
  AOI21_X1 U17142 ( .B1(n16074), .B2(n16606), .A(n16073), .ZN(n16075) );
  OAI211_X1 U17143 ( .C1(n16077), .C2(n16475), .A(n16076), .B(n16075), .ZN(
        n16110) );
  MUX2_X1 U17144 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n16110), .S(n16734), .Z(
        P1_U3546) );
  AOI22_X1 U17145 ( .A1(n16080), .A2(n16079), .B1(n16078), .B2(n16606), .ZN(
        n16081) );
  OAI211_X1 U17146 ( .C1(n16083), .C2(n16540), .A(n16082), .B(n16081), .ZN(
        n16111) );
  MUX2_X1 U17147 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n16111), .S(n16734), .Z(
        P1_U3545) );
  AOI21_X1 U17148 ( .B1(n16085), .B2(n16606), .A(n16084), .ZN(n16086) );
  OAI211_X1 U17149 ( .C1(n16088), .C2(n16540), .A(n16087), .B(n16086), .ZN(
        n16112) );
  MUX2_X1 U17150 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n16112), .S(n16734), .Z(
        P1_U3544) );
  AOI21_X1 U17151 ( .B1(n16090), .B2(n16606), .A(n16089), .ZN(n16091) );
  OAI21_X1 U17152 ( .B1(n16092), .B2(n16464), .A(n16091), .ZN(n16093) );
  AOI21_X1 U17153 ( .B1(n16094), .B2(n16561), .A(n16093), .ZN(n16095) );
  OAI21_X1 U17154 ( .B1(n16096), .B2(n16540), .A(n16095), .ZN(n16113) );
  MUX2_X1 U17155 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n16113), .S(n16734), .Z(
        P1_U3543) );
  MUX2_X1 U17156 ( .A(n16098), .B(P1_REG0_REG_30__SCAN_IN), .S(n16735), .Z(
        P1_U3526) );
  MUX2_X1 U17157 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n16099), .S(n16737), .Z(
        P1_U3525) );
  MUX2_X1 U17158 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n16100), .S(n16737), .Z(
        P1_U3524) );
  MUX2_X1 U17159 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n16101), .S(n16737), .Z(
        P1_U3523) );
  MUX2_X1 U17160 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n16102), .S(n16737), .Z(
        P1_U3522) );
  MUX2_X1 U17161 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n16103), .S(n16737), .Z(
        P1_U3521) );
  MUX2_X1 U17162 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n16104), .S(n16737), .Z(
        P1_U3520) );
  MUX2_X1 U17163 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n16105), .S(n16737), .Z(
        P1_U3519) );
  MUX2_X1 U17164 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n16106), .S(n16737), .Z(
        P1_U3518) );
  MUX2_X1 U17165 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n16107), .S(n16737), .Z(
        P1_U3517) );
  MUX2_X1 U17166 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n16108), .S(n16737), .Z(
        P1_U3516) );
  MUX2_X1 U17167 ( .A(n16109), .B(P1_REG0_REG_19__SCAN_IN), .S(n16735), .Z(
        P1_U3515) );
  MUX2_X1 U17168 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n16110), .S(n16737), .Z(
        P1_U3513) );
  MUX2_X1 U17169 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n16111), .S(n16737), .Z(
        P1_U3510) );
  MUX2_X1 U17170 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n16112), .S(n16737), .Z(
        P1_U3507) );
  MUX2_X1 U17171 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n16113), .S(n16737), .Z(
        P1_U3504) );
  MUX2_X1 U17172 ( .A(n16114), .B(P1_D_REG_0__SCAN_IN), .S(n16144), .Z(
        P1_U3445) );
  NAND3_X1 U17173 ( .A1(n16115), .A2(P1_IR_REG_31__SCAN_IN), .A3(
        P1_STATE_REG_SCAN_IN), .ZN(n16116) );
  OAI22_X1 U17174 ( .A1(n16117), .A2(n16116), .B1(n13501), .B2(n16139), .ZN(
        n16118) );
  AOI21_X1 U17175 ( .B1(n15519), .B2(n16135), .A(n16118), .ZN(n16119) );
  INV_X1 U17176 ( .A(n16119), .ZN(P1_U3324) );
  OAI222_X1 U17177 ( .A1(n11886), .A2(n16122), .B1(P1_U3086), .B2(n16120), 
        .C1(n16121), .C2(n16139), .ZN(P1_U3325) );
  OAI222_X1 U17178 ( .A1(P1_U3086), .A2(n7417), .B1(n11886), .B2(n16124), .C1(
        n16139), .C2(n16123), .ZN(P1_U3328) );
  OAI222_X1 U17179 ( .A1(P1_U3086), .A2(n16127), .B1(n11886), .B2(n16126), 
        .C1(n16125), .C2(n16139), .ZN(P1_U3329) );
  INV_X1 U17180 ( .A(n16128), .ZN(n16129) );
  OAI222_X1 U17181 ( .A1(n16139), .A2(n16131), .B1(n11886), .B2(n16130), .C1(
        P1_U3086), .C2(n16129), .ZN(P1_U3330) );
  OAI222_X1 U17182 ( .A1(n16139), .A2(n16134), .B1(n11886), .B2(n16133), .C1(
        P1_U3086), .C2(n16132), .ZN(P1_U3331) );
  NAND2_X1 U17183 ( .A1(n16136), .A2(n16135), .ZN(n16138) );
  OAI211_X1 U17184 ( .C1(n16140), .C2(n16139), .A(n16138), .B(n16137), .ZN(
        P1_U3332) );
  MUX2_X1 U17185 ( .A(n16141), .B(n13607), .S(P1_STATE_REG_SCAN_IN), .Z(
        P1_U3333) );
  INV_X1 U17186 ( .A(n16142), .ZN(n16143) );
  MUX2_X1 U17187 ( .A(n16143), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  AND2_X1 U17188 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n16144), .ZN(P1_U3323) );
  AND2_X1 U17189 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n16144), .ZN(P1_U3322) );
  AND2_X1 U17190 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n16144), .ZN(P1_U3321) );
  AND2_X1 U17191 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n16144), .ZN(P1_U3320) );
  AND2_X1 U17192 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n16144), .ZN(P1_U3319) );
  AND2_X1 U17193 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n16144), .ZN(P1_U3318) );
  AND2_X1 U17194 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n16144), .ZN(P1_U3317) );
  AND2_X1 U17195 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n16144), .ZN(P1_U3316) );
  AND2_X1 U17196 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n16144), .ZN(P1_U3315) );
  AND2_X1 U17197 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n16144), .ZN(P1_U3314) );
  AND2_X1 U17198 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n16144), .ZN(P1_U3313) );
  AND2_X1 U17199 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n16144), .ZN(P1_U3312) );
  AND2_X1 U17200 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n16144), .ZN(P1_U3311) );
  AND2_X1 U17201 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n16144), .ZN(P1_U3310) );
  AND2_X1 U17202 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n16144), .ZN(P1_U3309) );
  AND2_X1 U17203 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n16144), .ZN(P1_U3308) );
  AND2_X1 U17204 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n16144), .ZN(P1_U3307) );
  AND2_X1 U17205 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n16144), .ZN(P1_U3306) );
  AND2_X1 U17206 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n16144), .ZN(P1_U3305) );
  AND2_X1 U17207 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n16144), .ZN(P1_U3304) );
  AND2_X1 U17208 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n16144), .ZN(P1_U3303) );
  AND2_X1 U17209 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n16144), .ZN(P1_U3302) );
  AND2_X1 U17210 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n16144), .ZN(P1_U3301) );
  AND2_X1 U17211 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n16144), .ZN(P1_U3300) );
  AND2_X1 U17212 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n16144), .ZN(P1_U3299) );
  AND2_X1 U17213 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n16144), .ZN(P1_U3298) );
  AND2_X1 U17214 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n16144), .ZN(P1_U3297) );
  AND2_X1 U17215 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n16144), .ZN(P1_U3296) );
  AND2_X1 U17216 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n16144), .ZN(P1_U3295) );
  AND2_X1 U17217 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n16144), .ZN(P1_U3294) );
  INV_X1 U17218 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n16146) );
  AOI21_X1 U17219 ( .B1(n16146), .B2(n16152), .A(n16145), .ZN(P2_U3417) );
  AND2_X1 U17220 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n16149), .ZN(P2_U3295) );
  AND2_X1 U17221 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n16149), .ZN(P2_U3294) );
  AND2_X1 U17222 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n16149), .ZN(P2_U3293) );
  AND2_X1 U17223 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n16149), .ZN(P2_U3292) );
  AND2_X1 U17224 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n16149), .ZN(P2_U3291) );
  AND2_X1 U17225 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n16149), .ZN(P2_U3290) );
  AND2_X1 U17226 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n16149), .ZN(P2_U3289) );
  AND2_X1 U17227 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n16149), .ZN(P2_U3288) );
  AND2_X1 U17228 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n16149), .ZN(P2_U3287) );
  AND2_X1 U17229 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n16149), .ZN(P2_U3286) );
  AND2_X1 U17230 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n16149), .ZN(P2_U3285) );
  AND2_X1 U17231 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n16149), .ZN(P2_U3284) );
  AND2_X1 U17232 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n16149), .ZN(P2_U3283) );
  AND2_X1 U17233 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n16149), .ZN(P2_U3282) );
  AND2_X1 U17234 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n16149), .ZN(P2_U3281) );
  AND2_X1 U17235 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n16149), .ZN(P2_U3280) );
  AND2_X1 U17236 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n16149), .ZN(P2_U3279) );
  AND2_X1 U17237 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n16149), .ZN(P2_U3278) );
  AND2_X1 U17238 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n16149), .ZN(P2_U3277) );
  AND2_X1 U17239 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n16149), .ZN(P2_U3276) );
  AND2_X1 U17240 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n16149), .ZN(P2_U3275) );
  AND2_X1 U17241 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n16149), .ZN(P2_U3274) );
  AND2_X1 U17242 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n16149), .ZN(P2_U3273) );
  AND2_X1 U17243 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n16149), .ZN(P2_U3272) );
  AND2_X1 U17244 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n16149), .ZN(P2_U3271) );
  AND2_X1 U17245 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n16149), .ZN(P2_U3270) );
  AND2_X1 U17246 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n16149), .ZN(P2_U3269) );
  AND2_X1 U17247 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n16149), .ZN(P2_U3268) );
  AND2_X1 U17248 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n16149), .ZN(P2_U3267) );
  AND2_X1 U17249 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n16149), .ZN(P2_U3266) );
  NOR2_X1 U17250 ( .A1(n10096), .A2(P2_U3947), .ZN(P2_U3087) );
  NOR2_X1 U17251 ( .A1(P3_U3897), .A2(n16150), .ZN(P3_U3150) );
  INV_X1 U17252 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n16153) );
  AOI21_X1 U17253 ( .B1(n16153), .B2(n16152), .A(n16151), .ZN(P2_U3416) );
  AOI21_X1 U17254 ( .B1(n16233), .B2(P2_REG1_REG_0__SCAN_IN), .A(n16154), .ZN(
        n16159) );
  AOI22_X1 U17255 ( .A1(P2_REG3_REG_0__SCAN_IN), .A2(P2_U3088), .B1(
        P2_ADDR_REG_0__SCAN_IN), .B2(n10096), .ZN(n16158) );
  OAI22_X1 U17256 ( .A1(n16220), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n16190), .ZN(n16156) );
  OAI21_X1 U17257 ( .B1(n16231), .B2(n16156), .A(P2_IR_REG_0__SCAN_IN), .ZN(
        n16157) );
  OAI211_X1 U17258 ( .C1(P2_IR_REG_0__SCAN_IN), .C2(n16159), .A(n16158), .B(
        n16157), .ZN(P2_U3214) );
  AOI22_X1 U17259 ( .A1(n10096), .A2(P2_ADDR_REG_3__SCAN_IN), .B1(n16231), 
        .B2(n16160), .ZN(n16171) );
  NAND2_X1 U17260 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_U3088), .ZN(n16170) );
  NAND2_X1 U17261 ( .A1(n16162), .A2(n16161), .ZN(n16163) );
  NAND3_X1 U17262 ( .A1(n16233), .A2(n16164), .A3(n16163), .ZN(n16169) );
  OAI211_X1 U17263 ( .C1(n16167), .C2(n16166), .A(n16229), .B(n16165), .ZN(
        n16168) );
  NAND4_X1 U17264 ( .A1(n16171), .A2(n16170), .A3(n16169), .A4(n16168), .ZN(
        P2_U3217) );
  AOI22_X1 U17265 ( .A1(n10096), .A2(P2_ADDR_REG_7__SCAN_IN), .B1(n16231), 
        .B2(n16172), .ZN(n16183) );
  NAND2_X1 U17266 ( .A1(n16174), .A2(n16173), .ZN(n16175) );
  NAND3_X1 U17267 ( .A1(n16176), .A2(n16233), .A3(n16175), .ZN(n16181) );
  OAI211_X1 U17268 ( .C1(n16179), .C2(n16178), .A(n16229), .B(n16177), .ZN(
        n16180) );
  NAND4_X1 U17269 ( .A1(n16183), .A2(n16182), .A3(n16181), .A4(n16180), .ZN(
        P2_U3221) );
  AOI22_X1 U17270 ( .A1(n10096), .A2(P2_ADDR_REG_11__SCAN_IN), .B1(n16231), 
        .B2(n16184), .ZN(n16197) );
  OAI21_X1 U17271 ( .B1(n16187), .B2(n16186), .A(n16185), .ZN(n16188) );
  NAND2_X1 U17272 ( .A1(n16188), .A2(n16229), .ZN(n16195) );
  AOI211_X1 U17273 ( .C1(n16192), .C2(n16191), .A(n16190), .B(n16189), .ZN(
        n16193) );
  INV_X1 U17274 ( .A(n16193), .ZN(n16194) );
  NAND4_X1 U17275 ( .A1(n16197), .A2(n16196), .A3(n16195), .A4(n16194), .ZN(
        P2_U3225) );
  OAI21_X1 U17276 ( .B1(n16214), .B2(n16199), .A(n16198), .ZN(n16200) );
  AOI21_X1 U17277 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(n10096), .A(n16200), 
        .ZN(n16209) );
  XOR2_X1 U17278 ( .A(n16202), .B(n16201), .Z(n16203) );
  NAND2_X1 U17279 ( .A1(n16203), .A2(n16233), .ZN(n16208) );
  OAI211_X1 U17280 ( .C1(n16206), .C2(n16205), .A(n16229), .B(n16204), .ZN(
        n16207) );
  NAND3_X1 U17281 ( .A1(n16209), .A2(n16208), .A3(n16207), .ZN(P2_U3230) );
  AOI21_X1 U17282 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n16211), .A(n16210), 
        .ZN(n16221) );
  OAI21_X1 U17283 ( .B1(n16214), .B2(n16213), .A(n16212), .ZN(n16215) );
  AOI21_X1 U17284 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n10096), .A(n16215), 
        .ZN(n16219) );
  XOR2_X1 U17285 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n16216), .Z(n16217) );
  NAND2_X1 U17286 ( .A1(n16217), .A2(n16233), .ZN(n16218) );
  OAI211_X1 U17287 ( .C1(n16221), .C2(n16220), .A(n16219), .B(n16218), .ZN(
        P2_U3232) );
  INV_X1 U17288 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n16238) );
  INV_X1 U17289 ( .A(n16222), .ZN(n16223) );
  OAI21_X1 U17290 ( .B1(n16225), .B2(n16224), .A(n16223), .ZN(n16234) );
  NAND2_X1 U17291 ( .A1(n16226), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n16227) );
  NAND2_X1 U17292 ( .A1(n16228), .A2(n16227), .ZN(n16230) );
  AOI222_X1 U17293 ( .A1(n16234), .A2(n16233), .B1(n16232), .B2(n16231), .C1(
        n16230), .C2(n16229), .ZN(n16236) );
  OAI211_X1 U17294 ( .C1(n16238), .C2(n16237), .A(n16236), .B(n16235), .ZN(
        P2_U3226) );
  INV_X1 U17295 ( .A(n16239), .ZN(n16245) );
  NAND2_X1 U17296 ( .A1(n7417), .A2(n10258), .ZN(n16243) );
  NAND2_X1 U17297 ( .A1(n16241), .A2(n16243), .ZN(n16242) );
  MUX2_X1 U17298 ( .A(n16243), .B(n16242), .S(P1_IR_REG_0__SCAN_IN), .Z(n16244) );
  NAND2_X1 U17299 ( .A1(n16245), .A2(n16244), .ZN(n16248) );
  AOI22_X1 U17300 ( .A1(P1_REG3_REG_0__SCAN_IN), .A2(P1_U3086), .B1(
        P1_ADDR_REG_0__SCAN_IN), .B2(n16246), .ZN(n16247) );
  OAI21_X1 U17301 ( .B1(n16249), .B2(n16248), .A(n16247), .ZN(P1_U3243) );
  OAI21_X1 U17302 ( .B1(n16252), .B2(n16251), .A(n16250), .ZN(n16264) );
  INV_X1 U17303 ( .A(n16253), .ZN(n16258) );
  NAND3_X1 U17304 ( .A1(n16256), .A2(n16255), .A3(n16254), .ZN(n16257) );
  NAND2_X1 U17305 ( .A1(n16258), .A2(n16257), .ZN(n16260) );
  AOI222_X1 U17306 ( .A1(n16264), .A2(n16263), .B1(n16262), .B2(n16261), .C1(
        n16260), .C2(n16259), .ZN(n16266) );
  OAI211_X1 U17307 ( .C1(n7637), .C2(n16267), .A(n16266), .B(n16265), .ZN(
        P1_U3255) );
  AOI21_X1 U17308 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(n16274), .A(n16270), .ZN(
        n16269) );
  INV_X1 U17309 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n16268) );
  NOR2_X1 U17310 ( .A1(n16269), .A2(n16268), .ZN(n16417) );
  AOI21_X1 U17311 ( .B1(n16269), .B2(n16268), .A(n16417), .ZN(SUB_1596_U53) );
  XOR2_X1 U17312 ( .A(n16271), .B(P2_ADDR_REG_1__SCAN_IN), .Z(n16416) );
  XOR2_X1 U17313 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(n16283), .Z(n16275) );
  AND2_X1 U17314 ( .A1(n16276), .A2(n16275), .ZN(n16280) );
  NOR2_X1 U17315 ( .A1(n16280), .A2(n16278), .ZN(n16277) );
  XOR2_X1 U17316 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(n16277), .Z(SUB_1596_U61) );
  NOR2_X1 U17317 ( .A1(n16280), .A2(n16279), .ZN(n16289) );
  XNOR2_X1 U17318 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(n16285), .ZN(n16288) );
  XNOR2_X1 U17319 ( .A(n16289), .B(n16288), .ZN(n16290) );
  XNOR2_X1 U17320 ( .A(P2_ADDR_REG_3__SCAN_IN), .B(n16290), .ZN(SUB_1596_U60)
         );
  NOR2_X1 U17321 ( .A1(n16284), .A2(n8009), .ZN(n16287) );
  NOR2_X1 U17322 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(n16285), .ZN(n16286) );
  XOR2_X1 U17323 ( .A(n16298), .B(n16297), .Z(SUB_1596_U59) );
  NAND2_X1 U17324 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n16306), .ZN(n16291) );
  OAI21_X1 U17325 ( .B1(n16306), .B2(P1_ADDR_REG_5__SCAN_IN), .A(n16291), .ZN(
        n16295) );
  NOR2_X1 U17326 ( .A1(n16292), .A2(n8522), .ZN(n16294) );
  XNOR2_X1 U17327 ( .A(n16295), .B(n16308), .ZN(n16302) );
  NAND2_X1 U17328 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(n16296), .ZN(n16299) );
  NOR2_X1 U17329 ( .A1(n16302), .A2(n16301), .ZN(n16303) );
  AOI21_X1 U17330 ( .B1(n16302), .B2(n16301), .A(n16303), .ZN(n16300) );
  INV_X1 U17331 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n16305) );
  XNOR2_X1 U17332 ( .A(n16300), .B(n16305), .ZN(SUB_1596_U58) );
  INV_X1 U17333 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n16414) );
  NAND2_X1 U17334 ( .A1(n16302), .A2(n16301), .ZN(n16304) );
  NOR2_X1 U17335 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(n16311), .ZN(n16314) );
  AOI21_X1 U17336 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(n16311), .A(n16314), .ZN(
        n16309) );
  XNOR2_X1 U17337 ( .A(n16313), .B(n16309), .ZN(n16412) );
  NAND2_X1 U17338 ( .A1(n16413), .A2(n16412), .ZN(n16310) );
  NOR2_X1 U17339 ( .A1(n16413), .A2(n16412), .ZN(n16411) );
  NAND2_X1 U17340 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(n16311), .ZN(n16312) );
  XNOR2_X1 U17341 ( .A(n16316), .B(n16315), .ZN(n16317) );
  XNOR2_X1 U17342 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n16317), .ZN(n16322) );
  XNOR2_X1 U17343 ( .A(n16323), .B(n16322), .ZN(SUB_1596_U56) );
  NOR2_X1 U17344 ( .A1(n16316), .A2(n16315), .ZN(n16319) );
  NOR2_X1 U17345 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n16317), .ZN(n16318) );
  INV_X1 U17346 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n16320) );
  AOI22_X1 U17347 ( .A1(P3_ADDR_REG_8__SCAN_IN), .A2(n16320), .B1(
        P1_ADDR_REG_8__SCAN_IN), .B2(n11611), .ZN(n16329) );
  XOR2_X1 U17348 ( .A(n16328), .B(n16329), .Z(n16326) );
  NOR2_X1 U17349 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n16321), .ZN(n16324) );
  NOR2_X1 U17350 ( .A1(n16326), .A2(n16325), .ZN(n16334) );
  NOR2_X1 U17351 ( .A1(n16334), .A2(n16333), .ZN(n16327) );
  XOR2_X1 U17352 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n16327), .Z(SUB_1596_U55) );
  NAND2_X1 U17353 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n11611), .ZN(n16330) );
  NOR2_X1 U17354 ( .A1(P1_ADDR_REG_9__SCAN_IN), .A2(n16439), .ZN(n16331) );
  AOI21_X1 U17355 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(n16439), .A(n16331), .ZN(
        n16332) );
  XOR2_X1 U17356 ( .A(n16335), .B(n16332), .Z(n16337) );
  XOR2_X1 U17357 ( .A(n16339), .B(P2_ADDR_REG_9__SCAN_IN), .Z(SUB_1596_U54) );
  AND2_X1 U17358 ( .A1(n16439), .A2(P1_ADDR_REG_9__SCAN_IN), .ZN(n16336) );
  XNOR2_X1 U17359 ( .A(P3_ADDR_REG_10__SCAN_IN), .B(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n16346) );
  XNOR2_X1 U17360 ( .A(n16345), .B(n16346), .ZN(n16343) );
  NAND2_X1 U17361 ( .A1(n16338), .A2(n16337), .ZN(n16340) );
  OAI21_X1 U17362 ( .B1(n16343), .B2(n16342), .A(n16344), .ZN(n16341) );
  XNOR2_X1 U17363 ( .A(n16341), .B(P2_ADDR_REG_10__SCAN_IN), .ZN(SUB_1596_U70)
         );
  INV_X1 U17364 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n16348) );
  XOR2_X1 U17365 ( .A(P3_ADDR_REG_11__SCAN_IN), .B(P1_ADDR_REG_11__SCAN_IN), 
        .Z(n16353) );
  XOR2_X1 U17366 ( .A(n16352), .B(n16353), .Z(n16350) );
  XNOR2_X1 U17367 ( .A(P2_ADDR_REG_11__SCAN_IN), .B(n16351), .ZN(SUB_1596_U69)
         );
  INV_X1 U17368 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n16354) );
  XNOR2_X1 U17369 ( .A(P3_ADDR_REG_12__SCAN_IN), .B(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n16358) );
  XNOR2_X1 U17370 ( .A(n16359), .B(n16358), .ZN(n16355) );
  XNOR2_X1 U17371 ( .A(P2_ADDR_REG_12__SCAN_IN), .B(n16357), .ZN(SUB_1596_U68)
         );
  XOR2_X1 U17372 ( .A(P3_ADDR_REG_13__SCAN_IN), .B(P1_ADDR_REG_13__SCAN_IN), 
        .Z(n16360) );
  XOR2_X1 U17373 ( .A(n16367), .B(n16360), .Z(n16362) );
  OAI21_X1 U17374 ( .B1(n16363), .B2(n16362), .A(n16364), .ZN(n16361) );
  XNOR2_X1 U17375 ( .A(n16361), .B(P2_ADDR_REG_13__SCAN_IN), .ZN(SUB_1596_U67)
         );
  INV_X1 U17376 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n16368) );
  NAND2_X1 U17377 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(n16365), .ZN(n16366) );
  XOR2_X1 U17378 ( .A(P3_ADDR_REG_14__SCAN_IN), .B(P1_ADDR_REG_14__SCAN_IN), 
        .Z(n16373) );
  XNOR2_X1 U17379 ( .A(n16374), .B(n16373), .ZN(n16370) );
  OAI21_X1 U17380 ( .B1(n16371), .B2(n16370), .A(n16372), .ZN(n16369) );
  XNOR2_X1 U17381 ( .A(n16369), .B(P2_ADDR_REG_14__SCAN_IN), .ZN(SUB_1596_U66)
         );
  INV_X1 U17382 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n16375) );
  XNOR2_X1 U17383 ( .A(P3_ADDR_REG_15__SCAN_IN), .B(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n16377) );
  XOR2_X1 U17384 ( .A(n16378), .B(n16377), .Z(n16381) );
  NAND2_X1 U17385 ( .A1(n16381), .A2(n16380), .ZN(n16382) );
  OAI21_X1 U17386 ( .B1(n16380), .B2(n16381), .A(n16382), .ZN(n16376) );
  XNOR2_X1 U17387 ( .A(n16376), .B(P2_ADDR_REG_15__SCAN_IN), .ZN(SUB_1596_U65)
         );
  INV_X1 U17388 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n16379) );
  XOR2_X1 U17389 ( .A(P1_ADDR_REG_16__SCAN_IN), .B(n16385), .Z(n16386) );
  XNOR2_X1 U17390 ( .A(P3_ADDR_REG_16__SCAN_IN), .B(n16386), .ZN(n16388) );
  AOI21_X1 U17391 ( .B1(n16388), .B2(n16389), .A(n16390), .ZN(n16384) );
  INV_X1 U17392 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n16391) );
  XNOR2_X1 U17393 ( .A(n16384), .B(n16391), .ZN(SUB_1596_U64) );
  NOR2_X1 U17394 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(n16385), .ZN(n16387) );
  XOR2_X1 U17395 ( .A(n16398), .B(P2_ADDR_REG_17__SCAN_IN), .Z(n16400) );
  XOR2_X1 U17396 ( .A(n16400), .B(n16399), .Z(SUB_1596_U63) );
  NOR2_X1 U17397 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(n16392), .ZN(n16395) );
  AND2_X1 U17398 ( .A1(P3_ADDR_REG_17__SCAN_IN), .A2(n16393), .ZN(n16394) );
  NOR2_X1 U17399 ( .A1(n16395), .A2(n16394), .ZN(n16403) );
  NOR2_X1 U17400 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n16404), .ZN(n16396) );
  AOI21_X1 U17401 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n16404), .A(n16396), 
        .ZN(n16397) );
  XOR2_X1 U17402 ( .A(n16403), .B(n16397), .Z(n16408) );
  NAND2_X1 U17403 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(n16398), .ZN(n16401) );
  XNOR2_X1 U17404 ( .A(P2_ADDR_REG_18__SCAN_IN), .B(n16409), .ZN(SUB_1596_U62)
         );
  AND2_X1 U17405 ( .A1(n16404), .A2(P1_ADDR_REG_18__SCAN_IN), .ZN(n16402) );
  OAI22_X1 U17406 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n16404), .B1(n16403), 
        .B2(n16402), .ZN(n16407) );
  XNOR2_X1 U17407 ( .A(n16405), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n16406) );
  XNOR2_X1 U17408 ( .A(n16407), .B(n16406), .ZN(n16410) );
  AOI21_X1 U17409 ( .B1(n16413), .B2(n16412), .A(n16411), .ZN(n16415) );
  XNOR2_X1 U17410 ( .A(n16415), .B(n16414), .ZN(SUB_1596_U57) );
  XOR2_X1 U17411 ( .A(n16417), .B(n16416), .Z(SUB_1596_U5) );
  AOI21_X1 U17412 ( .B1(n16420), .B2(n16419), .A(n16418), .ZN(n16434) );
  AOI21_X1 U17413 ( .B1(n16422), .B2(n12046), .A(n16421), .ZN(n16424) );
  NOR2_X1 U17414 ( .A1(n16424), .A2(n16423), .ZN(n16432) );
  AOI21_X1 U17415 ( .B1(n16426), .B2(n9628), .A(n16425), .ZN(n16430) );
  OAI22_X1 U17416 ( .A1(n16430), .A2(n16429), .B1(n16428), .B2(n16427), .ZN(
        n16431) );
  AOI211_X1 U17417 ( .C1(n16434), .C2(n16433), .A(n16432), .B(n16431), .ZN(
        n16437) );
  INV_X1 U17418 ( .A(n16435), .ZN(n16436) );
  OAI211_X1 U17419 ( .C1(n16439), .C2(n16438), .A(n16437), .B(n16436), .ZN(
        P3_U3191) );
  INV_X1 U17420 ( .A(P1_RD_REG_SCAN_IN), .ZN(n16441) );
  INV_X1 U17421 ( .A(P3_RD_REG_SCAN_IN), .ZN(n16440) );
  OAI221_X1 U17422 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .C1(n8925), .C2(n16441), .A(n16440), .ZN(U29) );
  INV_X1 U17423 ( .A(n16442), .ZN(n16443) );
  AOI211_X1 U17424 ( .C1(n16660), .C2(n16445), .A(n16444), .B(n16443), .ZN(
        n16446) );
  AOI22_X1 U17425 ( .A1(n16734), .A2(n16446), .B1(n10258), .B2(n16732), .ZN(
        P1_U3528) );
  AOI22_X1 U17426 ( .A1(n16737), .A2(n16446), .B1(n10252), .B2(n16735), .ZN(
        P1_U3459) );
  INV_X1 U17427 ( .A(n16447), .ZN(n16452) );
  AOI222_X1 U17428 ( .A1(n16452), .A2(n16451), .B1(n16450), .B2(n16449), .C1(
        n16497), .C2(n16448), .ZN(n16453) );
  OAI21_X1 U17429 ( .B1(n16454), .B2(n11306), .A(n16453), .ZN(P3_U3172) );
  INV_X1 U17430 ( .A(n16455), .ZN(n16459) );
  INV_X1 U17431 ( .A(n16456), .ZN(n16458) );
  AOI211_X1 U17432 ( .C1(n16596), .C2(n16459), .A(n16458), .B(n16457), .ZN(
        n16460) );
  AOI22_X1 U17433 ( .A1(n16718), .A2(n16460), .B1(n9592), .B2(n16717), .ZN(
        P3_U3460) );
  AOI22_X1 U17434 ( .A1(n14891), .A2(n16460), .B1(n8959), .B2(n16719), .ZN(
        P3_U3393) );
  XNOR2_X1 U17435 ( .A(n16468), .B(n16461), .ZN(n16487) );
  INV_X1 U17436 ( .A(n16487), .ZN(n16474) );
  AND2_X1 U17437 ( .A1(n16463), .A2(n16462), .ZN(n16482) );
  AOI211_X1 U17438 ( .C1(n16465), .C2(n16466), .A(n16464), .B(n7458), .ZN(
        n16485) );
  XNOR2_X1 U17439 ( .A(n16468), .B(n16467), .ZN(n16470) );
  OAI21_X1 U17440 ( .B1(n16470), .B2(n16726), .A(n16469), .ZN(n16471) );
  AOI21_X1 U17441 ( .B1(n16472), .B2(n16487), .A(n16471), .ZN(n16490) );
  OAI211_X1 U17442 ( .C1(n16475), .C2(n16474), .A(n16473), .B(n16490), .ZN(
        n16476) );
  INV_X1 U17443 ( .A(n16476), .ZN(n16478) );
  AOI22_X1 U17444 ( .A1(n16734), .A2(n16478), .B1(n16477), .B2(n16732), .ZN(
        P1_U3529) );
  AOI22_X1 U17445 ( .A1(n16737), .A2(n16478), .B1(n10357), .B2(n16735), .ZN(
        P1_U3462) );
  INV_X1 U17446 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n16479) );
  OAI22_X1 U17447 ( .A1(n16481), .A2(n16480), .B1(n16622), .B2(n16479), .ZN(
        n16484) );
  MUX2_X1 U17448 ( .A(n16482), .B(P1_REG2_REG_1__SCAN_IN), .S(n7414), .Z(
        n16483) );
  NOR2_X1 U17449 ( .A1(n16484), .A2(n16483), .ZN(n16489) );
  AOI22_X1 U17450 ( .A1(n16633), .A2(n16487), .B1(n16486), .B2(n16485), .ZN(
        n16488) );
  OAI211_X1 U17451 ( .C1(n7414), .C2(n16490), .A(n16489), .B(n16488), .ZN(
        P1_U3292) );
  INV_X1 U17452 ( .A(n16491), .ZN(n16492) );
  AOI21_X1 U17453 ( .B1(n16493), .B2(n16499), .A(n16492), .ZN(n16505) );
  INV_X1 U17454 ( .A(n16505), .ZN(n16514) );
  NOR2_X1 U17455 ( .A1(n16494), .A2(n16711), .ZN(n16507) );
  AOI22_X1 U17456 ( .A1(n16498), .A2(n16497), .B1(n16496), .B2(n16495), .ZN(
        n16504) );
  XNOR2_X1 U17457 ( .A(n16500), .B(n16499), .ZN(n16502) );
  NAND2_X1 U17458 ( .A1(n16502), .A2(n16501), .ZN(n16503) );
  OAI211_X1 U17459 ( .C1(n16505), .C2(n16521), .A(n16504), .B(n16503), .ZN(
        n16512) );
  AOI211_X1 U17460 ( .C1(n16596), .C2(n16514), .A(n16507), .B(n16512), .ZN(
        n16506) );
  AOI22_X1 U17461 ( .A1(n16718), .A2(n16506), .B1(n9598), .B2(n16717), .ZN(
        P3_U3461) );
  AOI22_X1 U17462 ( .A1(n14891), .A2(n16506), .B1(n8363), .B2(n16719), .ZN(
        P3_U3396) );
  INV_X1 U17463 ( .A(n16507), .ZN(n16511) );
  OAI22_X1 U17464 ( .A1(n16511), .A2(n16510), .B1(n16509), .B2(n16508), .ZN(
        n16513) );
  AOI211_X1 U17465 ( .C1(n16515), .C2(n16514), .A(n16513), .B(n16512), .ZN(
        n16516) );
  AOI22_X1 U17466 ( .A1(n16517), .A2(n9670), .B1(n16516), .B2(n14352), .ZN(
        P3_U3231) );
  AOI22_X1 U17467 ( .A1(n16737), .A2(n16518), .B1(n10394), .B2(n16735), .ZN(
        P1_U3465) );
  INV_X1 U17468 ( .A(n16519), .ZN(n16523) );
  AOI21_X1 U17469 ( .B1(n16521), .B2(n16615), .A(n16520), .ZN(n16522) );
  AOI211_X1 U17470 ( .C1(n16524), .C2(n16652), .A(n16523), .B(n16522), .ZN(
        n16526) );
  AOI22_X1 U17471 ( .A1(n16718), .A2(n16526), .B1(n9603), .B2(n16717), .ZN(
        P3_U3462) );
  INV_X1 U17472 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n16525) );
  AOI22_X1 U17473 ( .A1(n14891), .A2(n16526), .B1(n16525), .B2(n16719), .ZN(
        P3_U3399) );
  AND2_X1 U17474 ( .A1(n16606), .A2(n16527), .ZN(n16536) );
  AOI22_X1 U17475 ( .A1(n16528), .A2(n16536), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(P1_U3086), .ZN(n16534) );
  XOR2_X1 U17476 ( .A(n7626), .B(n16529), .Z(n16532) );
  AOI22_X1 U17477 ( .A1(n16532), .A2(n16531), .B1(n16530), .B2(n16537), .ZN(
        n16533) );
  OAI211_X1 U17478 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n16535), .A(n16534), .B(
        n16533), .ZN(P1_U3218) );
  NOR2_X1 U17479 ( .A1(n16537), .A2(n16536), .ZN(n16539) );
  OAI211_X1 U17480 ( .C1(n16541), .C2(n16540), .A(n16539), .B(n16538), .ZN(
        n16542) );
  AOI21_X1 U17481 ( .B1(n16561), .B2(n16543), .A(n16542), .ZN(n16545) );
  AOI22_X1 U17482 ( .A1(n16734), .A2(n16545), .B1(n10419), .B2(n16732), .ZN(
        P1_U3531) );
  INV_X1 U17483 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n16544) );
  AOI22_X1 U17484 ( .A1(n16737), .A2(n16545), .B1(n16544), .B2(n16735), .ZN(
        P1_U3468) );
  INV_X1 U17485 ( .A(n16546), .ZN(n16550) );
  OAI21_X1 U17486 ( .B1(n16548), .B2(n16711), .A(n16547), .ZN(n16549) );
  AOI21_X1 U17487 ( .B1(n16550), .B2(n16647), .A(n16549), .ZN(n16551) );
  AOI22_X1 U17488 ( .A1(n16718), .A2(n16551), .B1(n9653), .B2(n16717), .ZN(
        P3_U3463) );
  AOI22_X1 U17489 ( .A1(n14891), .A2(n16551), .B1(n9007), .B2(n16719), .ZN(
        P3_U3402) );
  NAND2_X1 U17490 ( .A1(n16552), .A2(n16730), .ZN(n16558) );
  INV_X1 U17491 ( .A(n16553), .ZN(n16557) );
  NAND2_X1 U17492 ( .A1(n16606), .A2(n16554), .ZN(n16555) );
  NAND4_X1 U17493 ( .A1(n16558), .A2(n16557), .A3(n16556), .A4(n16555), .ZN(
        n16559) );
  AOI21_X1 U17494 ( .B1(n16561), .B2(n16560), .A(n16559), .ZN(n16563) );
  INV_X1 U17495 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n16562) );
  AOI22_X1 U17496 ( .A1(n16734), .A2(n16563), .B1(n16562), .B2(n16732), .ZN(
        P1_U3532) );
  AOI22_X1 U17497 ( .A1(n16737), .A2(n16563), .B1(n10697), .B2(n16735), .ZN(
        P1_U3471) );
  INV_X1 U17498 ( .A(n16564), .ZN(n16568) );
  OAI22_X1 U17499 ( .A1(n16566), .A2(n16713), .B1(n16565), .B2(n16711), .ZN(
        n16567) );
  NOR2_X1 U17500 ( .A1(n16568), .A2(n16567), .ZN(n16570) );
  AOI22_X1 U17501 ( .A1(n16718), .A2(n16570), .B1(n9024), .B2(n16717), .ZN(
        P3_U3464) );
  INV_X1 U17502 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n16569) );
  AOI22_X1 U17503 ( .A1(n14891), .A2(n16570), .B1(n16569), .B2(n16719), .ZN(
        P3_U3405) );
  OAI21_X1 U17504 ( .B1(n16572), .B2(n16725), .A(n16571), .ZN(n16574) );
  AOI211_X1 U17505 ( .C1(n16660), .C2(n16575), .A(n16574), .B(n16573), .ZN(
        n16577) );
  AOI22_X1 U17506 ( .A1(n16734), .A2(n16577), .B1(n10715), .B2(n16732), .ZN(
        P1_U3533) );
  INV_X1 U17507 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n16576) );
  AOI22_X1 U17508 ( .A1(n16737), .A2(n16577), .B1(n16576), .B2(n16735), .ZN(
        P1_U3474) );
  INV_X1 U17509 ( .A(n16578), .ZN(n16583) );
  OAI21_X1 U17510 ( .B1(n16596), .B2(n16620), .A(n16579), .ZN(n16582) );
  NAND2_X1 U17511 ( .A1(n16580), .A2(n16652), .ZN(n16581) );
  AND3_X1 U17512 ( .A1(n16583), .A2(n16582), .A3(n16581), .ZN(n16584) );
  AOI22_X1 U17513 ( .A1(n16718), .A2(n16584), .B1(n9616), .B2(n16717), .ZN(
        P3_U3465) );
  AOI22_X1 U17514 ( .A1(n14891), .A2(n16584), .B1(n9043), .B2(n16719), .ZN(
        P3_U3408) );
  AOI21_X1 U17515 ( .B1(n16740), .B2(n16586), .A(n16585), .ZN(n16587) );
  OAI211_X1 U17516 ( .C1(n16590), .C2(n16589), .A(n16588), .B(n16587), .ZN(
        n16591) );
  INV_X1 U17517 ( .A(n16591), .ZN(n16594) );
  AOI22_X1 U17518 ( .A1(n16747), .A2(n16594), .B1(n16592), .B2(n16746), .ZN(
        P2_U3505) );
  INV_X1 U17519 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n16593) );
  AOI22_X1 U17520 ( .A1(n16751), .A2(n16594), .B1(n16593), .B2(n16748), .ZN(
        P2_U3448) );
  AOI22_X1 U17521 ( .A1(n16597), .A2(n16596), .B1(n16595), .B2(n16652), .ZN(
        n16599) );
  NAND2_X1 U17522 ( .A1(n16597), .A2(n16620), .ZN(n16598) );
  AOI22_X1 U17523 ( .A1(n16718), .A2(n16602), .B1(n9620), .B2(n16717), .ZN(
        P3_U3466) );
  INV_X1 U17524 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n16601) );
  AOI22_X1 U17525 ( .A1(n14891), .A2(n16602), .B1(n16601), .B2(n16719), .ZN(
        P3_U3411) );
  INV_X1 U17526 ( .A(n16603), .ZN(n16605) );
  AOI211_X1 U17527 ( .C1(n16607), .C2(n16606), .A(n16605), .B(n16604), .ZN(
        n16608) );
  OAI21_X1 U17528 ( .B1(n16726), .B2(n16609), .A(n16608), .ZN(n16610) );
  AOI21_X1 U17529 ( .B1(n16730), .B2(n16611), .A(n16610), .ZN(n16613) );
  AOI22_X1 U17530 ( .A1(n16734), .A2(n16613), .B1(n10824), .B2(n16732), .ZN(
        P1_U3535) );
  INV_X1 U17531 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n16612) );
  AOI22_X1 U17532 ( .A1(n16737), .A2(n16613), .B1(n16612), .B2(n16735), .ZN(
        P1_U3480) );
  INV_X1 U17533 ( .A(n16616), .ZN(n16619) );
  OAI22_X1 U17534 ( .A1(n16616), .A2(n16615), .B1(n16614), .B2(n16711), .ZN(
        n16618) );
  AOI211_X1 U17535 ( .C1(n16620), .C2(n16619), .A(n16618), .B(n16617), .ZN(
        n16621) );
  AOI22_X1 U17536 ( .A1(n16718), .A2(n16621), .B1(n9090), .B2(n16717), .ZN(
        P3_U3467) );
  AOI22_X1 U17537 ( .A1(n14891), .A2(n16621), .B1(n9086), .B2(n16719), .ZN(
        P3_U3414) );
  OAI22_X1 U17538 ( .A1(n16625), .A2(n16624), .B1(n16623), .B2(n16622), .ZN(
        n16626) );
  AOI21_X1 U17539 ( .B1(n16628), .B2(n16627), .A(n16626), .ZN(n16629) );
  OAI21_X1 U17540 ( .B1(n16631), .B2(n16630), .A(n16629), .ZN(n16632) );
  AOI21_X1 U17541 ( .B1(n16634), .B2(n16633), .A(n16632), .ZN(n16635) );
  OAI21_X1 U17542 ( .B1(n7414), .B2(n16636), .A(n16635), .ZN(P1_U3285) );
  OAI211_X1 U17543 ( .C1(n16639), .C2(n16678), .A(n16638), .B(n16637), .ZN(
        n16640) );
  AOI21_X1 U17544 ( .B1(n16642), .B2(n16641), .A(n16640), .ZN(n16645) );
  AOI22_X1 U17545 ( .A1(n16747), .A2(n16645), .B1(n16643), .B2(n16746), .ZN(
        P2_U3507) );
  INV_X1 U17546 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n16644) );
  AOI22_X1 U17547 ( .A1(n16751), .A2(n16645), .B1(n16644), .B2(n16748), .ZN(
        P2_U3454) );
  AND3_X1 U17548 ( .A1(n16648), .A2(n16647), .A3(n16646), .ZN(n16650) );
  AOI211_X1 U17549 ( .C1(n16652), .C2(n16651), .A(n16650), .B(n16649), .ZN(
        n16654) );
  AOI22_X1 U17550 ( .A1(n16718), .A2(n16654), .B1(n9628), .B2(n16717), .ZN(
        P3_U3468) );
  INV_X1 U17551 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n16653) );
  AOI22_X1 U17552 ( .A1(n14891), .A2(n16654), .B1(n16653), .B2(n16719), .ZN(
        P3_U3417) );
  OAI21_X1 U17553 ( .B1(n16656), .B2(n16725), .A(n16655), .ZN(n16658) );
  AOI211_X1 U17554 ( .C1(n16660), .C2(n16659), .A(n16658), .B(n16657), .ZN(
        n16662) );
  AOI22_X1 U17555 ( .A1(n16734), .A2(n16662), .B1(n11549), .B2(n16732), .ZN(
        P1_U3537) );
  INV_X1 U17556 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n16661) );
  AOI22_X1 U17557 ( .A1(n16737), .A2(n16662), .B1(n16661), .B2(n16735), .ZN(
        P1_U3486) );
  OAI22_X1 U17558 ( .A1(n16664), .A2(n16713), .B1(n16663), .B2(n16711), .ZN(
        n16666) );
  NOR2_X1 U17559 ( .A1(n16666), .A2(n16665), .ZN(n16668) );
  INV_X1 U17560 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n16667) );
  AOI22_X1 U17561 ( .A1(n16718), .A2(n16668), .B1(n16667), .B2(n16717), .ZN(
        P3_U3469) );
  AOI22_X1 U17562 ( .A1(n14891), .A2(n16668), .B1(n9110), .B2(n16719), .ZN(
        P3_U3420) );
  OAI211_X1 U17563 ( .C1(n16671), .C2(n16725), .A(n16670), .B(n16669), .ZN(
        n16674) );
  NOR2_X1 U17564 ( .A1(n16672), .A2(n16726), .ZN(n16673) );
  AOI211_X1 U17565 ( .C1(n16730), .C2(n16675), .A(n16674), .B(n16673), .ZN(
        n16676) );
  AOI22_X1 U17566 ( .A1(n16734), .A2(n16676), .B1(n10601), .B2(n16732), .ZN(
        P1_U3538) );
  AOI22_X1 U17567 ( .A1(n16737), .A2(n16676), .B1(n11567), .B2(n16735), .ZN(
        P1_U3489) );
  OAI21_X1 U17568 ( .B1(n16679), .B2(n16678), .A(n16677), .ZN(n16681) );
  AOI211_X1 U17569 ( .C1(n16704), .C2(n16682), .A(n16681), .B(n16680), .ZN(
        n16685) );
  AOI22_X1 U17570 ( .A1(n16747), .A2(n16685), .B1(n16683), .B2(n16746), .ZN(
        P2_U3509) );
  INV_X1 U17571 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n16684) );
  AOI22_X1 U17572 ( .A1(n16751), .A2(n16685), .B1(n16684), .B2(n16748), .ZN(
        P2_U3460) );
  OAI22_X1 U17573 ( .A1(n16687), .A2(n16713), .B1(n16686), .B2(n16711), .ZN(
        n16688) );
  NOR2_X1 U17574 ( .A1(n16689), .A2(n16688), .ZN(n16692) );
  AOI22_X1 U17575 ( .A1(n16718), .A2(n16692), .B1(n16690), .B2(n16717), .ZN(
        P3_U3470) );
  INV_X1 U17576 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n16691) );
  AOI22_X1 U17577 ( .A1(n14891), .A2(n16692), .B1(n16691), .B2(n16719), .ZN(
        P3_U3423) );
  OAI21_X1 U17578 ( .B1(n16694), .B2(n16725), .A(n16693), .ZN(n16695) );
  AOI211_X1 U17579 ( .C1(n16697), .C2(n16730), .A(n16696), .B(n16695), .ZN(
        n16699) );
  AOI22_X1 U17580 ( .A1(n16734), .A2(n16699), .B1(n11575), .B2(n16732), .ZN(
        P1_U3539) );
  INV_X1 U17581 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n16698) );
  AOI22_X1 U17582 ( .A1(n16737), .A2(n16699), .B1(n16698), .B2(n16735), .ZN(
        P1_U3492) );
  NAND2_X1 U17583 ( .A1(n16700), .A2(n16740), .ZN(n16701) );
  NAND2_X1 U17584 ( .A1(n16702), .A2(n16701), .ZN(n16703) );
  AOI21_X1 U17585 ( .B1(n16705), .B2(n16704), .A(n16703), .ZN(n16706) );
  AND2_X1 U17586 ( .A1(n16707), .A2(n16706), .ZN(n16710) );
  AOI22_X1 U17587 ( .A1(n16747), .A2(n16710), .B1(n16708), .B2(n16746), .ZN(
        P2_U3511) );
  INV_X1 U17588 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n16709) );
  AOI22_X1 U17589 ( .A1(n16751), .A2(n16710), .B1(n16709), .B2(n16748), .ZN(
        P2_U3466) );
  OAI22_X1 U17590 ( .A1(n16714), .A2(n16713), .B1(n16712), .B2(n16711), .ZN(
        n16715) );
  NOR2_X1 U17591 ( .A1(n16716), .A2(n16715), .ZN(n16721) );
  AOI22_X1 U17592 ( .A1(n16718), .A2(n16721), .B1(n9155), .B2(n16717), .ZN(
        P3_U3472) );
  INV_X1 U17593 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n16720) );
  AOI22_X1 U17594 ( .A1(n14891), .A2(n16721), .B1(n16720), .B2(n16719), .ZN(
        P3_U3429) );
  OAI211_X1 U17595 ( .C1(n7730), .C2(n16725), .A(n16724), .B(n16723), .ZN(
        n16729) );
  NOR2_X1 U17596 ( .A1(n16727), .A2(n16726), .ZN(n16728) );
  AOI211_X1 U17597 ( .C1(n16731), .C2(n16730), .A(n16729), .B(n16728), .ZN(
        n16736) );
  AOI22_X1 U17598 ( .A1(n16734), .A2(n16736), .B1(n16733), .B2(n16732), .ZN(
        P1_U3541) );
  AOI22_X1 U17599 ( .A1(n16737), .A2(n16736), .B1(n12013), .B2(n16735), .ZN(
        P1_U3498) );
  OR2_X1 U17600 ( .A1(n16739), .A2(n16738), .ZN(n16745) );
  NAND2_X1 U17601 ( .A1(n16741), .A2(n16740), .ZN(n16742) );
  AND4_X1 U17602 ( .A1(n16745), .A2(n16744), .A3(n16743), .A4(n16742), .ZN(
        n16750) );
  AOI22_X1 U17603 ( .A1(n16747), .A2(n16750), .B1(n11807), .B2(n16746), .ZN(
        P2_U3513) );
  INV_X1 U17604 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n16749) );
  AOI22_X1 U17605 ( .A1(n16751), .A2(n16750), .B1(n16749), .B2(n16748), .ZN(
        P2_U3472) );
  AOI21_X1 U17606 ( .B1(P1_WR_REG_SCAN_IN), .B2(P2_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n16752) );
  OAI21_X1 U17607 ( .B1(P1_WR_REG_SCAN_IN), .B2(P2_WR_REG_SCAN_IN), .A(n16752), 
        .ZN(U28) );
  CLKBUF_X1 U7514 ( .A(n8980), .Z(n9308) );
  CLKBUF_X2 U8159 ( .A(n8984), .Z(n9644) );
  OAI21_X1 U8206 ( .B1(n14977), .B2(n7926), .A(n7924), .ZN(n14945) );
endmodule

