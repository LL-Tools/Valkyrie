

module b21_C_gen_AntiSAT_k_256_4 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2, 
        keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7, 
        keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12, 
        keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17, 
        keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22, 
        keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27, 
        keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32, 
        keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37, 
        keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42, 
        keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47, 
        keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52, 
        keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57, 
        keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62, 
        keyinput_f63, keyinput_f64, keyinput_f65, keyinput_f66, keyinput_f67, 
        keyinput_f68, keyinput_f69, keyinput_f70, keyinput_f71, keyinput_f72, 
        keyinput_f73, keyinput_f74, keyinput_f75, keyinput_f76, keyinput_f77, 
        keyinput_f78, keyinput_f79, keyinput_f80, keyinput_f81, keyinput_f82, 
        keyinput_f83, keyinput_f84, keyinput_f85, keyinput_f86, keyinput_f87, 
        keyinput_f88, keyinput_f89, keyinput_f90, keyinput_f91, keyinput_f92, 
        keyinput_f93, keyinput_f94, keyinput_f95, keyinput_f96, keyinput_f97, 
        keyinput_f98, keyinput_f99, keyinput_f100, keyinput_f101, 
        keyinput_f102, keyinput_f103, keyinput_f104, keyinput_f105, 
        keyinput_f106, keyinput_f107, keyinput_f108, keyinput_f109, 
        keyinput_f110, keyinput_f111, keyinput_f112, keyinput_f113, 
        keyinput_f114, keyinput_f115, keyinput_f116, keyinput_f117, 
        keyinput_f118, keyinput_f119, keyinput_f120, keyinput_f121, 
        keyinput_f122, keyinput_f123, keyinput_f124, keyinput_f125, 
        keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, keyinput_g2, 
        keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, 
        keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, 
        keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, 
        keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, 
        keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, 
        keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, 
        keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, 
        keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, 
        keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, 
        keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, 
        keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, 
        keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, 
        keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, keyinput_g67, 
        keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, keyinput_g72, 
        keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, keyinput_g77, 
        keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, keyinput_g82, 
        keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, keyinput_g87, 
        keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, keyinput_g92, 
        keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, keyinput_g97, 
        keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101, 
        keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105, 
        keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109, 
        keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113, 
        keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117, 
        keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121, 
        keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125, 
        keyinput_g126, keyinput_g127, ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, 
        ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, 
        ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, 
        ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, 
        ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, P1_U3352, P1_U3351, 
        P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, 
        P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, 
        P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, 
        P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, 
        P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, 
        P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, 
        P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, 
        P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, 
        P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, 
        P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, 
        P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, 
        P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, 
        P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, 
        P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, 
        P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, 
        P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, 
        P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, 
        P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, 
        P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, 
        P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, 
        P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, 
        P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, 
        P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, 
        P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, 
        P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, 
        P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, 
        P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, 
        P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, 
        P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, 
        P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, 
        P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, 
        P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, 
        P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, 
        P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, 
        P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, 
        P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, 
        P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, 
        P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, 
        P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, 
        P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, 
        P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, 
        P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, 
        P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, 
        P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, 
        P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, 
        P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, 
        P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, 
        P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3152, P2_U3151, P2_U3966 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2,
         keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7,
         keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12,
         keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17,
         keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22,
         keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27,
         keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32,
         keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37,
         keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42,
         keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47,
         keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52,
         keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57,
         keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62,
         keyinput_f63, keyinput_f64, keyinput_f65, keyinput_f66, keyinput_f67,
         keyinput_f68, keyinput_f69, keyinput_f70, keyinput_f71, keyinput_f72,
         keyinput_f73, keyinput_f74, keyinput_f75, keyinput_f76, keyinput_f77,
         keyinput_f78, keyinput_f79, keyinput_f80, keyinput_f81, keyinput_f82,
         keyinput_f83, keyinput_f84, keyinput_f85, keyinput_f86, keyinput_f87,
         keyinput_f88, keyinput_f89, keyinput_f90, keyinput_f91, keyinput_f92,
         keyinput_f93, keyinput_f94, keyinput_f95, keyinput_f96, keyinput_f97,
         keyinput_f98, keyinput_f99, keyinput_f100, keyinput_f101,
         keyinput_f102, keyinput_f103, keyinput_f104, keyinput_f105,
         keyinput_f106, keyinput_f107, keyinput_f108, keyinput_f109,
         keyinput_f110, keyinput_f111, keyinput_f112, keyinput_f113,
         keyinput_f114, keyinput_f115, keyinput_f116, keyinput_f117,
         keyinput_f118, keyinput_f119, keyinput_f120, keyinput_f121,
         keyinput_f122, keyinput_f123, keyinput_f124, keyinput_f125,
         keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, keyinput_g2,
         keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7,
         keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12,
         keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17,
         keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22,
         keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27,
         keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32,
         keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37,
         keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42,
         keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47,
         keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52,
         keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57,
         keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62,
         keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, keyinput_g67,
         keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, keyinput_g72,
         keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, keyinput_g77,
         keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, keyinput_g82,
         keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, keyinput_g87,
         keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, keyinput_g92,
         keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, keyinput_g97,
         keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101,
         keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105,
         keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109,
         keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113,
         keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117,
         keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121,
         keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125,
         keyinput_g126, keyinput_g127;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486,
         n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496,
         n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506,
         n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516,
         n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526,
         n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536,
         n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546,
         n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556,
         n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566,
         n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576,
         n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586,
         n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596,
         n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606,
         n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616,
         n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626,
         n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636,
         n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646,
         n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656,
         n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666,
         n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676,
         n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686,
         n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696,
         n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706,
         n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716,
         n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726,
         n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736,
         n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746,
         n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756,
         n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766,
         n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776,
         n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786,
         n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796,
         n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806,
         n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816,
         n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826,
         n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836,
         n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846,
         n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856,
         n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866,
         n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876,
         n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886,
         n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896,
         n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906,
         n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916,
         n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926,
         n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936,
         n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946,
         n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956,
         n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966,
         n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976,
         n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986,
         n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996,
         n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006,
         n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016,
         n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026,
         n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036,
         n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046,
         n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056,
         n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066,
         n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076,
         n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086,
         n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096,
         n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106,
         n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116,
         n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126,
         n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136,
         n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146,
         n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156,
         n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166,
         n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176,
         n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186,
         n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196,
         n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206,
         n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216,
         n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226,
         n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236,
         n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246,
         n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256,
         n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266,
         n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276,
         n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286,
         n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296,
         n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306,
         n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316,
         n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326,
         n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336,
         n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346,
         n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356,
         n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366,
         n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376,
         n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386,
         n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396,
         n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406,
         n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416,
         n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426,
         n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436,
         n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446,
         n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456,
         n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466,
         n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476,
         n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486,
         n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496,
         n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506,
         n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516,
         n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526,
         n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536,
         n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546,
         n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556,
         n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566,
         n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576,
         n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5586, n5587,
         n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597,
         n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607,
         n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617,
         n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627,
         n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637,
         n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647,
         n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657,
         n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667,
         n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677,
         n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687,
         n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697,
         n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707,
         n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717,
         n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727,
         n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737,
         n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747,
         n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757,
         n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767,
         n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777,
         n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787,
         n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797,
         n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807,
         n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817,
         n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827,
         n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837,
         n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847,
         n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857,
         n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867,
         n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877,
         n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887,
         n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897,
         n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907,
         n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917,
         n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927,
         n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937,
         n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947,
         n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957,
         n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967,
         n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977,
         n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987,
         n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997,
         n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007,
         n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017,
         n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027,
         n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037,
         n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047,
         n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057,
         n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067,
         n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077,
         n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087,
         n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097,
         n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107,
         n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117,
         n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127,
         n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137,
         n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147,
         n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157,
         n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167,
         n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177,
         n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187,
         n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197,
         n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207,
         n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217,
         n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227,
         n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237,
         n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247,
         n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257,
         n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267,
         n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277,
         n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287,
         n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297,
         n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307,
         n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317,
         n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327,
         n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337,
         n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347,
         n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357,
         n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367,
         n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377,
         n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387,
         n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397,
         n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407,
         n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417,
         n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427,
         n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437,
         n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447,
         n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457,
         n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467,
         n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477,
         n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487,
         n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497,
         n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507,
         n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517,
         n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527,
         n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537,
         n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547,
         n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557,
         n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567,
         n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577,
         n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587,
         n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597,
         n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607,
         n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617,
         n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627,
         n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637,
         n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647,
         n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657,
         n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667,
         n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677,
         n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687,
         n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697,
         n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707,
         n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717,
         n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727,
         n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737,
         n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747,
         n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757,
         n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767,
         n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777,
         n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787,
         n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797,
         n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807,
         n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817,
         n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827,
         n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837,
         n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847,
         n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857,
         n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867,
         n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877,
         n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887,
         n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897,
         n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907,
         n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917,
         n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927,
         n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937,
         n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947,
         n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957,
         n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967,
         n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977,
         n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987,
         n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997,
         n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007,
         n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017,
         n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027,
         n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037,
         n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047,
         n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057,
         n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067,
         n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077,
         n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087,
         n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097,
         n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107,
         n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117,
         n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127,
         n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137,
         n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147,
         n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157,
         n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167,
         n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177,
         n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187,
         n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197,
         n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207,
         n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217,
         n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227,
         n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237,
         n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247,
         n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257,
         n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267,
         n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277,
         n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287,
         n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297,
         n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307,
         n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317,
         n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327,
         n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337,
         n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347,
         n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357,
         n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367,
         n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377,
         n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387,
         n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397,
         n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407,
         n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417,
         n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427,
         n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437,
         n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447,
         n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457,
         n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467,
         n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477,
         n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487,
         n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497,
         n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507,
         n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517,
         n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527,
         n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537,
         n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547,
         n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557,
         n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567,
         n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577,
         n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587,
         n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597,
         n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607,
         n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617,
         n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627,
         n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637,
         n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647,
         n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657,
         n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667,
         n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677,
         n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687,
         n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697,
         n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707,
         n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717,
         n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727,
         n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737,
         n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747,
         n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757,
         n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767,
         n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777,
         n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787,
         n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797,
         n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807,
         n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817,
         n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827,
         n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837,
         n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847,
         n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857,
         n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867,
         n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877,
         n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887,
         n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897,
         n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907,
         n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917,
         n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927,
         n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937,
         n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947,
         n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957,
         n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967,
         n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977,
         n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987,
         n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997,
         n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007,
         n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017,
         n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027,
         n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037,
         n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047,
         n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057,
         n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067,
         n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077,
         n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087,
         n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097,
         n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107,
         n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117,
         n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127,
         n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137,
         n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147,
         n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157,
         n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167,
         n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177,
         n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187,
         n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197,
         n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207,
         n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217,
         n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227,
         n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237,
         n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247,
         n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257,
         n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267,
         n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277,
         n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287,
         n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297,
         n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307,
         n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317,
         n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327,
         n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337,
         n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347,
         n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357,
         n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367,
         n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377,
         n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387,
         n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397,
         n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407,
         n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417,
         n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427,
         n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437,
         n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447,
         n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457,
         n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467,
         n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477,
         n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487,
         n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497,
         n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507,
         n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517,
         n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527,
         n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537,
         n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547,
         n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557,
         n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567,
         n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577,
         n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587,
         n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597,
         n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607,
         n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617,
         n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627,
         n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637,
         n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647,
         n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657,
         n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667,
         n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677,
         n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687,
         n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697,
         n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707,
         n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8716, n8717, n8718,
         n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728,
         n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738,
         n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748,
         n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758,
         n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768,
         n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778,
         n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788,
         n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798,
         n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808,
         n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818,
         n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828,
         n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838,
         n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848,
         n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858,
         n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868,
         n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8879,
         n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889,
         n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899,
         n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909,
         n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919,
         n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929,
         n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939,
         n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949,
         n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959,
         n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969,
         n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979,
         n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989,
         n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999,
         n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009,
         n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019,
         n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029,
         n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039,
         n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049,
         n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059,
         n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069,
         n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079,
         n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089,
         n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099,
         n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109,
         n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119,
         n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129,
         n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139,
         n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149,
         n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159,
         n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169,
         n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179,
         n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189,
         n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199,
         n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209,
         n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219,
         n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229,
         n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239,
         n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249,
         n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259,
         n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269,
         n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279,
         n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289,
         n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299,
         n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309,
         n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319,
         n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329,
         n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339,
         n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349,
         n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359,
         n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369,
         n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379,
         n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389,
         n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399,
         n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409,
         n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419,
         n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429,
         n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439,
         n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449,
         n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459,
         n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469,
         n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479,
         n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489,
         n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499,
         n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509,
         n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519,
         n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529,
         n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539,
         n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549,
         n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559,
         n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569,
         n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579,
         n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589,
         n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599,
         n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609,
         n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619,
         n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629,
         n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639,
         n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649,
         n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659,
         n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669,
         n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679,
         n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689,
         n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699,
         n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709,
         n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719,
         n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729,
         n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739,
         n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749,
         n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759,
         n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769,
         n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779,
         n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789,
         n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799,
         n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809,
         n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819,
         n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829,
         n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839,
         n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849,
         n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859,
         n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869,
         n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879,
         n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889,
         n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899,
         n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909,
         n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919,
         n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929,
         n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939,
         n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949,
         n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959,
         n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969,
         n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979,
         n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989,
         n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999,
         n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553;

  AOI21_X1 U4982 ( .B1(n8844), .B2(n8810), .A(n8809), .ZN(n8811) );
  OR2_X1 U4983 ( .A1(n8001), .A2(n8000), .ZN(n8002) );
  NAND2_X1 U4984 ( .A1(n8574), .A2(n8534), .ZN(n8538) );
  INV_X2 U4985 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  NAND2_X1 U4986 ( .A1(n4880), .A2(n4879), .ZN(n8589) );
  NAND2_X1 U4987 ( .A1(n8642), .A2(n8628), .ZN(n8627) );
  NAND2_X1 U4988 ( .A1(n8767), .A2(n8674), .ZN(n8659) );
  NAND2_X1 U4989 ( .A1(n5026), .A2(n5028), .ZN(n7068) );
  OR2_X1 U4990 ( .A1(n7395), .A2(n7228), .ZN(n8307) );
  CLKBUF_X2 U4991 ( .A(n5268), .Z(n8016) );
  NAND2_X1 U4992 ( .A1(n6322), .A2(n9073), .ZN(n6319) );
  INV_X4 U4993 ( .A(n4484), .ZN(n7936) );
  CLKBUF_X2 U4994 ( .A(n7421), .Z(n4480) );
  CLKBUF_X2 U4995 ( .A(n6404), .Z(n9118) );
  CLKBUF_X2 U4996 ( .A(n5259), .Z(n5815) );
  CLKBUF_X1 U4997 ( .A(n5230), .Z(n5802) );
  NAND4_X1 U4998 ( .A1(n6142), .A2(n6141), .A3(n6140), .A4(n6139), .ZN(n9359)
         );
  NOR2_X1 U5000 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n5340) );
  INV_X1 U5001 ( .A(n6589), .ZN(n6576) );
  INV_X1 U5002 ( .A(n5263), .ZN(n8007) );
  INV_X1 U5003 ( .A(n5231), .ZN(n7673) );
  NOR2_X2 U5004 ( .A1(n8659), .A2(n8760), .ZN(n8642) );
  NAND2_X1 U5005 ( .A1(n7242), .A2(n7241), .ZN(n7396) );
  NAND2_X1 U5006 ( .A1(n5589), .A2(n8395), .ZN(n5212) );
  NAND2_X1 U5007 ( .A1(n8641), .A2(n8640), .ZN(n8761) );
  NAND2_X1 U5008 ( .A1(n5441), .A2(n5440), .ZN(n7395) );
  NAND2_X1 U5009 ( .A1(n5346), .A2(n5345), .ZN(n6960) );
  BUF_X1 U5010 ( .A(n6300), .Z(n6842) );
  INV_X1 U5011 ( .A(n9263), .ZN(n9338) );
  NAND2_X1 U5012 ( .A1(n6404), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n4824) );
  OAI211_X2 U5013 ( .C1(n6842), .C2(n6309), .A(n6308), .B(n6307), .ZN(n6310)
         );
  XNOR2_X1 U5014 ( .A(n6136), .B(P1_IR_REG_30__SCAN_IN), .ZN(n6138) );
  OAI21_X1 U5015 ( .B1(n7615), .B2(n5307), .A(n7613), .ZN(n7618) );
  AOI21_X1 U5016 ( .B1(n8773), .B2(n8810), .A(n8731), .ZN(n8732) );
  INV_X1 U5017 ( .A(n6042), .ZN(n7702) );
  INV_X1 U5019 ( .A(n9358), .ZN(n7603) );
  NAND4_X1 U5020 ( .A1(n6298), .A2(n6297), .A3(n6296), .A4(n6295), .ZN(n9357)
         );
  INV_X1 U5022 ( .A(n6138), .ZN(n9771) );
  AND3_X1 U5023 ( .A1(n4697), .A2(n5114), .A3(n4508), .ZN(n4477) );
  INV_X1 U5024 ( .A(n5257), .ZN(n4478) );
  AND2_X1 U5025 ( .A1(n5843), .A2(n7590), .ZN(n5257) );
  NOR2_X4 U5026 ( .A1(n4502), .A2(n8843), .ZN(n8674) );
  NAND2_X2 U5027 ( .A1(n5196), .A2(n5195), .ZN(n5294) );
  AOI21_X2 U5028 ( .B1(n8654), .B2(n8655), .A(n7637), .ZN(n8641) );
  XNOR2_X2 U5029 ( .A(n6118), .B(n6117), .ZN(n6945) );
  NOR3_X2 U5030 ( .A1(n9599), .A2(n9701), .A3(n4700), .ZN(n4698) );
  NAND2_X2 U5031 ( .A1(n8256), .A2(n6048), .ZN(n7112) );
  AOI21_X2 U5032 ( .B1(n7581), .B2(n8325), .A(n7580), .ZN(n7660) );
  OAI21_X2 U5033 ( .B1(n7542), .B2(n8241), .A(n8239), .ZN(n7581) );
  OR2_X2 U5034 ( .A1(n6409), .A2(n6306), .ZN(n6307) );
  OR2_X2 U5035 ( .A1(n8706), .A2(n8775), .ZN(n4502) );
  NOR2_X2 U5036 ( .A1(n5429), .A2(n5473), .ZN(n5454) );
  NAND2_X2 U5037 ( .A1(n5411), .A2(n5410), .ZN(n8722) );
  INV_X1 U5038 ( .A(n8426), .ZN(n6041) );
  NAND2_X2 U5039 ( .A1(n5237), .A2(n5236), .ZN(n8426) );
  INV_X2 U5040 ( .A(n4478), .ZN(n4479) );
  AND2_X2 U5041 ( .A1(n7620), .A2(n7619), .ZN(n8534) );
  AND2_X1 U5042 ( .A1(n7596), .A2(n9771), .ZN(n7421) );
  AOI21_X2 U5043 ( .B1(n7397), .B2(n4515), .A(n5076), .ZN(n7484) );
  NAND2_X2 U5044 ( .A1(n5393), .A2(n5392), .ZN(n7157) );
  NAND4_X4 U5045 ( .A1(n4826), .A2(n6270), .A3(n4825), .A4(n4824), .ZN(n9358)
         );
  NAND2_X2 U5046 ( .A1(n5055), .A2(n6945), .ZN(n6380) );
  INV_X2 U5047 ( .A(n6119), .ZN(n5055) );
  BUF_X4 U5048 ( .A(n4827), .Z(n4481) );
  XNOR2_X2 U5049 ( .A(n4738), .B(n5470), .ZN(n7372) );
  NAND2_X1 U5050 ( .A1(n5215), .A2(n5214), .ZN(n4482) );
  NAND2_X1 U5052 ( .A1(n8534), .A2(n8408), .ZN(n8227) );
  NAND2_X1 U5053 ( .A1(n7371), .A2(n7370), .ZN(n7705) );
  NAND2_X1 U5054 ( .A1(n4781), .A2(n7270), .ZN(n7327) );
  NOR3_X1 U5055 ( .A1(n9202), .A2(n9201), .A3(n9200), .ZN(n9204) );
  MUX2_X1 U5056 ( .A(n9153), .B(n9152), .S(n9256), .Z(n9156) );
  AND2_X2 U5057 ( .A1(n7468), .A2(n7467), .ZN(n7487) );
  NOR2_X2 U5058 ( .A1(n4496), .A2(n7462), .ZN(n7468) );
  INV_X4 U5059 ( .A(n10366), .ZN(n10362) );
  INV_X1 U5060 ( .A(n9356), .ZN(n6423) );
  INV_X2 U5061 ( .A(n6553), .ZN(n6566) );
  INV_X2 U5062 ( .A(n4484), .ZN(n7973) );
  CLKBUF_X2 U5063 ( .A(n6576), .Z(n7956) );
  NAND2_X1 U5064 ( .A1(n8254), .A2(n8257), .ZN(n6049) );
  INV_X1 U5065 ( .A(n8423), .ZN(n7608) );
  INV_X1 U5066 ( .A(n7890), .ZN(n4484) );
  NAND2_X1 U5067 ( .A1(n8426), .A2(n7702), .ZN(n6048) );
  BUF_X2 U5068 ( .A(n5313), .Z(n8189) );
  AND2_X1 U5069 ( .A1(n7596), .A2(n6138), .ZN(n6404) );
  INV_X1 U5070 ( .A(n7120), .ZN(n10465) );
  NAND2_X1 U5071 ( .A1(n5843), .A2(n8185), .ZN(n5295) );
  NOR2_X1 U5072 ( .A1(n8870), .A2(n5161), .ZN(n5230) );
  NAND2_X2 U5073 ( .A1(n5893), .A2(n5942), .ZN(n6300) );
  NOR2_X1 U5074 ( .A1(n8185), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8869) );
  NAND4_X1 U5075 ( .A1(n5136), .A2(n5135), .A3(n5218), .A4(n4609), .ZN(n5174)
         );
  INV_X4 U5076 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  NOR2_X1 U5077 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n5134) );
  NAND2_X1 U5078 ( .A1(n4815), .A2(n4814), .ZN(n5042) );
  AOI21_X1 U5079 ( .B1(n8195), .B2(n4582), .A(n4505), .ZN(n8406) );
  NAND2_X1 U5080 ( .A1(n9020), .A2(n9021), .ZN(n4816) );
  NAND2_X1 U5081 ( .A1(n8924), .A2(n7921), .ZN(n9020) );
  OR2_X1 U5082 ( .A1(n8397), .A2(n4717), .ZN(n4716) );
  OAI211_X1 U5083 ( .C1(n9001), .C2(n4555), .A(n4786), .B(n4785), .ZN(n8964)
         );
  NOR2_X1 U5084 ( .A1(n8737), .A2(n4513), .ZN(n8740) );
  AOI21_X1 U5085 ( .B1(n4575), .B2(n4574), .A(n4519), .ZN(n8193) );
  OR2_X1 U5086 ( .A1(n8743), .A2(n8742), .ZN(n8816) );
  OR2_X1 U5087 ( .A1(n7783), .A2(n7782), .ZN(n9010) );
  INV_X1 U5088 ( .A(n4894), .ZN(n4893) );
  NAND2_X1 U5089 ( .A1(n4807), .A2(n4806), .ZN(n7724) );
  NAND2_X1 U5090 ( .A1(n8233), .A2(n4896), .ZN(n4895) );
  NAND2_X1 U5091 ( .A1(n6916), .A2(n6915), .ZN(n6950) );
  NAND2_X1 U5092 ( .A1(n6948), .A2(n6947), .ZN(n6946) );
  NAND2_X1 U5093 ( .A1(n6914), .A2(n6913), .ZN(n6925) );
  MUX2_X1 U5094 ( .A(n9256), .B(n9145), .S(n9144), .Z(n9157) );
  AND2_X1 U5095 ( .A1(n5020), .A2(n5499), .ZN(n5019) );
  NAND2_X1 U5096 ( .A1(n7229), .A2(n8306), .ZN(n7397) );
  OR2_X1 U5097 ( .A1(n5022), .A2(n5021), .ZN(n5020) );
  OAI21_X1 U5098 ( .B1(n5704), .B2(n5703), .A(n5702), .ZN(n5725) );
  NAND2_X1 U5099 ( .A1(n6817), .A2(n6874), .ZN(n6868) );
  INV_X1 U5100 ( .A(n5066), .ZN(n7229) );
  AOI21_X1 U5101 ( .B1(n5040), .B2(n5039), .A(n6231), .ZN(n7615) );
  NAND2_X1 U5102 ( .A1(n5485), .A2(n5484), .ZN(n7462) );
  OR2_X1 U5103 ( .A1(n5713), .A2(n10069), .ZN(n5737) );
  OAI21_X1 U5104 ( .B1(n5454), .B2(n5471), .A(n5478), .ZN(n4738) );
  NAND2_X1 U5105 ( .A1(n6323), .A2(n9278), .ZN(n4823) );
  AND2_X2 U5106 ( .A1(n6821), .A2(n10208), .ZN(n10456) );
  NAND2_X1 U5107 ( .A1(n5269), .A2(n8059), .ZN(n8069) );
  OAI21_X1 U5108 ( .B1(n5359), .B2(n4742), .A(n4740), .ZN(n5477) );
  OAI21_X1 U5109 ( .B1(n6613), .B2(n6612), .A(n9555), .ZN(n9047) );
  INV_X2 U5110 ( .A(n10399), .ZN(n4483) );
  NAND2_X1 U5111 ( .A1(n9072), .A2(n9078), .ZN(n9276) );
  NAND2_X1 U5112 ( .A1(n7688), .A2(n7689), .ZN(n8058) );
  NAND2_X1 U5113 ( .A1(n5336), .A2(n5335), .ZN(n5359) );
  INV_X1 U5114 ( .A(n10444), .ZN(n6515) );
  NAND2_X1 U5115 ( .A1(n6462), .A2(n4612), .ZN(n8950) );
  XNOR2_X1 U5116 ( .A(n5217), .B(n5216), .ZN(n6411) );
  INV_X1 U5117 ( .A(n9515), .ZN(n9544) );
  CLKBUF_X1 U5118 ( .A(n5245), .Z(n7667) );
  NAND2_X1 U5119 ( .A1(n5257), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5240) );
  NAND2_X1 U5120 ( .A1(n5784), .A2(n4820), .ZN(n6618) );
  NOR2_X1 U5121 ( .A1(n7593), .A2(n8870), .ZN(n5246) );
  AND2_X1 U5122 ( .A1(n6134), .A2(n6133), .ZN(n6137) );
  AND2_X2 U5123 ( .A1(n8870), .A2(n7593), .ZN(n5245) );
  INV_X1 U5124 ( .A(n5161), .ZN(n7593) );
  OAI21_X1 U5125 ( .B1(n6126), .B2(n6125), .A(P1_IR_REG_29__SCAN_IN), .ZN(
        n6134) );
  NAND2_X1 U5126 ( .A1(n9766), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6136) );
  NAND2_X1 U5127 ( .A1(n5160), .A2(n4498), .ZN(n5161) );
  MUX2_X1 U5128 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5159), .S(
        P2_IR_REG_29__SCAN_IN), .Z(n5160) );
  XNOR2_X1 U5129 ( .A(n5158), .B(P2_IR_REG_30__SCAN_IN), .ZN(n8870) );
  NAND2_X1 U5130 ( .A1(n6130), .A2(n6129), .ZN(n9766) );
  MUX2_X1 U5131 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5201), .S(
        P2_IR_REG_27__SCAN_IN), .Z(n5202) );
  NAND2_X1 U5132 ( .A1(n4696), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5128) );
  NAND2_X1 U5133 ( .A1(n5082), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5158) );
  XNOR2_X1 U5134 ( .A(n5170), .B(n5169), .ZN(n8395) );
  OAI21_X1 U5135 ( .B1(n5168), .B2(P2_IR_REG_21__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5167) );
  NAND2_X1 U5136 ( .A1(n5168), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5170) );
  INV_X2 U5137 ( .A(n9768), .ZN(n9773) );
  NAND3_X1 U5138 ( .A1(n4695), .A2(n4694), .A3(n4477), .ZN(n4696) );
  NAND2_X2 U5139 ( .A1(n8185), .A2(P1_U3084), .ZN(n9774) );
  XNOR2_X1 U5140 ( .A(n5176), .B(n5175), .ZN(n8517) );
  AND3_X1 U5141 ( .A1(n4697), .A2(n4517), .A3(n5114), .ZN(n5096) );
  AND3_X1 U5142 ( .A1(n4987), .A2(n4517), .A3(n5099), .ZN(n4695) );
  AND2_X1 U5143 ( .A1(n5099), .A2(n4508), .ZN(n5113) );
  INV_X1 U5144 ( .A(n5778), .ZN(n5099) );
  AND2_X1 U5145 ( .A1(n4818), .A2(n5103), .ZN(n4697) );
  AND4_X1 U5146 ( .A1(n5133), .A2(n5459), .A3(n5341), .A4(n5509), .ZN(n5135)
         );
  NAND2_X1 U5147 ( .A1(n10175), .A2(n4968), .ZN(n4967) );
  AND2_X1 U5148 ( .A1(n5799), .A2(n5808), .ZN(n4818) );
  AND4_X1 U5149 ( .A1(n10097), .A2(n6023), .A3(n10108), .A4(n5100), .ZN(n5101)
         );
  AND3_X1 U5150 ( .A1(n4776), .A2(n4775), .A3(n6022), .ZN(n5102) );
  AND2_X2 U5151 ( .A1(n5258), .A2(n5134), .ZN(n5218) );
  AND2_X1 U5152 ( .A1(n5791), .A2(n10145), .ZN(n5114) );
  CLKBUF_X1 U5153 ( .A(P2_IR_REG_0__SCAN_IN), .Z(n10413) );
  NOR2_X2 U5154 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5258) );
  INV_X1 U5155 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5808) );
  INV_X1 U5156 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5341) );
  NOR2_X1 U5157 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n5132) );
  NOR2_X1 U5158 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n5131) );
  NOR2_X1 U5159 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n5130) );
  NOR2_X1 U5160 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n5133) );
  INV_X1 U5161 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5137) );
  INV_X1 U5162 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n10108) );
  INV_X1 U5163 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n10097) );
  INV_X1 U5164 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5509) );
  INV_X1 U5165 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5459) );
  INV_X1 U5166 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5775) );
  INV_X1 U5167 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5098) );
  AND2_X1 U5168 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5298) );
  INV_X1 U5169 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n6117) );
  INV_X1 U5170 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n6022) );
  INV_X1 U5171 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n6023) );
  NOR2_X1 U5172 ( .A1(P1_IR_REG_29__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n6131) );
  NOR2_X1 U5173 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n4776) );
  NOR2_X1 U5174 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n4775) );
  INV_X1 U5175 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n10145) );
  NOR2_X1 U5176 ( .A1(P1_ADDR_REG_19__SCAN_IN), .A2(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n10176) );
  INV_X1 U5177 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n9967) );
  INV_X1 U5178 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5121) );
  AND2_X1 U5179 ( .A1(P1_ADDR_REG_19__SCAN_IN), .A2(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n10175) );
  AOI21_X1 U5180 ( .B1(n9228), .B2(n9481), .A(n9227), .ZN(n9240) );
  NOR4_X2 U5182 ( .A1(n9157), .A2(n9156), .A3(n9155), .A4(n9154), .ZN(n9170)
         );
  INV_X2 U5183 ( .A(n5520), .ZN(n5284) );
  XNOR2_X2 U5184 ( .A(n7999), .B(n8000), .ZN(n7998) );
  AND2_X1 U5185 ( .A1(n6122), .A2(n6121), .ZN(n9515) );
  XNOR2_X2 U5186 ( .A(n5750), .B(n5751), .ZN(n5749) );
  OAI21_X2 U5187 ( .B1(n4585), .B2(n5037), .A(n5035), .ZN(n8155) );
  NAND2_X2 U5188 ( .A1(n8003), .A2(n8002), .ZN(n4585) );
  OR2_X2 U5189 ( .A1(n10204), .A2(n10227), .ZN(n4496) );
  NAND2_X2 U5190 ( .A1(n5206), .A2(n5205), .ZN(n5602) );
  NAND2_X2 U5191 ( .A1(n4587), .A2(n4586), .ZN(n5040) );
  NOR2_X2 U5192 ( .A1(n7161), .A2(n8722), .ZN(n7234) );
  NOR2_X1 U5193 ( .A1(n9655), .A2(n9407), .ZN(n9326) );
  INV_X1 U5194 ( .A(n7927), .ZN(n7926) );
  NAND2_X1 U5195 ( .A1(n4931), .A2(n4934), .ZN(n8171) );
  AOI21_X1 U5196 ( .B1(n4935), .B2(n7585), .A(n4563), .ZN(n4934) );
  NAND2_X1 U5197 ( .A1(n7569), .A2(n4932), .ZN(n4931) );
  OAI21_X1 U5198 ( .B1(n5538), .B2(n4955), .A(n4952), .ZN(n5629) );
  INV_X1 U5199 ( .A(n4956), .ZN(n4955) );
  AOI21_X1 U5200 ( .B1(n4956), .B2(n4954), .A(n4953), .ZN(n4952) );
  AND2_X1 U5201 ( .A1(n4957), .A2(n5555), .ZN(n4956) );
  AOI22_X1 U5202 ( .A1(n9357), .A2(n7320), .B1(n7890), .B2(n6690), .ZN(n6555)
         );
  NAND2_X1 U5203 ( .A1(n8348), .A2(n8354), .ZN(n4754) );
  INV_X1 U5204 ( .A(n5470), .ZN(n5479) );
  INV_X1 U5205 ( .A(n5495), .ZN(n5021) );
  NAND2_X1 U5206 ( .A1(n4506), .A2(n9655), .ZN(n9250) );
  NAND2_X1 U5207 ( .A1(n4611), .A2(n9354), .ZN(n9308) );
  INV_X1 U5208 ( .A(n8950), .ZN(n4611) );
  NOR2_X1 U5209 ( .A1(n5471), .A2(n5479), .ZN(n5474) );
  OAI21_X1 U5210 ( .B1(n5293), .B2(n4943), .A(n5310), .ZN(n4942) );
  OR2_X1 U5211 ( .A1(n8810), .A2(n8192), .ZN(n8388) );
  NOR2_X1 U5212 ( .A1(n10212), .A2(n5079), .ZN(n5078) );
  INV_X1 U5213 ( .A(n8307), .ZN(n5079) );
  OR2_X1 U5214 ( .A1(n8775), .A2(n8095), .ZN(n8350) );
  INV_X1 U5215 ( .A(n5174), .ZN(n5173) );
  INV_X1 U5216 ( .A(n7857), .ZN(n4789) );
  NOR2_X1 U5217 ( .A1(n9424), .A2(n4855), .ZN(n4854) );
  NAND2_X1 U5218 ( .A1(n4856), .A2(n9268), .ZN(n4855) );
  OR2_X1 U5219 ( .A1(n9671), .A2(n9415), .ZN(n9423) );
  OR2_X1 U5220 ( .A1(n9664), .A2(n9430), .ZN(n9241) );
  OAI21_X1 U5221 ( .B1(n4648), .B2(n4544), .A(n9478), .ZN(n4647) );
  NOR2_X1 U5222 ( .A1(n4544), .A2(n4644), .ZN(n4643) );
  INV_X1 U5223 ( .A(n8038), .ZN(n4644) );
  NAND2_X1 U5224 ( .A1(n9681), .A2(n9027), .ZN(n9231) );
  INV_X1 U5225 ( .A(n9209), .ZN(n4838) );
  AND2_X1 U5226 ( .A1(n9554), .A2(n9539), .ZN(n9274) );
  OAI21_X1 U5227 ( .B1(n7188), .B2(n4973), .A(n4971), .ZN(n10241) );
  INV_X1 U5228 ( .A(n4974), .ZN(n4973) );
  AOI21_X1 U5229 ( .B1(n4974), .B2(n4972), .A(n4551), .ZN(n4971) );
  NAND2_X1 U5230 ( .A1(n7527), .A2(n7526), .ZN(n7569) );
  OAI21_X1 U5231 ( .B1(n7505), .B2(n7504), .A(n7503), .ZN(n7525) );
  AND2_X1 U5232 ( .A1(n4990), .A2(n5108), .ZN(n4989) );
  AND2_X1 U5233 ( .A1(n5684), .A2(n5667), .ZN(n5682) );
  OAI21_X1 U5234 ( .B1(n5504), .B2(n5503), .A(n5502), .ZN(n5538) );
  INV_X1 U5235 ( .A(n5500), .ZN(n5503) );
  AND2_X1 U5236 ( .A1(n5404), .A2(n5363), .ZN(n5381) );
  NAND2_X1 U5237 ( .A1(n5337), .A2(n10147), .ZN(n5360) );
  INV_X1 U5238 ( .A(n5331), .ZN(n5332) );
  AOI21_X1 U5239 ( .B1(n4608), .B2(n8077), .A(n4546), .ZN(n4604) );
  INV_X1 U5240 ( .A(n8023), .ZN(n5010) );
  NAND2_X1 U5241 ( .A1(n5012), .A2(n5009), .ZN(n5008) );
  INV_X1 U5242 ( .A(n5295), .ZN(n5313) );
  NAND2_X1 U5243 ( .A1(n5151), .A2(n5084), .ZN(n5203) );
  INV_X1 U5244 ( .A(n5086), .ZN(n5084) );
  NAND2_X1 U5245 ( .A1(n4678), .A2(n4492), .ZN(n4675) );
  NOR2_X1 U5246 ( .A1(n8569), .A2(n8371), .ZN(n5074) );
  NAND2_X1 U5247 ( .A1(n8633), .A2(n7664), .ZN(n8615) );
  NAND2_X1 U5248 ( .A1(n8799), .A2(n8414), .ZN(n4918) );
  INV_X1 U5249 ( .A(n8325), .ZN(n7539) );
  AND2_X1 U5250 ( .A1(n8239), .A2(n7480), .ZN(n8321) );
  AND2_X1 U5251 ( .A1(n8297), .A2(n6964), .ZN(n4915) );
  AND2_X1 U5252 ( .A1(n8289), .A2(n8290), .ZN(n8286) );
  OR2_X1 U5253 ( .A1(n8783), .A2(n8686), .ZN(n7633) );
  NAND2_X1 U5254 ( .A1(n6555), .A2(n6554), .ZN(n6559) );
  INV_X1 U5255 ( .A(n6409), .ZN(n7785) );
  AND2_X1 U5256 ( .A1(n7871), .A2(n7870), .ZN(n8968) );
  OR2_X1 U5257 ( .A1(n7965), .A2(n7964), .ZN(n9433) );
  INV_X1 U5258 ( .A(n9344), .ZN(n9481) );
  AOI21_X1 U5259 ( .B1(n9606), .B2(n9728), .A(n9612), .ZN(n9598) );
  NAND2_X1 U5260 ( .A1(n8029), .A2(n8031), .ZN(n4660) );
  NAND2_X1 U5261 ( .A1(n4993), .A2(n4991), .ZN(n6714) );
  AND2_X1 U5262 ( .A1(n9282), .A2(n4992), .ZN(n4991) );
  INV_X1 U5263 ( .A(n5097), .ZN(n4992) );
  NAND2_X1 U5264 ( .A1(n6300), .A2(n7590), .ZN(n6715) );
  NOR2_X1 U5265 ( .A1(n7461), .A2(n7364), .ZN(n4820) );
  AND2_X1 U5266 ( .A1(n4542), .A2(n5093), .ZN(n5059) );
  INV_X1 U5267 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n6357) );
  AND2_X1 U5268 ( .A1(n4601), .A2(n4606), .ZN(n4599) );
  NAND2_X1 U5269 ( .A1(n8069), .A2(n5273), .ZN(n6183) );
  INV_X1 U5270 ( .A(n5271), .ZN(n5272) );
  OR2_X1 U5271 ( .A1(n8559), .A2(n7625), .ZN(n7630) );
  INV_X1 U5272 ( .A(n5042), .ZN(n5049) );
  NAND2_X1 U5273 ( .A1(n5047), .A2(n5046), .ZN(n5045) );
  INV_X1 U5274 ( .A(n8875), .ZN(n5046) );
  NOR2_X1 U5275 ( .A1(n9333), .A2(n6945), .ZN(n4951) );
  NAND2_X1 U5276 ( .A1(n4948), .A2(n4947), .ZN(n4946) );
  NAND2_X1 U5277 ( .A1(n9334), .A2(n6945), .ZN(n4944) );
  OAI21_X1 U5278 ( .B1(n9400), .B2(n9399), .A(n4768), .ZN(n4767) );
  AOI21_X1 U5279 ( .B1(n9401), .B2(n10332), .A(n10324), .ZN(n4768) );
  NAND2_X1 U5280 ( .A1(n4754), .A2(n8382), .ZN(n4753) );
  INV_X1 U5281 ( .A(n4734), .ZN(n4733) );
  INV_X1 U5282 ( .A(n10247), .ZN(n4866) );
  NOR2_X1 U5283 ( .A1(n9140), .A2(n9132), .ZN(n4846) );
  INV_X1 U5284 ( .A(n5380), .ZN(n5033) );
  INV_X1 U5285 ( .A(n5376), .ZN(n5030) );
  INV_X1 U5286 ( .A(n7104), .ZN(n5027) );
  AND2_X1 U5287 ( .A1(n4595), .A2(n5526), .ZN(n4589) );
  OR2_X1 U5288 ( .A1(n8833), .A2(n8638), .ZN(n8361) );
  NOR2_X1 U5289 ( .A1(n8799), .A2(n8794), .ZN(n4877) );
  OR2_X1 U5290 ( .A1(n8794), .A2(n8143), .ZN(n8236) );
  OR2_X1 U5291 ( .A1(n7462), .A2(n10218), .ZN(n4911) );
  NAND2_X1 U5292 ( .A1(n7397), .A2(n8302), .ZN(n5080) );
  OAI21_X1 U5293 ( .B1(n8297), .B2(n5062), .A(n8295), .ZN(n5061) );
  NAND2_X1 U5294 ( .A1(n5063), .A2(n8292), .ZN(n5062) );
  INV_X1 U5295 ( .A(n8266), .ZN(n5073) );
  NAND2_X1 U5296 ( .A1(n6284), .A2(n8254), .ZN(n6794) );
  INV_X1 U5297 ( .A(n6783), .ZN(n8263) );
  NAND2_X1 U5298 ( .A1(n5588), .A2(n5600), .ZN(n5268) );
  OR2_X1 U5299 ( .A1(n8534), .A2(n8408), .ZN(n8378) );
  OR2_X1 U5300 ( .A1(n8823), .A2(n8074), .ZN(n8369) );
  OR2_X1 U5301 ( .A1(n8828), .A2(n8586), .ZN(n8230) );
  NOR2_X1 U5302 ( .A1(n4883), .A2(n4504), .ZN(n4882) );
  INV_X1 U5303 ( .A(n4889), .ZN(n4883) );
  INV_X1 U5304 ( .A(n8901), .ZN(n4788) );
  NOR2_X1 U5305 ( .A1(n4555), .A2(n7856), .ZN(n4783) );
  INV_X1 U5306 ( .A(n8966), .ZN(n7900) );
  NAND2_X1 U5307 ( .A1(n8976), .A2(n6573), .ZN(n6747) );
  XNOR2_X1 U5308 ( .A(n9429), .B(n9422), .ZN(n4870) );
  NAND2_X1 U5309 ( .A1(n9069), .A2(n9268), .ZN(n4853) );
  NOR2_X1 U5310 ( .A1(n8047), .A2(n9065), .ZN(n4856) );
  NOR2_X1 U5311 ( .A1(n9681), .A2(n8039), .ZN(n4708) );
  NOR2_X1 U5312 ( .A1(n9674), .A2(n4707), .ZN(n4706) );
  INV_X1 U5313 ( .A(n4708), .ZN(n4707) );
  OR2_X1 U5314 ( .A1(n9674), .A2(n9481), .ZN(n9269) );
  OR2_X1 U5315 ( .A1(n9701), .A2(n9563), .ZN(n9211) );
  AND2_X1 U5316 ( .A1(n4535), .A2(n4629), .ZN(n4628) );
  NAND2_X1 U5317 ( .A1(n4630), .A2(n8032), .ZN(n4629) );
  AND2_X1 U5318 ( .A1(n9712), .A2(n9564), .ZN(n9203) );
  OR2_X1 U5319 ( .A1(n9715), .A2(n9573), .ZN(n9199) );
  NAND2_X1 U5320 ( .A1(n4866), .A2(n4863), .ZN(n4862) );
  INV_X1 U5321 ( .A(n10248), .ZN(n4863) );
  NAND2_X1 U5322 ( .A1(n7381), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n7419) );
  NAND2_X1 U5323 ( .A1(n7190), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n7289) );
  INV_X1 U5324 ( .A(n7192), .ZN(n7190) );
  OR2_X1 U5325 ( .A1(n7407), .A2(n7286), .ZN(n9161) );
  INV_X1 U5326 ( .A(n4846), .ZN(n4843) );
  AOI21_X1 U5327 ( .B1(n4488), .B2(n4618), .A(n4553), .ZN(n4617) );
  NAND2_X1 U5328 ( .A1(n4616), .A2(n4488), .ZN(n4615) );
  NAND2_X1 U5329 ( .A1(n6604), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n6729) );
  INV_X1 U5330 ( .A(n6606), .ZN(n6604) );
  INV_X1 U5331 ( .A(n9766), .ZN(n6132) );
  NAND2_X1 U5332 ( .A1(n7454), .A2(n7453), .ZN(n7505) );
  NAND2_X1 U5333 ( .A1(n7450), .A2(n7449), .ZN(n7454) );
  AOI21_X1 U5334 ( .B1(n4926), .B2(n4928), .A(n4924), .ZN(n4923) );
  INV_X1 U5335 ( .A(n5684), .ZN(n4924) );
  NAND2_X1 U5336 ( .A1(n4966), .A2(n4964), .ZN(n5504) );
  NOR2_X1 U5337 ( .A1(n5475), .A2(n4965), .ZN(n4964) );
  AND2_X1 U5338 ( .A1(n5474), .A2(n5473), .ZN(n5475) );
  AND2_X1 U5339 ( .A1(n5477), .A2(n5472), .ZN(n5429) );
  NAND2_X1 U5340 ( .A1(n5360), .A2(n5339), .ZN(n5358) );
  INV_X1 U5341 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5791) );
  OAI21_X1 U5342 ( .B1(n7590), .B2(n4579), .A(n4578), .ZN(n5194) );
  NAND2_X1 U5343 ( .A1(n7590), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n4578) );
  OAI21_X1 U5344 ( .B1(n7590), .B2(n4577), .A(n4576), .ZN(n5191) );
  INV_X1 U5345 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n4577) );
  NAND2_X1 U5346 ( .A1(n7590), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n4576) );
  INV_X1 U5347 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4968) );
  NAND2_X1 U5348 ( .A1(n7618), .A2(n4588), .ZN(n5613) );
  OR2_X1 U5349 ( .A1(n5308), .A2(n5309), .ZN(n4588) );
  XNOR2_X1 U5350 ( .A(n5252), .B(n5034), .ZN(n7688) );
  INV_X1 U5351 ( .A(n5251), .ZN(n5034) );
  INV_X1 U5352 ( .A(n5642), .ZN(n5017) );
  OR2_X1 U5353 ( .A1(n8139), .A2(n5017), .ZN(n5016) );
  INV_X1 U5354 ( .A(n8081), .ZN(n5014) );
  AND2_X1 U5355 ( .A1(n7173), .A2(n5453), .ZN(n5022) );
  NAND2_X1 U5356 ( .A1(n7068), .A2(n5449), .ZN(n7071) );
  NAND2_X1 U5357 ( .A1(n5268), .A2(n8426), .ZN(n5251) );
  NOR2_X1 U5358 ( .A1(n5593), .A2(n5024), .ZN(n5023) );
  INV_X1 U5359 ( .A(n5554), .ZN(n5024) );
  NAND2_X1 U5360 ( .A1(n5036), .A2(n8100), .ZN(n5035) );
  AND2_X1 U5361 ( .A1(n8101), .A2(n5038), .ZN(n5037) );
  INV_X1 U5362 ( .A(n8101), .ZN(n5036) );
  INV_X1 U5363 ( .A(n8584), .ZN(n8225) );
  NAND2_X1 U5364 ( .A1(n4677), .A2(n7700), .ZN(n4676) );
  INV_X1 U5365 ( .A(n4679), .ZN(n4677) );
  AND2_X1 U5366 ( .A1(n8434), .A2(n8435), .ZN(n8432) );
  OR2_X1 U5367 ( .A1(n5870), .A2(n5869), .ZN(n4687) );
  OR2_X1 U5368 ( .A1(n5881), .A2(n5880), .ZN(n4685) );
  AND2_X1 U5369 ( .A1(n4685), .A2(n4684), .ZN(n5919) );
  NAND2_X1 U5370 ( .A1(n5916), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n4684) );
  OR2_X1 U5371 ( .A1(n5919), .A2(n5918), .ZN(n4683) );
  NAND2_X1 U5372 ( .A1(n7554), .A2(n4667), .ZN(n8454) );
  OR2_X1 U5373 ( .A1(n7555), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n4667) );
  NOR2_X1 U5374 ( .A1(n8498), .A2(n4568), .ZN(n8500) );
  NAND2_X1 U5375 ( .A1(n8500), .A2(n8501), .ZN(n8511) );
  NAND2_X1 U5376 ( .A1(n8361), .A2(n8360), .ZN(n8613) );
  NAND2_X1 U5377 ( .A1(n5736), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5762) );
  INV_X1 U5378 ( .A(n5737), .ZN(n5736) );
  NOR2_X1 U5379 ( .A1(n8662), .A2(n8669), .ZN(n7637) );
  AND2_X1 U5380 ( .A1(n8236), .A2(n8238), .ZN(n8325) );
  OR2_X1 U5381 ( .A1(n7482), .A2(n8321), .ZN(n4919) );
  OAI21_X1 U5382 ( .B1(n5078), .B2(n5077), .A(n8313), .ZN(n5076) );
  INV_X1 U5383 ( .A(n7474), .ZN(n5077) );
  NAND2_X1 U5384 ( .A1(n4914), .A2(n10212), .ZN(n10203) );
  INV_X1 U5385 ( .A(n10201), .ZN(n4914) );
  NOR2_X1 U5386 ( .A1(n6874), .A2(n5069), .ZN(n5068) );
  INV_X1 U5387 ( .A(n8282), .ZN(n5069) );
  AND2_X1 U5388 ( .A1(n8279), .A2(n8282), .ZN(n8202) );
  NAND2_X1 U5389 ( .A1(n8064), .A2(n6792), .ZN(n8266) );
  NAND2_X1 U5390 ( .A1(n8266), .A2(n8273), .ZN(n6783) );
  NAND2_X1 U5391 ( .A1(n8175), .A2(n8174), .ZN(n8739) );
  INV_X1 U5392 ( .A(n4898), .ZN(n4897) );
  OAI21_X1 U5393 ( .B1(n4899), .B2(n4902), .A(n4903), .ZN(n4898) );
  NAND2_X1 U5394 ( .A1(n4904), .A2(n8586), .ZN(n4903) );
  NAND2_X1 U5395 ( .A1(n4901), .A2(n4900), .ZN(n4899) );
  NAND2_X1 U5396 ( .A1(n8623), .A2(n4902), .ZN(n4900) );
  NOR2_X1 U5397 ( .A1(n8833), .A2(n8410), .ZN(n4905) );
  INV_X1 U5398 ( .A(n8613), .ZN(n8623) );
  NOR2_X1 U5399 ( .A1(n8622), .A2(n8623), .ZN(n8621) );
  NAND2_X1 U5400 ( .A1(n5732), .A2(n5731), .ZN(n8760) );
  NOR2_X1 U5401 ( .A1(n7635), .A2(n4890), .ZN(n4889) );
  INV_X1 U5402 ( .A(n4497), .ZN(n4890) );
  NAND2_X1 U5403 ( .A1(n4887), .A2(n4891), .ZN(n4886) );
  INV_X1 U5404 ( .A(n8685), .ZN(n4887) );
  AOI21_X1 U5405 ( .B1(n4490), .B2(n8321), .A(n4528), .ZN(n4917) );
  OAI211_X2 U5406 ( .C1(n6411), .C2(n5295), .A(n5221), .B(n5220), .ZN(n6287)
         );
  AND2_X1 U5407 ( .A1(n5588), .A2(n8400), .ZN(n8803) );
  AND2_X1 U5408 ( .A1(n10435), .A2(n6872), .ZN(n10466) );
  NAND2_X1 U5409 ( .A1(n5203), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5204) );
  NAND2_X1 U5410 ( .A1(n5151), .A2(n5150), .ZN(n5200) );
  NOR2_X1 U5411 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n5018) );
  NAND2_X1 U5412 ( .A1(n5173), .A2(n5175), .ZN(n5171) );
  NAND2_X1 U5413 ( .A1(n4669), .A2(n10413), .ZN(n4668) );
  NAND2_X1 U5414 ( .A1(n4680), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4669) );
  INV_X1 U5415 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n4680) );
  OR2_X1 U5416 ( .A1(n7704), .A2(n7703), .ZN(n4813) );
  XNOR2_X1 U5417 ( .A(n6544), .B(n6576), .ZN(n6548) );
  AOI21_X1 U5418 ( .B1(n4808), .B2(n4810), .A(n4514), .ZN(n4806) );
  NAND2_X1 U5419 ( .A1(n7705), .A2(n4808), .ZN(n4807) );
  NAND2_X1 U5420 ( .A1(n4784), .A2(n7874), .ZN(n8899) );
  NAND2_X1 U5421 ( .A1(n4782), .A2(n8998), .ZN(n4784) );
  INV_X1 U5422 ( .A(n7272), .ZN(n4781) );
  NAND2_X1 U5423 ( .A1(n4778), .A2(n4777), .ZN(n6686) );
  AOI21_X1 U5424 ( .B1(n8879), .B2(n7984), .A(n7953), .ZN(n9415) );
  AND2_X1 U5425 ( .A1(n7913), .A2(n7912), .ZN(n9027) );
  NAND2_X1 U5426 ( .A1(n4827), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n4826) );
  INV_X1 U5427 ( .A(n5947), .ZN(n4756) );
  NAND2_X1 U5428 ( .A1(n6105), .A2(n6106), .ZN(n6104) );
  NOR2_X1 U5429 ( .A1(n7051), .A2(n4764), .ZN(n7250) );
  AND2_X1 U5430 ( .A1(n7373), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4764) );
  OR2_X1 U5431 ( .A1(n7053), .A2(n7054), .ZN(n7248) );
  OR2_X1 U5432 ( .A1(n7441), .A2(n7440), .ZN(n4763) );
  NOR2_X1 U5433 ( .A1(n9452), .A2(n9661), .ZN(n4693) );
  INV_X1 U5434 ( .A(n4693), .ZN(n9435) );
  INV_X1 U5435 ( .A(n4638), .ZN(n4635) );
  NAND2_X1 U5436 ( .A1(n4640), .A2(n4489), .ZN(n4639) );
  AND2_X1 U5437 ( .A1(n9241), .A2(n9427), .ZN(n9448) );
  AND2_X1 U5438 ( .A1(n7972), .A2(n7971), .ZN(n9430) );
  OAI21_X1 U5439 ( .B1(n9069), .B2(n4856), .A(n9268), .ZN(n4850) );
  OR2_X1 U5440 ( .A1(n9681), .A2(n9027), .ZN(n9467) );
  NAND2_X1 U5441 ( .A1(n9467), .A2(n9231), .ZN(n9478) );
  NOR2_X1 U5442 ( .A1(n8037), .A2(n4518), .ZN(n4648) );
  AOI21_X1 U5443 ( .B1(n4487), .B2(n4837), .A(n4521), .ZN(n4830) );
  NOR2_X1 U5444 ( .A1(n9064), .A2(n9065), .ZN(n9500) );
  AND2_X1 U5445 ( .A1(n7861), .A2(n7860), .ZN(n8049) );
  INV_X1 U5446 ( .A(n4836), .ZN(n4835) );
  OAI21_X1 U5447 ( .B1(n9538), .B2(n4837), .A(n9062), .ZN(n4836) );
  NAND2_X1 U5448 ( .A1(n8036), .A2(n4550), .ZN(n9506) );
  OR2_X1 U5449 ( .A1(n9693), .A2(n9540), .ZN(n8035) );
  NAND2_X1 U5450 ( .A1(n9537), .A2(n9538), .ZN(n9536) );
  NOR2_X1 U5451 ( .A1(n9534), .A2(n9693), .ZN(n9521) );
  INV_X1 U5452 ( .A(n4628), .ZN(n4626) );
  AND2_X1 U5453 ( .A1(n4625), .A2(n4977), .ZN(n4624) );
  OR2_X1 U5454 ( .A1(n4533), .A2(n4978), .ZN(n4977) );
  NAND2_X1 U5455 ( .A1(n4628), .A2(n4631), .ZN(n4625) );
  INV_X1 U5456 ( .A(n4985), .ZN(n4978) );
  INV_X1 U5457 ( .A(n9707), .ZN(n9554) );
  NOR2_X1 U5458 ( .A1(n4984), .A2(n8033), .ZN(n4983) );
  INV_X1 U5459 ( .A(n9591), .ZN(n4984) );
  AOI21_X1 U5460 ( .B1(n4982), .B2(n4503), .A(n4981), .ZN(n4980) );
  INV_X1 U5461 ( .A(n8033), .ZN(n4982) );
  NOR2_X1 U5462 ( .A1(n9580), .A2(n9564), .ZN(n4981) );
  NAND2_X1 U5463 ( .A1(n4627), .A2(n4630), .ZN(n9583) );
  OR2_X1 U5464 ( .A1(n9598), .A2(n8032), .ZN(n4627) );
  OR2_X1 U5465 ( .A1(n7419), .A2(n7418), .ZN(n7730) );
  OR2_X1 U5466 ( .A1(n9731), .A2(n9621), .ZN(n9614) );
  NAND2_X1 U5467 ( .A1(n4659), .A2(n4665), .ZN(n4657) );
  NAND2_X1 U5468 ( .A1(n8030), .A2(n4661), .ZN(n4656) );
  NOR2_X1 U5469 ( .A1(n9637), .A2(n4662), .ZN(n4661) );
  INV_X1 U5470 ( .A(n8031), .ZN(n4662) );
  NAND2_X1 U5471 ( .A1(n4664), .A2(n4666), .ZN(n4663) );
  INV_X1 U5472 ( .A(n8030), .ZN(n4664) );
  NOR2_X1 U5473 ( .A1(n9644), .A2(n9731), .ZN(n9645) );
  AND2_X1 U5474 ( .A1(n9614), .A2(n9181), .ZN(n9637) );
  NAND2_X1 U5475 ( .A1(n4976), .A2(n9154), .ZN(n7302) );
  INV_X1 U5476 ( .A(n7188), .ZN(n4976) );
  AND2_X1 U5477 ( .A1(n9289), .A2(n4975), .ZN(n4974) );
  NAND2_X1 U5478 ( .A1(n9287), .A2(n7301), .ZN(n4975) );
  NAND2_X1 U5479 ( .A1(n7188), .A2(n7301), .ZN(n4970) );
  AND2_X1 U5480 ( .A1(n9281), .A2(n6854), .ZN(n4998) );
  NAND2_X1 U5481 ( .A1(n6721), .A2(n9280), .ZN(n6855) );
  OAI211_X1 U5482 ( .C1(n6842), .C2(n6586), .A(n6585), .B(n6584), .ZN(n6707)
         );
  NOR2_X1 U5483 ( .A1(n4501), .A2(n4995), .ZN(n4994) );
  INV_X1 U5484 ( .A(n6458), .ZN(n4995) );
  NAND2_X1 U5485 ( .A1(n4614), .A2(n5974), .ZN(n4613) );
  INV_X1 U5486 ( .A(n10254), .ZN(n10350) );
  AND2_X1 U5487 ( .A1(n9264), .A2(n8071), .ZN(n10254) );
  NAND2_X1 U5488 ( .A1(n7749), .A2(n7748), .ZN(n9720) );
  OR2_X1 U5489 ( .A1(n6715), .A2(n6411), .ZN(n6412) );
  AND2_X1 U5490 ( .A1(n6337), .A2(n6336), .ZN(n10372) );
  AND2_X1 U5491 ( .A1(n4989), .A2(n4540), .ZN(n4987) );
  XNOR2_X1 U5492 ( .A(n8181), .B(n8180), .ZN(n8184) );
  XNOR2_X1 U5493 ( .A(n7505), .B(n7504), .ZN(n7902) );
  NAND2_X1 U5494 ( .A1(n5113), .A2(n4694), .ZN(n4986) );
  INV_X1 U5495 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5108) );
  NAND2_X1 U5496 ( .A1(n4925), .A2(n5662), .ZN(n5683) );
  NAND2_X1 U5497 ( .A1(n5648), .A2(n4929), .ZN(n4925) );
  NAND2_X1 U5498 ( .A1(n5648), .A2(n5647), .ZN(n5664) );
  INV_X1 U5499 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n6361) );
  XNOR2_X1 U5500 ( .A(n5386), .B(n5385), .ZN(n7001) );
  XNOR2_X1 U5501 ( .A(n5198), .B(n5197), .ZN(n5293) );
  OAI21_X1 U5502 ( .B1(n7590), .B2(n4715), .A(n4714), .ZN(n4713) );
  INV_X1 U5503 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n4715) );
  NAND2_X1 U5504 ( .A1(n7590), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4714) );
  AOI21_X1 U5505 ( .B1(n4604), .B2(n4602), .A(n4530), .ZN(n4601) );
  INV_X1 U5506 ( .A(n4608), .ZN(n4602) );
  INV_X1 U5507 ( .A(n4604), .ZN(n4603) );
  INV_X1 U5508 ( .A(n8416), .ZN(n7400) );
  AOI21_X1 U5509 ( .B1(n5006), .B2(n5089), .A(n5002), .ZN(n5001) );
  NAND2_X1 U5510 ( .A1(n5003), .A2(n8022), .ZN(n5002) );
  NAND2_X1 U5511 ( .A1(n5012), .A2(n8021), .ZN(n5005) );
  NOR2_X1 U5512 ( .A1(n5291), .A2(n6217), .ZN(n4586) );
  NAND2_X1 U5513 ( .A1(n5366), .A2(n5365), .ZN(n8116) );
  INV_X1 U5514 ( .A(n8167), .ZN(n8137) );
  NAND2_X1 U5515 ( .A1(n5213), .A2(n8517), .ZN(n8400) );
  NOR2_X1 U5516 ( .A1(n5847), .A2(n5846), .ZN(n5878) );
  NAND2_X1 U5517 ( .A1(n8553), .A2(n8552), .ZN(n8737) );
  OAI21_X1 U5518 ( .B1(n8547), .B2(n8546), .A(n10432), .ZN(n8553) );
  NAND2_X1 U5519 ( .A1(n6868), .A2(n6867), .ZN(n6870) );
  NAND2_X1 U5520 ( .A1(n8191), .A2(n8190), .ZN(n8810) );
  NAND2_X1 U5522 ( .A1(n7946), .A2(n8189), .ZN(n7651) );
  NAND2_X1 U5523 ( .A1(n6803), .A2(n6804), .ZN(n8975) );
  NAND2_X1 U5524 ( .A1(n6686), .A2(n6559), .ZN(n6803) );
  INV_X1 U5525 ( .A(n8874), .ZN(n4814) );
  NAND2_X1 U5526 ( .A1(n8877), .A2(n8875), .ZN(n4815) );
  NAND2_X1 U5527 ( .A1(n7960), .A2(n7959), .ZN(n9664) );
  NAND2_X1 U5528 ( .A1(n5044), .A2(n4545), .ZN(n5043) );
  INV_X1 U5529 ( .A(n6548), .ZN(n6676) );
  NAND2_X1 U5530 ( .A1(n7727), .A2(n7726), .ZN(n9728) );
  OAI211_X2 U5531 ( .C1(n6842), .C2(n6304), .A(n6303), .B(n6302), .ZN(n6690)
         );
  OR2_X1 U5532 ( .A1(n9463), .A2(n7929), .ZN(n7935) );
  AND2_X1 U5533 ( .A1(n5989), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n4772) );
  AND2_X1 U5534 ( .A1(n5943), .A2(n5899), .ZN(n10332) );
  OAI21_X1 U5535 ( .B1(n10337), .B2(n9404), .A(n9403), .ZN(n4770) );
  NAND2_X1 U5536 ( .A1(n9769), .A2(n6840), .ZN(n9117) );
  XNOR2_X1 U5537 ( .A(n4691), .B(n9655), .ZN(n9657) );
  NAND2_X1 U5538 ( .A1(n4693), .A2(n4692), .ZN(n4691) );
  INV_X1 U5539 ( .A(n10267), .ZN(n4692) );
  NAND2_X1 U5540 ( .A1(n9112), .A2(n9111), .ZN(n10267) );
  XNOR2_X1 U5541 ( .A(n10267), .B(n9435), .ZN(n10264) );
  NAND2_X1 U5542 ( .A1(n9662), .A2(n4653), .ZN(n9745) );
  NOR2_X1 U5543 ( .A1(n4654), .A2(n4493), .ZN(n4653) );
  AND2_X1 U5544 ( .A1(n6618), .A2(n5782), .ZN(n9762) );
  XNOR2_X1 U5545 ( .A(n5119), .B(n9967), .ZN(n9263) );
  NAND2_X1 U5546 ( .A1(n6121), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6118) );
  OAI211_X1 U5547 ( .C1(n9135), .C2(n9256), .A(n9139), .B(n4569), .ZN(n9149)
         );
  OR2_X1 U5548 ( .A1(n9134), .A2(n9251), .ZN(n4569) );
  NOR2_X1 U5549 ( .A1(n4737), .A2(n4736), .ZN(n4735) );
  INV_X1 U5550 ( .A(n8378), .ZN(n4736) );
  INV_X1 U5551 ( .A(n8376), .ZN(n4737) );
  NOR2_X1 U5552 ( .A1(n4596), .A2(n5021), .ZN(n4595) );
  INV_X1 U5553 ( .A(n5449), .ZN(n4596) );
  AOI21_X1 U5554 ( .B1(n4795), .B2(n4798), .A(n4794), .ZN(n4793) );
  INV_X1 U5555 ( .A(n8916), .ZN(n4794) );
  OR2_X1 U5556 ( .A1(n9246), .A2(n9256), .ZN(n5091) );
  AND2_X1 U5557 ( .A1(n4866), .A2(n9166), .ZN(n4864) );
  INV_X1 U5558 ( .A(n7301), .ZN(n4972) );
  NAND2_X1 U5559 ( .A1(n7138), .A2(n4620), .ZN(n4619) );
  INV_X1 U5560 ( .A(n4620), .ZN(n4618) );
  NOR2_X1 U5561 ( .A1(n4936), .A2(n4933), .ZN(n4932) );
  INV_X1 U5562 ( .A(n7585), .ZN(n4936) );
  INV_X1 U5563 ( .A(n7568), .ZN(n4933) );
  INV_X1 U5564 ( .A(n7570), .ZN(n4935) );
  AND2_X1 U5565 ( .A1(n4963), .A2(n5755), .ZN(n4962) );
  NAND2_X1 U5566 ( .A1(n5724), .A2(n5726), .ZN(n4963) );
  INV_X1 U5567 ( .A(n5726), .ZN(n4960) );
  INV_X1 U5568 ( .A(n4927), .ZN(n4926) );
  OAI21_X1 U5569 ( .B1(n4929), .B2(n4928), .A(n5682), .ZN(n4927) );
  INV_X1 U5570 ( .A(n5662), .ZN(n4928) );
  NAND2_X1 U5571 ( .A1(n5537), .A2(n5539), .ZN(n4957) );
  INV_X1 U5572 ( .A(n5557), .ZN(n4953) );
  INV_X1 U5573 ( .A(n5539), .ZN(n4954) );
  AND2_X1 U5574 ( .A1(n5472), .A2(n5474), .ZN(n5476) );
  NAND2_X1 U5575 ( .A1(n5480), .A2(n5481), .ZN(n4965) );
  AND2_X1 U5576 ( .A1(n5428), .A2(n5427), .ZN(n5473) );
  INV_X1 U5577 ( .A(P1_RD_REG_SCAN_IN), .ZN(n5177) );
  INV_X1 U5578 ( .A(n8015), .ZN(n5009) );
  AND2_X1 U5579 ( .A1(n7081), .A2(n5448), .ZN(n5449) );
  INV_X1 U5580 ( .A(n8100), .ZN(n5038) );
  OR2_X1 U5581 ( .A1(n5498), .A2(n5497), .ZN(n5499) );
  NAND2_X1 U5582 ( .A1(n4532), .A2(n4728), .ZN(n4727) );
  OR2_X1 U5583 ( .A1(n5463), .A2(n7222), .ZN(n5487) );
  OR2_X1 U5584 ( .A1(n8739), .A2(n8177), .ZN(n8385) );
  OR2_X1 U5585 ( .A1(n5369), .A2(n5368), .ZN(n5395) );
  INV_X1 U5586 ( .A(n8286), .ZN(n6869) );
  OR2_X1 U5587 ( .A1(n6047), .A2(n10465), .ZN(n6764) );
  OAI21_X1 U5588 ( .B1(n4897), .B2(n8582), .A(n4529), .ZN(n4894) );
  INV_X1 U5589 ( .A(n4899), .ZN(n4896) );
  INV_X1 U5590 ( .A(n4905), .ZN(n4902) );
  OR2_X1 U5591 ( .A1(n8662), .A2(n8639), .ZN(n8342) );
  NAND2_X1 U5592 ( .A1(n7487), .A2(n7518), .ZN(n7546) );
  NAND2_X1 U5593 ( .A1(n5080), .A2(n8307), .ZN(n10213) );
  AND2_X1 U5594 ( .A1(n8306), .A2(n8243), .ZN(n8207) );
  NAND2_X1 U5595 ( .A1(n5150), .A2(n5087), .ZN(n5086) );
  INV_X1 U5596 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5087) );
  AOI21_X1 U5597 ( .B1(n8908), .B2(n8907), .A(n4801), .ZN(n4800) );
  INV_X1 U5598 ( .A(n8987), .ZN(n4801) );
  NAND2_X1 U5599 ( .A1(n4809), .A2(n7710), .ZN(n4803) );
  INV_X1 U5600 ( .A(n4813), .ZN(n4809) );
  NAND2_X1 U5601 ( .A1(n9267), .A2(n9250), .ZN(n9302) );
  INV_X1 U5602 ( .A(n9270), .ZN(n4831) );
  NAND2_X1 U5603 ( .A1(n9554), .A2(n9572), .ZN(n4985) );
  NAND2_X1 U5604 ( .A1(n9580), .A2(n4703), .ZN(n4702) );
  NAND2_X1 U5605 ( .A1(n4701), .A2(n9554), .ZN(n4700) );
  INV_X1 U5606 ( .A(n4702), .ZN(n4701) );
  INV_X1 U5607 ( .A(n9618), .ZN(n4665) );
  INV_X1 U5608 ( .A(n4864), .ZN(n4858) );
  AND2_X1 U5609 ( .A1(n4862), .A2(n4536), .ZN(n4860) );
  NAND2_X1 U5610 ( .A1(n7417), .A2(n4864), .ZN(n4861) );
  OR2_X1 U5611 ( .A1(n7289), .A2(n7288), .ZN(n7383) );
  NOR2_X1 U5612 ( .A1(n7407), .A2(n7300), .ZN(n4712) );
  INV_X1 U5613 ( .A(n7017), .ZN(n7015) );
  OR2_X1 U5614 ( .A1(n6935), .A2(n6934), .ZN(n7017) );
  NAND2_X1 U5615 ( .A1(n6839), .A2(n4846), .ZN(n4845) );
  NAND2_X1 U5616 ( .A1(n7417), .A2(n9166), .ZN(n10249) );
  INV_X1 U5617 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5125) );
  AND2_X1 U5618 ( .A1(n7526), .A2(n7508), .ZN(n7524) );
  OAI21_X1 U5619 ( .B1(n5725), .B2(n4961), .A(n4958), .ZN(n7448) );
  AOI21_X1 U5620 ( .B1(n4962), .B2(n4960), .A(n4959), .ZN(n4958) );
  INV_X1 U5621 ( .A(n4962), .ZN(n4961) );
  INV_X1 U5622 ( .A(n5757), .ZN(n4959) );
  OAI21_X1 U5623 ( .B1(n6121), .B2(P1_IR_REG_20__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5122) );
  NOR2_X1 U5624 ( .A1(n5663), .A2(n4930), .ZN(n4929) );
  INV_X1 U5625 ( .A(n5647), .ZN(n4930) );
  NAND2_X1 U5626 ( .A1(n5645), .A2(n5644), .ZN(n5648) );
  NAND2_X1 U5627 ( .A1(n5506), .A2(n10114), .ZN(n5539) );
  AND2_X1 U5628 ( .A1(n5557), .A2(n5544), .ZN(n5555) );
  XNOR2_X1 U5629 ( .A(n5501), .B(n10068), .ZN(n5500) );
  AND2_X1 U5630 ( .A1(n5481), .A2(n5458), .ZN(n5470) );
  NAND2_X1 U5631 ( .A1(n5478), .A2(n5433), .ZN(n5471) );
  AOI21_X1 U5632 ( .B1(n4743), .B2(n4741), .A(n4531), .ZN(n4740) );
  INV_X1 U5633 ( .A(n4743), .ZN(n4742) );
  INV_X1 U5634 ( .A(n5360), .ZN(n4741) );
  AND2_X1 U5635 ( .A1(n4744), .A2(n5381), .ZN(n4743) );
  NAND2_X1 U5636 ( .A1(n5358), .A2(n5360), .ZN(n4744) );
  XNOR2_X1 U5637 ( .A(n5334), .B(SI_7_), .ZN(n5331) );
  NAND2_X1 U5638 ( .A1(n4939), .A2(n4938), .ZN(n5333) );
  AOI21_X1 U5639 ( .B1(n4941), .B2(n4943), .A(n4526), .ZN(n4938) );
  OAI21_X1 U5640 ( .B1(n7590), .B2(n4572), .A(n4571), .ZN(n5198) );
  NAND2_X1 U5641 ( .A1(n7590), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n4571) );
  AND2_X1 U5642 ( .A1(n5192), .A2(n5188), .ZN(n4724) );
  NAND2_X1 U5643 ( .A1(n4581), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n4580) );
  INV_X1 U5644 ( .A(n6143), .ZN(n4581) );
  NOR2_X1 U5645 ( .A1(n5322), .A2(n5321), .ZN(n5347) );
  INV_X1 U5646 ( .A(n8076), .ZN(n4607) );
  AOI21_X1 U5647 ( .B1(n8072), .B2(n8157), .A(n8156), .ZN(n4608) );
  NAND2_X1 U5648 ( .A1(n5012), .A2(n5004), .ZN(n5003) );
  NOR2_X1 U5649 ( .A1(n5011), .A2(n8015), .ZN(n5004) );
  NAND2_X1 U5650 ( .A1(n8110), .A2(n5376), .ZN(n8109) );
  NOR2_X1 U5651 ( .A1(n5395), .A2(n10062), .ZN(n5412) );
  NAND2_X1 U5652 ( .A1(n5029), .A2(n5032), .ZN(n5028) );
  AOI21_X1 U5653 ( .B1(n5031), .B2(n5030), .A(n5423), .ZN(n5029) );
  XNOR2_X1 U5654 ( .A(n5263), .B(n6287), .ZN(n6229) );
  INV_X1 U5655 ( .A(n8400), .ZN(n5600) );
  NAND2_X1 U5656 ( .A1(n4718), .A2(n5213), .ZN(n4717) );
  NAND2_X1 U5657 ( .A1(n8399), .A2(n5212), .ZN(n4718) );
  OR3_X1 U5658 ( .A1(n7367), .A2(n7513), .A3(n7458), .ZN(n5598) );
  INV_X1 U5659 ( .A(n7667), .ZN(n7625) );
  NOR2_X1 U5660 ( .A1(n7216), .A2(n4558), .ZN(n8448) );
  NAND2_X1 U5661 ( .A1(n8448), .A2(n8447), .ZN(n8446) );
  NAND2_X1 U5662 ( .A1(n8446), .A2(n4681), .ZN(n7219) );
  OR2_X1 U5663 ( .A1(n8440), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n4681) );
  NAND2_X1 U5664 ( .A1(n7219), .A2(n7220), .ZN(n7352) );
  NOR2_X1 U5665 ( .A1(n8457), .A2(n8456), .ZN(n8459) );
  XNOR2_X1 U5666 ( .A(n4688), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8515) );
  NAND2_X1 U5667 ( .A1(n8511), .A2(n4566), .ZN(n4688) );
  NAND2_X1 U5668 ( .A1(n4584), .A2(n4583), .ZN(n8530) );
  NAND2_X1 U5669 ( .A1(n5619), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5713) );
  NOR2_X1 U5670 ( .A1(n8783), .A2(n4875), .ZN(n4873) );
  INV_X1 U5671 ( .A(n5604), .ZN(n5603) );
  OR2_X1 U5672 ( .A1(n5564), .A2(n8478), .ZN(n5604) );
  NAND2_X1 U5673 ( .A1(n7487), .A2(n4877), .ZN(n7574) );
  NAND2_X1 U5674 ( .A1(n5514), .A2(n5513), .ZN(n8804) );
  AND2_X1 U5675 ( .A1(n8318), .A2(n8319), .ZN(n8317) );
  INV_X1 U5676 ( .A(n4908), .ZN(n4907) );
  OAI21_X1 U5677 ( .B1(n10212), .B2(n4909), .A(n4911), .ZN(n4908) );
  INV_X1 U5678 ( .A(n8317), .ZN(n8210) );
  NAND2_X1 U5679 ( .A1(n5080), .A2(n5078), .ZN(n10215) );
  AND2_X1 U5680 ( .A1(n8307), .A2(n8309), .ZN(n8208) );
  OAI21_X1 U5681 ( .B1(n10425), .B2(n5064), .A(n5060), .ZN(n5066) );
  NAND2_X1 U5682 ( .A1(n5065), .A2(n8292), .ZN(n5064) );
  NAND2_X1 U5683 ( .A1(n10424), .A2(n8292), .ZN(n7164) );
  NAND2_X1 U5684 ( .A1(n4872), .A2(n4871), .ZN(n7161) );
  INV_X1 U5685 ( .A(n10419), .ZN(n4872) );
  NAND2_X1 U5686 ( .A1(n10420), .A2(n10489), .ZN(n10419) );
  NAND2_X1 U5687 ( .A1(n10425), .A2(n10426), .ZN(n10424) );
  AND2_X1 U5688 ( .A1(n8203), .A2(n8274), .ZN(n5070) );
  NAND2_X1 U5689 ( .A1(n5071), .A2(n8274), .ZN(n6497) );
  AND2_X1 U5690 ( .A1(n8250), .A2(n6048), .ZN(n6051) );
  NAND2_X1 U5691 ( .A1(n6051), .A2(n6050), .ZN(n6284) );
  NAND2_X1 U5692 ( .A1(n6764), .A2(n8256), .ZN(n8250) );
  NAND2_X1 U5693 ( .A1(n8378), .A2(n8227), .ZN(n8535) );
  INV_X1 U5694 ( .A(n4885), .ZN(n4884) );
  OAI21_X1 U5695 ( .B1(n4886), .B2(n4504), .A(n7636), .ZN(n4885) );
  AND2_X1 U5696 ( .A1(n8333), .A2(n8683), .ZN(n8699) );
  NAND2_X1 U5697 ( .A1(n5563), .A2(n5562), .ZN(n8794) );
  OR2_X1 U5698 ( .A1(n5295), .A2(n6398), .ZN(n5282) );
  OR2_X1 U5699 ( .A1(n10472), .A2(n8517), .ZN(n6769) );
  NOR2_X1 U5700 ( .A1(n7513), .A2(n5573), .ZN(n10457) );
  AND2_X1 U5701 ( .A1(n7458), .A2(n5572), .ZN(n5573) );
  NOR2_X1 U5702 ( .A1(n5086), .A2(P2_IR_REG_28__SCAN_IN), .ZN(n5085) );
  INV_X1 U5703 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5083) );
  AND2_X1 U5704 ( .A1(n5218), .A2(n5154), .ZN(n5081) );
  INV_X1 U5705 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n4610) );
  AND3_X1 U5706 ( .A1(n5136), .A2(n5218), .A3(n5135), .ZN(n5147) );
  NAND2_X1 U5707 ( .A1(n8865), .A2(P2_IR_REG_1__SCAN_IN), .ZN(n4679) );
  AOI21_X1 U5708 ( .B1(n4800), .B2(n4797), .A(n4796), .ZN(n4795) );
  INV_X1 U5709 ( .A(n8988), .ZN(n4796) );
  INV_X1 U5710 ( .A(n4800), .ZN(n4798) );
  AND2_X1 U5711 ( .A1(n7745), .A2(n7723), .ZN(n5054) );
  AND2_X1 U5712 ( .A1(n7900), .A2(n4787), .ZN(n4786) );
  NAND2_X1 U5713 ( .A1(n4789), .A2(n4783), .ZN(n4785) );
  OR2_X1 U5714 ( .A1(n7873), .A2(n4788), .ZN(n4787) );
  AND2_X1 U5715 ( .A1(n7894), .A2(n7893), .ZN(n7896) );
  OR2_X1 U5716 ( .A1(n9497), .A2(n4484), .ZN(n7894) );
  NAND2_X1 U5717 ( .A1(n6727), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n6846) );
  INV_X1 U5718 ( .A(n6729), .ZN(n6727) );
  INV_X1 U5719 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n6845) );
  AOI21_X1 U5720 ( .B1(n6566), .B2(n9359), .A(n6147), .ZN(n6153) );
  NAND2_X1 U5721 ( .A1(n6152), .A2(n6151), .ZN(n6538) );
  NOR2_X1 U5722 ( .A1(n7330), .A2(n5058), .ZN(n5057) );
  INV_X1 U5723 ( .A(n7326), .ZN(n5058) );
  NAND2_X1 U5724 ( .A1(n7769), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n7789) );
  INV_X1 U5725 ( .A(n7771), .ZN(n7769) );
  NAND2_X1 U5726 ( .A1(n6465), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n6606) );
  NAND2_X1 U5727 ( .A1(n4804), .A2(n4802), .ZN(n4808) );
  NAND2_X1 U5728 ( .A1(n4499), .A2(n4805), .ZN(n4804) );
  NAND2_X1 U5729 ( .A1(n4803), .A2(n4509), .ZN(n4802) );
  AND2_X1 U5730 ( .A1(n4813), .A2(n4509), .ZN(n4805) );
  INV_X1 U5731 ( .A(n4811), .ZN(n4810) );
  AOI21_X1 U5732 ( .B1(n4499), .B2(n4813), .A(n4812), .ZN(n4811) );
  NAND2_X1 U5733 ( .A1(n9264), .A2(n4485), .ZN(n4949) );
  INV_X1 U5734 ( .A(n9266), .ZN(n4950) );
  NAND2_X1 U5735 ( .A1(n9266), .A2(n9265), .ZN(n4947) );
  AND2_X1 U5736 ( .A1(n4921), .A2(n9111), .ZN(n4920) );
  NAND2_X1 U5737 ( .A1(n9655), .A2(n9407), .ZN(n9267) );
  INV_X1 U5738 ( .A(n7984), .ZN(n7929) );
  NAND2_X1 U5739 ( .A1(n6064), .A2(n6154), .ZN(n6063) );
  OAI21_X1 U5740 ( .B1(n5985), .B2(n5984), .A(n5987), .ZN(n4774) );
  NOR2_X1 U5741 ( .A1(n4774), .A2(n4773), .ZN(n6091) );
  INV_X1 U5742 ( .A(n6094), .ZN(n4773) );
  AOI21_X1 U5743 ( .B1(n5994), .B2(n4760), .A(n4547), .ZN(n4759) );
  INV_X1 U5744 ( .A(n5992), .ZN(n4760) );
  OR2_X1 U5745 ( .A1(n5991), .A2(n4761), .ZN(n4758) );
  INV_X1 U5746 ( .A(n5994), .ZN(n4761) );
  NOR2_X1 U5747 ( .A1(n6445), .A2(n4765), .ZN(n6448) );
  AND2_X1 U5748 ( .A1(n7283), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n4765) );
  NOR2_X1 U5749 ( .A1(n6448), .A2(n6447), .ZN(n7051) );
  AND2_X1 U5750 ( .A1(n4763), .A2(n4762), .ZN(n9363) );
  NAND2_X1 U5751 ( .A1(n9366), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n4762) );
  NOR2_X1 U5752 ( .A1(n9363), .A2(n9362), .ZN(n9382) );
  NAND2_X1 U5753 ( .A1(n9053), .A2(n9052), .ZN(n9661) );
  INV_X1 U5754 ( .A(n4868), .ZN(n4867) );
  NAND2_X1 U5755 ( .A1(n4870), .A2(n10355), .ZN(n4869) );
  OAI22_X1 U5756 ( .A1(n9430), .A2(n10352), .B1(n9432), .B2(n9431), .ZN(n4868)
         );
  NOR2_X1 U5757 ( .A1(n4489), .A2(n9422), .ZN(n4636) );
  NOR2_X1 U5758 ( .A1(n5090), .A2(n4527), .ZN(n4638) );
  NAND2_X1 U5759 ( .A1(n4489), .A2(n9422), .ZN(n4633) );
  AND2_X1 U5760 ( .A1(n7966), .A2(n9433), .ZN(n9455) );
  NOR2_X1 U5761 ( .A1(n9671), .A2(n4705), .ZN(n4704) );
  INV_X1 U5762 ( .A(n4706), .ZN(n4705) );
  OR2_X1 U5763 ( .A1(n9454), .A2(n9664), .ZN(n9452) );
  INV_X1 U5764 ( .A(n4852), .ZN(n4851) );
  OAI21_X1 U5765 ( .B1(n9424), .B2(n4853), .A(n9423), .ZN(n4852) );
  AND2_X1 U5766 ( .A1(n9498), .A2(n4856), .ZN(n9469) );
  NAND2_X1 U5767 ( .A1(n9512), .A2(n4708), .ZN(n9482) );
  AND2_X1 U5768 ( .A1(n9269), .A2(n9268), .ZN(n9470) );
  INV_X1 U5769 ( .A(n4647), .ZN(n4646) );
  AND2_X1 U5770 ( .A1(n9521), .A2(n8049), .ZN(n9512) );
  NAND2_X1 U5771 ( .A1(n9512), .A2(n9497), .ZN(n9491) );
  INV_X1 U5772 ( .A(n7864), .ZN(n7862) );
  OR2_X1 U5773 ( .A1(n7845), .A2(n9003), .ZN(n7864) );
  NAND2_X1 U5774 ( .A1(n7805), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n7824) );
  INV_X1 U5775 ( .A(n7807), .ZN(n7805) );
  OR2_X1 U5776 ( .A1(n7789), .A2(n7788), .ZN(n7807) );
  NOR2_X1 U5777 ( .A1(n9599), .A2(n4702), .ZN(n9574) );
  AND4_X1 U5778 ( .A1(n7776), .A2(n7775), .A3(n7774), .A4(n7773), .ZN(n9573)
         );
  NOR2_X1 U5779 ( .A1(n9599), .A2(n9715), .ZN(n9584) );
  OR2_X1 U5780 ( .A1(n9623), .A2(n9720), .ZN(n9599) );
  NAND2_X1 U5781 ( .A1(n7728), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n7752) );
  AND2_X1 U5782 ( .A1(n9187), .A2(n9186), .ZN(n9618) );
  INV_X1 U5783 ( .A(n4865), .ZN(n9634) );
  OAI21_X1 U5784 ( .B1(n4859), .B2(n7417), .A(n4857), .ZN(n4865) );
  INV_X1 U5785 ( .A(n4860), .ZN(n4859) );
  AOI21_X1 U5786 ( .B1(n4860), .B2(n4858), .A(n9168), .ZN(n4857) );
  NAND2_X1 U5787 ( .A1(n4861), .A2(n4862), .ZN(n10246) );
  AND2_X1 U5788 ( .A1(n4861), .A2(n4860), .ZN(n8045) );
  NAND2_X1 U5789 ( .A1(n7202), .A2(n4710), .ZN(n9644) );
  AND2_X1 U5790 ( .A1(n4491), .A2(n4711), .ZN(n4710) );
  NAND2_X1 U5791 ( .A1(n7409), .A2(n9159), .ZN(n8030) );
  NAND2_X1 U5792 ( .A1(n7202), .A2(n4491), .ZN(n10243) );
  NAND2_X1 U5793 ( .A1(n7202), .A2(n4712), .ZN(n10242) );
  AND2_X1 U5794 ( .A1(n7202), .A2(n10281), .ZN(n7296) );
  NAND2_X1 U5795 ( .A1(n4841), .A2(n4839), .ZN(n7281) );
  AOI21_X1 U5796 ( .B1(n4842), .B2(n9147), .A(n4840), .ZN(n4839) );
  AOI21_X1 U5797 ( .B1(n4844), .B2(n4843), .A(n9150), .ZN(n4842) );
  OAI21_X1 U5798 ( .B1(n6721), .B2(n4997), .A(n4996), .ZN(n10338) );
  INV_X1 U5799 ( .A(n4998), .ZN(n4997) );
  AOI21_X1 U5800 ( .B1(n4998), .B2(n6726), .A(n4549), .ZN(n4996) );
  OR2_X1 U5801 ( .A1(n7145), .A2(n9350), .ZN(n4620) );
  OR2_X1 U5802 ( .A1(n10339), .A2(n7145), .ZN(n10340) );
  AND2_X1 U5803 ( .A1(n6844), .A2(n6843), .ZN(n6929) );
  NOR2_X1 U5804 ( .A1(n6704), .A2(n6707), .ZN(n6736) );
  AOI21_X1 U5805 ( .B1(n6725), .B2(n9312), .A(n9071), .ZN(n9136) );
  NAND2_X1 U5806 ( .A1(n5102), .A2(n5101), .ZN(n5118) );
  INV_X1 U5807 ( .A(n4524), .ZN(n4654) );
  NAND2_X1 U5808 ( .A1(n7844), .A2(n7843), .ZN(n9693) );
  NAND2_X1 U5809 ( .A1(n10358), .A2(n10375), .ZN(n10279) );
  INV_X1 U5810 ( .A(n6929), .ZN(n7136) );
  INV_X1 U5811 ( .A(n10372), .ZN(n10386) );
  XNOR2_X1 U5812 ( .A(n8184), .B(SI_30_), .ZN(n9110) );
  XNOR2_X1 U5813 ( .A(n7586), .B(n7585), .ZN(n7958) );
  NAND2_X1 U5814 ( .A1(n4937), .A2(n7570), .ZN(n7586) );
  NAND2_X1 U5815 ( .A1(n7569), .A2(n7568), .ZN(n4937) );
  XNOR2_X1 U5816 ( .A(n7569), .B(n7568), .ZN(n7946) );
  NAND2_X1 U5817 ( .A1(n5126), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5105) );
  AND2_X1 U5818 ( .A1(n5096), .A2(n4989), .ZN(n4817) );
  INV_X1 U5819 ( .A(n4986), .ZN(n4819) );
  NAND2_X1 U5820 ( .A1(n5120), .A2(n5056), .ZN(n6119) );
  OR2_X1 U5821 ( .A1(n5122), .A2(n5121), .ZN(n5056) );
  OAI21_X1 U5822 ( .B1(n5359), .B2(n5358), .A(n5360), .ZN(n5382) );
  XNOR2_X1 U5823 ( .A(n5312), .B(n10082), .ZN(n5310) );
  NOR2_X1 U5824 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5774) );
  NAND2_X1 U5825 ( .A1(n7172), .A2(n5495), .ZN(n7342) );
  AND2_X1 U5826 ( .A1(n8109), .A2(n5031), .ZN(n7105) );
  XOR2_X1 U5827 ( .A(n5552), .B(n5553), .Z(n7516) );
  CLKBUF_X1 U5828 ( .A(n7514), .Z(n7515) );
  XNOR2_X1 U5829 ( .A(n5292), .B(n6229), .ZN(n6217) );
  INV_X1 U5830 ( .A(n4587), .ZN(n6212) );
  AOI21_X1 U5831 ( .B1(n4511), .B2(n5017), .A(n5014), .ZN(n5013) );
  NAND2_X1 U5832 ( .A1(n5669), .A2(n5668), .ZN(n8775) );
  NOR2_X1 U5833 ( .A1(n5493), .A2(n4570), .ZN(n7173) );
  AND2_X1 U5834 ( .A1(n7337), .A2(n5469), .ZN(n4570) );
  NAND2_X1 U5835 ( .A1(n5251), .A2(n5252), .ZN(n5253) );
  NAND2_X1 U5836 ( .A1(n6229), .A2(n5292), .ZN(n5039) );
  AND2_X1 U5837 ( .A1(n7652), .A2(n7643), .ZN(n8590) );
  AND2_X1 U5838 ( .A1(n5601), .A2(n5600), .ZN(n10188) );
  AOI21_X1 U5839 ( .B1(n8529), .B2(n8178), .A(n8377), .ZN(n4574) );
  NAND2_X1 U5840 ( .A1(n4721), .A2(n4720), .ZN(n4719) );
  NAND2_X1 U5841 ( .A1(n8396), .A2(n8395), .ZN(n4720) );
  NAND2_X1 U5842 ( .A1(n8016), .A2(n5214), .ZN(n4582) );
  NAND2_X1 U5843 ( .A1(n5200), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5201) );
  NAND2_X1 U5844 ( .A1(n5834), .A2(n7700), .ZN(n4674) );
  INV_X1 U5845 ( .A(n4671), .ZN(n4670) );
  NOR2_X1 U5846 ( .A1(n8432), .A2(n4507), .ZN(n5870) );
  INV_X1 U5847 ( .A(n4687), .ZN(n5868) );
  AND2_X1 U5848 ( .A1(n4687), .A2(n4686), .ZN(n5847) );
  NAND2_X1 U5849 ( .A1(n5849), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n4686) );
  INV_X1 U5850 ( .A(n4685), .ZN(n5915) );
  INV_X1 U5851 ( .A(n4683), .ZN(n6163) );
  AND2_X1 U5852 ( .A1(n4683), .A2(n4682), .ZN(n6166) );
  NAND2_X1 U5853 ( .A1(n6168), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n4682) );
  NOR2_X1 U5854 ( .A1(n6343), .A2(n4690), .ZN(n6346) );
  AND2_X1 U5855 ( .A1(n6348), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n4690) );
  NOR2_X1 U5856 ( .A1(n6346), .A2(n6345), .ZN(n6645) );
  NOR2_X1 U5857 ( .A1(n6645), .A2(n4689), .ZN(n6648) );
  AND2_X1 U5858 ( .A1(n6650), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n4689) );
  NOR2_X1 U5859 ( .A1(n6648), .A2(n6647), .ZN(n7035) );
  XNOR2_X1 U5860 ( .A(n8454), .B(n8455), .ZN(n7557) );
  NOR2_X1 U5861 ( .A1(n7557), .A2(n7556), .ZN(n8456) );
  NAND2_X1 U5862 ( .A1(n5075), .A2(n8368), .ZN(n8568) );
  AND2_X1 U5863 ( .A1(n8620), .A2(n8619), .ZN(n8755) );
  NAND2_X1 U5864 ( .A1(n4919), .A2(n4490), .ZN(n7573) );
  AND2_X1 U5865 ( .A1(n4919), .A2(n4918), .ZN(n7540) );
  NAND2_X1 U5866 ( .A1(n10203), .A2(n4912), .ZN(n7464) );
  NAND2_X1 U5867 ( .A1(n10414), .A2(n6964), .ZN(n6965) );
  AND2_X1 U5868 ( .A1(n5067), .A2(n8284), .ZN(n6876) );
  NAND2_X1 U5869 ( .A1(n6818), .A2(n8282), .ZN(n6875) );
  OAI21_X1 U5870 ( .B1(n6461), .B2(n5295), .A(n5297), .ZN(n10444) );
  NAND2_X1 U5871 ( .A1(n10211), .A2(n10445), .ZN(n10439) );
  NAND2_X1 U5872 ( .A1(n6793), .A2(n8266), .ZN(n6483) );
  OR2_X1 U5873 ( .A1(n10458), .A2(n6769), .ZN(n10208) );
  INV_X1 U5874 ( .A(n8717), .ZN(n8723) );
  INV_X1 U5875 ( .A(n10439), .ZN(n10228) );
  AND2_X1 U5876 ( .A1(n8739), .A2(n8803), .ZN(n4573) );
  XOR2_X1 U5877 ( .A(n8535), .B(n8536), .Z(n8556) );
  OAI21_X1 U5878 ( .B1(n8622), .B2(n4899), .A(n4897), .ZN(n8581) );
  NOR2_X1 U5879 ( .A1(n8621), .A2(n4905), .ZN(n8600) );
  NAND2_X1 U5880 ( .A1(n5687), .A2(n5686), .ZN(n8843) );
  NAND2_X1 U5881 ( .A1(n4888), .A2(n4886), .ZN(n8665) );
  NAND2_X1 U5882 ( .A1(n7634), .A2(n4889), .ZN(n4888) );
  NAND2_X1 U5883 ( .A1(n7634), .A2(n4497), .ZN(n8681) );
  AND2_X1 U5884 ( .A1(n10496), .A2(n8803), .ZN(n8844) );
  NAND2_X1 U5885 ( .A1(n4678), .A2(n4679), .ZN(n6005) );
  NAND2_X1 U5886 ( .A1(n4821), .A2(n4565), .ZN(n6912) );
  OAI21_X1 U5887 ( .B1(n7705), .B2(n4499), .A(n4813), .ZN(n8889) );
  NAND2_X1 U5888 ( .A1(n7004), .A2(n7003), .ZN(n7183) );
  NAND2_X1 U5889 ( .A1(n7787), .A2(n7786), .ZN(n9712) );
  NAND2_X1 U5890 ( .A1(n4792), .A2(n4795), .ZN(n8917) );
  OR2_X1 U5891 ( .A1(n8910), .A2(n4798), .ZN(n4792) );
  NAND2_X1 U5892 ( .A1(n7327), .A2(n7326), .ZN(n7329) );
  NAND2_X1 U5893 ( .A1(n8898), .A2(n8901), .ZN(n7875) );
  AND2_X1 U5894 ( .A1(n8978), .A2(n8974), .ZN(n5053) );
  NOR2_X1 U5895 ( .A1(n6613), .A2(n6603), .ZN(n8977) );
  NAND2_X1 U5896 ( .A1(n4799), .A2(n8907), .ZN(n8990) );
  OR2_X1 U5897 ( .A1(n8910), .A2(n8908), .ZN(n4799) );
  NAND2_X1 U5898 ( .A1(n7804), .A2(n7803), .ZN(n9707) );
  NAND2_X1 U5899 ( .A1(n7269), .A2(n7268), .ZN(n7272) );
  NAND2_X1 U5900 ( .A1(n4780), .A2(n4779), .ZN(n6688) );
  NAND2_X1 U5901 ( .A1(n6558), .A2(n6559), .ZN(n6689) );
  INV_X1 U5902 ( .A(n9047), .ZN(n9019) );
  NAND2_X1 U5903 ( .A1(n7925), .A2(n7924), .ZN(n9674) );
  NAND2_X1 U5904 ( .A1(n7922), .A2(n6840), .ZN(n7925) );
  INV_X1 U5905 ( .A(n9019), .ZN(n9031) );
  NAND2_X1 U5906 ( .A1(n7716), .A2(n7715), .ZN(n9731) );
  INV_X1 U5907 ( .A(n9027), .ZN(n9501) );
  NAND2_X1 U5908 ( .A1(n6080), .A2(n6081), .ZN(n6079) );
  NAND2_X1 U5909 ( .A1(n6104), .A2(n5947), .ZN(n6080) );
  INV_X1 U5910 ( .A(n6081), .ZN(n4757) );
  AOI21_X1 U5911 ( .B1(n4756), .B2(n6081), .A(n4522), .ZN(n4755) );
  INV_X1 U5912 ( .A(n4774), .ZN(n6093) );
  NAND2_X1 U5913 ( .A1(n5991), .A2(n5992), .ZN(n5993) );
  XNOR2_X1 U5914 ( .A(n7250), .B(n7249), .ZN(n7053) );
  NOR2_X1 U5915 ( .A1(n7437), .A2(n4512), .ZN(n7441) );
  OAI211_X1 U5916 ( .C1(n4640), .C2(n4637), .A(n4634), .B(n4632), .ZN(n9658)
         );
  OR2_X1 U5917 ( .A1(n9461), .A2(n4633), .ZN(n4632) );
  NAND2_X1 U5918 ( .A1(n4638), .A2(n9428), .ZN(n4637) );
  OAI22_X1 U5919 ( .A1(n4636), .A2(n4635), .B1(n9422), .B2(n4638), .ZN(n4634)
         );
  AND2_X1 U5920 ( .A1(n4639), .A2(n4641), .ZN(n9451) );
  OAI21_X1 U5921 ( .B1(n9498), .B2(n9069), .A(n4849), .ZN(n9425) );
  INV_X1 U5922 ( .A(n4850), .ZN(n4849) );
  NAND2_X1 U5923 ( .A1(n7905), .A2(n7904), .ZN(n9681) );
  NAND2_X1 U5924 ( .A1(n7902), .A2(n6840), .ZN(n7905) );
  NAND2_X1 U5925 ( .A1(n9498), .A2(n9219), .ZN(n9479) );
  AOI21_X1 U5926 ( .B1(n4649), .B2(n4648), .A(n4544), .ZN(n4645) );
  AND2_X1 U5927 ( .A1(n4649), .A2(n4650), .ZN(n9490) );
  INV_X1 U5928 ( .A(n8049), .ZN(n9690) );
  NAND2_X1 U5929 ( .A1(n4832), .A2(n4835), .ZN(n9507) );
  NAND2_X1 U5930 ( .A1(n4834), .A2(n4833), .ZN(n4832) );
  NAND2_X1 U5931 ( .A1(n9536), .A2(n9209), .ZN(n9527) );
  NAND2_X1 U5932 ( .A1(n4623), .A2(n4622), .ZN(n9698) );
  AOI21_X1 U5933 ( .B1(n4624), .B2(n4626), .A(n9538), .ZN(n4622) );
  NAND2_X1 U5934 ( .A1(n4621), .A2(n4624), .ZN(n9546) );
  OR2_X1 U5935 ( .A1(n9598), .A2(n4626), .ZN(n4621) );
  NAND2_X1 U5936 ( .A1(n7823), .A2(n7822), .ZN(n9701) );
  NAND2_X1 U5937 ( .A1(n4979), .A2(n4980), .ZN(n9551) );
  NAND2_X1 U5938 ( .A1(n9583), .A2(n4983), .ZN(n4979) );
  INV_X1 U5939 ( .A(n9712), .ZN(n9580) );
  AOI21_X1 U5940 ( .B1(n9583), .B2(n9591), .A(n4503), .ZN(n9568) );
  AND2_X1 U5941 ( .A1(n4663), .A2(n4661), .ZN(n9640) );
  NAND2_X1 U5942 ( .A1(n4663), .A2(n8031), .ZN(n9638) );
  NAND2_X1 U5943 ( .A1(n4970), .A2(n4974), .ZN(n7408) );
  NAND2_X1 U5944 ( .A1(n7302), .A2(n7301), .ZN(n7303) );
  NAND2_X1 U5945 ( .A1(n6855), .A2(n4998), .ZN(n7137) );
  NOR2_X1 U5946 ( .A1(n6697), .A2(n5097), .ZN(n6698) );
  AND2_X1 U5947 ( .A1(n6463), .A2(n4613), .ZN(n4612) );
  INV_X1 U5948 ( .A(n8981), .ZN(n6631) );
  INV_X1 U5949 ( .A(n9648), .ZN(n10364) );
  OR2_X1 U5950 ( .A1(n6715), .A2(n6305), .ZN(n6308) );
  NAND2_X1 U5951 ( .A1(n6371), .A2(n9555), .ZN(n10366) );
  INV_X1 U5952 ( .A(n9555), .ZN(n10360) );
  INV_X1 U5953 ( .A(n9651), .ZN(n10343) );
  OAI21_X1 U5954 ( .B1(n9657), .B2(n10388), .A(n9656), .ZN(n9744) );
  AOI211_X1 U5955 ( .C1(n10372), .C2(n10267), .A(n10266), .B(n10265), .ZN(
        n10288) );
  INV_X1 U5956 ( .A(n4696), .ZN(n6130) );
  XNOR2_X1 U5957 ( .A(n8188), .B(n8187), .ZN(n9769) );
  OAI21_X1 U5958 ( .B1(n8184), .B2(n8183), .A(n8182), .ZN(n8188) );
  CLKBUF_X1 U5959 ( .A(n5893), .Z(n8071) );
  INV_X1 U5960 ( .A(n5784), .ZN(n7509) );
  NAND2_X1 U5961 ( .A1(n5096), .A2(n4990), .ZN(n4988) );
  XNOR2_X1 U5962 ( .A(n5756), .B(n5755), .ZN(n7858) );
  CLKBUF_X1 U5963 ( .A(n6119), .Z(n9327) );
  AND2_X1 U5964 ( .A1(n6363), .A2(n6441), .ZN(n9383) );
  INV_X1 U5965 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n9876) );
  INV_X1 U5966 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n9902) );
  OR2_X1 U5967 ( .A1(n5796), .A2(n5115), .ZN(n6586) );
  XNOR2_X1 U5968 ( .A(n5294), .B(n5293), .ZN(n6461) );
  NAND2_X1 U5969 ( .A1(n4725), .A2(n5192), .ZN(n5217) );
  NAND2_X1 U5970 ( .A1(n5099), .A2(n5098), .ZN(n5780) );
  XNOR2_X1 U5971 ( .A(n4771), .B(n10113), .ZN(n6309) );
  NAND2_X1 U5972 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n4771) );
  NOR2_X1 U5973 ( .A1(n9800), .A2(n10536), .ZN(n10535) );
  NAND2_X1 U5974 ( .A1(n4601), .A2(n4603), .ZN(n4600) );
  NAND2_X1 U5975 ( .A1(n5001), .A2(n5005), .ZN(n5000) );
  NAND2_X1 U5976 ( .A1(n5049), .A2(n4545), .ZN(n5048) );
  NAND2_X1 U5977 ( .A1(n4945), .A2(n4944), .ZN(n9341) );
  OAI211_X1 U5978 ( .C1(n9402), .C2(n4485), .A(n4769), .B(n4766), .ZN(P1_U3260) );
  INV_X1 U5979 ( .A(n4770), .ZN(n4769) );
  NAND2_X1 U5980 ( .A1(n4767), .A2(n4485), .ZN(n4766) );
  NAND2_X1 U5981 ( .A1(n4652), .A2(n4557), .ZN(P1_U3520) );
  NAND2_X1 U5982 ( .A1(n9745), .A2(n10396), .ZN(n4652) );
  INV_X1 U5983 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n4651) );
  NAND2_X1 U5984 ( .A1(n9506), .A2(n8038), .ZN(n4649) );
  AND2_X1 U5985 ( .A1(n4835), .A2(n4831), .ZN(n4487) );
  AND2_X2 U5986 ( .A1(n9263), .A2(n4485), .ZN(n9256) );
  AND2_X1 U5987 ( .A1(n7181), .A2(n4619), .ZN(n4488) );
  NAND2_X1 U5988 ( .A1(n9117), .A2(n5088), .ZN(n9655) );
  NOR2_X1 U5989 ( .A1(n9418), .A2(n9421), .ZN(n4489) );
  AND2_X1 U5990 ( .A1(n7539), .A2(n4918), .ZN(n4490) );
  INV_X1 U5991 ( .A(n4645), .ZN(n9477) );
  AND2_X1 U5992 ( .A1(n4712), .A2(n10269), .ZN(n4491) );
  INV_X1 U5993 ( .A(n6842), .ZN(n4614) );
  NAND2_X1 U5994 ( .A1(n4523), .A2(n4782), .ZN(n8898) );
  INV_X1 U5995 ( .A(n9147), .ZN(n4844) );
  NAND2_X1 U5996 ( .A1(n7285), .A2(n7284), .ZN(n7407) );
  NAND2_X1 U5997 ( .A1(n5653), .A2(n5652), .ZN(n8783) );
  INV_X1 U5998 ( .A(n8833), .ZN(n8628) );
  NAND2_X1 U5999 ( .A1(n5759), .A2(n5758), .ZN(n8833) );
  AND2_X1 U6000 ( .A1(n8013), .A2(n8012), .ZN(n8077) );
  AND2_X1 U6001 ( .A1(n4679), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n4492) );
  INV_X1 U6002 ( .A(n4837), .ZN(n4833) );
  OR2_X1 U6003 ( .A1(n9271), .A2(n4838), .ZN(n4837) );
  OR2_X1 U6004 ( .A1(n9660), .A2(n4548), .ZN(n4493) );
  INV_X1 U6005 ( .A(n8582), .ZN(n8233) );
  AND2_X1 U6006 ( .A1(n8369), .A2(n8368), .ZN(n8582) );
  AND2_X1 U6007 ( .A1(n5085), .A2(n5083), .ZN(n4494) );
  INV_X1 U6008 ( .A(n5063), .ZN(n10426) );
  NAND2_X1 U6009 ( .A1(n8294), .A2(n8292), .ZN(n5063) );
  INV_X1 U6010 ( .A(n8823), .ZN(n4879) );
  NAND2_X1 U6011 ( .A1(n7071), .A2(n5022), .ZN(n7172) );
  NAND2_X1 U6012 ( .A1(n7639), .A2(n7638), .ZN(n8828) );
  INV_X1 U6013 ( .A(n8828), .ZN(n4904) );
  NAND2_X1 U6014 ( .A1(n5710), .A2(n5709), .ZN(n8662) );
  INV_X1 U6015 ( .A(n7856), .ZN(n4790) );
  INV_X1 U6016 ( .A(n8297), .ZN(n5065) );
  AND2_X1 U6017 ( .A1(n6459), .A2(n6458), .ZN(n4495) );
  AND2_X1 U6018 ( .A1(n7416), .A2(n9094), .ZN(n9287) );
  INV_X1 U6019 ( .A(n6945), .ZN(n6316) );
  OR2_X1 U6020 ( .A1(n8395), .A2(n5213), .ZN(n5214) );
  INV_X2 U6021 ( .A(n6715), .ZN(n6840) );
  NAND2_X2 U6022 ( .A1(n6300), .A2(n8185), .ZN(n6409) );
  OR2_X1 U6023 ( .A1(n8713), .A2(n8126), .ZN(n4497) );
  OR2_X1 U6024 ( .A1(n5205), .A2(P2_IR_REG_29__SCAN_IN), .ZN(n4498) );
  AND2_X1 U6025 ( .A1(n7704), .A2(n7703), .ZN(n4499) );
  NAND2_X2 U6026 ( .A1(n6329), .A2(n6380), .ZN(n6589) );
  OR2_X1 U6027 ( .A1(n6091), .A2(n4772), .ZN(n4500) );
  AND2_X1 U6028 ( .A1(n9125), .A2(n9308), .ZN(n4501) );
  AND2_X1 U6029 ( .A1(n9715), .A2(n9607), .ZN(n4503) );
  INV_X1 U6030 ( .A(n10212), .ZN(n10200) );
  NOR2_X1 U6031 ( .A1(n8678), .A2(n8132), .ZN(n4504) );
  OR2_X1 U6032 ( .A1(n7157), .A2(n10428), .ZN(n8295) );
  AND2_X1 U6033 ( .A1(n4719), .A2(n4716), .ZN(n4505) );
  AND2_X1 U6034 ( .A1(n9112), .A2(n4920), .ZN(n4506) );
  AND2_X1 U6035 ( .A1(n8427), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n4507) );
  AND2_X1 U6036 ( .A1(n5098), .A2(n9983), .ZN(n4508) );
  INV_X1 U6037 ( .A(n9256), .ZN(n9251) );
  NAND2_X1 U6038 ( .A1(n7712), .A2(n8886), .ZN(n4509) );
  AND2_X1 U6039 ( .A1(n8534), .A2(n8389), .ZN(n4510) );
  AND2_X1 U6040 ( .A1(n5016), .A2(n8082), .ZN(n4511) );
  AND2_X1 U6041 ( .A1(n7438), .A2(n7714), .ZN(n4512) );
  NAND2_X1 U6042 ( .A1(n7375), .A2(n7374), .ZN(n9174) );
  INV_X1 U6043 ( .A(n9655), .ZN(n9409) );
  OR2_X1 U6044 ( .A1(n8738), .A2(n4573), .ZN(n4513) );
  AND2_X1 U6045 ( .A1(n9037), .A2(n7721), .ZN(n4514) );
  AND2_X1 U6046 ( .A1(n7474), .A2(n8302), .ZN(n4515) );
  OR2_X1 U6047 ( .A1(n4986), .A2(n4988), .ZN(n4516) );
  AND3_X1 U6048 ( .A1(n5121), .A2(n6117), .A3(n9967), .ZN(n4517) );
  OR2_X1 U6049 ( .A1(n5792), .A2(n5793), .ZN(n6464) );
  XNOR2_X1 U6050 ( .A(n8818), .B(n8225), .ZN(n8569) );
  NAND2_X1 U6051 ( .A1(n8173), .A2(n8172), .ZN(n8529) );
  INV_X1 U6052 ( .A(n8529), .ZN(n4583) );
  NAND2_X1 U6053 ( .A1(n5551), .A2(n5550), .ZN(n8799) );
  XNOR2_X1 U6054 ( .A(n4482), .B(n6042), .ZN(n5252) );
  NAND2_X1 U6055 ( .A1(n7641), .A2(n7640), .ZN(n8823) );
  NAND2_X1 U6056 ( .A1(n7186), .A2(n7185), .ZN(n7300) );
  NAND2_X1 U6057 ( .A1(n4789), .A2(n4790), .ZN(n8998) );
  NAND2_X1 U6058 ( .A1(n9512), .A2(n4706), .ZN(n4709) );
  INV_X1 U6059 ( .A(n8410), .ZN(n8638) );
  AND2_X1 U6060 ( .A1(n8039), .A2(n9345), .ZN(n4518) );
  AND2_X1 U6061 ( .A1(n8197), .A2(n8179), .ZN(n4519) );
  NAND2_X1 U6062 ( .A1(n9707), .A2(n9539), .ZN(n4520) );
  INV_X1 U6063 ( .A(n7710), .ZN(n4812) );
  INV_X1 U6064 ( .A(n9671), .ZN(n9416) );
  NAND2_X1 U6065 ( .A1(n7949), .A2(n7948), .ZN(n9671) );
  AND2_X1 U6066 ( .A1(n8039), .A2(n9511), .ZN(n9065) );
  AND2_X1 U6067 ( .A1(n9690), .A2(n8968), .ZN(n4521) );
  AND2_X1 U6068 ( .A1(n7879), .A2(n7878), .ZN(n9497) );
  INV_X1 U6069 ( .A(n9497), .ZN(n8039) );
  NOR2_X1 U6070 ( .A1(n6401), .A2(n5948), .ZN(n4522) );
  INV_X1 U6071 ( .A(n5032), .ZN(n5031) );
  OR2_X1 U6072 ( .A1(n7064), .A2(n5033), .ZN(n5032) );
  INV_X1 U6073 ( .A(n5007), .ZN(n5006) );
  NAND2_X1 U6074 ( .A1(n5010), .A2(n5008), .ZN(n5007) );
  NAND2_X1 U6075 ( .A1(n4819), .A2(n4817), .ZN(n5126) );
  AND2_X1 U6076 ( .A1(n8998), .A2(n7873), .ZN(n4523) );
  INV_X1 U6077 ( .A(n7635), .ZN(n4891) );
  AND2_X1 U6078 ( .A1(n8775), .A2(n8702), .ZN(n7635) );
  AND2_X1 U6079 ( .A1(n4869), .A2(n4867), .ZN(n4524) );
  OR2_X1 U6080 ( .A1(n5827), .A2(n5118), .ZN(n4525) );
  AND2_X1 U6081 ( .A1(n5312), .A2(SI_6_), .ZN(n4526) );
  NOR2_X1 U6082 ( .A1(n9457), .A2(n9430), .ZN(n4527) );
  INV_X1 U6083 ( .A(n4913), .ZN(n4912) );
  NOR2_X1 U6084 ( .A1(n10233), .A2(n7400), .ZN(n4913) );
  AND2_X1 U6085 ( .A1(n7551), .A2(n8143), .ZN(n4528) );
  INV_X1 U6086 ( .A(n4875), .ZN(n4874) );
  NAND2_X1 U6087 ( .A1(n4877), .A2(n4876), .ZN(n4875) );
  OR2_X1 U6088 ( .A1(n8409), .A2(n8823), .ZN(n4529) );
  AND2_X1 U6089 ( .A1(n4605), .A2(n4607), .ZN(n4530) );
  NAND2_X1 U6090 ( .A1(n5404), .A2(n5403), .ZN(n4531) );
  INV_X1 U6091 ( .A(n4659), .ZN(n4658) );
  OAI21_X1 U6092 ( .B1(n9637), .B2(n4660), .A(n4554), .ZN(n4659) );
  INV_X1 U6093 ( .A(n4880), .ZN(n8605) );
  AND2_X1 U6094 ( .A1(n4733), .A2(n4510), .ZN(n4532) );
  INV_X1 U6095 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n8865) );
  AND2_X1 U6096 ( .A1(n4980), .A2(n4520), .ZN(n4533) );
  AND2_X1 U6097 ( .A1(n5001), .A2(n5007), .ZN(n4534) );
  AND2_X1 U6098 ( .A1(n9423), .A2(n9237), .ZN(n9419) );
  AND2_X1 U6099 ( .A1(n4983), .A2(n4985), .ZN(n4535) );
  NOR2_X1 U6100 ( .A1(n9098), .A2(n9291), .ZN(n4536) );
  AND2_X1 U6101 ( .A1(n4665), .A2(n4661), .ZN(n4537) );
  AND2_X1 U6102 ( .A1(n5019), .A2(n4594), .ZN(n4538) );
  AND2_X1 U6103 ( .A1(n6869), .A2(n6867), .ZN(n4539) );
  INV_X1 U6104 ( .A(n4910), .ZN(n4909) );
  NOR2_X1 U6105 ( .A1(n7463), .A2(n4913), .ZN(n4910) );
  INV_X1 U6106 ( .A(n5090), .ZN(n4641) );
  AND2_X1 U6107 ( .A1(n5125), .A2(n5124), .ZN(n4540) );
  AND2_X1 U6108 ( .A1(n8286), .A2(n8284), .ZN(n4541) );
  NOR2_X1 U6109 ( .A1(n5118), .A2(P1_IR_REG_19__SCAN_IN), .ZN(n4542) );
  INV_X1 U6110 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5154) );
  INV_X1 U6111 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5799) );
  NAND2_X1 U6112 ( .A1(n5052), .A2(n6746), .ZN(n4543) );
  NAND2_X2 U6113 ( .A1(n9771), .A2(n6137), .ZN(n4828) );
  INV_X2 U6114 ( .A(n5520), .ZN(n7670) );
  AND2_X1 U6115 ( .A1(n9497), .A2(n9511), .ZN(n4544) );
  NAND2_X1 U6116 ( .A1(n5637), .A2(n5636), .ZN(n8788) );
  INV_X1 U6117 ( .A(n8788), .ZN(n4876) );
  AND2_X1 U6118 ( .A1(n7980), .A2(n8977), .ZN(n4545) );
  NOR3_X1 U6119 ( .A1(n8075), .A2(n8074), .A3(n8142), .ZN(n4546) );
  INV_X1 U6120 ( .A(n5246), .ZN(n5520) );
  AND2_X1 U6121 ( .A1(n7002), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4547) );
  NAND2_X1 U6122 ( .A1(n8145), .A2(n5642), .ZN(n8083) );
  OAI21_X1 U6123 ( .B1(n7705), .B2(n4810), .A(n4808), .ZN(n9035) );
  AND2_X1 U6124 ( .A1(n8230), .A2(n8231), .ZN(n8601) );
  INV_X1 U6125 ( .A(n8601), .ZN(n4901) );
  INV_X1 U6126 ( .A(n8907), .ZN(n4797) );
  INV_X1 U6127 ( .A(n9150), .ZN(n4847) );
  NAND2_X1 U6128 ( .A1(n7327), .A2(n5057), .ZN(n7371) );
  NAND2_X1 U6129 ( .A1(n7724), .A2(n7723), .ZN(n8934) );
  AND2_X1 U6130 ( .A1(n9661), .A2(n10372), .ZN(n4548) );
  NAND2_X1 U6131 ( .A1(n5147), .A2(n5137), .ZN(n5560) );
  NAND2_X1 U6132 ( .A1(n5638), .A2(n8139), .ZN(n8145) );
  NAND2_X1 U6133 ( .A1(n5025), .A2(n5554), .ZN(n5591) );
  OR2_X1 U6134 ( .A1(n7183), .A2(n10351), .ZN(n9144) );
  INV_X1 U6135 ( .A(n9144), .ZN(n4840) );
  INV_X1 U6136 ( .A(n4631), .ZN(n4630) );
  INV_X1 U6137 ( .A(n8669), .ZN(n8639) );
  AND2_X1 U6138 ( .A1(n7136), .A2(n9351), .ZN(n4549) );
  NAND2_X1 U6139 ( .A1(n7487), .A2(n4874), .ZN(n4878) );
  OR2_X1 U6140 ( .A1(n9525), .A2(n9510), .ZN(n4550) );
  INV_X1 U6141 ( .A(n4699), .ZN(n9552) );
  NOR2_X1 U6142 ( .A1(n9599), .A2(n4700), .ZN(n4699) );
  AND2_X1 U6143 ( .A1(n7407), .A2(n10253), .ZN(n4551) );
  AND2_X1 U6144 ( .A1(n4656), .A2(n4658), .ZN(n4552) );
  INV_X1 U6145 ( .A(n8021), .ZN(n5011) );
  NOR2_X1 U6146 ( .A1(n7183), .A2(n9349), .ZN(n4553) );
  NAND2_X1 U6147 ( .A1(n9731), .A2(n9346), .ZN(n4554) );
  AND2_X1 U6148 ( .A1(n7873), .A2(n4788), .ZN(n4555) );
  AND2_X1 U6149 ( .A1(n10329), .A2(n4759), .ZN(n4556) );
  INV_X1 U6150 ( .A(n4606), .ZN(n4605) );
  OAI21_X1 U6151 ( .B1(n8005), .B2(n4607), .A(n8077), .ZN(n4606) );
  INV_X1 U6152 ( .A(n8037), .ZN(n4650) );
  NAND2_X1 U6154 ( .A1(n7768), .A2(n7767), .ZN(n9715) );
  INV_X1 U6155 ( .A(n9715), .ZN(n4703) );
  OR2_X1 U6156 ( .A1(n10396), .A2(n4651), .ZN(n4557) );
  AND2_X1 U6157 ( .A1(n7217), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n4558) );
  AND2_X1 U6158 ( .A1(n4845), .A2(n4844), .ZN(n4559) );
  NAND2_X1 U6159 ( .A1(n5094), .A2(n5147), .ZN(n5153) );
  AND2_X1 U6160 ( .A1(n4758), .A2(n4759), .ZN(n4560) );
  INV_X1 U6161 ( .A(n4993), .ZN(n6697) );
  AND2_X1 U6162 ( .A1(n6855), .A2(n6854), .ZN(n4561) );
  NAND2_X1 U6163 ( .A1(n5993), .A2(n5994), .ZN(n4562) );
  NAND2_X1 U6164 ( .A1(n4615), .A2(n4617), .ZN(n7188) );
  INV_X1 U6165 ( .A(n8029), .ZN(n4666) );
  AND2_X1 U6166 ( .A1(n7589), .A2(n7588), .ZN(n4563) );
  INV_X1 U6167 ( .A(n9431), .ZN(n4921) );
  AND2_X1 U6168 ( .A1(n7071), .A2(n5453), .ZN(n4564) );
  NAND2_X1 U6169 ( .A1(n7413), .A2(n7412), .ZN(n9739) );
  INV_X1 U6170 ( .A(n9739), .ZN(n4711) );
  INV_X1 U6171 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n4990) );
  INV_X1 U6172 ( .A(n7157), .ZN(n4871) );
  NAND2_X1 U6173 ( .A1(n6594), .A2(n6593), .ZN(n4565) );
  INV_X1 U6174 ( .A(n5040), .ZN(n6228) );
  INV_X1 U6175 ( .A(n8398), .ZN(n5213) );
  OR2_X1 U6176 ( .A1(n8512), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n4566) );
  AND2_X1 U6177 ( .A1(n4670), .A2(n4675), .ZN(n4567) );
  AND2_X1 U6178 ( .A1(n8499), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n4568) );
  INV_X1 U6179 ( .A(n5268), .ZN(n8196) );
  INV_X1 U6180 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n4579) );
  INV_X1 U6181 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n4572) );
  MUX2_X1 U6182 ( .A(n9216), .B(n9215), .S(n9256), .Z(n9218) );
  MUX2_X2 U6183 ( .A(n9206), .B(n9205), .S(n9256), .Z(n9210) );
  NAND2_X1 U6184 ( .A1(n6426), .A2(n9072), .ZN(n9127) );
  INV_X1 U6185 ( .A(n4828), .ZN(n4827) );
  OAI21_X1 U6186 ( .B1(n9262), .B2(n9261), .A(n9260), .ZN(n9266) );
  NAND2_X1 U6187 ( .A1(n4951), .A2(n4946), .ZN(n4945) );
  AOI21_X1 U6188 ( .B1(n4950), .B2(n4949), .A(n9326), .ZN(n4948) );
  NAND2_X2 U6189 ( .A1(n8401), .A2(n5602), .ZN(n5843) );
  NAND2_X2 U6190 ( .A1(n5202), .A2(n5203), .ZN(n8401) );
  NAND2_X1 U6191 ( .A1(n8697), .A2(n7633), .ZN(n7634) );
  NAND2_X1 U6192 ( .A1(n6815), .A2(n6814), .ZN(n6817) );
  OAI21_X1 U6193 ( .B1(n8622), .B2(n4895), .A(n4893), .ZN(n4892) );
  OAI22_X1 U6194 ( .A1(n8567), .A2(n7659), .B1(n8818), .B2(n8584), .ZN(n8536)
         );
  OAI21_X1 U6195 ( .B1(n8804), .B2(n8415), .A(n7481), .ZN(n7482) );
  NAND2_X1 U6196 ( .A1(n7124), .A2(n6044), .ZN(n6045) );
  NAND2_X1 U6197 ( .A1(n6786), .A2(n6282), .ZN(n6283) );
  XNOR2_X1 U6198 ( .A(n8537), .B(n8544), .ZN(n8741) );
  OAI21_X2 U6199 ( .B1(n8645), .B2(n8411), .A(n8761), .ZN(n8622) );
  NAND2_X1 U6200 ( .A1(n7159), .A2(n7158), .ZN(n7240) );
  NAND2_X1 U6201 ( .A1(n7514), .A2(n7516), .ZN(n5025) );
  NAND2_X1 U6202 ( .A1(n5015), .A2(n5013), .ZN(n8124) );
  NAND2_X1 U6203 ( .A1(n7372), .A2(n8189), .ZN(n5462) );
  NOR2_X1 U6204 ( .A1(n5019), .A2(n4594), .ZN(n4592) );
  OAI21_X1 U6205 ( .B1(n8193), .B2(n8198), .A(n8387), .ZN(n8194) );
  INV_X1 U6206 ( .A(n8546), .ZN(n4575) );
  OAI21_X1 U6207 ( .B1(n4735), .B2(n8408), .A(n8379), .ZN(n4734) );
  INV_X1 U6208 ( .A(n5199), .ZN(n4943) );
  AOI21_X1 U6209 ( .B1(n4733), .B2(n8408), .A(n8382), .ZN(n4732) );
  NAND2_X1 U6210 ( .A1(n5477), .A2(n5476), .ZN(n4966) );
  INV_X1 U6211 ( .A(n4942), .ZN(n4941) );
  NAND2_X1 U6212 ( .A1(n8397), .A2(n8399), .ZN(n4722) );
  NAND2_X1 U6213 ( .A1(n4722), .A2(n5213), .ZN(n4721) );
  NAND2_X1 U6214 ( .A1(n6484), .A2(n8202), .ZN(n6818) );
  INV_X1 U6215 ( .A(n5061), .ZN(n5060) );
  NAND4_X2 U6216 ( .A1(n5081), .A2(n5094), .A3(n5136), .A4(n5135), .ZN(n5149)
         );
  NAND2_X1 U6217 ( .A1(n6967), .A2(n8290), .ZN(n10425) );
  NAND2_X1 U6218 ( .A1(n8698), .A2(n8699), .ZN(n8682) );
  AOI21_X2 U6219 ( .B1(n8596), .B2(n8601), .A(n7665), .ZN(n8583) );
  NAND2_X1 U6220 ( .A1(n4739), .A2(n4743), .ZN(n5405) );
  OAI21_X1 U6221 ( .B1(n8176), .B2(n8535), .A(n8227), .ZN(n8545) );
  OAI21_X1 U6222 ( .B1(n8650), .B2(n8655), .A(n8342), .ZN(n8635) );
  OAI211_X1 U6223 ( .C1(n5274), .C2(n4726), .A(n4723), .B(n5216), .ZN(n5196)
         );
  OR2_X1 U6225 ( .A1(n8522), .A2(n10472), .ZN(n8730) );
  MUX2_X1 U6226 ( .A(n10413), .B(n8873), .S(n5843), .Z(n7120) );
  NAND2_X1 U6227 ( .A1(n5243), .A2(n4580), .ZN(n5181) );
  NAND2_X1 U6228 ( .A1(n6818), .A2(n5068), .ZN(n5067) );
  NAND2_X1 U6229 ( .A1(n7485), .A2(n8319), .ZN(n7542) );
  NAND2_X1 U6230 ( .A1(n5075), .A2(n5074), .ZN(n8571) );
  NAND2_X1 U6231 ( .A1(n5275), .A2(n5274), .ZN(n4725) );
  NAND2_X1 U6232 ( .A1(n5238), .A2(n4713), .ZN(n5183) );
  AND3_X2 U6233 ( .A1(n7702), .A2(n8063), .A3(n10465), .ZN(n6790) );
  NAND2_X1 U6234 ( .A1(n6793), .A2(n5072), .ZN(n5071) );
  NAND2_X1 U6235 ( .A1(n8424), .A2(n7088), .ZN(n8274) );
  NAND2_X1 U6236 ( .A1(n8267), .A2(n8274), .ZN(n8199) );
  NOR2_X2 U6237 ( .A1(n8538), .A2(n8739), .ZN(n4584) );
  XNOR2_X1 U6238 ( .A(n4585), .B(n8102), .ZN(n8108) );
  OR2_X2 U6239 ( .A1(n6183), .A2(n6184), .ZN(n4587) );
  AOI21_X2 U6240 ( .B1(n5029), .B2(n8110), .A(n5027), .ZN(n5026) );
  OAI21_X2 U6241 ( .B1(n6667), .B2(n5357), .A(n6666), .ZN(n8110) );
  NOR2_X2 U6242 ( .A1(n5613), .A2(n5612), .ZN(n6667) );
  NAND2_X1 U6243 ( .A1(n7068), .A2(n4595), .ZN(n4597) );
  AND2_X1 U6244 ( .A1(n7068), .A2(n4589), .ZN(n4593) );
  NAND2_X1 U6245 ( .A1(n4591), .A2(n4590), .ZN(n10189) );
  NAND2_X1 U6246 ( .A1(n4597), .A2(n4538), .ZN(n4590) );
  NOR2_X1 U6247 ( .A1(n4593), .A2(n4592), .ZN(n4591) );
  OAI21_X2 U6248 ( .B1(n10189), .B2(n10190), .A(n5528), .ZN(n7514) );
  NAND2_X1 U6249 ( .A1(n4597), .A2(n5019), .ZN(n5527) );
  INV_X1 U6250 ( .A(n5526), .ZN(n4594) );
  NAND2_X1 U6251 ( .A1(n8006), .A2(n4599), .ZN(n4598) );
  OAI211_X1 U6252 ( .C1(n8006), .C2(n4600), .A(n4598), .B(n8080), .ZN(P2_U3216) );
  NAND2_X1 U6253 ( .A1(n8006), .A2(n8005), .ZN(n8158) );
  AND2_X1 U6254 ( .A1(n5137), .A2(n4610), .ZN(n4609) );
  INV_X1 U6255 ( .A(n10338), .ZN(n4616) );
  OAI21_X1 U6256 ( .B1(n10338), .B2(n7138), .A(n4620), .ZN(n7182) );
  NAND2_X1 U6257 ( .A1(n9598), .A2(n4624), .ZN(n4623) );
  NOR2_X1 U6258 ( .A1(n9603), .A2(n9622), .ZN(n4631) );
  INV_X1 U6259 ( .A(n9461), .ZN(n4640) );
  NAND2_X1 U6260 ( .A1(n9506), .A2(n4643), .ZN(n4642) );
  NAND2_X1 U6261 ( .A1(n4642), .A2(n4646), .ZN(n8041) );
  NAND2_X1 U6262 ( .A1(n8030), .A2(n4537), .ZN(n4655) );
  NAND2_X1 U6263 ( .A1(n4655), .A2(n4657), .ZN(n9612) );
  OAI21_X1 U6264 ( .B1(P2_IR_REG_1__SCAN_IN), .B2(n10413), .A(n4668), .ZN(
        n4678) );
  OAI21_X1 U6265 ( .B1(n4678), .B2(P2_REG1_REG_1__SCAN_IN), .A(n4676), .ZN(
        n4671) );
  OAI21_X1 U6266 ( .B1(n4675), .B2(n6002), .A(n4672), .ZN(n6001) );
  INV_X1 U6267 ( .A(n4673), .ZN(n4672) );
  OAI22_X1 U6268 ( .A1(n4678), .A2(n4674), .B1(n6002), .B2(n4676), .ZN(n4673)
         );
  INV_X1 U6269 ( .A(n5118), .ZN(n4694) );
  INV_X1 U6270 ( .A(n4698), .ZN(n9534) );
  NAND2_X1 U6271 ( .A1(n9512), .A2(n4704), .ZN(n9454) );
  INV_X1 U6272 ( .A(n4709), .ZN(n9462) );
  XNOR2_X1 U6273 ( .A(n5238), .B(n4713), .ZN(n6305) );
  NAND2_X1 U6274 ( .A1(n5189), .A2(n4724), .ZN(n4723) );
  INV_X1 U6275 ( .A(n5192), .ZN(n4726) );
  NAND2_X1 U6276 ( .A1(n5189), .A2(n5188), .ZN(n5275) );
  NAND2_X1 U6277 ( .A1(n8375), .A2(n4735), .ZN(n8380) );
  NAND2_X1 U6278 ( .A1(n4729), .A2(n4727), .ZN(n8386) );
  OR2_X1 U6279 ( .A1(n8375), .A2(n8408), .ZN(n4728) );
  NAND2_X1 U6280 ( .A1(n8381), .A2(n4730), .ZN(n4729) );
  NAND2_X1 U6281 ( .A1(n4731), .A2(n4732), .ZN(n4730) );
  NAND2_X1 U6282 ( .A1(n8375), .A2(n4733), .ZN(n4731) );
  NAND2_X1 U6283 ( .A1(n5359), .A2(n5360), .ZN(n4739) );
  NAND2_X1 U6284 ( .A1(n4745), .A2(n8317), .ZN(n8322) );
  NAND2_X1 U6285 ( .A1(n4746), .A2(n8315), .ZN(n4745) );
  NAND3_X1 U6286 ( .A1(n4749), .A2(n4747), .A3(n7463), .ZN(n4746) );
  NAND2_X1 U6287 ( .A1(n4748), .A2(n8389), .ZN(n4747) );
  NAND2_X1 U6288 ( .A1(n8305), .A2(n8304), .ZN(n4748) );
  NAND2_X1 U6289 ( .A1(n4750), .A2(n8382), .ZN(n4749) );
  NAND2_X1 U6290 ( .A1(n8312), .A2(n8311), .ZN(n4750) );
  AOI21_X1 U6291 ( .B1(n4751), .B2(n8359), .A(n8358), .ZN(n8365) );
  NAND3_X1 U6292 ( .A1(n4753), .A2(n8355), .A3(n4752), .ZN(n4751) );
  NAND3_X1 U6293 ( .A1(n8353), .A2(n8354), .A3(n8389), .ZN(n4752) );
  OAI21_X1 U6294 ( .B1(n4757), .B2(n6104), .A(n4755), .ZN(n6191) );
  NAND2_X1 U6295 ( .A1(n4758), .A2(n4556), .ZN(n10328) );
  INV_X1 U6296 ( .A(n4763), .ZN(n9360) );
  MUX2_X1 U6297 ( .A(n5944), .B(P1_REG2_REG_1__SCAN_IN), .S(n6309), .Z(n6064)
         );
  INV_X1 U6298 ( .A(n6689), .ZN(n4777) );
  INV_X1 U6299 ( .A(n6688), .ZN(n4778) );
  NAND2_X1 U6300 ( .A1(n6549), .A2(n6676), .ZN(n4779) );
  NAND2_X1 U6301 ( .A1(n6547), .A2(n6674), .ZN(n4780) );
  CLKBUF_X1 U6302 ( .A(n9001), .Z(n4782) );
  NAND2_X1 U6303 ( .A1(n8997), .A2(n8996), .ZN(n9001) );
  NAND2_X1 U6304 ( .A1(n4791), .A2(n4793), .ZN(n7840) );
  NAND2_X1 U6305 ( .A1(n8910), .A2(n4795), .ZN(n4791) );
  NAND2_X2 U6306 ( .A1(n4816), .A2(n9022), .ZN(n8877) );
  INV_X2 U6307 ( .A(n7891), .ZN(n7961) );
  NAND2_X2 U6308 ( .A1(n6618), .A2(n6380), .ZN(n7891) );
  NAND3_X1 U6309 ( .A1(n4543), .A2(n4822), .A3(n5050), .ZN(n4821) );
  NAND3_X1 U6310 ( .A1(n8975), .A2(n8978), .A3(n5051), .ZN(n4822) );
  NAND2_X1 U6311 ( .A1(n8956), .A2(n7765), .ZN(n7783) );
  NAND2_X1 U6312 ( .A1(n7840), .A2(n7839), .ZN(n7857) );
  NAND2_X1 U6313 ( .A1(n8957), .A2(n8958), .ZN(n8956) );
  NAND2_X1 U6314 ( .A1(n8925), .A2(n8926), .ZN(n8924) );
  INV_X2 U6315 ( .A(n6553), .ZN(n7320) );
  INV_X1 U6316 ( .A(n6745), .ZN(n5050) );
  NAND2_X1 U6317 ( .A1(n4940), .A2(n5199), .ZN(n5311) );
  NAND2_X1 U6318 ( .A1(n6153), .A2(n6538), .ZN(n6540) );
  NAND2_X1 U6319 ( .A1(n9010), .A2(n9013), .ZN(n8910) );
  NOR2_X4 U6320 ( .A1(n10340), .A2(n7183), .ZN(n7202) );
  NAND2_X1 U6321 ( .A1(n10176), .A2(n5177), .ZN(n4969) );
  INV_X1 U6322 ( .A(n6538), .ZN(n6539) );
  INV_X1 U6323 ( .A(n8877), .ZN(n5047) );
  INV_X1 U6324 ( .A(n5045), .ZN(n5044) );
  NAND2_X1 U6325 ( .A1(n8935), .A2(n7746), .ZN(n8957) );
  NAND2_X1 U6326 ( .A1(n7000), .A2(n6999), .ZN(n7267) );
  NAND2_X1 U6327 ( .A1(n8964), .A2(n7901), .ZN(n8925) );
  NAND2_X2 U6328 ( .A1(n4823), .A2(n6424), .ZN(n9306) );
  OAI21_X1 U6329 ( .B1(n6323), .B2(n9278), .A(n4823), .ZN(n6332) );
  AND2_X2 U6330 ( .A1(n6137), .A2(n6138), .ZN(n7984) );
  NAND3_X1 U6331 ( .A1(n6137), .A2(n6138), .A3(P1_REG3_REG_1__SCAN_IN), .ZN(
        n4825) );
  INV_X1 U6332 ( .A(n9537), .ZN(n4834) );
  NAND2_X1 U6333 ( .A1(n4829), .A2(n4830), .ZN(n9499) );
  NAND2_X1 U6334 ( .A1(n9537), .A2(n4487), .ZN(n4829) );
  NAND2_X1 U6335 ( .A1(n6839), .A2(n4842), .ZN(n4841) );
  NAND2_X1 U6336 ( .A1(n6839), .A2(n9137), .ZN(n7139) );
  INV_X1 U6337 ( .A(n4845), .ZN(n10347) );
  NAND2_X1 U6338 ( .A1(n9498), .A2(n4854), .ZN(n4848) );
  NAND2_X1 U6339 ( .A1(n4848), .A2(n4851), .ZN(n9441) );
  OAI21_X2 U6340 ( .B1(n9127), .B2(n9309), .A(n9307), .ZN(n6725) );
  NOR2_X2 U6341 ( .A1(n6873), .A2(n6960), .ZN(n10420) );
  NAND2_X1 U6342 ( .A1(n7487), .A2(n4873), .ZN(n8706) );
  INV_X1 U6343 ( .A(n4878), .ZN(n8705) );
  NAND2_X1 U6344 ( .A1(n7634), .A2(n4882), .ZN(n4881) );
  NAND2_X1 U6345 ( .A1(n4881), .A2(n4884), .ZN(n8654) );
  INV_X1 U6346 ( .A(n4892), .ZN(n8567) );
  NAND2_X1 U6347 ( .A1(n10201), .A2(n4910), .ZN(n4906) );
  NAND2_X1 U6348 ( .A1(n4906), .A2(n4907), .ZN(n7466) );
  NAND2_X1 U6349 ( .A1(n10414), .A2(n4915), .ZN(n7159) );
  NAND2_X1 U6350 ( .A1(n6868), .A2(n4539), .ZN(n6962) );
  NAND2_X1 U6351 ( .A1(n7482), .A2(n4490), .ZN(n4916) );
  NAND2_X1 U6352 ( .A1(n4916), .A2(n4917), .ZN(n7632) );
  INV_X1 U6353 ( .A(n4919), .ZN(n7538) );
  INV_X2 U6354 ( .A(n5149), .ZN(n5151) );
  NAND2_X1 U6355 ( .A1(n5648), .A2(n4926), .ZN(n4922) );
  NAND2_X1 U6356 ( .A1(n4922), .A2(n4923), .ZN(n5704) );
  NAND2_X1 U6357 ( .A1(n5294), .A2(n4941), .ZN(n4939) );
  NAND2_X1 U6358 ( .A1(n5294), .A2(n5293), .ZN(n4940) );
  OAI21_X1 U6359 ( .B1(n5538), .B2(n5537), .A(n5539), .ZN(n5556) );
  OAI21_X1 U6360 ( .B1(n5725), .B2(n5724), .A(n5726), .ZN(n5756) );
  INV_X2 U6361 ( .A(n5180), .ZN(n8185) );
  NAND2_X2 U6362 ( .A1(n4969), .A2(n4967), .ZN(n5180) );
  NAND3_X1 U6363 ( .A1(n4694), .A2(n5113), .A3(n5096), .ZN(n5110) );
  NAND2_X1 U6364 ( .A1(n6459), .A2(n4994), .ZN(n4993) );
  NAND2_X1 U6365 ( .A1(n8158), .A2(n4534), .ZN(n4999) );
  OAI211_X1 U6366 ( .C1(n8158), .C2(n5000), .A(n8028), .B(n4999), .ZN(P2_U3222) );
  INV_X1 U6367 ( .A(n5089), .ZN(n5012) );
  NAND2_X1 U6368 ( .A1(n5638), .A2(n4511), .ZN(n5015) );
  NAND2_X1 U6369 ( .A1(n5173), .A2(n5018), .ZN(n5168) );
  NAND2_X1 U6370 ( .A1(n5025), .A2(n5023), .ZN(n5628) );
  NAND2_X1 U6371 ( .A1(n8109), .A2(n5380), .ZN(n7063) );
  INV_X2 U6372 ( .A(n8155), .ZN(n8006) );
  NAND2_X1 U6373 ( .A1(n6540), .A2(n6541), .ZN(n6675) );
  NAND4_X1 U6374 ( .A1(n5048), .A2(n5043), .A3(n5041), .A4(n7995), .ZN(
        P1_U3218) );
  NAND3_X1 U6375 ( .A1(n5045), .A2(n5042), .A3(n7982), .ZN(n5041) );
  AND2_X1 U6376 ( .A1(n6746), .A2(n8974), .ZN(n5051) );
  INV_X1 U6377 ( .A(n6573), .ZN(n5052) );
  NAND2_X1 U6378 ( .A1(n5053), .A2(n8975), .ZN(n8976) );
  NAND2_X1 U6379 ( .A1(n7724), .A2(n5054), .ZN(n8935) );
  INV_X2 U6380 ( .A(n7891), .ZN(n7750) );
  NAND3_X1 U6381 ( .A1(n6946), .A2(n6931), .A3(n6950), .ZN(n7000) );
  NAND2_X1 U6382 ( .A1(n5117), .A2(n5093), .ZN(n5827) );
  NAND2_X1 U6383 ( .A1(n5117), .A2(n5059), .ZN(n6121) );
  NAND3_X1 U6384 ( .A1(n5099), .A2(n4508), .A3(n5114), .ZN(n5795) );
  NAND2_X1 U6385 ( .A1(n7875), .A2(n8899), .ZN(n8967) );
  NAND2_X1 U6386 ( .A1(n5067), .A2(n4541), .ZN(n6967) );
  NAND2_X1 U6387 ( .A1(n5070), .A2(n5071), .ZN(n6499) );
  NOR2_X1 U6388 ( .A1(n8199), .A2(n5073), .ZN(n5072) );
  NAND2_X1 U6389 ( .A1(n8583), .A2(n8582), .ZN(n5075) );
  NAND2_X1 U6390 ( .A1(n5151), .A2(n5085), .ZN(n5205) );
  NAND2_X1 U6391 ( .A1(n5151), .A2(n4494), .ZN(n5082) );
  OR2_X2 U6392 ( .A1(n8635), .A2(n8640), .ZN(n8633) );
  OAI21_X2 U6393 ( .B1(n8667), .B2(n8666), .A(n8344), .ZN(n8650) );
  NAND2_X1 U6394 ( .A1(n4640), .A2(n8042), .ZN(n9445) );
  XNOR2_X1 U6395 ( .A(n8171), .B(n7592), .ZN(n9051) );
  XNOR2_X1 U6396 ( .A(n8043), .B(n9424), .ZN(n9673) );
  NAND2_X1 U6397 ( .A1(n9445), .A2(n9420), .ZN(n8043) );
  NAND2_X1 U6398 ( .A1(n7603), .A2(n6310), .ZN(n6322) );
  OAI21_X1 U6399 ( .B1(n8171), .B2(n8170), .A(n8169), .ZN(n8181) );
  OAI21_X1 U6400 ( .B1(n7590), .B2(n5185), .A(n5184), .ZN(n5187) );
  NAND2_X1 U6401 ( .A1(n7590), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5184) );
  XNOR2_X1 U6402 ( .A(n5128), .B(n6127), .ZN(n5942) );
  NAND2_X1 U6403 ( .A1(n5128), .A2(n5127), .ZN(n6126) );
  NOR2_X1 U6404 ( .A1(n6132), .A2(n6131), .ZN(n6133) );
  XNOR2_X1 U6405 ( .A(n6126), .B(P1_IR_REG_28__SCAN_IN), .ZN(n5893) );
  AND2_X1 U6406 ( .A1(n9451), .A2(n9450), .ZN(n9663) );
  NOR2_X2 U6407 ( .A1(n6789), .A2(n6287), .ZN(n6503) );
  AND2_X1 U6408 ( .A1(n5231), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5232) );
  NAND2_X1 U6409 ( .A1(n7525), .A2(n7524), .ZN(n7527) );
  XNOR2_X1 U6410 ( .A(n7525), .B(n7524), .ZN(n7922) );
  INV_X1 U6411 ( .A(n5807), .ZN(n5117) );
  NAND2_X1 U6412 ( .A1(n5115), .A2(n5799), .ZN(n5807) );
  NAND2_X1 U6413 ( .A1(n5527), .A2(n5526), .ZN(n5528) );
  AND2_X1 U6414 ( .A1(n5230), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5233) );
  CLKBUF_X1 U6415 ( .A(n5802), .Z(n7669) );
  AND2_X1 U6416 ( .A1(n8545), .A2(n8544), .ZN(n8547) );
  OR2_X1 U6417 ( .A1(n6409), .A2(n5910), .ZN(n5088) );
  NOR2_X1 U6418 ( .A1(n8014), .A2(n8077), .ZN(n5089) );
  NOR2_X1 U6419 ( .A1(n9421), .A2(n9444), .ZN(n5090) );
  OR2_X1 U6420 ( .A1(n8034), .A2(n9563), .ZN(n5092) );
  AND2_X1 U6421 ( .A1(n5116), .A2(n5808), .ZN(n5093) );
  AND4_X1 U6422 ( .A1(n5146), .A2(n5145), .A3(n5144), .A4(n5143), .ZN(n5094)
         );
  INV_X1 U6423 ( .A(n6404), .ZN(n7811) );
  INV_X1 U6424 ( .A(n5795), .ZN(n5115) );
  INV_X1 U6425 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n6135) );
  INV_X1 U6426 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5368) );
  AND2_X1 U6427 ( .A1(n5214), .A2(n8399), .ZN(n8637) );
  INV_X1 U6428 ( .A(n8637), .ZN(n10432) );
  NOR2_X1 U6429 ( .A1(n8395), .A2(n8517), .ZN(n5095) );
  AND2_X1 U6430 ( .A1(n7889), .A2(n7888), .ZN(n9511) );
  INV_X1 U6431 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n5185) );
  AND2_X1 U6432 ( .A1(n9354), .A2(n8950), .ZN(n5097) );
  OR2_X1 U6433 ( .A1(n5452), .A2(n5451), .ZN(n5453) );
  OR2_X1 U6434 ( .A1(n6766), .A2(n6208), .ZN(n10494) );
  NAND2_X1 U6435 ( .A1(n9442), .A2(n9256), .ZN(n9244) );
  INV_X1 U6436 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5100) );
  OAI21_X1 U6437 ( .B1(n9302), .B2(n5091), .A(n9244), .ZN(n9249) );
  AND2_X1 U6438 ( .A1(n9424), .A2(n9420), .ZN(n9444) );
  INV_X1 U6439 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5124) );
  INV_X1 U6440 ( .A(n5670), .ZN(n5618) );
  INV_X1 U6441 ( .A(n5711), .ZN(n5619) );
  OAI22_X1 U6442 ( .A1(n7396), .A2(n8208), .B1(n10217), .B2(n7395), .ZN(n10201) );
  INV_X1 U6443 ( .A(n7882), .ZN(n7880) );
  INV_X1 U6444 ( .A(n7730), .ZN(n7728) );
  INV_X1 U6445 ( .A(n7383), .ZN(n7381) );
  INV_X1 U6446 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n6934) );
  INV_X1 U6447 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n6124) );
  INV_X1 U6448 ( .A(n7448), .ZN(n7450) );
  INV_X1 U6449 ( .A(n5643), .ZN(n5644) );
  INV_X1 U6450 ( .A(n5629), .ZN(n5631) );
  OR2_X1 U6451 ( .A1(n5479), .A2(n5478), .ZN(n5480) );
  AND2_X1 U6452 ( .A1(n5425), .A2(n5428), .ZN(n5472) );
  AND2_X1 U6453 ( .A1(n7346), .A2(n5494), .ZN(n5495) );
  NAND2_X1 U6454 ( .A1(n5270), .A2(n5272), .ZN(n5273) );
  OR2_X1 U6455 ( .A1(n5688), .A2(n8093), .ZN(n5711) );
  NAND2_X1 U6456 ( .A1(n5618), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5688) );
  NAND2_X1 U6457 ( .A1(n5298), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5322) );
  OAI22_X1 U6458 ( .A1(n8550), .A2(n10429), .B1(n8549), .B2(n8548), .ZN(n8551)
         );
  OR2_X1 U6459 ( .A1(n5762), .A2(n8104), .ZN(n7642) );
  NAND2_X1 U6460 ( .A1(n5603), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5654) );
  AND2_X1 U6461 ( .A1(n5412), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5442) );
  INV_X1 U6462 ( .A(n8662), .ZN(n8767) );
  INV_X1 U6463 ( .A(n8937), .ZN(n7745) );
  NAND2_X1 U6464 ( .A1(n7880), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n7906) );
  NAND2_X1 U6465 ( .A1(n6146), .A2(n6145), .ZN(n6147) );
  NAND2_X1 U6466 ( .A1(n7015), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n7192) );
  NAND2_X1 U6467 ( .A1(n7926), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n7965) );
  NAND2_X1 U6468 ( .A1(n7862), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n7882) );
  OR2_X1 U6469 ( .A1(n7824), .A2(n8918), .ZN(n7845) );
  NAND2_X1 U6470 ( .A1(n6313), .A2(n6312), .ZN(n6396) );
  XNOR2_X1 U6471 ( .A(n5263), .B(n8063), .ZN(n5271) );
  OR2_X1 U6472 ( .A1(n7642), .A2(n10151), .ZN(n7652) );
  NOR2_X1 U6473 ( .A1(n5487), .A2(n5486), .ZN(n5515) );
  OR2_X1 U6474 ( .A1(n5654), .A2(n8085), .ZN(n5670) );
  INV_X1 U6475 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n10062) );
  NAND2_X1 U6476 ( .A1(n5442), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5463) );
  AND2_X1 U6477 ( .A1(n8402), .A2(n8249), .ZN(n6035) );
  AND2_X1 U6478 ( .A1(n7981), .A2(n8977), .ZN(n7982) );
  OR2_X1 U6479 ( .A1(n7906), .A2(n8928), .ZN(n7927) );
  OR2_X1 U6480 ( .A1(n7752), .A2(n7751), .ZN(n7771) );
  INV_X1 U6481 ( .A(n9349), .ZN(n10351) );
  OR2_X1 U6482 ( .A1(n6846), .A2(n6845), .ZN(n6935) );
  NAND2_X1 U6483 ( .A1(n6557), .A2(n6556), .ZN(n6558) );
  OR2_X1 U6484 ( .A1(n6622), .A2(n6602), .ZN(n6613) );
  OR2_X1 U6485 ( .A1(n9494), .A2(n7929), .ZN(n7889) );
  INV_X1 U6486 ( .A(n9346), .ZN(n9621) );
  AND2_X1 U6487 ( .A1(n10345), .A2(n9148), .ZN(n6856) );
  NAND2_X1 U6488 ( .A1(n6415), .A2(n9275), .ZN(n6459) );
  OR2_X1 U6489 ( .A1(n6328), .A2(n8071), .ZN(n10352) );
  NAND2_X1 U6490 ( .A1(n10393), .A2(n6370), .ZN(n9555) );
  AND2_X1 U6491 ( .A1(n6318), .A2(n6317), .ZN(n9620) );
  AND2_X1 U6492 ( .A1(n5785), .A2(n5784), .ZN(n9761) );
  AND2_X1 U6493 ( .A1(n5757), .A2(n5730), .ZN(n5755) );
  NAND2_X1 U6494 ( .A1(n5634), .A2(n5633), .ZN(n5645) );
  NAND2_X1 U6495 ( .A1(n5539), .A2(n5508), .ZN(n5537) );
  NOR2_X1 U6496 ( .A1(n5827), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n6025) );
  INV_X1 U6497 ( .A(n8618), .ZN(n8586) );
  AND2_X1 U6498 ( .A1(n5626), .A2(n5625), .ZN(n8411) );
  AND4_X1 U6499 ( .A1(n5525), .A2(n5524), .A3(n5523), .A4(n5522), .ZN(n7465)
         );
  NAND2_X1 U6500 ( .A1(n5231), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5287) );
  AND2_X1 U6501 ( .A1(n5862), .A2(n5861), .ZN(n10403) );
  OR2_X1 U6502 ( .A1(n5212), .A2(n8398), .ZN(n10472) );
  NAND2_X1 U6503 ( .A1(n8385), .A2(n8379), .ZN(n8544) );
  AND2_X1 U6504 ( .A1(n6035), .A2(n7571), .ZN(n10216) );
  AND2_X1 U6505 ( .A1(n10499), .A2(n8803), .ZN(n8773) );
  NAND2_X1 U6506 ( .A1(n8342), .A2(n8345), .ZN(n8655) );
  AND2_X1 U6507 ( .A1(n8332), .A2(n8331), .ZN(n8213) );
  AND2_X1 U6508 ( .A1(n10224), .A2(n10223), .ZN(n10237) );
  INV_X1 U6509 ( .A(n10466), .ZN(n10485) );
  AND2_X1 U6510 ( .A1(n7927), .A2(n7907), .ZN(n9484) );
  AND2_X1 U6511 ( .A1(n6614), .A2(n8071), .ZN(n9030) );
  AND2_X1 U6512 ( .A1(n7831), .A2(n7830), .ZN(n9563) );
  AND2_X1 U6513 ( .A1(n5951), .A2(n9335), .ZN(n10331) );
  AND2_X1 U6514 ( .A1(n5951), .A2(n8071), .ZN(n10324) );
  INV_X1 U6515 ( .A(n9419), .ZN(n9424) );
  INV_X1 U6516 ( .A(n10352), .ZN(n10252) );
  INV_X1 U6517 ( .A(n9620), .ZN(n10355) );
  AND2_X1 U6518 ( .A1(n10366), .A2(n6623), .ZN(n9648) );
  OR2_X1 U6519 ( .A1(n6373), .A2(n6316), .ZN(n10388) );
  INV_X1 U6520 ( .A(n10279), .ZN(n9742) );
  AND2_X1 U6521 ( .A1(n9256), .A2(n6945), .ZN(n10393) );
  AND2_X1 U6522 ( .A1(n6058), .A2(n5969), .ZN(n7283) );
  AND2_X1 U6523 ( .A1(n5810), .A2(n5820), .ZN(n10300) );
  XNOR2_X1 U6524 ( .A(n5194), .B(n5193), .ZN(n5216) );
  NOR2_X1 U6525 ( .A1(n6043), .A2(n8196), .ZN(n6102) );
  NAND2_X1 U6526 ( .A1(n5601), .A2(n5590), .ZN(n8156) );
  OR2_X1 U6527 ( .A1(n5832), .A2(n5814), .ZN(n8412) );
  INV_X1 U6528 ( .A(n10499), .ZN(n10504) );
  AND2_X1 U6529 ( .A1(n10237), .A2(n10236), .ZN(n10240) );
  OR2_X1 U6530 ( .A1(n10458), .A2(n10457), .ZN(n10461) );
  XNOR2_X1 U6531 ( .A(n5142), .B(n5141), .ZN(n7367) );
  INV_X1 U6532 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6062) );
  INV_X1 U6533 ( .A(n9693), .ZN(n9525) );
  INV_X1 U6534 ( .A(n8977), .ZN(n9049) );
  NAND2_X1 U6535 ( .A1(n7935), .A2(n7934), .ZN(n9344) );
  OR2_X1 U6536 ( .A1(P1_U3083), .A2(n5892), .ZN(n10337) );
  INV_X1 U6537 ( .A(n10370), .ZN(n10371) );
  INV_X1 U6538 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n9943) );
  INV_X1 U6539 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n10063) );
  NOR2_X1 U6540 ( .A1(n10535), .A2(n10534), .ZN(n10533) );
  NAND2_X1 U6541 ( .A1(n5774), .A2(n5775), .ZN(n5778) );
  NOR2_X1 U6542 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n5103) );
  NAND2_X1 U6543 ( .A1(n5105), .A2(n5124), .ZN(n5107) );
  NAND2_X1 U6544 ( .A1(n5107), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5104) );
  XNOR2_X1 U6545 ( .A(n5104), .B(P1_IR_REG_26__SCAN_IN), .ZN(n5784) );
  OR2_X1 U6546 ( .A1(n5105), .A2(n5124), .ZN(n5106) );
  NAND2_X1 U6547 ( .A1(n5107), .A2(n5106), .ZN(n7461) );
  NAND2_X1 U6548 ( .A1(n4516), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5109) );
  XNOR2_X1 U6549 ( .A(n5109), .B(n5108), .ZN(n7364) );
  NAND2_X1 U6550 ( .A1(n5110), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5111) );
  XNOR2_X1 U6551 ( .A(n5111), .B(n4990), .ZN(n7246) );
  INV_X1 U6552 ( .A(n7246), .ZN(n5112) );
  NOR2_X1 U6553 ( .A1(n6618), .A2(n5112), .ZN(n5892) );
  AND2_X2 U6554 ( .A1(n5892), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U4006) );
  INV_X1 U6555 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n5116) );
  NAND2_X1 U6556 ( .A1(n5122), .A2(n5121), .ZN(n5120) );
  NAND2_X1 U6557 ( .A1(n5120), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5119) );
  NAND2_X1 U6558 ( .A1(n9338), .A2(n5055), .ZN(n6328) );
  NAND2_X1 U6559 ( .A1(n6328), .A2(n6618), .ZN(n5123) );
  NAND2_X1 U6560 ( .A1(n5123), .A2(n7246), .ZN(n5943) );
  NAND2_X1 U6561 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), 
        .ZN(n5127) );
  INV_X1 U6562 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n6127) );
  NAND2_X1 U6563 ( .A1(n5943), .A2(n6842), .ZN(n5129) );
  NAND2_X1 U6564 ( .A1(n5129), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  AND4_X2 U6565 ( .A1(n5340), .A2(n5132), .A3(n5131), .A4(n5130), .ZN(n5136)
         );
  INV_X1 U6566 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5175) );
  INV_X1 U6567 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5166) );
  NAND2_X1 U6568 ( .A1(n5167), .A2(n5166), .ZN(n5138) );
  NAND2_X1 U6569 ( .A1(n5138), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5157) );
  INV_X1 U6570 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5139) );
  NAND2_X1 U6571 ( .A1(n5157), .A2(n5139), .ZN(n5140) );
  NAND2_X1 U6572 ( .A1(n5140), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5142) );
  INV_X1 U6573 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5141) );
  NOR2_X1 U6574 ( .A1(P2_IR_REG_23__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), .ZN(
        n5146) );
  NOR2_X1 U6575 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n5145) );
  NOR2_X1 U6576 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n5144) );
  NOR2_X1 U6577 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .ZN(
        n5143) );
  NAND2_X1 U6578 ( .A1(n5149), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5148) );
  MUX2_X1 U6579 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5148), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n5152) );
  INV_X1 U6580 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5150) );
  NAND2_X1 U6581 ( .A1(n5152), .A2(n5200), .ZN(n7513) );
  NAND2_X1 U6582 ( .A1(n5153), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5155) );
  MUX2_X1 U6583 ( .A(n5155), .B(P2_IR_REG_31__SCAN_IN), .S(n5154), .Z(n5156)
         );
  NAND2_X1 U6584 ( .A1(n5156), .A2(n5149), .ZN(n7458) );
  OR2_X1 U6585 ( .A1(n5598), .A2(P2_U3152), .ZN(n5832) );
  XNOR2_X1 U6586 ( .A(n5157), .B(P2_IR_REG_23__SCAN_IN), .ZN(n5814) );
  INV_X2 U6587 ( .A(n8412), .ZN(P2_U3966) );
  NAND2_X1 U6588 ( .A1(n5205), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5159) );
  AND2_X2 U6589 ( .A1(n8870), .A2(n5161), .ZN(n5231) );
  NAND2_X1 U6590 ( .A1(n5231), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5165) );
  NAND2_X1 U6591 ( .A1(n5802), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5164) );
  XNOR2_X1 U6592 ( .A(n5322), .B(P2_REG3_REG_6__SCAN_IN), .ZN(n7604) );
  NAND2_X1 U6593 ( .A1(n5245), .A2(n7604), .ZN(n5163) );
  NAND2_X1 U6594 ( .A1(n7670), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5162) );
  NAND4_X1 U6595 ( .A1(n5165), .A2(n5164), .A3(n5163), .A4(n5162), .ZN(n8422)
         );
  XNOR2_X1 U6596 ( .A(n5167), .B(n5166), .ZN(n5589) );
  INV_X1 U6597 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5169) );
  INV_X1 U6598 ( .A(n5212), .ZN(n5588) );
  NAND2_X1 U6599 ( .A1(n5171), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5172) );
  XNOR2_X1 U6600 ( .A(n5172), .B(P2_IR_REG_20__SCAN_IN), .ZN(n8398) );
  NAND2_X1 U6601 ( .A1(n5174), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5176) );
  NAND2_X1 U6602 ( .A1(n8422), .A2(n8016), .ZN(n5306) );
  INV_X1 U6603 ( .A(n5306), .ZN(n5309) );
  NAND2_X1 U6604 ( .A1(n5180), .A2(SI_0_), .ZN(n6143) );
  AND2_X1 U6605 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n5178) );
  NAND2_X1 U6606 ( .A1(n8185), .A2(n5178), .ZN(n5243) );
  INV_X1 U6607 ( .A(SI_1_), .ZN(n5179) );
  XNOR2_X1 U6608 ( .A(n5181), .B(n5179), .ZN(n5238) );
  BUF_X8 U6609 ( .A(n5180), .Z(n7590) );
  NAND2_X1 U6610 ( .A1(n5181), .A2(SI_1_), .ZN(n5182) );
  NAND2_X1 U6611 ( .A1(n5183), .A2(n5182), .ZN(n5255) );
  INV_X1 U6612 ( .A(SI_2_), .ZN(n5186) );
  XNOR2_X1 U6613 ( .A(n5187), .B(n5186), .ZN(n5254) );
  NAND2_X1 U6614 ( .A1(n5255), .A2(n5254), .ZN(n5189) );
  NAND2_X1 U6615 ( .A1(n5187), .A2(SI_2_), .ZN(n5188) );
  INV_X1 U6616 ( .A(SI_3_), .ZN(n5190) );
  XNOR2_X1 U6617 ( .A(n5191), .B(n5190), .ZN(n5274) );
  NAND2_X1 U6618 ( .A1(n5191), .A2(SI_3_), .ZN(n5192) );
  INV_X1 U6619 ( .A(SI_4_), .ZN(n5193) );
  NAND2_X1 U6620 ( .A1(n5194), .A2(SI_4_), .ZN(n5195) );
  INV_X1 U6621 ( .A(SI_5_), .ZN(n5197) );
  NAND2_X1 U6622 ( .A1(n5198), .A2(SI_5_), .ZN(n5199) );
  MUX2_X1 U6623 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n7590), .Z(n5312) );
  INV_X1 U6624 ( .A(SI_6_), .ZN(n10082) );
  XNOR2_X1 U6625 ( .A(n5311), .B(n5310), .ZN(n6583) );
  MUX2_X2 U6626 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5204), .S(
        P2_IR_REG_28__SCAN_IN), .Z(n5206) );
  OR2_X1 U6627 ( .A1(n6583), .A2(n5295), .ZN(n5211) );
  INV_X1 U6628 ( .A(n5843), .ZN(n5259) );
  INV_X1 U6629 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5207) );
  NAND2_X1 U6630 ( .A1(n5218), .A2(n5207), .ZN(n5343) );
  NAND2_X1 U6631 ( .A1(n5343), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5296) );
  INV_X1 U6632 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5208) );
  NAND2_X1 U6633 ( .A1(n5296), .A2(n5208), .ZN(n5209) );
  NAND2_X1 U6634 ( .A1(n5209), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5315) );
  XNOR2_X1 U6635 ( .A(n5315), .B(P2_IR_REG_6__SCAN_IN), .ZN(n5916) );
  AOI22_X1 U6636 ( .A1(n4479), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n5815), .B2(
        n5916), .ZN(n5210) );
  NAND2_X1 U6637 ( .A1(n5211), .A2(n5210), .ZN(n6813) );
  NAND2_X1 U6638 ( .A1(n5212), .A2(n8517), .ZN(n6037) );
  NAND2_X1 U6639 ( .A1(n6037), .A2(n8395), .ZN(n5215) );
  XNOR2_X1 U6640 ( .A(n6813), .B(n8007), .ZN(n5308) );
  OR2_X1 U6641 ( .A1(n5218), .A2(n8865), .ZN(n5219) );
  XNOR2_X1 U6642 ( .A(n5219), .B(P2_IR_REG_4__SCAN_IN), .ZN(n5849) );
  NAND2_X1 U6643 ( .A1(n5815), .A2(n5849), .ZN(n5221) );
  NAND2_X1 U6644 ( .A1(n4479), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n5220) );
  NAND2_X1 U6645 ( .A1(n5802), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5229) );
  INV_X1 U6646 ( .A(n5298), .ZN(n5224) );
  INV_X1 U6647 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n5283) );
  INV_X1 U6648 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n5222) );
  NAND2_X1 U6649 ( .A1(n5283), .A2(n5222), .ZN(n5223) );
  NAND2_X1 U6650 ( .A1(n5224), .A2(n5223), .ZN(n7083) );
  INV_X1 U6651 ( .A(n7083), .ZN(n5225) );
  NAND2_X1 U6652 ( .A1(n5245), .A2(n5225), .ZN(n5228) );
  NAND2_X1 U6653 ( .A1(n5284), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5227) );
  NAND2_X1 U6654 ( .A1(n5231), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5226) );
  NAND4_X1 U6655 ( .A1(n5229), .A2(n5228), .A3(n5227), .A4(n5226), .ZN(n8424)
         );
  NAND2_X1 U6656 ( .A1(n8424), .A2(n8016), .ZN(n5292) );
  NOR2_X1 U6657 ( .A1(n5233), .A2(n5232), .ZN(n5237) );
  NAND2_X1 U6658 ( .A1(n5245), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n5235) );
  NAND2_X1 U6659 ( .A1(n5246), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5234) );
  AND2_X1 U6660 ( .A1(n5235), .A2(n5234), .ZN(n5236) );
  NAND2_X1 U6661 ( .A1(n5259), .A2(n6005), .ZN(n5239) );
  OAI211_X2 U6662 ( .C1(n5295), .C2(n6305), .A(n5240), .B(n5239), .ZN(n6042)
         );
  NAND2_X1 U6663 ( .A1(n8185), .A2(SI_0_), .ZN(n5242) );
  INV_X1 U6664 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5241) );
  NAND2_X1 U6665 ( .A1(n5242), .A2(n5241), .ZN(n5244) );
  AND2_X1 U6666 ( .A1(n5244), .A2(n5243), .ZN(n8873) );
  NAND2_X1 U6667 ( .A1(n5245), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n5250) );
  NAND2_X1 U6668 ( .A1(n5230), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5249) );
  NAND2_X1 U6669 ( .A1(n5246), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5248) );
  NAND2_X1 U6670 ( .A1(n5231), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5247) );
  NAND4_X1 U6671 ( .A1(n5250), .A2(n5249), .A3(n5248), .A4(n5247), .ZN(n6047)
         );
  NAND2_X1 U6672 ( .A1(n6047), .A2(n7120), .ZN(n6043) );
  AOI21_X1 U6673 ( .B1(n5263), .B2(n10465), .A(n6102), .ZN(n7689) );
  INV_X1 U6674 ( .A(n5252), .ZN(n8056) );
  NAND2_X1 U6675 ( .A1(n8058), .A2(n5253), .ZN(n5269) );
  XNOR2_X1 U6676 ( .A(n5254), .B(n5255), .ZN(n6301) );
  INV_X1 U6677 ( .A(n6301), .ZN(n5256) );
  NAND2_X1 U6678 ( .A1(n5313), .A2(n5256), .ZN(n5262) );
  NAND2_X1 U6679 ( .A1(n4479), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n5261) );
  OR2_X1 U6680 ( .A1(n5258), .A2(n8865), .ZN(n5277) );
  XNOR2_X1 U6681 ( .A(n5277), .B(P2_IR_REG_2__SCAN_IN), .ZN(n5855) );
  NAND2_X1 U6682 ( .A1(n5259), .A2(n5855), .ZN(n5260) );
  AND3_X2 U6683 ( .A1(n5262), .A2(n5261), .A3(n5260), .ZN(n8063) );
  NAND2_X1 U6684 ( .A1(n5245), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n5267) );
  NAND2_X1 U6685 ( .A1(n5802), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5266) );
  NAND2_X1 U6686 ( .A1(n5284), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5265) );
  NAND2_X1 U6687 ( .A1(n5231), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5264) );
  NAND4_X2 U6688 ( .A1(n5267), .A2(n5266), .A3(n5265), .A4(n5264), .ZN(n6179)
         );
  NAND2_X1 U6689 ( .A1(n6179), .A2(n5268), .ZN(n5270) );
  XNOR2_X1 U6690 ( .A(n5271), .B(n5270), .ZN(n8059) );
  XNOR2_X1 U6691 ( .A(n5275), .B(n5274), .ZN(n6398) );
  NAND2_X1 U6692 ( .A1(n4479), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n5281) );
  INV_X1 U6693 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5276) );
  NAND2_X1 U6694 ( .A1(n5277), .A2(n5276), .ZN(n5278) );
  NAND2_X1 U6695 ( .A1(n5278), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5279) );
  XNOR2_X1 U6696 ( .A(n5279), .B(P2_IR_REG_3__SCAN_IN), .ZN(n8427) );
  NAND2_X1 U6697 ( .A1(n5815), .A2(n8427), .ZN(n5280) );
  AND3_X2 U6698 ( .A1(n5282), .A2(n5281), .A3(n5280), .ZN(n10471) );
  XNOR2_X1 U6699 ( .A(n5263), .B(n10471), .ZN(n6216) );
  NAND2_X1 U6700 ( .A1(n5802), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5288) );
  NAND2_X1 U6701 ( .A1(n5245), .A2(n5283), .ZN(n5286) );
  NAND2_X1 U6702 ( .A1(n5284), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5285) );
  NAND4_X1 U6703 ( .A1(n5288), .A2(n5287), .A3(n5286), .A4(n5285), .ZN(n8425)
         );
  AND2_X1 U6704 ( .A1(n8425), .A2(n8016), .ZN(n5289) );
  NAND2_X1 U6705 ( .A1(n6216), .A2(n5289), .ZN(n5290) );
  OAI21_X1 U6706 ( .B1(n6216), .B2(n5289), .A(n5290), .ZN(n6184) );
  INV_X1 U6707 ( .A(n5290), .ZN(n5291) );
  XNOR2_X1 U6708 ( .A(n5296), .B(P2_IR_REG_5__SCAN_IN), .ZN(n5884) );
  AOI22_X1 U6709 ( .A1(n4479), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n5815), .B2(
        n5884), .ZN(n5297) );
  XNOR2_X1 U6710 ( .A(n10444), .B(n5263), .ZN(n5303) );
  NAND2_X1 U6711 ( .A1(n5231), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5302) );
  NAND2_X1 U6712 ( .A1(n5802), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5301) );
  OAI21_X1 U6713 ( .B1(n5298), .B2(P2_REG3_REG_5__SCAN_IN), .A(n5322), .ZN(
        n6225) );
  INV_X1 U6714 ( .A(n6225), .ZN(n10446) );
  NAND2_X1 U6715 ( .A1(n5245), .A2(n10446), .ZN(n5300) );
  NAND2_X1 U6716 ( .A1(n5284), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5299) );
  NAND4_X1 U6717 ( .A1(n5302), .A2(n5301), .A3(n5300), .A4(n5299), .ZN(n8423)
         );
  NAND2_X1 U6718 ( .A1(n8423), .A2(n8016), .ZN(n5304) );
  XNOR2_X1 U6719 ( .A(n5303), .B(n5304), .ZN(n6231) );
  INV_X1 U6720 ( .A(n5303), .ZN(n7612) );
  INV_X1 U6721 ( .A(n5304), .ZN(n5305) );
  NOR2_X1 U6722 ( .A1(n7612), .A2(n5305), .ZN(n5307) );
  XNOR2_X1 U6723 ( .A(n5308), .B(n5306), .ZN(n7613) );
  MUX2_X1 U6724 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n7590), .Z(n5334) );
  XNOR2_X1 U6725 ( .A(n5333), .B(n5331), .ZN(n6716) );
  NAND2_X1 U6726 ( .A1(n6716), .A2(n8189), .ZN(n5319) );
  INV_X1 U6727 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5314) );
  NAND2_X1 U6728 ( .A1(n5315), .A2(n5314), .ZN(n5316) );
  NAND2_X1 U6729 ( .A1(n5316), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5317) );
  XNOR2_X1 U6730 ( .A(n5317), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6168) );
  AOI22_X1 U6731 ( .A1(n4479), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n5815), .B2(
        n6168), .ZN(n5318) );
  NAND2_X1 U6732 ( .A1(n5319), .A2(n5318), .ZN(n6866) );
  XNOR2_X1 U6733 ( .A(n6866), .B(n8007), .ZN(n6665) );
  INV_X1 U6734 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6820) );
  OR2_X1 U6735 ( .A1(n7673), .A2(n6820), .ZN(n5328) );
  NAND2_X1 U6736 ( .A1(n5802), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5327) );
  INV_X1 U6737 ( .A(n5322), .ZN(n5320) );
  AOI21_X1 U6738 ( .B1(n5320), .B2(P2_REG3_REG_6__SCAN_IN), .A(
        P2_REG3_REG_7__SCAN_IN), .ZN(n5323) );
  NAND2_X1 U6739 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(P2_REG3_REG_6__SCAN_IN), 
        .ZN(n5321) );
  OR2_X1 U6740 ( .A1(n5323), .A2(n5347), .ZN(n6824) );
  INV_X1 U6741 ( .A(n6824), .ZN(n5324) );
  NAND2_X1 U6742 ( .A1(n5245), .A2(n5324), .ZN(n5326) );
  NAND2_X1 U6743 ( .A1(n5284), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5325) );
  NAND4_X1 U6744 ( .A1(n5328), .A2(n5327), .A3(n5326), .A4(n5325), .ZN(n8421)
         );
  AND2_X1 U6745 ( .A1(n8421), .A2(n8016), .ZN(n5329) );
  NAND2_X1 U6746 ( .A1(n6665), .A2(n5329), .ZN(n5330) );
  OAI21_X1 U6747 ( .B1(n6665), .B2(n5329), .A(n5330), .ZN(n5612) );
  INV_X1 U6748 ( .A(n5330), .ZN(n5357) );
  NAND2_X1 U6749 ( .A1(n5333), .A2(n5332), .ZN(n5336) );
  NAND2_X1 U6750 ( .A1(n5334), .A2(SI_7_), .ZN(n5335) );
  INV_X1 U6751 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n5813) );
  INV_X1 U6752 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n5811) );
  MUX2_X1 U6753 ( .A(n5813), .B(n5811), .S(n7590), .Z(n5337) );
  INV_X1 U6754 ( .A(SI_8_), .ZN(n10147) );
  INV_X1 U6755 ( .A(n5337), .ZN(n5338) );
  NAND2_X1 U6756 ( .A1(n5338), .A2(SI_8_), .ZN(n5339) );
  XNOR2_X1 U6757 ( .A(n5359), .B(n5358), .ZN(n6841) );
  NAND2_X1 U6758 ( .A1(n6841), .A2(n8189), .ZN(n5346) );
  NAND2_X1 U6759 ( .A1(n5340), .A2(n5341), .ZN(n5342) );
  OR2_X1 U6760 ( .A1(n5343), .A2(n5342), .ZN(n5364) );
  NAND2_X1 U6761 ( .A1(n5364), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5344) );
  XNOR2_X1 U6762 ( .A(n5344), .B(P2_IR_REG_8__SCAN_IN), .ZN(n6348) );
  AOI22_X1 U6763 ( .A1(n4479), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n5815), .B2(
        n6348), .ZN(n5345) );
  XNOR2_X1 U6764 ( .A(n6960), .B(n8007), .ZN(n5353) );
  INV_X1 U6765 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n6898) );
  OR2_X1 U6766 ( .A1(n7673), .A2(n6898), .ZN(n5352) );
  NAND2_X1 U6767 ( .A1(n5802), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5351) );
  NAND2_X1 U6768 ( .A1(n5347), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5369) );
  OR2_X1 U6769 ( .A1(n5347), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5348) );
  AND2_X1 U6770 ( .A1(n5369), .A2(n5348), .ZN(n6659) );
  NAND2_X1 U6771 ( .A1(n5245), .A2(n6659), .ZN(n5350) );
  NAND2_X1 U6772 ( .A1(n7670), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5349) );
  NAND4_X1 U6773 ( .A1(n5352), .A2(n5351), .A3(n5350), .A4(n5349), .ZN(n8420)
         );
  AND2_X1 U6774 ( .A1(n8420), .A2(n8016), .ZN(n5354) );
  NAND2_X1 U6775 ( .A1(n5353), .A2(n5354), .ZN(n5375) );
  INV_X1 U6776 ( .A(n5353), .ZN(n8118) );
  INV_X1 U6777 ( .A(n5354), .ZN(n5355) );
  NAND2_X1 U6778 ( .A1(n8118), .A2(n5355), .ZN(n5356) );
  AND2_X1 U6779 ( .A1(n5375), .A2(n5356), .ZN(n6666) );
  INV_X1 U6780 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n5824) );
  MUX2_X1 U6781 ( .A(n5824), .B(n9902), .S(n7590), .Z(n5361) );
  INV_X1 U6782 ( .A(SI_9_), .ZN(n9892) );
  NAND2_X1 U6783 ( .A1(n5361), .A2(n9892), .ZN(n5404) );
  INV_X1 U6784 ( .A(n5361), .ZN(n5362) );
  NAND2_X1 U6785 ( .A1(n5362), .A2(SI_9_), .ZN(n5363) );
  XNOR2_X1 U6786 ( .A(n5382), .B(n5381), .ZN(n6906) );
  NAND2_X1 U6787 ( .A1(n6906), .A2(n8189), .ZN(n5366) );
  NOR2_X1 U6788 ( .A1(n5364), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n5438) );
  OR2_X1 U6789 ( .A1(n5438), .A2(n8865), .ZN(n5388) );
  XNOR2_X1 U6790 ( .A(n5388), .B(P2_IR_REG_9__SCAN_IN), .ZN(n6650) );
  AOI22_X1 U6791 ( .A1(n4479), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n5815), .B2(
        n6650), .ZN(n5365) );
  XNOR2_X1 U6792 ( .A(n8116), .B(n8007), .ZN(n5379) );
  INV_X1 U6793 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n5367) );
  OR2_X1 U6794 ( .A1(n7673), .A2(n5367), .ZN(n5374) );
  NAND2_X1 U6795 ( .A1(n5802), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5373) );
  NAND2_X1 U6796 ( .A1(n5369), .A2(n5368), .ZN(n5370) );
  AND2_X1 U6797 ( .A1(n5395), .A2(n5370), .ZN(n10437) );
  NAND2_X1 U6798 ( .A1(n5245), .A2(n10437), .ZN(n5372) );
  NAND2_X1 U6799 ( .A1(n7670), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5371) );
  NAND4_X1 U6800 ( .A1(n5374), .A2(n5373), .A3(n5372), .A4(n5371), .ZN(n8419)
         );
  NAND2_X1 U6801 ( .A1(n8419), .A2(n8016), .ZN(n5377) );
  XNOR2_X1 U6802 ( .A(n5379), .B(n5377), .ZN(n8117) );
  AND2_X1 U6803 ( .A1(n8117), .A2(n5375), .ZN(n5376) );
  INV_X1 U6804 ( .A(n5377), .ZN(n5378) );
  OR2_X1 U6805 ( .A1(n5379), .A2(n5378), .ZN(n5380) );
  NAND2_X1 U6806 ( .A1(n5405), .A2(n5404), .ZN(n5386) );
  INV_X1 U6807 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n5831) );
  MUX2_X1 U6808 ( .A(n5831), .B(n10063), .S(n7590), .Z(n5383) );
  INV_X1 U6809 ( .A(SI_10_), .ZN(n10080) );
  NAND2_X1 U6810 ( .A1(n5383), .A2(n10080), .ZN(n5403) );
  INV_X1 U6811 ( .A(n5383), .ZN(n5384) );
  NAND2_X1 U6812 ( .A1(n5384), .A2(SI_10_), .ZN(n5425) );
  AND2_X1 U6813 ( .A1(n5403), .A2(n5425), .ZN(n5385) );
  NAND2_X1 U6814 ( .A1(n7001), .A2(n8189), .ZN(n5393) );
  INV_X1 U6815 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5436) );
  AOI21_X1 U6816 ( .B1(n5388), .B2(n5436), .A(n8865), .ZN(n5389) );
  NAND2_X1 U6817 ( .A1(n5389), .A2(P2_IR_REG_10__SCAN_IN), .ZN(n5391) );
  INV_X1 U6818 ( .A(n5389), .ZN(n5390) );
  INV_X1 U6819 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5435) );
  NAND2_X1 U6820 ( .A1(n5390), .A2(n5435), .ZN(n5408) );
  AND2_X1 U6821 ( .A1(n5391), .A2(n5408), .ZN(n7036) );
  AOI22_X1 U6822 ( .A1(n5387), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n5815), .B2(
        n7036), .ZN(n5392) );
  XNOR2_X1 U6823 ( .A(n7157), .B(n8007), .ZN(n7103) );
  INV_X1 U6824 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n5394) );
  OR2_X1 U6825 ( .A1(n7673), .A2(n5394), .ZN(n5400) );
  NAND2_X1 U6826 ( .A1(n5802), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5399) );
  AND2_X1 U6827 ( .A1(n5395), .A2(n10062), .ZN(n5396) );
  NOR2_X1 U6828 ( .A1(n5412), .A2(n5396), .ZN(n7058) );
  NAND2_X1 U6829 ( .A1(n5245), .A2(n7058), .ZN(n5398) );
  NAND2_X1 U6830 ( .A1(n7670), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5397) );
  NAND4_X1 U6831 ( .A1(n5400), .A2(n5399), .A3(n5398), .A4(n5397), .ZN(n8418)
         );
  AND2_X1 U6832 ( .A1(n8418), .A2(n8016), .ZN(n5401) );
  NAND2_X1 U6833 ( .A1(n7103), .A2(n5401), .ZN(n5402) );
  OAI21_X1 U6834 ( .B1(n7103), .B2(n5401), .A(n5402), .ZN(n7064) );
  INV_X1 U6835 ( .A(n5402), .ZN(n5423) );
  AND2_X1 U6836 ( .A1(n5477), .A2(n5425), .ZN(n5407) );
  MUX2_X1 U6837 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .S(n7590), .Z(n5424) );
  INV_X1 U6838 ( .A(SI_11_), .ZN(n5406) );
  XNOR2_X1 U6839 ( .A(n5424), .B(n5406), .ZN(n5426) );
  XNOR2_X1 U6840 ( .A(n5407), .B(n5426), .ZN(n7184) );
  NAND2_X1 U6841 ( .A1(n7184), .A2(n8189), .ZN(n5411) );
  NAND2_X1 U6842 ( .A1(n5408), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5409) );
  XNOR2_X1 U6843 ( .A(n5409), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7217) );
  AOI22_X1 U6844 ( .A1(n5387), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n5815), .B2(
        n7217), .ZN(n5410) );
  XNOR2_X1 U6845 ( .A(n8722), .B(n8007), .ZN(n5419) );
  NAND2_X1 U6846 ( .A1(n5231), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n5418) );
  NAND2_X1 U6847 ( .A1(n5802), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5417) );
  NOR2_X1 U6848 ( .A1(n5412), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5413) );
  OR2_X1 U6849 ( .A1(n5442), .A2(n5413), .ZN(n8719) );
  INV_X1 U6850 ( .A(n8719), .ZN(n5414) );
  NAND2_X1 U6851 ( .A1(n7667), .A2(n5414), .ZN(n5416) );
  NAND2_X1 U6852 ( .A1(n7670), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5415) );
  NAND4_X1 U6853 ( .A1(n5418), .A2(n5417), .A3(n5416), .A4(n5415), .ZN(n8417)
         );
  AND2_X1 U6854 ( .A1(n8417), .A2(n8016), .ZN(n5420) );
  NAND2_X1 U6855 ( .A1(n5419), .A2(n5420), .ZN(n5448) );
  INV_X1 U6856 ( .A(n5419), .ZN(n7069) );
  INV_X1 U6857 ( .A(n5420), .ZN(n5421) );
  NAND2_X1 U6858 ( .A1(n7069), .A2(n5421), .ZN(n5422) );
  AND2_X1 U6859 ( .A1(n5448), .A2(n5422), .ZN(n7104) );
  NAND2_X1 U6860 ( .A1(n5424), .A2(SI_11_), .ZN(n5428) );
  INV_X1 U6861 ( .A(n5426), .ZN(n5427) );
  INV_X1 U6862 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n5430) );
  MUX2_X1 U6863 ( .A(n5430), .B(n9876), .S(n7590), .Z(n5431) );
  INV_X1 U6864 ( .A(SI_12_), .ZN(n10150) );
  NAND2_X1 U6865 ( .A1(n5431), .A2(n10150), .ZN(n5478) );
  INV_X1 U6866 ( .A(n5431), .ZN(n5432) );
  NAND2_X1 U6867 ( .A1(n5432), .A2(SI_12_), .ZN(n5433) );
  XNOR2_X1 U6868 ( .A(n5454), .B(n5471), .ZN(n7282) );
  NAND2_X1 U6869 ( .A1(n7282), .A2(n8189), .ZN(n5441) );
  INV_X1 U6870 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5434) );
  AND3_X1 U6871 ( .A1(n5436), .A2(n5435), .A3(n5434), .ZN(n5437) );
  AND2_X1 U6872 ( .A1(n5438), .A2(n5437), .ZN(n5460) );
  OR2_X1 U6873 ( .A1(n5460), .A2(n8865), .ZN(n5439) );
  XNOR2_X1 U6874 ( .A(n5439), .B(P2_IR_REG_12__SCAN_IN), .ZN(n8440) );
  AOI22_X1 U6875 ( .A1(n5387), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n5815), .B2(
        n8440), .ZN(n5440) );
  XNOR2_X1 U6876 ( .A(n7395), .B(n8007), .ZN(n5452) );
  INV_X1 U6877 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7237) );
  OR2_X1 U6878 ( .A1(n7673), .A2(n7237), .ZN(n5447) );
  NAND2_X1 U6879 ( .A1(n7669), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5446) );
  OR2_X1 U6880 ( .A1(n5442), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5443) );
  AND2_X1 U6881 ( .A1(n5463), .A2(n5443), .ZN(n7233) );
  NAND2_X1 U6882 ( .A1(n7667), .A2(n7233), .ZN(n5445) );
  NAND2_X1 U6883 ( .A1(n5284), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5444) );
  NAND4_X1 U6884 ( .A1(n5447), .A2(n5446), .A3(n5445), .A4(n5444), .ZN(n10217)
         );
  NAND2_X1 U6885 ( .A1(n10217), .A2(n8016), .ZN(n5450) );
  XNOR2_X1 U6886 ( .A(n5452), .B(n5450), .ZN(n7081) );
  INV_X1 U6887 ( .A(n5450), .ZN(n5451) );
  MUX2_X1 U6888 ( .A(n6062), .B(n9943), .S(n7590), .Z(n5456) );
  INV_X1 U6889 ( .A(SI_13_), .ZN(n5455) );
  NAND2_X1 U6890 ( .A1(n5456), .A2(n5455), .ZN(n5481) );
  INV_X1 U6891 ( .A(n5456), .ZN(n5457) );
  NAND2_X1 U6892 ( .A1(n5457), .A2(SI_13_), .ZN(n5458) );
  NAND2_X1 U6893 ( .A1(n5460), .A2(n5459), .ZN(n5548) );
  NAND2_X1 U6894 ( .A1(n5548), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5482) );
  XNOR2_X1 U6895 ( .A(n5482), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7353) );
  AOI22_X1 U6896 ( .A1(n5387), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n5815), .B2(
        n7353), .ZN(n5461) );
  NAND2_X2 U6897 ( .A1(n5462), .A2(n5461), .ZN(n10227) );
  XNOR2_X1 U6898 ( .A(n10227), .B(n5263), .ZN(n7337) );
  INV_X1 U6899 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n10210) );
  OR2_X1 U6900 ( .A1(n7673), .A2(n10210), .ZN(n5468) );
  NAND2_X1 U6901 ( .A1(n5802), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n5467) );
  INV_X1 U6902 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n7222) );
  NAND2_X1 U6903 ( .A1(n5463), .A2(n7222), .ZN(n5464) );
  AND2_X1 U6904 ( .A1(n5487), .A2(n5464), .ZN(n7174) );
  NAND2_X1 U6905 ( .A1(n7667), .A2(n7174), .ZN(n5466) );
  NAND2_X1 U6906 ( .A1(n5284), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5465) );
  NAND4_X1 U6907 ( .A1(n5468), .A2(n5467), .A3(n5466), .A4(n5465), .ZN(n8416)
         );
  NAND2_X1 U6908 ( .A1(n8416), .A2(n8016), .ZN(n5469) );
  NOR2_X1 U6909 ( .A1(n7337), .A2(n5469), .ZN(n5493) );
  MUX2_X1 U6910 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n7590), .Z(n5501) );
  INV_X1 U6911 ( .A(SI_14_), .ZN(n10068) );
  XNOR2_X1 U6912 ( .A(n5504), .B(n5500), .ZN(n7410) );
  NAND2_X1 U6913 ( .A1(n7410), .A2(n8189), .ZN(n5485) );
  INV_X1 U6914 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5546) );
  NAND2_X1 U6915 ( .A1(n5482), .A2(n5546), .ZN(n5483) );
  NAND2_X1 U6916 ( .A1(n5483), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5510) );
  XNOR2_X1 U6917 ( .A(n5510), .B(P2_IR_REG_14__SCAN_IN), .ZN(n7555) );
  AOI22_X1 U6918 ( .A1(n5387), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n5815), .B2(
        n7555), .ZN(n5484) );
  XNOR2_X1 U6919 ( .A(n7462), .B(n8007), .ZN(n5498) );
  NAND2_X1 U6920 ( .A1(n7669), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n5492) );
  INV_X1 U6921 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n5486) );
  AND2_X1 U6922 ( .A1(n5487), .A2(n5486), .ZN(n5488) );
  OR2_X1 U6923 ( .A1(n5515), .A2(n5488), .ZN(n7341) );
  INV_X1 U6924 ( .A(n7341), .ZN(n7401) );
  NAND2_X1 U6925 ( .A1(n7667), .A2(n7401), .ZN(n5491) );
  NAND2_X1 U6926 ( .A1(n5284), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5490) );
  NAND2_X1 U6927 ( .A1(n5231), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n5489) );
  NAND4_X1 U6928 ( .A1(n5492), .A2(n5491), .A3(n5490), .A4(n5489), .ZN(n10218)
         );
  NAND2_X1 U6929 ( .A1(n10218), .A2(n8016), .ZN(n5496) );
  XNOR2_X1 U6930 ( .A(n5498), .B(n5496), .ZN(n7346) );
  INV_X1 U6931 ( .A(n5493), .ZN(n5494) );
  INV_X1 U6932 ( .A(n5496), .ZN(n5497) );
  NAND2_X1 U6933 ( .A1(n5501), .A2(SI_14_), .ZN(n5502) );
  INV_X1 U6934 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6189) );
  INV_X1 U6935 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n5505) );
  MUX2_X1 U6936 ( .A(n6189), .B(n5505), .S(n7590), .Z(n5506) );
  INV_X1 U6937 ( .A(n5506), .ZN(n5507) );
  NAND2_X1 U6938 ( .A1(n5507), .A2(SI_15_), .ZN(n5508) );
  XNOR2_X1 U6939 ( .A(n5538), .B(n5537), .ZN(n7713) );
  NAND2_X1 U6940 ( .A1(n7713), .A2(n8189), .ZN(n5514) );
  NAND2_X1 U6941 ( .A1(n5510), .A2(n5509), .ZN(n5511) );
  NAND2_X1 U6942 ( .A1(n5511), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5512) );
  XNOR2_X1 U6943 ( .A(n5512), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8464) );
  AOI22_X1 U6944 ( .A1(n5815), .A2(n8464), .B1(n5387), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n5513) );
  XNOR2_X1 U6945 ( .A(n8804), .B(n5263), .ZN(n5526) );
  NAND2_X1 U6946 ( .A1(n7669), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n5525) );
  NAND2_X1 U6947 ( .A1(n5515), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5530) );
  INV_X1 U6948 ( .A(n5515), .ZN(n5517) );
  INV_X1 U6949 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n5516) );
  NAND2_X1 U6950 ( .A1(n5517), .A2(n5516), .ZN(n5518) );
  NAND2_X1 U6951 ( .A1(n5530), .A2(n5518), .ZN(n10198) );
  INV_X1 U6952 ( .A(n10198), .ZN(n5519) );
  NAND2_X1 U6953 ( .A1(n7667), .A2(n5519), .ZN(n5524) );
  INV_X1 U6954 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n5521) );
  OR2_X1 U6955 ( .A1(n5520), .A2(n5521), .ZN(n5523) );
  INV_X1 U6956 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n7470) );
  OR2_X1 U6957 ( .A1(n7673), .A2(n7470), .ZN(n5522) );
  NOR2_X1 U6958 ( .A1(n7465), .A2(n8196), .ZN(n10190) );
  INV_X1 U6959 ( .A(n5530), .ZN(n5529) );
  NAND2_X1 U6960 ( .A1(n5529), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5564) );
  INV_X1 U6961 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n8461) );
  NAND2_X1 U6962 ( .A1(n5530), .A2(n8461), .ZN(n5531) );
  AND2_X1 U6963 ( .A1(n5564), .A2(n5531), .ZN(n7521) );
  NAND2_X1 U6964 ( .A1(n7521), .A2(n7667), .ZN(n5536) );
  INV_X1 U6965 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n5532) );
  OR2_X1 U6966 ( .A1(n7673), .A2(n5532), .ZN(n5535) );
  NAND2_X1 U6967 ( .A1(n7669), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n5534) );
  NAND2_X1 U6968 ( .A1(n7670), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5533) );
  NAND4_X1 U6969 ( .A1(n5536), .A2(n5535), .A3(n5534), .A4(n5533), .ZN(n8414)
         );
  NAND2_X1 U6970 ( .A1(n8414), .A2(n8016), .ZN(n5552) );
  INV_X1 U6971 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n5541) );
  INV_X1 U6972 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n5540) );
  MUX2_X1 U6973 ( .A(n5541), .B(n5540), .S(n7590), .Z(n5542) );
  INV_X1 U6974 ( .A(SI_16_), .ZN(n10133) );
  NAND2_X1 U6975 ( .A1(n5542), .A2(n10133), .ZN(n5557) );
  INV_X1 U6976 ( .A(n5542), .ZN(n5543) );
  NAND2_X1 U6977 ( .A1(n5543), .A2(SI_16_), .ZN(n5544) );
  XNOR2_X1 U6978 ( .A(n5556), .B(n5555), .ZN(n7725) );
  NAND2_X1 U6979 ( .A1(n7725), .A2(n8189), .ZN(n5551) );
  INV_X1 U6980 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5545) );
  NAND3_X1 U6981 ( .A1(n5546), .A2(n5509), .A3(n5545), .ZN(n5547) );
  OAI21_X1 U6982 ( .B1(n5548), .B2(n5547), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n5549) );
  XNOR2_X1 U6983 ( .A(n5549), .B(P2_IR_REG_16__SCAN_IN), .ZN(n8480) );
  AOI22_X1 U6984 ( .A1(n5387), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n5815), .B2(
        n8480), .ZN(n5550) );
  XNOR2_X1 U6985 ( .A(n8799), .B(n5263), .ZN(n5553) );
  NAND2_X1 U6986 ( .A1(n5553), .A2(n5552), .ZN(n5554) );
  MUX2_X1 U6987 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(P2_DATAO_REG_17__SCAN_IN), 
        .S(n7590), .Z(n5632) );
  INV_X1 U6988 ( .A(SI_17_), .ZN(n9906) );
  XNOR2_X1 U6989 ( .A(n5632), .B(n9906), .ZN(n5630) );
  XNOR2_X1 U6990 ( .A(n5629), .B(n5630), .ZN(n7747) );
  NAND2_X1 U6991 ( .A1(n7747), .A2(n8189), .ZN(n5563) );
  INV_X1 U6992 ( .A(n5147), .ZN(n5558) );
  NAND2_X1 U6993 ( .A1(n5558), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5559) );
  MUX2_X1 U6994 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5559), .S(
        P2_IR_REG_17__SCAN_IN), .Z(n5561) );
  NAND2_X1 U6995 ( .A1(n5561), .A2(n5560), .ZN(n8493) );
  INV_X1 U6996 ( .A(n8493), .ZN(n8499) );
  AOI22_X1 U6997 ( .A1(n5387), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n5815), .B2(
        n8499), .ZN(n5562) );
  XNOR2_X1 U6998 ( .A(n8794), .B(n8007), .ZN(n8141) );
  INV_X1 U6999 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8478) );
  NAND2_X1 U7000 ( .A1(n5564), .A2(n8478), .ZN(n5565) );
  NAND2_X1 U7001 ( .A1(n5604), .A2(n5565), .ZN(n7547) );
  INV_X1 U7002 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8494) );
  OR2_X1 U7003 ( .A1(n7673), .A2(n8494), .ZN(n5567) );
  NAND2_X1 U7004 ( .A1(n7669), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n5566) );
  AND2_X1 U7005 ( .A1(n5567), .A2(n5566), .ZN(n5569) );
  NAND2_X1 U7006 ( .A1(n7670), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5568) );
  OAI211_X1 U7007 ( .C1(n7547), .C2(n7625), .A(n5569), .B(n5568), .ZN(n8413)
         );
  AND2_X1 U7008 ( .A1(n8413), .A2(n8016), .ZN(n5570) );
  NAND2_X1 U7009 ( .A1(n8141), .A2(n5570), .ZN(n5627) );
  OAI21_X1 U7010 ( .B1(n8141), .B2(n5570), .A(n5627), .ZN(n5593) );
  INV_X1 U7011 ( .A(P2_B_REG_SCAN_IN), .ZN(n5571) );
  XOR2_X1 U7012 ( .A(n7367), .B(n5571), .Z(n5572) );
  INV_X1 U7013 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n10459) );
  AND2_X1 U7014 ( .A1(n7367), .A2(n7513), .ZN(n10460) );
  AOI21_X1 U7015 ( .B1(n10457), .B2(n10459), .A(n10460), .ZN(n6206) );
  NOR4_X1 U7016 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n5577) );
  NOR4_X1 U7017 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n5576) );
  NOR4_X1 U7018 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n5575) );
  NOR4_X1 U7019 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n5574) );
  NAND4_X1 U7020 ( .A1(n5577), .A2(n5576), .A3(n5575), .A4(n5574), .ZN(n5583)
         );
  NOR2_X1 U7021 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .ZN(
        n5581) );
  NOR4_X1 U7022 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n5580) );
  NOR4_X1 U7023 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n5579) );
  NOR4_X1 U7024 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n5578) );
  NAND4_X1 U7025 ( .A1(n5581), .A2(n5580), .A3(n5579), .A4(n5578), .ZN(n5582)
         );
  OAI21_X1 U7026 ( .B1(n5583), .B2(n5582), .A(n10457), .ZN(n6204) );
  INV_X1 U7027 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n10462) );
  AND2_X1 U7028 ( .A1(n7513), .A2(n7458), .ZN(n10464) );
  AOI21_X1 U7029 ( .B1(n10457), .B2(n10462), .A(n10464), .ZN(n6767) );
  AND2_X1 U7030 ( .A1(n6204), .A2(n6767), .ZN(n5584) );
  NAND2_X1 U7031 ( .A1(n6206), .A2(n5584), .ZN(n5596) );
  INV_X1 U7032 ( .A(n5596), .ZN(n5587) );
  NOR2_X1 U7033 ( .A1(n5814), .A2(P2_U3152), .ZN(n10463) );
  NAND2_X1 U7034 ( .A1(n5598), .A2(n10463), .ZN(n10458) );
  INV_X1 U7035 ( .A(n10458), .ZN(n5586) );
  NAND2_X1 U7036 ( .A1(n5587), .A2(n5586), .ZN(n5595) );
  INV_X1 U7037 ( .A(n5595), .ZN(n5601) );
  INV_X1 U7038 ( .A(n8803), .ZN(n10488) );
  INV_X1 U7039 ( .A(n4486), .ZN(n8402) );
  INV_X1 U7040 ( .A(n8395), .ZN(n8249) );
  INV_X1 U7041 ( .A(n6035), .ZN(n5817) );
  AND2_X1 U7042 ( .A1(n10488), .A2(n5817), .ZN(n5590) );
  INV_X1 U7043 ( .A(n5628), .ZN(n5592) );
  AOI211_X1 U7044 ( .C1(n5591), .C2(n5593), .A(n8156), .B(n5592), .ZN(n5611)
         );
  INV_X1 U7045 ( .A(n8794), .ZN(n7551) );
  OR2_X1 U7046 ( .A1(n10458), .A2(n8398), .ZN(n5594) );
  NAND2_X1 U7047 ( .A1(n5595), .A2(n5594), .ZN(n10192) );
  NAND2_X1 U7048 ( .A1(n10192), .A2(n8803), .ZN(n8167) );
  NOR2_X1 U7049 ( .A1(n7551), .A2(n8167), .ZN(n5610) );
  NAND2_X1 U7050 ( .A1(n5596), .A2(n6769), .ZN(n6099) );
  AOI21_X1 U7051 ( .B1(n6035), .B2(n8400), .A(n5814), .ZN(n5597) );
  AND2_X1 U7052 ( .A1(n5598), .A2(n5597), .ZN(n6098) );
  NAND2_X1 U7053 ( .A1(n6099), .A2(n6098), .ZN(n5599) );
  NAND2_X1 U7054 ( .A1(n5599), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10199) );
  OAI22_X1 U7055 ( .A1(n10199), .A2(n7547), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8478), .ZN(n5609) );
  INV_X1 U7056 ( .A(n8414), .ZN(n7544) );
  INV_X1 U7057 ( .A(n5602), .ZN(n7571) );
  NAND2_X1 U7058 ( .A1(n10188), .A2(n10216), .ZN(n8160) );
  AND2_X1 U7059 ( .A1(n6035), .A2(n5602), .ZN(n8701) );
  INV_X1 U7060 ( .A(n8701), .ZN(n10427) );
  NAND2_X1 U7061 ( .A1(n10188), .A2(n8701), .ZN(n8161) );
  INV_X1 U7062 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n8858) );
  INV_X1 U7063 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n8496) );
  NAND2_X1 U7064 ( .A1(n5604), .A2(n8496), .ZN(n5605) );
  NAND2_X1 U7065 ( .A1(n5654), .A2(n5605), .ZN(n8148) );
  OR2_X1 U7066 ( .A1(n8148), .A2(n7625), .ZN(n5607) );
  AOI22_X1 U7067 ( .A1(n5231), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n7669), .B2(
        P2_REG1_REG_18__SCAN_IN), .ZN(n5606) );
  OAI211_X1 U7068 ( .C1(n5520), .C2(n8858), .A(n5607), .B(n5606), .ZN(n8700)
         );
  INV_X1 U7069 ( .A(n8700), .ZN(n8086) );
  OAI22_X1 U7070 ( .A1(n7544), .A2(n8160), .B1(n8161), .B2(n8086), .ZN(n5608)
         );
  OR4_X1 U7071 ( .A1(n5611), .A2(n5610), .A3(n5609), .A4(n5608), .ZN(P2_U3230)
         );
  AOI211_X1 U7072 ( .C1(n5613), .C2(n5612), .A(n8156), .B(n6667), .ZN(n5617)
         );
  INV_X1 U7073 ( .A(n8422), .ZN(n6482) );
  NOR2_X1 U7074 ( .A1(n8160), .A2(n6482), .ZN(n5616) );
  INV_X1 U7075 ( .A(n8420), .ZN(n10430) );
  INV_X1 U7076 ( .A(n6866), .ZN(n10480) );
  OAI22_X1 U7077 ( .A1(n8161), .A2(n10430), .B1(n10480), .B2(n8167), .ZN(n5615) );
  INV_X1 U7078 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n9929) );
  OAI22_X1 U7079 ( .A1(n10199), .A2(n6824), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9929), .ZN(n5614) );
  OR4_X1 U7080 ( .A1(n5617), .A2(n5616), .A3(n5615), .A4(n5614), .ZN(P2_U3215)
         );
  OR2_X1 U7081 ( .A1(n8156), .A2(n8196), .ZN(n8142) );
  INV_X1 U7082 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n8085) );
  INV_X1 U7083 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n8093) );
  INV_X1 U7084 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n10069) );
  NAND2_X1 U7085 ( .A1(n5713), .A2(n10069), .ZN(n5620) );
  AND2_X1 U7086 ( .A1(n5737), .A2(n5620), .ZN(n8643) );
  NAND2_X1 U7087 ( .A1(n8643), .A2(n7667), .ZN(n5626) );
  INV_X1 U7088 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n5623) );
  NAND2_X1 U7089 ( .A1(n7670), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n5622) );
  NAND2_X1 U7090 ( .A1(n7669), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n5621) );
  OAI211_X1 U7091 ( .C1(n7673), .C2(n5623), .A(n5622), .B(n5621), .ZN(n5624)
         );
  INV_X1 U7092 ( .A(n5624), .ZN(n5625) );
  NOR2_X1 U7093 ( .A1(n8142), .A2(n8411), .ZN(n5734) );
  NOR2_X1 U7094 ( .A1(n8411), .A2(n8196), .ZN(n5748) );
  NOR2_X1 U7095 ( .A1(n5748), .A2(n8156), .ZN(n5733) );
  NAND2_X1 U7096 ( .A1(n5628), .A2(n5627), .ZN(n5638) );
  NAND2_X1 U7097 ( .A1(n5631), .A2(n5630), .ZN(n5634) );
  NAND2_X1 U7098 ( .A1(n5632), .A2(SI_17_), .ZN(n5633) );
  MUX2_X1 U7099 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n7590), .Z(n5646) );
  XNOR2_X1 U7100 ( .A(n5646), .B(SI_18_), .ZN(n5643) );
  XNOR2_X1 U7101 ( .A(n5645), .B(n5643), .ZN(n7766) );
  NAND2_X1 U7102 ( .A1(n7766), .A2(n8189), .ZN(n5637) );
  NAND2_X1 U7103 ( .A1(n5560), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5635) );
  XNOR2_X1 U7104 ( .A(n5635), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8512) );
  AOI22_X1 U7105 ( .A1(n5387), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n5815), .B2(
        n8512), .ZN(n5636) );
  XNOR2_X1 U7106 ( .A(n8788), .B(n8007), .ZN(n5641) );
  NAND2_X1 U7107 ( .A1(n8700), .A2(n8016), .ZN(n5639) );
  XNOR2_X1 U7108 ( .A(n5641), .B(n5639), .ZN(n8139) );
  INV_X1 U7109 ( .A(n5639), .ZN(n5640) );
  NAND2_X1 U7110 ( .A1(n5641), .A2(n5640), .ZN(n5642) );
  NAND2_X1 U7111 ( .A1(n5646), .A2(SI_18_), .ZN(n5647) );
  INV_X1 U7112 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n6684) );
  INV_X1 U7113 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n9907) );
  MUX2_X1 U7114 ( .A(n6684), .B(n9907), .S(n7590), .Z(n5649) );
  INV_X1 U7115 ( .A(SI_19_), .ZN(n10083) );
  NAND2_X1 U7116 ( .A1(n5649), .A2(n10083), .ZN(n5662) );
  INV_X1 U7117 ( .A(n5649), .ZN(n5650) );
  NAND2_X1 U7118 ( .A1(n5650), .A2(SI_19_), .ZN(n5651) );
  NAND2_X1 U7119 ( .A1(n5662), .A2(n5651), .ZN(n5663) );
  XNOR2_X1 U7120 ( .A(n5664), .B(n5663), .ZN(n7784) );
  NAND2_X1 U7121 ( .A1(n7784), .A2(n8189), .ZN(n5653) );
  INV_X1 U7122 ( .A(n8517), .ZN(n10449) );
  AOI22_X1 U7123 ( .A1(n5387), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n5815), .B2(
        n10449), .ZN(n5652) );
  XNOR2_X1 U7124 ( .A(n8783), .B(n5263), .ZN(n5658) );
  NAND2_X1 U7125 ( .A1(n5654), .A2(n8085), .ZN(n5655) );
  NAND2_X1 U7126 ( .A1(n5670), .A2(n5655), .ZN(n8709) );
  AOI22_X1 U7127 ( .A1(n5231), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n7669), .B2(
        P2_REG1_REG_19__SCAN_IN), .ZN(n5657) );
  NAND2_X1 U7128 ( .A1(n7670), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n5656) );
  OAI211_X1 U7129 ( .C1(n8709), .C2(n7625), .A(n5657), .B(n5656), .ZN(n8686)
         );
  NAND2_X1 U7130 ( .A1(n8686), .A2(n8016), .ZN(n5659) );
  NAND2_X1 U7131 ( .A1(n5658), .A2(n5659), .ZN(n8082) );
  INV_X1 U7132 ( .A(n5658), .ZN(n5661) );
  INV_X1 U7133 ( .A(n5659), .ZN(n5660) );
  NAND2_X1 U7134 ( .A1(n5661), .A2(n5660), .ZN(n8081) );
  INV_X1 U7135 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n6988) );
  INV_X1 U7136 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n10077) );
  MUX2_X1 U7137 ( .A(n6988), .B(n10077), .S(n7590), .Z(n5665) );
  INV_X1 U7138 ( .A(SI_20_), .ZN(n10135) );
  NAND2_X1 U7139 ( .A1(n5665), .A2(n10135), .ZN(n5684) );
  INV_X1 U7140 ( .A(n5665), .ZN(n5666) );
  NAND2_X1 U7141 ( .A1(n5666), .A2(SI_20_), .ZN(n5667) );
  XNOR2_X1 U7142 ( .A(n5683), .B(n5682), .ZN(n7802) );
  NAND2_X1 U7143 ( .A1(n7802), .A2(n8189), .ZN(n5669) );
  NAND2_X1 U7144 ( .A1(n5387), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n5668) );
  XNOR2_X1 U7145 ( .A(n8775), .B(n8007), .ZN(n5679) );
  INV_X1 U7146 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n9901) );
  NAND2_X1 U7147 ( .A1(n5670), .A2(n9901), .ZN(n5671) );
  NAND2_X1 U7148 ( .A1(n5688), .A2(n5671), .ZN(n8690) );
  OR2_X1 U7149 ( .A1(n8690), .A2(n7625), .ZN(n5676) );
  INV_X1 U7150 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8691) );
  NAND2_X1 U7151 ( .A1(n7669), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n5673) );
  NAND2_X1 U7152 ( .A1(n7670), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n5672) );
  OAI211_X1 U7153 ( .C1(n7673), .C2(n8691), .A(n5673), .B(n5672), .ZN(n5674)
         );
  INV_X1 U7154 ( .A(n5674), .ZN(n5675) );
  NAND2_X1 U7155 ( .A1(n5676), .A2(n5675), .ZN(n8702) );
  NAND2_X1 U7156 ( .A1(n8702), .A2(n8016), .ZN(n5677) );
  XNOR2_X1 U7157 ( .A(n5679), .B(n5677), .ZN(n8125) );
  NAND2_X1 U7158 ( .A1(n8124), .A2(n8125), .ZN(n5681) );
  INV_X1 U7159 ( .A(n5677), .ZN(n5678) );
  NAND2_X1 U7160 ( .A1(n5679), .A2(n5678), .ZN(n5680) );
  NAND2_X1 U7161 ( .A1(n5681), .A2(n5680), .ZN(n8091) );
  MUX2_X1 U7162 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n7590), .Z(n5701) );
  INV_X1 U7163 ( .A(SI_21_), .ZN(n5685) );
  XNOR2_X1 U7164 ( .A(n5701), .B(n5685), .ZN(n5700) );
  XNOR2_X1 U7165 ( .A(n5704), .B(n5700), .ZN(n7821) );
  NAND2_X1 U7166 ( .A1(n7821), .A2(n8189), .ZN(n5687) );
  NAND2_X1 U7167 ( .A1(n5387), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n5686) );
  XNOR2_X1 U7168 ( .A(n8843), .B(n8007), .ZN(n5696) );
  NAND2_X1 U7169 ( .A1(n5688), .A2(n8093), .ZN(n5689) );
  AND2_X1 U7170 ( .A1(n5711), .A2(n5689), .ZN(n8675) );
  NAND2_X1 U7171 ( .A1(n8675), .A2(n7667), .ZN(n5695) );
  INV_X1 U7172 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n5692) );
  NAND2_X1 U7173 ( .A1(n7670), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n5691) );
  NAND2_X1 U7174 ( .A1(n7669), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n5690) );
  OAI211_X1 U7175 ( .C1(n7673), .C2(n5692), .A(n5691), .B(n5690), .ZN(n5693)
         );
  INV_X1 U7176 ( .A(n5693), .ZN(n5694) );
  NAND2_X1 U7177 ( .A1(n5695), .A2(n5694), .ZN(n8687) );
  NAND2_X1 U7178 ( .A1(n8687), .A2(n8016), .ZN(n5697) );
  XNOR2_X1 U7179 ( .A(n5696), .B(n5697), .ZN(n8092) );
  INV_X1 U7180 ( .A(n5696), .ZN(n5698) );
  NOR2_X1 U7181 ( .A1(n5698), .A2(n5697), .ZN(n5699) );
  AOI21_X2 U7182 ( .B1(n8091), .B2(n8092), .A(n5699), .ZN(n5720) );
  INV_X1 U7183 ( .A(n5700), .ZN(n5703) );
  NAND2_X1 U7184 ( .A1(n5701), .A2(SI_21_), .ZN(n5702) );
  INV_X1 U7185 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7156) );
  INV_X1 U7186 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7842) );
  MUX2_X1 U7187 ( .A(n7156), .B(n7842), .S(n7590), .Z(n5706) );
  INV_X1 U7188 ( .A(SI_22_), .ZN(n5705) );
  NAND2_X1 U7189 ( .A1(n5706), .A2(n5705), .ZN(n5726) );
  INV_X1 U7190 ( .A(n5706), .ZN(n5707) );
  NAND2_X1 U7191 ( .A1(n5707), .A2(SI_22_), .ZN(n5708) );
  NAND2_X1 U7192 ( .A1(n5726), .A2(n5708), .ZN(n5724) );
  XNOR2_X1 U7193 ( .A(n5725), .B(n5724), .ZN(n7841) );
  NAND2_X1 U7194 ( .A1(n7841), .A2(n8189), .ZN(n5710) );
  NAND2_X1 U7195 ( .A1(n5387), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n5709) );
  XNOR2_X1 U7196 ( .A(n8662), .B(n8007), .ZN(n5721) );
  XNOR2_X1 U7197 ( .A(n5720), .B(n5721), .ZN(n8134) );
  INV_X1 U7198 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n9962) );
  NAND2_X1 U7199 ( .A1(n5711), .A2(n9962), .ZN(n5712) );
  NAND2_X1 U7200 ( .A1(n5713), .A2(n5712), .ZN(n8657) );
  OR2_X1 U7201 ( .A1(n8657), .A2(n7625), .ZN(n5718) );
  INV_X1 U7202 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n8658) );
  NAND2_X1 U7203 ( .A1(n7670), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n5715) );
  NAND2_X1 U7204 ( .A1(n7669), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n5714) );
  OAI211_X1 U7205 ( .C1(n7673), .C2(n8658), .A(n5715), .B(n5714), .ZN(n5716)
         );
  INV_X1 U7206 ( .A(n5716), .ZN(n5717) );
  NAND2_X1 U7207 ( .A1(n5718), .A2(n5717), .ZN(n8669) );
  NAND2_X1 U7208 ( .A1(n8669), .A2(n8016), .ZN(n5719) );
  NAND2_X1 U7209 ( .A1(n8134), .A2(n5719), .ZN(n8131) );
  INV_X1 U7210 ( .A(n5721), .ZN(n5722) );
  NAND2_X1 U7211 ( .A1(n5720), .A2(n5722), .ZN(n5723) );
  NAND2_X2 U7212 ( .A1(n8131), .A2(n5723), .ZN(n5750) );
  INV_X1 U7213 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n5727) );
  INV_X1 U7214 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7859) );
  MUX2_X1 U7215 ( .A(n5727), .B(n7859), .S(n7590), .Z(n5728) );
  INV_X1 U7216 ( .A(SI_23_), .ZN(n9961) );
  NAND2_X1 U7217 ( .A1(n5728), .A2(n9961), .ZN(n5757) );
  INV_X1 U7218 ( .A(n5728), .ZN(n5729) );
  NAND2_X1 U7219 ( .A1(n5729), .A2(SI_23_), .ZN(n5730) );
  NAND2_X1 U7220 ( .A1(n7858), .A2(n8189), .ZN(n5732) );
  NAND2_X1 U7221 ( .A1(n5387), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n5731) );
  XNOR2_X1 U7222 ( .A(n8760), .B(n8007), .ZN(n5751) );
  MUX2_X1 U7223 ( .A(n5734), .B(n5733), .S(n5749), .Z(n5747) );
  INV_X1 U7224 ( .A(n8760), .ZN(n8645) );
  NOR2_X1 U7225 ( .A1(n8645), .A2(n8167), .ZN(n5746) );
  INV_X1 U7226 ( .A(n8643), .ZN(n5735) );
  OAI22_X1 U7227 ( .A1(n10199), .A2(n5735), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10069), .ZN(n5745) );
  INV_X1 U7228 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n10144) );
  NAND2_X1 U7229 ( .A1(n5737), .A2(n10144), .ZN(n5738) );
  NAND2_X1 U7230 ( .A1(n5762), .A2(n5738), .ZN(n8625) );
  OR2_X1 U7231 ( .A1(n8625), .A2(n7625), .ZN(n5743) );
  INV_X1 U7232 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n8626) );
  NAND2_X1 U7233 ( .A1(n7669), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n5740) );
  NAND2_X1 U7234 ( .A1(n7670), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n5739) );
  OAI211_X1 U7235 ( .C1(n7673), .C2(n8626), .A(n5740), .B(n5739), .ZN(n5741)
         );
  INV_X1 U7236 ( .A(n5741), .ZN(n5742) );
  NAND2_X1 U7237 ( .A1(n5743), .A2(n5742), .ZN(n8410) );
  OAI22_X1 U7238 ( .A1(n8638), .A2(n8161), .B1(n8160), .B2(n8639), .ZN(n5744)
         );
  OR4_X1 U7239 ( .A1(n5747), .A2(n5746), .A3(n5745), .A4(n5744), .ZN(P2_U3218)
         );
  NOR2_X1 U7240 ( .A1(n8142), .A2(n8638), .ZN(n5761) );
  AND2_X1 U7241 ( .A1(n8410), .A2(n8016), .ZN(n7997) );
  NOR2_X1 U7242 ( .A1(n7997), .A2(n8156), .ZN(n5760) );
  NAND2_X1 U7243 ( .A1(n5749), .A2(n5748), .ZN(n5754) );
  INV_X1 U7244 ( .A(n5750), .ZN(n5752) );
  NAND2_X1 U7245 ( .A1(n5752), .A2(n5751), .ZN(n5753) );
  NAND2_X2 U7246 ( .A1(n5754), .A2(n5753), .ZN(n7999) );
  INV_X1 U7247 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7365) );
  INV_X1 U7248 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7877) );
  MUX2_X1 U7249 ( .A(n7365), .B(n7877), .S(n7590), .Z(n7451) );
  XNOR2_X1 U7250 ( .A(n7451), .B(SI_24_), .ZN(n7449) );
  XNOR2_X1 U7251 ( .A(n7448), .B(n7449), .ZN(n7876) );
  NAND2_X1 U7252 ( .A1(n7876), .A2(n8189), .ZN(n5759) );
  NAND2_X1 U7253 ( .A1(n5387), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n5758) );
  XNOR2_X1 U7254 ( .A(n8833), .B(n5263), .ZN(n8000) );
  MUX2_X1 U7255 ( .A(n5761), .B(n5760), .S(n7998), .Z(n5772) );
  NOR2_X1 U7256 ( .A1(n8628), .A2(n8167), .ZN(n5771) );
  OAI22_X1 U7257 ( .A1(n10199), .A2(n8625), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10144), .ZN(n5770) );
  INV_X1 U7258 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8104) );
  NAND2_X1 U7259 ( .A1(n5762), .A2(n8104), .ZN(n5763) );
  NAND2_X1 U7260 ( .A1(n7642), .A2(n5763), .ZN(n8603) );
  OR2_X1 U7261 ( .A1(n8603), .A2(n7625), .ZN(n5768) );
  INV_X1 U7262 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n8604) );
  NAND2_X1 U7263 ( .A1(n7670), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n5765) );
  NAND2_X1 U7264 ( .A1(n7669), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n5764) );
  OAI211_X1 U7265 ( .C1(n7673), .C2(n8604), .A(n5765), .B(n5764), .ZN(n5766)
         );
  INV_X1 U7266 ( .A(n5766), .ZN(n5767) );
  NAND2_X1 U7267 ( .A1(n5768), .A2(n5767), .ZN(n8618) );
  OAI22_X1 U7268 ( .A1(n8586), .A2(n8161), .B1(n8160), .B2(n8411), .ZN(n5769)
         );
  OR4_X1 U7269 ( .A1(n5772), .A2(n5771), .A3(n5770), .A4(n5769), .ZN(P2_U3231)
         );
  XNOR2_X1 U7270 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  NAND2_X1 U7271 ( .A1(n8185), .A2(P2_U3152), .ZN(n7595) );
  CLKBUF_X1 U7272 ( .A(n7595), .Z(n8872) );
  AOI22_X1 U7273 ( .A1(n8869), .A2(P1_DATAO_REG_1__SCAN_IN), .B1(n6005), .B2(
        P2_STATE_REG_SCAN_IN), .ZN(n5773) );
  OAI21_X1 U7274 ( .B1(n6305), .B2(n8872), .A(n5773), .ZN(P2_U3357) );
  INV_X1 U7275 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6306) );
  NOR2_X1 U7276 ( .A1(n8185), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9768) );
  INV_X1 U7277 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n10113) );
  OAI222_X1 U7278 ( .A1(n9774), .A2(n6306), .B1(n9773), .B2(n6305), .C1(n6309), 
        .C2(P1_U3084), .ZN(P1_U3352) );
  INV_X1 U7279 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6299) );
  INV_X1 U7280 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n6027) );
  OR2_X1 U7281 ( .A1(n5774), .A2(n6027), .ZN(n5776) );
  XNOR2_X1 U7282 ( .A(n5776), .B(n5775), .ZN(n6304) );
  OAI222_X1 U7283 ( .A1(n9774), .A2(n6299), .B1(n9773), .B2(n6301), .C1(n6304), 
        .C2(P1_U3084), .ZN(P1_U3351) );
  AOI22_X1 U7284 ( .A1(n8427), .A2(P2_STATE_REG_SCAN_IN), .B1(n8869), .B2(
        P1_DATAO_REG_3__SCAN_IN), .ZN(n5777) );
  OAI21_X1 U7285 ( .B1(n6398), .B2(n7595), .A(n5777), .ZN(P2_U3355) );
  INV_X1 U7286 ( .A(n8869), .ZN(n7510) );
  INV_X1 U7287 ( .A(n5855), .ZN(n5939) );
  OAI222_X1 U7288 ( .A1(n7510), .A2(n5185), .B1(n8872), .B2(n6301), .C1(
        P2_U3152), .C2(n5939), .ZN(P2_U3356) );
  INV_X1 U7289 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6397) );
  NAND2_X1 U7290 ( .A1(n5778), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5779) );
  XNOR2_X1 U7291 ( .A(n5779), .B(n5098), .ZN(n6401) );
  OAI222_X1 U7292 ( .A1(n9774), .A2(n6397), .B1(n9773), .B2(n6398), .C1(n6401), 
        .C2(P1_U3084), .ZN(P1_U3350) );
  INV_X1 U7293 ( .A(n5849), .ZN(n5877) );
  OAI222_X1 U7294 ( .A1(n7510), .A2(n4579), .B1(n8872), .B2(n6411), .C1(
        P2_U3152), .C2(n5877), .ZN(P2_U3354) );
  INV_X1 U7295 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6410) );
  NAND2_X1 U7296 ( .A1(n5780), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5781) );
  INV_X1 U7297 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n9983) );
  XNOR2_X1 U7298 ( .A(n5781), .B(n9983), .ZN(n6414) );
  OAI222_X1 U7299 ( .A1(n9774), .A2(n6410), .B1(n9773), .B2(n6411), .C1(n6414), 
        .C2(P1_U3084), .ZN(P1_U3349) );
  AND2_X1 U7300 ( .A1(n7246), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5782) );
  INV_X1 U7301 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n5789) );
  NAND2_X1 U7302 ( .A1(n7461), .A2(P1_B_REG_SCAN_IN), .ZN(n5783) );
  MUX2_X1 U7303 ( .A(P1_B_REG_SCAN_IN), .B(n5783), .S(n7364), .Z(n5785) );
  NAND2_X1 U7304 ( .A1(n9761), .A2(n5789), .ZN(n5787) );
  NAND2_X1 U7305 ( .A1(n7509), .A2(n7461), .ZN(n5786) );
  NAND2_X1 U7306 ( .A1(n5787), .A2(n5786), .ZN(n6367) );
  INV_X1 U7307 ( .A(n6367), .ZN(n6601) );
  NAND2_X1 U7308 ( .A1(n6601), .A2(n9762), .ZN(n5788) );
  OAI21_X1 U7309 ( .B1(n9762), .B2(n5789), .A(n5788), .ZN(P1_U3441) );
  INV_X1 U7310 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6460) );
  NOR2_X1 U7311 ( .A1(n5113), .A2(n6027), .ZN(n5790) );
  MUX2_X1 U7312 ( .A(n6027), .B(n5790), .S(P1_IR_REG_5__SCAN_IN), .Z(n5792) );
  AND2_X1 U7313 ( .A1(n5113), .A2(n5791), .ZN(n5793) );
  OAI222_X1 U7314 ( .A1(n9774), .A2(n6460), .B1(n9773), .B2(n6461), .C1(n6464), 
        .C2(P1_U3084), .ZN(P1_U3348) );
  INV_X1 U7315 ( .A(n5884), .ZN(n5867) );
  OAI222_X1 U7316 ( .A1(n7510), .A2(n4572), .B1(n8872), .B2(n6461), .C1(
        P2_U3152), .C2(n5867), .ZN(P2_U3353) );
  NOR2_X1 U7317 ( .A1(n5793), .A2(n6027), .ZN(n5794) );
  MUX2_X1 U7318 ( .A(n6027), .B(n5794), .S(P1_IR_REG_6__SCAN_IN), .Z(n5796) );
  INV_X1 U7319 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n9930) );
  OAI222_X1 U7320 ( .A1(n6586), .A2(P1_U3084), .B1(n9773), .B2(n6583), .C1(
        n9930), .C2(n9774), .ZN(P1_U3347) );
  INV_X1 U7321 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n5797) );
  INV_X1 U7322 ( .A(n5916), .ZN(n5923) );
  OAI222_X1 U7323 ( .A1(n7510), .A2(n5797), .B1(n8872), .B2(n6583), .C1(
        P2_U3152), .C2(n5923), .ZN(P2_U3352) );
  INV_X1 U7324 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n5798) );
  INV_X1 U7325 ( .A(n6716), .ZN(n5801) );
  INV_X1 U7326 ( .A(n6168), .ZN(n5929) );
  OAI222_X1 U7327 ( .A1(n7510), .A2(n5798), .B1(n8872), .B2(n5801), .C1(
        P2_U3152), .C2(n5929), .ZN(P2_U3351) );
  INV_X1 U7328 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6717) );
  NAND2_X1 U7329 ( .A1(n5795), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5800) );
  XNOR2_X1 U7330 ( .A(n5800), .B(n5799), .ZN(n6720) );
  OAI222_X1 U7331 ( .A1(n9774), .A2(n6717), .B1(n9773), .B2(n5801), .C1(n6720), 
        .C2(P1_U3084), .ZN(P1_U3346) );
  NAND2_X1 U7332 ( .A1(n5231), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n5805) );
  NAND2_X1 U7333 ( .A1(n7669), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n5804) );
  NAND2_X1 U7334 ( .A1(n7670), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n5803) );
  AND3_X1 U7335 ( .A1(n5805), .A2(n5804), .A3(n5803), .ZN(n8548) );
  NAND2_X1 U7336 ( .A1(n8412), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n5806) );
  OAI21_X1 U7337 ( .B1(n8412), .B2(n8548), .A(n5806), .ZN(P2_U3582) );
  INV_X1 U7338 ( .A(n6841), .ZN(n5812) );
  NAND2_X1 U7339 ( .A1(n5807), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5809) );
  OR2_X1 U7340 ( .A1(n5809), .A2(n5808), .ZN(n5810) );
  NAND2_X1 U7341 ( .A1(n5809), .A2(n5808), .ZN(n5820) );
  INV_X1 U7342 ( .A(n10300), .ZN(n5976) );
  OAI222_X1 U7343 ( .A1(n9774), .A2(n5811), .B1(n9773), .B2(n5812), .C1(n5976), 
        .C2(P1_U3084), .ZN(P1_U3345) );
  INV_X1 U7344 ( .A(n6348), .ZN(n6176) );
  OAI222_X1 U7345 ( .A1(n7510), .A2(n5813), .B1(n8872), .B2(n5812), .C1(
        P2_U3152), .C2(n6176), .ZN(P2_U3350) );
  NAND2_X1 U7346 ( .A1(n5814), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8405) );
  NAND2_X1 U7347 ( .A1(n10458), .A2(n8405), .ZN(n5816) );
  NAND2_X1 U7348 ( .A1(n5816), .A2(n5815), .ZN(n5819) );
  OR2_X1 U7349 ( .A1(n10458), .A2(n5817), .ZN(n5818) );
  NAND2_X1 U7350 ( .A1(n5819), .A2(n5818), .ZN(n10404) );
  NOR2_X1 U7351 ( .A1(n10404), .A2(P2_U3966), .ZN(P2_U3151) );
  NAND2_X1 U7352 ( .A1(n5820), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5821) );
  XNOR2_X1 U7353 ( .A(n5821), .B(P1_IR_REG_9__SCAN_IN), .ZN(n10309) );
  INV_X1 U7354 ( .A(n10309), .ZN(n5822) );
  INV_X1 U7355 ( .A(n6906), .ZN(n5823) );
  OAI222_X1 U7356 ( .A1(P1_U3084), .A2(n5822), .B1(n9773), .B2(n5823), .C1(
        n9902), .C2(n9774), .ZN(P1_U3344) );
  INV_X1 U7357 ( .A(n6650), .ZN(n6356) );
  OAI222_X1 U7358 ( .A1(n7510), .A2(n5824), .B1(n8872), .B2(n5823), .C1(n6356), 
        .C2(P2_U3152), .ZN(P2_U3349) );
  INV_X1 U7359 ( .A(n7001), .ZN(n5830) );
  NAND2_X1 U7360 ( .A1(n5827), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5825) );
  MUX2_X1 U7361 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5825), .S(
        P1_IR_REG_10__SCAN_IN), .Z(n5826) );
  INV_X1 U7362 ( .A(n5826), .ZN(n5828) );
  NOR2_X1 U7363 ( .A1(n5828), .A2(n6025), .ZN(n7002) );
  INV_X1 U7364 ( .A(n7002), .ZN(n5829) );
  OAI222_X1 U7365 ( .A1(n9774), .A2(n10063), .B1(n9773), .B2(n5830), .C1(
        P1_U3084), .C2(n5829), .ZN(P1_U3343) );
  INV_X1 U7366 ( .A(n7036), .ZN(n6658) );
  OAI222_X1 U7367 ( .A1(n7510), .A2(n5831), .B1(n8872), .B2(n5830), .C1(n6658), 
        .C2(P2_U3152), .ZN(P2_U3348) );
  OAI211_X1 U7368 ( .C1(n10458), .C2(n6035), .A(n8405), .B(n5832), .ZN(n5845)
         );
  NAND2_X1 U7369 ( .A1(n5845), .A2(n5843), .ZN(n5833) );
  NAND2_X1 U7370 ( .A1(n8412), .A2(n5833), .ZN(n5862) );
  NAND2_X1 U7371 ( .A1(n5862), .A2(n5602), .ZN(n10406) );
  INV_X1 U7372 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n10092) );
  NOR2_X1 U7373 ( .A1(n10092), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6223) );
  INV_X1 U7374 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n7700) );
  NAND2_X1 U7375 ( .A1(n10413), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6002) );
  INV_X1 U7376 ( .A(n6002), .ZN(n5834) );
  INV_X1 U7377 ( .A(n6001), .ZN(n5836) );
  NAND2_X1 U7378 ( .A1(n6005), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5835) );
  NAND2_X1 U7379 ( .A1(n5836), .A2(n5835), .ZN(n5935) );
  INV_X1 U7380 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n5837) );
  XNOR2_X1 U7381 ( .A(n5855), .B(n5837), .ZN(n5936) );
  NAND2_X1 U7382 ( .A1(n5935), .A2(n5936), .ZN(n5934) );
  NAND2_X1 U7383 ( .A1(n5855), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5838) );
  NAND2_X1 U7384 ( .A1(n5934), .A2(n5838), .ZN(n8434) );
  OR2_X1 U7385 ( .A1(n8427), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5840) );
  NAND2_X1 U7386 ( .A1(n8427), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5839) );
  AND2_X1 U7387 ( .A1(n5840), .A2(n5839), .ZN(n8435) );
  NAND2_X1 U7388 ( .A1(n5849), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5841) );
  OAI21_X1 U7389 ( .B1(n5849), .B2(P2_REG1_REG_4__SCAN_IN), .A(n5841), .ZN(
        n5869) );
  NAND2_X1 U7390 ( .A1(n5884), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5842) );
  OAI21_X1 U7391 ( .B1(n5884), .B2(P2_REG1_REG_5__SCAN_IN), .A(n5842), .ZN(
        n5846) );
  AND2_X1 U7392 ( .A1(n5843), .A2(n8401), .ZN(n5844) );
  NAND2_X1 U7393 ( .A1(n5845), .A2(n5844), .ZN(n10407) );
  AOI211_X1 U7394 ( .C1(n5847), .C2(n5846), .A(n5878), .B(n10407), .ZN(n5848)
         );
  AOI211_X1 U7395 ( .C1(P2_ADDR_REG_5__SCAN_IN), .C2(n10404), .A(n6223), .B(
        n5848), .ZN(n5866) );
  NAND2_X1 U7396 ( .A1(n5849), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5859) );
  INV_X1 U7397 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n5850) );
  MUX2_X1 U7398 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n5850), .S(n5849), .Z(n5873)
         );
  NAND2_X1 U7399 ( .A1(n8427), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5858) );
  INV_X1 U7400 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n5851) );
  MUX2_X1 U7401 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n5851), .S(n6005), .Z(n5852)
         );
  NAND3_X1 U7402 ( .A1(n5852), .A2(P2_REG2_REG_0__SCAN_IN), .A3(n10413), .ZN(
        n6007) );
  INV_X1 U7403 ( .A(n6007), .ZN(n5853) );
  AOI21_X1 U7404 ( .B1(n6005), .B2(P2_REG2_REG_1__SCAN_IN), .A(n5853), .ZN(
        n5933) );
  INV_X1 U7405 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n5854) );
  MUX2_X1 U7406 ( .A(n5854), .B(P2_REG2_REG_2__SCAN_IN), .S(n5855), .Z(n5932)
         );
  NOR2_X1 U7407 ( .A1(n5933), .A2(n5932), .ZN(n5931) );
  AOI21_X1 U7408 ( .B1(n5855), .B2(P2_REG2_REG_2__SCAN_IN), .A(n5931), .ZN(
        n8429) );
  INV_X1 U7409 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n5856) );
  MUX2_X1 U7410 ( .A(n5856), .B(P2_REG2_REG_3__SCAN_IN), .S(n8427), .Z(n8430)
         );
  OR2_X1 U7411 ( .A1(n8429), .A2(n8430), .ZN(n5857) );
  NAND2_X1 U7412 ( .A1(n5858), .A2(n5857), .ZN(n5874) );
  NAND2_X1 U7413 ( .A1(n5873), .A2(n5874), .ZN(n5872) );
  NAND2_X1 U7414 ( .A1(n5859), .A2(n5872), .ZN(n5864) );
  INV_X1 U7415 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n5860) );
  MUX2_X1 U7416 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n5860), .S(n5884), .Z(n5863)
         );
  NOR2_X1 U7417 ( .A1(n5602), .A2(n8401), .ZN(n5861) );
  NAND2_X1 U7418 ( .A1(n5863), .A2(n5864), .ZN(n5885) );
  OAI211_X1 U7419 ( .C1(n5864), .C2(n5863), .A(n10403), .B(n5885), .ZN(n5865)
         );
  OAI211_X1 U7420 ( .C1(n10406), .C2(n5867), .A(n5866), .B(n5865), .ZN(
        P2_U3250) );
  NOR2_X1 U7421 ( .A1(n5222), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6213) );
  AOI211_X1 U7422 ( .C1(n5870), .C2(n5869), .A(n5868), .B(n10407), .ZN(n5871)
         );
  AOI211_X1 U7423 ( .C1(P2_ADDR_REG_4__SCAN_IN), .C2(n10404), .A(n6213), .B(
        n5871), .ZN(n5876) );
  OAI211_X1 U7424 ( .C1(n5874), .C2(n5873), .A(n10403), .B(n5872), .ZN(n5875)
         );
  OAI211_X1 U7425 ( .C1(n10406), .C2(n5877), .A(n5876), .B(n5875), .ZN(
        P2_U3249) );
  NAND2_X1 U7426 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3152), .ZN(n7605) );
  INV_X1 U7427 ( .A(n7605), .ZN(n5883) );
  AOI21_X1 U7428 ( .B1(n5884), .B2(P2_REG1_REG_5__SCAN_IN), .A(n5878), .ZN(
        n5881) );
  INV_X1 U7429 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n5879) );
  MUX2_X1 U7430 ( .A(n5879), .B(P2_REG1_REG_6__SCAN_IN), .S(n5916), .Z(n5880)
         );
  AOI211_X1 U7431 ( .C1(n5881), .C2(n5880), .A(n5915), .B(n10407), .ZN(n5882)
         );
  AOI211_X1 U7432 ( .C1(P2_ADDR_REG_6__SCAN_IN), .C2(n10404), .A(n5883), .B(
        n5882), .ZN(n5891) );
  NAND2_X1 U7433 ( .A1(n5884), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5886) );
  NAND2_X1 U7434 ( .A1(n5886), .A2(n5885), .ZN(n5889) );
  INV_X1 U7435 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n5887) );
  MUX2_X1 U7436 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n5887), .S(n5916), .Z(n5888)
         );
  NAND2_X1 U7437 ( .A1(n5888), .A2(n5889), .ZN(n5922) );
  OAI211_X1 U7438 ( .C1(n5889), .C2(n5888), .A(n10403), .B(n5922), .ZN(n5890)
         );
  OAI211_X1 U7439 ( .C1(n10406), .C2(n5923), .A(n5891), .B(n5890), .ZN(
        P2_U3251) );
  INV_X1 U7440 ( .A(n10337), .ZN(n10299) );
  INV_X1 U7441 ( .A(n5943), .ZN(n5903) );
  NOR2_X1 U7442 ( .A1(n5942), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5894) );
  NOR2_X1 U7443 ( .A1(n5894), .A2(n8071), .ZN(n6156) );
  INV_X1 U7444 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n5895) );
  XNOR2_X1 U7445 ( .A(n6156), .B(n5895), .ZN(n5897) );
  INV_X1 U7446 ( .A(n5942), .ZN(n9405) );
  OR2_X1 U7447 ( .A1(n8071), .A2(n9405), .ZN(n5898) );
  INV_X1 U7448 ( .A(n5898), .ZN(n6158) );
  INV_X1 U7449 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n6273) );
  NAND2_X1 U7450 ( .A1(n6158), .A2(n6273), .ZN(n5896) );
  NAND4_X1 U7451 ( .A1(n5897), .A2(P1_STATE_REG_SCAN_IN), .A3(n6842), .A4(
        n5896), .ZN(n5902) );
  NOR2_X1 U7452 ( .A1(n5898), .A2(P1_U3084), .ZN(n5899) );
  NAND3_X1 U7453 ( .A1(n10332), .A2(P1_IR_REG_0__SCAN_IN), .A3(n6273), .ZN(
        n5901) );
  NAND2_X1 U7454 ( .A1(P1_U3084), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5900) );
  OAI211_X1 U7455 ( .C1(n5903), .C2(n5902), .A(n5901), .B(n5900), .ZN(n5904)
         );
  AOI21_X1 U7456 ( .B1(n10299), .B2(P1_ADDR_REG_0__SCAN_IN), .A(n5904), .ZN(
        n5905) );
  INV_X1 U7457 ( .A(n5905), .ZN(P1_U3241) );
  INV_X1 U7458 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n5910) );
  NAND2_X1 U7459 ( .A1(n7669), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n5908) );
  NAND2_X1 U7460 ( .A1(n5231), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n5907) );
  NAND2_X1 U7461 ( .A1(n7670), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n5906) );
  NAND3_X1 U7462 ( .A1(n5908), .A2(n5907), .A3(n5906), .ZN(n8526) );
  NAND2_X1 U7463 ( .A1(P2_U3966), .A2(n8526), .ZN(n5909) );
  OAI21_X1 U7464 ( .B1(P2_U3966), .B2(n5910), .A(n5909), .ZN(P2_U3583) );
  OR2_X1 U7465 ( .A1(n6025), .A2(n6027), .ZN(n5911) );
  XNOR2_X1 U7466 ( .A(n5911), .B(P1_IR_REG_11__SCAN_IN), .ZN(n10323) );
  INV_X1 U7467 ( .A(n10323), .ZN(n6244) );
  INV_X1 U7468 ( .A(n7184), .ZN(n5914) );
  INV_X1 U7469 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n5912) );
  OAI222_X1 U7470 ( .A1(P1_U3084), .A2(n6244), .B1(n9773), .B2(n5914), .C1(
        n5912), .C2(n9774), .ZN(P1_U3342) );
  INV_X1 U7471 ( .A(n7217), .ZN(n7211) );
  INV_X1 U7472 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n5913) );
  OAI222_X1 U7473 ( .A1(P2_U3152), .A2(n7211), .B1(n8872), .B2(n5914), .C1(
        n5913), .C2(n7510), .ZN(P2_U3347) );
  NOR2_X1 U7474 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9929), .ZN(n5921) );
  NAND2_X1 U7475 ( .A1(n6168), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5917) );
  OAI21_X1 U7476 ( .B1(n6168), .B2(P2_REG1_REG_7__SCAN_IN), .A(n5917), .ZN(
        n5918) );
  AOI211_X1 U7477 ( .C1(n5919), .C2(n5918), .A(n6163), .B(n10407), .ZN(n5920)
         );
  AOI211_X1 U7478 ( .C1(P2_ADDR_REG_7__SCAN_IN), .C2(n10404), .A(n5921), .B(
        n5920), .ZN(n5928) );
  OAI21_X1 U7479 ( .B1(n5923), .B2(n5887), .A(n5922), .ZN(n5926) );
  MUX2_X1 U7480 ( .A(n6820), .B(P2_REG2_REG_7__SCAN_IN), .S(n6168), .Z(n5924)
         );
  INV_X1 U7481 ( .A(n5924), .ZN(n5925) );
  NAND2_X1 U7482 ( .A1(n5925), .A2(n5926), .ZN(n6169) );
  OAI211_X1 U7483 ( .C1(n5926), .C2(n5925), .A(n10403), .B(n6169), .ZN(n5927)
         );
  OAI211_X1 U7484 ( .C1(n10406), .C2(n5929), .A(n5928), .B(n5927), .ZN(
        P2_U3252) );
  INV_X1 U7485 ( .A(n7282), .ZN(n5970) );
  AOI22_X1 U7486 ( .A1(n8440), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_12__SCAN_IN), .B2(n8869), .ZN(n5930) );
  OAI21_X1 U7487 ( .B1(n5970), .B2(n8872), .A(n5930), .ZN(P2_U3346) );
  INV_X1 U7488 ( .A(n10403), .ZN(n10405) );
  AOI211_X1 U7489 ( .C1(n5933), .C2(n5932), .A(n5931), .B(n10405), .ZN(n5941)
         );
  AOI22_X1 U7490 ( .A1(n10404), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n5938) );
  INV_X1 U7491 ( .A(n10407), .ZN(n10402) );
  OAI211_X1 U7492 ( .C1(n5936), .C2(n5935), .A(n10402), .B(n5934), .ZN(n5937)
         );
  OAI211_X1 U7493 ( .C1(n10406), .C2(n5939), .A(n5938), .B(n5937), .ZN(n5940)
         );
  OR2_X1 U7494 ( .A1(n5941), .A2(n5940), .ZN(P2_U3247) );
  NOR2_X1 U7495 ( .A1(n5942), .A2(P1_U3084), .ZN(n7534) );
  NAND2_X1 U7496 ( .A1(n5943), .A2(n7534), .ZN(n9399) );
  INV_X1 U7497 ( .A(n9399), .ZN(n5951) );
  INV_X1 U7498 ( .A(n8071), .ZN(n9335) );
  INV_X1 U7499 ( .A(n10331), .ZN(n9385) );
  INV_X1 U7500 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n5944) );
  AND2_X1 U7501 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n6154) );
  INV_X1 U7502 ( .A(n6309), .ZN(n5945) );
  NAND2_X1 U7503 ( .A1(n5945), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5946) );
  NAND2_X1 U7504 ( .A1(n6063), .A2(n5946), .ZN(n6105) );
  XNOR2_X1 U7505 ( .A(n6304), .B(P1_REG2_REG_2__SCAN_IN), .ZN(n6106) );
  INV_X1 U7506 ( .A(n6304), .ZN(n6107) );
  NAND2_X1 U7507 ( .A1(n6107), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5947) );
  XNOR2_X1 U7508 ( .A(n6401), .B(P1_REG2_REG_3__SCAN_IN), .ZN(n6081) );
  INV_X1 U7509 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n5948) );
  INV_X1 U7510 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n5949) );
  XNOR2_X1 U7511 ( .A(n6414), .B(n5949), .ZN(n6192) );
  NOR2_X1 U7512 ( .A1(n6191), .A2(n6192), .ZN(n6190) );
  AND2_X1 U7513 ( .A1(n6414), .A2(n5949), .ZN(n5950) );
  NOR2_X1 U7514 ( .A1(n6190), .A2(n5950), .ZN(n5985) );
  XNOR2_X1 U7515 ( .A(n6464), .B(P1_REG2_REG_5__SCAN_IN), .ZN(n5983) );
  XNOR2_X1 U7516 ( .A(n5985), .B(n5983), .ZN(n5966) );
  INV_X1 U7517 ( .A(n6464), .ZN(n5974) );
  AND2_X1 U7518 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n8949) );
  INV_X1 U7519 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n5952) );
  MUX2_X1 U7520 ( .A(n5952), .B(P1_REG1_REG_1__SCAN_IN), .S(n6309), .Z(n6066)
         );
  AND2_X1 U7521 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n6067) );
  NAND2_X1 U7522 ( .A1(n6066), .A2(n6067), .ZN(n6109) );
  OR2_X1 U7523 ( .A1(n6309), .A2(n5952), .ZN(n6108) );
  NAND2_X1 U7524 ( .A1(n6109), .A2(n6108), .ZN(n5955) );
  INV_X1 U7525 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n5953) );
  MUX2_X1 U7526 ( .A(n5953), .B(P1_REG1_REG_2__SCAN_IN), .S(n6304), .Z(n5954)
         );
  NAND2_X1 U7527 ( .A1(n5955), .A2(n5954), .ZN(n6112) );
  NAND2_X1 U7528 ( .A1(n6107), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6074) );
  NAND2_X1 U7529 ( .A1(n6112), .A2(n6074), .ZN(n5957) );
  INV_X1 U7530 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n5958) );
  MUX2_X1 U7531 ( .A(n5958), .B(P1_REG1_REG_3__SCAN_IN), .S(n6401), .Z(n5956)
         );
  NAND2_X1 U7532 ( .A1(n5957), .A2(n5956), .ZN(n6076) );
  OR2_X1 U7533 ( .A1(n6401), .A2(n5958), .ZN(n5959) );
  AND2_X1 U7534 ( .A1(n6076), .A2(n5959), .ZN(n6195) );
  INV_X1 U7535 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6439) );
  MUX2_X1 U7536 ( .A(n6439), .B(P1_REG1_REG_4__SCAN_IN), .S(n6414), .Z(n6194)
         );
  NAND2_X1 U7537 ( .A1(n6195), .A2(n6194), .ZN(n6193) );
  NAND2_X1 U7538 ( .A1(n6414), .A2(n6439), .ZN(n5960) );
  NAND2_X1 U7539 ( .A1(n6193), .A2(n5960), .ZN(n5962) );
  INV_X1 U7540 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6481) );
  MUX2_X1 U7541 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n6481), .S(n6464), .Z(n5961)
         );
  NOR2_X1 U7542 ( .A1(n5962), .A2(n5961), .ZN(n5973) );
  INV_X1 U7543 ( .A(n10332), .ZN(n9367) );
  AOI211_X1 U7544 ( .C1(n5962), .C2(n5961), .A(n5973), .B(n9367), .ZN(n5963)
         );
  AOI211_X1 U7545 ( .C1(n10324), .C2(n5974), .A(n8949), .B(n5963), .ZN(n5965)
         );
  NAND2_X1 U7546 ( .A1(n10299), .A2(P1_ADDR_REG_5__SCAN_IN), .ZN(n5964) );
  OAI211_X1 U7547 ( .C1(n9385), .C2(n5966), .A(n5965), .B(n5964), .ZN(P1_U3246) );
  NAND2_X1 U7548 ( .A1(n6025), .A2(n6023), .ZN(n5967) );
  NAND2_X1 U7549 ( .A1(n5967), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5968) );
  NAND2_X1 U7550 ( .A1(n5968), .A2(n6022), .ZN(n6058) );
  OR2_X1 U7551 ( .A1(n5968), .A2(n6022), .ZN(n5969) );
  INV_X1 U7552 ( .A(n7283), .ZN(n6242) );
  OAI222_X1 U7553 ( .A1(n9774), .A2(n9876), .B1(n9773), .B2(n5970), .C1(n6242), 
        .C2(P1_U3084), .ZN(P1_U3341) );
  NOR2_X1 U7554 ( .A1(n10309), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5971) );
  AOI21_X1 U7555 ( .B1(P1_REG1_REG_9__SCAN_IN), .B2(n10309), .A(n5971), .ZN(
        n10317) );
  INV_X1 U7556 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n5972) );
  NOR2_X1 U7557 ( .A1(n5976), .A2(n5972), .ZN(n5977) );
  INV_X1 U7558 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n5975) );
  INV_X1 U7559 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6835) );
  AOI21_X1 U7560 ( .B1(P1_REG1_REG_5__SCAN_IN), .B2(n5974), .A(n5973), .ZN(
        n6088) );
  MUX2_X1 U7561 ( .A(n6835), .B(P1_REG1_REG_6__SCAN_IN), .S(n6586), .Z(n6087)
         );
  AND2_X1 U7562 ( .A1(n6088), .A2(n6087), .ZN(n6085) );
  AOI21_X1 U7563 ( .B1(n6586), .B2(n6835), .A(n6085), .ZN(n6014) );
  MUX2_X1 U7564 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n5975), .S(n6720), .Z(n6015)
         );
  NOR2_X1 U7565 ( .A1(n6014), .A2(n6015), .ZN(n6013) );
  AOI21_X1 U7566 ( .B1(n6720), .B2(n5975), .A(n6013), .ZN(n10303) );
  NAND2_X1 U7567 ( .A1(n5976), .A2(n5972), .ZN(n10302) );
  OAI21_X1 U7568 ( .B1(n5977), .B2(n10303), .A(n10302), .ZN(n10318) );
  NAND2_X1 U7569 ( .A1(n10317), .A2(n10318), .ZN(n10316) );
  OAI21_X1 U7570 ( .B1(n10309), .B2(P1_REG1_REG_9__SCAN_IN), .A(n10316), .ZN(
        n5980) );
  INV_X1 U7571 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n5978) );
  MUX2_X1 U7572 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n5978), .S(n7002), .Z(n5979)
         );
  NAND2_X1 U7573 ( .A1(n5980), .A2(n5979), .ZN(n6236) );
  OAI21_X1 U7574 ( .B1(n5980), .B2(n5979), .A(n6236), .ZN(n5999) );
  INV_X1 U7575 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n5997) );
  NOR2_X1 U7576 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6934), .ZN(n7023) );
  AOI21_X1 U7577 ( .B1(n10324), .B2(n7002), .A(n7023), .ZN(n5996) );
  INV_X1 U7578 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n5981) );
  XNOR2_X1 U7579 ( .A(n7002), .B(n5981), .ZN(n5994) );
  NAND2_X1 U7580 ( .A1(n10309), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5992) );
  NOR2_X1 U7581 ( .A1(n10300), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5982) );
  AOI21_X1 U7582 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n10300), .A(n5982), .ZN(
        n10296) );
  XOR2_X1 U7583 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n6720), .Z(n6012) );
  INV_X1 U7584 ( .A(n6586), .ZN(n5989) );
  INV_X1 U7585 ( .A(n5983), .ZN(n5984) );
  INV_X1 U7586 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n5986) );
  NAND2_X1 U7587 ( .A1(n6464), .A2(n5986), .ZN(n5987) );
  INV_X1 U7588 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n5988) );
  MUX2_X1 U7589 ( .A(n5988), .B(P1_REG2_REG_6__SCAN_IN), .S(n6586), .Z(n6094)
         );
  INV_X1 U7590 ( .A(n6720), .ZN(n6016) );
  OAI22_X1 U7591 ( .A1(n6012), .A2(n4500), .B1(P1_REG2_REG_7__SCAN_IN), .B2(
        n6016), .ZN(n10297) );
  NAND2_X1 U7592 ( .A1(n10296), .A2(n10297), .ZN(n10295) );
  OAI21_X1 U7593 ( .B1(n10300), .B2(P1_REG2_REG_8__SCAN_IN), .A(n10295), .ZN(
        n10311) );
  OR2_X1 U7594 ( .A1(n10309), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5990) );
  NAND2_X1 U7595 ( .A1(n5990), .A2(n5992), .ZN(n10312) );
  NOR2_X1 U7596 ( .A1(n10311), .A2(n10312), .ZN(n10310) );
  INV_X1 U7597 ( .A(n10310), .ZN(n5991) );
  OAI211_X1 U7598 ( .C1(n5994), .C2(n5993), .A(n10331), .B(n4562), .ZN(n5995)
         );
  OAI211_X1 U7599 ( .C1(n5997), .C2(n10337), .A(n5996), .B(n5995), .ZN(n5998)
         );
  AOI21_X1 U7600 ( .B1(n5999), .B2(n10332), .A(n5998), .ZN(n6000) );
  INV_X1 U7601 ( .A(n6000), .ZN(P1_U3251) );
  INV_X1 U7602 ( .A(n10406), .ZN(n8491) );
  INV_X1 U7603 ( .A(n10404), .ZN(n7359) );
  INV_X1 U7604 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10511) );
  INV_X1 U7605 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n7685) );
  OAI22_X1 U7606 ( .A1(n7359), .A2(n10511), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7685), .ZN(n6004) );
  AOI211_X1 U7607 ( .C1(n6002), .C2(n4567), .A(n6001), .B(n10407), .ZN(n6003)
         );
  AOI211_X1 U7608 ( .C1(n8491), .C2(n6005), .A(n6004), .B(n6003), .ZN(n6011)
         );
  AND2_X1 U7609 ( .A1(n10413), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6009) );
  MUX2_X1 U7610 ( .A(n5851), .B(P2_REG2_REG_1__SCAN_IN), .S(n6005), .Z(n6006)
         );
  INV_X1 U7611 ( .A(n6006), .ZN(n6008) );
  OAI211_X1 U7612 ( .C1(n6009), .C2(n6008), .A(n10403), .B(n6007), .ZN(n6010)
         );
  NAND2_X1 U7613 ( .A1(n6011), .A2(n6010), .ZN(P2_U3246) );
  INV_X1 U7614 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n9793) );
  XNOR2_X1 U7615 ( .A(n6012), .B(n4500), .ZN(n6020) );
  AOI21_X1 U7616 ( .B1(n6015), .B2(n6014), .A(n6013), .ZN(n6018) );
  NAND2_X1 U7617 ( .A1(n10324), .A2(n6016), .ZN(n6017) );
  NAND2_X1 U7618 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n6754) );
  OAI211_X1 U7619 ( .C1(n6018), .C2(n9367), .A(n6017), .B(n6754), .ZN(n6019)
         );
  AOI21_X1 U7620 ( .B1(n10331), .B2(n6020), .A(n6019), .ZN(n6021) );
  OAI21_X1 U7621 ( .B1(n9793), .B2(n10337), .A(n6021), .ZN(P1_U3248) );
  INV_X1 U7622 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10121) );
  INV_X1 U7623 ( .A(n7410), .ZN(n6031) );
  INV_X1 U7624 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n10123) );
  AND3_X1 U7625 ( .A1(n6023), .A2(n6022), .A3(n10123), .ZN(n6024) );
  AND2_X1 U7626 ( .A1(n6025), .A2(n6024), .ZN(n6028) );
  NOR2_X1 U7627 ( .A1(n6028), .A2(n6027), .ZN(n6026) );
  MUX2_X1 U7628 ( .A(n6027), .B(n6026), .S(P1_IR_REG_14__SCAN_IN), .Z(n6030)
         );
  NAND2_X1 U7629 ( .A1(n6028), .A2(n10097), .ZN(n6252) );
  INV_X1 U7630 ( .A(n6252), .ZN(n6029) );
  NOR2_X1 U7631 ( .A1(n6030), .A2(n6029), .ZN(n7411) );
  INV_X1 U7632 ( .A(n7411), .ZN(n7249) );
  OAI222_X1 U7633 ( .A1(n9774), .A2(n10121), .B1(n9773), .B2(n6031), .C1(
        P1_U3084), .C2(n7249), .ZN(P1_U3339) );
  INV_X1 U7634 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6032) );
  INV_X1 U7635 ( .A(n7555), .ZN(n7560) );
  OAI222_X1 U7636 ( .A1(n7510), .A2(n6032), .B1(n8872), .B2(n6031), .C1(n7560), 
        .C2(P2_U3152), .ZN(P2_U3344) );
  INV_X1 U7637 ( .A(n6767), .ZN(n6207) );
  AND4_X1 U7638 ( .A1(n6098), .A2(P2_STATE_REG_SCAN_IN), .A3(n6207), .A4(n6769), .ZN(n6033) );
  AND2_X1 U7639 ( .A1(n6204), .A2(n6033), .ZN(n6034) );
  AND2_X2 U7640 ( .A1(n6206), .A2(n6034), .ZN(n10499) );
  MUX2_X1 U7641 ( .A(n4486), .B(n6035), .S(n5213), .Z(n6036) );
  INV_X1 U7642 ( .A(n6036), .ZN(n6039) );
  INV_X1 U7643 ( .A(n6037), .ZN(n6038) );
  NAND2_X1 U7644 ( .A1(n6039), .A2(n6038), .ZN(n10435) );
  NOR2_X1 U7645 ( .A1(n8398), .A2(n8517), .ZN(n6040) );
  NAND2_X1 U7646 ( .A1(n4486), .A2(n6040), .ZN(n6872) );
  NAND2_X1 U7647 ( .A1(n6041), .A2(n6042), .ZN(n8256) );
  NAND2_X1 U7648 ( .A1(n7112), .A2(n6043), .ZN(n7124) );
  NAND2_X1 U7649 ( .A1(n6041), .A2(n7702), .ZN(n6044) );
  OR2_X2 U7650 ( .A1(n6179), .A2(n8063), .ZN(n8254) );
  NAND2_X1 U7651 ( .A1(n6179), .A2(n8063), .ZN(n8257) );
  NAND2_X1 U7652 ( .A1(n6045), .A2(n6049), .ZN(n6281) );
  OAI21_X1 U7653 ( .B1(n6045), .B2(n6049), .A(n6281), .ZN(n6046) );
  INV_X1 U7654 ( .A(n6046), .ZN(n6782) );
  OR2_X1 U7655 ( .A1(n4486), .A2(n8517), .ZN(n8399) );
  INV_X1 U7656 ( .A(n6049), .ZN(n6050) );
  OAI21_X1 U7657 ( .B1(n6051), .B2(n6050), .A(n6284), .ZN(n6052) );
  AOI222_X1 U7658 ( .A1(n10432), .A2(n6052), .B1(n8425), .B2(n8701), .C1(n8426), .C2(n10216), .ZN(n6779) );
  NOR2_X1 U7659 ( .A1(n6042), .A2(n7120), .ZN(n6054) );
  INV_X1 U7660 ( .A(n6790), .ZN(n6053) );
  OAI21_X1 U7661 ( .B1(n8063), .B2(n6054), .A(n6053), .ZN(n6776) );
  INV_X1 U7662 ( .A(n6776), .ZN(n6055) );
  INV_X1 U7663 ( .A(n10472), .ZN(n10418) );
  INV_X1 U7664 ( .A(n8063), .ZN(n6778) );
  AOI22_X1 U7665 ( .A1(n6055), .A2(n10418), .B1(n8803), .B2(n6778), .ZN(n6056)
         );
  OAI211_X1 U7666 ( .C1(n10466), .C2(n6782), .A(n6779), .B(n6056), .ZN(n6209)
         );
  NAND2_X1 U7667 ( .A1(n6209), .A2(n10499), .ZN(n6057) );
  OAI21_X1 U7668 ( .B1(n10499), .B2(n5837), .A(n6057), .ZN(P2_U3522) );
  INV_X1 U7669 ( .A(n7372), .ZN(n6061) );
  NAND2_X1 U7670 ( .A1(n6058), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6059) );
  XNOR2_X1 U7671 ( .A(n6059), .B(P1_IR_REG_13__SCAN_IN), .ZN(n7373) );
  INV_X1 U7672 ( .A(n7373), .ZN(n6060) );
  OAI222_X1 U7673 ( .A1(n9774), .A2(n9943), .B1(n9773), .B2(n6061), .C1(
        P1_U3084), .C2(n6060), .ZN(P1_U3340) );
  INV_X1 U7674 ( .A(n7353), .ZN(n7215) );
  OAI222_X1 U7675 ( .A1(n7510), .A2(n6062), .B1(n8872), .B2(n6061), .C1(n7215), 
        .C2(P2_U3152), .ZN(P2_U3345) );
  INV_X1 U7676 ( .A(n10324), .ZN(n7444) );
  OAI211_X1 U7677 ( .C1(n6064), .C2(n6154), .A(n10331), .B(n6063), .ZN(n6065)
         );
  OAI21_X1 U7678 ( .B1(n7444), .B2(n6309), .A(n6065), .ZN(n6071) );
  INV_X1 U7679 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n6069) );
  OAI211_X1 U7680 ( .C1(n6067), .C2(n6066), .A(n10332), .B(n6109), .ZN(n6068)
         );
  OAI21_X1 U7681 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n6069), .A(n6068), .ZN(n6070) );
  AOI211_X1 U7682 ( .C1(n10299), .C2(P1_ADDR_REG_1__SCAN_IN), .A(n6071), .B(
        n6070), .ZN(n6072) );
  INV_X1 U7683 ( .A(n6072), .ZN(P1_U3242) );
  INV_X1 U7684 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n6084) );
  NAND2_X1 U7685 ( .A1(P1_U3084), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n6805) );
  MUX2_X1 U7686 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n5958), .S(n6401), .Z(n6073)
         );
  NAND3_X1 U7687 ( .A1(n6112), .A2(n6074), .A3(n6073), .ZN(n6075) );
  NAND3_X1 U7688 ( .A1(n10332), .A2(n6076), .A3(n6075), .ZN(n6077) );
  OAI211_X1 U7689 ( .C1(n7444), .C2(n6401), .A(n6805), .B(n6077), .ZN(n6078)
         );
  INV_X1 U7690 ( .A(n6078), .ZN(n6083) );
  OAI211_X1 U7691 ( .C1(n6081), .C2(n6080), .A(n10331), .B(n6079), .ZN(n6082)
         );
  OAI211_X1 U7692 ( .C1(n6084), .C2(n10337), .A(n6083), .B(n6082), .ZN(
        P1_U3244) );
  INV_X1 U7693 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n6097) );
  INV_X1 U7694 ( .A(n6085), .ZN(n6086) );
  OAI21_X1 U7695 ( .B1(n6088), .B2(n6087), .A(n6086), .ZN(n6090) );
  INV_X1 U7696 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6466) );
  NOR2_X1 U7697 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6466), .ZN(n6617) );
  NOR2_X1 U7698 ( .A1(n7444), .A2(n6586), .ZN(n6089) );
  AOI211_X1 U7699 ( .C1(n10332), .C2(n6090), .A(n6617), .B(n6089), .ZN(n6096)
         );
  INV_X1 U7700 ( .A(n6091), .ZN(n6092) );
  OAI211_X1 U7701 ( .C1(n6094), .C2(n6093), .A(n10331), .B(n6092), .ZN(n6095)
         );
  OAI211_X1 U7702 ( .C1(n6097), .C2(n10337), .A(n6096), .B(n6095), .ZN(
        P1_U3247) );
  INV_X1 U7703 ( .A(n8142), .ZN(n8057) );
  INV_X1 U7704 ( .A(n8156), .ZN(n10194) );
  AOI22_X1 U7705 ( .A1(n8057), .A2(n6047), .B1(n7120), .B2(n10194), .ZN(n6103)
         );
  INV_X1 U7706 ( .A(n8161), .ZN(n7611) );
  AND2_X1 U7707 ( .A1(n6098), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6203) );
  AND2_X1 U7708 ( .A1(n6099), .A2(n6203), .ZN(n8062) );
  INV_X1 U7709 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n10148) );
  OAI22_X1 U7710 ( .A1(n8167), .A2(n10465), .B1(n8062), .B2(n10148), .ZN(n6100) );
  AOI21_X1 U7711 ( .B1(n7611), .B2(n8426), .A(n6100), .ZN(n6101) );
  OAI21_X1 U7712 ( .B1(n6103), .B2(n6102), .A(n6101), .ZN(P2_U3234) );
  OAI211_X1 U7713 ( .C1(n6106), .C2(n6105), .A(n10331), .B(n6104), .ZN(n6116)
         );
  NAND2_X1 U7714 ( .A1(n10324), .A2(n6107), .ZN(n6115) );
  NAND2_X1 U7715 ( .A1(P1_U3084), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n6114) );
  MUX2_X1 U7716 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n5953), .S(n6304), .Z(n6110)
         );
  NAND3_X1 U7717 ( .A1(n6110), .A2(n6109), .A3(n6108), .ZN(n6111) );
  NAND3_X1 U7718 ( .A1(n10332), .A2(n6112), .A3(n6111), .ZN(n6113) );
  NAND4_X1 U7719 ( .A1(n6116), .A2(n6115), .A3(n6114), .A4(n6113), .ZN(n6160)
         );
  NAND2_X1 U7720 ( .A1(n4525), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6120) );
  MUX2_X1 U7721 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6120), .S(
        P1_IR_REG_19__SCAN_IN), .Z(n6122) );
  AND2_X1 U7722 ( .A1(n6945), .A2(n9544), .ZN(n6335) );
  NAND2_X1 U7723 ( .A1(n9263), .A2(n6335), .ZN(n6123) );
  NAND2_X2 U7724 ( .A1(n7750), .A2(n6123), .ZN(n6553) );
  AND2_X1 U7725 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), .ZN(
        n6125) );
  INV_X1 U7726 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n6128) );
  AND3_X1 U7727 ( .A1(n6128), .A2(n6127), .A3(n6124), .ZN(n6129) );
  NAND2_X1 U7728 ( .A1(n7984), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n6142) );
  NAND2_X1 U7729 ( .A1(n4827), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6141) );
  INV_X1 U7730 ( .A(n6137), .ZN(n7596) );
  NAND2_X1 U7731 ( .A1(n6404), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6140) );
  NAND2_X1 U7732 ( .A1(n7421), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n6139) );
  XNOR2_X1 U7733 ( .A(n6143), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n9775) );
  MUX2_X1 U7734 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9775), .S(n6300), .Z(n7599) );
  INV_X1 U7735 ( .A(n6380), .ZN(n6144) );
  AND2_X2 U7736 ( .A1(n6144), .A2(n6618), .ZN(n7890) );
  NAND2_X1 U7737 ( .A1(n7599), .A2(n7890), .ZN(n6146) );
  INV_X1 U7738 ( .A(n6618), .ZN(n6148) );
  NAND2_X1 U7739 ( .A1(n6148), .A2(P1_IR_REG_0__SCAN_IN), .ZN(n6145) );
  NAND2_X1 U7740 ( .A1(n9359), .A2(n7890), .ZN(n6152) );
  INV_X1 U7741 ( .A(n7599), .ZN(n6333) );
  NAND2_X1 U7742 ( .A1(n6148), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6149) );
  OAI21_X1 U7743 ( .B1(n6333), .B2(n7891), .A(n6149), .ZN(n6150) );
  INV_X1 U7744 ( .A(n6150), .ZN(n6151) );
  OAI21_X1 U7745 ( .B1(n6153), .B2(n6538), .A(n6540), .ZN(n7600) );
  INV_X1 U7746 ( .A(n7600), .ZN(n6159) );
  NAND3_X1 U7747 ( .A1(n9335), .A2(n9405), .A3(n6154), .ZN(n6155) );
  OAI211_X1 U7748 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n6156), .A(P1_U4006), .B(
        n6155), .ZN(n6157) );
  AOI21_X1 U7749 ( .B1(n6159), .B2(n6158), .A(n6157), .ZN(n6201) );
  AOI211_X1 U7750 ( .C1(n10299), .C2(P1_ADDR_REG_2__SCAN_IN), .A(n6160), .B(
        n6201), .ZN(n6161) );
  INV_X1 U7751 ( .A(n6161), .ZN(P1_U3243) );
  INV_X1 U7752 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n6162) );
  NOR2_X1 U7753 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6162), .ZN(n6662) );
  NAND2_X1 U7754 ( .A1(n6348), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n6164) );
  OAI21_X1 U7755 ( .B1(n6348), .B2(P2_REG1_REG_8__SCAN_IN), .A(n6164), .ZN(
        n6165) );
  NOR2_X1 U7756 ( .A1(n6166), .A2(n6165), .ZN(n6343) );
  AOI211_X1 U7757 ( .C1(n6166), .C2(n6165), .A(n6343), .B(n10407), .ZN(n6167)
         );
  AOI211_X1 U7758 ( .C1(P2_ADDR_REG_8__SCAN_IN), .C2(n10404), .A(n6662), .B(
        n6167), .ZN(n6175) );
  NAND2_X1 U7759 ( .A1(n6168), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6170) );
  NAND2_X1 U7760 ( .A1(n6170), .A2(n6169), .ZN(n6173) );
  MUX2_X1 U7761 ( .A(n6898), .B(P2_REG2_REG_8__SCAN_IN), .S(n6348), .Z(n6171)
         );
  INV_X1 U7762 ( .A(n6171), .ZN(n6172) );
  NAND2_X1 U7763 ( .A1(n6172), .A2(n6173), .ZN(n6349) );
  OAI211_X1 U7764 ( .C1(n6173), .C2(n6172), .A(n10403), .B(n6349), .ZN(n6174)
         );
  OAI211_X1 U7765 ( .C1(n10406), .C2(n6176), .A(n6175), .B(n6174), .ZN(
        P2_U3253) );
  INV_X1 U7766 ( .A(n7713), .ZN(n6188) );
  NAND2_X1 U7767 ( .A1(n6252), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6177) );
  XNOR2_X1 U7768 ( .A(n6177), .B(P1_IR_REG_15__SCAN_IN), .ZN(n7714) );
  INV_X1 U7769 ( .A(n9774), .ZN(n7535) );
  AOI22_X1 U7770 ( .A1(n7714), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n7535), .ZN(n6178) );
  OAI21_X1 U7771 ( .B1(n6188), .B2(n9773), .A(n6178), .ZN(P1_U3338) );
  INV_X1 U7772 ( .A(n10471), .ZN(n6792) );
  NAND2_X1 U7773 ( .A1(n6179), .A2(n10216), .ZN(n6181) );
  NAND2_X1 U7774 ( .A1(n8424), .A2(n8701), .ZN(n6180) );
  NAND2_X1 U7775 ( .A1(n6181), .A2(n6180), .ZN(n6795) );
  AOI22_X1 U7776 ( .A1(n10188), .A2(n6795), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        P2_U3152), .ZN(n6182) );
  OAI21_X1 U7777 ( .B1(n10199), .B2(P2_REG3_REG_3__SCAN_IN), .A(n6182), .ZN(
        n6186) );
  AOI211_X1 U7778 ( .C1(n6184), .C2(n6183), .A(n8156), .B(n6212), .ZN(n6185)
         );
  AOI211_X1 U7779 ( .C1(n8137), .C2(n6792), .A(n6186), .B(n6185), .ZN(n6187)
         );
  INV_X1 U7780 ( .A(n6187), .ZN(P2_U3220) );
  INV_X1 U7781 ( .A(n8464), .ZN(n8455) );
  OAI222_X1 U7782 ( .A1(n7510), .A2(n6189), .B1(n8872), .B2(n6188), .C1(
        P2_U3152), .C2(n8455), .ZN(P2_U3343) );
  AOI21_X1 U7783 ( .B1(n6192), .B2(n6191), .A(n6190), .ZN(n6199) );
  OAI21_X1 U7784 ( .B1(n6195), .B2(n6194), .A(n6193), .ZN(n6197) );
  AND2_X1 U7785 ( .A1(P1_U3084), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n8980) );
  NOR2_X1 U7786 ( .A1(n7444), .A2(n6414), .ZN(n6196) );
  AOI211_X1 U7787 ( .C1(n10332), .C2(n6197), .A(n8980), .B(n6196), .ZN(n6198)
         );
  OAI21_X1 U7788 ( .B1(n6199), .B2(n9385), .A(n6198), .ZN(n6200) );
  AOI211_X1 U7789 ( .C1(n10299), .C2(P1_ADDR_REG_4__SCAN_IN), .A(n6201), .B(
        n6200), .ZN(n6202) );
  INV_X1 U7790 ( .A(n6202), .ZN(P1_U3245) );
  NAND2_X1 U7791 ( .A1(n6204), .A2(n6203), .ZN(n6205) );
  OR2_X1 U7792 ( .A1(n6206), .A2(n6205), .ZN(n6766) );
  NAND2_X1 U7793 ( .A1(n6769), .A2(n6207), .ZN(n6208) );
  INV_X2 U7794 ( .A(n10494), .ZN(n10496) );
  INV_X1 U7795 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n6211) );
  NAND2_X1 U7796 ( .A1(n6209), .A2(n10496), .ZN(n6210) );
  OAI21_X1 U7797 ( .B1(n10496), .B2(n6211), .A(n6210), .ZN(P2_U3457) );
  AOI21_X1 U7798 ( .B1(n6217), .B2(n6212), .A(n6228), .ZN(n6222) );
  AOI22_X1 U7799 ( .A1(n7611), .A2(n8423), .B1(n8137), .B2(n6287), .ZN(n6215)
         );
  INV_X1 U7800 ( .A(n6213), .ZN(n6214) );
  OAI211_X1 U7801 ( .C1(n7083), .C2(n10199), .A(n6215), .B(n6214), .ZN(n6220)
         );
  NAND3_X1 U7802 ( .A1(n8057), .A2(n6217), .A3(n6216), .ZN(n6218) );
  INV_X1 U7803 ( .A(n8425), .ZN(n8064) );
  AOI21_X1 U7804 ( .B1(n6218), .B2(n8160), .A(n8064), .ZN(n6219) );
  NOR2_X1 U7805 ( .A1(n6220), .A2(n6219), .ZN(n6221) );
  OAI21_X1 U7806 ( .B1(n6222), .B2(n8156), .A(n6221), .ZN(P2_U3232) );
  INV_X1 U7807 ( .A(n7615), .ZN(n6234) );
  INV_X1 U7808 ( .A(n6223), .ZN(n6224) );
  OAI21_X1 U7809 ( .B1(n10199), .B2(n6225), .A(n6224), .ZN(n6227) );
  INV_X1 U7810 ( .A(n8424), .ZN(n6487) );
  OAI22_X1 U7811 ( .A1(n8160), .A2(n6487), .B1(n6515), .B2(n8167), .ZN(n6226)
         );
  AOI211_X1 U7812 ( .C1(n7611), .C2(n8422), .A(n6227), .B(n6226), .ZN(n6233)
         );
  OAI22_X1 U7813 ( .A1(n8142), .A2(n6487), .B1(n6229), .B2(n8156), .ZN(n6230)
         );
  NAND3_X1 U7814 ( .A1(n5040), .A2(n6231), .A3(n6230), .ZN(n6232) );
  OAI211_X1 U7815 ( .C1(n6234), .C2(n8156), .A(n6233), .B(n6232), .ZN(P2_U3229) );
  NAND2_X1 U7816 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_U3084), .ZN(n6241) );
  INV_X1 U7817 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n6235) );
  MUX2_X1 U7818 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n6235), .S(n7283), .Z(n6238)
         );
  INV_X1 U7819 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n10286) );
  AOI22_X1 U7820 ( .A1(P1_REG1_REG_11__SCAN_IN), .A2(n10323), .B1(n6244), .B2(
        n10286), .ZN(n10326) );
  OAI21_X1 U7821 ( .B1(P1_REG1_REG_10__SCAN_IN), .B2(n7002), .A(n6236), .ZN(
        n10327) );
  NAND2_X1 U7822 ( .A1(n10326), .A2(n10327), .ZN(n10325) );
  OAI21_X1 U7823 ( .B1(n10323), .B2(P1_REG1_REG_11__SCAN_IN), .A(n10325), .ZN(
        n6237) );
  NAND2_X1 U7824 ( .A1(n6238), .A2(n6237), .ZN(n6451) );
  OAI21_X1 U7825 ( .B1(n6238), .B2(n6237), .A(n6451), .ZN(n6239) );
  NAND2_X1 U7826 ( .A1(n10332), .A2(n6239), .ZN(n6240) );
  OAI211_X1 U7827 ( .C1(n7444), .C2(n6242), .A(n6241), .B(n6240), .ZN(n6249)
         );
  INV_X1 U7828 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n6243) );
  AOI22_X1 U7829 ( .A1(P1_REG2_REG_11__SCAN_IN), .A2(n10323), .B1(n6244), .B2(
        n6243), .ZN(n10329) );
  OAI21_X1 U7830 ( .B1(n10323), .B2(P1_REG2_REG_11__SCAN_IN), .A(n10328), .ZN(
        n6247) );
  NAND2_X1 U7831 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n7283), .ZN(n6245) );
  OAI21_X1 U7832 ( .B1(n7283), .B2(P1_REG2_REG_12__SCAN_IN), .A(n6245), .ZN(
        n6246) );
  NOR2_X1 U7833 ( .A1(n6246), .A2(n6247), .ZN(n6445) );
  AOI211_X1 U7834 ( .C1(n6247), .C2(n6246), .A(n6445), .B(n9385), .ZN(n6248)
         );
  AOI211_X1 U7835 ( .C1(P1_ADDR_REG_12__SCAN_IN), .C2(n10299), .A(n6249), .B(
        n6248), .ZN(n6250) );
  INV_X1 U7836 ( .A(n6250), .ZN(P1_U3253) );
  INV_X1 U7837 ( .A(n7725), .ZN(n6255) );
  AOI22_X1 U7838 ( .A1(n8480), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n8869), .ZN(n6251) );
  OAI21_X1 U7839 ( .B1(n6255), .B2(n8872), .A(n6251), .ZN(P2_U3342) );
  OR2_X1 U7840 ( .A1(n6252), .A2(P1_IR_REG_15__SCAN_IN), .ZN(n6253) );
  NAND2_X1 U7841 ( .A1(n6253), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6358) );
  XNOR2_X1 U7842 ( .A(n6358), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9366) );
  AOI22_X1 U7843 ( .A1(n9366), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n7535), .ZN(n6254) );
  OAI21_X1 U7844 ( .B1(n6255), .B2(n9773), .A(n6254), .ZN(P1_U3337) );
  NOR2_X1 U7845 ( .A1(P1_D_REG_3__SCAN_IN), .A2(P1_D_REG_4__SCAN_IN), .ZN(
        n6259) );
  NOR4_X1 U7846 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_2__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n6258) );
  NOR4_X1 U7847 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n6257) );
  NOR4_X1 U7848 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n6256) );
  NAND4_X1 U7849 ( .A1(n6259), .A2(n6258), .A3(n6257), .A4(n6256), .ZN(n6265)
         );
  NOR4_X1 U7850 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n6263) );
  NOR4_X1 U7851 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n6262) );
  NOR4_X1 U7852 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n6261) );
  NOR4_X1 U7853 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n6260) );
  NAND4_X1 U7854 ( .A1(n6263), .A2(n6262), .A3(n6261), .A4(n6260), .ZN(n6264)
         );
  OAI21_X1 U7855 ( .B1(n6265), .B2(n6264), .A(n9761), .ZN(n6599) );
  NAND2_X1 U7856 ( .A1(n6367), .A2(n6599), .ZN(n6266) );
  AOI21_X1 U7857 ( .B1(n10393), .B2(n9327), .A(n6266), .ZN(n6275) );
  OR2_X1 U7858 ( .A1(n6328), .A2(n6335), .ZN(n6619) );
  NAND2_X1 U7859 ( .A1(n6619), .A2(n9762), .ZN(n6365) );
  INV_X1 U7860 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n10107) );
  NAND2_X1 U7861 ( .A1(n9761), .A2(n10107), .ZN(n6267) );
  NAND2_X1 U7862 ( .A1(n7509), .A2(n7364), .ZN(n9764) );
  NAND2_X1 U7863 ( .A1(n6267), .A2(n9764), .ZN(n6366) );
  NOR2_X1 U7864 ( .A1(n6365), .A2(n6366), .ZN(n6268) );
  NAND2_X1 U7865 ( .A1(n6275), .A2(n6268), .ZN(n10399) );
  NAND2_X1 U7866 ( .A1(n9263), .A2(n9327), .ZN(n6373) );
  NOR2_X1 U7867 ( .A1(n9359), .A2(n6333), .ZN(n6320) );
  INV_X1 U7868 ( .A(n6320), .ZN(n6382) );
  NAND2_X1 U7869 ( .A1(n9359), .A2(n6333), .ZN(n9074) );
  NAND2_X1 U7870 ( .A1(n6382), .A2(n9074), .ZN(n9277) );
  NOR2_X1 U7871 ( .A1(n6380), .A2(n4485), .ZN(n6269) );
  NAND2_X1 U7872 ( .A1(n6269), .A2(n9338), .ZN(n6636) );
  INV_X1 U7873 ( .A(n6636), .ZN(n9336) );
  INV_X1 U7874 ( .A(n6373), .ZN(n6337) );
  NOR2_X1 U7875 ( .A1(n9336), .A2(n6337), .ZN(n6271) );
  INV_X1 U7876 ( .A(n6328), .ZN(n9264) );
  NAND2_X1 U7877 ( .A1(n7421), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n6270) );
  AOI22_X1 U7878 ( .A1(n9277), .A2(n6271), .B1(n10254), .B2(n9358), .ZN(n6376)
         );
  OAI21_X1 U7879 ( .B1(n6333), .B2(n6373), .A(n6376), .ZN(n6276) );
  NAND2_X1 U7880 ( .A1(n6276), .A2(n4483), .ZN(n6272) );
  OAI21_X1 U7881 ( .B1(n4483), .B2(n6273), .A(n6272), .ZN(P1_U3523) );
  INV_X1 U7882 ( .A(n6366), .ZN(n6600) );
  NOR2_X1 U7883 ( .A1(n6365), .A2(n6600), .ZN(n6274) );
  NAND2_X1 U7884 ( .A1(n6275), .A2(n6274), .ZN(n10394) );
  INV_X2 U7885 ( .A(n10394), .ZN(n10396) );
  INV_X1 U7886 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6278) );
  NAND2_X1 U7887 ( .A1(n6276), .A2(n10396), .ZN(n6277) );
  OAI21_X1 U7888 ( .B1(n10396), .B2(n6278), .A(n6277), .ZN(P1_U3454) );
  INV_X1 U7889 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n6291) );
  INV_X1 U7890 ( .A(n6179), .ZN(n6279) );
  NAND2_X1 U7891 ( .A1(n6279), .A2(n8063), .ZN(n6280) );
  NAND2_X1 U7892 ( .A1(n6281), .A2(n6280), .ZN(n6784) );
  NAND2_X1 U7893 ( .A1(n8425), .A2(n10471), .ZN(n8273) );
  NAND2_X1 U7894 ( .A1(n6784), .A2(n6783), .ZN(n6786) );
  NAND2_X1 U7895 ( .A1(n8064), .A2(n10471), .ZN(n6282) );
  INV_X1 U7896 ( .A(n6287), .ZN(n7088) );
  OR2_X1 U7897 ( .A1(n8424), .A2(n7088), .ZN(n8267) );
  NAND2_X1 U7898 ( .A1(n6283), .A2(n8199), .ZN(n6489) );
  OAI21_X1 U7899 ( .B1(n6283), .B2(n8199), .A(n6489), .ZN(n7090) );
  INV_X1 U7900 ( .A(n7090), .ZN(n6289) );
  NAND2_X1 U7901 ( .A1(n6794), .A2(n8263), .ZN(n6793) );
  XOR2_X1 U7902 ( .A(n8199), .B(n6483), .Z(n6285) );
  AOI222_X1 U7903 ( .A1(n10432), .A2(n6285), .B1(n8423), .B2(n8701), .C1(n8425), .C2(n10216), .ZN(n7092) );
  NAND2_X1 U7904 ( .A1(n6790), .A2(n10471), .ZN(n6789) );
  AND2_X1 U7905 ( .A1(n6789), .A2(n6287), .ZN(n6286) );
  NOR2_X1 U7906 ( .A1(n6503), .A2(n6286), .ZN(n7085) );
  AOI22_X1 U7907 ( .A1(n7085), .A2(n10418), .B1(n8803), .B2(n6287), .ZN(n6288)
         );
  OAI211_X1 U7908 ( .C1(n10466), .C2(n6289), .A(n7092), .B(n6288), .ZN(n6292)
         );
  NAND2_X1 U7909 ( .A1(n6292), .A2(n10496), .ZN(n6290) );
  OAI21_X1 U7910 ( .B1(n10496), .B2(n6291), .A(n6290), .ZN(P2_U3463) );
  INV_X1 U7911 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6294) );
  NAND2_X1 U7912 ( .A1(n6292), .A2(n10499), .ZN(n6293) );
  OAI21_X1 U7913 ( .B1(n10499), .B2(n6294), .A(n6293), .ZN(P2_U3524) );
  NAND2_X1 U7914 ( .A1(n7984), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n6298) );
  NAND2_X1 U7915 ( .A1(n4827), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6297) );
  NAND2_X1 U7916 ( .A1(n6404), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6296) );
  NAND2_X1 U7917 ( .A1(n7421), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n6295) );
  OR2_X1 U7918 ( .A1(n6409), .A2(n6299), .ZN(n6303) );
  OR2_X1 U7919 ( .A1(n6715), .A2(n6301), .ZN(n6302) );
  XNOR2_X2 U7920 ( .A(n9357), .B(n6690), .ZN(n9278) );
  INV_X1 U7921 ( .A(n6310), .ZN(n6334) );
  NAND2_X1 U7922 ( .A1(n9358), .A2(n6334), .ZN(n9073) );
  AND2_X1 U7923 ( .A1(n9359), .A2(n7599), .ZN(n6377) );
  NAND2_X1 U7924 ( .A1(n6319), .A2(n6377), .ZN(n6379) );
  NAND2_X1 U7925 ( .A1(n9358), .A2(n6310), .ZN(n6311) );
  NAND2_X1 U7926 ( .A1(n6379), .A2(n6311), .ZN(n6315) );
  INV_X1 U7927 ( .A(n6315), .ZN(n6313) );
  INV_X1 U7928 ( .A(n9278), .ZN(n6312) );
  INV_X1 U7929 ( .A(n6396), .ZN(n6314) );
  AOI21_X1 U7930 ( .B1(n9278), .B2(n6315), .A(n6314), .ZN(n6990) );
  INV_X1 U7931 ( .A(n10393), .ZN(n10375) );
  NAND2_X1 U7932 ( .A1(n9338), .A2(n4485), .ZN(n6318) );
  NAND2_X1 U7933 ( .A1(n5055), .A2(n6316), .ZN(n6317) );
  INV_X1 U7934 ( .A(n6319), .ZN(n6321) );
  NAND2_X1 U7935 ( .A1(n6321), .A2(n6320), .ZN(n6384) );
  NAND2_X1 U7936 ( .A1(n6384), .A2(n6322), .ZN(n6323) );
  INV_X1 U7937 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n6532) );
  NAND2_X1 U7938 ( .A1(n7984), .A2(n6532), .ZN(n6327) );
  NAND2_X1 U7939 ( .A1(n4481), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6326) );
  NAND2_X1 U7940 ( .A1(n6404), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6325) );
  NAND2_X1 U7941 ( .A1(n7421), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n6324) );
  NAND4_X1 U7942 ( .A1(n6327), .A2(n6326), .A3(n6325), .A4(n6324), .ZN(n9356)
         );
  OAI22_X1 U7943 ( .A1(n6423), .A2(n10350), .B1(n7603), .B2(n10352), .ZN(n6331) );
  NAND2_X1 U7944 ( .A1(n9338), .A2(n9544), .ZN(n6329) );
  NAND3_X1 U7945 ( .A1(n6636), .A2(n6589), .A3(n9544), .ZN(n10358) );
  NOR2_X1 U7946 ( .A1(n6990), .A2(n10358), .ZN(n6330) );
  AOI211_X1 U7947 ( .C1(n10355), .C2(n6332), .A(n6331), .B(n6330), .ZN(n6995)
         );
  NAND2_X1 U7948 ( .A1(n6334), .A2(n6333), .ZN(n6388) );
  OR2_X1 U7949 ( .A1(n6388), .A2(n6690), .ZN(n6430) );
  INV_X1 U7950 ( .A(n6430), .ZN(n6531) );
  AOI21_X1 U7951 ( .B1(n6690), .B2(n6388), .A(n6531), .ZN(n6993) );
  INV_X1 U7952 ( .A(n10388), .ZN(n9721) );
  INV_X1 U7953 ( .A(n6335), .ZN(n6336) );
  AOI22_X1 U7954 ( .A1(n6993), .A2(n9721), .B1(n10372), .B2(n6690), .ZN(n6338)
         );
  OAI211_X1 U7955 ( .C1(n6990), .C2(n10375), .A(n6995), .B(n6338), .ZN(n6340)
         );
  NAND2_X1 U7956 ( .A1(n6340), .A2(n4483), .ZN(n6339) );
  OAI21_X1 U7957 ( .B1(n4483), .B2(n5953), .A(n6339), .ZN(P1_U3525) );
  INV_X1 U7958 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n6342) );
  NAND2_X1 U7959 ( .A1(n6340), .A2(n10396), .ZN(n6341) );
  OAI21_X1 U7960 ( .B1(n10396), .B2(n6342), .A(n6341), .ZN(P1_U3460) );
  NOR2_X1 U7961 ( .A1(n5368), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8112) );
  NAND2_X1 U7962 ( .A1(n6650), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n6344) );
  OAI21_X1 U7963 ( .B1(n6650), .B2(P2_REG1_REG_9__SCAN_IN), .A(n6344), .ZN(
        n6345) );
  AOI211_X1 U7964 ( .C1(n6346), .C2(n6345), .A(n6645), .B(n10407), .ZN(n6347)
         );
  AOI211_X1 U7965 ( .C1(P2_ADDR_REG_9__SCAN_IN), .C2(n10404), .A(n8112), .B(
        n6347), .ZN(n6355) );
  NAND2_X1 U7966 ( .A1(n6348), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n6350) );
  NAND2_X1 U7967 ( .A1(n6350), .A2(n6349), .ZN(n6353) );
  MUX2_X1 U7968 ( .A(n5367), .B(P2_REG2_REG_9__SCAN_IN), .S(n6650), .Z(n6351)
         );
  INV_X1 U7969 ( .A(n6351), .ZN(n6352) );
  NAND2_X1 U7970 ( .A1(n6352), .A2(n6353), .ZN(n6651) );
  OAI211_X1 U7971 ( .C1(n6353), .C2(n6352), .A(n10403), .B(n6651), .ZN(n6354)
         );
  OAI211_X1 U7972 ( .C1(n10406), .C2(n6356), .A(n6355), .B(n6354), .ZN(
        P2_U3254) );
  INV_X1 U7973 ( .A(n7747), .ZN(n6393) );
  NAND2_X1 U7974 ( .A1(n6358), .A2(n6357), .ZN(n6359) );
  NAND2_X1 U7975 ( .A1(n6359), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6362) );
  INV_X1 U7976 ( .A(n6362), .ZN(n6360) );
  NAND2_X1 U7977 ( .A1(n6360), .A2(P1_IR_REG_17__SCAN_IN), .ZN(n6363) );
  NAND2_X1 U7978 ( .A1(n6362), .A2(n6361), .ZN(n6441) );
  AOI22_X1 U7979 ( .A1(n9383), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n7535), .ZN(n6364) );
  OAI21_X1 U7980 ( .B1(n6393), .B2(n9773), .A(n6364), .ZN(P1_U3336) );
  INV_X1 U7981 ( .A(n6365), .ZN(n6679) );
  NAND2_X1 U7982 ( .A1(n6366), .A2(n6599), .ZN(n6368) );
  NOR2_X1 U7983 ( .A1(n6368), .A2(n6367), .ZN(n6369) );
  NAND2_X1 U7984 ( .A1(n6679), .A2(n6369), .ZN(n6371) );
  AND2_X1 U7985 ( .A1(n9762), .A2(n9327), .ZN(n6370) );
  AOI22_X1 U7986 ( .A1(n10362), .A2(P1_REG2_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(n10360), .ZN(n6375) );
  NOR2_X1 U7987 ( .A1(n6371), .A2(n4485), .ZN(n9626) );
  INV_X1 U7988 ( .A(n9626), .ZN(n6372) );
  OR2_X1 U7989 ( .A1(n6372), .A2(n10388), .ZN(n9651) );
  NOR2_X1 U7990 ( .A1(n6373), .A2(n6945), .ZN(n6623) );
  OAI21_X1 U7991 ( .B1(n10343), .B2(n9648), .A(n7599), .ZN(n6374) );
  OAI211_X1 U7992 ( .C1(n6376), .C2(n10362), .A(n6375), .B(n6374), .ZN(
        P1_U3291) );
  OR2_X1 U7993 ( .A1(n6319), .A2(n6377), .ZN(n6378) );
  NAND2_X1 U7994 ( .A1(n6379), .A2(n6378), .ZN(n10376) );
  NOR2_X1 U7995 ( .A1(n6380), .A2(n9544), .ZN(n6381) );
  AND2_X1 U7996 ( .A1(n10366), .A2(n6381), .ZN(n10344) );
  INV_X1 U7997 ( .A(n10344), .ZN(n7154) );
  AOI22_X1 U7998 ( .A1(n10252), .A2(n9359), .B1(n9357), .B2(n10254), .ZN(n6387) );
  NAND2_X1 U7999 ( .A1(n6382), .A2(n6319), .ZN(n6383) );
  NAND2_X1 U8000 ( .A1(n6384), .A2(n6383), .ZN(n6385) );
  NAND2_X1 U8001 ( .A1(n6385), .A2(n10355), .ZN(n6386) );
  OAI211_X1 U8002 ( .C1(n10376), .C2(n10358), .A(n6387), .B(n6386), .ZN(n10378) );
  AOI21_X1 U8003 ( .B1(n6310), .B2(n7599), .A(n10388), .ZN(n6389) );
  NAND2_X1 U8004 ( .A1(n6389), .A2(n6388), .ZN(n10374) );
  OAI22_X1 U8005 ( .A1(n10374), .A2(n4485), .B1(n9555), .B2(n6069), .ZN(n6390)
         );
  OAI21_X1 U8006 ( .B1(n10378), .B2(n6390), .A(n10366), .ZN(n6392) );
  AOI22_X1 U8007 ( .A1(n9648), .A2(n6310), .B1(n10362), .B2(
        P1_REG2_REG_1__SCAN_IN), .ZN(n6391) );
  OAI211_X1 U8008 ( .C1(n10376), .C2(n7154), .A(n6392), .B(n6391), .ZN(
        P1_U3290) );
  INV_X1 U8009 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n6394) );
  OAI222_X1 U8010 ( .A1(n7510), .A2(n6394), .B1(n8872), .B2(n6393), .C1(n8493), 
        .C2(P2_U3152), .ZN(P2_U3341) );
  INV_X1 U8011 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n6436) );
  INV_X1 U8012 ( .A(n9357), .ZN(n6525) );
  INV_X1 U8013 ( .A(n6690), .ZN(n9076) );
  NAND2_X1 U8014 ( .A1(n6525), .A2(n9076), .ZN(n6395) );
  NAND2_X1 U8015 ( .A1(n6396), .A2(n6395), .ZN(n6524) );
  OR2_X1 U8016 ( .A1(n6409), .A2(n6397), .ZN(n6400) );
  OR2_X1 U8017 ( .A1(n6715), .A2(n6398), .ZN(n6399) );
  OAI211_X1 U8018 ( .C1(n6842), .C2(n6401), .A(n6400), .B(n6399), .ZN(n6807)
         );
  NAND2_X1 U8019 ( .A1(n6423), .A2(n6807), .ZN(n9072) );
  INV_X1 U8020 ( .A(n6807), .ZN(n10380) );
  NAND2_X1 U8021 ( .A1(n9356), .A2(n10380), .ZN(n9078) );
  NAND2_X1 U8022 ( .A1(n6524), .A2(n9276), .ZN(n6523) );
  NAND2_X1 U8023 ( .A1(n6423), .A2(n10380), .ZN(n6402) );
  NAND2_X1 U8024 ( .A1(n6523), .A2(n6402), .ZN(n6415) );
  NAND2_X1 U8025 ( .A1(n4481), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6408) );
  INV_X1 U8026 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n6403) );
  XNOR2_X1 U8027 ( .A(n6403), .B(P1_REG3_REG_3__SCAN_IN), .ZN(n8982) );
  NAND2_X1 U8028 ( .A1(n7984), .A2(n8982), .ZN(n6407) );
  NAND2_X1 U8029 ( .A1(n6404), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6406) );
  NAND2_X1 U8030 ( .A1(n4480), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n6405) );
  NAND4_X1 U8031 ( .A1(n6408), .A2(n6407), .A3(n6406), .A4(n6405), .ZN(n9355)
         );
  INV_X1 U8032 ( .A(n9355), .ZN(n6526) );
  OR2_X1 U8033 ( .A1(n6409), .A2(n6410), .ZN(n6413) );
  OAI211_X1 U8034 ( .C1(n6842), .C2(n6414), .A(n6413), .B(n6412), .ZN(n8981)
         );
  NAND2_X1 U8035 ( .A1(n6526), .A2(n8981), .ZN(n9079) );
  NAND2_X1 U8036 ( .A1(n9355), .A2(n6631), .ZN(n9307) );
  NAND2_X1 U8037 ( .A1(n9079), .A2(n9307), .ZN(n9275) );
  OAI21_X1 U8038 ( .B1(n6415), .B2(n9275), .A(n6459), .ZN(n6633) );
  INV_X1 U8039 ( .A(n6633), .ZN(n6434) );
  INV_X1 U8040 ( .A(n10358), .ZN(n6699) );
  NAND2_X1 U8041 ( .A1(n4481), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6422) );
  NAND3_X1 U8042 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n6467) );
  INV_X1 U8043 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n6417) );
  NAND2_X1 U8044 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n6416) );
  NAND2_X1 U8045 ( .A1(n6417), .A2(n6416), .ZN(n6418) );
  AND2_X1 U8046 ( .A1(n6467), .A2(n6418), .ZN(n8951) );
  NAND2_X1 U8047 ( .A1(n7984), .A2(n8951), .ZN(n6421) );
  NAND2_X1 U8048 ( .A1(n4480), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n6420) );
  NAND2_X1 U8049 ( .A1(n6404), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6419) );
  NAND4_X1 U8050 ( .A1(n6422), .A2(n6421), .A3(n6420), .A4(n6419), .ZN(n9354)
         );
  INV_X1 U8051 ( .A(n9354), .ZN(n6615) );
  OAI22_X1 U8052 ( .A1(n6423), .A2(n10352), .B1(n6615), .B2(n10350), .ZN(n6429) );
  NAND2_X1 U8053 ( .A1(n6525), .A2(n6690), .ZN(n6424) );
  INV_X1 U8054 ( .A(n9276), .ZN(n6425) );
  NAND2_X1 U8055 ( .A1(n9306), .A2(n6425), .ZN(n6426) );
  XNOR2_X1 U8056 ( .A(n9127), .B(n9275), .ZN(n6427) );
  NOR2_X1 U8057 ( .A1(n6427), .A2(n9620), .ZN(n6428) );
  AOI211_X1 U8058 ( .C1(n6699), .C2(n6633), .A(n6429), .B(n6428), .ZN(n6635)
         );
  NOR2_X1 U8059 ( .A1(n6430), .A2(n6807), .ZN(n6431) );
  INV_X1 U8060 ( .A(n6431), .ZN(n6530) );
  NAND2_X1 U8061 ( .A1(n6431), .A2(n6631), .ZN(n6474) );
  INV_X1 U8062 ( .A(n6474), .ZN(n6432) );
  AOI21_X1 U8063 ( .B1(n8981), .B2(n6530), .A(n6432), .ZN(n6628) );
  AOI22_X1 U8064 ( .A1(n6628), .A2(n9721), .B1(n10372), .B2(n8981), .ZN(n6433)
         );
  OAI211_X1 U8065 ( .C1(n6434), .C2(n10375), .A(n6635), .B(n6433), .ZN(n6437)
         );
  NAND2_X1 U8066 ( .A1(n6437), .A2(n10396), .ZN(n6435) );
  OAI21_X1 U8067 ( .B1(n10396), .B2(n6436), .A(n6435), .ZN(P1_U3466) );
  NAND2_X1 U8068 ( .A1(n6437), .A2(n4483), .ZN(n6438) );
  OAI21_X1 U8069 ( .B1(n4483), .B2(n6439), .A(n6438), .ZN(P1_U3527) );
  INV_X1 U8070 ( .A(n7766), .ZN(n6444) );
  AOI22_X1 U8071 ( .A1(n8512), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n8869), .ZN(n6440) );
  OAI21_X1 U8072 ( .B1(n6444), .B2(n8872), .A(n6440), .ZN(P2_U3340) );
  NAND2_X1 U8073 ( .A1(n6441), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6442) );
  XNOR2_X1 U8074 ( .A(n6442), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9395) );
  AOI22_X1 U8075 ( .A1(n9395), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n7535), .ZN(n6443) );
  OAI21_X1 U8076 ( .B1(n6444), .B2(n9773), .A(n6443), .ZN(P1_U3335) );
  INV_X1 U8077 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n6457) );
  NAND2_X1 U8078 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n7373), .ZN(n6446) );
  OAI21_X1 U8079 ( .B1(n7373), .B2(P1_REG2_REG_13__SCAN_IN), .A(n6446), .ZN(
        n6447) );
  AOI211_X1 U8080 ( .C1(n6448), .C2(n6447), .A(n7051), .B(n9385), .ZN(n6449)
         );
  AOI21_X1 U8081 ( .B1(n10324), .B2(n7373), .A(n6449), .ZN(n6456) );
  INV_X1 U8082 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n6450) );
  MUX2_X1 U8083 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n6450), .S(n7373), .Z(n6453)
         );
  OAI21_X1 U8084 ( .B1(n7283), .B2(P1_REG1_REG_12__SCAN_IN), .A(n6451), .ZN(
        n6452) );
  NAND2_X1 U8085 ( .A1(n6453), .A2(n6452), .ZN(n7046) );
  OAI21_X1 U8086 ( .B1(n6453), .B2(n6452), .A(n7046), .ZN(n6454) );
  AND2_X1 U8087 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n7389) );
  AOI21_X1 U8088 ( .B1(n10332), .B2(n6454), .A(n7389), .ZN(n6455) );
  OAI211_X1 U8089 ( .C1(n10337), .C2(n6457), .A(n6456), .B(n6455), .ZN(
        P1_U3254) );
  INV_X1 U8090 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n6478) );
  NAND2_X1 U8091 ( .A1(n6526), .A2(n6631), .ZN(n6458) );
  OR2_X1 U8092 ( .A1(n6409), .A2(n6460), .ZN(n6463) );
  OR2_X1 U8093 ( .A1(n6715), .A2(n6461), .ZN(n6462) );
  NAND2_X1 U8094 ( .A1(n6615), .A2(n8950), .ZN(n9125) );
  INV_X1 U8095 ( .A(n4501), .ZN(n6694) );
  OAI21_X1 U8096 ( .B1(n4495), .B2(n6694), .A(n4993), .ZN(n6644) );
  INV_X1 U8097 ( .A(n9079), .ZN(n9309) );
  XNOR2_X1 U8098 ( .A(n6725), .B(n6694), .ZN(n6473) );
  NAND2_X1 U8099 ( .A1(n4481), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6472) );
  INV_X1 U8100 ( .A(n6467), .ZN(n6465) );
  NAND2_X1 U8101 ( .A1(n6467), .A2(n6466), .ZN(n6468) );
  AND2_X1 U8102 ( .A1(n6606), .A2(n6468), .ZN(n6706) );
  NAND2_X1 U8103 ( .A1(n7984), .A2(n6706), .ZN(n6471) );
  NAND2_X1 U8104 ( .A1(n4480), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n6470) );
  NAND2_X1 U8105 ( .A1(n9118), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6469) );
  NAND4_X1 U8106 ( .A1(n6472), .A2(n6471), .A3(n6470), .A4(n6469), .ZN(n9353)
         );
  AOI222_X1 U8107 ( .A1(n10355), .A2(n6473), .B1(n9353), .B2(n10254), .C1(
        n9355), .C2(n10252), .ZN(n6640) );
  AOI21_X1 U8108 ( .B1(n6474), .B2(n8950), .A(n10388), .ZN(n6475) );
  OR2_X1 U8109 ( .A1(n6474), .A2(n8950), .ZN(n6704) );
  AND2_X1 U8110 ( .A1(n6475), .A2(n6704), .ZN(n6638) );
  AOI21_X1 U8111 ( .B1(n10372), .B2(n8950), .A(n6638), .ZN(n6476) );
  OAI211_X1 U8112 ( .C1(n9742), .C2(n6644), .A(n6640), .B(n6476), .ZN(n6479)
         );
  NAND2_X1 U8113 ( .A1(n6479), .A2(n10396), .ZN(n6477) );
  OAI21_X1 U8114 ( .B1(n10396), .B2(n6478), .A(n6477), .ZN(P1_U3469) );
  NAND2_X1 U8115 ( .A1(n6479), .A2(n4483), .ZN(n6480) );
  OAI21_X1 U8116 ( .B1(n4483), .B2(n6481), .A(n6480), .ZN(P1_U3528) );
  OR2_X1 U8117 ( .A1(n6482), .A2(n6813), .ZN(n8279) );
  NAND2_X1 U8118 ( .A1(n6482), .A2(n6813), .ZN(n8282) );
  NAND2_X1 U8119 ( .A1(n7608), .A2(n10444), .ZN(n8268) );
  NAND2_X1 U8120 ( .A1(n6515), .A2(n8423), .ZN(n8275) );
  NAND2_X1 U8121 ( .A1(n8268), .A2(n8275), .ZN(n8201) );
  NAND2_X1 U8122 ( .A1(n6499), .A2(n8268), .ZN(n6484) );
  OAI21_X1 U8123 ( .B1(n8202), .B2(n6484), .A(n6818), .ZN(n6485) );
  AOI222_X1 U8124 ( .A1(n10432), .A2(n6485), .B1(n8421), .B2(n8701), .C1(n8423), .C2(n10216), .ZN(n6486) );
  INV_X1 U8125 ( .A(n6486), .ZN(n7095) );
  NAND2_X1 U8126 ( .A1(n6503), .A2(n6515), .ZN(n6504) );
  OR2_X1 U8127 ( .A1(n6504), .A2(n6813), .ZN(n6822) );
  INV_X1 U8128 ( .A(n6822), .ZN(n6823) );
  AOI211_X1 U8129 ( .C1(n6813), .C2(n6504), .A(n10472), .B(n6823), .ZN(n7093)
         );
  NOR2_X1 U8130 ( .A1(n7095), .A2(n7093), .ZN(n6522) );
  NAND2_X1 U8131 ( .A1(n10496), .A2(n10485), .ZN(n8860) );
  INV_X1 U8132 ( .A(n8860), .ZN(n6512) );
  NAND2_X1 U8133 ( .A1(n6487), .A2(n7088), .ZN(n6488) );
  NAND2_X1 U8134 ( .A1(n6489), .A2(n6488), .ZN(n6507) );
  NAND2_X1 U8135 ( .A1(n6507), .A2(n8201), .ZN(n6509) );
  NAND2_X1 U8136 ( .A1(n7608), .A2(n6515), .ZN(n6490) );
  NAND2_X1 U8137 ( .A1(n6509), .A2(n6490), .ZN(n6492) );
  INV_X1 U8138 ( .A(n8202), .ZN(n6491) );
  NAND2_X1 U8139 ( .A1(n6492), .A2(n6491), .ZN(n6815) );
  OR2_X1 U8140 ( .A1(n6492), .A2(n6491), .ZN(n6493) );
  NAND2_X1 U8141 ( .A1(n6815), .A2(n6493), .ZN(n7098) );
  INV_X1 U8142 ( .A(n8844), .ZN(n8847) );
  INV_X1 U8143 ( .A(n6813), .ZN(n7607) );
  INV_X1 U8144 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n6494) );
  OAI22_X1 U8145 ( .A1(n8847), .A2(n7607), .B1(n10496), .B2(n6494), .ZN(n6495)
         );
  AOI21_X1 U8146 ( .B1(n6512), .B2(n7098), .A(n6495), .ZN(n6496) );
  OAI21_X1 U8147 ( .B1(n6522), .B2(n10494), .A(n6496), .ZN(P2_U3469) );
  NAND2_X1 U8148 ( .A1(n6497), .A2(n8201), .ZN(n6498) );
  NAND2_X1 U8149 ( .A1(n6499), .A2(n6498), .ZN(n6500) );
  NAND2_X1 U8150 ( .A1(n6500), .A2(n10432), .ZN(n6502) );
  AOI22_X1 U8151 ( .A1(n10216), .A2(n8424), .B1(n8422), .B2(n8701), .ZN(n6501)
         );
  NAND2_X1 U8152 ( .A1(n6502), .A2(n6501), .ZN(n10452) );
  INV_X1 U8153 ( .A(n6503), .ZN(n6506) );
  INV_X1 U8154 ( .A(n6504), .ZN(n6505) );
  AOI211_X1 U8155 ( .C1(n10444), .C2(n6506), .A(n10472), .B(n6505), .ZN(n10443) );
  NOR2_X1 U8156 ( .A1(n10452), .A2(n10443), .ZN(n6518) );
  OR2_X1 U8157 ( .A1(n6507), .A2(n8201), .ZN(n6508) );
  NAND2_X1 U8158 ( .A1(n6509), .A2(n6508), .ZN(n10453) );
  INV_X1 U8159 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n6510) );
  OAI22_X1 U8160 ( .A1(n8847), .A2(n6515), .B1(n10496), .B2(n6510), .ZN(n6511)
         );
  AOI21_X1 U8161 ( .B1(n6512), .B2(n10453), .A(n6511), .ZN(n6513) );
  OAI21_X1 U8162 ( .B1(n6518), .B2(n10494), .A(n6513), .ZN(P2_U3466) );
  NAND2_X1 U8163 ( .A1(n10499), .A2(n10485), .ZN(n8791) );
  INV_X1 U8164 ( .A(n8791), .ZN(n6520) );
  INV_X1 U8165 ( .A(n8773), .ZN(n8776) );
  INV_X1 U8166 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6514) );
  OAI22_X1 U8167 ( .A1(n8776), .A2(n6515), .B1(n10499), .B2(n6514), .ZN(n6516)
         );
  AOI21_X1 U8168 ( .B1(n6520), .B2(n10453), .A(n6516), .ZN(n6517) );
  OAI21_X1 U8169 ( .B1(n6518), .B2(n10504), .A(n6517), .ZN(P2_U3525) );
  OAI22_X1 U8170 ( .A1(n8776), .A2(n7607), .B1(n10499), .B2(n5879), .ZN(n6519)
         );
  AOI21_X1 U8171 ( .B1(n7098), .B2(n6520), .A(n6519), .ZN(n6521) );
  OAI21_X1 U8172 ( .B1(n6522), .B2(n10504), .A(n6521), .ZN(P2_U3526) );
  XNOR2_X1 U8173 ( .A(n9306), .B(n9276), .ZN(n6529) );
  OAI21_X1 U8174 ( .B1(n6524), .B2(n9276), .A(n6523), .ZN(n10384) );
  OAI22_X1 U8175 ( .A1(n6526), .A2(n10350), .B1(n6525), .B2(n10352), .ZN(n6527) );
  AOI21_X1 U8176 ( .B1(n10384), .B2(n6699), .A(n6527), .ZN(n6528) );
  OAI21_X1 U8177 ( .B1(n9620), .B2(n6529), .A(n6528), .ZN(n10382) );
  INV_X1 U8178 ( .A(n10382), .ZN(n6537) );
  OAI21_X1 U8179 ( .B1(n10380), .B2(n6531), .A(n6530), .ZN(n10381) );
  AOI22_X1 U8180 ( .A1(n10362), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n10360), .B2(
        n6532), .ZN(n6534) );
  NAND2_X1 U8181 ( .A1(n9648), .A2(n6807), .ZN(n6533) );
  OAI211_X1 U8182 ( .C1(n10381), .C2(n9651), .A(n6534), .B(n6533), .ZN(n6535)
         );
  AOI21_X1 U8183 ( .B1(n10384), .B2(n10344), .A(n6535), .ZN(n6536) );
  OAI21_X1 U8184 ( .B1(n6537), .B2(n10362), .A(n6536), .ZN(P1_U3288) );
  NAND2_X1 U8185 ( .A1(n6539), .A2(n6589), .ZN(n6541) );
  NAND2_X1 U8186 ( .A1(n9358), .A2(n7890), .ZN(n6543) );
  NAND2_X1 U8187 ( .A1(n6310), .A2(n7961), .ZN(n6542) );
  NAND2_X1 U8188 ( .A1(n6543), .A2(n6542), .ZN(n6544) );
  NAND2_X1 U8189 ( .A1(n6675), .A2(n6548), .ZN(n6547) );
  NAND2_X1 U8190 ( .A1(n9358), .A2(n7320), .ZN(n6546) );
  NAND2_X1 U8191 ( .A1(n6310), .A2(n7973), .ZN(n6545) );
  NAND2_X1 U8192 ( .A1(n6546), .A2(n6545), .ZN(n6674) );
  INV_X1 U8193 ( .A(n6675), .ZN(n6549) );
  NAND2_X1 U8194 ( .A1(n9357), .A2(n7890), .ZN(n6551) );
  NAND2_X1 U8195 ( .A1(n6690), .A2(n7750), .ZN(n6550) );
  NAND2_X1 U8196 ( .A1(n6551), .A2(n6550), .ZN(n6552) );
  XNOR2_X1 U8197 ( .A(n6552), .B(n6576), .ZN(n6554) );
  INV_X1 U8198 ( .A(n6554), .ZN(n6557) );
  INV_X1 U8199 ( .A(n6555), .ZN(n6556) );
  NAND2_X1 U8200 ( .A1(n9356), .A2(n7973), .ZN(n6561) );
  NAND2_X1 U8201 ( .A1(n6807), .A2(n7961), .ZN(n6560) );
  NAND2_X1 U8202 ( .A1(n6561), .A2(n6560), .ZN(n6562) );
  XNOR2_X1 U8203 ( .A(n6562), .B(n6589), .ZN(n6567) );
  AOI22_X1 U8204 ( .A1(n9356), .A2(n7320), .B1(n7936), .B2(n6807), .ZN(n6568)
         );
  XNOR2_X1 U8205 ( .A(n6567), .B(n6568), .ZN(n6804) );
  NAND2_X1 U8206 ( .A1(n9355), .A2(n7973), .ZN(n6564) );
  NAND2_X1 U8207 ( .A1(n8981), .A2(n7961), .ZN(n6563) );
  NAND2_X1 U8208 ( .A1(n6564), .A2(n6563), .ZN(n6565) );
  XNOR2_X1 U8209 ( .A(n6565), .B(n6589), .ZN(n6572) );
  AOI22_X1 U8210 ( .A1(n9355), .A2(n7320), .B1(n7936), .B2(n8981), .ZN(n6570)
         );
  XNOR2_X1 U8211 ( .A(n6572), .B(n6570), .ZN(n8978) );
  INV_X1 U8212 ( .A(n6567), .ZN(n6569) );
  NAND2_X1 U8213 ( .A1(n6569), .A2(n6568), .ZN(n8974) );
  INV_X1 U8214 ( .A(n6570), .ZN(n6571) );
  NAND2_X1 U8215 ( .A1(n6572), .A2(n6571), .ZN(n6573) );
  NAND2_X1 U8216 ( .A1(n9354), .A2(n7936), .ZN(n6575) );
  NAND2_X1 U8217 ( .A1(n8950), .A2(n7750), .ZN(n6574) );
  NAND2_X1 U8218 ( .A1(n6575), .A2(n6574), .ZN(n6577) );
  XNOR2_X1 U8219 ( .A(n6577), .B(n7956), .ZN(n6744) );
  INV_X1 U8220 ( .A(n6744), .ZN(n6578) );
  NOR2_X1 U8221 ( .A1(n6747), .A2(n6578), .ZN(n6581) );
  AOI21_X1 U8222 ( .B1(n6747), .B2(n6578), .A(n6581), .ZN(n8946) );
  NAND2_X1 U8223 ( .A1(n9354), .A2(n7320), .ZN(n6580) );
  NAND2_X1 U8224 ( .A1(n8950), .A2(n7936), .ZN(n6579) );
  AND2_X1 U8225 ( .A1(n6580), .A2(n6579), .ZN(n8947) );
  NAND2_X1 U8226 ( .A1(n8946), .A2(n8947), .ZN(n8945) );
  INV_X1 U8227 ( .A(n6581), .ZN(n6582) );
  NAND2_X1 U8228 ( .A1(n8945), .A2(n6582), .ZN(n6598) );
  NAND2_X1 U8229 ( .A1(n9353), .A2(n7936), .ZN(n6588) );
  OR2_X1 U8230 ( .A1(n6715), .A2(n6583), .ZN(n6585) );
  OR2_X1 U8231 ( .A1(n6409), .A2(n9930), .ZN(n6584) );
  NAND2_X1 U8232 ( .A1(n6707), .A2(n7961), .ZN(n6587) );
  NAND2_X1 U8233 ( .A1(n6588), .A2(n6587), .ZN(n6590) );
  XNOR2_X1 U8234 ( .A(n6590), .B(n6589), .ZN(n6596) );
  INV_X1 U8235 ( .A(n6596), .ZN(n6594) );
  NAND2_X1 U8236 ( .A1(n9353), .A2(n7320), .ZN(n6592) );
  NAND2_X1 U8237 ( .A1(n6707), .A2(n7936), .ZN(n6591) );
  NAND2_X1 U8238 ( .A1(n6592), .A2(n6591), .ZN(n6595) );
  INV_X1 U8239 ( .A(n6595), .ZN(n6593) );
  NAND2_X1 U8240 ( .A1(n6596), .A2(n6595), .ZN(n6743) );
  NAND2_X1 U8241 ( .A1(n4565), .A2(n6743), .ZN(n6597) );
  XNOR2_X1 U8242 ( .A(n6598), .B(n6597), .ZN(n6627) );
  NAND3_X1 U8243 ( .A1(n6601), .A2(n6600), .A3(n6599), .ZN(n6622) );
  INV_X1 U8244 ( .A(n9762), .ZN(n6602) );
  OR2_X1 U8245 ( .A1(n10372), .A2(n9264), .ZN(n6603) );
  NOR2_X1 U8246 ( .A1(n6613), .A2(n6636), .ZN(n6614) );
  NAND2_X1 U8247 ( .A1(n4481), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6611) );
  INV_X1 U8248 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n6605) );
  NAND2_X1 U8249 ( .A1(n6606), .A2(n6605), .ZN(n6607) );
  AND2_X1 U8250 ( .A1(n6729), .A2(n6607), .ZN(n6978) );
  NAND2_X1 U8251 ( .A1(n7984), .A2(n6978), .ZN(n6610) );
  NAND2_X1 U8252 ( .A1(n4480), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n6609) );
  NAND2_X1 U8253 ( .A1(n9118), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6608) );
  NAND4_X1 U8254 ( .A1(n6611), .A2(n6610), .A3(n6609), .A4(n6608), .ZN(n9352)
         );
  INV_X1 U8255 ( .A(n6623), .ZN(n6612) );
  INV_X1 U8256 ( .A(n6707), .ZN(n6829) );
  NAND2_X1 U8257 ( .A1(n6614), .A2(n9335), .ZN(n9026) );
  OAI22_X1 U8258 ( .A1(n9019), .A2(n6829), .B1(n9026), .B2(n6615), .ZN(n6616)
         );
  AOI211_X1 U8259 ( .C1(n9030), .C2(n9352), .A(n6617), .B(n6616), .ZN(n6626)
         );
  AND3_X1 U8260 ( .A1(n6619), .A2(n6618), .A3(n7246), .ZN(n6620) );
  NAND2_X1 U8261 ( .A1(n6622), .A2(n10386), .ZN(n6678) );
  NAND2_X1 U8262 ( .A1(n6620), .A2(n6678), .ZN(n6621) );
  NAND2_X1 U8263 ( .A1(n6621), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6624) );
  NAND3_X1 U8264 ( .A1(n6623), .A2(n6622), .A3(n9762), .ZN(n6680) );
  NAND2_X1 U8265 ( .A1(n6624), .A2(n6680), .ZN(n9042) );
  NAND2_X1 U8266 ( .A1(n9042), .A2(n6706), .ZN(n6625) );
  OAI211_X1 U8267 ( .C1(n6627), .C2(n9049), .A(n6626), .B(n6625), .ZN(P1_U3237) );
  NAND2_X1 U8268 ( .A1(n6628), .A2(n10343), .ZN(n6630) );
  AOI22_X1 U8269 ( .A1(n10362), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n8982), .B2(
        n10360), .ZN(n6629) );
  OAI211_X1 U8270 ( .C1(n6631), .C2(n10364), .A(n6630), .B(n6629), .ZN(n6632)
         );
  AOI21_X1 U8271 ( .B1(n6633), .B2(n10344), .A(n6632), .ZN(n6634) );
  OAI21_X1 U8272 ( .B1(n6635), .B2(n10362), .A(n6634), .ZN(P1_U3287) );
  AND2_X1 U8273 ( .A1(n6636), .A2(n6589), .ZN(n6637) );
  NAND2_X1 U8274 ( .A1(n10366), .A2(n6637), .ZN(n9633) );
  AOI22_X1 U8275 ( .A1(n6638), .A2(n9544), .B1(n10360), .B2(n8951), .ZN(n6639)
         );
  AOI21_X1 U8276 ( .B1(n6640), .B2(n6639), .A(n10362), .ZN(n6641) );
  INV_X1 U8277 ( .A(n6641), .ZN(n6643) );
  AOI22_X1 U8278 ( .A1(n9648), .A2(n8950), .B1(n10362), .B2(
        P1_REG2_REG_5__SCAN_IN), .ZN(n6642) );
  OAI211_X1 U8279 ( .C1(n6644), .C2(n9633), .A(n6643), .B(n6642), .ZN(P1_U3286) );
  NOR2_X1 U8280 ( .A1(n10062), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7059) );
  INV_X1 U8281 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n6646) );
  MUX2_X1 U8282 ( .A(n6646), .B(P2_REG1_REG_10__SCAN_IN), .S(n7036), .Z(n6647)
         );
  AOI211_X1 U8283 ( .C1(n6648), .C2(n6647), .A(n7035), .B(n10407), .ZN(n6649)
         );
  AOI211_X1 U8284 ( .C1(P2_ADDR_REG_10__SCAN_IN), .C2(n10404), .A(n7059), .B(
        n6649), .ZN(n6657) );
  NAND2_X1 U8285 ( .A1(n6650), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6652) );
  NAND2_X1 U8286 ( .A1(n6652), .A2(n6651), .ZN(n6655) );
  MUX2_X1 U8287 ( .A(n5394), .B(P2_REG2_REG_10__SCAN_IN), .S(n7036), .Z(n6653)
         );
  INV_X1 U8288 ( .A(n6653), .ZN(n6654) );
  NAND2_X1 U8289 ( .A1(n6654), .A2(n6655), .ZN(n7029) );
  OAI211_X1 U8290 ( .C1(n6655), .C2(n6654), .A(n10403), .B(n7029), .ZN(n6656)
         );
  OAI211_X1 U8291 ( .C1(n10406), .C2(n6658), .A(n6657), .B(n6656), .ZN(
        P2_U3255) );
  INV_X1 U8292 ( .A(n6659), .ZN(n6897) );
  NAND2_X1 U8293 ( .A1(n8421), .A2(n10216), .ZN(n6661) );
  NAND2_X1 U8294 ( .A1(n8419), .A2(n8701), .ZN(n6660) );
  NAND2_X1 U8295 ( .A1(n6661), .A2(n6660), .ZN(n6877) );
  NAND2_X1 U8296 ( .A1(n10188), .A2(n6877), .ZN(n6664) );
  INV_X1 U8297 ( .A(n6662), .ZN(n6663) );
  OAI211_X1 U8298 ( .C1(n10199), .C2(n6897), .A(n6664), .B(n6663), .ZN(n6672)
         );
  NAND3_X1 U8299 ( .A1(n8057), .A2(n6665), .A3(n8421), .ZN(n6670) );
  OAI21_X1 U8300 ( .B1(n6667), .B2(n6666), .A(n10194), .ZN(n6669) );
  INV_X1 U8301 ( .A(n8110), .ZN(n6668) );
  AOI21_X1 U8302 ( .B1(n6670), .B2(n6669), .A(n6668), .ZN(n6671) );
  AOI211_X1 U8303 ( .C1(n8137), .C2(n6960), .A(n6672), .B(n6671), .ZN(n6673)
         );
  INV_X1 U8304 ( .A(n6673), .ZN(P2_U3223) );
  XNOR2_X1 U8305 ( .A(n6675), .B(n6674), .ZN(n6677) );
  XNOR2_X1 U8306 ( .A(n6677), .B(n6676), .ZN(n6683) );
  NAND3_X1 U8307 ( .A1(n6680), .A2(n6679), .A3(n6678), .ZN(n7598) );
  AOI22_X1 U8308 ( .A1(n9031), .A2(n6310), .B1(n7598), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n6682) );
  INV_X1 U8309 ( .A(n9026), .ZN(n9041) );
  AOI22_X1 U8310 ( .A1(n9041), .A2(n9359), .B1(n9030), .B2(n9357), .ZN(n6681)
         );
  OAI211_X1 U8311 ( .C1(n6683), .C2(n9049), .A(n6682), .B(n6681), .ZN(P1_U3220) );
  INV_X1 U8312 ( .A(n7784), .ZN(n6685) );
  OAI222_X1 U8313 ( .A1(n7510), .A2(n6684), .B1(n7595), .B2(n6685), .C1(n8517), 
        .C2(P2_U3152), .ZN(P2_U3339) );
  OAI222_X1 U8314 ( .A1(P1_U3084), .A2(n9544), .B1(n9773), .B2(n6685), .C1(
        n9907), .C2(n9774), .ZN(P1_U3334) );
  INV_X1 U8315 ( .A(n6686), .ZN(n6687) );
  AOI21_X1 U8316 ( .B1(n6689), .B2(n6688), .A(n6687), .ZN(n6693) );
  AOI22_X1 U8317 ( .A1(n9031), .A2(n6690), .B1(n7598), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n6692) );
  AOI22_X1 U8318 ( .A1(n9041), .A2(n9358), .B1(n9030), .B2(n9356), .ZN(n6691)
         );
  OAI211_X1 U8319 ( .C1(n6693), .C2(n9049), .A(n6692), .B(n6691), .ZN(P1_U3235) );
  OR2_X1 U8320 ( .A1(n6725), .A2(n6694), .ZN(n6695) );
  NAND2_X1 U8321 ( .A1(n6695), .A2(n9125), .ZN(n6696) );
  INV_X1 U8322 ( .A(n9353), .ZN(n6712) );
  NAND2_X1 U8323 ( .A1(n6712), .A2(n6707), .ZN(n9129) );
  NAND2_X1 U8324 ( .A1(n9353), .A2(n6829), .ZN(n9314) );
  NAND2_X1 U8325 ( .A1(n9129), .A2(n9314), .ZN(n9282) );
  XNOR2_X1 U8326 ( .A(n6696), .B(n9282), .ZN(n6702) );
  OAI21_X1 U8327 ( .B1(n6698), .B2(n9282), .A(n6714), .ZN(n6833) );
  NAND2_X1 U8328 ( .A1(n6833), .A2(n6699), .ZN(n6701) );
  AOI22_X1 U8329 ( .A1(n10254), .A2(n9352), .B1(n9354), .B2(n10252), .ZN(n6700) );
  OAI211_X1 U8330 ( .C1(n9620), .C2(n6702), .A(n6701), .B(n6700), .ZN(n6831)
         );
  MUX2_X1 U8331 ( .A(n6831), .B(P1_REG2_REG_6__SCAN_IN), .S(n10362), .Z(n6703)
         );
  INV_X1 U8332 ( .A(n6703), .ZN(n6711) );
  AND2_X1 U8333 ( .A1(n6704), .A2(n6707), .ZN(n6705) );
  OR2_X1 U8334 ( .A1(n6705), .A2(n6736), .ZN(n6830) );
  AOI22_X1 U8335 ( .A1(n9648), .A2(n6707), .B1(n6706), .B2(n10360), .ZN(n6708)
         );
  OAI21_X1 U8336 ( .B1(n6830), .B2(n9651), .A(n6708), .ZN(n6709) );
  AOI21_X1 U8337 ( .B1(n6833), .B2(n10344), .A(n6709), .ZN(n6710) );
  NAND2_X1 U8338 ( .A1(n6711), .A2(n6710), .ZN(P1_U3285) );
  INV_X1 U8339 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n6740) );
  NAND2_X1 U8340 ( .A1(n6712), .A2(n6829), .ZN(n6713) );
  NAND2_X1 U8341 ( .A1(n6714), .A2(n6713), .ZN(n6721) );
  INV_X1 U8342 ( .A(n9352), .ZN(n6853) );
  NAND2_X1 U8343 ( .A1(n6716), .A2(n6840), .ZN(n6719) );
  OR2_X1 U8344 ( .A1(n6409), .A2(n6717), .ZN(n6718) );
  OAI211_X1 U8345 ( .C1(n6842), .C2(n6720), .A(n6719), .B(n6718), .ZN(n6756)
         );
  NAND2_X1 U8346 ( .A1(n6853), .A2(n6756), .ZN(n9137) );
  INV_X1 U8347 ( .A(n6756), .ZN(n6980) );
  NAND2_X1 U8348 ( .A1(n9352), .A2(n6980), .ZN(n9134) );
  NAND2_X1 U8349 ( .A1(n9137), .A2(n9134), .ZN(n9280) );
  OAI21_X1 U8350 ( .B1(n6721), .B2(n9280), .A(n6855), .ZN(n6722) );
  INV_X1 U8351 ( .A(n6722), .ZN(n6986) );
  INV_X1 U8352 ( .A(n9280), .ZN(n6726) );
  AND2_X1 U8353 ( .A1(n9129), .A2(n9125), .ZN(n9312) );
  INV_X1 U8354 ( .A(n9308), .ZN(n6723) );
  NAND2_X1 U8355 ( .A1(n9129), .A2(n6723), .ZN(n6724) );
  NAND2_X1 U8356 ( .A1(n6724), .A2(n9314), .ZN(n9071) );
  NAND2_X1 U8357 ( .A1(n9136), .A2(n6726), .ZN(n6839) );
  OAI21_X1 U8358 ( .B1(n6726), .B2(n9136), .A(n6839), .ZN(n6735) );
  NAND2_X1 U8359 ( .A1(n4481), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6734) );
  INV_X1 U8360 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n6728) );
  NAND2_X1 U8361 ( .A1(n6729), .A2(n6728), .ZN(n6730) );
  AND2_X1 U8362 ( .A1(n6846), .A2(n6730), .ZN(n6953) );
  NAND2_X1 U8363 ( .A1(n7984), .A2(n6953), .ZN(n6733) );
  NAND2_X1 U8364 ( .A1(n4480), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n6732) );
  NAND2_X1 U8365 ( .A1(n9118), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6731) );
  NAND4_X1 U8366 ( .A1(n6734), .A2(n6733), .A3(n6732), .A4(n6731), .ZN(n9351)
         );
  AOI222_X1 U8367 ( .A1(n10355), .A2(n6735), .B1(n9353), .B2(n10252), .C1(
        n9351), .C2(n10254), .ZN(n6981) );
  INV_X1 U8368 ( .A(n6736), .ZN(n6737) );
  AND2_X1 U8369 ( .A1(n6736), .A2(n6980), .ZN(n6860) );
  AOI211_X1 U8370 ( .C1(n6756), .C2(n6737), .A(n10388), .B(n6860), .ZN(n6984)
         );
  AOI21_X1 U8371 ( .B1(n10372), .B2(n6756), .A(n6984), .ZN(n6738) );
  OAI211_X1 U8372 ( .C1(n9742), .C2(n6986), .A(n6981), .B(n6738), .ZN(n6741)
         );
  NAND2_X1 U8373 ( .A1(n6741), .A2(n10396), .ZN(n6739) );
  OAI21_X1 U8374 ( .B1(n10396), .B2(n6740), .A(n6739), .ZN(P1_U3475) );
  NAND2_X1 U8375 ( .A1(n6741), .A2(n4483), .ZN(n6742) );
  OAI21_X1 U8376 ( .B1(n4483), .B2(n5975), .A(n6742), .ZN(P1_U3530) );
  NAND2_X1 U8377 ( .A1(n6744), .A2(n8947), .ZN(n6746) );
  OAI21_X1 U8378 ( .B1(n6744), .B2(n8947), .A(n6743), .ZN(n6745) );
  NAND2_X1 U8379 ( .A1(n9352), .A2(n7936), .ZN(n6749) );
  NAND2_X1 U8380 ( .A1(n6756), .A2(n7961), .ZN(n6748) );
  NAND2_X1 U8381 ( .A1(n6749), .A2(n6748), .ZN(n6750) );
  XNOR2_X1 U8382 ( .A(n6750), .B(n7956), .ZN(n6921) );
  NAND2_X1 U8383 ( .A1(n9352), .A2(n7320), .ZN(n6752) );
  NAND2_X1 U8384 ( .A1(n6756), .A2(n7936), .ZN(n6751) );
  AND2_X1 U8385 ( .A1(n6752), .A2(n6751), .ZN(n6909) );
  INV_X1 U8386 ( .A(n6909), .ZN(n6913) );
  XNOR2_X1 U8387 ( .A(n6921), .B(n6913), .ZN(n6753) );
  XNOR2_X1 U8388 ( .A(n6912), .B(n6753), .ZN(n6762) );
  INV_X1 U8389 ( .A(n6754), .ZN(n6755) );
  AOI21_X1 U8390 ( .B1(n9041), .B2(n9353), .A(n6755), .ZN(n6760) );
  NAND2_X1 U8391 ( .A1(n9031), .A2(n6756), .ZN(n6759) );
  NAND2_X1 U8392 ( .A1(n9042), .A2(n6978), .ZN(n6758) );
  NAND2_X1 U8393 ( .A1(n9030), .A2(n9351), .ZN(n6757) );
  NAND4_X1 U8394 ( .A1(n6760), .A2(n6759), .A3(n6758), .A4(n6757), .ZN(n6761)
         );
  AOI21_X1 U8395 ( .B1(n6762), .B2(n8977), .A(n6761), .ZN(n6763) );
  INV_X1 U8396 ( .A(n6763), .ZN(P1_U3211) );
  INV_X1 U8397 ( .A(n6764), .ZN(n7113) );
  NAND2_X1 U8398 ( .A1(n6047), .A2(n10465), .ZN(n8253) );
  INV_X1 U8399 ( .A(n8253), .ZN(n6765) );
  NOR2_X1 U8400 ( .A1(n7113), .A2(n6765), .ZN(n10467) );
  INV_X1 U8401 ( .A(n6766), .ZN(n6768) );
  NAND2_X1 U8402 ( .A1(n6768), .A2(n6767), .ZN(n6821) );
  NAND2_X1 U8403 ( .A1(n5095), .A2(n5213), .ZN(n6787) );
  NAND2_X1 U8404 ( .A1(n10435), .A2(n6787), .ZN(n10454) );
  NAND2_X1 U8405 ( .A1(n10211), .A2(n10454), .ZN(n8717) );
  INV_X1 U8406 ( .A(n10208), .ZN(n10447) );
  OAI22_X1 U8407 ( .A1(n10467), .A2(n8637), .B1(n6041), .B2(n10427), .ZN(
        n10469) );
  AOI21_X1 U8408 ( .B1(n10447), .B2(P2_REG3_REG_0__SCAN_IN), .A(n10469), .ZN(
        n6770) );
  NOR2_X1 U8409 ( .A1(n10456), .A2(n6770), .ZN(n6771) );
  AOI21_X1 U8410 ( .B1(n10456), .B2(P2_REG2_REG_0__SCAN_IN), .A(n6771), .ZN(
        n6774) );
  NOR2_X1 U8411 ( .A1(n5212), .A2(n5213), .ZN(n10445) );
  INV_X1 U8412 ( .A(n6821), .ZN(n6772) );
  NAND2_X1 U8413 ( .A1(n6772), .A2(n8196), .ZN(n7121) );
  INV_X1 U8414 ( .A(n7121), .ZN(n7086) );
  OAI21_X1 U8415 ( .B1(n10228), .B2(n7086), .A(n7120), .ZN(n6773) );
  OAI211_X1 U8416 ( .C1(n10467), .C2(n8717), .A(n6774), .B(n6773), .ZN(
        P2_U3296) );
  INV_X1 U8417 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n6775) );
  OAI22_X1 U8418 ( .A1(n7121), .A2(n6776), .B1(n6775), .B2(n10208), .ZN(n6777)
         );
  AOI21_X1 U8419 ( .B1(n10228), .B2(n6778), .A(n6777), .ZN(n6781) );
  MUX2_X1 U8420 ( .A(n5854), .B(n6779), .S(n10211), .Z(n6780) );
  OAI211_X1 U8421 ( .C1(n6782), .C2(n8717), .A(n6781), .B(n6780), .ZN(P2_U3294) );
  OR2_X1 U8422 ( .A1(n6784), .A2(n6783), .ZN(n6785) );
  NAND2_X1 U8423 ( .A1(n6786), .A2(n6785), .ZN(n10477) );
  INV_X1 U8424 ( .A(n10477), .ZN(n6802) );
  INV_X1 U8425 ( .A(n6787), .ZN(n6788) );
  NAND2_X1 U8426 ( .A1(n10211), .A2(n6788), .ZN(n10417) );
  OAI21_X1 U8427 ( .B1(n6790), .B2(n10471), .A(n6789), .ZN(n10473) );
  OAI22_X1 U8428 ( .A1(n7121), .A2(n10473), .B1(n10208), .B2(
        P2_REG3_REG_3__SCAN_IN), .ZN(n6791) );
  AOI21_X1 U8429 ( .B1(n10228), .B2(n6792), .A(n6791), .ZN(n6801) );
  OAI21_X1 U8430 ( .B1(n8263), .B2(n6794), .A(n6793), .ZN(n6796) );
  AOI21_X1 U8431 ( .B1(n6796), .B2(n10432), .A(n6795), .ZN(n6799) );
  INV_X1 U8432 ( .A(n10435), .ZN(n6797) );
  NAND2_X1 U8433 ( .A1(n10477), .A2(n6797), .ZN(n6798) );
  AND2_X1 U8434 ( .A1(n6799), .A2(n6798), .ZN(n10474) );
  MUX2_X1 U8435 ( .A(n10474), .B(n5856), .S(n10456), .Z(n6800) );
  OAI211_X1 U8436 ( .C1(n6802), .C2(n10417), .A(n6801), .B(n6800), .ZN(
        P2_U3293) );
  OAI21_X1 U8437 ( .B1(n6804), .B2(n6803), .A(n8975), .ZN(n6811) );
  INV_X1 U8438 ( .A(n9042), .ZN(n9024) );
  AOI22_X1 U8439 ( .A1(n9041), .A2(n9357), .B1(n9030), .B2(n9355), .ZN(n6809)
         );
  INV_X1 U8440 ( .A(n6805), .ZN(n6806) );
  AOI21_X1 U8441 ( .B1(n9031), .B2(n6807), .A(n6806), .ZN(n6808) );
  OAI211_X1 U8442 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n9024), .A(n6809), .B(
        n6808), .ZN(n6810) );
  AOI21_X1 U8443 ( .B1(n6811), .B2(n8977), .A(n6810), .ZN(n6812) );
  INV_X1 U8444 ( .A(n6812), .ZN(P1_U3216) );
  OR2_X1 U8445 ( .A1(n8422), .A2(n6813), .ZN(n6814) );
  INV_X1 U8446 ( .A(n8421), .ZN(n6816) );
  OR2_X1 U8447 ( .A1(n6866), .A2(n6816), .ZN(n8284) );
  NAND2_X1 U8448 ( .A1(n6866), .A2(n6816), .ZN(n8283) );
  NAND2_X1 U8449 ( .A1(n8284), .A2(n8283), .ZN(n6874) );
  OAI21_X1 U8450 ( .B1(n6817), .B2(n6874), .A(n6868), .ZN(n10484) );
  INV_X1 U8451 ( .A(n10484), .ZN(n6828) );
  INV_X1 U8452 ( .A(n6874), .ZN(n8281) );
  XNOR2_X1 U8453 ( .A(n6875), .B(n8281), .ZN(n6819) );
  AOI222_X1 U8454 ( .A1(n10432), .A2(n6819), .B1(n8422), .B2(n10216), .C1(
        n8420), .C2(n8701), .ZN(n10481) );
  MUX2_X1 U8455 ( .A(n6820), .B(n10481), .S(n10211), .Z(n6827) );
  NOR2_X2 U8456 ( .A1(n6821), .A2(n10449), .ZN(n10422) );
  INV_X1 U8457 ( .A(n10422), .ZN(n10206) );
  OR2_X1 U8458 ( .A1(n6822), .A2(n6866), .ZN(n6873) );
  OAI211_X1 U8459 ( .C1(n6823), .C2(n10480), .A(n10418), .B(n6873), .ZN(n10479) );
  OAI22_X1 U8460 ( .A1(n10206), .A2(n10479), .B1(n6824), .B2(n10208), .ZN(
        n6825) );
  AOI21_X1 U8461 ( .B1(n10228), .B2(n6866), .A(n6825), .ZN(n6826) );
  OAI211_X1 U8462 ( .C1(n6828), .C2(n8717), .A(n6827), .B(n6826), .ZN(P2_U3289) );
  OAI22_X1 U8463 ( .A1(n6830), .A2(n10388), .B1(n6829), .B2(n10386), .ZN(n6832) );
  AOI211_X1 U8464 ( .C1(n10393), .C2(n6833), .A(n6832), .B(n6831), .ZN(n6836)
         );
  OR2_X1 U8465 ( .A1(n6836), .A2(n10399), .ZN(n6834) );
  OAI21_X1 U8466 ( .B1(n4483), .B2(n6835), .A(n6834), .ZN(P1_U3529) );
  INV_X1 U8467 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n6838) );
  OR2_X1 U8468 ( .A1(n6836), .A2(n10394), .ZN(n6837) );
  OAI21_X1 U8469 ( .B1(n10396), .B2(n6838), .A(n6837), .ZN(P1_U3472) );
  NAND2_X1 U8470 ( .A1(n6841), .A2(n6840), .ZN(n6844) );
  AOI22_X1 U8471 ( .A1(n7785), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n4614), .B2(
        n10300), .ZN(n6843) );
  NAND2_X1 U8472 ( .A1(n6929), .A2(n9351), .ZN(n10345) );
  INV_X1 U8473 ( .A(n9351), .ZN(n10353) );
  NAND2_X1 U8474 ( .A1(n10353), .A2(n7136), .ZN(n9148) );
  XNOR2_X1 U8475 ( .A(n7139), .B(n6856), .ZN(n6852) );
  NAND2_X1 U8476 ( .A1(n6846), .A2(n6845), .ZN(n6847) );
  AND2_X1 U8477 ( .A1(n6935), .A2(n6847), .ZN(n10361) );
  NAND2_X1 U8478 ( .A1(n7984), .A2(n10361), .ZN(n6851) );
  NAND2_X1 U8479 ( .A1(n4481), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6850) );
  NAND2_X1 U8480 ( .A1(n9118), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6849) );
  NAND2_X1 U8481 ( .A1(n4480), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n6848) );
  NAND4_X1 U8482 ( .A1(n6851), .A2(n6850), .A3(n6849), .A4(n6848), .ZN(n9350)
         );
  AOI222_X1 U8483 ( .A1(n10355), .A2(n6852), .B1(n9350), .B2(n10254), .C1(
        n9352), .C2(n10252), .ZN(n6890) );
  NAND2_X1 U8484 ( .A1(n6853), .A2(n6980), .ZN(n6854) );
  INV_X1 U8485 ( .A(n6856), .ZN(n9281) );
  OAI21_X1 U8486 ( .B1(n4561), .B2(n9281), .A(n7137), .ZN(n6891) );
  INV_X1 U8487 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n6858) );
  INV_X1 U8488 ( .A(n6953), .ZN(n6857) );
  OAI22_X1 U8489 ( .A1(n10366), .A2(n6858), .B1(n6857), .B2(n9555), .ZN(n6859)
         );
  AOI21_X1 U8490 ( .B1(n9648), .B2(n7136), .A(n6859), .ZN(n6863) );
  NAND2_X1 U8491 ( .A1(n6860), .A2(n6929), .ZN(n10339) );
  OR2_X1 U8492 ( .A1(n6860), .A2(n6929), .ZN(n6861) );
  AND2_X1 U8493 ( .A1(n10339), .A2(n6861), .ZN(n6888) );
  NAND2_X1 U8494 ( .A1(n6888), .A2(n10343), .ZN(n6862) );
  OAI211_X1 U8495 ( .C1(n6891), .C2(n9633), .A(n6863), .B(n6862), .ZN(n6864)
         );
  INV_X1 U8496 ( .A(n6864), .ZN(n6865) );
  OAI21_X1 U8497 ( .B1(n10362), .B2(n6890), .A(n6865), .ZN(P1_U3283) );
  OR2_X1 U8498 ( .A1(n6866), .A2(n8421), .ZN(n6867) );
  OR2_X1 U8499 ( .A1(n6960), .A2(n10430), .ZN(n8289) );
  NAND2_X1 U8500 ( .A1(n6960), .A2(n10430), .ZN(n8290) );
  NAND2_X1 U8501 ( .A1(n6870), .A2(n8286), .ZN(n6871) );
  NAND2_X1 U8502 ( .A1(n6962), .A2(n6871), .ZN(n6905) );
  INV_X1 U8503 ( .A(n6905), .ZN(n6880) );
  INV_X1 U8504 ( .A(n6872), .ZN(n10493) );
  AOI211_X1 U8505 ( .C1(n6960), .C2(n6873), .A(n10472), .B(n10420), .ZN(n6902)
         );
  OAI21_X1 U8506 ( .B1(n6876), .B2(n8286), .A(n6967), .ZN(n6878) );
  AOI21_X1 U8507 ( .B1(n6878), .B2(n10432), .A(n6877), .ZN(n6879) );
  OAI21_X1 U8508 ( .B1(n10435), .B2(n6905), .A(n6879), .ZN(n6896) );
  AOI211_X1 U8509 ( .C1(n6880), .C2(n10493), .A(n6902), .B(n6896), .ZN(n6887)
         );
  INV_X1 U8510 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n6881) );
  NOR2_X1 U8511 ( .A1(n10496), .A2(n6881), .ZN(n6882) );
  AOI21_X1 U8512 ( .B1(n8844), .B2(n6960), .A(n6882), .ZN(n6883) );
  OAI21_X1 U8513 ( .B1(n6887), .B2(n10494), .A(n6883), .ZN(P2_U3475) );
  INV_X1 U8514 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6884) );
  NOR2_X1 U8515 ( .A1(n10499), .A2(n6884), .ZN(n6885) );
  AOI21_X1 U8516 ( .B1(n8773), .B2(n6960), .A(n6885), .ZN(n6886) );
  OAI21_X1 U8517 ( .B1(n6887), .B2(n10504), .A(n6886), .ZN(P2_U3528) );
  INV_X1 U8518 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n6893) );
  AOI22_X1 U8519 ( .A1(n6888), .A2(n9721), .B1(n10372), .B2(n7136), .ZN(n6889)
         );
  OAI211_X1 U8520 ( .C1(n9742), .C2(n6891), .A(n6890), .B(n6889), .ZN(n6894)
         );
  NAND2_X1 U8521 ( .A1(n6894), .A2(n10396), .ZN(n6892) );
  OAI21_X1 U8522 ( .B1(n10396), .B2(n6893), .A(n6892), .ZN(P1_U3478) );
  NAND2_X1 U8523 ( .A1(n6894), .A2(n4483), .ZN(n6895) );
  OAI21_X1 U8524 ( .B1(n4483), .B2(n5972), .A(n6895), .ZN(P1_U3531) );
  NAND2_X1 U8525 ( .A1(n6896), .A2(n10211), .ZN(n6904) );
  OAI22_X1 U8526 ( .A1(n10211), .A2(n6898), .B1(n6897), .B2(n10208), .ZN(n6901) );
  INV_X1 U8527 ( .A(n6960), .ZN(n6899) );
  NOR2_X1 U8528 ( .A1(n10439), .A2(n6899), .ZN(n6900) );
  AOI211_X1 U8529 ( .C1(n6902), .C2(n10422), .A(n6901), .B(n6900), .ZN(n6903)
         );
  OAI211_X1 U8530 ( .C1(n6905), .C2(n10417), .A(n6904), .B(n6903), .ZN(
        P2_U3288) );
  NAND2_X1 U8531 ( .A1(n6906), .A2(n6840), .ZN(n6908) );
  AOI22_X1 U8532 ( .A1(n7785), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n4614), .B2(
        n10309), .ZN(n6907) );
  NAND2_X1 U8533 ( .A1(n6908), .A2(n6907), .ZN(n7145) );
  INV_X1 U8534 ( .A(n7145), .ZN(n10387) );
  NAND2_X1 U8535 ( .A1(n6912), .A2(n6909), .ZN(n6923) );
  OR2_X1 U8536 ( .A1(n6929), .A2(n4484), .ZN(n6911) );
  NAND2_X1 U8537 ( .A1(n9351), .A2(n7320), .ZN(n6910) );
  NAND2_X1 U8538 ( .A1(n6911), .A2(n6910), .ZN(n6924) );
  AND2_X1 U8539 ( .A1(n6923), .A2(n6924), .ZN(n6916) );
  INV_X1 U8540 ( .A(n6912), .ZN(n6914) );
  NAND2_X1 U8541 ( .A1(n6925), .A2(n6921), .ZN(n6915) );
  NAND2_X1 U8542 ( .A1(n7145), .A2(n7750), .ZN(n6918) );
  NAND2_X1 U8543 ( .A1(n9350), .A2(n7936), .ZN(n6917) );
  NAND2_X1 U8544 ( .A1(n6918), .A2(n6917), .ZN(n6919) );
  XNOR2_X1 U8545 ( .A(n6919), .B(n6589), .ZN(n6996) );
  AND2_X1 U8546 ( .A1(n9350), .A2(n7320), .ZN(n6920) );
  AOI21_X1 U8547 ( .B1(n7145), .B2(n7936), .A(n6920), .ZN(n6997) );
  XNOR2_X1 U8548 ( .A(n6996), .B(n6997), .ZN(n6931) );
  INV_X1 U8549 ( .A(n6921), .ZN(n6922) );
  NAND2_X1 U8550 ( .A1(n6923), .A2(n6922), .ZN(n6927) );
  INV_X1 U8551 ( .A(n6924), .ZN(n6926) );
  NAND3_X1 U8552 ( .A1(n6927), .A2(n6926), .A3(n6925), .ZN(n6948) );
  NAND2_X1 U8553 ( .A1(n9351), .A2(n7936), .ZN(n6928) );
  OAI21_X1 U8554 ( .B1(n6929), .B2(n7891), .A(n6928), .ZN(n6930) );
  XNOR2_X1 U8555 ( .A(n6930), .B(n6589), .ZN(n6947) );
  INV_X1 U8556 ( .A(n7000), .ZN(n6933) );
  AOI21_X1 U8557 ( .B1(n6946), .B2(n6950), .A(n6931), .ZN(n6932) );
  OAI21_X1 U8558 ( .B1(n6933), .B2(n6932), .A(n8977), .ZN(n6944) );
  NAND2_X1 U8559 ( .A1(n4481), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6940) );
  NAND2_X1 U8560 ( .A1(n6935), .A2(n6934), .ZN(n6936) );
  AND2_X1 U8561 ( .A1(n7017), .A2(n6936), .ZN(n7148) );
  NAND2_X1 U8562 ( .A1(n7984), .A2(n7148), .ZN(n6939) );
  NAND2_X1 U8563 ( .A1(n4480), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n6938) );
  NAND2_X1 U8564 ( .A1(n9118), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6937) );
  NAND4_X1 U8565 ( .A1(n6940), .A2(n6939), .A3(n6938), .A4(n6937), .ZN(n9349)
         );
  INV_X1 U8566 ( .A(n9030), .ZN(n9045) );
  AND2_X1 U8567 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n10308) );
  AOI21_X1 U8568 ( .B1(n9041), .B2(n9351), .A(n10308), .ZN(n6941) );
  OAI21_X1 U8569 ( .B1(n10351), .B2(n9045), .A(n6941), .ZN(n6942) );
  AOI21_X1 U8570 ( .B1(n10361), .B2(n9042), .A(n6942), .ZN(n6943) );
  OAI211_X1 U8571 ( .C1(n10387), .C2(n9019), .A(n6944), .B(n6943), .ZN(
        P1_U3229) );
  INV_X1 U8572 ( .A(n7802), .ZN(n6987) );
  OAI222_X1 U8573 ( .A1(n6945), .A2(P1_U3084), .B1(n9773), .B2(n6987), .C1(
        n10077), .C2(n9774), .ZN(P1_U3333) );
  INV_X1 U8574 ( .A(n6946), .ZN(n6951) );
  AOI21_X1 U8575 ( .B1(n6950), .B2(n6948), .A(n6947), .ZN(n6949) );
  AOI211_X1 U8576 ( .C1(n6951), .C2(n6950), .A(n9049), .B(n6949), .ZN(n6959)
         );
  NAND2_X1 U8577 ( .A1(P1_U3084), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n10306) );
  INV_X1 U8578 ( .A(n10306), .ZN(n6952) );
  AOI21_X1 U8579 ( .B1(n9041), .B2(n9352), .A(n6952), .ZN(n6957) );
  NAND2_X1 U8580 ( .A1(n9031), .A2(n7136), .ZN(n6956) );
  NAND2_X1 U8581 ( .A1(n9042), .A2(n6953), .ZN(n6955) );
  NAND2_X1 U8582 ( .A1(n9030), .A2(n9350), .ZN(n6954) );
  NAND4_X1 U8583 ( .A1(n6957), .A2(n6956), .A3(n6955), .A4(n6954), .ZN(n6958)
         );
  OR2_X1 U8584 ( .A1(n6959), .A2(n6958), .ZN(P1_U3219) );
  NAND2_X1 U8585 ( .A1(n6960), .A2(n8420), .ZN(n6961) );
  NAND2_X1 U8586 ( .A1(n6962), .A2(n6961), .ZN(n10416) );
  INV_X1 U8587 ( .A(n10416), .ZN(n6963) );
  INV_X1 U8588 ( .A(n8419), .ZN(n6968) );
  OR2_X1 U8589 ( .A1(n8116), .A2(n6968), .ZN(n8294) );
  NAND2_X1 U8590 ( .A1(n8116), .A2(n6968), .ZN(n8292) );
  NAND2_X1 U8591 ( .A1(n6963), .A2(n5063), .ZN(n10414) );
  OR2_X1 U8592 ( .A1(n8116), .A2(n8419), .ZN(n6964) );
  INV_X1 U8593 ( .A(n8418), .ZN(n10428) );
  NAND2_X1 U8594 ( .A1(n7157), .A2(n10428), .ZN(n8244) );
  NAND2_X1 U8595 ( .A1(n8295), .A2(n8244), .ZN(n8297) );
  NAND2_X1 U8596 ( .A1(n6965), .A2(n5065), .ZN(n6966) );
  NAND2_X1 U8597 ( .A1(n7159), .A2(n6966), .ZN(n7127) );
  XNOR2_X1 U8598 ( .A(n7164), .B(n5065), .ZN(n6970) );
  INV_X1 U8599 ( .A(n8417), .ZN(n7160) );
  INV_X1 U8600 ( .A(n10216), .ZN(n10429) );
  OAI22_X1 U8601 ( .A1(n7160), .A2(n10427), .B1(n6968), .B2(n10429), .ZN(n6969) );
  AOI21_X1 U8602 ( .B1(n6970), .B2(n10432), .A(n6969), .ZN(n6971) );
  OAI21_X1 U8603 ( .B1(n7127), .B2(n10435), .A(n6971), .ZN(n7128) );
  NAND2_X1 U8604 ( .A1(n7128), .A2(n10211), .ZN(n6977) );
  INV_X1 U8605 ( .A(n8116), .ZN(n10489) );
  AOI21_X1 U8606 ( .B1(n10419), .B2(n7157), .A(n10472), .ZN(n6972) );
  AND2_X1 U8607 ( .A1(n6972), .A2(n7161), .ZN(n7129) );
  NAND2_X1 U8608 ( .A1(n10456), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6974) );
  NAND2_X1 U8609 ( .A1(n10447), .A2(n7058), .ZN(n6973) );
  OAI211_X1 U8610 ( .C1(n10439), .C2(n4871), .A(n6974), .B(n6973), .ZN(n6975)
         );
  AOI21_X1 U8611 ( .B1(n10422), .B2(n7129), .A(n6975), .ZN(n6976) );
  OAI211_X1 U8612 ( .C1(n7127), .C2(n10417), .A(n6977), .B(n6976), .ZN(
        P2_U3286) );
  AOI22_X1 U8613 ( .A1(n10362), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n6978), .B2(
        n10360), .ZN(n6979) );
  OAI21_X1 U8614 ( .B1(n10364), .B2(n6980), .A(n6979), .ZN(n6983) );
  NOR2_X1 U8615 ( .A1(n6981), .A2(n10362), .ZN(n6982) );
  AOI211_X1 U8616 ( .C1(n6984), .C2(n9626), .A(n6983), .B(n6982), .ZN(n6985)
         );
  OAI21_X1 U8617 ( .B1(n6986), .B2(n9633), .A(n6985), .ZN(P1_U3284) );
  OAI222_X1 U8618 ( .A1(n7510), .A2(n6988), .B1(P2_U3152), .B2(n5213), .C1(
        n8872), .C2(n6987), .ZN(P2_U3338) );
  AOI22_X1 U8619 ( .A1(n10362), .A2(P1_REG2_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n10360), .ZN(n6989) );
  OAI21_X1 U8620 ( .B1(n10364), .B2(n9076), .A(n6989), .ZN(n6992) );
  NOR2_X1 U8621 ( .A1(n6990), .A2(n7154), .ZN(n6991) );
  AOI211_X1 U8622 ( .C1(n6993), .C2(n10343), .A(n6992), .B(n6991), .ZN(n6994)
         );
  OAI21_X1 U8623 ( .B1(n6995), .B2(n10362), .A(n6994), .ZN(P1_U3289) );
  INV_X1 U8624 ( .A(n6996), .ZN(n6998) );
  NAND2_X1 U8625 ( .A1(n6998), .A2(n6997), .ZN(n6999) );
  NAND2_X1 U8626 ( .A1(n7001), .A2(n6840), .ZN(n7004) );
  AOI22_X1 U8627 ( .A1(n7785), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n4614), .B2(
        n7002), .ZN(n7003) );
  NAND2_X1 U8628 ( .A1(n7183), .A2(n7961), .ZN(n7006) );
  NAND2_X1 U8629 ( .A1(n9349), .A2(n7936), .ZN(n7005) );
  NAND2_X1 U8630 ( .A1(n7006), .A2(n7005), .ZN(n7007) );
  XNOR2_X1 U8631 ( .A(n7007), .B(n6589), .ZN(n7010) );
  NAND2_X1 U8632 ( .A1(n7183), .A2(n7936), .ZN(n7009) );
  NAND2_X1 U8633 ( .A1(n9349), .A2(n7320), .ZN(n7008) );
  NAND2_X1 U8634 ( .A1(n7009), .A2(n7008), .ZN(n7011) );
  NAND2_X1 U8635 ( .A1(n7010), .A2(n7011), .ZN(n7266) );
  INV_X1 U8636 ( .A(n7010), .ZN(n7013) );
  INV_X1 U8637 ( .A(n7011), .ZN(n7012) );
  NAND2_X1 U8638 ( .A1(n7013), .A2(n7012), .ZN(n7268) );
  NAND2_X1 U8639 ( .A1(n7266), .A2(n7268), .ZN(n7014) );
  XNOR2_X1 U8640 ( .A(n7267), .B(n7014), .ZN(n7028) );
  INV_X1 U8641 ( .A(n9350), .ZN(n7141) );
  NAND2_X1 U8642 ( .A1(n4481), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n7022) );
  INV_X1 U8643 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n7016) );
  NAND2_X1 U8644 ( .A1(n7017), .A2(n7016), .ZN(n7018) );
  AND2_X1 U8645 ( .A1(n7192), .A2(n7018), .ZN(n7274) );
  NAND2_X1 U8646 ( .A1(n7984), .A2(n7274), .ZN(n7021) );
  NAND2_X1 U8647 ( .A1(n4480), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n7020) );
  NAND2_X1 U8648 ( .A1(n9118), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n7019) );
  NAND4_X1 U8649 ( .A1(n7022), .A2(n7021), .A3(n7020), .A4(n7019), .ZN(n9348)
         );
  AOI21_X1 U8650 ( .B1(n9030), .B2(n9348), .A(n7023), .ZN(n7025) );
  NAND2_X1 U8651 ( .A1(n9042), .A2(n7148), .ZN(n7024) );
  OAI211_X1 U8652 ( .C1(n7141), .C2(n9026), .A(n7025), .B(n7024), .ZN(n7026)
         );
  AOI21_X1 U8653 ( .B1(n7183), .B2(n9031), .A(n7026), .ZN(n7027) );
  OAI21_X1 U8654 ( .B1(n7028), .B2(n9049), .A(n7027), .ZN(P1_U3215) );
  NAND2_X1 U8655 ( .A1(n7036), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n7030) );
  NAND2_X1 U8656 ( .A1(n7030), .A2(n7029), .ZN(n7032) );
  INV_X1 U8657 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n8720) );
  MUX2_X1 U8658 ( .A(n8720), .B(P2_REG2_REG_11__SCAN_IN), .S(n7217), .Z(n7031)
         );
  NOR2_X1 U8659 ( .A1(n7032), .A2(n7031), .ZN(n7210) );
  AOI21_X1 U8660 ( .B1(n7032), .B2(n7031), .A(n7210), .ZN(n7044) );
  INV_X1 U8661 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n10066) );
  NOR2_X1 U8662 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10066), .ZN(n7033) );
  AOI21_X1 U8663 ( .B1(n10404), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n7033), .ZN(
        n7041) );
  INV_X1 U8664 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n7034) );
  MUX2_X1 U8665 ( .A(n7034), .B(P2_REG1_REG_11__SCAN_IN), .S(n7217), .Z(n7038)
         );
  AOI21_X1 U8666 ( .B1(n7036), .B2(P2_REG1_REG_10__SCAN_IN), .A(n7035), .ZN(
        n7037) );
  NOR2_X1 U8667 ( .A1(n7037), .A2(n7038), .ZN(n7216) );
  AOI21_X1 U8668 ( .B1(n7038), .B2(n7037), .A(n7216), .ZN(n7039) );
  NAND2_X1 U8669 ( .A1(n10402), .A2(n7039), .ZN(n7040) );
  OAI211_X1 U8670 ( .C1(n10406), .C2(n7211), .A(n7041), .B(n7040), .ZN(n7042)
         );
  INV_X1 U8671 ( .A(n7042), .ZN(n7043) );
  OAI21_X1 U8672 ( .B1(n7044), .B2(n10405), .A(n7043), .ZN(P2_U3256) );
  NAND2_X1 U8673 ( .A1(P1_U3084), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n8890) );
  INV_X1 U8674 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n7045) );
  MUX2_X1 U8675 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n7045), .S(n7411), .Z(n7048)
         );
  OAI21_X1 U8676 ( .B1(n7373), .B2(P1_REG1_REG_13__SCAN_IN), .A(n7046), .ZN(
        n7047) );
  NAND2_X1 U8677 ( .A1(n7048), .A2(n7047), .ZN(n7253) );
  OAI21_X1 U8678 ( .B1(n7048), .B2(n7047), .A(n7253), .ZN(n7049) );
  NAND2_X1 U8679 ( .A1(n7049), .A2(n10332), .ZN(n7050) );
  OAI211_X1 U8680 ( .C1(n7444), .C2(n7249), .A(n8890), .B(n7050), .ZN(n7056)
         );
  INV_X1 U8681 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7054) );
  INV_X1 U8682 ( .A(n7248), .ZN(n7052) );
  AOI211_X1 U8683 ( .C1(n7054), .C2(n7053), .A(n7052), .B(n9385), .ZN(n7055)
         );
  AOI211_X1 U8684 ( .C1(n10299), .C2(P1_ADDR_REG_14__SCAN_IN), .A(n7056), .B(
        n7055), .ZN(n7057) );
  INV_X1 U8685 ( .A(n7057), .ZN(P1_U3255) );
  INV_X1 U8686 ( .A(n7058), .ZN(n7062) );
  INV_X1 U8687 ( .A(n8160), .ZN(n8119) );
  AOI22_X1 U8688 ( .A1(n7611), .A2(n8417), .B1(n8119), .B2(n8419), .ZN(n7061)
         );
  INV_X1 U8689 ( .A(n7059), .ZN(n7060) );
  OAI211_X1 U8690 ( .C1(n7062), .C2(n10199), .A(n7061), .B(n7060), .ZN(n7066)
         );
  AOI211_X1 U8691 ( .C1(n7064), .C2(n7063), .A(n8156), .B(n7105), .ZN(n7065)
         );
  AOI211_X1 U8692 ( .C1(n8137), .C2(n7157), .A(n7066), .B(n7065), .ZN(n7067)
         );
  INV_X1 U8693 ( .A(n7067), .ZN(P2_U3219) );
  INV_X1 U8694 ( .A(n7068), .ZN(n7106) );
  NOR3_X1 U8695 ( .A1(n7069), .A2(n8142), .A3(n7160), .ZN(n7070) );
  AOI21_X1 U8696 ( .B1(n7106), .B2(n10194), .A(n7070), .ZN(n7082) );
  INV_X1 U8697 ( .A(n7071), .ZN(n7079) );
  INV_X1 U8698 ( .A(n7233), .ZN(n7077) );
  NAND2_X1 U8699 ( .A1(n8417), .A2(n10216), .ZN(n7073) );
  NAND2_X1 U8700 ( .A1(n8416), .A2(n8701), .ZN(n7072) );
  AND2_X1 U8701 ( .A1(n7073), .A2(n7072), .ZN(n7231) );
  INV_X1 U8702 ( .A(n7231), .ZN(n7074) );
  AOI22_X1 U8703 ( .A1(n10188), .A2(n7074), .B1(P2_REG3_REG_12__SCAN_IN), .B2(
        P2_U3152), .ZN(n7076) );
  NAND2_X1 U8704 ( .A1(n8137), .A2(n7395), .ZN(n7075) );
  OAI211_X1 U8705 ( .C1(n10199), .C2(n7077), .A(n7076), .B(n7075), .ZN(n7078)
         );
  AOI21_X1 U8706 ( .B1(n7079), .B2(n10194), .A(n7078), .ZN(n7080) );
  OAI21_X1 U8707 ( .B1(n7082), .B2(n7081), .A(n7080), .ZN(P2_U3226) );
  OAI22_X1 U8708 ( .A1(n5850), .A2(n10211), .B1(n7083), .B2(n10208), .ZN(n7084) );
  AOI21_X1 U8709 ( .B1(n7086), .B2(n7085), .A(n7084), .ZN(n7087) );
  OAI21_X1 U8710 ( .B1(n7088), .B2(n10439), .A(n7087), .ZN(n7089) );
  AOI21_X1 U8711 ( .B1(n8723), .B2(n7090), .A(n7089), .ZN(n7091) );
  OAI21_X1 U8712 ( .B1(n10456), .B2(n7092), .A(n7091), .ZN(P2_U3292) );
  AOI22_X1 U8713 ( .A1(n7093), .A2(n10422), .B1(n7604), .B2(n10447), .ZN(n7094) );
  OAI21_X1 U8714 ( .B1(n7607), .B2(n10439), .A(n7094), .ZN(n7097) );
  MUX2_X1 U8715 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n7095), .S(n10211), .Z(n7096)
         );
  AOI211_X1 U8716 ( .C1(n8723), .C2(n7098), .A(n7097), .B(n7096), .ZN(n7099)
         );
  INV_X1 U8717 ( .A(n7099), .ZN(P2_U3290) );
  INV_X1 U8718 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7100) );
  INV_X1 U8719 ( .A(n7821), .ZN(n7996) );
  OAI222_X1 U8720 ( .A1(n7510), .A2(n7100), .B1(P2_U3152), .B2(n8395), .C1(
        n7595), .C2(n7996), .ZN(P2_U3337) );
  AOI22_X1 U8721 ( .A1(n10216), .A2(n8418), .B1(n10217), .B2(n8701), .ZN(n7165) );
  INV_X1 U8722 ( .A(n7165), .ZN(n7101) );
  AOI22_X1 U8723 ( .A1(n10188), .A2(n7101), .B1(P2_REG3_REG_11__SCAN_IN), .B2(
        P2_U3152), .ZN(n7102) );
  OAI21_X1 U8724 ( .B1(n8719), .B2(n10199), .A(n7102), .ZN(n7110) );
  NAND3_X1 U8725 ( .A1(n8057), .A2(n7103), .A3(n8418), .ZN(n7108) );
  OAI21_X1 U8726 ( .B1(n7105), .B2(n7104), .A(n10194), .ZN(n7107) );
  AOI21_X1 U8727 ( .B1(n7108), .B2(n7107), .A(n7106), .ZN(n7109) );
  AOI211_X1 U8728 ( .C1(n8137), .C2(n8722), .A(n7110), .B(n7109), .ZN(n7111)
         );
  INV_X1 U8729 ( .A(n7111), .ZN(P2_U3238) );
  INV_X1 U8730 ( .A(n6048), .ZN(n7115) );
  NAND2_X1 U8731 ( .A1(n7112), .A2(n7113), .ZN(n7114) );
  OAI211_X1 U8732 ( .C1(n8250), .C2(n7115), .A(n7114), .B(n10432), .ZN(n7119)
         );
  NAND2_X1 U8733 ( .A1(n6047), .A2(n10216), .ZN(n7117) );
  NAND2_X1 U8734 ( .A1(n6179), .A2(n8701), .ZN(n7116) );
  NAND2_X1 U8735 ( .A1(n7117), .A2(n7116), .ZN(n7687) );
  INV_X1 U8736 ( .A(n7687), .ZN(n7118) );
  NAND2_X1 U8737 ( .A1(n7119), .A2(n7118), .ZN(n7694) );
  NOR2_X1 U8739 ( .A1(n10211), .A2(n5851), .ZN(n7123) );
  XNOR2_X1 U8740 ( .A(n6042), .B(n7120), .ZN(n7693) );
  OAI22_X1 U8741 ( .A1(n7121), .A2(n7693), .B1(n7685), .B2(n10208), .ZN(n7122)
         );
  AOI211_X1 U8742 ( .C1(n10211), .C2(n7694), .A(n7123), .B(n7122), .ZN(n7126)
         );
  OAI21_X1 U8743 ( .B1(n7112), .B2(n6043), .A(n7124), .ZN(n7696) );
  AOI22_X1 U8744 ( .A1(n8723), .A2(n7696), .B1(n10228), .B2(n6042), .ZN(n7125)
         );
  NAND2_X1 U8745 ( .A1(n7126), .A2(n7125), .ZN(P2_U3295) );
  INV_X1 U8746 ( .A(n7127), .ZN(n7130) );
  AOI211_X1 U8747 ( .C1(n7130), .C2(n10493), .A(n7129), .B(n7128), .ZN(n7135)
         );
  AOI22_X1 U8748 ( .A1(n8773), .A2(n7157), .B1(n10504), .B2(
        P2_REG1_REG_10__SCAN_IN), .ZN(n7131) );
  OAI21_X1 U8749 ( .B1(n7135), .B2(n10504), .A(n7131), .ZN(P2_U3530) );
  INV_X1 U8750 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n7132) );
  NOR2_X1 U8751 ( .A1(n10496), .A2(n7132), .ZN(n7133) );
  AOI21_X1 U8752 ( .B1(n8844), .B2(n7157), .A(n7133), .ZN(n7134) );
  OAI21_X1 U8753 ( .B1(n7135), .B2(n10494), .A(n7134), .ZN(P2_U3481) );
  AND2_X1 U8754 ( .A1(n7145), .A2(n9350), .ZN(n7138) );
  NAND2_X1 U8755 ( .A1(n7183), .A2(n10351), .ZN(n9146) );
  NAND2_X1 U8756 ( .A1(n9144), .A2(n9146), .ZN(n7181) );
  INV_X1 U8757 ( .A(n7181), .ZN(n9286) );
  XNOR2_X1 U8758 ( .A(n7182), .B(n9286), .ZN(n10179) );
  INV_X1 U8759 ( .A(n9148), .ZN(n9140) );
  NAND2_X1 U8760 ( .A1(n10387), .A2(n9350), .ZN(n9284) );
  NAND2_X1 U8761 ( .A1(n9284), .A2(n10345), .ZN(n9147) );
  NAND2_X1 U8762 ( .A1(n7145), .A2(n7141), .ZN(n9285) );
  INV_X1 U8763 ( .A(n9285), .ZN(n9141) );
  NOR2_X1 U8764 ( .A1(n4559), .A2(n9141), .ZN(n7140) );
  XNOR2_X1 U8765 ( .A(n7140), .B(n7181), .ZN(n7143) );
  INV_X1 U8766 ( .A(n9348), .ZN(n7187) );
  OAI22_X1 U8767 ( .A1(n7141), .A2(n10352), .B1(n7187), .B2(n10350), .ZN(n7142) );
  AOI21_X1 U8768 ( .B1(n7143), .B2(n10355), .A(n7142), .ZN(n7144) );
  OAI21_X1 U8769 ( .B1(n10179), .B2(n10358), .A(n7144), .ZN(n10182) );
  NAND2_X1 U8770 ( .A1(n10182), .A2(n10366), .ZN(n7153) );
  INV_X1 U8771 ( .A(n7183), .ZN(n10181) );
  INV_X1 U8772 ( .A(n10340), .ZN(n7147) );
  INV_X1 U8773 ( .A(n7202), .ZN(n7146) );
  OAI211_X1 U8774 ( .C1(n10181), .C2(n7147), .A(n7146), .B(n9721), .ZN(n10180)
         );
  INV_X1 U8775 ( .A(n10180), .ZN(n7151) );
  AOI22_X1 U8776 ( .A1(n10362), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n7148), .B2(
        n10360), .ZN(n7149) );
  OAI21_X1 U8777 ( .B1(n10181), .B2(n10364), .A(n7149), .ZN(n7150) );
  AOI21_X1 U8778 ( .B1(n7151), .B2(n9626), .A(n7150), .ZN(n7152) );
  OAI211_X1 U8779 ( .C1(n10179), .C2(n7154), .A(n7153), .B(n7152), .ZN(
        P1_U3281) );
  INV_X1 U8780 ( .A(n7841), .ZN(n7155) );
  OAI222_X1 U8781 ( .A1(P1_U3084), .A2(n9263), .B1(n9773), .B2(n7155), .C1(
        n7842), .C2(n9774), .ZN(P1_U3331) );
  OAI222_X1 U8782 ( .A1(n7510), .A2(n7156), .B1(n7595), .B2(n7155), .C1(n4486), 
        .C2(P2_U3152), .ZN(P2_U3336) );
  NAND2_X1 U8783 ( .A1(n7157), .A2(n8418), .ZN(n7158) );
  OR2_X1 U8784 ( .A1(n8722), .A2(n7160), .ZN(n8306) );
  NAND2_X1 U8785 ( .A1(n8722), .A2(n7160), .ZN(n8243) );
  XNOR2_X1 U8786 ( .A(n7240), .B(n8207), .ZN(n8724) );
  NAND2_X1 U8787 ( .A1(n7161), .A2(n8722), .ZN(n7162) );
  NAND2_X1 U8788 ( .A1(n7162), .A2(n10418), .ZN(n7163) );
  NOR2_X1 U8789 ( .A1(n7234), .A2(n7163), .ZN(n8725) );
  INV_X1 U8790 ( .A(n8207), .ZN(n7239) );
  XNOR2_X1 U8791 ( .A(n7229), .B(n7239), .ZN(n7166) );
  OAI21_X1 U8792 ( .B1(n7166), .B2(n8637), .A(n7165), .ZN(n8718) );
  AOI211_X1 U8793 ( .C1(n8724), .C2(n10485), .A(n8725), .B(n8718), .ZN(n7171)
         );
  INV_X1 U8794 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n7167) );
  NOR2_X1 U8795 ( .A1(n10496), .A2(n7167), .ZN(n7168) );
  AOI21_X1 U8796 ( .B1(n8844), .B2(n8722), .A(n7168), .ZN(n7169) );
  OAI21_X1 U8797 ( .B1(n7171), .B2(n10494), .A(n7169), .ZN(P2_U3484) );
  AOI22_X1 U8798 ( .A1(n8773), .A2(n8722), .B1(n10504), .B2(
        P2_REG1_REG_11__SCAN_IN), .ZN(n7170) );
  OAI21_X1 U8799 ( .B1(n7171), .B2(n10504), .A(n7170), .ZN(P2_U3531) );
  OAI211_X1 U8800 ( .C1(n7173), .C2(n4564), .A(n7172), .B(n10194), .ZN(n7178)
         );
  INV_X1 U8801 ( .A(n7174), .ZN(n10209) );
  OAI22_X1 U8802 ( .A1(n10199), .A2(n10209), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7222), .ZN(n7176) );
  INV_X1 U8803 ( .A(n10217), .ZN(n7228) );
  INV_X1 U8804 ( .A(n10218), .ZN(n7475) );
  OAI22_X1 U8805 ( .A1(n7228), .A2(n8160), .B1(n8161), .B2(n7475), .ZN(n7175)
         );
  AOI211_X1 U8806 ( .C1(n8137), .C2(n10227), .A(n7176), .B(n7175), .ZN(n7177)
         );
  NAND2_X1 U8807 ( .A1(n7178), .A2(n7177), .ZN(P2_U3236) );
  INV_X1 U8808 ( .A(n7858), .ZN(n7180) );
  NAND2_X1 U8809 ( .A1(n8869), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n7179) );
  OAI211_X1 U8810 ( .C1(n7180), .C2(n8872), .A(n8405), .B(n7179), .ZN(P2_U3335) );
  NAND2_X1 U8811 ( .A1(n7184), .A2(n6840), .ZN(n7186) );
  AOI22_X1 U8812 ( .A1(n7785), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n4614), .B2(
        n10323), .ZN(n7185) );
  OR2_X1 U8813 ( .A1(n7300), .A2(n7187), .ZN(n7416) );
  NAND2_X1 U8814 ( .A1(n7300), .A2(n7187), .ZN(n9094) );
  NAND2_X1 U8815 ( .A1(n7188), .A2(n9287), .ZN(n7189) );
  NAND2_X1 U8816 ( .A1(n7302), .A2(n7189), .ZN(n7201) );
  NAND2_X1 U8817 ( .A1(n9146), .A2(n9285), .ZN(n9150) );
  INV_X1 U8818 ( .A(n9287), .ZN(n9154) );
  XNOR2_X1 U8819 ( .A(n7281), .B(n9154), .ZN(n7199) );
  NAND2_X1 U8820 ( .A1(n4481), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n7197) );
  INV_X1 U8821 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n7191) );
  NAND2_X1 U8822 ( .A1(n7192), .A2(n7191), .ZN(n7193) );
  AND2_X1 U8823 ( .A1(n7289), .A2(n7193), .ZN(n7331) );
  NAND2_X1 U8824 ( .A1(n7984), .A2(n7331), .ZN(n7196) );
  NAND2_X1 U8825 ( .A1(n4480), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n7195) );
  NAND2_X1 U8826 ( .A1(n9118), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n7194) );
  NAND4_X1 U8827 ( .A1(n7197), .A2(n7196), .A3(n7195), .A4(n7194), .ZN(n10253)
         );
  INV_X1 U8828 ( .A(n10253), .ZN(n7286) );
  OAI22_X1 U8829 ( .A1(n10351), .A2(n10352), .B1(n7286), .B2(n10350), .ZN(
        n7198) );
  AOI21_X1 U8830 ( .B1(n7199), .B2(n10355), .A(n7198), .ZN(n7200) );
  OAI21_X1 U8831 ( .B1(n7201), .B2(n10358), .A(n7200), .ZN(n10283) );
  INV_X1 U8832 ( .A(n10283), .ZN(n7208) );
  INV_X1 U8833 ( .A(n7201), .ZN(n10285) );
  INV_X1 U8834 ( .A(n7300), .ZN(n10281) );
  NOR2_X1 U8835 ( .A1(n7202), .A2(n10281), .ZN(n7203) );
  OR2_X1 U8836 ( .A1(n7296), .A2(n7203), .ZN(n10282) );
  AOI22_X1 U8837 ( .A1(n10362), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n7274), .B2(
        n10360), .ZN(n7205) );
  NAND2_X1 U8838 ( .A1(n7300), .A2(n9648), .ZN(n7204) );
  OAI211_X1 U8839 ( .C1(n10282), .C2(n9651), .A(n7205), .B(n7204), .ZN(n7206)
         );
  AOI21_X1 U8840 ( .B1(n10285), .B2(n10344), .A(n7206), .ZN(n7207) );
  OAI21_X1 U8841 ( .B1(n7208), .B2(n10362), .A(n7207), .ZN(P1_U3280) );
  NAND2_X1 U8842 ( .A1(n8440), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n7212) );
  MUX2_X1 U8843 ( .A(n7237), .B(P2_REG2_REG_12__SCAN_IN), .S(n8440), .Z(n7209)
         );
  INV_X1 U8844 ( .A(n7209), .ZN(n8442) );
  AOI21_X1 U8845 ( .B1(n7211), .B2(n8720), .A(n7210), .ZN(n8443) );
  NAND2_X1 U8846 ( .A1(n8442), .A2(n8443), .ZN(n8441) );
  NAND2_X1 U8847 ( .A1(n7212), .A2(n8441), .ZN(n7214) );
  AOI22_X1 U8848 ( .A1(n7353), .A2(n10210), .B1(P2_REG2_REG_13__SCAN_IN), .B2(
        n7215), .ZN(n7213) );
  NOR2_X1 U8849 ( .A1(n7214), .A2(n7213), .ZN(n7348) );
  AOI21_X1 U8850 ( .B1(n7214), .B2(n7213), .A(n7348), .ZN(n7227) );
  INV_X1 U8851 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n10238) );
  AOI22_X1 U8852 ( .A1(n7353), .A2(P2_REG1_REG_13__SCAN_IN), .B1(n10238), .B2(
        n7215), .ZN(n7220) );
  INV_X1 U8853 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7218) );
  MUX2_X1 U8854 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n7218), .S(n8440), .Z(n8447)
         );
  OAI21_X1 U8855 ( .B1(n7220), .B2(n7219), .A(n7352), .ZN(n7221) );
  NAND2_X1 U8856 ( .A1(n7221), .A2(n10402), .ZN(n7226) );
  INV_X1 U8857 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n7223) );
  OAI22_X1 U8858 ( .A1(n7359), .A2(n7223), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7222), .ZN(n7224) );
  AOI21_X1 U8859 ( .B1(n8491), .B2(n7353), .A(n7224), .ZN(n7225) );
  OAI211_X1 U8860 ( .C1(n7227), .C2(n10405), .A(n7226), .B(n7225), .ZN(
        P2_U3258) );
  NAND2_X1 U8861 ( .A1(n7395), .A2(n7228), .ZN(n8309) );
  NAND2_X1 U8862 ( .A1(n7397), .A2(n8243), .ZN(n7230) );
  XOR2_X1 U8863 ( .A(n8208), .B(n7230), .Z(n7232) );
  OAI21_X1 U8864 ( .B1(n7232), .B2(n8637), .A(n7231), .ZN(n7308) );
  AOI21_X1 U8865 ( .B1(n7233), .B2(n10447), .A(n7308), .ZN(n7245) );
  INV_X1 U8866 ( .A(n7234), .ZN(n7236) );
  INV_X1 U8867 ( .A(n7395), .ZN(n7312) );
  NAND2_X1 U8868 ( .A1(n7234), .A2(n7312), .ZN(n10204) );
  INV_X1 U8869 ( .A(n10204), .ZN(n7235) );
  AOI211_X1 U8870 ( .C1(n7395), .C2(n7236), .A(n10472), .B(n7235), .ZN(n7309)
         );
  OAI22_X1 U8871 ( .A1(n10439), .A2(n7312), .B1(n7237), .B2(n10211), .ZN(n7238) );
  AOI21_X1 U8872 ( .B1(n7309), .B2(n10422), .A(n7238), .ZN(n7244) );
  NAND2_X1 U8873 ( .A1(n7240), .A2(n7239), .ZN(n7242) );
  NAND2_X1 U8874 ( .A1(n8722), .A2(n8417), .ZN(n7241) );
  XNOR2_X1 U8875 ( .A(n7396), .B(n8208), .ZN(n7310) );
  NAND2_X1 U8876 ( .A1(n7310), .A2(n8723), .ZN(n7243) );
  OAI211_X1 U8877 ( .C1(n7245), .C2(n10456), .A(n7244), .B(n7243), .ZN(
        P2_U3284) );
  NAND2_X1 U8878 ( .A1(n7858), .A2(n9768), .ZN(n7247) );
  OR2_X1 U8879 ( .A1(n7246), .A2(P1_U3084), .ZN(n9340) );
  OAI211_X1 U8880 ( .C1(n7859), .C2(n9774), .A(n7247), .B(n9340), .ZN(P1_U3330) );
  INV_X1 U8881 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n7252) );
  OAI21_X1 U8882 ( .B1(n7250), .B2(n7249), .A(n7248), .ZN(n7438) );
  XNOR2_X1 U8883 ( .A(n7438), .B(n7714), .ZN(n7251) );
  NOR2_X1 U8884 ( .A1(n7251), .A2(n7252), .ZN(n7437) );
  AOI211_X1 U8885 ( .C1(n7252), .C2(n7251), .A(n9385), .B(n7437), .ZN(n7261)
         );
  INV_X1 U8886 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n7256) );
  OAI21_X1 U8887 ( .B1(n7411), .B2(P1_REG1_REG_14__SCAN_IN), .A(n7253), .ZN(
        n7432) );
  XNOR2_X1 U8888 ( .A(n7432), .B(n7714), .ZN(n7254) );
  INV_X1 U8889 ( .A(n7254), .ZN(n7255) );
  AND2_X1 U8890 ( .A1(n7254), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n7433) );
  AOI211_X1 U8891 ( .C1(n7256), .C2(n7255), .A(n9367), .B(n7433), .ZN(n7260)
         );
  INV_X1 U8892 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n7258) );
  NAND2_X1 U8893 ( .A1(n10324), .A2(n7714), .ZN(n7257) );
  NAND2_X1 U8894 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9039) );
  OAI211_X1 U8895 ( .C1(n10337), .C2(n7258), .A(n7257), .B(n9039), .ZN(n7259)
         );
  OR3_X1 U8896 ( .A1(n7261), .A2(n7260), .A3(n7259), .ZN(P1_U3256) );
  NAND2_X1 U8897 ( .A1(n7300), .A2(n7961), .ZN(n7263) );
  NAND2_X1 U8898 ( .A1(n9348), .A2(n7936), .ZN(n7262) );
  NAND2_X1 U8899 ( .A1(n7263), .A2(n7262), .ZN(n7264) );
  XNOR2_X1 U8900 ( .A(n7264), .B(n7956), .ZN(n7322) );
  AND2_X1 U8901 ( .A1(n9348), .A2(n6566), .ZN(n7265) );
  AOI21_X1 U8902 ( .B1(n7300), .B2(n7936), .A(n7265), .ZN(n7323) );
  XNOR2_X1 U8903 ( .A(n7322), .B(n7323), .ZN(n7273) );
  NAND2_X1 U8904 ( .A1(n7267), .A2(n7266), .ZN(n7269) );
  INV_X1 U8905 ( .A(n7273), .ZN(n7270) );
  INV_X1 U8906 ( .A(n7327), .ZN(n7271) );
  AOI211_X1 U8907 ( .C1(n7273), .C2(n7272), .A(n9049), .B(n7271), .ZN(n7280)
         );
  NAND2_X1 U8908 ( .A1(n7300), .A2(n9047), .ZN(n7278) );
  AND2_X1 U8909 ( .A1(P1_U3084), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n10322) );
  AOI21_X1 U8910 ( .B1(n9041), .B2(n9349), .A(n10322), .ZN(n7277) );
  NAND2_X1 U8911 ( .A1(n9042), .A2(n7274), .ZN(n7276) );
  NAND2_X1 U8912 ( .A1(n9030), .A2(n10253), .ZN(n7275) );
  NAND4_X1 U8913 ( .A1(n7278), .A2(n7277), .A3(n7276), .A4(n7275), .ZN(n7279)
         );
  OR2_X1 U8914 ( .A1(n7280), .A2(n7279), .ZN(P1_U3234) );
  NAND2_X1 U8915 ( .A1(n7281), .A2(n9094), .ZN(n7417) );
  NAND2_X1 U8916 ( .A1(n7417), .A2(n7416), .ZN(n7287) );
  NAND2_X1 U8917 ( .A1(n7282), .A2(n6840), .ZN(n7285) );
  AOI22_X1 U8918 ( .A1(n7785), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n4614), .B2(
        n7283), .ZN(n7284) );
  NAND2_X1 U8919 ( .A1(n7407), .A2(n7286), .ZN(n10248) );
  NAND2_X1 U8920 ( .A1(n9161), .A2(n10248), .ZN(n9289) );
  XNOR2_X1 U8921 ( .A(n7287), .B(n9289), .ZN(n7295) );
  NAND2_X1 U8922 ( .A1(n4481), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n7294) );
  INV_X1 U8923 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n7288) );
  NAND2_X1 U8924 ( .A1(n7289), .A2(n7288), .ZN(n7290) );
  AND2_X1 U8925 ( .A1(n7383), .A2(n7290), .ZN(n10258) );
  NAND2_X1 U8926 ( .A1(n7984), .A2(n10258), .ZN(n7293) );
  NAND2_X1 U8927 ( .A1(n4480), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n7292) );
  NAND2_X1 U8928 ( .A1(n9118), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n7291) );
  NAND4_X1 U8929 ( .A1(n7294), .A2(n7293), .A3(n7292), .A4(n7291), .ZN(n9347)
         );
  AOI222_X1 U8930 ( .A1(n10355), .A2(n7295), .B1(n9347), .B2(n10254), .C1(
        n9348), .C2(n10252), .ZN(n10276) );
  INV_X1 U8931 ( .A(n7407), .ZN(n10277) );
  OAI211_X1 U8932 ( .C1(n7296), .C2(n10277), .A(n9721), .B(n10242), .ZN(n10275) );
  INV_X1 U8933 ( .A(n10275), .ZN(n7299) );
  AOI22_X1 U8934 ( .A1(n10362), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n7331), .B2(
        n10360), .ZN(n7297) );
  OAI21_X1 U8935 ( .B1(n10277), .B2(n10364), .A(n7297), .ZN(n7298) );
  AOI21_X1 U8936 ( .B1(n7299), .B2(n9626), .A(n7298), .ZN(n7307) );
  NOR2_X1 U8937 ( .A1(n10362), .A2(n10358), .ZN(n7305) );
  NAND2_X1 U8938 ( .A1(n7300), .A2(n9348), .ZN(n7301) );
  OAI21_X1 U8939 ( .B1(n7303), .B2(n9289), .A(n7408), .ZN(n7304) );
  INV_X1 U8940 ( .A(n7304), .ZN(n10280) );
  OAI21_X1 U8941 ( .B1(n10344), .B2(n7305), .A(n10280), .ZN(n7306) );
  OAI211_X1 U8942 ( .C1(n10276), .C2(n10362), .A(n7307), .B(n7306), .ZN(
        P1_U3279) );
  AOI211_X1 U8943 ( .C1(n7310), .C2(n10485), .A(n7309), .B(n7308), .ZN(n7316)
         );
  INV_X1 U8944 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n7311) );
  OAI22_X1 U8945 ( .A1(n7312), .A2(n8847), .B1(n10496), .B2(n7311), .ZN(n7313)
         );
  INV_X1 U8946 ( .A(n7313), .ZN(n7314) );
  OAI21_X1 U8947 ( .B1(n7316), .B2(n10494), .A(n7314), .ZN(P2_U3487) );
  AOI22_X1 U8948 ( .A1(n7395), .A2(n8773), .B1(n10504), .B2(
        P2_REG1_REG_12__SCAN_IN), .ZN(n7315) );
  OAI21_X1 U8949 ( .B1(n7316), .B2(n10504), .A(n7315), .ZN(P2_U3532) );
  NAND2_X1 U8950 ( .A1(n7407), .A2(n7750), .ZN(n7318) );
  NAND2_X1 U8951 ( .A1(n10253), .A2(n7973), .ZN(n7317) );
  NAND2_X1 U8952 ( .A1(n7318), .A2(n7317), .ZN(n7319) );
  XNOR2_X1 U8953 ( .A(n7319), .B(n7956), .ZN(n7369) );
  AND2_X1 U8954 ( .A1(n10253), .A2(n7320), .ZN(n7321) );
  AOI21_X1 U8955 ( .B1(n7407), .B2(n7936), .A(n7321), .ZN(n7368) );
  XNOR2_X1 U8956 ( .A(n7369), .B(n7368), .ZN(n7330) );
  INV_X1 U8957 ( .A(n7322), .ZN(n7325) );
  INV_X1 U8958 ( .A(n7323), .ZN(n7324) );
  NAND2_X1 U8959 ( .A1(n7325), .A2(n7324), .ZN(n7326) );
  INV_X1 U8960 ( .A(n7371), .ZN(n7328) );
  AOI21_X1 U8961 ( .B1(n7330), .B2(n7329), .A(n7328), .ZN(n7336) );
  INV_X1 U8962 ( .A(n9347), .ZN(n9172) );
  AOI22_X1 U8963 ( .A1(n9041), .A2(n9348), .B1(P1_REG3_REG_12__SCAN_IN), .B2(
        P1_U3084), .ZN(n7333) );
  NAND2_X1 U8964 ( .A1(n9042), .A2(n7331), .ZN(n7332) );
  OAI211_X1 U8965 ( .C1(n9172), .C2(n9045), .A(n7333), .B(n7332), .ZN(n7334)
         );
  AOI21_X1 U8966 ( .B1(n7407), .B2(n9047), .A(n7334), .ZN(n7335) );
  OAI21_X1 U8967 ( .B1(n7336), .B2(n9049), .A(n7335), .ZN(P1_U3222) );
  INV_X1 U8968 ( .A(n7172), .ZN(n7339) );
  NOR3_X1 U8969 ( .A1(n7337), .A2(n7400), .A3(n8142), .ZN(n7338) );
  AOI21_X1 U8970 ( .B1(n7339), .B2(n10194), .A(n7338), .ZN(n7347) );
  INV_X1 U8971 ( .A(n7465), .ZN(n8415) );
  AOI22_X1 U8972 ( .A1(n8119), .A2(n8416), .B1(n7611), .B2(n8415), .ZN(n7340)
         );
  NAND2_X1 U8973 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3152), .ZN(n7357) );
  OAI211_X1 U8974 ( .C1(n7341), .C2(n10199), .A(n7340), .B(n7357), .ZN(n7344)
         );
  NOR2_X1 U8975 ( .A1(n7342), .A2(n8156), .ZN(n7343) );
  AOI211_X1 U8976 ( .C1(n8137), .C2(n7462), .A(n7344), .B(n7343), .ZN(n7345)
         );
  OAI21_X1 U8977 ( .B1(n7347), .B2(n7346), .A(n7345), .ZN(P2_U3217) );
  NOR2_X1 U8978 ( .A1(n7353), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n7349) );
  NOR2_X1 U8979 ( .A1(n7349), .A2(n7348), .ZN(n7351) );
  INV_X1 U8980 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n7559) );
  AOI22_X1 U8981 ( .A1(n7555), .A2(n7559), .B1(P2_REG2_REG_14__SCAN_IN), .B2(
        n7560), .ZN(n7350) );
  NOR2_X1 U8982 ( .A1(n7351), .A2(n7350), .ZN(n7558) );
  AOI21_X1 U8983 ( .B1(n7351), .B2(n7350), .A(n7558), .ZN(n7363) );
  INV_X1 U8984 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n7500) );
  AOI22_X1 U8985 ( .A1(n7555), .A2(P2_REG1_REG_14__SCAN_IN), .B1(n7500), .B2(
        n7560), .ZN(n7355) );
  OAI21_X1 U8986 ( .B1(n7353), .B2(P2_REG1_REG_13__SCAN_IN), .A(n7352), .ZN(
        n7354) );
  NAND2_X1 U8987 ( .A1(n7355), .A2(n7354), .ZN(n7554) );
  OAI21_X1 U8988 ( .B1(n7355), .B2(n7354), .A(n7554), .ZN(n7356) );
  NAND2_X1 U8989 ( .A1(n7356), .A2(n10402), .ZN(n7362) );
  INV_X1 U8990 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7358) );
  OAI21_X1 U8991 ( .B1(n7359), .B2(n7358), .A(n7357), .ZN(n7360) );
  AOI21_X1 U8992 ( .B1(n8491), .B2(n7555), .A(n7360), .ZN(n7361) );
  OAI211_X1 U8993 ( .C1(n7363), .C2(n10405), .A(n7362), .B(n7361), .ZN(
        P2_U3259) );
  INV_X1 U8994 ( .A(n7876), .ZN(n7366) );
  OAI222_X1 U8995 ( .A1(n7364), .A2(P1_U3084), .B1(n9773), .B2(n7366), .C1(
        n7877), .C2(n9774), .ZN(P1_U3329) );
  OAI222_X1 U8996 ( .A1(P2_U3152), .A2(n7367), .B1(n7595), .B2(n7366), .C1(
        n7365), .C2(n7510), .ZN(P2_U3334) );
  NAND2_X1 U8997 ( .A1(n7369), .A2(n7368), .ZN(n7370) );
  NAND2_X1 U8998 ( .A1(n7372), .A2(n6840), .ZN(n7375) );
  AOI22_X1 U8999 ( .A1(n7785), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n4614), .B2(
        n7373), .ZN(n7374) );
  NAND2_X1 U9000 ( .A1(n9174), .A2(n7961), .ZN(n7377) );
  NAND2_X1 U9001 ( .A1(n9347), .A2(n7936), .ZN(n7376) );
  NAND2_X1 U9002 ( .A1(n7377), .A2(n7376), .ZN(n7378) );
  XNOR2_X1 U9003 ( .A(n7378), .B(n7956), .ZN(n7704) );
  AND2_X1 U9004 ( .A1(n9347), .A2(n7320), .ZN(n7379) );
  AOI21_X1 U9005 ( .B1(n9174), .B2(n7936), .A(n7379), .ZN(n7703) );
  XNOR2_X1 U9006 ( .A(n7704), .B(n7703), .ZN(n7380) );
  XNOR2_X1 U9007 ( .A(n7705), .B(n7380), .ZN(n7394) );
  NAND2_X1 U9008 ( .A1(n4481), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n7388) );
  INV_X1 U9009 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n7382) );
  NAND2_X1 U9010 ( .A1(n7383), .A2(n7382), .ZN(n7384) );
  AND2_X1 U9011 ( .A1(n7419), .A2(n7384), .ZN(n8892) );
  NAND2_X1 U9012 ( .A1(n7984), .A2(n8892), .ZN(n7387) );
  NAND2_X1 U9013 ( .A1(n4480), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n7386) );
  NAND2_X1 U9014 ( .A1(n9118), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n7385) );
  NAND4_X1 U9015 ( .A1(n7388), .A2(n7387), .A3(n7386), .A4(n7385), .ZN(n10255)
         );
  INV_X1 U9016 ( .A(n10255), .ZN(n9636) );
  AOI21_X1 U9017 ( .B1(n9041), .B2(n10253), .A(n7389), .ZN(n7391) );
  NAND2_X1 U9018 ( .A1(n9042), .A2(n10258), .ZN(n7390) );
  OAI211_X1 U9019 ( .C1(n9636), .C2(n9045), .A(n7391), .B(n7390), .ZN(n7392)
         );
  AOI21_X1 U9020 ( .B1(n9174), .B2(n9047), .A(n7392), .ZN(n7393) );
  OAI21_X1 U9021 ( .B1(n7394), .B2(n9049), .A(n7393), .ZN(P1_U3232) );
  INV_X1 U9022 ( .A(n10227), .ZN(n10233) );
  OR2_X1 U9023 ( .A1(n10227), .A2(n7400), .ZN(n8311) );
  NAND2_X1 U9024 ( .A1(n10227), .A2(n7400), .ZN(n8304) );
  NAND2_X1 U9025 ( .A1(n8311), .A2(n8304), .ZN(n10212) );
  OR2_X1 U9026 ( .A1(n7462), .A2(n7475), .ZN(n8313) );
  NAND2_X1 U9027 ( .A1(n7462), .A2(n7475), .ZN(n8314) );
  NAND2_X1 U9028 ( .A1(n8313), .A2(n8314), .ZN(n8316) );
  INV_X1 U9029 ( .A(n8316), .ZN(n7463) );
  XNOR2_X1 U9030 ( .A(n7464), .B(n7463), .ZN(n7496) );
  INV_X1 U9031 ( .A(n7496), .ZN(n7406) );
  AND2_X1 U9032 ( .A1(n8309), .A2(n8243), .ZN(n8302) );
  NAND2_X1 U9033 ( .A1(n10215), .A2(n8304), .ZN(n7398) );
  XNOR2_X1 U9034 ( .A(n7398), .B(n8316), .ZN(n7399) );
  OAI222_X1 U9035 ( .A1(n10427), .A2(n7465), .B1(n10429), .B2(n7400), .C1(
        n7399), .C2(n8637), .ZN(n7494) );
  INV_X1 U9036 ( .A(n7462), .ZN(n7502) );
  AOI211_X1 U9037 ( .C1(n7462), .C2(n4496), .A(n10472), .B(n7468), .ZN(n7495)
         );
  NAND2_X1 U9038 ( .A1(n7495), .A2(n10422), .ZN(n7403) );
  AOI22_X1 U9039 ( .A1(n10456), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n7401), .B2(
        n10447), .ZN(n7402) );
  OAI211_X1 U9040 ( .C1(n7502), .C2(n10439), .A(n7403), .B(n7402), .ZN(n7404)
         );
  AOI21_X1 U9041 ( .B1(n7494), .B2(n10211), .A(n7404), .ZN(n7405) );
  OAI21_X1 U9042 ( .B1(n8717), .B2(n7406), .A(n7405), .ZN(P2_U3282) );
  OR2_X1 U9043 ( .A1(n9174), .A2(n9347), .ZN(n9160) );
  NAND2_X1 U9044 ( .A1(n10241), .A2(n9160), .ZN(n7409) );
  NAND2_X1 U9045 ( .A1(n9174), .A2(n9347), .ZN(n9159) );
  NAND2_X1 U9046 ( .A1(n7410), .A2(n6840), .ZN(n7413) );
  AOI22_X1 U9047 ( .A1(n7785), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n4614), .B2(
        n7411), .ZN(n7412) );
  OR2_X1 U9048 ( .A1(n9739), .A2(n9636), .ZN(n8044) );
  NAND2_X1 U9049 ( .A1(n9739), .A2(n9636), .ZN(n9158) );
  NAND2_X1 U9050 ( .A1(n8044), .A2(n9158), .ZN(n9291) );
  XNOR2_X1 U9051 ( .A(n8030), .B(n9291), .ZN(n9743) );
  INV_X1 U9052 ( .A(n9644), .ZN(n7414) );
  AOI211_X1 U9053 ( .C1(n9739), .C2(n10243), .A(n10388), .B(n7414), .ZN(n9738)
         );
  AOI22_X1 U9054 ( .A1(n10362), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n8892), .B2(
        n10360), .ZN(n7415) );
  OAI21_X1 U9055 ( .B1(n4711), .B2(n10364), .A(n7415), .ZN(n7430) );
  AND2_X1 U9056 ( .A1(n9161), .A2(n7416), .ZN(n9166) );
  OR2_X1 U9057 ( .A1(n9174), .A2(n9172), .ZN(n9099) );
  NAND2_X1 U9058 ( .A1(n9174), .A2(n9172), .ZN(n9087) );
  NAND2_X1 U9059 ( .A1(n9099), .A2(n9087), .ZN(n10247) );
  INV_X1 U9060 ( .A(n9087), .ZN(n9098) );
  NOR2_X1 U9061 ( .A1(n8045), .A2(n9620), .ZN(n7428) );
  OAI21_X1 U9062 ( .B1(n10246), .B2(n9098), .A(n9291), .ZN(n7427) );
  NAND2_X1 U9063 ( .A1(n4481), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n7425) );
  INV_X1 U9064 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n7418) );
  NAND2_X1 U9065 ( .A1(n7419), .A2(n7418), .ZN(n7420) );
  AND2_X1 U9066 ( .A1(n7730), .A2(n7420), .ZN(n9647) );
  NAND2_X1 U9067 ( .A1(n7984), .A2(n9647), .ZN(n7424) );
  NAND2_X1 U9068 ( .A1(n4480), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n7423) );
  NAND2_X1 U9069 ( .A1(n9118), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n7422) );
  NAND4_X1 U9070 ( .A1(n7425), .A2(n7424), .A3(n7423), .A4(n7422), .ZN(n9346)
         );
  OAI22_X1 U9071 ( .A1(n9172), .A2(n10352), .B1(n9621), .B2(n10350), .ZN(n7426) );
  AOI21_X1 U9072 ( .B1(n7428), .B2(n7427), .A(n7426), .ZN(n9741) );
  NOR2_X1 U9073 ( .A1(n9741), .A2(n10362), .ZN(n7429) );
  AOI211_X1 U9074 ( .C1(n9626), .C2(n9738), .A(n7430), .B(n7429), .ZN(n7431)
         );
  OAI21_X1 U9075 ( .B1(n9633), .B2(n9743), .A(n7431), .ZN(P1_U3277) );
  INV_X1 U9076 ( .A(n7432), .ZN(n7434) );
  AOI21_X1 U9077 ( .B1(n7434), .B2(n7714), .A(n7433), .ZN(n7436) );
  XNOR2_X1 U9078 ( .A(n9366), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n7435) );
  NOR2_X1 U9079 ( .A1(n7436), .A2(n7435), .ZN(n9365) );
  AOI211_X1 U9080 ( .C1(n7436), .C2(n7435), .A(n9365), .B(n9367), .ZN(n7447)
         );
  NAND2_X1 U9081 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n9366), .ZN(n7439) );
  OAI21_X1 U9082 ( .B1(n9366), .B2(P1_REG2_REG_16__SCAN_IN), .A(n7439), .ZN(
        n7440) );
  AOI211_X1 U9083 ( .C1(n7441), .C2(n7440), .A(n9360), .B(n9385), .ZN(n7446)
         );
  INV_X1 U9084 ( .A(n9366), .ZN(n7443) );
  NAND2_X1 U9085 ( .A1(n10299), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n7442) );
  NAND2_X1 U9086 ( .A1(P1_U3084), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n8938) );
  OAI211_X1 U9087 ( .C1(n7444), .C2(n7443), .A(n7442), .B(n8938), .ZN(n7445)
         );
  OR3_X1 U9088 ( .A1(n7447), .A2(n7446), .A3(n7445), .ZN(P1_U3257) );
  INV_X1 U9089 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7459) );
  INV_X1 U9090 ( .A(n7451), .ZN(n7452) );
  NAND2_X1 U9091 ( .A1(n7452), .A2(SI_24_), .ZN(n7453) );
  INV_X1 U9092 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7903) );
  MUX2_X1 U9093 ( .A(n7459), .B(n7903), .S(n7590), .Z(n7455) );
  INV_X1 U9094 ( .A(SI_25_), .ZN(n10091) );
  NAND2_X1 U9095 ( .A1(n7455), .A2(n10091), .ZN(n7503) );
  INV_X1 U9096 ( .A(n7455), .ZN(n7456) );
  NAND2_X1 U9097 ( .A1(n7456), .A2(SI_25_), .ZN(n7457) );
  NAND2_X1 U9098 ( .A1(n7503), .A2(n7457), .ZN(n7504) );
  INV_X1 U9099 ( .A(n7902), .ZN(n7460) );
  OAI222_X1 U9100 ( .A1(n7510), .A2(n7459), .B1(n7595), .B2(n7460), .C1(
        P2_U3152), .C2(n7458), .ZN(P2_U3333) );
  OAI222_X1 U9101 ( .A1(P1_U3084), .A2(n7461), .B1(n9773), .B2(n7460), .C1(
        n7903), .C2(n9774), .ZN(P1_U3328) );
  OR2_X1 U9102 ( .A1(n8804), .A2(n7465), .ZN(n8318) );
  NAND2_X1 U9103 ( .A1(n8804), .A2(n7465), .ZN(n8319) );
  NAND2_X1 U9104 ( .A1(n7466), .A2(n8210), .ZN(n7481) );
  OAI21_X1 U9105 ( .B1(n7466), .B2(n8210), .A(n7481), .ZN(n8802) );
  INV_X1 U9106 ( .A(n8804), .ZN(n7467) );
  OAI21_X1 U9107 ( .B1(n7468), .B2(n7467), .A(n10418), .ZN(n7469) );
  OR2_X1 U9108 ( .A1(n7469), .A2(n7487), .ZN(n8805) );
  OAI22_X1 U9109 ( .A1(n10211), .A2(n7470), .B1(n10198), .B2(n10208), .ZN(
        n7471) );
  AOI21_X1 U9110 ( .B1(n8804), .B2(n10228), .A(n7471), .ZN(n7472) );
  OAI21_X1 U9111 ( .B1(n8805), .B2(n10206), .A(n7472), .ZN(n7478) );
  INV_X1 U9112 ( .A(n8304), .ZN(n7473) );
  NOR2_X1 U9113 ( .A1(n8316), .A2(n7473), .ZN(n7474) );
  XNOR2_X1 U9114 ( .A(n7484), .B(n8317), .ZN(n7476) );
  OAI22_X1 U9115 ( .A1(n7475), .A2(n10429), .B1(n7544), .B2(n10427), .ZN(
        n10187) );
  AOI21_X1 U9116 ( .B1(n7476), .B2(n10432), .A(n10187), .ZN(n8806) );
  NOR2_X1 U9117 ( .A1(n8806), .A2(n10456), .ZN(n7477) );
  AOI211_X1 U9118 ( .C1(n8723), .C2(n8802), .A(n7478), .B(n7477), .ZN(n7479)
         );
  INV_X1 U9119 ( .A(n7479), .ZN(P2_U3281) );
  OR2_X1 U9120 ( .A1(n8799), .A2(n7544), .ZN(n8239) );
  AND2_X1 U9121 ( .A1(n8799), .A2(n7544), .ZN(n8241) );
  INV_X1 U9122 ( .A(n8241), .ZN(n7480) );
  AOI21_X1 U9123 ( .B1(n8321), .B2(n7482), .A(n7538), .ZN(n7483) );
  INV_X1 U9124 ( .A(n7483), .ZN(n8801) );
  NAND2_X1 U9125 ( .A1(n7484), .A2(n8318), .ZN(n7485) );
  INV_X1 U9126 ( .A(n8321), .ZN(n8211) );
  XNOR2_X1 U9127 ( .A(n7542), .B(n8211), .ZN(n7486) );
  AOI22_X1 U9128 ( .A1(n8415), .A2(n10216), .B1(n8413), .B2(n8701), .ZN(n7517)
         );
  OAI21_X1 U9129 ( .B1(n7486), .B2(n8637), .A(n7517), .ZN(n8797) );
  INV_X1 U9130 ( .A(n8799), .ZN(n7518) );
  INV_X1 U9131 ( .A(n7487), .ZN(n7489) );
  INV_X1 U9132 ( .A(n7546), .ZN(n7488) );
  AOI211_X1 U9133 ( .C1(n8799), .C2(n7489), .A(n10472), .B(n7488), .ZN(n8798)
         );
  NAND2_X1 U9134 ( .A1(n8798), .A2(n10422), .ZN(n7491) );
  AOI22_X1 U9135 ( .A1(n10456), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n7521), .B2(
        n10447), .ZN(n7490) );
  OAI211_X1 U9136 ( .C1(n7518), .C2(n10439), .A(n7491), .B(n7490), .ZN(n7492)
         );
  AOI21_X1 U9137 ( .B1(n8797), .B2(n10211), .A(n7492), .ZN(n7493) );
  OAI21_X1 U9138 ( .B1(n8801), .B2(n8717), .A(n7493), .ZN(P2_U3280) );
  INV_X1 U9139 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n7497) );
  AOI211_X1 U9140 ( .C1(n7496), .C2(n10485), .A(n7495), .B(n7494), .ZN(n7499)
         );
  MUX2_X1 U9141 ( .A(n7497), .B(n7499), .S(n10496), .Z(n7498) );
  OAI21_X1 U9142 ( .B1(n7502), .B2(n8847), .A(n7498), .ZN(P2_U3493) );
  MUX2_X1 U9143 ( .A(n7500), .B(n7499), .S(n10499), .Z(n7501) );
  OAI21_X1 U9144 ( .B1(n7502), .B2(n8776), .A(n7501), .ZN(P2_U3534) );
  INV_X1 U9145 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7511) );
  INV_X1 U9146 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7923) );
  MUX2_X1 U9147 ( .A(n7511), .B(n7923), .S(n7590), .Z(n7506) );
  INV_X1 U9148 ( .A(SI_26_), .ZN(n10124) );
  NAND2_X1 U9149 ( .A1(n7506), .A2(n10124), .ZN(n7526) );
  INV_X1 U9150 ( .A(n7506), .ZN(n7507) );
  NAND2_X1 U9151 ( .A1(n7507), .A2(SI_26_), .ZN(n7508) );
  INV_X1 U9152 ( .A(n7922), .ZN(n7512) );
  OAI222_X1 U9153 ( .A1(n7509), .A2(P1_U3084), .B1(n9773), .B2(n7512), .C1(
        n7923), .C2(n9774), .ZN(P1_U3327) );
  OAI222_X1 U9154 ( .A1(P2_U3152), .A2(n7513), .B1(n8872), .B2(n7512), .C1(
        n7511), .C2(n7510), .ZN(P2_U3332) );
  XOR2_X1 U9155 ( .A(n7515), .B(n7516), .Z(n7523) );
  INV_X1 U9156 ( .A(n10199), .ZN(n8164) );
  INV_X1 U9157 ( .A(n10188), .ZN(n8150) );
  OAI22_X1 U9158 ( .A1(n8150), .A2(n7517), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8461), .ZN(n7520) );
  NOR2_X1 U9159 ( .A1(n7518), .A2(n8167), .ZN(n7519) );
  AOI211_X1 U9160 ( .C1(n8164), .C2(n7521), .A(n7520), .B(n7519), .ZN(n7522)
         );
  OAI21_X1 U9161 ( .B1(n7523), .B2(n8156), .A(n7522), .ZN(P2_U3228) );
  INV_X1 U9162 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n7528) );
  INV_X1 U9163 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n7947) );
  MUX2_X1 U9164 ( .A(n7528), .B(n7947), .S(n7590), .Z(n7530) );
  INV_X1 U9165 ( .A(SI_27_), .ZN(n7529) );
  NAND2_X1 U9166 ( .A1(n7530), .A2(n7529), .ZN(n7570) );
  INV_X1 U9167 ( .A(n7530), .ZN(n7531) );
  NAND2_X1 U9168 ( .A1(n7531), .A2(SI_27_), .ZN(n7532) );
  AND2_X1 U9169 ( .A1(n7570), .A2(n7532), .ZN(n7568) );
  INV_X1 U9170 ( .A(n7946), .ZN(n7537) );
  INV_X1 U9171 ( .A(n8401), .ZN(n8523) );
  AOI22_X1 U9172 ( .A1(n8523), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_27__SCAN_IN), .B2(n8869), .ZN(n7533) );
  OAI21_X1 U9173 ( .B1(n7537), .B2(n7595), .A(n7533), .ZN(P2_U3331) );
  AOI21_X1 U9174 ( .B1(n7535), .B2(P2_DATAO_REG_27__SCAN_IN), .A(n7534), .ZN(
        n7536) );
  OAI21_X1 U9175 ( .B1(n7537), .B2(n9773), .A(n7536), .ZN(P1_U3326) );
  INV_X1 U9176 ( .A(n8413), .ZN(n8143) );
  NAND2_X1 U9177 ( .A1(n8794), .A2(n8143), .ZN(n8238) );
  OAI21_X1 U9178 ( .B1(n7540), .B2(n7539), .A(n7573), .ZN(n7541) );
  INV_X1 U9179 ( .A(n7541), .ZN(n8796) );
  XNOR2_X1 U9180 ( .A(n7581), .B(n8325), .ZN(n7543) );
  OAI222_X1 U9181 ( .A1(n10427), .A2(n8086), .B1(n10429), .B2(n7544), .C1(
        n8637), .C2(n7543), .ZN(n8792) );
  INV_X1 U9182 ( .A(n7574), .ZN(n7545) );
  AOI211_X1 U9183 ( .C1(n8794), .C2(n7546), .A(n10472), .B(n7545), .ZN(n8793)
         );
  NAND2_X1 U9184 ( .A1(n10211), .A2(n8517), .ZN(n8607) );
  INV_X1 U9185 ( .A(n8607), .ZN(n8708) );
  NAND2_X1 U9186 ( .A1(n8793), .A2(n8708), .ZN(n7550) );
  INV_X1 U9187 ( .A(n7547), .ZN(n7548) );
  AOI22_X1 U9188 ( .A1(n10456), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n7548), .B2(
        n10447), .ZN(n7549) );
  OAI211_X1 U9189 ( .C1(n7551), .C2(n10439), .A(n7550), .B(n7549), .ZN(n7552)
         );
  AOI21_X1 U9190 ( .B1(n8792), .B2(n10211), .A(n7552), .ZN(n7553) );
  OAI21_X1 U9191 ( .B1(n8796), .B2(n8717), .A(n7553), .ZN(P2_U3279) );
  INV_X1 U9192 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n7556) );
  AOI211_X1 U9193 ( .C1(n7557), .C2(n7556), .A(n8456), .B(n10407), .ZN(n7567)
         );
  AOI21_X1 U9194 ( .B1(n7560), .B2(n7559), .A(n7558), .ZN(n8463) );
  XNOR2_X1 U9195 ( .A(n8463), .B(n8464), .ZN(n7561) );
  NOR2_X1 U9196 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n7561), .ZN(n8465) );
  AOI21_X1 U9197 ( .B1(n7561), .B2(P2_REG2_REG_15__SCAN_IN), .A(n8465), .ZN(
        n7562) );
  NOR2_X1 U9198 ( .A1(n7562), .A2(n10405), .ZN(n7566) );
  AND2_X1 U9199 ( .A1(P2_U3152), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n7563) );
  AOI21_X1 U9200 ( .B1(n10404), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n7563), .ZN(
        n7564) );
  OAI21_X1 U9201 ( .B1(n10406), .B2(n8455), .A(n7564), .ZN(n7565) );
  OR3_X1 U9202 ( .A1(n7567), .A2(n7566), .A3(n7565), .ZN(P2_U3260) );
  MUX2_X1 U9203 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n7590), .Z(n7587) );
  INV_X1 U9204 ( .A(SI_28_), .ZN(n7588) );
  XNOR2_X1 U9205 ( .A(n7587), .B(n7588), .ZN(n7585) );
  INV_X1 U9206 ( .A(n7958), .ZN(n8070) );
  AOI22_X1 U9207 ( .A1(n7571), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_28__SCAN_IN), .B2(n8869), .ZN(n7572) );
  OAI21_X1 U9208 ( .B1(n8070), .B2(n7595), .A(n7572), .ZN(P2_U3330) );
  OR2_X1 U9209 ( .A1(n8788), .A2(n8086), .ZN(n8332) );
  NAND2_X1 U9210 ( .A1(n8788), .A2(n8086), .ZN(n8331) );
  XNOR2_X1 U9211 ( .A(n7632), .B(n8213), .ZN(n8861) );
  NAND2_X1 U9212 ( .A1(n8788), .A2(n7574), .ZN(n7575) );
  NAND2_X1 U9213 ( .A1(n7575), .A2(n10418), .ZN(n7576) );
  NOR2_X1 U9214 ( .A1(n8705), .A2(n7576), .ZN(n8787) );
  NAND2_X1 U9215 ( .A1(n8788), .A2(n10228), .ZN(n7578) );
  NAND2_X1 U9216 ( .A1(n10456), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n7577) );
  OAI211_X1 U9217 ( .C1(n10208), .C2(n8148), .A(n7578), .B(n7577), .ZN(n7579)
         );
  AOI21_X1 U9218 ( .B1(n8787), .B2(n10422), .A(n7579), .ZN(n7584) );
  INV_X1 U9219 ( .A(n8236), .ZN(n7580) );
  XOR2_X1 U9220 ( .A(n7660), .B(n8213), .Z(n7582) );
  AOI22_X1 U9221 ( .A1(n8686), .A2(n8701), .B1(n10216), .B2(n8413), .ZN(n8149)
         );
  OAI21_X1 U9222 ( .B1(n7582), .B2(n8637), .A(n8149), .ZN(n8786) );
  NAND2_X1 U9223 ( .A1(n8786), .A2(n10211), .ZN(n7583) );
  OAI211_X1 U9224 ( .C1(n8861), .C2(n8717), .A(n7584), .B(n7583), .ZN(P2_U3278) );
  INV_X1 U9225 ( .A(n7587), .ZN(n7589) );
  MUX2_X1 U9226 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .S(n7590), .Z(n8168) );
  INV_X1 U9227 ( .A(SI_29_), .ZN(n7591) );
  XNOR2_X1 U9228 ( .A(n8168), .B(n7591), .ZN(n7592) );
  INV_X1 U9229 ( .A(n9051), .ZN(n7597) );
  AOI22_X1 U9230 ( .A1(n7593), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n8869), .ZN(n7594) );
  OAI21_X1 U9231 ( .B1(n7597), .B2(n7595), .A(n7594), .ZN(P2_U3329) );
  INV_X1 U9232 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n10079) );
  OAI222_X1 U9233 ( .A1(n9773), .A2(n7597), .B1(n7596), .B2(P1_U3084), .C1(
        n10079), .C2(n9774), .ZN(P1_U3324) );
  AOI22_X1 U9234 ( .A1(n9031), .A2(n7599), .B1(n7598), .B2(
        P1_REG3_REG_0__SCAN_IN), .ZN(n7602) );
  NAND2_X1 U9235 ( .A1(n7600), .A2(n8977), .ZN(n7601) );
  OAI211_X1 U9236 ( .C1(n9045), .C2(n7603), .A(n7602), .B(n7601), .ZN(P1_U3230) );
  INV_X1 U9237 ( .A(n7604), .ZN(n7606) );
  OAI21_X1 U9238 ( .B1(n10199), .B2(n7606), .A(n7605), .ZN(n7610) );
  OAI22_X1 U9239 ( .A1(n8160), .A2(n7608), .B1(n7607), .B2(n8167), .ZN(n7609)
         );
  AOI211_X1 U9240 ( .C1(n7611), .C2(n8421), .A(n7610), .B(n7609), .ZN(n7617)
         );
  AOI22_X1 U9241 ( .A1(n8057), .A2(n8423), .B1(n10194), .B2(n7612), .ZN(n7614)
         );
  OR3_X1 U9242 ( .A1(n7615), .A2(n7614), .A3(n7613), .ZN(n7616) );
  OAI211_X1 U9243 ( .C1(n7618), .C2(n8156), .A(n7617), .B(n7616), .ZN(P2_U3241) );
  NAND2_X1 U9244 ( .A1(n7958), .A2(n8189), .ZN(n7620) );
  NAND2_X1 U9245 ( .A1(n5387), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n7619) );
  INV_X1 U9246 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n10151) );
  INV_X1 U9247 ( .A(n7652), .ZN(n7622) );
  AND2_X1 U9248 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(P2_REG3_REG_28__SCAN_IN), 
        .ZN(n7621) );
  NAND2_X1 U9249 ( .A1(n7622), .A2(n7621), .ZN(n8541) );
  INV_X1 U9250 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n9904) );
  INV_X1 U9251 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n7623) );
  OAI21_X1 U9252 ( .B1(n7652), .B2(n9904), .A(n7623), .ZN(n7624) );
  NAND2_X1 U9253 ( .A1(n8541), .A2(n7624), .ZN(n8559) );
  INV_X1 U9254 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n8558) );
  NAND2_X1 U9255 ( .A1(n7670), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n7627) );
  NAND2_X1 U9256 ( .A1(n7669), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n7626) );
  OAI211_X1 U9257 ( .C1(n7673), .C2(n8558), .A(n7627), .B(n7626), .ZN(n7628)
         );
  INV_X1 U9258 ( .A(n7628), .ZN(n7629) );
  NAND2_X1 U9259 ( .A1(n7630), .A2(n7629), .ZN(n8408) );
  NAND2_X1 U9260 ( .A1(n8788), .A2(n8700), .ZN(n7631) );
  AOI22_X1 U9261 ( .A1(n7632), .A2(n7631), .B1(n4876), .B2(n8086), .ZN(n8697)
         );
  INV_X1 U9262 ( .A(n8783), .ZN(n8713) );
  INV_X1 U9263 ( .A(n8686), .ZN(n8126) );
  INV_X1 U9264 ( .A(n8702), .ZN(n8095) );
  NAND2_X1 U9265 ( .A1(n8775), .A2(n8095), .ZN(n8340) );
  NAND2_X1 U9266 ( .A1(n8350), .A2(n8340), .ZN(n8685) );
  INV_X1 U9267 ( .A(n8843), .ZN(n8678) );
  INV_X1 U9268 ( .A(n8687), .ZN(n8132) );
  NAND2_X1 U9269 ( .A1(n8678), .A2(n8132), .ZN(n7636) );
  NAND2_X1 U9270 ( .A1(n8662), .A2(n8639), .ZN(n8345) );
  OR2_X1 U9271 ( .A1(n8760), .A2(n8411), .ZN(n8356) );
  NAND2_X1 U9272 ( .A1(n8760), .A2(n8411), .ZN(n8612) );
  NAND2_X1 U9273 ( .A1(n8356), .A2(n8612), .ZN(n8640) );
  NAND2_X1 U9274 ( .A1(n8833), .A2(n8638), .ZN(n8360) );
  NAND2_X1 U9275 ( .A1(n7902), .A2(n8189), .ZN(n7639) );
  NAND2_X1 U9276 ( .A1(n5387), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n7638) );
  NAND2_X1 U9277 ( .A1(n8828), .A2(n8586), .ZN(n8231) );
  NAND2_X1 U9278 ( .A1(n7922), .A2(n8189), .ZN(n7641) );
  NAND2_X1 U9279 ( .A1(n5387), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n7640) );
  NAND2_X1 U9280 ( .A1(n7642), .A2(n10151), .ZN(n7643) );
  NAND2_X1 U9281 ( .A1(n8590), .A2(n7667), .ZN(n7649) );
  INV_X1 U9282 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n7646) );
  NAND2_X1 U9283 ( .A1(n7670), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n7645) );
  NAND2_X1 U9284 ( .A1(n7669), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n7644) );
  OAI211_X1 U9285 ( .C1(n7673), .C2(n7646), .A(n7645), .B(n7644), .ZN(n7647)
         );
  INV_X1 U9286 ( .A(n7647), .ZN(n7648) );
  NAND2_X1 U9287 ( .A1(n7649), .A2(n7648), .ZN(n8409) );
  INV_X1 U9288 ( .A(n8409), .ZN(n8074) );
  NAND2_X1 U9289 ( .A1(n8823), .A2(n8074), .ZN(n8368) );
  NAND2_X1 U9290 ( .A1(n5387), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n7650) );
  XNOR2_X1 U9291 ( .A(n7652), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n8575) );
  NAND2_X1 U9292 ( .A1(n8575), .A2(n7667), .ZN(n7658) );
  INV_X1 U9293 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n7655) );
  NAND2_X1 U9294 ( .A1(n7669), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n7654) );
  NAND2_X1 U9295 ( .A1(n7670), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n7653) );
  OAI211_X1 U9296 ( .C1(n7655), .C2(n7673), .A(n7654), .B(n7653), .ZN(n7656)
         );
  INV_X1 U9297 ( .A(n7656), .ZN(n7657) );
  NAND2_X1 U9298 ( .A1(n7658), .A2(n7657), .ZN(n8584) );
  INV_X1 U9299 ( .A(n8569), .ZN(n7659) );
  NAND2_X1 U9300 ( .A1(n7660), .A2(n8332), .ZN(n7661) );
  NAND2_X1 U9301 ( .A1(n7661), .A2(n8331), .ZN(n8698) );
  OR2_X1 U9302 ( .A1(n8783), .A2(n8126), .ZN(n8333) );
  NAND2_X1 U9303 ( .A1(n8783), .A2(n8126), .ZN(n8683) );
  AND2_X1 U9304 ( .A1(n8340), .A2(n8683), .ZN(n8328) );
  NAND2_X1 U9305 ( .A1(n8682), .A2(n8328), .ZN(n7662) );
  NAND2_X1 U9306 ( .A1(n7662), .A2(n8350), .ZN(n8667) );
  OR2_X1 U9307 ( .A1(n8843), .A2(n8132), .ZN(n8341) );
  NAND2_X1 U9308 ( .A1(n8843), .A2(n8132), .ZN(n8344) );
  NAND2_X1 U9309 ( .A1(n8341), .A2(n8344), .ZN(n8666) );
  INV_X1 U9310 ( .A(n8612), .ZN(n7663) );
  NOR2_X1 U9311 ( .A1(n8613), .A2(n7663), .ZN(n7664) );
  NAND2_X1 U9312 ( .A1(n8615), .A2(n8361), .ZN(n8596) );
  INV_X1 U9313 ( .A(n8230), .ZN(n7665) );
  OR2_X1 U9314 ( .A1(n8818), .A2(n8225), .ZN(n8226) );
  AND2_X2 U9315 ( .A1(n8571), .A2(n8226), .ZN(n8176) );
  INV_X1 U9316 ( .A(n8535), .ZN(n7666) );
  XNOR2_X1 U9317 ( .A(n8176), .B(n7666), .ZN(n7679) );
  NAND2_X1 U9318 ( .A1(n8584), .A2(n10216), .ZN(n7678) );
  INV_X1 U9319 ( .A(n8541), .ZN(n7668) );
  NAND2_X1 U9320 ( .A1(n7668), .A2(n7667), .ZN(n7676) );
  INV_X1 U9321 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n8540) );
  NAND2_X1 U9322 ( .A1(n7669), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n7672) );
  NAND2_X1 U9323 ( .A1(n7670), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n7671) );
  OAI211_X1 U9324 ( .C1(n8540), .C2(n7673), .A(n7672), .B(n7671), .ZN(n7674)
         );
  INV_X1 U9325 ( .A(n7674), .ZN(n7675) );
  NAND2_X1 U9326 ( .A1(n7676), .A2(n7675), .ZN(n8407) );
  NAND2_X1 U9327 ( .A1(n8407), .A2(n8701), .ZN(n7677) );
  NAND2_X1 U9328 ( .A1(n7678), .A2(n7677), .ZN(n8024) );
  AOI21_X1 U9329 ( .B1(n7679), .B2(n10432), .A(n8024), .ZN(n8566) );
  OAI211_X1 U9330 ( .C1(n8534), .C2(n8574), .A(n10418), .B(n8538), .ZN(n8560)
         );
  OAI211_X1 U9331 ( .C1(n8534), .C2(n10488), .A(n8566), .B(n8560), .ZN(n7682)
         );
  MUX2_X1 U9332 ( .A(n7682), .B(P2_REG0_REG_28__SCAN_IN), .S(n10494), .Z(n7680) );
  INV_X1 U9333 ( .A(n7680), .ZN(n7681) );
  OAI21_X1 U9334 ( .B1(n8556), .B2(n8860), .A(n7681), .ZN(P2_U3516) );
  MUX2_X1 U9335 ( .A(n7682), .B(P2_REG1_REG_28__SCAN_IN), .S(n10504), .Z(n7683) );
  INV_X1 U9336 ( .A(n7683), .ZN(n7684) );
  OAI21_X1 U9337 ( .B1(n8556), .B2(n8791), .A(n7684), .ZN(P2_U3548) );
  INV_X1 U9338 ( .A(n8062), .ZN(n7686) );
  AOI22_X1 U9339 ( .A1(n10188), .A2(n7687), .B1(n7686), .B2(
        P2_REG3_REG_1__SCAN_IN), .ZN(n7692) );
  OAI21_X1 U9340 ( .B1(n7689), .B2(n7688), .A(n8058), .ZN(n7690) );
  NAND2_X1 U9341 ( .A1(n10194), .A2(n7690), .ZN(n7691) );
  OAI211_X1 U9342 ( .C1(n7702), .C2(n8167), .A(n7692), .B(n7691), .ZN(P2_U3224) );
  INV_X1 U9343 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n7697) );
  NOR2_X1 U9344 ( .A1(n7693), .A2(n10472), .ZN(n7695) );
  AOI211_X1 U9345 ( .C1(n10485), .C2(n7696), .A(n7695), .B(n7694), .ZN(n7699)
         );
  MUX2_X1 U9346 ( .A(n7697), .B(n7699), .S(n10496), .Z(n7698) );
  OAI21_X1 U9347 ( .B1(n8847), .B2(n7702), .A(n7698), .ZN(P2_U3454) );
  MUX2_X1 U9348 ( .A(n7700), .B(n7699), .S(n10499), .Z(n7701) );
  OAI21_X1 U9349 ( .B1(n8776), .B2(n7702), .A(n7701), .ZN(P2_U3521) );
  NAND2_X1 U9350 ( .A1(n9739), .A2(n7961), .ZN(n7707) );
  NAND2_X1 U9351 ( .A1(n10255), .A2(n7973), .ZN(n7706) );
  NAND2_X1 U9352 ( .A1(n7707), .A2(n7706), .ZN(n7708) );
  XNOR2_X1 U9353 ( .A(n7708), .B(n7956), .ZN(n8887) );
  AND2_X1 U9354 ( .A1(n10255), .A2(n7320), .ZN(n7709) );
  AOI21_X1 U9355 ( .B1(n9739), .B2(n7936), .A(n7709), .ZN(n7711) );
  NAND2_X1 U9356 ( .A1(n8887), .A2(n7711), .ZN(n7710) );
  INV_X1 U9357 ( .A(n8887), .ZN(n7712) );
  INV_X1 U9358 ( .A(n7711), .ZN(n8886) );
  NAND2_X1 U9359 ( .A1(n7713), .A2(n6840), .ZN(n7716) );
  AOI22_X1 U9360 ( .A1(n7785), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n4614), .B2(
        n7714), .ZN(n7715) );
  NAND2_X1 U9361 ( .A1(n9731), .A2(n7750), .ZN(n7718) );
  NAND2_X1 U9362 ( .A1(n9346), .A2(n7973), .ZN(n7717) );
  NAND2_X1 U9363 ( .A1(n7718), .A2(n7717), .ZN(n7719) );
  XNOR2_X1 U9364 ( .A(n7719), .B(n7956), .ZN(n9037) );
  AND2_X1 U9365 ( .A1(n9346), .A2(n7320), .ZN(n7720) );
  AOI21_X1 U9366 ( .B1(n9731), .B2(n7973), .A(n7720), .ZN(n7721) );
  INV_X1 U9367 ( .A(n9037), .ZN(n7722) );
  INV_X1 U9368 ( .A(n7721), .ZN(n9036) );
  NAND2_X1 U9369 ( .A1(n7722), .A2(n9036), .ZN(n7723) );
  NAND2_X1 U9370 ( .A1(n7725), .A2(n6840), .ZN(n7727) );
  AOI22_X1 U9371 ( .A1(n7785), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n9366), .B2(
        n4614), .ZN(n7726) );
  NAND2_X1 U9372 ( .A1(n9728), .A2(n7961), .ZN(n7737) );
  NAND2_X1 U9373 ( .A1(n4481), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n7735) );
  INV_X1 U9374 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n7729) );
  NAND2_X1 U9375 ( .A1(n7730), .A2(n7729), .ZN(n7731) );
  AND2_X1 U9376 ( .A1(n7752), .A2(n7731), .ZN(n9627) );
  NAND2_X1 U9377 ( .A1(n7984), .A2(n9627), .ZN(n7734) );
  NAND2_X1 U9378 ( .A1(n4480), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n7733) );
  NAND2_X1 U9379 ( .A1(n9118), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n7732) );
  NAND4_X1 U9380 ( .A1(n7735), .A2(n7734), .A3(n7733), .A4(n7732), .ZN(n9606)
         );
  NAND2_X1 U9381 ( .A1(n9606), .A2(n7936), .ZN(n7736) );
  NAND2_X1 U9382 ( .A1(n7737), .A2(n7736), .ZN(n7738) );
  XNOR2_X1 U9383 ( .A(n7738), .B(n7956), .ZN(n7740) );
  AND2_X1 U9384 ( .A1(n9606), .A2(n7320), .ZN(n7739) );
  AOI21_X1 U9385 ( .B1(n9728), .B2(n7973), .A(n7739), .ZN(n7741) );
  NAND2_X1 U9386 ( .A1(n7740), .A2(n7741), .ZN(n7746) );
  INV_X1 U9387 ( .A(n7740), .ZN(n7743) );
  INV_X1 U9388 ( .A(n7741), .ZN(n7742) );
  NAND2_X1 U9389 ( .A1(n7743), .A2(n7742), .ZN(n7744) );
  NAND2_X1 U9390 ( .A1(n7746), .A2(n7744), .ZN(n8937) );
  NAND2_X1 U9391 ( .A1(n7747), .A2(n6840), .ZN(n7749) );
  AOI22_X1 U9392 ( .A1(n9383), .A2(n4614), .B1(n7785), .B2(
        P2_DATAO_REG_17__SCAN_IN), .ZN(n7748) );
  NAND2_X1 U9393 ( .A1(n9720), .A2(n7750), .ZN(n7759) );
  NAND2_X1 U9394 ( .A1(n4481), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n7757) );
  INV_X1 U9395 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n7751) );
  NAND2_X1 U9396 ( .A1(n7752), .A2(n7751), .ZN(n7753) );
  AND2_X1 U9397 ( .A1(n7771), .A2(n7753), .ZN(n9601) );
  NAND2_X1 U9398 ( .A1(n7984), .A2(n9601), .ZN(n7756) );
  NAND2_X1 U9399 ( .A1(n9118), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n7755) );
  NAND2_X1 U9400 ( .A1(n4480), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n7754) );
  NAND4_X1 U9401 ( .A1(n7757), .A2(n7756), .A3(n7755), .A4(n7754), .ZN(n9593)
         );
  NAND2_X1 U9402 ( .A1(n9593), .A2(n7936), .ZN(n7758) );
  NAND2_X1 U9403 ( .A1(n7759), .A2(n7758), .ZN(n7760) );
  XNOR2_X1 U9404 ( .A(n7760), .B(n6589), .ZN(n7762) );
  AND2_X1 U9405 ( .A1(n9593), .A2(n6566), .ZN(n7761) );
  AOI21_X1 U9406 ( .B1(n9720), .B2(n7973), .A(n7761), .ZN(n7763) );
  XNOR2_X1 U9407 ( .A(n7762), .B(n7763), .ZN(n8958) );
  INV_X1 U9408 ( .A(n7762), .ZN(n7764) );
  NAND2_X1 U9409 ( .A1(n7764), .A2(n7763), .ZN(n7765) );
  NAND2_X1 U9410 ( .A1(n7766), .A2(n6840), .ZN(n7768) );
  AOI22_X1 U9411 ( .A1(n9395), .A2(n4614), .B1(n7785), .B2(
        P2_DATAO_REG_18__SCAN_IN), .ZN(n7767) );
  NAND2_X1 U9412 ( .A1(n9715), .A2(n7961), .ZN(n7778) );
  INV_X1 U9413 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n7770) );
  NAND2_X1 U9414 ( .A1(n7771), .A2(n7770), .ZN(n7772) );
  AND2_X1 U9415 ( .A1(n7789), .A2(n7772), .ZN(n9585) );
  NAND2_X1 U9416 ( .A1(n9585), .A2(n7984), .ZN(n7776) );
  NAND2_X1 U9417 ( .A1(n4481), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n7775) );
  NAND2_X1 U9418 ( .A1(n4480), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n7774) );
  NAND2_X1 U9419 ( .A1(n9118), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n7773) );
  INV_X1 U9420 ( .A(n9573), .ZN(n9607) );
  NAND2_X1 U9421 ( .A1(n9607), .A2(n7936), .ZN(n7777) );
  NAND2_X1 U9422 ( .A1(n7778), .A2(n7777), .ZN(n7779) );
  XNOR2_X1 U9423 ( .A(n7779), .B(n7956), .ZN(n7782) );
  NAND2_X1 U9424 ( .A1(n7783), .A2(n7782), .ZN(n9009) );
  NAND2_X1 U9425 ( .A1(n9715), .A2(n7890), .ZN(n7781) );
  OR2_X1 U9426 ( .A1(n9573), .A2(n6553), .ZN(n7780) );
  NAND2_X1 U9427 ( .A1(n7781), .A2(n7780), .ZN(n9008) );
  NAND2_X1 U9428 ( .A1(n9009), .A2(n9008), .ZN(n9013) );
  NAND2_X1 U9429 ( .A1(n7784), .A2(n6840), .ZN(n7787) );
  AOI22_X1 U9430 ( .A1(n7785), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n4485), .B2(
        n4614), .ZN(n7786) );
  NAND2_X1 U9431 ( .A1(n9712), .A2(n7961), .ZN(n7794) );
  INV_X1 U9432 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n7788) );
  NAND2_X1 U9433 ( .A1(n7789), .A2(n7788), .ZN(n7790) );
  NAND2_X1 U9434 ( .A1(n7807), .A2(n7790), .ZN(n9576) );
  AOI22_X1 U9435 ( .A1(n4481), .A2(P1_REG1_REG_19__SCAN_IN), .B1(n4480), .B2(
        P1_REG0_REG_19__SCAN_IN), .ZN(n7792) );
  NAND2_X1 U9436 ( .A1(n9118), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n7791) );
  OAI211_X1 U9437 ( .C1(n9576), .C2(n7929), .A(n7792), .B(n7791), .ZN(n9592)
         );
  NAND2_X1 U9438 ( .A1(n9592), .A2(n7936), .ZN(n7793) );
  NAND2_X1 U9439 ( .A1(n7794), .A2(n7793), .ZN(n7795) );
  XNOR2_X1 U9440 ( .A(n7795), .B(n6589), .ZN(n7798) );
  NAND2_X1 U9441 ( .A1(n9712), .A2(n7973), .ZN(n7797) );
  NAND2_X1 U9442 ( .A1(n9592), .A2(n7320), .ZN(n7796) );
  NAND2_X1 U9443 ( .A1(n7797), .A2(n7796), .ZN(n7799) );
  AND2_X1 U9444 ( .A1(n7798), .A2(n7799), .ZN(n8908) );
  INV_X1 U9445 ( .A(n7798), .ZN(n7801) );
  INV_X1 U9446 ( .A(n7799), .ZN(n7800) );
  NAND2_X1 U9447 ( .A1(n7801), .A2(n7800), .ZN(n8907) );
  NAND2_X1 U9448 ( .A1(n7802), .A2(n6840), .ZN(n7804) );
  OR2_X1 U9449 ( .A1(n6409), .A2(n10077), .ZN(n7803) );
  NAND2_X1 U9450 ( .A1(n9707), .A2(n7961), .ZN(n7813) );
  INV_X1 U9451 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n9557) );
  INV_X1 U9452 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n7806) );
  NAND2_X1 U9453 ( .A1(n7807), .A2(n7806), .ZN(n7808) );
  NAND2_X1 U9454 ( .A1(n7824), .A2(n7808), .ZN(n9556) );
  OR2_X1 U9455 ( .A1(n9556), .A2(n7929), .ZN(n7810) );
  AOI22_X1 U9456 ( .A1(n4481), .A2(P1_REG1_REG_20__SCAN_IN), .B1(n4480), .B2(
        P1_REG0_REG_20__SCAN_IN), .ZN(n7809) );
  OAI211_X1 U9457 ( .C1(n7811), .C2(n9557), .A(n7810), .B(n7809), .ZN(n9539)
         );
  NAND2_X1 U9458 ( .A1(n9539), .A2(n7936), .ZN(n7812) );
  NAND2_X1 U9459 ( .A1(n7813), .A2(n7812), .ZN(n7814) );
  XNOR2_X1 U9460 ( .A(n7814), .B(n6589), .ZN(n7817) );
  NAND2_X1 U9461 ( .A1(n9707), .A2(n7936), .ZN(n7816) );
  NAND2_X1 U9462 ( .A1(n9539), .A2(n6566), .ZN(n7815) );
  NAND2_X1 U9463 ( .A1(n7816), .A2(n7815), .ZN(n7818) );
  NAND2_X1 U9464 ( .A1(n7817), .A2(n7818), .ZN(n8987) );
  INV_X1 U9465 ( .A(n7817), .ZN(n7820) );
  INV_X1 U9466 ( .A(n7818), .ZN(n7819) );
  NAND2_X1 U9467 ( .A1(n7820), .A2(n7819), .ZN(n8988) );
  NAND2_X1 U9468 ( .A1(n7821), .A2(n6840), .ZN(n7823) );
  INV_X1 U9469 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n10065) );
  OR2_X1 U9470 ( .A1(n6409), .A2(n10065), .ZN(n7822) );
  NAND2_X1 U9471 ( .A1(n9701), .A2(n7961), .ZN(n7833) );
  INV_X1 U9472 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n8918) );
  NAND2_X1 U9473 ( .A1(n7824), .A2(n8918), .ZN(n7825) );
  NAND2_X1 U9474 ( .A1(n7845), .A2(n7825), .ZN(n9535) );
  OR2_X1 U9475 ( .A1(n9535), .A2(n7929), .ZN(n7831) );
  INV_X1 U9476 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n7828) );
  NAND2_X1 U9477 ( .A1(n4480), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n7827) );
  NAND2_X1 U9478 ( .A1(n9118), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n7826) );
  OAI211_X1 U9479 ( .C1(n4828), .C2(n7828), .A(n7827), .B(n7826), .ZN(n7829)
         );
  INV_X1 U9480 ( .A(n7829), .ZN(n7830) );
  INV_X1 U9481 ( .A(n9563), .ZN(n9528) );
  NAND2_X1 U9482 ( .A1(n9528), .A2(n7890), .ZN(n7832) );
  NAND2_X1 U9483 ( .A1(n7833), .A2(n7832), .ZN(n7834) );
  XNOR2_X1 U9484 ( .A(n7834), .B(n6589), .ZN(n7836) );
  NOR2_X1 U9485 ( .A1(n9563), .A2(n6553), .ZN(n7835) );
  AOI21_X1 U9486 ( .B1(n9701), .B2(n7973), .A(n7835), .ZN(n7837) );
  XNOR2_X1 U9487 ( .A(n7836), .B(n7837), .ZN(n8916) );
  INV_X1 U9488 ( .A(n7836), .ZN(n7838) );
  NAND2_X1 U9489 ( .A1(n7838), .A2(n7837), .ZN(n7839) );
  NAND2_X1 U9490 ( .A1(n7841), .A2(n6840), .ZN(n7844) );
  OR2_X1 U9491 ( .A1(n6409), .A2(n7842), .ZN(n7843) );
  INV_X1 U9492 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9003) );
  NAND2_X1 U9493 ( .A1(n7845), .A2(n9003), .ZN(n7846) );
  NAND2_X1 U9494 ( .A1(n7864), .A2(n7846), .ZN(n9522) );
  INV_X1 U9495 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n7849) );
  NAND2_X1 U9496 ( .A1(n4480), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n7848) );
  NAND2_X1 U9497 ( .A1(n9118), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n7847) );
  OAI211_X1 U9498 ( .C1(n4828), .C2(n7849), .A(n7848), .B(n7847), .ZN(n7850)
         );
  INV_X1 U9499 ( .A(n7850), .ZN(n7851) );
  OAI21_X1 U9500 ( .B1(n9522), .B2(n7929), .A(n7851), .ZN(n9540) );
  AND2_X1 U9501 ( .A1(n9540), .A2(n7320), .ZN(n7852) );
  AOI21_X1 U9502 ( .B1(n9693), .B2(n7936), .A(n7852), .ZN(n7856) );
  NAND2_X1 U9503 ( .A1(n7857), .A2(n7856), .ZN(n8997) );
  NAND2_X1 U9504 ( .A1(n9693), .A2(n7961), .ZN(n7854) );
  NAND2_X1 U9505 ( .A1(n9540), .A2(n7890), .ZN(n7853) );
  NAND2_X1 U9506 ( .A1(n7854), .A2(n7853), .ZN(n7855) );
  XNOR2_X1 U9507 ( .A(n7855), .B(n6589), .ZN(n8996) );
  NAND2_X1 U9508 ( .A1(n7858), .A2(n6840), .ZN(n7861) );
  OR2_X1 U9509 ( .A1(n6409), .A2(n7859), .ZN(n7860) );
  INV_X1 U9510 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n7863) );
  NAND2_X1 U9511 ( .A1(n7864), .A2(n7863), .ZN(n7865) );
  NAND2_X1 U9512 ( .A1(n7882), .A2(n7865), .ZN(n9514) );
  OR2_X1 U9513 ( .A1(n9514), .A2(n7929), .ZN(n7871) );
  INV_X1 U9514 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n7868) );
  NAND2_X1 U9515 ( .A1(n4480), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n7867) );
  NAND2_X1 U9516 ( .A1(n9118), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n7866) );
  OAI211_X1 U9517 ( .C1(n4828), .C2(n7868), .A(n7867), .B(n7866), .ZN(n7869)
         );
  INV_X1 U9518 ( .A(n7869), .ZN(n7870) );
  OAI22_X1 U9519 ( .A1(n8049), .A2(n7891), .B1(n8968), .B2(n4484), .ZN(n7872)
         );
  XNOR2_X1 U9520 ( .A(n7872), .B(n7956), .ZN(n7873) );
  OAI22_X1 U9521 ( .A1(n8049), .A2(n4484), .B1(n8968), .B2(n6553), .ZN(n8901)
         );
  INV_X1 U9522 ( .A(n7873), .ZN(n7874) );
  NAND2_X1 U9523 ( .A1(n7876), .A2(n6840), .ZN(n7879) );
  OR2_X1 U9524 ( .A1(n6409), .A2(n7877), .ZN(n7878) );
  INV_X1 U9525 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n7881) );
  NAND2_X1 U9526 ( .A1(n7882), .A2(n7881), .ZN(n7883) );
  NAND2_X1 U9527 ( .A1(n7906), .A2(n7883), .ZN(n9494) );
  INV_X1 U9528 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n7886) );
  NAND2_X1 U9529 ( .A1(n4480), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n7885) );
  NAND2_X1 U9530 ( .A1(n9118), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n7884) );
  OAI211_X1 U9531 ( .C1(n4828), .C2(n7886), .A(n7885), .B(n7884), .ZN(n7887)
         );
  INV_X1 U9532 ( .A(n7887), .ZN(n7888) );
  OAI22_X1 U9533 ( .A1(n9497), .A2(n7891), .B1(n9511), .B2(n4484), .ZN(n7892)
         );
  XNOR2_X1 U9534 ( .A(n7892), .B(n7956), .ZN(n7895) );
  INV_X1 U9535 ( .A(n9511), .ZN(n9345) );
  NAND2_X1 U9536 ( .A1(n9345), .A2(n7320), .ZN(n7893) );
  NAND2_X1 U9537 ( .A1(n7895), .A2(n7896), .ZN(n7901) );
  INV_X1 U9538 ( .A(n7895), .ZN(n7898) );
  INV_X1 U9539 ( .A(n7896), .ZN(n7897) );
  NAND2_X1 U9540 ( .A1(n7898), .A2(n7897), .ZN(n7899) );
  NAND2_X1 U9541 ( .A1(n7901), .A2(n7899), .ZN(n8966) );
  OR2_X1 U9542 ( .A1(n6409), .A2(n7903), .ZN(n7904) );
  NAND2_X1 U9543 ( .A1(n9681), .A2(n7961), .ZN(n7915) );
  INV_X1 U9544 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n8928) );
  NAND2_X1 U9545 ( .A1(n7906), .A2(n8928), .ZN(n7907) );
  NAND2_X1 U9546 ( .A1(n9484), .A2(n7984), .ZN(n7913) );
  INV_X1 U9547 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n7910) );
  NAND2_X1 U9548 ( .A1(n9118), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n7909) );
  NAND2_X1 U9549 ( .A1(n4480), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n7908) );
  OAI211_X1 U9550 ( .C1(n4828), .C2(n7910), .A(n7909), .B(n7908), .ZN(n7911)
         );
  INV_X1 U9551 ( .A(n7911), .ZN(n7912) );
  NAND2_X1 U9552 ( .A1(n9501), .A2(n7890), .ZN(n7914) );
  NAND2_X1 U9553 ( .A1(n7915), .A2(n7914), .ZN(n7916) );
  XNOR2_X1 U9554 ( .A(n7916), .B(n6589), .ZN(n7918) );
  NOR2_X1 U9555 ( .A1(n9027), .A2(n6553), .ZN(n7917) );
  AOI21_X1 U9556 ( .B1(n9681), .B2(n7936), .A(n7917), .ZN(n7919) );
  XNOR2_X1 U9557 ( .A(n7918), .B(n7919), .ZN(n8926) );
  INV_X1 U9558 ( .A(n7918), .ZN(n7920) );
  NAND2_X1 U9559 ( .A1(n7920), .A2(n7919), .ZN(n7921) );
  OR2_X1 U9560 ( .A1(n6409), .A2(n7923), .ZN(n7924) );
  NAND2_X1 U9561 ( .A1(n9674), .A2(n7961), .ZN(n7938) );
  INV_X1 U9562 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n9025) );
  NAND2_X1 U9563 ( .A1(n7927), .A2(n9025), .ZN(n7928) );
  NAND2_X1 U9564 ( .A1(n7965), .A2(n7928), .ZN(n9463) );
  INV_X1 U9565 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n7932) );
  NAND2_X1 U9566 ( .A1(n4480), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n7931) );
  NAND2_X1 U9567 ( .A1(n9118), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n7930) );
  OAI211_X1 U9568 ( .C1(n4828), .C2(n7932), .A(n7931), .B(n7930), .ZN(n7933)
         );
  INV_X1 U9569 ( .A(n7933), .ZN(n7934) );
  NAND2_X1 U9570 ( .A1(n9344), .A2(n7936), .ZN(n7937) );
  NAND2_X1 U9571 ( .A1(n7938), .A2(n7937), .ZN(n7939) );
  XNOR2_X1 U9572 ( .A(n7939), .B(n6589), .ZN(n7942) );
  NAND2_X1 U9573 ( .A1(n9674), .A2(n7890), .ZN(n7941) );
  NAND2_X1 U9574 ( .A1(n9344), .A2(n6566), .ZN(n7940) );
  NAND2_X1 U9575 ( .A1(n7941), .A2(n7940), .ZN(n7943) );
  NAND2_X1 U9576 ( .A1(n7942), .A2(n7943), .ZN(n9021) );
  INV_X1 U9577 ( .A(n7942), .ZN(n7945) );
  INV_X1 U9578 ( .A(n7943), .ZN(n7944) );
  NAND2_X1 U9579 ( .A1(n7945), .A2(n7944), .ZN(n9022) );
  NAND2_X1 U9580 ( .A1(n7946), .A2(n6840), .ZN(n7949) );
  OR2_X1 U9581 ( .A1(n6409), .A2(n7947), .ZN(n7948) );
  NAND2_X1 U9582 ( .A1(n9671), .A2(n7961), .ZN(n7955) );
  XNOR2_X1 U9583 ( .A(n7965), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n8879) );
  INV_X1 U9584 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n7952) );
  NAND2_X1 U9585 ( .A1(n4480), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n7951) );
  NAND2_X1 U9586 ( .A1(n9118), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n7950) );
  OAI211_X1 U9587 ( .C1(n4828), .C2(n7952), .A(n7951), .B(n7950), .ZN(n7953)
         );
  OR2_X1 U9588 ( .A1(n9415), .A2(n4484), .ZN(n7954) );
  NAND2_X1 U9589 ( .A1(n7955), .A2(n7954), .ZN(n7957) );
  XNOR2_X1 U9590 ( .A(n7957), .B(n7956), .ZN(n8875) );
  NAND2_X1 U9591 ( .A1(n7958), .A2(n6840), .ZN(n7960) );
  INV_X1 U9592 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n10120) );
  OR2_X1 U9593 ( .A1(n6409), .A2(n10120), .ZN(n7959) );
  NAND2_X1 U9594 ( .A1(n9664), .A2(n7961), .ZN(n7975) );
  INV_X1 U9595 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n7963) );
  INV_X1 U9596 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n7962) );
  OAI21_X1 U9597 ( .B1(n7965), .B2(n7963), .A(n7962), .ZN(n7966) );
  NAND2_X1 U9598 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n7964) );
  NAND2_X1 U9599 ( .A1(n9455), .A2(n7984), .ZN(n7972) );
  INV_X1 U9600 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n7969) );
  NAND2_X1 U9601 ( .A1(n9118), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n7968) );
  NAND2_X1 U9602 ( .A1(n4480), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n7967) );
  OAI211_X1 U9603 ( .C1(n4828), .C2(n7969), .A(n7968), .B(n7967), .ZN(n7970)
         );
  INV_X1 U9604 ( .A(n7970), .ZN(n7971) );
  INV_X1 U9605 ( .A(n9430), .ZN(n9343) );
  NAND2_X1 U9606 ( .A1(n9343), .A2(n7973), .ZN(n7974) );
  NAND2_X1 U9607 ( .A1(n7975), .A2(n7974), .ZN(n7976) );
  XNOR2_X1 U9608 ( .A(n7976), .B(n6589), .ZN(n7979) );
  NOR2_X1 U9609 ( .A1(n9430), .A2(n6553), .ZN(n7977) );
  AOI21_X1 U9610 ( .B1(n9664), .B2(n7890), .A(n7977), .ZN(n7978) );
  XNOR2_X1 U9611 ( .A(n7979), .B(n7978), .ZN(n7981) );
  INV_X1 U9612 ( .A(n7981), .ZN(n7980) );
  NOR2_X1 U9613 ( .A1(n9415), .A2(n6553), .ZN(n7983) );
  AOI21_X1 U9614 ( .B1(n9671), .B2(n7890), .A(n7983), .ZN(n8874) );
  AOI22_X1 U9615 ( .A1(n9455), .A2(n9042), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n7993) );
  INV_X1 U9616 ( .A(n9433), .ZN(n7985) );
  NAND2_X1 U9617 ( .A1(n7985), .A2(n7984), .ZN(n7991) );
  INV_X1 U9618 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n7988) );
  NAND2_X1 U9619 ( .A1(n4480), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n7987) );
  NAND2_X1 U9620 ( .A1(n9118), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n7986) );
  OAI211_X1 U9621 ( .C1(n4828), .C2(n7988), .A(n7987), .B(n7986), .ZN(n7989)
         );
  INV_X1 U9622 ( .A(n7989), .ZN(n7990) );
  NAND2_X1 U9623 ( .A1(n7991), .A2(n7990), .ZN(n9442) );
  NAND2_X1 U9624 ( .A1(n9442), .A2(n9030), .ZN(n7992) );
  OAI211_X1 U9625 ( .C1(n9415), .C2(n9026), .A(n7993), .B(n7992), .ZN(n7994)
         );
  AOI21_X1 U9626 ( .B1(n9664), .B2(n9047), .A(n7994), .ZN(n7995) );
  OAI222_X1 U9627 ( .A1(n9327), .A2(P1_U3084), .B1(n9773), .B2(n7996), .C1(
        n10065), .C2(n9774), .ZN(P1_U3332) );
  NAND2_X1 U9628 ( .A1(n7998), .A2(n7997), .ZN(n8003) );
  INV_X1 U9629 ( .A(n7999), .ZN(n8001) );
  XOR2_X1 U9630 ( .A(n5263), .B(n8828), .Z(n8101) );
  NAND2_X1 U9631 ( .A1(n8618), .A2(n8016), .ZN(n8100) );
  XNOR2_X1 U9632 ( .A(n8823), .B(n8007), .ZN(n8073) );
  AND2_X1 U9633 ( .A1(n8409), .A2(n8016), .ZN(n8004) );
  NAND2_X1 U9634 ( .A1(n8073), .A2(n8004), .ZN(n8076) );
  OAI21_X1 U9635 ( .B1(n8073), .B2(n8004), .A(n8076), .ZN(n8157) );
  INV_X1 U9636 ( .A(n8157), .ZN(n8005) );
  XNOR2_X1 U9637 ( .A(n8818), .B(n8007), .ZN(n8008) );
  AND2_X1 U9638 ( .A1(n8584), .A2(n8016), .ZN(n8009) );
  NAND2_X1 U9639 ( .A1(n8008), .A2(n8009), .ZN(n8013) );
  AND2_X1 U9640 ( .A1(n8076), .A2(n8013), .ZN(n8015) );
  INV_X1 U9641 ( .A(n8013), .ZN(n8014) );
  INV_X1 U9642 ( .A(n8008), .ZN(n8011) );
  INV_X1 U9643 ( .A(n8009), .ZN(n8010) );
  NAND2_X1 U9644 ( .A1(n8011), .A2(n8010), .ZN(n8012) );
  INV_X1 U9645 ( .A(n8534), .ZN(n8563) );
  NOR2_X1 U9646 ( .A1(n8534), .A2(n8803), .ZN(n8020) );
  INV_X1 U9647 ( .A(n8020), .ZN(n8018) );
  NAND2_X1 U9648 ( .A1(n8408), .A2(n8016), .ZN(n8017) );
  XNOR2_X1 U9649 ( .A(n8017), .B(n5263), .ZN(n8019) );
  MUX2_X1 U9650 ( .A(n8563), .B(n8018), .S(n8019), .Z(n8023) );
  MUX2_X1 U9651 ( .A(n8020), .B(n8534), .S(n8019), .Z(n8021) );
  OAI21_X1 U9652 ( .B1(n8534), .B2(n8167), .A(n8156), .ZN(n8022) );
  NAND2_X1 U9653 ( .A1(n8024), .A2(n10188), .ZN(n8027) );
  INV_X1 U9654 ( .A(n8559), .ZN(n8025) );
  AOI22_X1 U9655 ( .A1(n8025), .A2(n8164), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3152), .ZN(n8026) );
  AND2_X1 U9656 ( .A1(n8027), .A2(n8026), .ZN(n8028) );
  INV_X1 U9657 ( .A(n9539), .ZN(n9572) );
  AND2_X1 U9658 ( .A1(n9739), .A2(n10255), .ZN(n8029) );
  OR2_X1 U9659 ( .A1(n9739), .A2(n10255), .ZN(n8031) );
  NAND2_X1 U9660 ( .A1(n9731), .A2(n9621), .ZN(n9181) );
  INV_X1 U9661 ( .A(n9606), .ZN(n9635) );
  OR2_X1 U9662 ( .A1(n9728), .A2(n9635), .ZN(n9187) );
  NAND2_X1 U9663 ( .A1(n9728), .A2(n9635), .ZN(n9186) );
  NOR2_X1 U9664 ( .A1(n9720), .A2(n9593), .ZN(n8032) );
  INV_X1 U9665 ( .A(n9593), .ZN(n9622) );
  INV_X1 U9666 ( .A(n9720), .ZN(n9603) );
  NAND2_X1 U9667 ( .A1(n9715), .A2(n9573), .ZN(n9093) );
  NAND2_X1 U9668 ( .A1(n9199), .A2(n9093), .ZN(n9591) );
  NOR2_X1 U9669 ( .A1(n9712), .A2(n9592), .ZN(n8033) );
  INV_X1 U9670 ( .A(n9592), .ZN(n9564) );
  NAND2_X1 U9671 ( .A1(n9701), .A2(n9563), .ZN(n9209) );
  NAND2_X1 U9672 ( .A1(n9211), .A2(n9209), .ZN(n9545) );
  INV_X1 U9673 ( .A(n9701), .ZN(n8034) );
  NAND2_X1 U9674 ( .A1(n9698), .A2(n5092), .ZN(n9520) );
  NAND2_X1 U9675 ( .A1(n9520), .A2(n8035), .ZN(n8036) );
  INV_X1 U9676 ( .A(n9540), .ZN(n9510) );
  NAND2_X1 U9677 ( .A1(n8049), .A2(n8968), .ZN(n8038) );
  NOR2_X1 U9678 ( .A1(n8049), .A2(n8968), .ZN(n8037) );
  INV_X1 U9679 ( .A(n9681), .ZN(n8933) );
  NAND2_X1 U9680 ( .A1(n8933), .A2(n9027), .ZN(n8040) );
  NAND2_X1 U9681 ( .A1(n8041), .A2(n8040), .ZN(n9461) );
  NOR2_X1 U9682 ( .A1(n9674), .A2(n9344), .ZN(n9418) );
  INV_X1 U9683 ( .A(n9418), .ZN(n8042) );
  NAND2_X1 U9684 ( .A1(n9674), .A2(n9344), .ZN(n9420) );
  NAND2_X1 U9685 ( .A1(n9671), .A2(n9415), .ZN(n9237) );
  AOI22_X1 U9686 ( .A1(n9671), .A2(n9648), .B1(P1_REG2_REG_27__SCAN_IN), .B2(
        n10362), .ZN(n8055) );
  INV_X1 U9687 ( .A(n8044), .ZN(n9168) );
  INV_X1 U9688 ( .A(n9181), .ZN(n8046) );
  NOR2_X1 U9689 ( .A1(n9634), .A2(n8046), .ZN(n9616) );
  NAND2_X1 U9690 ( .A1(n9187), .A2(n9614), .ZN(n9092) );
  OAI21_X1 U9691 ( .B1(n9616), .B2(n9092), .A(n9186), .ZN(n9604) );
  AND2_X1 U9692 ( .A1(n9720), .A2(n9622), .ZN(n9082) );
  NOR2_X1 U9693 ( .A1(n9604), .A2(n9082), .ZN(n9589) );
  OR2_X1 U9694 ( .A1(n9720), .A2(n9622), .ZN(n9587) );
  NAND2_X1 U9695 ( .A1(n9199), .A2(n9587), .ZN(n9192) );
  OAI21_X1 U9696 ( .B1(n9589), .B2(n9192), .A(n9093), .ZN(n9570) );
  NOR2_X1 U9697 ( .A1(n9712), .A2(n9564), .ZN(n9201) );
  NOR2_X1 U9698 ( .A1(n9201), .A2(n9203), .ZN(n9567) );
  AOI21_X1 U9699 ( .B1(n9570), .B2(n9567), .A(n9203), .ZN(n9561) );
  NAND2_X1 U9700 ( .A1(n9707), .A2(n9572), .ZN(n9055) );
  OAI21_X1 U9701 ( .B1(n9561), .B2(n9274), .A(n9055), .ZN(n9537) );
  INV_X1 U9702 ( .A(n9545), .ZN(n9538) );
  AND2_X1 U9703 ( .A1(n9693), .A2(n9510), .ZN(n9271) );
  NAND2_X1 U9704 ( .A1(n9525), .A2(n9540), .ZN(n9062) );
  NOR2_X1 U9705 ( .A1(n9690), .A2(n8968), .ZN(n9270) );
  NOR2_X1 U9706 ( .A1(n8039), .A2(n9511), .ZN(n9064) );
  NAND2_X1 U9707 ( .A1(n9499), .A2(n9500), .ZN(n9498) );
  INV_X1 U9708 ( .A(n9065), .ZN(n9219) );
  INV_X1 U9709 ( .A(n9231), .ZN(n8047) );
  NAND2_X1 U9710 ( .A1(n9269), .A2(n9467), .ZN(n9069) );
  NAND2_X1 U9711 ( .A1(n9674), .A2(n9481), .ZN(n9268) );
  XNOR2_X1 U9712 ( .A(n9425), .B(n9424), .ZN(n8048) );
  OAI222_X1 U9713 ( .A1(n10350), .A2(n9430), .B1(n10352), .B2(n9481), .C1(
        n8048), .C2(n9620), .ZN(n9669) );
  INV_X1 U9714 ( .A(n9728), .ZN(n9630) );
  NAND2_X1 U9715 ( .A1(n9645), .A2(n9630), .ZN(n9623) );
  INV_X1 U9716 ( .A(n9454), .ZN(n8050) );
  AOI211_X1 U9717 ( .C1(n9671), .C2(n4709), .A(n10388), .B(n8050), .ZN(n9670)
         );
  INV_X1 U9718 ( .A(n9670), .ZN(n8052) );
  INV_X1 U9719 ( .A(n8879), .ZN(n8051) );
  OAI22_X1 U9720 ( .A1(n8052), .A2(n4485), .B1(n9555), .B2(n8051), .ZN(n8053)
         );
  OAI21_X1 U9721 ( .B1(n9669), .B2(n8053), .A(n10366), .ZN(n8054) );
  OAI211_X1 U9722 ( .C1(n9673), .C2(n9633), .A(n8055), .B(n8054), .ZN(P1_U3264) );
  AOI22_X1 U9723 ( .A1(n8057), .A2(n8426), .B1(n10194), .B2(n8056), .ZN(n8061)
         );
  INV_X1 U9724 ( .A(n8058), .ZN(n8060) );
  NOR3_X1 U9725 ( .A1(n8061), .A2(n8060), .A3(n8059), .ZN(n8067) );
  OAI22_X1 U9726 ( .A1(n8167), .A2(n8063), .B1(n6775), .B2(n8062), .ZN(n8066)
         );
  OAI22_X1 U9727 ( .A1(n6041), .A2(n8160), .B1(n8161), .B2(n8064), .ZN(n8065)
         );
  NOR3_X1 U9728 ( .A1(n8067), .A2(n8066), .A3(n8065), .ZN(n8068) );
  OAI21_X1 U9729 ( .B1(n8069), .B2(n8156), .A(n8068), .ZN(P2_U3239) );
  OAI222_X1 U9730 ( .A1(n9774), .A2(n10120), .B1(P1_U3084), .B2(n8071), .C1(
        n8070), .C2(n9773), .ZN(P1_U3325) );
  INV_X1 U9731 ( .A(n8077), .ZN(n8072) );
  INV_X1 U9732 ( .A(n8073), .ZN(n8075) );
  AOI22_X1 U9733 ( .A1(n8408), .A2(n8701), .B1(n10216), .B2(n8409), .ZN(n8572)
         );
  AOI22_X1 U9734 ( .A1(n8575), .A2(n8164), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3152), .ZN(n8078) );
  OAI21_X1 U9735 ( .B1(n8572), .B2(n8150), .A(n8078), .ZN(n8079) );
  AOI21_X1 U9736 ( .B1(n8818), .B2(n8137), .A(n8079), .ZN(n8080) );
  NAND2_X1 U9737 ( .A1(n8082), .A2(n8081), .ZN(n8084) );
  XOR2_X1 U9738 ( .A(n8084), .B(n8083), .Z(n8090) );
  OAI22_X1 U9739 ( .A1(n10199), .A2(n8709), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8085), .ZN(n8088) );
  OAI22_X1 U9740 ( .A1(n8086), .A2(n8160), .B1(n8161), .B2(n8095), .ZN(n8087)
         );
  AOI211_X1 U9741 ( .C1(n8783), .C2(n8137), .A(n8088), .B(n8087), .ZN(n8089)
         );
  OAI21_X1 U9742 ( .B1(n8090), .B2(n8156), .A(n8089), .ZN(P2_U3221) );
  XNOR2_X1 U9743 ( .A(n8091), .B(n8092), .ZN(n8099) );
  INV_X1 U9744 ( .A(n8675), .ZN(n8094) );
  OAI22_X1 U9745 ( .A1(n10199), .A2(n8094), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8093), .ZN(n8097) );
  OAI22_X1 U9746 ( .A1(n8095), .A2(n8160), .B1(n8161), .B2(n8639), .ZN(n8096)
         );
  AOI211_X1 U9747 ( .C1(n8843), .C2(n8137), .A(n8097), .B(n8096), .ZN(n8098)
         );
  OAI21_X1 U9748 ( .B1(n8099), .B2(n8156), .A(n8098), .ZN(P2_U3225) );
  XNOR2_X1 U9749 ( .A(n8101), .B(n8100), .ZN(n8102) );
  NOR2_X1 U9750 ( .A1(n10199), .A2(n8603), .ZN(n8106) );
  AND2_X1 U9751 ( .A1(n8410), .A2(n10216), .ZN(n8103) );
  AOI21_X1 U9752 ( .B1(n8409), .B2(n8701), .A(n8103), .ZN(n8597) );
  OAI22_X1 U9753 ( .A1(n8597), .A2(n8150), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8104), .ZN(n8105) );
  AOI211_X1 U9754 ( .C1(n8828), .C2(n8137), .A(n8106), .B(n8105), .ZN(n8107)
         );
  OAI21_X1 U9755 ( .B1(n8108), .B2(n8156), .A(n8107), .ZN(P2_U3227) );
  OAI21_X1 U9756 ( .B1(n8117), .B2(n8110), .A(n8109), .ZN(n8111) );
  NAND2_X1 U9757 ( .A1(n8111), .A2(n10194), .ZN(n8123) );
  INV_X1 U9758 ( .A(n8112), .ZN(n8114) );
  NAND2_X1 U9759 ( .A1(n8164), .A2(n10437), .ZN(n8113) );
  OAI211_X1 U9760 ( .C1(n8161), .C2(n10428), .A(n8114), .B(n8113), .ZN(n8115)
         );
  AOI21_X1 U9761 ( .B1(n8137), .B2(n8116), .A(n8115), .ZN(n8122) );
  NOR3_X1 U9762 ( .A1(n8142), .A2(n8118), .A3(n8117), .ZN(n8120) );
  OAI21_X1 U9763 ( .B1(n8120), .B2(n8119), .A(n8420), .ZN(n8121) );
  NAND3_X1 U9764 ( .A1(n8123), .A2(n8122), .A3(n8121), .ZN(P2_U3233) );
  XNOR2_X1 U9765 ( .A(n8124), .B(n8125), .ZN(n8130) );
  OAI22_X1 U9766 ( .A1(n10199), .A2(n8690), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9901), .ZN(n8128) );
  OAI22_X1 U9767 ( .A1(n8126), .A2(n8160), .B1(n8161), .B2(n8132), .ZN(n8127)
         );
  AOI211_X1 U9768 ( .C1(n8775), .C2(n8137), .A(n8128), .B(n8127), .ZN(n8129)
         );
  OAI21_X1 U9769 ( .B1(n8130), .B2(n8156), .A(n8129), .ZN(P2_U3235) );
  OAI22_X1 U9770 ( .A1(n8411), .A2(n10427), .B1(n8132), .B2(n10429), .ZN(n8652) );
  AOI22_X1 U9771 ( .A1(n8652), .A2(n10188), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3152), .ZN(n8133) );
  OAI21_X1 U9772 ( .B1(n8657), .B2(n10199), .A(n8133), .ZN(n8136) );
  NOR3_X1 U9773 ( .A1(n8134), .A2(n8639), .A3(n8142), .ZN(n8135) );
  AOI211_X1 U9774 ( .C1(n8137), .C2(n8662), .A(n8136), .B(n8135), .ZN(n8138)
         );
  OAI21_X1 U9775 ( .B1(n8131), .B2(n8156), .A(n8138), .ZN(P2_U3237) );
  INV_X1 U9776 ( .A(n8139), .ZN(n8140) );
  AOI21_X1 U9777 ( .B1(n5628), .B2(n8140), .A(n8156), .ZN(n8147) );
  INV_X1 U9778 ( .A(n8141), .ZN(n8144) );
  NOR3_X1 U9779 ( .A1(n8144), .A2(n8143), .A3(n8142), .ZN(n8146) );
  OAI21_X1 U9780 ( .B1(n8147), .B2(n8146), .A(n8145), .ZN(n8154) );
  INV_X1 U9781 ( .A(n8148), .ZN(n8152) );
  OAI22_X1 U9782 ( .A1(n8150), .A2(n8149), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8496), .ZN(n8151) );
  AOI21_X1 U9783 ( .B1(n8152), .B2(n8164), .A(n8151), .ZN(n8153) );
  OAI211_X1 U9784 ( .C1(n4876), .C2(n8167), .A(n8154), .B(n8153), .ZN(P2_U3240) );
  AOI21_X1 U9785 ( .B1(n8155), .B2(n8157), .A(n8156), .ZN(n8159) );
  NAND2_X1 U9786 ( .A1(n8159), .A2(n8158), .ZN(n8166) );
  NOR2_X1 U9787 ( .A1(n10151), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8163) );
  OAI22_X1 U9788 ( .A1(n8225), .A2(n8161), .B1(n8586), .B2(n8160), .ZN(n8162)
         );
  AOI211_X1 U9789 ( .C1(n8164), .C2(n8590), .A(n8163), .B(n8162), .ZN(n8165)
         );
  OAI211_X1 U9790 ( .C1(n4879), .C2(n8167), .A(n8166), .B(n8165), .ZN(P2_U3242) );
  NOR2_X1 U9791 ( .A1(n8168), .A2(SI_29_), .ZN(n8170) );
  NAND2_X1 U9792 ( .A1(n8168), .A2(SI_29_), .ZN(n8169) );
  MUX2_X1 U9793 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n8185), .Z(n8180) );
  NAND2_X1 U9794 ( .A1(n9110), .A2(n8189), .ZN(n8173) );
  NAND2_X1 U9795 ( .A1(n4479), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n8172) );
  NOR2_X1 U9796 ( .A1(n8529), .A2(n8548), .ZN(n8197) );
  NOR2_X1 U9797 ( .A1(n8526), .A2(n8395), .ZN(n8178) );
  INV_X1 U9798 ( .A(n8178), .ZN(n8179) );
  NAND2_X1 U9799 ( .A1(n9051), .A2(n8189), .ZN(n8175) );
  NAND2_X1 U9800 ( .A1(n5387), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n8174) );
  INV_X1 U9801 ( .A(n8407), .ZN(n8177) );
  NAND2_X1 U9802 ( .A1(n8739), .A2(n8177), .ZN(n8379) );
  INV_X1 U9803 ( .A(n8379), .ZN(n8377) );
  NOR2_X1 U9804 ( .A1(n8545), .A2(n8544), .ZN(n8546) );
  INV_X1 U9805 ( .A(SI_30_), .ZN(n8183) );
  NAND2_X1 U9806 ( .A1(n8181), .A2(n8180), .ZN(n8182) );
  MUX2_X1 U9807 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n8185), .Z(n8186) );
  XNOR2_X1 U9808 ( .A(n8186), .B(SI_31_), .ZN(n8187) );
  NAND2_X1 U9809 ( .A1(n9769), .A2(n8189), .ZN(n8191) );
  NAND2_X1 U9810 ( .A1(n5387), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n8190) );
  INV_X1 U9811 ( .A(n8526), .ZN(n8192) );
  NAND2_X1 U9812 ( .A1(n8529), .A2(n8548), .ZN(n8383) );
  NAND2_X1 U9813 ( .A1(n8388), .A2(n8383), .ZN(n8198) );
  NAND2_X1 U9814 ( .A1(n8810), .A2(n8192), .ZN(n8387) );
  XNOR2_X1 U9815 ( .A(n8194), .B(n10449), .ZN(n8195) );
  INV_X1 U9816 ( .A(n8197), .ZN(n8384) );
  NAND2_X1 U9817 ( .A1(n8387), .A2(n8384), .ZN(n8221) );
  INV_X1 U9818 ( .A(n8221), .ZN(n8219) );
  INV_X1 U9819 ( .A(n8544), .ZN(n8218) );
  INV_X1 U9820 ( .A(n8198), .ZN(n8224) );
  INV_X1 U9821 ( .A(n8640), .ZN(n8355) );
  NAND3_X1 U9822 ( .A1(n10467), .A2(n8398), .A3(n8263), .ZN(n8200) );
  NOR4_X1 U9823 ( .A1(n8200), .A2(n8199), .A3(n6049), .A4(n7112), .ZN(n8204)
         );
  INV_X1 U9824 ( .A(n8201), .ZN(n8203) );
  NAND4_X1 U9825 ( .A1(n8204), .A2(n8203), .A3(n8202), .A4(n8281), .ZN(n8205)
         );
  NOR4_X1 U9826 ( .A1(n8297), .A2(n8205), .A3(n5063), .A4(n6869), .ZN(n8206)
         );
  NAND4_X1 U9827 ( .A1(n10200), .A2(n8208), .A3(n8207), .A4(n8206), .ZN(n8209)
         );
  NOR4_X1 U9828 ( .A1(n8211), .A2(n8210), .A3(n8316), .A4(n8209), .ZN(n8212)
         );
  NAND4_X1 U9829 ( .A1(n8699), .A2(n8325), .A3(n8213), .A4(n8212), .ZN(n8214)
         );
  NOR4_X1 U9830 ( .A1(n8655), .A2(n8666), .A3(n8685), .A4(n8214), .ZN(n8215)
         );
  NAND4_X1 U9831 ( .A1(n8601), .A2(n8355), .A3(n8623), .A4(n8215), .ZN(n8216)
         );
  NOR4_X1 U9832 ( .A1(n8535), .A2(n8569), .A3(n8233), .A4(n8216), .ZN(n8217)
         );
  NAND4_X1 U9833 ( .A1(n8219), .A2(n8218), .A3(n8224), .A4(n8217), .ZN(n8220)
         );
  XNOR2_X1 U9834 ( .A(n8220), .B(n10449), .ZN(n8396) );
  INV_X1 U9835 ( .A(n8385), .ZN(n8222) );
  AOI21_X1 U9836 ( .B1(n8222), .B2(n8383), .A(n8221), .ZN(n8223) );
  NAND2_X1 U9837 ( .A1(n5095), .A2(n4486), .ZN(n8389) );
  MUX2_X1 U9838 ( .A(n8224), .B(n8223), .S(n8389), .Z(n8394) );
  NAND2_X1 U9839 ( .A1(n8818), .A2(n8225), .ZN(n8229) );
  AND2_X1 U9840 ( .A1(n8227), .A2(n8226), .ZN(n8228) );
  INV_X1 U9841 ( .A(n8389), .ZN(n8382) );
  MUX2_X1 U9842 ( .A(n8229), .B(n8228), .S(n8382), .Z(n8376) );
  AND2_X1 U9843 ( .A1(n8369), .A2(n8230), .ZN(n8235) );
  INV_X1 U9844 ( .A(n8231), .ZN(n8232) );
  NOR2_X1 U9845 ( .A1(n8233), .A2(n8232), .ZN(n8234) );
  MUX2_X1 U9846 ( .A(n8235), .B(n8234), .S(n8389), .Z(n8367) );
  AND2_X1 U9847 ( .A1(n8332), .A2(n8236), .ZN(n8237) );
  MUX2_X1 U9848 ( .A(n8238), .B(n8237), .S(n8389), .Z(n8327) );
  INV_X1 U9849 ( .A(n8239), .ZN(n8240) );
  MUX2_X1 U9850 ( .A(n8241), .B(n8240), .S(n8382), .Z(n8242) );
  INV_X1 U9851 ( .A(n8242), .ZN(n8324) );
  NAND2_X1 U9852 ( .A1(n8243), .A2(n8244), .ZN(n8247) );
  INV_X1 U9853 ( .A(n8244), .ZN(n8245) );
  OAI211_X1 U9854 ( .C1(n8245), .C2(n8294), .A(n8306), .B(n8295), .ZN(n8246)
         );
  MUX2_X1 U9855 ( .A(n8247), .B(n8246), .S(n8389), .Z(n8248) );
  INV_X1 U9856 ( .A(n8248), .ZN(n8301) );
  AND2_X1 U9857 ( .A1(n8253), .A2(n8249), .ZN(n8251) );
  OAI211_X1 U9858 ( .C1(n8251), .C2(n8250), .A(n6048), .B(n8257), .ZN(n8252)
         );
  NAND2_X1 U9859 ( .A1(n8252), .A2(n8254), .ZN(n8260) );
  NAND2_X1 U9860 ( .A1(n6048), .A2(n8253), .ZN(n8255) );
  NAND3_X1 U9861 ( .A1(n8256), .A2(n8255), .A3(n8254), .ZN(n8258) );
  NAND2_X1 U9862 ( .A1(n8258), .A2(n8257), .ZN(n8259) );
  MUX2_X1 U9863 ( .A(n8260), .B(n8259), .S(n8382), .Z(n8264) );
  AND2_X1 U9864 ( .A1(n8268), .A2(n8267), .ZN(n8262) );
  AND2_X1 U9865 ( .A1(n8275), .A2(n8274), .ZN(n8261) );
  MUX2_X1 U9866 ( .A(n8262), .B(n8261), .S(n8389), .Z(n8265) );
  NAND3_X1 U9867 ( .A1(n8264), .A2(n8265), .A3(n8263), .ZN(n8272) );
  INV_X1 U9868 ( .A(n8265), .ZN(n8277) );
  AND2_X1 U9869 ( .A1(n8267), .A2(n8266), .ZN(n8269) );
  OAI211_X1 U9870 ( .C1(n8277), .C2(n8269), .A(n8282), .B(n8268), .ZN(n8270)
         );
  NAND2_X1 U9871 ( .A1(n8270), .A2(n8389), .ZN(n8271) );
  NAND2_X1 U9872 ( .A1(n8272), .A2(n8271), .ZN(n8280) );
  AND2_X1 U9873 ( .A1(n8274), .A2(n8273), .ZN(n8276) );
  OAI211_X1 U9874 ( .C1(n8277), .C2(n8276), .A(n8275), .B(n8279), .ZN(n8278)
         );
  AOI22_X1 U9875 ( .A1(n8280), .A2(n8279), .B1(n8382), .B2(n8278), .ZN(n8288)
         );
  OAI21_X1 U9876 ( .B1(n8282), .B2(n8389), .A(n8281), .ZN(n8287) );
  MUX2_X1 U9877 ( .A(n8284), .B(n8283), .S(n8389), .Z(n8285) );
  OAI211_X1 U9878 ( .C1(n8288), .C2(n8287), .A(n8286), .B(n8285), .ZN(n8293)
         );
  MUX2_X1 U9879 ( .A(n8290), .B(n8289), .S(n8389), .Z(n8291) );
  NAND3_X1 U9880 ( .A1(n8293), .A2(n8292), .A3(n8291), .ZN(n8299) );
  NAND3_X1 U9881 ( .A1(n8295), .A2(n8382), .A3(n8294), .ZN(n8296) );
  OAI21_X1 U9882 ( .B1(n8297), .B2(n5063), .A(n8296), .ZN(n8298) );
  NAND2_X1 U9883 ( .A1(n8299), .A2(n8298), .ZN(n8300) );
  NAND2_X1 U9884 ( .A1(n8301), .A2(n8300), .ZN(n8308) );
  NAND2_X1 U9885 ( .A1(n8308), .A2(n8302), .ZN(n8303) );
  NAND3_X1 U9886 ( .A1(n10200), .A2(n8307), .A3(n8303), .ZN(n8305) );
  NAND3_X1 U9887 ( .A1(n8308), .A2(n8307), .A3(n8306), .ZN(n8310) );
  NAND3_X1 U9888 ( .A1(n10200), .A2(n8310), .A3(n8309), .ZN(n8312) );
  MUX2_X1 U9889 ( .A(n8314), .B(n8313), .S(n8389), .Z(n8315) );
  MUX2_X1 U9890 ( .A(n8319), .B(n8318), .S(n8389), .Z(n8320) );
  NAND3_X1 U9891 ( .A1(n8322), .A2(n8321), .A3(n8320), .ZN(n8323) );
  NAND3_X1 U9892 ( .A1(n8325), .A2(n8324), .A3(n8323), .ZN(n8326) );
  NAND2_X1 U9893 ( .A1(n8327), .A2(n8326), .ZN(n8335) );
  NAND2_X1 U9894 ( .A1(n8335), .A2(n8331), .ZN(n8330) );
  INV_X1 U9895 ( .A(n8328), .ZN(n8329) );
  AOI21_X1 U9896 ( .B1(n8333), .B2(n8330), .A(n8329), .ZN(n8339) );
  INV_X1 U9897 ( .A(n8331), .ZN(n8334) );
  OAI211_X1 U9898 ( .C1(n8335), .C2(n8334), .A(n8333), .B(n8332), .ZN(n8337)
         );
  INV_X1 U9899 ( .A(n8350), .ZN(n8336) );
  AOI21_X1 U9900 ( .B1(n8337), .B2(n8683), .A(n8336), .ZN(n8338) );
  MUX2_X1 U9901 ( .A(n8339), .B(n8338), .S(n8382), .Z(n8349) );
  INV_X1 U9902 ( .A(n8340), .ZN(n8343) );
  AND2_X1 U9903 ( .A1(n8342), .A2(n8341), .ZN(n8351) );
  OAI21_X1 U9904 ( .B1(n8349), .B2(n8343), .A(n8351), .ZN(n8348) );
  INV_X1 U9905 ( .A(n8344), .ZN(n8347) );
  INV_X1 U9906 ( .A(n8345), .ZN(n8346) );
  AOI21_X1 U9907 ( .B1(n8351), .B2(n8347), .A(n8346), .ZN(n8354) );
  INV_X1 U9908 ( .A(n8349), .ZN(n8352) );
  NAND3_X1 U9909 ( .A1(n8352), .A2(n8351), .A3(n8350), .ZN(n8353) );
  INV_X1 U9910 ( .A(n8356), .ZN(n8357) );
  OAI21_X1 U9911 ( .B1(n8613), .B2(n8357), .A(n8382), .ZN(n8359) );
  INV_X1 U9912 ( .A(n8360), .ZN(n8358) );
  AOI21_X1 U9913 ( .B1(n8360), .B2(n8612), .A(n8382), .ZN(n8364) );
  INV_X1 U9914 ( .A(n8361), .ZN(n8362) );
  NAND2_X1 U9915 ( .A1(n8362), .A2(n8389), .ZN(n8363) );
  OAI211_X1 U9916 ( .C1(n8365), .C2(n8364), .A(n8601), .B(n8363), .ZN(n8366)
         );
  NAND2_X1 U9917 ( .A1(n8367), .A2(n8366), .ZN(n8374) );
  INV_X1 U9918 ( .A(n8368), .ZN(n8371) );
  INV_X1 U9919 ( .A(n8369), .ZN(n8370) );
  MUX2_X1 U9920 ( .A(n8371), .B(n8370), .S(n8389), .Z(n8372) );
  NOR2_X1 U9921 ( .A1(n8569), .A2(n8372), .ZN(n8373) );
  NAND2_X1 U9922 ( .A1(n8374), .A2(n8373), .ZN(n8375) );
  INV_X1 U9923 ( .A(n8408), .ZN(n8550) );
  NAND3_X1 U9924 ( .A1(n8380), .A2(n8379), .A3(n8378), .ZN(n8381) );
  NAND4_X1 U9925 ( .A1(n8386), .A2(n8385), .A3(n8384), .A4(n8383), .ZN(n8393)
         );
  INV_X1 U9926 ( .A(n8387), .ZN(n8391) );
  INV_X1 U9927 ( .A(n8388), .ZN(n8390) );
  MUX2_X1 U9928 ( .A(n8391), .B(n8390), .S(n8389), .Z(n8392) );
  AOI21_X1 U9929 ( .B1(n8394), .B2(n8393), .A(n8392), .ZN(n8397) );
  NOR4_X1 U9930 ( .A1(n10458), .A2(n10429), .A3(n8401), .A4(n8400), .ZN(n8404)
         );
  OAI21_X1 U9931 ( .B1(n8405), .B2(n8402), .A(P2_B_REG_SCAN_IN), .ZN(n8403) );
  OAI22_X1 U9932 ( .A1(n8406), .A2(n8405), .B1(n8404), .B2(n8403), .ZN(
        P2_U3244) );
  MUX2_X1 U9933 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n8407), .S(P2_U3966), .Z(
        P2_U3581) );
  MUX2_X1 U9934 ( .A(n8408), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8412), .Z(
        P2_U3580) );
  MUX2_X1 U9935 ( .A(n8584), .B(P2_DATAO_REG_27__SCAN_IN), .S(n8412), .Z(
        P2_U3579) );
  MUX2_X1 U9936 ( .A(n8409), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8412), .Z(
        P2_U3578) );
  MUX2_X1 U9937 ( .A(n8618), .B(P2_DATAO_REG_25__SCAN_IN), .S(n8412), .Z(
        P2_U3577) );
  MUX2_X1 U9938 ( .A(n8410), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8412), .Z(
        P2_U3576) );
  INV_X1 U9939 ( .A(n8411), .ZN(n8617) );
  MUX2_X1 U9940 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n8617), .S(P2_U3966), .Z(
        P2_U3575) );
  MUX2_X1 U9941 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8669), .S(P2_U3966), .Z(
        P2_U3574) );
  MUX2_X1 U9942 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8687), .S(P2_U3966), .Z(
        P2_U3573) );
  MUX2_X1 U9943 ( .A(n8702), .B(P2_DATAO_REG_20__SCAN_IN), .S(n8412), .Z(
        P2_U3572) );
  MUX2_X1 U9944 ( .A(n8686), .B(P2_DATAO_REG_19__SCAN_IN), .S(n8412), .Z(
        P2_U3571) );
  MUX2_X1 U9945 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8700), .S(P2_U3966), .Z(
        P2_U3570) );
  MUX2_X1 U9946 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8413), .S(P2_U3966), .Z(
        P2_U3569) );
  MUX2_X1 U9947 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8414), .S(P2_U3966), .Z(
        P2_U3568) );
  MUX2_X1 U9948 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8415), .S(P2_U3966), .Z(
        P2_U3567) );
  MUX2_X1 U9949 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n10218), .S(P2_U3966), .Z(
        P2_U3566) );
  MUX2_X1 U9950 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n8416), .S(P2_U3966), .Z(
        P2_U3565) );
  MUX2_X1 U9951 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n10217), .S(P2_U3966), .Z(
        P2_U3564) );
  MUX2_X1 U9952 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n8417), .S(P2_U3966), .Z(
        P2_U3563) );
  MUX2_X1 U9953 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n8418), .S(P2_U3966), .Z(
        P2_U3562) );
  MUX2_X1 U9954 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n8419), .S(P2_U3966), .Z(
        P2_U3561) );
  MUX2_X1 U9955 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n8420), .S(P2_U3966), .Z(
        P2_U3560) );
  MUX2_X1 U9956 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n8421), .S(P2_U3966), .Z(
        P2_U3559) );
  MUX2_X1 U9957 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n8422), .S(P2_U3966), .Z(
        P2_U3558) );
  MUX2_X1 U9958 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n8423), .S(P2_U3966), .Z(
        P2_U3557) );
  MUX2_X1 U9959 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n8424), .S(P2_U3966), .Z(
        P2_U3556) );
  MUX2_X1 U9960 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n8425), .S(P2_U3966), .Z(
        P2_U3555) );
  MUX2_X1 U9961 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n6179), .S(P2_U3966), .Z(
        P2_U3554) );
  MUX2_X1 U9962 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n8426), .S(P2_U3966), .Z(
        P2_U3553) );
  MUX2_X1 U9963 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n6047), .S(P2_U3966), .Z(
        P2_U3552) );
  NAND2_X1 U9964 ( .A1(n8491), .A2(n8427), .ZN(n8439) );
  NOR2_X1 U9965 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5283), .ZN(n8428) );
  AOI21_X1 U9966 ( .B1(n10404), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n8428), .ZN(
        n8438) );
  XOR2_X1 U9967 ( .A(n8430), .B(n8429), .Z(n8431) );
  NAND2_X1 U9968 ( .A1(n10403), .A2(n8431), .ZN(n8437) );
  INV_X1 U9969 ( .A(n8432), .ZN(n8433) );
  OAI211_X1 U9970 ( .C1(n8435), .C2(n8434), .A(n10402), .B(n8433), .ZN(n8436)
         );
  NAND4_X1 U9971 ( .A1(n8439), .A2(n8438), .A3(n8437), .A4(n8436), .ZN(
        P2_U3248) );
  NAND2_X1 U9972 ( .A1(n8491), .A2(n8440), .ZN(n8453) );
  OAI211_X1 U9973 ( .C1(n8443), .C2(n8442), .A(n10403), .B(n8441), .ZN(n8452)
         );
  INV_X1 U9974 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n8444) );
  NOR2_X1 U9975 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8444), .ZN(n8445) );
  AOI21_X1 U9976 ( .B1(n10404), .B2(P2_ADDR_REG_12__SCAN_IN), .A(n8445), .ZN(
        n8451) );
  OAI21_X1 U9977 ( .B1(n8448), .B2(n8447), .A(n8446), .ZN(n8449) );
  NAND2_X1 U9978 ( .A1(n10402), .A2(n8449), .ZN(n8450) );
  NAND4_X1 U9979 ( .A1(n8453), .A2(n8452), .A3(n8451), .A4(n8450), .ZN(
        P2_U3257) );
  NOR2_X1 U9980 ( .A1(n8455), .A2(n8454), .ZN(n8457) );
  XOR2_X1 U9981 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n8480), .Z(n8458) );
  NAND2_X1 U9982 ( .A1(n8458), .A2(n8459), .ZN(n8481) );
  OAI21_X1 U9983 ( .B1(n8459), .B2(n8458), .A(n8481), .ZN(n8460) );
  NAND2_X1 U9984 ( .A1(n8460), .A2(n10402), .ZN(n8473) );
  NOR2_X1 U9985 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8461), .ZN(n8462) );
  AOI21_X1 U9986 ( .B1(n10404), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n8462), .ZN(
        n8472) );
  NOR2_X1 U9987 ( .A1(n8464), .A2(n8463), .ZN(n8466) );
  NOR2_X1 U9988 ( .A1(n8466), .A2(n8465), .ZN(n8469) );
  MUX2_X1 U9989 ( .A(n5532), .B(P2_REG2_REG_16__SCAN_IN), .S(n8480), .Z(n8467)
         );
  INV_X1 U9990 ( .A(n8467), .ZN(n8468) );
  NAND2_X1 U9991 ( .A1(n8468), .A2(n8469), .ZN(n8474) );
  OAI211_X1 U9992 ( .C1(n8469), .C2(n8468), .A(n10403), .B(n8474), .ZN(n8471)
         );
  NAND2_X1 U9993 ( .A1(n8491), .A2(n8480), .ZN(n8470) );
  NAND4_X1 U9994 ( .A1(n8473), .A2(n8472), .A3(n8471), .A4(n8470), .ZN(
        P2_U3261) );
  NAND2_X1 U9995 ( .A1(n8480), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n8475) );
  NAND2_X1 U9996 ( .A1(n8475), .A2(n8474), .ZN(n8477) );
  XNOR2_X1 U9997 ( .A(n8493), .B(P2_REG2_REG_17__SCAN_IN), .ZN(n8476) );
  NAND2_X1 U9998 ( .A1(n8476), .A2(n8477), .ZN(n8492) );
  OAI211_X1 U9999 ( .C1(n8477), .C2(n8476), .A(n10403), .B(n8492), .ZN(n8490)
         );
  NOR2_X1 U10000 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8478), .ZN(n8479) );
  AOI21_X1 U10001 ( .B1(n10404), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n8479), .ZN(
        n8489) );
  OR2_X1 U10002 ( .A1(n10406), .A2(n8493), .ZN(n8488) );
  OR2_X1 U10003 ( .A1(n8480), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n8482) );
  NAND2_X1 U10004 ( .A1(n8482), .A2(n8481), .ZN(n8485) );
  INV_X1 U10005 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8483) );
  XNOR2_X1 U10006 ( .A(n8493), .B(n8483), .ZN(n8484) );
  NOR2_X1 U10007 ( .A1(n8484), .A2(n8485), .ZN(n8498) );
  AOI21_X1 U10008 ( .B1(n8485), .B2(n8484), .A(n8498), .ZN(n8486) );
  NAND2_X1 U10009 ( .A1(n10402), .A2(n8486), .ZN(n8487) );
  NAND4_X1 U10010 ( .A1(n8490), .A2(n8489), .A3(n8488), .A4(n8487), .ZN(
        P2_U3262) );
  NAND2_X1 U10011 ( .A1(n8491), .A2(n8512), .ZN(n8506) );
  OAI21_X1 U10012 ( .B1(n8494), .B2(n8493), .A(n8492), .ZN(n8507) );
  XOR2_X1 U10013 ( .A(n8507), .B(n8512), .Z(n8495) );
  NAND2_X1 U10014 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n8495), .ZN(n8509) );
  OAI211_X1 U10015 ( .C1(P2_REG2_REG_18__SCAN_IN), .C2(n8495), .A(n10403), .B(
        n8509), .ZN(n8505) );
  NOR2_X1 U10016 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8496), .ZN(n8497) );
  AOI21_X1 U10017 ( .B1(n10404), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n8497), .ZN(
        n8504) );
  INV_X1 U10018 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8789) );
  XNOR2_X1 U10019 ( .A(n8512), .B(n8789), .ZN(n8501) );
  OAI21_X1 U10020 ( .B1(n8501), .B2(n8500), .A(n8511), .ZN(n8502) );
  NAND2_X1 U10021 ( .A1(n10402), .A2(n8502), .ZN(n8503) );
  NAND4_X1 U10022 ( .A1(n8506), .A2(n8505), .A3(n8504), .A4(n8503), .ZN(
        P2_U3263) );
  NAND2_X1 U10023 ( .A1(n8512), .A2(n8507), .ZN(n8508) );
  NAND2_X1 U10024 ( .A1(n8509), .A2(n8508), .ZN(n8510) );
  XOR2_X1 U10025 ( .A(n8510), .B(P2_REG2_REG_19__SCAN_IN), .Z(n8516) );
  INV_X1 U10026 ( .A(n8516), .ZN(n8514) );
  INV_X1 U10027 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8784) );
  OAI21_X1 U10028 ( .B1(n8515), .B2(n10407), .A(n10406), .ZN(n8513) );
  AOI21_X1 U10029 ( .B1(n10403), .B2(n8514), .A(n8513), .ZN(n8519) );
  AOI22_X1 U10030 ( .A1(n8516), .A2(n10403), .B1(n10402), .B2(n8515), .ZN(
        n8518) );
  MUX2_X1 U10031 ( .A(n8519), .B(n8518), .S(n8517), .Z(n8521) );
  NAND2_X1 U10032 ( .A1(n10404), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n8520) );
  OAI211_X1 U10033 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n8085), .A(n8521), .B(
        n8520), .ZN(P2_U3264) );
  XNOR2_X1 U10034 ( .A(n8810), .B(n8530), .ZN(n8522) );
  NAND2_X1 U10035 ( .A1(n8523), .A2(P2_B_REG_SCAN_IN), .ZN(n8524) );
  NAND2_X1 U10036 ( .A1(n8701), .A2(n8524), .ZN(n8549) );
  INV_X1 U10037 ( .A(n8549), .ZN(n8525) );
  NAND2_X1 U10038 ( .A1(n8526), .A2(n8525), .ZN(n8733) );
  NOR2_X1 U10039 ( .A1(n10456), .A2(n8733), .ZN(n8532) );
  AOI21_X1 U10040 ( .B1(n10456), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8532), .ZN(
        n8528) );
  NAND2_X1 U10041 ( .A1(n8810), .A2(n10228), .ZN(n8527) );
  OAI211_X1 U10042 ( .C1(n8730), .C2(n10206), .A(n8528), .B(n8527), .ZN(
        P2_U3265) );
  OAI211_X1 U10043 ( .C1(n4583), .C2(n4584), .A(n10418), .B(n8530), .ZN(n8734)
         );
  NOR2_X1 U10044 ( .A1(n4583), .A2(n10439), .ZN(n8531) );
  AOI211_X1 U10045 ( .C1(n10456), .C2(P2_REG2_REG_30__SCAN_IN), .A(n8532), .B(
        n8531), .ZN(n8533) );
  OAI21_X1 U10046 ( .B1(n10206), .B2(n8734), .A(n8533), .ZN(P2_U3266) );
  AOI22_X1 U10047 ( .A1(n8536), .A2(n8535), .B1(n8550), .B2(n8534), .ZN(n8537)
         );
  AOI211_X1 U10048 ( .C1(n8739), .C2(n8538), .A(n10472), .B(n4584), .ZN(n8738)
         );
  INV_X1 U10049 ( .A(n8739), .ZN(n8539) );
  NOR2_X1 U10050 ( .A1(n8539), .A2(n10439), .ZN(n8543) );
  OAI22_X1 U10051 ( .A1(n8541), .A2(n10208), .B1(n8540), .B2(n10211), .ZN(
        n8542) );
  AOI211_X1 U10052 ( .C1(n8738), .C2(n10422), .A(n8543), .B(n8542), .ZN(n8555)
         );
  INV_X1 U10053 ( .A(n8551), .ZN(n8552) );
  NAND2_X1 U10054 ( .A1(n8737), .A2(n10211), .ZN(n8554) );
  OAI211_X1 U10055 ( .C1(n8741), .C2(n8717), .A(n8555), .B(n8554), .ZN(
        P2_U3267) );
  INV_X1 U10056 ( .A(n8556), .ZN(n8557) );
  NAND2_X1 U10057 ( .A1(n8557), .A2(n8723), .ZN(n8565) );
  OAI22_X1 U10058 ( .A1(n8559), .A2(n10208), .B1(n8558), .B2(n10211), .ZN(
        n8562) );
  NOR2_X1 U10059 ( .A1(n8560), .A2(n10206), .ZN(n8561) );
  AOI211_X1 U10060 ( .C1(n10228), .C2(n8563), .A(n8562), .B(n8561), .ZN(n8564)
         );
  OAI211_X1 U10061 ( .C1(n10456), .C2(n8566), .A(n8565), .B(n8564), .ZN(
        P2_U3268) );
  XNOR2_X1 U10062 ( .A(n8567), .B(n8569), .ZN(n8820) );
  NAND2_X1 U10063 ( .A1(n8568), .A2(n8569), .ZN(n8570) );
  NAND3_X1 U10064 ( .A1(n8571), .A2(n10432), .A3(n8570), .ZN(n8573) );
  NAND2_X1 U10065 ( .A1(n8573), .A2(n8572), .ZN(n8743) );
  INV_X1 U10066 ( .A(n8818), .ZN(n8578) );
  AOI211_X1 U10067 ( .C1(n8818), .C2(n8589), .A(n10472), .B(n8574), .ZN(n8742)
         );
  NAND2_X1 U10068 ( .A1(n8742), .A2(n10422), .ZN(n8577) );
  AOI22_X1 U10069 ( .A1(n8575), .A2(n10447), .B1(P2_REG2_REG_27__SCAN_IN), 
        .B2(n10456), .ZN(n8576) );
  OAI211_X1 U10070 ( .C1(n8578), .C2(n10439), .A(n8577), .B(n8576), .ZN(n8579)
         );
  AOI21_X1 U10071 ( .B1(n8743), .B2(n10211), .A(n8579), .ZN(n8580) );
  OAI21_X1 U10072 ( .B1(n8820), .B2(n8717), .A(n8580), .ZN(P2_U3269) );
  XNOR2_X1 U10073 ( .A(n8581), .B(n8582), .ZN(n8825) );
  XNOR2_X1 U10074 ( .A(n8583), .B(n8582), .ZN(n8588) );
  NAND2_X1 U10075 ( .A1(n8584), .A2(n8701), .ZN(n8585) );
  OAI21_X1 U10076 ( .B1(n8586), .B2(n10429), .A(n8585), .ZN(n8587) );
  AOI21_X1 U10077 ( .B1(n8588), .B2(n10432), .A(n8587), .ZN(n8747) );
  INV_X1 U10078 ( .A(n8747), .ZN(n8594) );
  OAI211_X1 U10079 ( .C1(n4879), .C2(n4880), .A(n8589), .B(n10418), .ZN(n8746)
         );
  AOI22_X1 U10080 ( .A1(n8590), .A2(n10447), .B1(n10456), .B2(
        P2_REG2_REG_26__SCAN_IN), .ZN(n8592) );
  NAND2_X1 U10081 ( .A1(n8823), .A2(n10228), .ZN(n8591) );
  OAI211_X1 U10082 ( .C1(n8746), .C2(n8607), .A(n8592), .B(n8591), .ZN(n8593)
         );
  AOI21_X1 U10083 ( .B1(n8594), .B2(n10211), .A(n8593), .ZN(n8595) );
  OAI21_X1 U10084 ( .B1(n8825), .B2(n8717), .A(n8595), .ZN(P2_U3270) );
  XNOR2_X1 U10085 ( .A(n8596), .B(n4901), .ZN(n8599) );
  INV_X1 U10086 ( .A(n8597), .ZN(n8598) );
  AOI21_X1 U10087 ( .B1(n8599), .B2(n10432), .A(n8598), .ZN(n8751) );
  XOR2_X1 U10088 ( .A(n8601), .B(n8600), .Z(n8830) );
  INV_X1 U10089 ( .A(n8830), .ZN(n8602) );
  NAND2_X1 U10090 ( .A1(n8602), .A2(n8723), .ZN(n8611) );
  OAI22_X1 U10091 ( .A1(n10211), .A2(n8604), .B1(n8603), .B2(n10208), .ZN(
        n8609) );
  INV_X1 U10092 ( .A(n8627), .ZN(n8606) );
  OAI211_X1 U10093 ( .C1(n4904), .C2(n8606), .A(n10418), .B(n8605), .ZN(n8750)
         );
  NOR2_X1 U10094 ( .A1(n8750), .A2(n8607), .ZN(n8608) );
  AOI211_X1 U10095 ( .C1(n10228), .C2(n8828), .A(n8609), .B(n8608), .ZN(n8610)
         );
  OAI211_X1 U10096 ( .C1(n10456), .C2(n8751), .A(n8611), .B(n8610), .ZN(
        P2_U3271) );
  NAND2_X1 U10097 ( .A1(n8633), .A2(n8612), .ZN(n8614) );
  NAND2_X1 U10098 ( .A1(n8614), .A2(n8613), .ZN(n8616) );
  NAND3_X1 U10099 ( .A1(n8616), .A2(n8615), .A3(n10432), .ZN(n8620) );
  AOI22_X1 U10100 ( .A1(n8618), .A2(n8701), .B1(n8617), .B2(n10216), .ZN(n8619) );
  AOI21_X1 U10101 ( .B1(n8623), .B2(n8622), .A(n8621), .ZN(n8835) );
  INV_X1 U10102 ( .A(n8835), .ZN(n8624) );
  NAND2_X1 U10103 ( .A1(n8624), .A2(n8723), .ZN(n8632) );
  OAI22_X1 U10104 ( .A1(n10211), .A2(n8626), .B1(n8625), .B2(n10208), .ZN(
        n8630) );
  OAI211_X1 U10105 ( .C1(n8628), .C2(n8642), .A(n10418), .B(n8627), .ZN(n8754)
         );
  NOR2_X1 U10106 ( .A1(n8754), .A2(n10206), .ZN(n8629) );
  AOI211_X1 U10107 ( .C1(n10228), .C2(n8833), .A(n8630), .B(n8629), .ZN(n8631)
         );
  OAI211_X1 U10108 ( .C1(n10456), .C2(n8755), .A(n8632), .B(n8631), .ZN(
        P2_U3272) );
  INV_X1 U10109 ( .A(n8633), .ZN(n8634) );
  AOI21_X1 U10110 ( .B1(n8635), .B2(n8640), .A(n8634), .ZN(n8636) );
  OAI222_X1 U10111 ( .A1(n10429), .A2(n8639), .B1(n10427), .B2(n8638), .C1(
        n8637), .C2(n8636), .ZN(n8758) );
  INV_X1 U10112 ( .A(n8758), .ZN(n8649) );
  OR2_X1 U10113 ( .A1(n8641), .A2(n8640), .ZN(n8762) );
  NAND3_X1 U10114 ( .A1(n8762), .A2(n8761), .A3(n8723), .ZN(n8648) );
  AOI211_X1 U10115 ( .C1(n8760), .C2(n8659), .A(n10472), .B(n8642), .ZN(n8759)
         );
  AOI22_X1 U10116 ( .A1(n10456), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n8643), 
        .B2(n10447), .ZN(n8644) );
  OAI21_X1 U10117 ( .B1(n8645), .B2(n10439), .A(n8644), .ZN(n8646) );
  AOI21_X1 U10118 ( .B1(n8759), .B2(n10422), .A(n8646), .ZN(n8647) );
  OAI211_X1 U10119 ( .C1(n10456), .C2(n8649), .A(n8648), .B(n8647), .ZN(
        P2_U3273) );
  INV_X1 U10120 ( .A(n8655), .ZN(n8651) );
  XNOR2_X1 U10121 ( .A(n8650), .B(n8651), .ZN(n8653) );
  AOI21_X1 U10122 ( .B1(n8653), .B2(n10432), .A(n8652), .ZN(n8766) );
  XOR2_X1 U10123 ( .A(n8655), .B(n8654), .Z(n8840) );
  INV_X1 U10124 ( .A(n8840), .ZN(n8656) );
  NAND2_X1 U10125 ( .A1(n8656), .A2(n8723), .ZN(n8664) );
  OAI22_X1 U10126 ( .A1(n10211), .A2(n8658), .B1(n8657), .B2(n10208), .ZN(
        n8661) );
  OAI211_X1 U10127 ( .C1(n8767), .C2(n8674), .A(n10418), .B(n8659), .ZN(n8765)
         );
  NOR2_X1 U10128 ( .A1(n8765), .A2(n10206), .ZN(n8660) );
  AOI211_X1 U10129 ( .C1(n10228), .C2(n8662), .A(n8661), .B(n8660), .ZN(n8663)
         );
  OAI211_X1 U10130 ( .C1(n10456), .C2(n8766), .A(n8664), .B(n8663), .ZN(
        P2_U3274) );
  XOR2_X1 U10131 ( .A(n8665), .B(n8666), .Z(n8846) );
  XNOR2_X1 U10132 ( .A(n8667), .B(n8666), .ZN(n8668) );
  NAND2_X1 U10133 ( .A1(n8668), .A2(n10432), .ZN(n8671) );
  AOI22_X1 U10134 ( .A1(n8669), .A2(n8701), .B1(n10216), .B2(n8702), .ZN(n8670) );
  NAND2_X1 U10135 ( .A1(n8671), .A2(n8670), .ZN(n8771) );
  NAND2_X1 U10136 ( .A1(n8843), .A2(n4502), .ZN(n8672) );
  NAND2_X1 U10137 ( .A1(n8672), .A2(n10418), .ZN(n8673) );
  NOR2_X1 U10138 ( .A1(n8674), .A2(n8673), .ZN(n8770) );
  NAND2_X1 U10139 ( .A1(n8770), .A2(n10422), .ZN(n8677) );
  AOI22_X1 U10140 ( .A1(n10456), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8675), 
        .B2(n10447), .ZN(n8676) );
  OAI211_X1 U10141 ( .C1(n8678), .C2(n10439), .A(n8677), .B(n8676), .ZN(n8679)
         );
  AOI21_X1 U10142 ( .B1(n8771), .B2(n10211), .A(n8679), .ZN(n8680) );
  OAI21_X1 U10143 ( .B1(n8846), .B2(n8717), .A(n8680), .ZN(P2_U3275) );
  XNOR2_X1 U10144 ( .A(n8681), .B(n8685), .ZN(n8849) );
  NAND2_X1 U10145 ( .A1(n8682), .A2(n8683), .ZN(n8684) );
  XOR2_X1 U10146 ( .A(n8685), .B(n8684), .Z(n8688) );
  AOI222_X1 U10147 ( .A1(n10432), .A2(n8688), .B1(n8687), .B2(n8701), .C1(
        n8686), .C2(n10216), .ZN(n8778) );
  INV_X1 U10148 ( .A(n8778), .ZN(n8695) );
  NAND2_X1 U10149 ( .A1(n8706), .A2(n8775), .ZN(n8689) );
  NAND3_X1 U10150 ( .A1(n4502), .A2(n10418), .A3(n8689), .ZN(n8777) );
  OAI22_X1 U10151 ( .A1(n10211), .A2(n8691), .B1(n8690), .B2(n10208), .ZN(
        n8692) );
  AOI21_X1 U10152 ( .B1(n8775), .B2(n10228), .A(n8692), .ZN(n8693) );
  OAI21_X1 U10153 ( .B1(n8777), .B2(n10206), .A(n8693), .ZN(n8694) );
  AOI21_X1 U10154 ( .B1(n8695), .B2(n10211), .A(n8694), .ZN(n8696) );
  OAI21_X1 U10155 ( .B1(n8849), .B2(n8717), .A(n8696), .ZN(P2_U3276) );
  XOR2_X1 U10156 ( .A(n8697), .B(n8699), .Z(n8856) );
  OAI21_X1 U10157 ( .B1(n8699), .B2(n8698), .A(n8682), .ZN(n8703) );
  AOI222_X1 U10158 ( .A1(n10432), .A2(n8703), .B1(n8702), .B2(n8701), .C1(
        n8700), .C2(n10216), .ZN(n8704) );
  INV_X1 U10159 ( .A(n8704), .ZN(n8781) );
  INV_X1 U10160 ( .A(n8706), .ZN(n8707) );
  AOI211_X1 U10161 ( .C1(n8783), .C2(n4878), .A(n10472), .B(n8707), .ZN(n8782)
         );
  NAND2_X1 U10162 ( .A1(n8782), .A2(n8708), .ZN(n8712) );
  INV_X1 U10163 ( .A(n8709), .ZN(n8710) );
  AOI22_X1 U10164 ( .A1(n10456), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n8710), 
        .B2(n10447), .ZN(n8711) );
  OAI211_X1 U10165 ( .C1(n8713), .C2(n10439), .A(n8712), .B(n8711), .ZN(n8714)
         );
  AOI21_X1 U10166 ( .B1(n8781), .B2(n10211), .A(n8714), .ZN(n8716) );
  OAI21_X1 U10167 ( .B1(n8856), .B2(n8717), .A(n8716), .ZN(P2_U3277) );
  NAND2_X1 U10168 ( .A1(n8718), .A2(n10211), .ZN(n8729) );
  OAI22_X1 U10169 ( .A1(n10211), .A2(n8720), .B1(n8719), .B2(n10208), .ZN(
        n8721) );
  AOI21_X1 U10170 ( .B1(n10228), .B2(n8722), .A(n8721), .ZN(n8728) );
  NAND2_X1 U10171 ( .A1(n8724), .A2(n8723), .ZN(n8727) );
  NAND2_X1 U10172 ( .A1(n8725), .A2(n10422), .ZN(n8726) );
  NAND4_X1 U10173 ( .A1(n8729), .A2(n8728), .A3(n8727), .A4(n8726), .ZN(
        P2_U3285) );
  NAND2_X1 U10174 ( .A1(n8730), .A2(n8733), .ZN(n8808) );
  MUX2_X1 U10175 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n8808), .S(n10499), .Z(
        n8731) );
  INV_X1 U10176 ( .A(n8732), .ZN(P2_U3551) );
  AND2_X1 U10177 ( .A1(n8734), .A2(n8733), .ZN(n8813) );
  INV_X1 U10178 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n8735) );
  MUX2_X1 U10179 ( .A(n8813), .B(n8735), .S(n10504), .Z(n8736) );
  OAI21_X1 U10180 ( .B1(n4583), .B2(n8776), .A(n8736), .ZN(P2_U3550) );
  OAI21_X1 U10181 ( .B1(n8741), .B2(n10466), .A(n8740), .ZN(n8815) );
  MUX2_X1 U10182 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n8815), .S(n10499), .Z(
        P2_U3549) );
  MUX2_X1 U10183 ( .A(n8816), .B(P2_REG1_REG_27__SCAN_IN), .S(n10504), .Z(
        n8744) );
  AOI21_X1 U10184 ( .B1(n8773), .B2(n8818), .A(n8744), .ZN(n8745) );
  OAI21_X1 U10185 ( .B1(n8820), .B2(n8791), .A(n8745), .ZN(P2_U3547) );
  NAND2_X1 U10186 ( .A1(n8747), .A2(n8746), .ZN(n8821) );
  MUX2_X1 U10187 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n8821), .S(n10499), .Z(
        n8748) );
  AOI21_X1 U10188 ( .B1(n8773), .B2(n8823), .A(n8748), .ZN(n8749) );
  OAI21_X1 U10189 ( .B1(n8825), .B2(n8791), .A(n8749), .ZN(P2_U3546) );
  NAND2_X1 U10190 ( .A1(n8751), .A2(n8750), .ZN(n8826) );
  MUX2_X1 U10191 ( .A(n8826), .B(P2_REG1_REG_25__SCAN_IN), .S(n10504), .Z(
        n8752) );
  AOI21_X1 U10192 ( .B1(n8773), .B2(n8828), .A(n8752), .ZN(n8753) );
  OAI21_X1 U10193 ( .B1(n8830), .B2(n8791), .A(n8753), .ZN(P2_U3545) );
  NAND2_X1 U10194 ( .A1(n8755), .A2(n8754), .ZN(n8831) );
  MUX2_X1 U10195 ( .A(n8831), .B(P2_REG1_REG_24__SCAN_IN), .S(n10504), .Z(
        n8756) );
  AOI21_X1 U10196 ( .B1(n8773), .B2(n8833), .A(n8756), .ZN(n8757) );
  OAI21_X1 U10197 ( .B1(n8835), .B2(n8791), .A(n8757), .ZN(P2_U3544) );
  AOI211_X1 U10198 ( .C1(n8803), .C2(n8760), .A(n8759), .B(n8758), .ZN(n8764)
         );
  NAND3_X1 U10199 ( .A1(n8762), .A2(n8761), .A3(n10485), .ZN(n8763) );
  NAND2_X1 U10200 ( .A1(n8764), .A2(n8763), .ZN(n8836) );
  MUX2_X1 U10201 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n8836), .S(n10499), .Z(
        P2_U3543) );
  OAI211_X1 U10202 ( .C1(n8767), .C2(n10488), .A(n8766), .B(n8765), .ZN(n8837)
         );
  MUX2_X1 U10203 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n8837), .S(n10499), .Z(
        n8768) );
  INV_X1 U10204 ( .A(n8768), .ZN(n8769) );
  OAI21_X1 U10205 ( .B1(n8840), .B2(n8791), .A(n8769), .ZN(P2_U3542) );
  OR2_X1 U10206 ( .A1(n8771), .A2(n8770), .ZN(n8841) );
  MUX2_X1 U10207 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n8841), .S(n10499), .Z(
        n8772) );
  AOI21_X1 U10208 ( .B1(n8773), .B2(n8843), .A(n8772), .ZN(n8774) );
  OAI21_X1 U10209 ( .B1(n8846), .B2(n8791), .A(n8774), .ZN(P2_U3541) );
  INV_X1 U10210 ( .A(n8775), .ZN(n8848) );
  OAI22_X1 U10211 ( .A1(n8849), .A2(n8791), .B1(n8848), .B2(n8776), .ZN(n8780)
         );
  NAND2_X1 U10212 ( .A1(n8778), .A2(n8777), .ZN(n8850) );
  MUX2_X1 U10213 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n8850), .S(n10499), .Z(
        n8779) );
  OR2_X1 U10214 ( .A1(n8780), .A2(n8779), .ZN(P2_U3540) );
  AOI211_X1 U10215 ( .C1(n8803), .C2(n8783), .A(n8782), .B(n8781), .ZN(n8853)
         );
  MUX2_X1 U10216 ( .A(n8784), .B(n8853), .S(n10499), .Z(n8785) );
  OAI21_X1 U10217 ( .B1(n8856), .B2(n8791), .A(n8785), .ZN(P2_U3539) );
  AOI211_X1 U10218 ( .C1(n8803), .C2(n8788), .A(n8787), .B(n8786), .ZN(n8857)
         );
  MUX2_X1 U10219 ( .A(n8789), .B(n8857), .S(n10499), .Z(n8790) );
  OAI21_X1 U10220 ( .B1(n8861), .B2(n8791), .A(n8790), .ZN(P2_U3538) );
  AOI211_X1 U10221 ( .C1(n8803), .C2(n8794), .A(n8793), .B(n8792), .ZN(n8795)
         );
  OAI21_X1 U10222 ( .B1(n8796), .B2(n10466), .A(n8795), .ZN(n8862) );
  MUX2_X1 U10223 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n8862), .S(n10499), .Z(
        P2_U3537) );
  AOI211_X1 U10224 ( .C1(n8803), .C2(n8799), .A(n8798), .B(n8797), .ZN(n8800)
         );
  OAI21_X1 U10225 ( .B1(n8801), .B2(n10466), .A(n8800), .ZN(n8863) );
  MUX2_X1 U10226 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n8863), .S(n10499), .Z(
        P2_U3536) );
  NAND2_X1 U10227 ( .A1(n8802), .A2(n10485), .ZN(n8807) );
  NAND2_X1 U10228 ( .A1(n8804), .A2(n8803), .ZN(n10191) );
  NAND4_X1 U10229 ( .A1(n8807), .A2(n8806), .A3(n10191), .A4(n8805), .ZN(n8864) );
  MUX2_X1 U10230 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n8864), .S(n10499), .Z(
        P2_U3535) );
  MUX2_X1 U10231 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n8808), .S(n10496), .Z(
        n8809) );
  INV_X1 U10232 ( .A(n8811), .ZN(P2_U3519) );
  INV_X1 U10233 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n8812) );
  MUX2_X1 U10234 ( .A(n8813), .B(n8812), .S(n10494), .Z(n8814) );
  OAI21_X1 U10235 ( .B1(n4583), .B2(n8847), .A(n8814), .ZN(P2_U3518) );
  MUX2_X1 U10236 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n8815), .S(n10496), .Z(
        P2_U3517) );
  MUX2_X1 U10237 ( .A(n8816), .B(P2_REG0_REG_27__SCAN_IN), .S(n10494), .Z(
        n8817) );
  AOI21_X1 U10238 ( .B1(n8844), .B2(n8818), .A(n8817), .ZN(n8819) );
  OAI21_X1 U10239 ( .B1(n8820), .B2(n8860), .A(n8819), .ZN(P2_U3515) );
  MUX2_X1 U10240 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n8821), .S(n10496), .Z(
        n8822) );
  AOI21_X1 U10241 ( .B1(n8844), .B2(n8823), .A(n8822), .ZN(n8824) );
  OAI21_X1 U10242 ( .B1(n8825), .B2(n8860), .A(n8824), .ZN(P2_U3514) );
  MUX2_X1 U10243 ( .A(n8826), .B(P2_REG0_REG_25__SCAN_IN), .S(n10494), .Z(
        n8827) );
  AOI21_X1 U10244 ( .B1(n8844), .B2(n8828), .A(n8827), .ZN(n8829) );
  OAI21_X1 U10245 ( .B1(n8830), .B2(n8860), .A(n8829), .ZN(P2_U3513) );
  MUX2_X1 U10246 ( .A(n8831), .B(P2_REG0_REG_24__SCAN_IN), .S(n10494), .Z(
        n8832) );
  AOI21_X1 U10247 ( .B1(n8844), .B2(n8833), .A(n8832), .ZN(n8834) );
  OAI21_X1 U10248 ( .B1(n8835), .B2(n8860), .A(n8834), .ZN(P2_U3512) );
  MUX2_X1 U10249 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n8836), .S(n10496), .Z(
        P2_U3511) );
  MUX2_X1 U10250 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n8837), .S(n10496), .Z(
        n8838) );
  INV_X1 U10251 ( .A(n8838), .ZN(n8839) );
  OAI21_X1 U10252 ( .B1(n8840), .B2(n8860), .A(n8839), .ZN(P2_U3510) );
  MUX2_X1 U10253 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n8841), .S(n10496), .Z(
        n8842) );
  AOI21_X1 U10254 ( .B1(n8844), .B2(n8843), .A(n8842), .ZN(n8845) );
  OAI21_X1 U10255 ( .B1(n8846), .B2(n8860), .A(n8845), .ZN(P2_U3509) );
  OAI22_X1 U10256 ( .A1(n8849), .A2(n8860), .B1(n8848), .B2(n8847), .ZN(n8852)
         );
  MUX2_X1 U10257 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n8850), .S(n10496), .Z(
        n8851) );
  OR2_X1 U10258 ( .A1(n8852), .A2(n8851), .ZN(P2_U3508) );
  INV_X1 U10259 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n8854) );
  MUX2_X1 U10260 ( .A(n8854), .B(n8853), .S(n10496), .Z(n8855) );
  OAI21_X1 U10261 ( .B1(n8856), .B2(n8860), .A(n8855), .ZN(P2_U3507) );
  MUX2_X1 U10262 ( .A(n8858), .B(n8857), .S(n10496), .Z(n8859) );
  OAI21_X1 U10263 ( .B1(n8861), .B2(n8860), .A(n8859), .ZN(P2_U3505) );
  MUX2_X1 U10264 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n8862), .S(n10496), .Z(
        P2_U3502) );
  MUX2_X1 U10265 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n8863), .S(n10496), .Z(
        P2_U3499) );
  MUX2_X1 U10266 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n8864), .S(n10496), .Z(
        P2_U3496) );
  INV_X1 U10267 ( .A(n9769), .ZN(n8868) );
  NOR4_X1 U10268 ( .A1(n4498), .A2(P2_IR_REG_30__SCAN_IN), .A3(n8865), .A4(
        P2_U3152), .ZN(n8866) );
  AOI21_X1 U10269 ( .B1(n8869), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n8866), .ZN(
        n8867) );
  OAI21_X1 U10270 ( .B1(n8868), .B2(n8872), .A(n8867), .ZN(P2_U3327) );
  INV_X1 U10271 ( .A(n9110), .ZN(n9772) );
  AOI22_X1 U10272 ( .A1(n8870), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n8869), .ZN(n8871) );
  OAI21_X1 U10273 ( .B1(n9772), .B2(n8872), .A(n8871), .ZN(P2_U3328) );
  MUX2_X1 U10274 ( .A(n8873), .B(n10413), .S(P2_STATE_REG_SCAN_IN), .Z(
        P2_U3358) );
  XNOR2_X1 U10275 ( .A(n8875), .B(n8874), .ZN(n8876) );
  XNOR2_X1 U10276 ( .A(n8877), .B(n8876), .ZN(n8885) );
  NAND2_X1 U10277 ( .A1(P1_U3084), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n8881) );
  NAND2_X1 U10278 ( .A1(n8879), .A2(n9042), .ZN(n8880) );
  OAI211_X1 U10279 ( .C1(n9481), .C2(n9026), .A(n8881), .B(n8880), .ZN(n8882)
         );
  AOI21_X1 U10280 ( .B1(n9343), .B2(n9030), .A(n8882), .ZN(n8884) );
  NAND2_X1 U10281 ( .A1(n9671), .A2(n9047), .ZN(n8883) );
  OAI211_X1 U10282 ( .C1(n8885), .C2(n9049), .A(n8884), .B(n8883), .ZN(
        P1_U3212) );
  XNOR2_X1 U10283 ( .A(n8887), .B(n8886), .ZN(n8888) );
  XNOR2_X1 U10284 ( .A(n8889), .B(n8888), .ZN(n8897) );
  INV_X1 U10285 ( .A(n8890), .ZN(n8891) );
  AOI21_X1 U10286 ( .B1(n9041), .B2(n9347), .A(n8891), .ZN(n8894) );
  NAND2_X1 U10287 ( .A1(n9042), .A2(n8892), .ZN(n8893) );
  OAI211_X1 U10288 ( .C1(n9621), .C2(n9045), .A(n8894), .B(n8893), .ZN(n8895)
         );
  AOI21_X1 U10289 ( .B1(n9739), .B2(n9031), .A(n8895), .ZN(n8896) );
  OAI21_X1 U10290 ( .B1(n8897), .B2(n9049), .A(n8896), .ZN(P1_U3213) );
  NAND2_X1 U10291 ( .A1(n8899), .A2(n8898), .ZN(n8900) );
  XOR2_X1 U10292 ( .A(n8901), .B(n8900), .Z(n8906) );
  AOI22_X1 U10293 ( .A1(n9345), .A2(n9030), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3084), .ZN(n8903) );
  NAND2_X1 U10294 ( .A1(n9041), .A2(n9540), .ZN(n8902) );
  OAI211_X1 U10295 ( .C1(n9024), .C2(n9514), .A(n8903), .B(n8902), .ZN(n8904)
         );
  AOI21_X1 U10296 ( .B1(n9690), .B2(n9031), .A(n8904), .ZN(n8905) );
  OAI21_X1 U10297 ( .B1(n8906), .B2(n9049), .A(n8905), .ZN(P1_U3214) );
  NOR2_X1 U10298 ( .A1(n4797), .A2(n8908), .ZN(n8909) );
  XNOR2_X1 U10299 ( .A(n8910), .B(n8909), .ZN(n8915) );
  NAND2_X1 U10300 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9403) );
  OAI21_X1 U10301 ( .B1(n9045), .B2(n9572), .A(n9403), .ZN(n8911) );
  AOI21_X1 U10302 ( .B1(n9041), .B2(n9607), .A(n8911), .ZN(n8912) );
  OAI21_X1 U10303 ( .B1(n9024), .B2(n9576), .A(n8912), .ZN(n8913) );
  AOI21_X1 U10304 ( .B1(n9712), .B2(n9047), .A(n8913), .ZN(n8914) );
  OAI21_X1 U10305 ( .B1(n8915), .B2(n9049), .A(n8914), .ZN(P1_U3217) );
  XOR2_X1 U10306 ( .A(n8917), .B(n8916), .Z(n8923) );
  OAI22_X1 U10307 ( .A1(n9026), .A2(n9572), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8918), .ZN(n8919) );
  AOI21_X1 U10308 ( .B1(n9030), .B2(n9540), .A(n8919), .ZN(n8920) );
  OAI21_X1 U10309 ( .B1(n9024), .B2(n9535), .A(n8920), .ZN(n8921) );
  AOI21_X1 U10310 ( .B1(n9701), .B2(n9047), .A(n8921), .ZN(n8922) );
  OAI21_X1 U10311 ( .B1(n8923), .B2(n9049), .A(n8922), .ZN(P1_U3221) );
  OAI21_X1 U10312 ( .B1(n8926), .B2(n8925), .A(n8924), .ZN(n8927) );
  NAND2_X1 U10313 ( .A1(n8927), .A2(n8977), .ZN(n8932) );
  OAI22_X1 U10314 ( .A1(n9511), .A2(n9026), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8928), .ZN(n8930) );
  NOR2_X1 U10315 ( .A1(n9481), .A2(n9045), .ZN(n8929) );
  AOI211_X1 U10316 ( .C1(n9484), .C2(n9042), .A(n8930), .B(n8929), .ZN(n8931)
         );
  OAI211_X1 U10317 ( .C1(n8933), .C2(n9019), .A(n8932), .B(n8931), .ZN(
        P1_U3223) );
  INV_X1 U10318 ( .A(n8935), .ZN(n8936) );
  AOI21_X1 U10319 ( .B1(n8934), .B2(n8937), .A(n8936), .ZN(n8944) );
  INV_X1 U10320 ( .A(n8938), .ZN(n8939) );
  AOI21_X1 U10321 ( .B1(n9030), .B2(n9593), .A(n8939), .ZN(n8941) );
  NAND2_X1 U10322 ( .A1(n9042), .A2(n9627), .ZN(n8940) );
  OAI211_X1 U10323 ( .C1(n9621), .C2(n9026), .A(n8941), .B(n8940), .ZN(n8942)
         );
  AOI21_X1 U10324 ( .B1(n9728), .B2(n9047), .A(n8942), .ZN(n8943) );
  OAI21_X1 U10325 ( .B1(n8944), .B2(n9049), .A(n8943), .ZN(P1_U3224) );
  OAI21_X1 U10326 ( .B1(n8947), .B2(n8946), .A(n8945), .ZN(n8948) );
  NAND2_X1 U10327 ( .A1(n8948), .A2(n8977), .ZN(n8955) );
  AOI21_X1 U10328 ( .B1(n9031), .B2(n8950), .A(n8949), .ZN(n8954) );
  AOI22_X1 U10329 ( .A1(n9041), .A2(n9355), .B1(n9030), .B2(n9353), .ZN(n8953)
         );
  NAND2_X1 U10330 ( .A1(n9042), .A2(n8951), .ZN(n8952) );
  NAND4_X1 U10331 ( .A1(n8955), .A2(n8954), .A3(n8953), .A4(n8952), .ZN(
        P1_U3225) );
  OAI21_X1 U10332 ( .B1(n8958), .B2(n8957), .A(n8956), .ZN(n8959) );
  NAND2_X1 U10333 ( .A1(n8959), .A2(n8977), .ZN(n8963) );
  NAND2_X1 U10334 ( .A1(n9030), .A2(n9607), .ZN(n8960) );
  NAND2_X1 U10335 ( .A1(P1_U3084), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9370) );
  OAI211_X1 U10336 ( .C1(n9635), .C2(n9026), .A(n8960), .B(n9370), .ZN(n8961)
         );
  AOI21_X1 U10337 ( .B1(n9601), .B2(n9042), .A(n8961), .ZN(n8962) );
  OAI211_X1 U10338 ( .C1(n9603), .C2(n9019), .A(n8963), .B(n8962), .ZN(
        P1_U3226) );
  INV_X1 U10339 ( .A(n8964), .ZN(n8965) );
  AOI21_X1 U10340 ( .B1(n8967), .B2(n8966), .A(n8965), .ZN(n8973) );
  NAND2_X1 U10341 ( .A1(n9501), .A2(n9030), .ZN(n8970) );
  INV_X1 U10342 ( .A(n8968), .ZN(n9529) );
  AOI22_X1 U10343 ( .A1(n9529), .A2(n9041), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3084), .ZN(n8969) );
  OAI211_X1 U10344 ( .C1(n9024), .C2(n9494), .A(n8970), .B(n8969), .ZN(n8971)
         );
  AOI21_X1 U10345 ( .B1(n8039), .B2(n9047), .A(n8971), .ZN(n8972) );
  OAI21_X1 U10346 ( .B1(n8973), .B2(n9049), .A(n8972), .ZN(P1_U3227) );
  AND2_X1 U10347 ( .A1(n8975), .A2(n8974), .ZN(n8979) );
  OAI211_X1 U10348 ( .C1(n8979), .C2(n8978), .A(n8977), .B(n8976), .ZN(n8986)
         );
  AOI21_X1 U10349 ( .B1(n9031), .B2(n8981), .A(n8980), .ZN(n8985) );
  AOI22_X1 U10350 ( .A1(n9041), .A2(n9356), .B1(n9030), .B2(n9354), .ZN(n8984)
         );
  NAND2_X1 U10351 ( .A1(n9042), .A2(n8982), .ZN(n8983) );
  NAND4_X1 U10352 ( .A1(n8986), .A2(n8985), .A3(n8984), .A4(n8983), .ZN(
        P1_U3228) );
  NAND2_X1 U10353 ( .A1(n8988), .A2(n8987), .ZN(n8989) );
  XNOR2_X1 U10354 ( .A(n8990), .B(n8989), .ZN(n8995) );
  AOI22_X1 U10355 ( .A1(n9528), .A2(n9030), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3084), .ZN(n8992) );
  NAND2_X1 U10356 ( .A1(n9041), .A2(n9592), .ZN(n8991) );
  OAI211_X1 U10357 ( .C1(n9024), .C2(n9556), .A(n8992), .B(n8991), .ZN(n8993)
         );
  AOI21_X1 U10358 ( .B1(n9707), .B2(n9047), .A(n8993), .ZN(n8994) );
  OAI21_X1 U10359 ( .B1(n8995), .B2(n9049), .A(n8994), .ZN(P1_U3231) );
  INV_X1 U10360 ( .A(n8998), .ZN(n9002) );
  AOI21_X1 U10361 ( .B1(n8998), .B2(n8997), .A(n8996), .ZN(n8999) );
  NOR2_X1 U10362 ( .A1(n8999), .A2(n9049), .ZN(n9000) );
  OAI21_X1 U10363 ( .B1(n9002), .B2(n9001), .A(n9000), .ZN(n9007) );
  OAI22_X1 U10364 ( .A1(n9026), .A2(n9563), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9003), .ZN(n9005) );
  NOR2_X1 U10365 ( .A1(n9024), .A2(n9522), .ZN(n9004) );
  AOI211_X1 U10366 ( .C1(n9030), .C2(n9529), .A(n9005), .B(n9004), .ZN(n9006)
         );
  OAI211_X1 U10367 ( .C1(n9525), .C2(n9019), .A(n9007), .B(n9006), .ZN(
        P1_U3233) );
  INV_X1 U10368 ( .A(n9010), .ZN(n9014) );
  AOI21_X1 U10369 ( .B1(n9010), .B2(n9009), .A(n9008), .ZN(n9011) );
  NOR2_X1 U10370 ( .A1(n9011), .A2(n9049), .ZN(n9012) );
  OAI21_X1 U10371 ( .B1(n9014), .B2(n9013), .A(n9012), .ZN(n9018) );
  AOI22_X1 U10372 ( .A1(n9030), .A2(n9592), .B1(P1_REG3_REG_18__SCAN_IN), .B2(
        P1_U3084), .ZN(n9015) );
  OAI21_X1 U10373 ( .B1(n9622), .B2(n9026), .A(n9015), .ZN(n9016) );
  AOI21_X1 U10374 ( .B1(n9585), .B2(n9042), .A(n9016), .ZN(n9017) );
  OAI211_X1 U10375 ( .C1(n4703), .C2(n9019), .A(n9018), .B(n9017), .ZN(
        P1_U3236) );
  NAND2_X1 U10376 ( .A1(n9022), .A2(n9021), .ZN(n9023) );
  XNOR2_X1 U10377 ( .A(n9020), .B(n9023), .ZN(n9034) );
  INV_X1 U10378 ( .A(n9415), .ZN(n9472) );
  NOR2_X1 U10379 ( .A1(n9463), .A2(n9024), .ZN(n9029) );
  OAI22_X1 U10380 ( .A1(n9027), .A2(n9026), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9025), .ZN(n9028) );
  AOI211_X1 U10381 ( .C1(n9472), .C2(n9030), .A(n9029), .B(n9028), .ZN(n9033)
         );
  NAND2_X1 U10382 ( .A1(n9674), .A2(n9031), .ZN(n9032) );
  OAI211_X1 U10383 ( .C1(n9034), .C2(n9049), .A(n9033), .B(n9032), .ZN(
        P1_U3238) );
  XNOR2_X1 U10384 ( .A(n9037), .B(n9036), .ZN(n9038) );
  XNOR2_X1 U10385 ( .A(n9035), .B(n9038), .ZN(n9050) );
  INV_X1 U10386 ( .A(n9039), .ZN(n9040) );
  AOI21_X1 U10387 ( .B1(n9041), .B2(n10255), .A(n9040), .ZN(n9044) );
  NAND2_X1 U10388 ( .A1(n9042), .A2(n9647), .ZN(n9043) );
  OAI211_X1 U10389 ( .C1(n9635), .C2(n9045), .A(n9044), .B(n9043), .ZN(n9046)
         );
  AOI21_X1 U10390 ( .B1(n9731), .B2(n9047), .A(n9046), .ZN(n9048) );
  OAI21_X1 U10391 ( .B1(n9050), .B2(n9049), .A(n9048), .ZN(P1_U3239) );
  NAND2_X1 U10392 ( .A1(n9051), .A2(n6840), .ZN(n9053) );
  OR2_X1 U10393 ( .A1(n6409), .A2(n10079), .ZN(n9052) );
  INV_X1 U10394 ( .A(n9661), .ZN(n9246) );
  INV_X1 U10395 ( .A(n9241), .ZN(n9426) );
  AOI21_X1 U10396 ( .B1(n9246), .B2(n9442), .A(n9426), .ZN(n9303) );
  INV_X1 U10397 ( .A(n9423), .ZN(n9230) );
  NAND2_X1 U10398 ( .A1(n9664), .A2(n9430), .ZN(n9427) );
  OAI211_X1 U10399 ( .C1(n9230), .C2(n9268), .A(n9427), .B(n9237), .ZN(n9054)
         );
  INV_X1 U10400 ( .A(n9442), .ZN(n9252) );
  AOI22_X1 U10401 ( .A1(n9303), .A2(n9054), .B1(n9252), .B2(n9661), .ZN(n9323)
         );
  INV_X1 U10402 ( .A(n9055), .ZN(n9273) );
  NAND2_X1 U10403 ( .A1(n9211), .A2(n9273), .ZN(n9056) );
  NAND2_X1 U10404 ( .A1(n9056), .A2(n9209), .ZN(n9057) );
  NOR2_X1 U10405 ( .A1(n9271), .A2(n9057), .ZN(n9207) );
  INV_X1 U10406 ( .A(n9192), .ZN(n9061) );
  INV_X1 U10407 ( .A(n9093), .ZN(n9058) );
  NOR2_X1 U10408 ( .A1(n9203), .A2(n9058), .ZN(n9197) );
  INV_X1 U10409 ( .A(n9197), .ZN(n9060) );
  OR2_X1 U10410 ( .A1(n9274), .A2(n9201), .ZN(n9196) );
  INV_X1 U10411 ( .A(n9196), .ZN(n9059) );
  OAI211_X1 U10412 ( .C1(n9061), .C2(n9060), .A(n9059), .B(n9211), .ZN(n9063)
         );
  INV_X1 U10413 ( .A(n9062), .ZN(n9272) );
  OR2_X1 U10414 ( .A1(n9064), .A2(n9270), .ZN(n9220) );
  AOI211_X1 U10415 ( .C1(n9207), .C2(n9063), .A(n9272), .B(n9220), .ZN(n9068)
         );
  INV_X1 U10416 ( .A(n9064), .ZN(n9066) );
  OR2_X1 U10417 ( .A1(n9065), .A2(n4521), .ZN(n9217) );
  NAND2_X1 U10418 ( .A1(n9066), .A2(n9217), .ZN(n9067) );
  NAND2_X1 U10419 ( .A1(n9067), .A2(n9231), .ZN(n9222) );
  NOR2_X1 U10420 ( .A1(n9068), .A2(n9222), .ZN(n9070) );
  NOR2_X1 U10421 ( .A1(n9070), .A2(n9069), .ZN(n9319) );
  INV_X1 U10422 ( .A(n9071), .ZN(n9091) );
  INV_X1 U10423 ( .A(n9072), .ZN(n9310) );
  NAND2_X1 U10424 ( .A1(n9073), .A2(n9074), .ZN(n9075) );
  AOI211_X1 U10425 ( .C1(n9076), .C2(n9357), .A(n9327), .B(n9075), .ZN(n9077)
         );
  NOR3_X1 U10426 ( .A1(n9306), .A2(n9310), .A3(n9077), .ZN(n9081) );
  AND2_X1 U10427 ( .A1(n9307), .A2(n9078), .ZN(n9305) );
  INV_X1 U10428 ( .A(n9305), .ZN(n9080) );
  OAI211_X1 U10429 ( .C1(n9081), .C2(n9080), .A(n9312), .B(n9079), .ZN(n9090)
         );
  INV_X1 U10430 ( .A(n9082), .ZN(n9185) );
  NAND2_X1 U10431 ( .A1(n9093), .A2(n9185), .ZN(n9191) );
  NAND3_X1 U10432 ( .A1(n9186), .A2(n9181), .A3(n9158), .ZN(n9083) );
  NOR2_X1 U10433 ( .A1(n9191), .A2(n9083), .ZN(n9101) );
  INV_X1 U10434 ( .A(n9101), .ZN(n9089) );
  NAND2_X1 U10435 ( .A1(n10248), .A2(n9094), .ZN(n9162) );
  INV_X1 U10436 ( .A(n9162), .ZN(n9086) );
  NAND2_X1 U10437 ( .A1(n9148), .A2(n9137), .ZN(n9084) );
  NOR2_X1 U10438 ( .A1(n9150), .A2(n9084), .ZN(n9085) );
  NAND3_X1 U10439 ( .A1(n9087), .A2(n9086), .A3(n9085), .ZN(n9088) );
  OR2_X1 U10440 ( .A1(n9089), .A2(n9088), .ZN(n9304) );
  AOI21_X1 U10441 ( .B1(n9091), .B2(n9090), .A(n9304), .ZN(n9108) );
  NAND4_X1 U10442 ( .A1(n9093), .A2(n9185), .A3(n9186), .A4(n9092), .ZN(n9104)
         );
  INV_X1 U10443 ( .A(n9094), .ZN(n9096) );
  AOI21_X1 U10444 ( .B1(n4847), .B2(n9147), .A(n4840), .ZN(n9095) );
  OAI21_X1 U10445 ( .B1(n9096), .B2(n9095), .A(n9166), .ZN(n9097) );
  NAND2_X1 U10446 ( .A1(n9097), .A2(n10248), .ZN(n9100) );
  AOI21_X1 U10447 ( .B1(n9100), .B2(n9099), .A(n9098), .ZN(n9102) );
  OAI21_X1 U10448 ( .B1(n9168), .B2(n9102), .A(n9101), .ZN(n9103) );
  OAI211_X1 U10449 ( .C1(n9304), .C2(n9134), .A(n9104), .B(n9103), .ZN(n9316)
         );
  INV_X1 U10450 ( .A(n9222), .ZN(n9106) );
  INV_X1 U10451 ( .A(n9203), .ZN(n9105) );
  NAND3_X1 U10452 ( .A1(n9106), .A2(n9207), .A3(n9105), .ZN(n9320) );
  INV_X1 U10453 ( .A(n9320), .ZN(n9107) );
  OAI21_X1 U10454 ( .B1(n9108), .B2(n9316), .A(n9107), .ZN(n9109) );
  NAND4_X1 U10455 ( .A1(n9303), .A2(n9419), .A3(n9319), .A4(n9109), .ZN(n9116)
         );
  NAND2_X1 U10456 ( .A1(n9110), .A2(n6840), .ZN(n9112) );
  INV_X1 U10457 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n9890) );
  OR2_X1 U10458 ( .A1(n6409), .A2(n9890), .ZN(n9111) );
  NAND2_X1 U10459 ( .A1(n4481), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n9115) );
  NAND2_X1 U10460 ( .A1(n9118), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n9114) );
  NAND2_X1 U10461 ( .A1(n4480), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n9113) );
  AND3_X1 U10462 ( .A1(n9115), .A2(n9114), .A3(n9113), .ZN(n9431) );
  AOI21_X1 U10463 ( .B1(n9323), .B2(n9116), .A(n4506), .ZN(n9123) );
  NAND2_X1 U10464 ( .A1(n4481), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n9121) );
  NAND2_X1 U10465 ( .A1(n9118), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n9120) );
  NAND2_X1 U10466 ( .A1(n4480), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n9119) );
  AND3_X1 U10467 ( .A1(n9121), .A2(n9120), .A3(n9119), .ZN(n9407) );
  AOI21_X1 U10468 ( .B1(n9431), .B2(n10267), .A(n9326), .ZN(n9300) );
  INV_X1 U10469 ( .A(n9300), .ZN(n9122) );
  OAI21_X1 U10470 ( .B1(n9123), .B2(n9122), .A(n9267), .ZN(n9124) );
  XNOR2_X1 U10471 ( .A(n9124), .B(n9544), .ZN(n9334) );
  INV_X1 U10472 ( .A(n9125), .ZN(n9126) );
  AOI211_X1 U10473 ( .C1(n9127), .C2(n9307), .A(n9126), .B(n9309), .ZN(n9131)
         );
  INV_X1 U10474 ( .A(n9282), .ZN(n9128) );
  NAND2_X1 U10475 ( .A1(n9128), .A2(n9308), .ZN(n9130) );
  OAI21_X1 U10476 ( .B1(n9131), .B2(n9130), .A(n9129), .ZN(n9133) );
  INV_X1 U10477 ( .A(n9137), .ZN(n9132) );
  AOI21_X1 U10478 ( .B1(n9133), .B2(n9134), .A(n9132), .ZN(n9135) );
  INV_X1 U10479 ( .A(n9136), .ZN(n9138) );
  NAND3_X1 U10480 ( .A1(n9138), .A2(n9256), .A3(n9137), .ZN(n9139) );
  AOI211_X1 U10481 ( .C1(n9149), .C2(n10345), .A(n9141), .B(n9140), .ZN(n9143)
         );
  INV_X1 U10482 ( .A(n9284), .ZN(n9142) );
  NOR3_X1 U10483 ( .A1(n9143), .A2(n9142), .A3(n9256), .ZN(n9145) );
  NAND2_X1 U10484 ( .A1(n10248), .A2(n9146), .ZN(n9153) );
  AOI21_X1 U10485 ( .B1(n9149), .B2(n9148), .A(n9147), .ZN(n9151) );
  NOR2_X1 U10486 ( .A1(n9151), .A2(n9150), .ZN(n9152) );
  INV_X1 U10487 ( .A(n9161), .ZN(n9155) );
  INV_X1 U10488 ( .A(n9158), .ZN(n9169) );
  NAND2_X1 U10489 ( .A1(n10248), .A2(n9251), .ZN(n9165) );
  NAND2_X1 U10490 ( .A1(n9160), .A2(n9159), .ZN(n9164) );
  NAND3_X1 U10491 ( .A1(n9162), .A2(n9256), .A3(n9161), .ZN(n9163) );
  OAI211_X1 U10492 ( .C1(n9166), .C2(n9165), .A(n9164), .B(n9163), .ZN(n9167)
         );
  NOR4_X1 U10493 ( .A1(n9170), .A2(n9169), .A3(n9168), .A4(n9167), .ZN(n9184)
         );
  INV_X1 U10494 ( .A(n9174), .ZN(n10269) );
  NAND2_X1 U10495 ( .A1(n9347), .A2(n9256), .ZN(n9173) );
  INV_X1 U10496 ( .A(n9173), .ZN(n9171) );
  AOI22_X1 U10497 ( .A1(n10269), .A2(n9171), .B1(n9256), .B2(n10255), .ZN(
        n9180) );
  NAND2_X1 U10498 ( .A1(n9172), .A2(n9251), .ZN(n9175) );
  OAI22_X1 U10499 ( .A1(n10269), .A2(n9175), .B1(n9256), .B2(n10255), .ZN(
        n9178) );
  OAI21_X1 U10500 ( .B1(n9636), .B2(n9173), .A(n10269), .ZN(n9177) );
  OAI21_X1 U10501 ( .B1(n10255), .B2(n9175), .A(n9174), .ZN(n9176) );
  AOI22_X1 U10502 ( .A1(n9178), .A2(n9739), .B1(n9177), .B2(n9176), .ZN(n9179)
         );
  OAI211_X1 U10503 ( .C1(n9180), .C2(n9739), .A(n9637), .B(n9179), .ZN(n9183)
         );
  MUX2_X1 U10504 ( .A(n9614), .B(n9181), .S(n9256), .Z(n9182) );
  OAI211_X1 U10505 ( .C1(n9184), .C2(n9183), .A(n9618), .B(n9182), .ZN(n9195)
         );
  NAND2_X1 U10506 ( .A1(n9185), .A2(n9587), .ZN(n9605) );
  INV_X1 U10507 ( .A(n9186), .ZN(n9189) );
  INV_X1 U10508 ( .A(n9187), .ZN(n9188) );
  MUX2_X1 U10509 ( .A(n9189), .B(n9188), .S(n9256), .Z(n9190) );
  NOR2_X1 U10510 ( .A1(n9605), .A2(n9190), .ZN(n9194) );
  MUX2_X1 U10511 ( .A(n9192), .B(n9191), .S(n9256), .Z(n9193) );
  AOI21_X1 U10512 ( .B1(n9195), .B2(n9194), .A(n9193), .ZN(n9202) );
  INV_X1 U10513 ( .A(n9202), .ZN(n9198) );
  AOI21_X1 U10514 ( .B1(n9198), .B2(n9197), .A(n9196), .ZN(n9206) );
  INV_X1 U10515 ( .A(n9199), .ZN(n9200) );
  NOR3_X1 U10516 ( .A1(n9204), .A2(n9203), .A3(n9273), .ZN(n9205) );
  NAND2_X1 U10517 ( .A1(n9210), .A2(n9211), .ZN(n9208) );
  AOI21_X1 U10518 ( .B1(n9208), .B2(n9207), .A(n9272), .ZN(n9216) );
  OAI21_X1 U10519 ( .B1(n9210), .B2(n9274), .A(n9209), .ZN(n9214) );
  INV_X1 U10520 ( .A(n9211), .ZN(n9212) );
  NOR2_X1 U10521 ( .A1(n9272), .A2(n9212), .ZN(n9213) );
  AOI21_X1 U10522 ( .B1(n9214), .B2(n9213), .A(n9271), .ZN(n9215) );
  NOR3_X1 U10523 ( .A1(n9218), .A2(n9220), .A3(n9217), .ZN(n9225) );
  NAND2_X1 U10524 ( .A1(n9220), .A2(n9219), .ZN(n9221) );
  NAND2_X1 U10525 ( .A1(n9221), .A2(n9467), .ZN(n9223) );
  MUX2_X1 U10526 ( .A(n9223), .B(n9222), .S(n9256), .Z(n9224) );
  OR2_X1 U10527 ( .A1(n9225), .A2(n9224), .ZN(n9229) );
  OAI22_X1 U10528 ( .A1(n9229), .A2(n9674), .B1(n9256), .B2(n9231), .ZN(n9228)
         );
  OAI21_X1 U10529 ( .B1(n9674), .B2(n9467), .A(n9481), .ZN(n9226) );
  MUX2_X1 U10530 ( .A(n9674), .B(n9226), .S(n9256), .Z(n9227) );
  INV_X1 U10531 ( .A(n9229), .ZN(n9236) );
  AOI21_X1 U10532 ( .B1(n9231), .B2(n9344), .A(n9230), .ZN(n9234) );
  INV_X1 U10533 ( .A(n9237), .ZN(n9232) );
  AOI21_X1 U10534 ( .B1(n9467), .B2(n9674), .A(n9232), .ZN(n9233) );
  MUX2_X1 U10535 ( .A(n9234), .B(n9233), .S(n9256), .Z(n9235) );
  AOI21_X1 U10536 ( .B1(n9236), .B2(n9419), .A(n9235), .ZN(n9239) );
  MUX2_X1 U10537 ( .A(n9237), .B(n9423), .S(n9256), .Z(n9238) );
  OAI211_X1 U10538 ( .C1(n9240), .C2(n9239), .A(n9448), .B(n9238), .ZN(n9243)
         );
  MUX2_X1 U10539 ( .A(n9241), .B(n9427), .S(n9256), .Z(n9242) );
  NAND2_X1 U10540 ( .A1(n9243), .A2(n9242), .ZN(n9262) );
  INV_X1 U10541 ( .A(n9407), .ZN(n9342) );
  NAND2_X1 U10542 ( .A1(n4921), .A2(n9342), .ZN(n9245) );
  NAND2_X1 U10543 ( .A1(n10267), .A2(n9245), .ZN(n9322) );
  NAND2_X1 U10544 ( .A1(n9252), .A2(n9251), .ZN(n9253) );
  NAND3_X1 U10545 ( .A1(n9322), .A2(n9256), .A3(n9246), .ZN(n9247) );
  AOI21_X1 U10546 ( .B1(n9253), .B2(n9247), .A(n9302), .ZN(n9248) );
  AOI21_X1 U10547 ( .B1(n9249), .B2(n9322), .A(n9248), .ZN(n9261) );
  INV_X1 U10548 ( .A(n9250), .ZN(n9258) );
  NOR3_X1 U10549 ( .A1(n9661), .A2(n9252), .A3(n9251), .ZN(n9255) );
  INV_X1 U10550 ( .A(n9253), .ZN(n9254) );
  AOI22_X1 U10551 ( .A1(n9322), .A2(n9255), .B1(n9254), .B2(n9661), .ZN(n9257)
         );
  OAI22_X1 U10552 ( .A1(n9258), .A2(n9257), .B1(n9256), .B2(n9322), .ZN(n9259)
         );
  AOI22_X1 U10553 ( .A1(n9259), .A2(n9267), .B1(n9256), .B2(n9302), .ZN(n9260)
         );
  NAND2_X1 U10554 ( .A1(n9263), .A2(n5055), .ZN(n9265) );
  INV_X1 U10555 ( .A(n9267), .ZN(n9299) );
  XNOR2_X1 U10556 ( .A(n9661), .B(n9442), .ZN(n9422) );
  INV_X1 U10557 ( .A(n9422), .ZN(n9428) );
  INV_X1 U10558 ( .A(n9500), .ZN(n9296) );
  OR2_X1 U10559 ( .A1(n9270), .A2(n4521), .ZN(n9508) );
  NOR2_X1 U10560 ( .A1(n9272), .A2(n9271), .ZN(n9526) );
  NOR2_X1 U10561 ( .A1(n9274), .A2(n9273), .ZN(n9560) );
  INV_X1 U10562 ( .A(n9567), .ZN(n9569) );
  NOR4_X1 U10563 ( .A1(n9277), .A2(n9276), .A3(n9275), .A4(n6319), .ZN(n9279)
         );
  NAND3_X1 U10564 ( .A1(n9279), .A2(n4501), .A3(n9278), .ZN(n9283) );
  NOR4_X1 U10565 ( .A1(n9283), .A2(n9282), .A3(n9281), .A4(n9280), .ZN(n9288)
         );
  AND2_X1 U10566 ( .A1(n9285), .A2(n9284), .ZN(n10348) );
  NAND4_X1 U10567 ( .A1(n9288), .A2(n9287), .A3(n9286), .A4(n10348), .ZN(n9290) );
  NOR4_X1 U10568 ( .A1(n9291), .A2(n9290), .A3(n10247), .A4(n9289), .ZN(n9292)
         );
  NAND3_X1 U10569 ( .A1(n9618), .A2(n9637), .A3(n9292), .ZN(n9293) );
  NOR4_X1 U10570 ( .A1(n9569), .A2(n9605), .A3(n9591), .A4(n9293), .ZN(n9294)
         );
  NAND4_X1 U10571 ( .A1(n9526), .A2(n9538), .A3(n9560), .A4(n9294), .ZN(n9295)
         );
  NOR4_X1 U10572 ( .A1(n9296), .A2(n9478), .A3(n9508), .A4(n9295), .ZN(n9297)
         );
  NAND4_X1 U10573 ( .A1(n9448), .A2(n9419), .A3(n9470), .A4(n9297), .ZN(n9298)
         );
  NOR4_X1 U10574 ( .A1(n9299), .A2(n4506), .A3(n9428), .A4(n9298), .ZN(n9301)
         );
  AOI21_X1 U10575 ( .B1(n9301), .B2(n9300), .A(n5055), .ZN(n9332) );
  INV_X1 U10576 ( .A(n9302), .ZN(n9329) );
  INV_X1 U10577 ( .A(n9303), .ZN(n9325) );
  INV_X1 U10578 ( .A(n9304), .ZN(n9318) );
  NAND3_X1 U10579 ( .A1(n9306), .A2(n9305), .A3(n9308), .ZN(n9313) );
  OAI211_X1 U10580 ( .C1(n9310), .C2(n9309), .A(n9308), .B(n9307), .ZN(n9311)
         );
  NAND3_X1 U10581 ( .A1(n9313), .A2(n9312), .A3(n9311), .ZN(n9315) );
  NAND2_X1 U10582 ( .A1(n9315), .A2(n9314), .ZN(n9317) );
  AOI21_X1 U10583 ( .B1(n9318), .B2(n9317), .A(n9316), .ZN(n9321) );
  OAI211_X1 U10584 ( .C1(n9321), .C2(n9320), .A(n9319), .B(n9423), .ZN(n9324)
         );
  OAI211_X1 U10585 ( .C1(n9325), .C2(n9324), .A(n9323), .B(n9322), .ZN(n9328)
         );
  AOI211_X1 U10586 ( .C1(n9329), .C2(n9328), .A(n9327), .B(n9326), .ZN(n9330)
         );
  NOR2_X1 U10587 ( .A1(n9332), .A2(n9330), .ZN(n9331) );
  MUX2_X1 U10588 ( .A(n9332), .B(n9331), .S(n9544), .Z(n9333) );
  NAND4_X1 U10589 ( .A1(n9336), .A2(n9762), .A3(n9405), .A4(n9335), .ZN(n9337)
         );
  OAI211_X1 U10590 ( .C1(n9338), .C2(n9340), .A(n9337), .B(P1_B_REG_SCAN_IN), 
        .ZN(n9339) );
  OAI21_X1 U10591 ( .B1(n9341), .B2(n9340), .A(n9339), .ZN(P1_U3240) );
  MUX2_X1 U10592 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n9342), .S(P1_U4006), .Z(
        P1_U3586) );
  MUX2_X1 U10593 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n4921), .S(P1_U4006), .Z(
        P1_U3585) );
  MUX2_X1 U10594 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9442), .S(P1_U4006), .Z(
        P1_U3584) );
  MUX2_X1 U10595 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9343), .S(P1_U4006), .Z(
        P1_U3583) );
  MUX2_X1 U10596 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9472), .S(P1_U4006), .Z(
        P1_U3582) );
  MUX2_X1 U10597 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9344), .S(P1_U4006), .Z(
        P1_U3581) );
  MUX2_X1 U10598 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9501), .S(P1_U4006), .Z(
        P1_U3580) );
  MUX2_X1 U10599 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9345), .S(P1_U4006), .Z(
        P1_U3579) );
  MUX2_X1 U10600 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9529), .S(P1_U4006), .Z(
        P1_U3578) );
  MUX2_X1 U10601 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9540), .S(P1_U4006), .Z(
        P1_U3577) );
  MUX2_X1 U10602 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9528), .S(P1_U4006), .Z(
        P1_U3576) );
  MUX2_X1 U10603 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9539), .S(P1_U4006), .Z(
        P1_U3575) );
  MUX2_X1 U10604 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9592), .S(P1_U4006), .Z(
        P1_U3574) );
  MUX2_X1 U10605 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9607), .S(P1_U4006), .Z(
        P1_U3573) );
  MUX2_X1 U10606 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9593), .S(P1_U4006), .Z(
        P1_U3572) );
  MUX2_X1 U10607 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9606), .S(P1_U4006), .Z(
        P1_U3571) );
  MUX2_X1 U10608 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9346), .S(P1_U4006), .Z(
        P1_U3570) );
  MUX2_X1 U10609 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n10255), .S(P1_U4006), .Z(
        P1_U3569) );
  MUX2_X1 U10610 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9347), .S(P1_U4006), .Z(
        P1_U3568) );
  MUX2_X1 U10611 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n10253), .S(P1_U4006), .Z(
        P1_U3567) );
  MUX2_X1 U10612 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9348), .S(P1_U4006), .Z(
        P1_U3566) );
  MUX2_X1 U10613 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9349), .S(P1_U4006), .Z(
        P1_U3565) );
  MUX2_X1 U10614 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9350), .S(P1_U4006), .Z(
        P1_U3564) );
  MUX2_X1 U10615 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9351), .S(P1_U4006), .Z(
        P1_U3563) );
  MUX2_X1 U10616 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9352), .S(P1_U4006), .Z(
        P1_U3562) );
  MUX2_X1 U10617 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9353), .S(P1_U4006), .Z(
        P1_U3561) );
  MUX2_X1 U10618 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9354), .S(P1_U4006), .Z(
        P1_U3560) );
  MUX2_X1 U10619 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9355), .S(P1_U4006), .Z(
        P1_U3559) );
  MUX2_X1 U10620 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9356), .S(P1_U4006), .Z(
        P1_U3558) );
  MUX2_X1 U10621 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n9357), .S(P1_U4006), .Z(
        P1_U3557) );
  MUX2_X1 U10622 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n9358), .S(P1_U4006), .Z(
        P1_U3556) );
  MUX2_X1 U10623 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n9359), .S(P1_U4006), .Z(
        P1_U3555) );
  INV_X1 U10624 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9375) );
  NAND2_X1 U10625 ( .A1(P1_REG2_REG_17__SCAN_IN), .A2(n9383), .ZN(n9361) );
  OAI21_X1 U10626 ( .B1(n9383), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9361), .ZN(
        n9362) );
  AOI211_X1 U10627 ( .C1(n9363), .C2(n9362), .A(n9382), .B(n9385), .ZN(n9364)
         );
  AOI21_X1 U10628 ( .B1(n10324), .B2(n9383), .A(n9364), .ZN(n9374) );
  AOI21_X1 U10629 ( .B1(n9366), .B2(P1_REG1_REG_16__SCAN_IN), .A(n9365), .ZN(
        n9369) );
  XNOR2_X1 U10630 ( .A(n9383), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n9368) );
  NOR2_X1 U10631 ( .A1(n9369), .A2(n9368), .ZN(n9376) );
  AOI211_X1 U10632 ( .C1(n9369), .C2(n9368), .A(n9376), .B(n9367), .ZN(n9372)
         );
  INV_X1 U10633 ( .A(n9370), .ZN(n9371) );
  NOR2_X1 U10634 ( .A1(n9372), .A2(n9371), .ZN(n9373) );
  OAI211_X1 U10635 ( .C1(n10337), .C2(n9375), .A(n9374), .B(n9373), .ZN(
        P1_U3258) );
  XOR2_X1 U10636 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9395), .Z(n9378) );
  AOI21_X1 U10637 ( .B1(n9383), .B2(P1_REG1_REG_17__SCAN_IN), .A(n9376), .ZN(
        n9377) );
  NAND2_X1 U10638 ( .A1(n9378), .A2(n9377), .ZN(n9394) );
  OAI21_X1 U10639 ( .B1(n9378), .B2(n9377), .A(n9394), .ZN(n9390) );
  INV_X1 U10640 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n9381) );
  NAND2_X1 U10641 ( .A1(n10324), .A2(n9395), .ZN(n9380) );
  NAND2_X1 U10642 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_U3084), .ZN(n9379) );
  OAI211_X1 U10643 ( .C1(n10337), .C2(n9381), .A(n9380), .B(n9379), .ZN(n9389)
         );
  AOI21_X1 U10644 ( .B1(n9383), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9382), .ZN(
        n9387) );
  NAND2_X1 U10645 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n9395), .ZN(n9384) );
  OAI21_X1 U10646 ( .B1(n9395), .B2(P1_REG2_REG_18__SCAN_IN), .A(n9384), .ZN(
        n9386) );
  NOR2_X1 U10647 ( .A1(n9387), .A2(n9386), .ZN(n9392) );
  AOI211_X1 U10648 ( .C1(n9387), .C2(n9386), .A(n9392), .B(n9385), .ZN(n9388)
         );
  AOI211_X1 U10649 ( .C1(n10332), .C2(n9390), .A(n9389), .B(n9388), .ZN(n9391)
         );
  INV_X1 U10650 ( .A(n9391), .ZN(P1_U3259) );
  INV_X1 U10651 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n9404) );
  AOI21_X1 U10652 ( .B1(n9395), .B2(P1_REG2_REG_18__SCAN_IN), .A(n9392), .ZN(
        n9393) );
  XNOR2_X1 U10653 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n9393), .ZN(n9400) );
  OAI21_X1 U10654 ( .B1(P1_REG1_REG_18__SCAN_IN), .B2(n9395), .A(n9394), .ZN(
        n9397) );
  INV_X1 U10655 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9396) );
  XOR2_X1 U10656 ( .A(n9397), .B(n9396), .Z(n9398) );
  AOI22_X1 U10657 ( .A1(n9400), .A2(n10331), .B1(n10332), .B2(n9398), .ZN(
        n9402) );
  INV_X1 U10658 ( .A(n9398), .ZN(n9401) );
  NAND2_X1 U10659 ( .A1(n9405), .A2(P1_B_REG_SCAN_IN), .ZN(n9406) );
  NAND2_X1 U10660 ( .A1(n10254), .A2(n9406), .ZN(n9432) );
  NOR2_X1 U10661 ( .A1(n9407), .A2(n9432), .ZN(n10266) );
  INV_X1 U10662 ( .A(n10266), .ZN(n9408) );
  NOR2_X1 U10663 ( .A1(n9408), .A2(n10362), .ZN(n9412) );
  NOR2_X1 U10664 ( .A1(n9409), .A2(n10364), .ZN(n9410) );
  AOI211_X1 U10665 ( .C1(n10362), .C2(P1_REG2_REG_31__SCAN_IN), .A(n9412), .B(
        n9410), .ZN(n9411) );
  OAI21_X1 U10666 ( .B1(n9657), .B2(n9651), .A(n9411), .ZN(P1_U3261) );
  AOI21_X1 U10667 ( .B1(n10362), .B2(P1_REG2_REG_30__SCAN_IN), .A(n9412), .ZN(
        n9414) );
  NAND2_X1 U10668 ( .A1(n10267), .A2(n9648), .ZN(n9413) );
  OAI211_X1 U10669 ( .C1(n10264), .C2(n9651), .A(n9414), .B(n9413), .ZN(
        P1_U3262) );
  INV_X1 U10670 ( .A(n9664), .ZN(n9457) );
  INV_X1 U10671 ( .A(n9448), .ZN(n9417) );
  NAND2_X1 U10672 ( .A1(n9416), .A2(n9415), .ZN(n9446) );
  NAND2_X1 U10673 ( .A1(n9417), .A2(n9446), .ZN(n9421) );
  INV_X1 U10674 ( .A(n9658), .ZN(n9440) );
  AOI21_X1 U10675 ( .B1(n9441), .B2(n9427), .A(n9426), .ZN(n9429) );
  OAI21_X1 U10676 ( .B1(n9433), .B2(n9555), .A(n4524), .ZN(n9438) );
  NAND2_X1 U10677 ( .A1(n9661), .A2(n9452), .ZN(n9434) );
  NAND2_X1 U10678 ( .A1(n9435), .A2(n9434), .ZN(n9659) );
  AOI22_X1 U10679 ( .A1(n9661), .A2(n9648), .B1(P1_REG2_REG_29__SCAN_IN), .B2(
        n10362), .ZN(n9436) );
  OAI21_X1 U10680 ( .B1(n9659), .B2(n9651), .A(n9436), .ZN(n9437) );
  AOI21_X1 U10681 ( .B1(n9438), .B2(n10366), .A(n9437), .ZN(n9439) );
  OAI21_X1 U10682 ( .B1(n9440), .B2(n9633), .A(n9439), .ZN(P1_U3355) );
  XOR2_X1 U10683 ( .A(n9448), .B(n9441), .Z(n9443) );
  AOI222_X1 U10684 ( .A1(n10355), .A2(n9443), .B1(n9442), .B2(n10254), .C1(
        n9472), .C2(n10252), .ZN(n9667) );
  NAND2_X1 U10685 ( .A1(n9445), .A2(n9444), .ZN(n9447) );
  NAND2_X1 U10686 ( .A1(n9447), .A2(n9446), .ZN(n9449) );
  NAND2_X1 U10687 ( .A1(n9449), .A2(n9448), .ZN(n9450) );
  INV_X1 U10688 ( .A(n9633), .ZN(n9547) );
  NAND2_X1 U10689 ( .A1(n9663), .A2(n9547), .ZN(n9460) );
  INV_X1 U10690 ( .A(n9452), .ZN(n9453) );
  AOI21_X1 U10691 ( .B1(n9664), .B2(n9454), .A(n9453), .ZN(n9665) );
  AOI22_X1 U10692 ( .A1(n9455), .A2(n10360), .B1(P1_REG2_REG_28__SCAN_IN), 
        .B2(n10362), .ZN(n9456) );
  OAI21_X1 U10693 ( .B1(n9457), .B2(n10364), .A(n9456), .ZN(n9458) );
  AOI21_X1 U10694 ( .B1(n9665), .B2(n10343), .A(n9458), .ZN(n9459) );
  OAI211_X1 U10695 ( .C1(n10362), .C2(n9667), .A(n9460), .B(n9459), .ZN(
        P1_U3263) );
  XNOR2_X1 U10696 ( .A(n9461), .B(n9470), .ZN(n9678) );
  AOI21_X1 U10697 ( .B1(n9674), .B2(n9482), .A(n9462), .ZN(n9675) );
  INV_X1 U10698 ( .A(n9674), .ZN(n9466) );
  INV_X1 U10699 ( .A(n9463), .ZN(n9464) );
  AOI22_X1 U10700 ( .A1(n9464), .A2(n10360), .B1(P1_REG2_REG_26__SCAN_IN), 
        .B2(n10362), .ZN(n9465) );
  OAI21_X1 U10701 ( .B1(n9466), .B2(n10364), .A(n9465), .ZN(n9475) );
  INV_X1 U10702 ( .A(n9467), .ZN(n9468) );
  NOR2_X1 U10703 ( .A1(n9469), .A2(n9468), .ZN(n9471) );
  XNOR2_X1 U10704 ( .A(n9471), .B(n9470), .ZN(n9473) );
  AOI222_X1 U10705 ( .A1(n10355), .A2(n9473), .B1(n9472), .B2(n10254), .C1(
        n9501), .C2(n10252), .ZN(n9677) );
  NOR2_X1 U10706 ( .A1(n9677), .A2(n10362), .ZN(n9474) );
  AOI211_X1 U10707 ( .C1(n9675), .C2(n10343), .A(n9475), .B(n9474), .ZN(n9476)
         );
  OAI21_X1 U10708 ( .B1(n9678), .B2(n9633), .A(n9476), .ZN(P1_U3265) );
  XOR2_X1 U10709 ( .A(n9478), .B(n9477), .Z(n9683) );
  AOI22_X1 U10710 ( .A1(n9681), .A2(n9648), .B1(P1_REG2_REG_25__SCAN_IN), .B2(
        n10362), .ZN(n9489) );
  XNOR2_X1 U10711 ( .A(n9479), .B(n9478), .ZN(n9480) );
  OAI222_X1 U10712 ( .A1(n10352), .A2(n9511), .B1(n10350), .B2(n9481), .C1(
        n9480), .C2(n9620), .ZN(n9679) );
  INV_X1 U10713 ( .A(n9482), .ZN(n9483) );
  AOI211_X1 U10714 ( .C1(n9681), .C2(n9491), .A(n10388), .B(n9483), .ZN(n9680)
         );
  INV_X1 U10715 ( .A(n9680), .ZN(n9486) );
  INV_X1 U10716 ( .A(n9484), .ZN(n9485) );
  OAI22_X1 U10717 ( .A1(n9486), .A2(n4485), .B1(n9555), .B2(n9485), .ZN(n9487)
         );
  OAI21_X1 U10718 ( .B1(n9679), .B2(n9487), .A(n10366), .ZN(n9488) );
  OAI211_X1 U10719 ( .C1(n9683), .C2(n9633), .A(n9489), .B(n9488), .ZN(
        P1_U3266) );
  XNOR2_X1 U10720 ( .A(n9490), .B(n9500), .ZN(n9687) );
  INV_X1 U10721 ( .A(n9512), .ZN(n9493) );
  INV_X1 U10722 ( .A(n9491), .ZN(n9492) );
  AOI211_X1 U10723 ( .C1(n8039), .C2(n9493), .A(n10388), .B(n9492), .ZN(n9684)
         );
  INV_X1 U10724 ( .A(n9494), .ZN(n9495) );
  AOI22_X1 U10725 ( .A1(n9495), .A2(n10360), .B1(P1_REG2_REG_24__SCAN_IN), 
        .B2(n10362), .ZN(n9496) );
  OAI21_X1 U10726 ( .B1(n9497), .B2(n10364), .A(n9496), .ZN(n9504) );
  OAI21_X1 U10727 ( .B1(n9500), .B2(n9499), .A(n9498), .ZN(n9502) );
  AOI222_X1 U10728 ( .A1(n10355), .A2(n9502), .B1(n9501), .B2(n10254), .C1(
        n9529), .C2(n10252), .ZN(n9686) );
  NOR2_X1 U10729 ( .A1(n9686), .A2(n10362), .ZN(n9503) );
  AOI211_X1 U10730 ( .C1(n9684), .C2(n9626), .A(n9504), .B(n9503), .ZN(n9505)
         );
  OAI21_X1 U10731 ( .B1(n9687), .B2(n9633), .A(n9505), .ZN(P1_U3267) );
  XNOR2_X1 U10732 ( .A(n9506), .B(n9508), .ZN(n9692) );
  AOI22_X1 U10733 ( .A1(n9690), .A2(n9648), .B1(P1_REG2_REG_23__SCAN_IN), .B2(
        n10362), .ZN(n9519) );
  XOR2_X1 U10734 ( .A(n9508), .B(n9507), .Z(n9509) );
  OAI222_X1 U10735 ( .A1(n10350), .A2(n9511), .B1(n10352), .B2(n9510), .C1(
        n9620), .C2(n9509), .ZN(n9688) );
  INV_X1 U10736 ( .A(n9521), .ZN(n9513) );
  AOI211_X1 U10737 ( .C1(n9690), .C2(n9513), .A(n10388), .B(n9512), .ZN(n9689)
         );
  INV_X1 U10738 ( .A(n9689), .ZN(n9516) );
  OAI22_X1 U10739 ( .A1(n9516), .A2(n4485), .B1(n9555), .B2(n9514), .ZN(n9517)
         );
  OAI21_X1 U10740 ( .B1(n9688), .B2(n9517), .A(n10366), .ZN(n9518) );
  OAI211_X1 U10741 ( .C1(n9692), .C2(n9633), .A(n9519), .B(n9518), .ZN(
        P1_U3268) );
  XOR2_X1 U10742 ( .A(n9520), .B(n9526), .Z(n9697) );
  AOI21_X1 U10743 ( .B1(n9693), .B2(n9534), .A(n9521), .ZN(n9694) );
  INV_X1 U10744 ( .A(n9522), .ZN(n9523) );
  AOI22_X1 U10745 ( .A1(n9523), .A2(n10360), .B1(n10362), .B2(
        P1_REG2_REG_22__SCAN_IN), .ZN(n9524) );
  OAI21_X1 U10746 ( .B1(n9525), .B2(n10364), .A(n9524), .ZN(n9532) );
  XNOR2_X1 U10747 ( .A(n9527), .B(n9526), .ZN(n9530) );
  AOI222_X1 U10748 ( .A1(n10355), .A2(n9530), .B1(n9529), .B2(n10254), .C1(
        n9528), .C2(n10252), .ZN(n9696) );
  NOR2_X1 U10749 ( .A1(n9696), .A2(n10362), .ZN(n9531) );
  AOI211_X1 U10750 ( .C1(n9694), .C2(n10343), .A(n9532), .B(n9531), .ZN(n9533)
         );
  OAI21_X1 U10751 ( .B1(n9697), .B2(n9633), .A(n9533), .ZN(P1_U3269) );
  AOI211_X1 U10752 ( .C1(n9701), .C2(n9552), .A(n10388), .B(n4698), .ZN(n9700)
         );
  NOR2_X1 U10753 ( .A1(n9535), .A2(n9555), .ZN(n9543) );
  OAI21_X1 U10754 ( .B1(n9538), .B2(n9537), .A(n9536), .ZN(n9541) );
  AOI222_X1 U10755 ( .A1(n10355), .A2(n9541), .B1(n9540), .B2(n10254), .C1(
        n9539), .C2(n10252), .ZN(n9703) );
  INV_X1 U10756 ( .A(n9703), .ZN(n9542) );
  AOI211_X1 U10757 ( .C1(n9700), .C2(n9544), .A(n9543), .B(n9542), .ZN(n9550)
         );
  AOI22_X1 U10758 ( .A1(n9701), .A2(n9648), .B1(P1_REG2_REG_21__SCAN_IN), .B2(
        n10362), .ZN(n9549) );
  OR2_X1 U10759 ( .A1(n9546), .A2(n9545), .ZN(n9699) );
  NAND3_X1 U10760 ( .A1(n9699), .A2(n9698), .A3(n9547), .ZN(n9548) );
  OAI211_X1 U10761 ( .C1(n9550), .C2(n10362), .A(n9549), .B(n9548), .ZN(
        P1_U3270) );
  XOR2_X1 U10762 ( .A(n9560), .B(n9551), .Z(n9709) );
  INV_X1 U10763 ( .A(n9574), .ZN(n9553) );
  AOI211_X1 U10764 ( .C1(n9707), .C2(n9553), .A(n10388), .B(n4699), .ZN(n9706)
         );
  NOR2_X1 U10765 ( .A1(n9554), .A2(n10364), .ZN(n9559) );
  OAI22_X1 U10766 ( .A1(n10366), .A2(n9557), .B1(n9556), .B2(n9555), .ZN(n9558) );
  AOI211_X1 U10767 ( .C1(n9706), .C2(n9626), .A(n9559), .B(n9558), .ZN(n9566)
         );
  XNOR2_X1 U10768 ( .A(n9561), .B(n9560), .ZN(n9562) );
  OAI222_X1 U10769 ( .A1(n10352), .A2(n9564), .B1(n10350), .B2(n9563), .C1(
        n9562), .C2(n9620), .ZN(n9705) );
  NAND2_X1 U10770 ( .A1(n9705), .A2(n10366), .ZN(n9565) );
  OAI211_X1 U10771 ( .C1(n9709), .C2(n9633), .A(n9566), .B(n9565), .ZN(
        P1_U3271) );
  XNOR2_X1 U10772 ( .A(n9568), .B(n9567), .ZN(n9714) );
  XNOR2_X1 U10773 ( .A(n9570), .B(n9569), .ZN(n9571) );
  OAI222_X1 U10774 ( .A1(n10352), .A2(n9573), .B1(n10350), .B2(n9572), .C1(
        n9571), .C2(n9620), .ZN(n9710) );
  INV_X1 U10775 ( .A(n9584), .ZN(n9575) );
  AOI211_X1 U10776 ( .C1(n9712), .C2(n9575), .A(n10388), .B(n9574), .ZN(n9711)
         );
  NAND2_X1 U10777 ( .A1(n9711), .A2(n9626), .ZN(n9579) );
  INV_X1 U10778 ( .A(n9576), .ZN(n9577) );
  AOI22_X1 U10779 ( .A1(n10362), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9577), 
        .B2(n10360), .ZN(n9578) );
  OAI211_X1 U10780 ( .C1(n9580), .C2(n10364), .A(n9579), .B(n9578), .ZN(n9581)
         );
  AOI21_X1 U10781 ( .B1(n9710), .B2(n10366), .A(n9581), .ZN(n9582) );
  OAI21_X1 U10782 ( .B1(n9714), .B2(n9633), .A(n9582), .ZN(P1_U3272) );
  XNOR2_X1 U10783 ( .A(n9583), .B(n9591), .ZN(n9719) );
  AOI21_X1 U10784 ( .B1(n9715), .B2(n9599), .A(n9584), .ZN(n9716) );
  AOI22_X1 U10785 ( .A1(n10362), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9585), 
        .B2(n10360), .ZN(n9586) );
  OAI21_X1 U10786 ( .B1(n4703), .B2(n10364), .A(n9586), .ZN(n9596) );
  INV_X1 U10787 ( .A(n9587), .ZN(n9588) );
  NOR2_X1 U10788 ( .A1(n9589), .A2(n9588), .ZN(n9590) );
  XOR2_X1 U10789 ( .A(n9591), .B(n9590), .Z(n9594) );
  AOI222_X1 U10790 ( .A1(n10355), .A2(n9594), .B1(n9593), .B2(n10252), .C1(
        n9592), .C2(n10254), .ZN(n9718) );
  NOR2_X1 U10791 ( .A1(n9718), .A2(n10362), .ZN(n9595) );
  AOI211_X1 U10792 ( .C1(n9716), .C2(n10343), .A(n9596), .B(n9595), .ZN(n9597)
         );
  OAI21_X1 U10793 ( .B1(n9633), .B2(n9719), .A(n9597), .ZN(P1_U3273) );
  XOR2_X1 U10794 ( .A(n9605), .B(n9598), .Z(n9725) );
  INV_X1 U10795 ( .A(n9599), .ZN(n9600) );
  AOI21_X1 U10796 ( .B1(n9720), .B2(n9623), .A(n9600), .ZN(n9722) );
  AOI22_X1 U10797 ( .A1(n10362), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9601), 
        .B2(n10360), .ZN(n9602) );
  OAI21_X1 U10798 ( .B1(n9603), .B2(n10364), .A(n9602), .ZN(n9610) );
  XOR2_X1 U10799 ( .A(n9605), .B(n9604), .Z(n9608) );
  AOI222_X1 U10800 ( .A1(n10355), .A2(n9608), .B1(n9607), .B2(n10254), .C1(
        n9606), .C2(n10252), .ZN(n9724) );
  NOR2_X1 U10801 ( .A1(n9724), .A2(n10362), .ZN(n9609) );
  AOI211_X1 U10802 ( .C1(n9722), .C2(n10343), .A(n9610), .B(n9609), .ZN(n9611)
         );
  OAI21_X1 U10803 ( .B1(n9633), .B2(n9725), .A(n9611), .ZN(P1_U3274) );
  AOI21_X1 U10804 ( .B1(n4552), .B2(n9618), .A(n9612), .ZN(n9613) );
  INV_X1 U10805 ( .A(n9613), .ZN(n9730) );
  INV_X1 U10806 ( .A(n9614), .ZN(n9615) );
  NOR2_X1 U10807 ( .A1(n9616), .A2(n9615), .ZN(n9617) );
  XOR2_X1 U10808 ( .A(n9618), .B(n9617), .Z(n9619) );
  OAI222_X1 U10809 ( .A1(n10350), .A2(n9622), .B1(n10352), .B2(n9621), .C1(
        n9620), .C2(n9619), .ZN(n9726) );
  INV_X1 U10810 ( .A(n9645), .ZN(n9625) );
  INV_X1 U10811 ( .A(n9623), .ZN(n9624) );
  AOI211_X1 U10812 ( .C1(n9728), .C2(n9625), .A(n10388), .B(n9624), .ZN(n9727)
         );
  NAND2_X1 U10813 ( .A1(n9727), .A2(n9626), .ZN(n9629) );
  AOI22_X1 U10814 ( .A1(n10362), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9627), 
        .B2(n10360), .ZN(n9628) );
  OAI211_X1 U10815 ( .C1(n9630), .C2(n10364), .A(n9629), .B(n9628), .ZN(n9631)
         );
  AOI21_X1 U10816 ( .B1(n9726), .B2(n10366), .A(n9631), .ZN(n9632) );
  OAI21_X1 U10817 ( .B1(n9633), .B2(n9730), .A(n9632), .ZN(P1_U3275) );
  XNOR2_X1 U10818 ( .A(n9634), .B(n9637), .ZN(n9643) );
  OAI22_X1 U10819 ( .A1(n9636), .A2(n10352), .B1(n9635), .B2(n10350), .ZN(
        n9642) );
  AND2_X1 U10820 ( .A1(n9638), .A2(n9637), .ZN(n9639) );
  OR2_X1 U10821 ( .A1(n9640), .A2(n9639), .ZN(n9737) );
  NOR2_X1 U10822 ( .A1(n9737), .A2(n10358), .ZN(n9641) );
  AOI211_X1 U10823 ( .C1(n10355), .C2(n9643), .A(n9642), .B(n9641), .ZN(n9736)
         );
  INV_X1 U10824 ( .A(n9737), .ZN(n9653) );
  AND2_X1 U10825 ( .A1(n9644), .A2(n9731), .ZN(n9646) );
  OR2_X1 U10826 ( .A1(n9646), .A2(n9645), .ZN(n9733) );
  AOI22_X1 U10827 ( .A1(n10362), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n9647), 
        .B2(n10360), .ZN(n9650) );
  NAND2_X1 U10828 ( .A1(n9731), .A2(n9648), .ZN(n9649) );
  OAI211_X1 U10829 ( .C1(n9733), .C2(n9651), .A(n9650), .B(n9649), .ZN(n9652)
         );
  AOI21_X1 U10830 ( .B1(n9653), .B2(n10344), .A(n9652), .ZN(n9654) );
  OAI21_X1 U10831 ( .B1(n9736), .B2(n10362), .A(n9654), .ZN(P1_U3276) );
  AOI21_X1 U10832 ( .B1(n9655), .B2(n10372), .A(n10266), .ZN(n9656) );
  MUX2_X1 U10833 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9744), .S(n4483), .Z(
        P1_U3554) );
  NAND2_X1 U10834 ( .A1(n9658), .A2(n10279), .ZN(n9662) );
  NOR2_X1 U10835 ( .A1(n9659), .A2(n10388), .ZN(n9660) );
  MUX2_X1 U10836 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9745), .S(n4483), .Z(
        P1_U3552) );
  NAND2_X1 U10837 ( .A1(n9663), .A2(n10279), .ZN(n9668) );
  AOI22_X1 U10838 ( .A1(n9665), .A2(n9721), .B1(n10372), .B2(n9664), .ZN(n9666) );
  NAND3_X1 U10839 ( .A1(n9668), .A2(n9667), .A3(n9666), .ZN(n9746) );
  MUX2_X1 U10840 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9746), .S(n4483), .Z(
        P1_U3551) );
  AOI211_X1 U10841 ( .C1(n10372), .C2(n9671), .A(n9670), .B(n9669), .ZN(n9672)
         );
  OAI21_X1 U10842 ( .B1(n9673), .B2(n9742), .A(n9672), .ZN(n9747) );
  MUX2_X1 U10843 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9747), .S(n4483), .Z(
        P1_U3550) );
  AOI22_X1 U10844 ( .A1(n9675), .A2(n9721), .B1(n10372), .B2(n9674), .ZN(n9676) );
  OAI211_X1 U10845 ( .C1(n9678), .C2(n9742), .A(n9677), .B(n9676), .ZN(n9748)
         );
  MUX2_X1 U10846 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9748), .S(n4483), .Z(
        P1_U3549) );
  AOI211_X1 U10847 ( .C1(n10372), .C2(n9681), .A(n9680), .B(n9679), .ZN(n9682)
         );
  OAI21_X1 U10848 ( .B1(n9683), .B2(n9742), .A(n9682), .ZN(n9749) );
  MUX2_X1 U10849 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9749), .S(n4483), .Z(
        P1_U3548) );
  AOI21_X1 U10850 ( .B1(n10372), .B2(n8039), .A(n9684), .ZN(n9685) );
  OAI211_X1 U10851 ( .C1(n9687), .C2(n9742), .A(n9686), .B(n9685), .ZN(n9750)
         );
  MUX2_X1 U10852 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9750), .S(n4483), .Z(
        P1_U3547) );
  AOI211_X1 U10853 ( .C1(n10372), .C2(n9690), .A(n9689), .B(n9688), .ZN(n9691)
         );
  OAI21_X1 U10854 ( .B1(n9692), .B2(n9742), .A(n9691), .ZN(n9751) );
  MUX2_X1 U10855 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9751), .S(n4483), .Z(
        P1_U3546) );
  AOI22_X1 U10856 ( .A1(n9694), .A2(n9721), .B1(n10372), .B2(n9693), .ZN(n9695) );
  OAI211_X1 U10857 ( .C1(n9697), .C2(n9742), .A(n9696), .B(n9695), .ZN(n9752)
         );
  MUX2_X1 U10858 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9752), .S(n4483), .Z(
        P1_U3545) );
  NAND3_X1 U10859 ( .A1(n9699), .A2(n9698), .A3(n10279), .ZN(n9704) );
  AOI21_X1 U10860 ( .B1(n10372), .B2(n9701), .A(n9700), .ZN(n9702) );
  NAND3_X1 U10861 ( .A1(n9704), .A2(n9703), .A3(n9702), .ZN(n9753) );
  MUX2_X1 U10862 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9753), .S(n4483), .Z(
        P1_U3544) );
  AOI211_X1 U10863 ( .C1(n10372), .C2(n9707), .A(n9706), .B(n9705), .ZN(n9708)
         );
  OAI21_X1 U10864 ( .B1(n9709), .B2(n9742), .A(n9708), .ZN(n9754) );
  MUX2_X1 U10865 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9754), .S(n4483), .Z(
        P1_U3543) );
  AOI211_X1 U10866 ( .C1(n10372), .C2(n9712), .A(n9711), .B(n9710), .ZN(n9713)
         );
  OAI21_X1 U10867 ( .B1(n9714), .B2(n9742), .A(n9713), .ZN(n9755) );
  MUX2_X1 U10868 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9755), .S(n4483), .Z(
        P1_U3542) );
  AOI22_X1 U10869 ( .A1(n9716), .A2(n9721), .B1(n10372), .B2(n9715), .ZN(n9717) );
  OAI211_X1 U10870 ( .C1(n9719), .C2(n9742), .A(n9718), .B(n9717), .ZN(n9756)
         );
  MUX2_X1 U10871 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9756), .S(n4483), .Z(
        P1_U3541) );
  AOI22_X1 U10872 ( .A1(n9722), .A2(n9721), .B1(n10372), .B2(n9720), .ZN(n9723) );
  OAI211_X1 U10873 ( .C1(n9725), .C2(n9742), .A(n9724), .B(n9723), .ZN(n9757)
         );
  MUX2_X1 U10874 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9757), .S(n4483), .Z(
        P1_U3540) );
  AOI211_X1 U10875 ( .C1(n10372), .C2(n9728), .A(n9727), .B(n9726), .ZN(n9729)
         );
  OAI21_X1 U10876 ( .B1(n9742), .B2(n9730), .A(n9729), .ZN(n9758) );
  MUX2_X1 U10877 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9758), .S(n4483), .Z(
        P1_U3539) );
  INV_X1 U10878 ( .A(n9731), .ZN(n9732) );
  OAI22_X1 U10879 ( .A1(n9733), .A2(n10388), .B1(n9732), .B2(n10386), .ZN(
        n9734) );
  INV_X1 U10880 ( .A(n9734), .ZN(n9735) );
  OAI211_X1 U10881 ( .C1(n10375), .C2(n9737), .A(n9736), .B(n9735), .ZN(n9759)
         );
  MUX2_X1 U10882 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n9759), .S(n4483), .Z(
        P1_U3538) );
  AOI21_X1 U10883 ( .B1(n10372), .B2(n9739), .A(n9738), .ZN(n9740) );
  OAI211_X1 U10884 ( .C1(n9743), .C2(n9742), .A(n9741), .B(n9740), .ZN(n9760)
         );
  MUX2_X1 U10885 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n9760), .S(n4483), .Z(
        P1_U3537) );
  MUX2_X1 U10886 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9744), .S(n10396), .Z(
        P1_U3522) );
  MUX2_X1 U10887 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9746), .S(n10396), .Z(
        P1_U3519) );
  MUX2_X1 U10888 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9747), .S(n10396), .Z(
        P1_U3518) );
  MUX2_X1 U10889 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9748), .S(n10396), .Z(
        P1_U3517) );
  MUX2_X1 U10890 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9749), .S(n10396), .Z(
        P1_U3516) );
  MUX2_X1 U10891 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9750), .S(n10396), .Z(
        P1_U3515) );
  MUX2_X1 U10892 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9751), .S(n10396), .Z(
        P1_U3514) );
  MUX2_X1 U10893 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9752), .S(n10396), .Z(
        P1_U3513) );
  MUX2_X1 U10894 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9753), .S(n10396), .Z(
        P1_U3512) );
  MUX2_X1 U10895 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9754), .S(n10396), .Z(
        P1_U3511) );
  MUX2_X1 U10896 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9755), .S(n10396), .Z(
        P1_U3510) );
  MUX2_X1 U10897 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9756), .S(n10396), .Z(
        P1_U3508) );
  MUX2_X1 U10898 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9757), .S(n10396), .Z(
        P1_U3505) );
  MUX2_X1 U10899 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9758), .S(n10396), .Z(
        P1_U3502) );
  MUX2_X1 U10900 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n9759), .S(n10396), .Z(
        P1_U3499) );
  MUX2_X1 U10901 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n9760), .S(n10396), .Z(
        P1_U3496) );
  INV_X1 U10902 ( .A(n9761), .ZN(n9763) );
  AND2_X1 U10903 ( .A1(n9763), .A2(n9762), .ZN(n10370) );
  MUX2_X1 U10904 ( .A(P1_D_REG_0__SCAN_IN), .B(n9764), .S(n10370), .Z(P1_U3440) );
  NAND3_X1 U10905 ( .A1(n6135), .A2(P1_STATE_REG_SCAN_IN), .A3(
        P1_IR_REG_31__SCAN_IN), .ZN(n9765) );
  OAI22_X1 U10906 ( .A1(n9766), .A2(n9765), .B1(n5910), .B2(n9774), .ZN(n9767)
         );
  AOI21_X1 U10907 ( .B1(n9769), .B2(n9768), .A(n9767), .ZN(n9770) );
  INV_X1 U10908 ( .A(n9770), .ZN(P1_U3322) );
  OAI222_X1 U10909 ( .A1(n9774), .A2(n9890), .B1(n9773), .B2(n9772), .C1(
        P1_U3084), .C2(n9771), .ZN(P1_U3323) );
  MUX2_X1 U10910 ( .A(n9775), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  NOR2_X1 U10911 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n9776) );
  AOI21_X1 U10912 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n9776), .ZN(n10514) );
  NOR2_X1 U10913 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n9777) );
  AOI21_X1 U10914 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n9777), .ZN(n10517) );
  NOR2_X1 U10915 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n9778) );
  AOI21_X1 U10916 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n9778), .ZN(n10520) );
  NOR2_X1 U10917 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n9779) );
  AOI21_X1 U10918 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n9779), .ZN(n10523) );
  NOR2_X1 U10919 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n9780) );
  AOI21_X1 U10920 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n9780), .ZN(n10526) );
  NOR2_X1 U10921 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n9786) );
  XNOR2_X1 U10922 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10553) );
  NAND2_X1 U10923 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n9784) );
  XOR2_X1 U10924 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10551) );
  NAND2_X1 U10925 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n9782) );
  XOR2_X1 U10926 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(P1_ADDR_REG_2__SCAN_IN), .Z(
        n10541) );
  AOI21_X1 U10927 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10507) );
  NAND3_X1 U10928 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n10509) );
  OAI21_X1 U10929 ( .B1(n10507), .B2(n10511), .A(n10509), .ZN(n10540) );
  NAND2_X1 U10930 ( .A1(n10541), .A2(n10540), .ZN(n9781) );
  NAND2_X1 U10931 ( .A1(n9782), .A2(n9781), .ZN(n10550) );
  NAND2_X1 U10932 ( .A1(n10551), .A2(n10550), .ZN(n9783) );
  NAND2_X1 U10933 ( .A1(n9784), .A2(n9783), .ZN(n10552) );
  NOR2_X1 U10934 ( .A1(n10553), .A2(n10552), .ZN(n9785) );
  NOR2_X1 U10935 ( .A1(n9786), .A2(n9785), .ZN(n9787) );
  NOR2_X1 U10936 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n9787), .ZN(n10543) );
  AND2_X1 U10937 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n9787), .ZN(n10542) );
  NOR2_X1 U10938 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10542), .ZN(n9788) );
  NOR2_X1 U10939 ( .A1(n10543), .A2(n9788), .ZN(n9789) );
  NAND2_X1 U10940 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(n9789), .ZN(n9791) );
  XOR2_X1 U10941 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(n9789), .Z(n10549) );
  NAND2_X1 U10942 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(n10549), .ZN(n9790) );
  NAND2_X1 U10943 ( .A1(n9791), .A2(n9790), .ZN(n9792) );
  NAND2_X1 U10944 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n9792), .ZN(n9795) );
  XNOR2_X1 U10945 ( .A(n9793), .B(n9792), .ZN(n10539) );
  NAND2_X1 U10946 ( .A1(n10539), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n9794) );
  NAND2_X1 U10947 ( .A1(n9795), .A2(n9794), .ZN(n9796) );
  NAND2_X1 U10948 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n9796), .ZN(n9798) );
  XOR2_X1 U10949 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n9796), .Z(n10548) );
  NAND2_X1 U10950 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n10548), .ZN(n9797) );
  NAND2_X1 U10951 ( .A1(n9798), .A2(n9797), .ZN(n9799) );
  AND2_X1 U10952 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n9799), .ZN(n9800) );
  XNOR2_X1 U10953 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n9799), .ZN(n10538) );
  INV_X1 U10954 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10537) );
  NOR2_X1 U10955 ( .A1(n10538), .A2(n10537), .ZN(n10536) );
  NAND2_X1 U10956 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n9801) );
  OAI21_X1 U10957 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n9801), .ZN(n10534) );
  AOI21_X1 U10958 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10533), .ZN(n10532) );
  NAND2_X1 U10959 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n9802) );
  OAI21_X1 U10960 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n9802), .ZN(n10531) );
  NOR2_X1 U10961 ( .A1(n10532), .A2(n10531), .ZN(n10530) );
  AOI21_X1 U10962 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10530), .ZN(n10529) );
  NOR2_X1 U10963 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n9803) );
  AOI21_X1 U10964 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n9803), .ZN(n10528) );
  NAND2_X1 U10965 ( .A1(n10529), .A2(n10528), .ZN(n10527) );
  OAI21_X1 U10966 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10527), .ZN(n10525) );
  NAND2_X1 U10967 ( .A1(n10526), .A2(n10525), .ZN(n10524) );
  OAI21_X1 U10968 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10524), .ZN(n10522) );
  NAND2_X1 U10969 ( .A1(n10523), .A2(n10522), .ZN(n10521) );
  OAI21_X1 U10970 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10521), .ZN(n10519) );
  NAND2_X1 U10971 ( .A1(n10520), .A2(n10519), .ZN(n10518) );
  OAI21_X1 U10972 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10518), .ZN(n10516) );
  NAND2_X1 U10973 ( .A1(n10517), .A2(n10516), .ZN(n10515) );
  OAI21_X1 U10974 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10515), .ZN(n10513) );
  NAND2_X1 U10975 ( .A1(n10514), .A2(n10513), .ZN(n10512) );
  OAI21_X1 U10976 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10512), .ZN(n10546) );
  NOR2_X1 U10977 ( .A1(n9381), .A2(n10546), .ZN(n9804) );
  NAND2_X1 U10978 ( .A1(n9381), .A2(n10546), .ZN(n10545) );
  OAI21_X1 U10979 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n9804), .A(n10545), .ZN(
        n10174) );
  OAI22_X1 U10980 ( .A1(P1_D_REG_2__SCAN_IN), .A2(keyinput_g125), .B1(
        keyinput_g33), .B2(P2_RD_REG_SCAN_IN), .ZN(n9805) );
  AOI221_X1 U10981 ( .B1(P1_D_REG_2__SCAN_IN), .B2(keyinput_g125), .C1(
        P2_RD_REG_SCAN_IN), .C2(keyinput_g33), .A(n9805), .ZN(n9812) );
  OAI22_X1 U10982 ( .A1(P2_DATAO_REG_24__SCAN_IN), .A2(keyinput_g72), .B1(
        SI_8_), .B2(keyinput_g24), .ZN(n9806) );
  AOI221_X1 U10983 ( .B1(P2_DATAO_REG_24__SCAN_IN), .B2(keyinput_g72), .C1(
        keyinput_g24), .C2(SI_8_), .A(n9806), .ZN(n9811) );
  OAI22_X1 U10984 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(keyinput_g112), .B1(
        P2_REG3_REG_21__SCAN_IN), .B2(keyinput_g45), .ZN(n9807) );
  AOI221_X1 U10985 ( .B1(P1_IR_REG_21__SCAN_IN), .B2(keyinput_g112), .C1(
        keyinput_g45), .C2(P2_REG3_REG_21__SCAN_IN), .A(n9807), .ZN(n9810) );
  OAI22_X1 U10986 ( .A1(P2_DATAO_REG_8__SCAN_IN), .A2(keyinput_g88), .B1(
        keyinput_g25), .B2(SI_7_), .ZN(n9808) );
  AOI221_X1 U10987 ( .B1(P2_DATAO_REG_8__SCAN_IN), .B2(keyinput_g88), .C1(
        SI_7_), .C2(keyinput_g25), .A(n9808), .ZN(n9809) );
  NAND4_X1 U10988 ( .A1(n9812), .A2(n9811), .A3(n9810), .A4(n9809), .ZN(n9840)
         );
  OAI22_X1 U10989 ( .A1(P1_IR_REG_29__SCAN_IN), .A2(keyinput_g120), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(keyinput_g54), .ZN(n9813) );
  AOI221_X1 U10990 ( .B1(P1_IR_REG_29__SCAN_IN), .B2(keyinput_g120), .C1(
        keyinput_g54), .C2(P2_REG3_REG_0__SCAN_IN), .A(n9813), .ZN(n9820) );
  OAI22_X1 U10991 ( .A1(SI_27_), .A2(keyinput_g5), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(keyinput_g70), .ZN(n9814) );
  AOI221_X1 U10992 ( .B1(SI_27_), .B2(keyinput_g5), .C1(keyinput_g70), .C2(
        P2_DATAO_REG_26__SCAN_IN), .A(n9814), .ZN(n9819) );
  OAI22_X1 U10993 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(keyinput_g79), .B1(
        P2_REG3_REG_15__SCAN_IN), .B2(keyinput_g63), .ZN(n9815) );
  AOI221_X1 U10994 ( .B1(P2_DATAO_REG_17__SCAN_IN), .B2(keyinput_g79), .C1(
        keyinput_g63), .C2(P2_REG3_REG_15__SCAN_IN), .A(n9815), .ZN(n9818) );
  OAI22_X1 U10995 ( .A1(SI_11_), .A2(keyinput_g21), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(keyinput_g86), .ZN(n9816) );
  AOI221_X1 U10996 ( .B1(SI_11_), .B2(keyinput_g21), .C1(keyinput_g86), .C2(
        P2_DATAO_REG_10__SCAN_IN), .A(n9816), .ZN(n9817) );
  NAND4_X1 U10997 ( .A1(n9820), .A2(n9819), .A3(n9818), .A4(n9817), .ZN(n9839)
         );
  OAI22_X1 U10998 ( .A1(P1_D_REG_4__SCAN_IN), .A2(keyinput_g127), .B1(
        P2_REG3_REG_19__SCAN_IN), .B2(keyinput_g41), .ZN(n9821) );
  AOI221_X1 U10999 ( .B1(P1_D_REG_4__SCAN_IN), .B2(keyinput_g127), .C1(
        keyinput_g41), .C2(P2_REG3_REG_19__SCAN_IN), .A(n9821), .ZN(n9828) );
  OAI22_X1 U11000 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(keyinput_g102), .B1(
        keyinput_g99), .B2(P1_IR_REG_8__SCAN_IN), .ZN(n9822) );
  AOI221_X1 U11001 ( .B1(P1_IR_REG_11__SCAN_IN), .B2(keyinput_g102), .C1(
        P1_IR_REG_8__SCAN_IN), .C2(keyinput_g99), .A(n9822), .ZN(n9827) );
  OAI22_X1 U11002 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(keyinput_g115), .B1(
        P2_REG3_REG_13__SCAN_IN), .B2(keyinput_g56), .ZN(n9823) );
  AOI221_X1 U11003 ( .B1(P1_IR_REG_24__SCAN_IN), .B2(keyinput_g115), .C1(
        keyinput_g56), .C2(P2_REG3_REG_13__SCAN_IN), .A(n9823), .ZN(n9826) );
  OAI22_X1 U11004 ( .A1(SI_20_), .A2(keyinput_g12), .B1(keyinput_g46), .B2(
        P2_REG3_REG_12__SCAN_IN), .ZN(n9824) );
  AOI221_X1 U11005 ( .B1(SI_20_), .B2(keyinput_g12), .C1(
        P2_REG3_REG_12__SCAN_IN), .C2(keyinput_g46), .A(n9824), .ZN(n9825) );
  NAND4_X1 U11006 ( .A1(n9828), .A2(n9827), .A3(n9826), .A4(n9825), .ZN(n9838)
         );
  OAI22_X1 U11007 ( .A1(SI_6_), .A2(keyinput_g26), .B1(SI_5_), .B2(
        keyinput_g27), .ZN(n9829) );
  AOI221_X1 U11008 ( .B1(SI_6_), .B2(keyinput_g26), .C1(keyinput_g27), .C2(
        SI_5_), .A(n9829), .ZN(n9836) );
  OAI22_X1 U11009 ( .A1(SI_25_), .A2(keyinput_g7), .B1(keyinput_g18), .B2(
        SI_14_), .ZN(n9830) );
  AOI221_X1 U11010 ( .B1(SI_25_), .B2(keyinput_g7), .C1(SI_14_), .C2(
        keyinput_g18), .A(n9830), .ZN(n9835) );
  OAI22_X1 U11011 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(keyinput_g100), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(keyinput_g82), .ZN(n9831) );
  AOI221_X1 U11012 ( .B1(P1_IR_REG_9__SCAN_IN), .B2(keyinput_g100), .C1(
        keyinput_g82), .C2(P2_DATAO_REG_14__SCAN_IN), .A(n9831), .ZN(n9834) );
  OAI22_X1 U11013 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(keyinput_g69), .B1(
        P2_REG3_REG_6__SCAN_IN), .B2(keyinput_g61), .ZN(n9832) );
  AOI221_X1 U11014 ( .B1(P2_DATAO_REG_27__SCAN_IN), .B2(keyinput_g69), .C1(
        keyinput_g61), .C2(P2_REG3_REG_6__SCAN_IN), .A(n9832), .ZN(n9833) );
  NAND4_X1 U11015 ( .A1(n9836), .A2(n9835), .A3(n9834), .A4(n9833), .ZN(n9837)
         );
  NOR4_X1 U11016 ( .A1(n9840), .A2(n9839), .A3(n9838), .A4(n9837), .ZN(n10172)
         );
  OAI22_X1 U11017 ( .A1(SI_21_), .A2(keyinput_g11), .B1(P2_STATE_REG_SCAN_IN), 
        .B2(keyinput_g34), .ZN(n9841) );
  AOI221_X1 U11018 ( .B1(SI_21_), .B2(keyinput_g11), .C1(keyinput_g34), .C2(
        P2_STATE_REG_SCAN_IN), .A(n9841), .ZN(n9848) );
  OAI22_X1 U11019 ( .A1(P2_DATAO_REG_11__SCAN_IN), .A2(keyinput_g85), .B1(
        keyinput_g42), .B2(P2_REG3_REG_28__SCAN_IN), .ZN(n9842) );
  AOI221_X1 U11020 ( .B1(P2_DATAO_REG_11__SCAN_IN), .B2(keyinput_g85), .C1(
        P2_REG3_REG_28__SCAN_IN), .C2(keyinput_g42), .A(n9842), .ZN(n9847) );
  OAI22_X1 U11021 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(keyinput_g110), .B1(SI_15_), .B2(keyinput_g17), .ZN(n9843) );
  AOI221_X1 U11022 ( .B1(P1_IR_REG_19__SCAN_IN), .B2(keyinput_g110), .C1(
        keyinput_g17), .C2(SI_15_), .A(n9843), .ZN(n9846) );
  OAI22_X1 U11023 ( .A1(P2_REG3_REG_23__SCAN_IN), .A2(keyinput_g38), .B1(
        P2_REG3_REG_16__SCAN_IN), .B2(keyinput_g48), .ZN(n9844) );
  AOI221_X1 U11024 ( .B1(P2_REG3_REG_23__SCAN_IN), .B2(keyinput_g38), .C1(
        keyinput_g48), .C2(P2_REG3_REG_16__SCAN_IN), .A(n9844), .ZN(n9845) );
  NAND4_X1 U11025 ( .A1(n9848), .A2(n9847), .A3(n9846), .A4(n9845), .ZN(n9979)
         );
  AOI22_X1 U11026 ( .A1(SI_30_), .A2(keyinput_g2), .B1(P2_B_REG_SCAN_IN), .B2(
        keyinput_g64), .ZN(n9849) );
  OAI221_X1 U11027 ( .B1(SI_30_), .B2(keyinput_g2), .C1(P2_B_REG_SCAN_IN), 
        .C2(keyinput_g64), .A(n9849), .ZN(n9856) );
  AOI22_X1 U11028 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(keyinput_g49), .B1(
        P2_REG3_REG_11__SCAN_IN), .B2(keyinput_g58), .ZN(n9850) );
  OAI221_X1 U11029 ( .B1(P2_REG3_REG_5__SCAN_IN), .B2(keyinput_g49), .C1(
        P2_REG3_REG_11__SCAN_IN), .C2(keyinput_g58), .A(n9850), .ZN(n9855) );
  AOI22_X1 U11030 ( .A1(P2_REG3_REG_2__SCAN_IN), .A2(keyinput_g59), .B1(SI_28_), .B2(keyinput_g4), .ZN(n9851) );
  OAI221_X1 U11031 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(keyinput_g59), .C1(
        SI_28_), .C2(keyinput_g4), .A(n9851), .ZN(n9854) );
  AOI22_X1 U11032 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(keyinput_g43), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(keyinput_g75), .ZN(n9852) );
  OAI221_X1 U11033 ( .B1(P2_REG3_REG_8__SCAN_IN), .B2(keyinput_g43), .C1(
        P2_DATAO_REG_21__SCAN_IN), .C2(keyinput_g75), .A(n9852), .ZN(n9853) );
  NOR4_X1 U11034 ( .A1(n9856), .A2(n9855), .A3(n9854), .A4(n9853), .ZN(n9874)
         );
  AOI22_X1 U11035 ( .A1(P2_DATAO_REG_22__SCAN_IN), .A2(keyinput_g74), .B1(
        P1_D_REG_1__SCAN_IN), .B2(keyinput_g124), .ZN(n9857) );
  OAI221_X1 U11036 ( .B1(P2_DATAO_REG_22__SCAN_IN), .B2(keyinput_g74), .C1(
        P1_D_REG_1__SCAN_IN), .C2(keyinput_g124), .A(n9857), .ZN(n9864) );
  AOI22_X1 U11037 ( .A1(P2_WR_REG_SCAN_IN), .A2(keyinput_g0), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(keyinput_g80), .ZN(n9858) );
  OAI221_X1 U11038 ( .B1(P2_WR_REG_SCAN_IN), .B2(keyinput_g0), .C1(
        P2_DATAO_REG_16__SCAN_IN), .C2(keyinput_g80), .A(n9858), .ZN(n9863) );
  AOI22_X1 U11039 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(keyinput_g60), .B1(
        P1_IR_REG_0__SCAN_IN), .B2(keyinput_g91), .ZN(n9859) );
  OAI221_X1 U11040 ( .B1(P2_REG3_REG_18__SCAN_IN), .B2(keyinput_g60), .C1(
        P1_IR_REG_0__SCAN_IN), .C2(keyinput_g91), .A(n9859), .ZN(n9862) );
  AOI22_X1 U11041 ( .A1(P2_DATAO_REG_31__SCAN_IN), .A2(keyinput_g65), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(keyinput_g68), .ZN(n9860) );
  OAI221_X1 U11042 ( .B1(P2_DATAO_REG_31__SCAN_IN), .B2(keyinput_g65), .C1(
        P2_DATAO_REG_28__SCAN_IN), .C2(keyinput_g68), .A(n9860), .ZN(n9861) );
  NOR4_X1 U11043 ( .A1(n9864), .A2(n9863), .A3(n9862), .A4(n9861), .ZN(n9873)
         );
  OAI22_X1 U11044 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(keyinput_g108), .B1(
        P2_REG3_REG_24__SCAN_IN), .B2(keyinput_g51), .ZN(n9865) );
  AOI221_X1 U11045 ( .B1(P1_IR_REG_17__SCAN_IN), .B2(keyinput_g108), .C1(
        keyinput_g51), .C2(P2_REG3_REG_24__SCAN_IN), .A(n9865), .ZN(n9871) );
  OAI22_X1 U11046 ( .A1(P1_D_REG_0__SCAN_IN), .A2(keyinput_g123), .B1(
        keyinput_g30), .B2(SI_2_), .ZN(n9866) );
  AOI221_X1 U11047 ( .B1(P1_D_REG_0__SCAN_IN), .B2(keyinput_g123), .C1(SI_2_), 
        .C2(keyinput_g30), .A(n9866), .ZN(n9870) );
  OAI22_X1 U11048 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(keyinput_g103), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(keyinput_g78), .ZN(n9867) );
  AOI221_X1 U11049 ( .B1(P1_IR_REG_12__SCAN_IN), .B2(keyinput_g103), .C1(
        keyinput_g78), .C2(P2_DATAO_REG_18__SCAN_IN), .A(n9867), .ZN(n9869) );
  XNOR2_X1 U11050 ( .A(P1_IR_REG_30__SCAN_IN), .B(keyinput_g121), .ZN(n9868)
         );
  AND4_X1 U11051 ( .A1(n9871), .A2(n9870), .A3(n9869), .A4(n9868), .ZN(n9872)
         );
  NAND3_X1 U11052 ( .A1(n9874), .A2(n9873), .A3(n9872), .ZN(n9978) );
  AOI22_X1 U11053 ( .A1(n9876), .A2(keyinput_g84), .B1(keyinput_g39), .B2(
        n10062), .ZN(n9875) );
  OAI221_X1 U11054 ( .B1(n9876), .B2(keyinput_g84), .C1(n10062), .C2(
        keyinput_g39), .A(n9875), .ZN(n9879) );
  AOI22_X1 U11055 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(keyinput_g94), .B1(
        P1_IR_REG_18__SCAN_IN), .B2(keyinput_g109), .ZN(n9877) );
  OAI221_X1 U11056 ( .B1(P1_IR_REG_3__SCAN_IN), .B2(keyinput_g94), .C1(
        P1_IR_REG_18__SCAN_IN), .C2(keyinput_g109), .A(n9877), .ZN(n9878) );
  NOR2_X1 U11057 ( .A1(n9879), .A2(n9878), .ZN(n9886) );
  INV_X1 U11058 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n10369) );
  INV_X1 U11059 ( .A(keyinput_g126), .ZN(n9880) );
  XNOR2_X1 U11060 ( .A(n10369), .B(n9880), .ZN(n9885) );
  XNOR2_X1 U11061 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput_g122), .ZN(n9884)
         );
  AOI22_X1 U11062 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(keyinput_g117), .B1(
        P1_IR_REG_13__SCAN_IN), .B2(keyinput_g104), .ZN(n9881) );
  OAI221_X1 U11063 ( .B1(P1_IR_REG_26__SCAN_IN), .B2(keyinput_g117), .C1(
        P1_IR_REG_13__SCAN_IN), .C2(keyinput_g104), .A(n9881), .ZN(n9882) );
  INV_X1 U11064 ( .A(n9882), .ZN(n9883) );
  AND4_X1 U11065 ( .A1(n9886), .A2(n9885), .A3(n9884), .A4(n9883), .ZN(n9927)
         );
  AOI22_X1 U11066 ( .A1(n8104), .A2(keyinput_g47), .B1(keyinput_g3), .B2(n7591), .ZN(n9887) );
  OAI221_X1 U11067 ( .B1(n8104), .B2(keyinput_g47), .C1(n7591), .C2(
        keyinput_g3), .A(n9887), .ZN(n9899) );
  INV_X1 U11068 ( .A(SI_31_), .ZN(n9889) );
  AOI22_X1 U11069 ( .A1(n9890), .A2(keyinput_g66), .B1(n9889), .B2(keyinput_g1), .ZN(n9888) );
  OAI221_X1 U11070 ( .B1(n9890), .B2(keyinput_g66), .C1(n9889), .C2(
        keyinput_g1), .A(n9888), .ZN(n9898) );
  INV_X1 U11071 ( .A(SI_18_), .ZN(n9893) );
  AOI22_X1 U11072 ( .A1(n9893), .A2(keyinput_g14), .B1(keyinput_g23), .B2(
        n9892), .ZN(n9891) );
  OAI221_X1 U11073 ( .B1(n9893), .B2(keyinput_g14), .C1(n9892), .C2(
        keyinput_g23), .A(n9891), .ZN(n9897) );
  XNOR2_X1 U11074 ( .A(P1_IR_REG_23__SCAN_IN), .B(keyinput_g114), .ZN(n9895)
         );
  XNOR2_X1 U11075 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(keyinput_g89), .ZN(n9894)
         );
  NAND2_X1 U11076 ( .A1(n9895), .A2(n9894), .ZN(n9896) );
  NOR4_X1 U11077 ( .A1(n9899), .A2(n9898), .A3(n9897), .A4(n9896), .ZN(n9926)
         );
  AOI22_X1 U11078 ( .A1(n9902), .A2(keyinput_g87), .B1(keyinput_g55), .B2(
        n9901), .ZN(n9900) );
  OAI221_X1 U11079 ( .B1(n9902), .B2(keyinput_g87), .C1(n9901), .C2(
        keyinput_g55), .A(n9900), .ZN(n9913) );
  AOI22_X1 U11080 ( .A1(n5368), .A2(keyinput_g53), .B1(n9904), .B2(
        keyinput_g36), .ZN(n9903) );
  OAI221_X1 U11081 ( .B1(n5368), .B2(keyinput_g53), .C1(n9904), .C2(
        keyinput_g36), .A(n9903), .ZN(n9912) );
  AOI22_X1 U11082 ( .A1(n9907), .A2(keyinput_g77), .B1(keyinput_g15), .B2(
        n9906), .ZN(n9905) );
  OAI221_X1 U11083 ( .B1(n9907), .B2(keyinput_g77), .C1(n9906), .C2(
        keyinput_g15), .A(n9905), .ZN(n9911) );
  XNOR2_X1 U11084 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput_g92), .ZN(n9909) );
  XNOR2_X1 U11085 ( .A(SI_10_), .B(keyinput_g22), .ZN(n9908) );
  NAND2_X1 U11086 ( .A1(n9909), .A2(n9908), .ZN(n9910) );
  NOR4_X1 U11087 ( .A1(n9913), .A2(n9912), .A3(n9911), .A4(n9910), .ZN(n9925)
         );
  XNOR2_X1 U11088 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput_g111), .ZN(n9917)
         );
  XNOR2_X1 U11089 ( .A(SI_13_), .B(keyinput_g19), .ZN(n9916) );
  XNOR2_X1 U11090 ( .A(P1_IR_REG_10__SCAN_IN), .B(keyinput_g101), .ZN(n9915)
         );
  XNOR2_X1 U11091 ( .A(P2_REG3_REG_14__SCAN_IN), .B(keyinput_g37), .ZN(n9914)
         );
  NAND4_X1 U11092 ( .A1(n9917), .A2(n9916), .A3(n9915), .A4(n9914), .ZN(n9923)
         );
  XNOR2_X1 U11093 ( .A(P1_IR_REG_25__SCAN_IN), .B(keyinput_g116), .ZN(n9921)
         );
  XNOR2_X1 U11094 ( .A(SI_4_), .B(keyinput_g28), .ZN(n9920) );
  XNOR2_X1 U11095 ( .A(P1_IR_REG_27__SCAN_IN), .B(keyinput_g118), .ZN(n9919)
         );
  XNOR2_X1 U11096 ( .A(SI_22_), .B(keyinput_g10), .ZN(n9918) );
  NAND4_X1 U11097 ( .A1(n9921), .A2(n9920), .A3(n9919), .A4(n9918), .ZN(n9922)
         );
  NOR2_X1 U11098 ( .A1(n9923), .A2(n9922), .ZN(n9924) );
  NAND4_X1 U11099 ( .A1(n9927), .A2(n9926), .A3(n9925), .A4(n9924), .ZN(n9977)
         );
  AOI22_X1 U11100 ( .A1(n9930), .A2(keyinput_g90), .B1(keyinput_g35), .B2(
        n9929), .ZN(n9928) );
  OAI221_X1 U11101 ( .B1(n9930), .B2(keyinput_g90), .C1(n9929), .C2(
        keyinput_g35), .A(n9928), .ZN(n9938) );
  AOI22_X1 U11102 ( .A1(n5283), .A2(keyinput_g40), .B1(n10150), .B2(
        keyinput_g20), .ZN(n9931) );
  OAI221_X1 U11103 ( .B1(n5283), .B2(keyinput_g40), .C1(n10150), .C2(
        keyinput_g20), .A(n9931), .ZN(n9937) );
  AOI22_X1 U11104 ( .A1(n10079), .A2(keyinput_g67), .B1(n10083), .B2(
        keyinput_g13), .ZN(n9932) );
  OAI221_X1 U11105 ( .B1(n10079), .B2(keyinput_g67), .C1(n10083), .C2(
        keyinput_g13), .A(n9932), .ZN(n9936) );
  XNOR2_X1 U11106 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput_g119), .ZN(n9934)
         );
  XNOR2_X1 U11107 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(keyinput_g73), .ZN(n9933)
         );
  NAND2_X1 U11108 ( .A1(n9934), .A2(n9933), .ZN(n9935) );
  NOR4_X1 U11109 ( .A1(n9938), .A2(n9937), .A3(n9936), .A4(n9935), .ZN(n9975)
         );
  INV_X1 U11110 ( .A(SI_24_), .ZN(n9940) );
  AOI22_X1 U11111 ( .A1(n9940), .A2(keyinput_g8), .B1(keyinput_g76), .B2(
        n10077), .ZN(n9939) );
  OAI221_X1 U11112 ( .B1(n9940), .B2(keyinput_g8), .C1(n10077), .C2(
        keyinput_g76), .A(n9939), .ZN(n9949) );
  AOI22_X1 U11113 ( .A1(n10133), .A2(keyinput_g16), .B1(keyinput_g62), .B2(
        n10151), .ZN(n9941) );
  OAI221_X1 U11114 ( .B1(n10133), .B2(keyinput_g16), .C1(n10151), .C2(
        keyinput_g62), .A(n9941), .ZN(n9948) );
  AOI22_X1 U11115 ( .A1(n9943), .A2(keyinput_g83), .B1(n10145), .B2(
        keyinput_g97), .ZN(n9942) );
  OAI221_X1 U11116 ( .B1(n9943), .B2(keyinput_g83), .C1(n10145), .C2(
        keyinput_g97), .A(n9942), .ZN(n9947) );
  XNOR2_X1 U11117 ( .A(P1_IR_REG_15__SCAN_IN), .B(keyinput_g106), .ZN(n9945)
         );
  XNOR2_X1 U11118 ( .A(keyinput_g44), .B(P2_REG3_REG_1__SCAN_IN), .ZN(n9944)
         );
  NAND2_X1 U11119 ( .A1(n9945), .A2(n9944), .ZN(n9946) );
  NOR4_X1 U11120 ( .A1(n9949), .A2(n9948), .A3(n9947), .A4(n9946), .ZN(n9974)
         );
  XNOR2_X1 U11121 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput_g98), .ZN(n9953) );
  XNOR2_X1 U11122 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput_g95), .ZN(n9952) );
  XNOR2_X1 U11123 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(keyinput_g71), .ZN(n9951)
         );
  XNOR2_X1 U11124 ( .A(SI_0_), .B(keyinput_g32), .ZN(n9950) );
  NAND4_X1 U11125 ( .A1(n9953), .A2(n9952), .A3(n9951), .A4(n9950), .ZN(n9959)
         );
  XNOR2_X1 U11126 ( .A(P2_REG3_REG_17__SCAN_IN), .B(keyinput_g50), .ZN(n9957)
         );
  XNOR2_X1 U11127 ( .A(SI_3_), .B(keyinput_g29), .ZN(n9956) );
  XNOR2_X1 U11128 ( .A(P1_IR_REG_16__SCAN_IN), .B(keyinput_g107), .ZN(n9955)
         );
  XNOR2_X1 U11129 ( .A(SI_1_), .B(keyinput_g31), .ZN(n9954) );
  NAND4_X1 U11130 ( .A1(n9957), .A2(n9956), .A3(n9955), .A4(n9954), .ZN(n9958)
         );
  NOR2_X1 U11131 ( .A1(n9959), .A2(n9958), .ZN(n9973) );
  AOI22_X1 U11132 ( .A1(n9962), .A2(keyinput_g57), .B1(n9961), .B2(keyinput_g9), .ZN(n9960) );
  OAI221_X1 U11133 ( .B1(n9962), .B2(keyinput_g57), .C1(n9961), .C2(
        keyinput_g9), .A(n9960), .ZN(n9971) );
  XNOR2_X1 U11134 ( .A(SI_26_), .B(keyinput_g6), .ZN(n9966) );
  XNOR2_X1 U11135 ( .A(P1_IR_REG_14__SCAN_IN), .B(keyinput_g105), .ZN(n9965)
         );
  XNOR2_X1 U11136 ( .A(P1_IR_REG_2__SCAN_IN), .B(keyinput_g93), .ZN(n9964) );
  XNOR2_X1 U11137 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput_g96), .ZN(n9963) );
  NAND4_X1 U11138 ( .A1(n9966), .A2(n9965), .A3(n9964), .A4(n9963), .ZN(n9970)
         );
  XNOR2_X1 U11139 ( .A(n9967), .B(keyinput_g113), .ZN(n9969) );
  XNOR2_X1 U11140 ( .A(keyinput_g52), .B(n5222), .ZN(n9968) );
  NOR4_X1 U11141 ( .A1(n9971), .A2(n9970), .A3(n9969), .A4(n9968), .ZN(n9972)
         );
  NAND4_X1 U11142 ( .A1(n9975), .A2(n9974), .A3(n9973), .A4(n9972), .ZN(n9976)
         );
  NOR4_X1 U11143 ( .A1(n9979), .A2(n9978), .A3(n9977), .A4(n9976), .ZN(n10171)
         );
  AOI22_X1 U11144 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(keyinput_f56), .B1(
        P2_REG3_REG_27__SCAN_IN), .B2(keyinput_f36), .ZN(n9980) );
  OAI221_X1 U11145 ( .B1(P2_REG3_REG_13__SCAN_IN), .B2(keyinput_f56), .C1(
        P2_REG3_REG_27__SCAN_IN), .C2(keyinput_f36), .A(n9980), .ZN(n9987) );
  AOI22_X1 U11146 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(keyinput_f66), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(keyinput_f83), .ZN(n9981) );
  OAI221_X1 U11147 ( .B1(P2_DATAO_REG_30__SCAN_IN), .B2(keyinput_f66), .C1(
        P2_DATAO_REG_13__SCAN_IN), .C2(keyinput_f83), .A(n9981), .ZN(n9986) );
  AOI22_X1 U11148 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(keyinput_f48), .B1(
        P1_IR_REG_29__SCAN_IN), .B2(keyinput_f120), .ZN(n9982) );
  OAI221_X1 U11149 ( .B1(P2_REG3_REG_16__SCAN_IN), .B2(keyinput_f48), .C1(
        P1_IR_REG_29__SCAN_IN), .C2(keyinput_f120), .A(n9982), .ZN(n9985) );
  XNOR2_X1 U11150 ( .A(n9983), .B(keyinput_f95), .ZN(n9984) );
  NOR4_X1 U11151 ( .A1(n9987), .A2(n9986), .A3(n9985), .A4(n9984), .ZN(n10015)
         );
  AOI22_X1 U11152 ( .A1(P2_DATAO_REG_12__SCAN_IN), .A2(keyinput_f84), .B1(
        SI_22_), .B2(keyinput_f10), .ZN(n9988) );
  OAI221_X1 U11153 ( .B1(P2_DATAO_REG_12__SCAN_IN), .B2(keyinput_f84), .C1(
        SI_22_), .C2(keyinput_f10), .A(n9988), .ZN(n9995) );
  AOI22_X1 U11154 ( .A1(P1_D_REG_3__SCAN_IN), .A2(keyinput_f126), .B1(
        P1_IR_REG_22__SCAN_IN), .B2(keyinput_f113), .ZN(n9989) );
  OAI221_X1 U11155 ( .B1(P1_D_REG_3__SCAN_IN), .B2(keyinput_f126), .C1(
        P1_IR_REG_22__SCAN_IN), .C2(keyinput_f113), .A(n9989), .ZN(n9994) );
  AOI22_X1 U11156 ( .A1(SI_31_), .A2(keyinput_f1), .B1(P2_REG3_REG_7__SCAN_IN), 
        .B2(keyinput_f35), .ZN(n9990) );
  OAI221_X1 U11157 ( .B1(SI_31_), .B2(keyinput_f1), .C1(P2_REG3_REG_7__SCAN_IN), .C2(keyinput_f35), .A(n9990), .ZN(n9993) );
  AOI22_X1 U11158 ( .A1(P1_D_REG_1__SCAN_IN), .A2(keyinput_f124), .B1(
        P1_IR_REG_12__SCAN_IN), .B2(keyinput_f103), .ZN(n9991) );
  OAI221_X1 U11159 ( .B1(P1_D_REG_1__SCAN_IN), .B2(keyinput_f124), .C1(
        P1_IR_REG_12__SCAN_IN), .C2(keyinput_f103), .A(n9991), .ZN(n9992) );
  NOR4_X1 U11160 ( .A1(n9995), .A2(n9994), .A3(n9993), .A4(n9992), .ZN(n10014)
         );
  AOI22_X1 U11161 ( .A1(P2_REG3_REG_28__SCAN_IN), .A2(keyinput_f42), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(keyinput_f69), .ZN(n9996) );
  OAI221_X1 U11162 ( .B1(P2_REG3_REG_28__SCAN_IN), .B2(keyinput_f42), .C1(
        P2_DATAO_REG_27__SCAN_IN), .C2(keyinput_f69), .A(n9996), .ZN(n10003)
         );
  AOI22_X1 U11163 ( .A1(SI_11_), .A2(keyinput_f21), .B1(P1_IR_REG_17__SCAN_IN), 
        .B2(keyinput_f108), .ZN(n9997) );
  OAI221_X1 U11164 ( .B1(SI_11_), .B2(keyinput_f21), .C1(P1_IR_REG_17__SCAN_IN), .C2(keyinput_f108), .A(n9997), .ZN(n10002) );
  AOI22_X1 U11165 ( .A1(P2_REG3_REG_1__SCAN_IN), .A2(keyinput_f44), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(keyinput_f70), .ZN(n9998) );
  OAI221_X1 U11166 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(keyinput_f44), .C1(
        P2_DATAO_REG_26__SCAN_IN), .C2(keyinput_f70), .A(n9998), .ZN(n10001)
         );
  AOI22_X1 U11167 ( .A1(keyinput_f0), .A2(P2_WR_REG_SCAN_IN), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(keyinput_f77), .ZN(n9999) );
  OAI221_X1 U11168 ( .B1(keyinput_f0), .B2(P2_WR_REG_SCAN_IN), .C1(
        P2_DATAO_REG_19__SCAN_IN), .C2(keyinput_f77), .A(n9999), .ZN(n10000)
         );
  NOR4_X1 U11169 ( .A1(n10003), .A2(n10002), .A3(n10001), .A4(n10000), .ZN(
        n10013) );
  AOI22_X1 U11170 ( .A1(SI_27_), .A2(keyinput_f5), .B1(P1_IR_REG_9__SCAN_IN), 
        .B2(keyinput_f100), .ZN(n10004) );
  OAI221_X1 U11171 ( .B1(SI_27_), .B2(keyinput_f5), .C1(P1_IR_REG_9__SCAN_IN), 
        .C2(keyinput_f100), .A(n10004), .ZN(n10011) );
  AOI22_X1 U11172 ( .A1(SI_13_), .A2(keyinput_f19), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(keyinput_f71), .ZN(n10005) );
  OAI221_X1 U11173 ( .B1(SI_13_), .B2(keyinput_f19), .C1(
        P2_DATAO_REG_25__SCAN_IN), .C2(keyinput_f71), .A(n10005), .ZN(n10010)
         );
  AOI22_X1 U11174 ( .A1(SI_30_), .A2(keyinput_f2), .B1(SI_18_), .B2(
        keyinput_f14), .ZN(n10006) );
  OAI221_X1 U11175 ( .B1(SI_30_), .B2(keyinput_f2), .C1(SI_18_), .C2(
        keyinput_f14), .A(n10006), .ZN(n10009) );
  AOI22_X1 U11176 ( .A1(P2_REG3_REG_22__SCAN_IN), .A2(keyinput_f57), .B1(
        P1_D_REG_4__SCAN_IN), .B2(keyinput_f127), .ZN(n10007) );
  OAI221_X1 U11177 ( .B1(P2_REG3_REG_22__SCAN_IN), .B2(keyinput_f57), .C1(
        P1_D_REG_4__SCAN_IN), .C2(keyinput_f127), .A(n10007), .ZN(n10008) );
  NOR4_X1 U11178 ( .A1(n10011), .A2(n10010), .A3(n10009), .A4(n10008), .ZN(
        n10012) );
  NAND4_X1 U11179 ( .A1(n10015), .A2(n10014), .A3(n10013), .A4(n10012), .ZN(
        n10165) );
  AOI22_X1 U11180 ( .A1(P2_DATAO_REG_31__SCAN_IN), .A2(keyinput_f65), .B1(
        P2_REG3_REG_17__SCAN_IN), .B2(keyinput_f50), .ZN(n10016) );
  OAI221_X1 U11181 ( .B1(P2_DATAO_REG_31__SCAN_IN), .B2(keyinput_f65), .C1(
        P2_REG3_REG_17__SCAN_IN), .C2(keyinput_f50), .A(n10016), .ZN(n10023)
         );
  AOI22_X1 U11182 ( .A1(SI_29_), .A2(keyinput_f3), .B1(P2_REG3_REG_15__SCAN_IN), .B2(keyinput_f63), .ZN(n10017) );
  OAI221_X1 U11183 ( .B1(SI_29_), .B2(keyinput_f3), .C1(
        P2_REG3_REG_15__SCAN_IN), .C2(keyinput_f63), .A(n10017), .ZN(n10022)
         );
  AOI22_X1 U11184 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(keyinput_f117), .B1(
        P1_IR_REG_21__SCAN_IN), .B2(keyinput_f112), .ZN(n10018) );
  OAI221_X1 U11185 ( .B1(P1_IR_REG_26__SCAN_IN), .B2(keyinput_f117), .C1(
        P1_IR_REG_21__SCAN_IN), .C2(keyinput_f112), .A(n10018), .ZN(n10021) );
  AOI22_X1 U11186 ( .A1(SI_23_), .A2(keyinput_f9), .B1(P1_IR_REG_23__SCAN_IN), 
        .B2(keyinput_f114), .ZN(n10019) );
  OAI221_X1 U11187 ( .B1(SI_23_), .B2(keyinput_f9), .C1(P1_IR_REG_23__SCAN_IN), 
        .C2(keyinput_f114), .A(n10019), .ZN(n10020) );
  NOR4_X1 U11188 ( .A1(n10023), .A2(n10022), .A3(n10021), .A4(n10020), .ZN(
        n10051) );
  AOI22_X1 U11189 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(keyinput_f41), .B1(
        P1_IR_REG_16__SCAN_IN), .B2(keyinput_f107), .ZN(n10024) );
  OAI221_X1 U11190 ( .B1(P2_REG3_REG_19__SCAN_IN), .B2(keyinput_f41), .C1(
        P1_IR_REG_16__SCAN_IN), .C2(keyinput_f107), .A(n10024), .ZN(n10031) );
  AOI22_X1 U11191 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(keyinput_f52), .B1(
        P2_REG3_REG_6__SCAN_IN), .B2(keyinput_f61), .ZN(n10025) );
  OAI221_X1 U11192 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(keyinput_f52), .C1(
        P2_REG3_REG_6__SCAN_IN), .C2(keyinput_f61), .A(n10025), .ZN(n10030) );
  AOI22_X1 U11193 ( .A1(SI_17_), .A2(keyinput_f15), .B1(P1_IR_REG_19__SCAN_IN), 
        .B2(keyinput_f110), .ZN(n10026) );
  OAI221_X1 U11194 ( .B1(SI_17_), .B2(keyinput_f15), .C1(P1_IR_REG_19__SCAN_IN), .C2(keyinput_f110), .A(n10026), .ZN(n10029) );
  AOI22_X1 U11195 ( .A1(SI_24_), .A2(keyinput_f8), .B1(P1_D_REG_2__SCAN_IN), 
        .B2(keyinput_f125), .ZN(n10027) );
  OAI221_X1 U11196 ( .B1(SI_24_), .B2(keyinput_f8), .C1(P1_D_REG_2__SCAN_IN), 
        .C2(keyinput_f125), .A(n10027), .ZN(n10028) );
  NOR4_X1 U11197 ( .A1(n10031), .A2(n10030), .A3(n10029), .A4(n10028), .ZN(
        n10050) );
  AOI22_X1 U11198 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(keyinput_f118), .B1(
        P1_IR_REG_24__SCAN_IN), .B2(keyinput_f115), .ZN(n10032) );
  OAI221_X1 U11199 ( .B1(P1_IR_REG_27__SCAN_IN), .B2(keyinput_f118), .C1(
        P1_IR_REG_24__SCAN_IN), .C2(keyinput_f115), .A(n10032), .ZN(n10039) );
  AOI22_X1 U11200 ( .A1(SI_7_), .A2(keyinput_f25), .B1(P1_IR_REG_3__SCAN_IN), 
        .B2(keyinput_f94), .ZN(n10033) );
  OAI221_X1 U11201 ( .B1(SI_7_), .B2(keyinput_f25), .C1(P1_IR_REG_3__SCAN_IN), 
        .C2(keyinput_f94), .A(n10033), .ZN(n10038) );
  AOI22_X1 U11202 ( .A1(SI_21_), .A2(keyinput_f11), .B1(P1_IR_REG_0__SCAN_IN), 
        .B2(keyinput_f91), .ZN(n10034) );
  OAI221_X1 U11203 ( .B1(SI_21_), .B2(keyinput_f11), .C1(P1_IR_REG_0__SCAN_IN), 
        .C2(keyinput_f91), .A(n10034), .ZN(n10037) );
  AOI22_X1 U11204 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(keyinput_f60), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(keyinput_f90), .ZN(n10035) );
  OAI221_X1 U11205 ( .B1(P2_REG3_REG_18__SCAN_IN), .B2(keyinput_f60), .C1(
        P2_DATAO_REG_6__SCAN_IN), .C2(keyinput_f90), .A(n10035), .ZN(n10036)
         );
  NOR4_X1 U11206 ( .A1(n10039), .A2(n10038), .A3(n10037), .A4(n10036), .ZN(
        n10049) );
  AOI22_X1 U11207 ( .A1(P2_DATAO_REG_8__SCAN_IN), .A2(keyinput_f88), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(keyinput_f72), .ZN(n10040) );
  OAI221_X1 U11208 ( .B1(P2_DATAO_REG_8__SCAN_IN), .B2(keyinput_f88), .C1(
        P2_DATAO_REG_24__SCAN_IN), .C2(keyinput_f72), .A(n10040), .ZN(n10047)
         );
  AOI22_X1 U11209 ( .A1(P2_DATAO_REG_11__SCAN_IN), .A2(keyinput_f85), .B1(
        P1_IR_REG_28__SCAN_IN), .B2(keyinput_f119), .ZN(n10041) );
  OAI221_X1 U11210 ( .B1(P2_DATAO_REG_11__SCAN_IN), .B2(keyinput_f85), .C1(
        P1_IR_REG_28__SCAN_IN), .C2(keyinput_f119), .A(n10041), .ZN(n10046) );
  AOI22_X1 U11211 ( .A1(P2_DATAO_REG_7__SCAN_IN), .A2(keyinput_f89), .B1(
        P1_IR_REG_11__SCAN_IN), .B2(keyinput_f102), .ZN(n10042) );
  OAI221_X1 U11212 ( .B1(P2_DATAO_REG_7__SCAN_IN), .B2(keyinput_f89), .C1(
        P1_IR_REG_11__SCAN_IN), .C2(keyinput_f102), .A(n10042), .ZN(n10045) );
  AOI22_X1 U11213 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(keyinput_f40), .B1(
        P2_REG3_REG_14__SCAN_IN), .B2(keyinput_f37), .ZN(n10043) );
  OAI221_X1 U11214 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(keyinput_f40), .C1(
        P2_REG3_REG_14__SCAN_IN), .C2(keyinput_f37), .A(n10043), .ZN(n10044)
         );
  NOR4_X1 U11215 ( .A1(n10047), .A2(n10046), .A3(n10045), .A4(n10044), .ZN(
        n10048) );
  NAND4_X1 U11216 ( .A1(n10051), .A2(n10050), .A3(n10049), .A4(n10048), .ZN(
        n10164) );
  AOI22_X1 U11217 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(keyinput_f46), .B1(SI_1_), .B2(keyinput_f31), .ZN(n10052) );
  OAI221_X1 U11218 ( .B1(P2_REG3_REG_12__SCAN_IN), .B2(keyinput_f46), .C1(
        SI_1_), .C2(keyinput_f31), .A(n10052), .ZN(n10060) );
  AOI22_X1 U11219 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(keyinput_f43), .B1(
        P1_IR_REG_25__SCAN_IN), .B2(keyinput_f116), .ZN(n10053) );
  OAI221_X1 U11220 ( .B1(P2_REG3_REG_8__SCAN_IN), .B2(keyinput_f43), .C1(
        P1_IR_REG_25__SCAN_IN), .C2(keyinput_f116), .A(n10053), .ZN(n10059) );
  AOI22_X1 U11221 ( .A1(SI_4_), .A2(keyinput_f28), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(keyinput_f80), .ZN(n10054) );
  OAI221_X1 U11222 ( .B1(SI_4_), .B2(keyinput_f28), .C1(
        P2_DATAO_REG_16__SCAN_IN), .C2(keyinput_f80), .A(n10054), .ZN(n10058)
         );
  XNOR2_X1 U11223 ( .A(P1_IR_REG_15__SCAN_IN), .B(keyinput_f106), .ZN(n10056)
         );
  XNOR2_X1 U11224 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(keyinput_f79), .ZN(n10055) );
  NAND2_X1 U11225 ( .A1(n10056), .A2(n10055), .ZN(n10057) );
  NOR4_X1 U11226 ( .A1(n10060), .A2(n10059), .A3(n10058), .A4(n10057), .ZN(
        n10105) );
  AOI22_X1 U11227 ( .A1(n10063), .A2(keyinput_f86), .B1(keyinput_f39), .B2(
        n10062), .ZN(n10061) );
  OAI221_X1 U11228 ( .B1(n10063), .B2(keyinput_f86), .C1(n10062), .C2(
        keyinput_f39), .A(n10061), .ZN(n10075) );
  AOI22_X1 U11229 ( .A1(n10066), .A2(keyinput_f58), .B1(n10065), .B2(
        keyinput_f75), .ZN(n10064) );
  OAI221_X1 U11230 ( .B1(n10066), .B2(keyinput_f58), .C1(n10065), .C2(
        keyinput_f75), .A(n10064), .ZN(n10074) );
  AOI22_X1 U11231 ( .A1(n10069), .A2(keyinput_f38), .B1(n10068), .B2(
        keyinput_f18), .ZN(n10067) );
  OAI221_X1 U11232 ( .B1(n10069), .B2(keyinput_f38), .C1(n10068), .C2(
        keyinput_f18), .A(n10067), .ZN(n10073) );
  XNOR2_X1 U11233 ( .A(P1_IR_REG_8__SCAN_IN), .B(keyinput_f99), .ZN(n10071) );
  XNOR2_X1 U11234 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput_f96), .ZN(n10070) );
  NAND2_X1 U11235 ( .A1(n10071), .A2(n10070), .ZN(n10072) );
  NOR4_X1 U11236 ( .A1(n10075), .A2(n10074), .A3(n10073), .A4(n10072), .ZN(
        n10104) );
  AOI22_X1 U11237 ( .A1(n10077), .A2(keyinput_f76), .B1(keyinput_f53), .B2(
        n5368), .ZN(n10076) );
  OAI221_X1 U11238 ( .B1(n10077), .B2(keyinput_f76), .C1(n5368), .C2(
        keyinput_f53), .A(n10076), .ZN(n10089) );
  AOI22_X1 U11239 ( .A1(n10080), .A2(keyinput_f22), .B1(keyinput_f67), .B2(
        n10079), .ZN(n10078) );
  OAI221_X1 U11240 ( .B1(n10080), .B2(keyinput_f22), .C1(n10079), .C2(
        keyinput_f67), .A(n10078), .ZN(n10088) );
  AOI22_X1 U11241 ( .A1(n10083), .A2(keyinput_f13), .B1(keyinput_f26), .B2(
        n10082), .ZN(n10081) );
  OAI221_X1 U11242 ( .B1(n10083), .B2(keyinput_f13), .C1(n10082), .C2(
        keyinput_f26), .A(n10081), .ZN(n10087) );
  XNOR2_X1 U11243 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput_f111), .ZN(n10085)
         );
  XNOR2_X1 U11244 ( .A(P2_B_REG_SCAN_IN), .B(keyinput_f64), .ZN(n10084) );
  NAND2_X1 U11245 ( .A1(n10085), .A2(n10084), .ZN(n10086) );
  NOR4_X1 U11246 ( .A1(n10089), .A2(n10088), .A3(n10087), .A4(n10086), .ZN(
        n10103) );
  AOI22_X1 U11247 ( .A1(n10092), .A2(keyinput_f49), .B1(n10091), .B2(
        keyinput_f7), .ZN(n10090) );
  OAI221_X1 U11248 ( .B1(n10092), .B2(keyinput_f49), .C1(n10091), .C2(
        keyinput_f7), .A(n10090), .ZN(n10101) );
  XNOR2_X1 U11249 ( .A(P1_IR_REG_2__SCAN_IN), .B(keyinput_f93), .ZN(n10096) );
  XNOR2_X1 U11250 ( .A(P2_STATE_REG_SCAN_IN), .B(keyinput_f34), .ZN(n10095) );
  XNOR2_X1 U11251 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(keyinput_f74), .ZN(n10094) );
  XNOR2_X1 U11252 ( .A(SI_0_), .B(keyinput_f32), .ZN(n10093) );
  NAND4_X1 U11253 ( .A1(n10096), .A2(n10095), .A3(n10094), .A4(n10093), .ZN(
        n10100) );
  XNOR2_X1 U11254 ( .A(n10097), .B(keyinput_f105), .ZN(n10099) );
  XNOR2_X1 U11255 ( .A(keyinput_f4), .B(n7588), .ZN(n10098) );
  NOR4_X1 U11256 ( .A1(n10101), .A2(n10100), .A3(n10099), .A4(n10098), .ZN(
        n10102) );
  NAND4_X1 U11257 ( .A1(n10105), .A2(n10104), .A3(n10103), .A4(n10102), .ZN(
        n10163) );
  AOI22_X1 U11258 ( .A1(n10108), .A2(keyinput_f109), .B1(keyinput_f123), .B2(
        n10107), .ZN(n10106) );
  OAI221_X1 U11259 ( .B1(n10108), .B2(keyinput_f109), .C1(n10107), .C2(
        keyinput_f123), .A(n10106), .ZN(n10118) );
  XNOR2_X1 U11260 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput_f122), .ZN(n10112)
         );
  XNOR2_X1 U11261 ( .A(P2_REG3_REG_21__SCAN_IN), .B(keyinput_f45), .ZN(n10111)
         );
  XNOR2_X1 U11262 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(keyinput_f87), .ZN(n10110)
         );
  XNOR2_X1 U11263 ( .A(SI_3_), .B(keyinput_f29), .ZN(n10109) );
  NAND4_X1 U11264 ( .A1(n10112), .A2(n10111), .A3(n10110), .A4(n10109), .ZN(
        n10117) );
  XNOR2_X1 U11265 ( .A(n10113), .B(keyinput_f92), .ZN(n10116) );
  INV_X1 U11266 ( .A(SI_15_), .ZN(n10114) );
  XNOR2_X1 U11267 ( .A(keyinput_f17), .B(n10114), .ZN(n10115) );
  NOR4_X1 U11268 ( .A1(n10118), .A2(n10117), .A3(n10116), .A4(n10115), .ZN(
        n10161) );
  AOI22_X1 U11269 ( .A1(n10121), .A2(keyinput_f82), .B1(keyinput_f68), .B2(
        n10120), .ZN(n10119) );
  OAI221_X1 U11270 ( .B1(n10121), .B2(keyinput_f82), .C1(n10120), .C2(
        keyinput_f68), .A(n10119), .ZN(n10131) );
  AOI22_X1 U11271 ( .A1(n10124), .A2(keyinput_f6), .B1(n10123), .B2(
        keyinput_f104), .ZN(n10122) );
  OAI221_X1 U11272 ( .B1(n10124), .B2(keyinput_f6), .C1(n10123), .C2(
        keyinput_f104), .A(n10122), .ZN(n10130) );
  XNOR2_X1 U11273 ( .A(SI_9_), .B(keyinput_f23), .ZN(n10128) );
  XNOR2_X1 U11274 ( .A(SI_2_), .B(keyinput_f30), .ZN(n10127) );
  XNOR2_X1 U11275 ( .A(P1_IR_REG_10__SCAN_IN), .B(keyinput_f101), .ZN(n10126)
         );
  XNOR2_X1 U11276 ( .A(P2_REG3_REG_20__SCAN_IN), .B(keyinput_f55), .ZN(n10125)
         );
  NAND4_X1 U11277 ( .A1(n10128), .A2(n10127), .A3(n10126), .A4(n10125), .ZN(
        n10129) );
  NOR3_X1 U11278 ( .A1(n10131), .A2(n10130), .A3(n10129), .ZN(n10160) );
  AOI22_X1 U11279 ( .A1(n8104), .A2(keyinput_f47), .B1(n10133), .B2(
        keyinput_f16), .ZN(n10132) );
  OAI221_X1 U11280 ( .B1(n8104), .B2(keyinput_f47), .C1(n10133), .C2(
        keyinput_f16), .A(n10132), .ZN(n10142) );
  AOI22_X1 U11281 ( .A1(n6775), .A2(keyinput_f59), .B1(n10135), .B2(
        keyinput_f12), .ZN(n10134) );
  OAI221_X1 U11282 ( .B1(n6775), .B2(keyinput_f59), .C1(n10135), .C2(
        keyinput_f12), .A(n10134), .ZN(n10141) );
  XNOR2_X1 U11283 ( .A(SI_5_), .B(keyinput_f27), .ZN(n10139) );
  XNOR2_X1 U11284 ( .A(P1_IR_REG_30__SCAN_IN), .B(keyinput_f121), .ZN(n10138)
         );
  XNOR2_X1 U11285 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput_f98), .ZN(n10137) );
  XNOR2_X1 U11286 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(keyinput_f73), .ZN(n10136) );
  NAND4_X1 U11287 ( .A1(n10139), .A2(n10138), .A3(n10137), .A4(n10136), .ZN(
        n10140) );
  NOR3_X1 U11288 ( .A1(n10142), .A2(n10141), .A3(n10140), .ZN(n10159) );
  AOI22_X1 U11289 ( .A1(n10145), .A2(keyinput_f97), .B1(keyinput_f51), .B2(
        n10144), .ZN(n10143) );
  OAI221_X1 U11290 ( .B1(n10145), .B2(keyinput_f97), .C1(n10144), .C2(
        keyinput_f51), .A(n10143), .ZN(n10157) );
  AOI22_X1 U11291 ( .A1(n10148), .A2(keyinput_f54), .B1(n10147), .B2(
        keyinput_f24), .ZN(n10146) );
  OAI221_X1 U11292 ( .B1(n10148), .B2(keyinput_f54), .C1(n10147), .C2(
        keyinput_f24), .A(n10146), .ZN(n10156) );
  AOI22_X1 U11293 ( .A1(n10151), .A2(keyinput_f62), .B1(n10150), .B2(
        keyinput_f20), .ZN(n10149) );
  OAI221_X1 U11294 ( .B1(n10151), .B2(keyinput_f62), .C1(n10150), .C2(
        keyinput_f20), .A(n10149), .ZN(n10155) );
  XNOR2_X1 U11295 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(keyinput_f78), .ZN(n10153) );
  XNOR2_X1 U11296 ( .A(P2_RD_REG_SCAN_IN), .B(keyinput_f33), .ZN(n10152) );
  NAND2_X1 U11297 ( .A1(n10153), .A2(n10152), .ZN(n10154) );
  NOR4_X1 U11298 ( .A1(n10157), .A2(n10156), .A3(n10155), .A4(n10154), .ZN(
        n10158) );
  NAND4_X1 U11299 ( .A1(n10161), .A2(n10160), .A3(n10159), .A4(n10158), .ZN(
        n10162) );
  OR4_X1 U11300 ( .A1(n10165), .A2(n10164), .A3(n10163), .A4(n10162), .ZN(
        n10167) );
  AOI21_X1 U11301 ( .B1(keyinput_f81), .B2(n10167), .A(keyinput_g81), .ZN(
        n10169) );
  INV_X1 U11302 ( .A(keyinput_f81), .ZN(n10166) );
  AOI21_X1 U11303 ( .B1(n10167), .B2(n10166), .A(P2_DATAO_REG_15__SCAN_IN), 
        .ZN(n10168) );
  AOI22_X1 U11304 ( .A1(P2_DATAO_REG_15__SCAN_IN), .A2(n10169), .B1(
        keyinput_g81), .B2(n10168), .ZN(n10170) );
  AOI21_X1 U11305 ( .B1(n10172), .B2(n10171), .A(n10170), .ZN(n10173) );
  XNOR2_X1 U11306 ( .A(n10174), .B(n10173), .ZN(n10178) );
  NOR2_X1 U11307 ( .A1(n10176), .A2(n10175), .ZN(n10177) );
  XOR2_X1 U11308 ( .A(n10178), .B(n10177), .Z(ADD_1071_U4) );
  INV_X1 U11309 ( .A(n10179), .ZN(n10184) );
  OAI21_X1 U11310 ( .B1(n10181), .B2(n10386), .A(n10180), .ZN(n10183) );
  AOI211_X1 U11311 ( .C1(n10393), .C2(n10184), .A(n10183), .B(n10182), .ZN(
        n10186) );
  INV_X1 U11312 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n10185) );
  AOI22_X1 U11313 ( .A1(n10396), .A2(n10186), .B1(n10185), .B2(n10394), .ZN(
        P1_U3484) );
  AOI22_X1 U11314 ( .A1(n4483), .A2(n10186), .B1(n5978), .B2(n10399), .ZN(
        P1_U3533) );
  AOI22_X1 U11315 ( .A1(n10188), .A2(n10187), .B1(P2_REG3_REG_15__SCAN_IN), 
        .B2(P2_U3152), .ZN(n10197) );
  XNOR2_X1 U11316 ( .A(n10189), .B(n10190), .ZN(n10195) );
  INV_X1 U11317 ( .A(n10191), .ZN(n10193) );
  AOI22_X1 U11318 ( .A1(n10195), .A2(n10194), .B1(n10193), .B2(n10192), .ZN(
        n10196) );
  OAI211_X1 U11319 ( .C1(n10199), .C2(n10198), .A(n10197), .B(n10196), .ZN(
        P2_U3243) );
  NAND2_X1 U11320 ( .A1(n10201), .A2(n10200), .ZN(n10202) );
  NAND2_X1 U11321 ( .A1(n10203), .A2(n10202), .ZN(n10231) );
  AOI21_X1 U11322 ( .B1(n10204), .B2(n10227), .A(n10472), .ZN(n10205) );
  NAND2_X1 U11323 ( .A1(n10205), .A2(n4496), .ZN(n10232) );
  OAI22_X1 U11324 ( .A1(n10231), .A2(n10417), .B1(n10206), .B2(n10232), .ZN(
        n10207) );
  INV_X1 U11325 ( .A(n10207), .ZN(n10230) );
  OAI22_X1 U11326 ( .A1(n10211), .A2(n10210), .B1(n10209), .B2(n10208), .ZN(
        n10226) );
  OR2_X1 U11327 ( .A1(n10231), .A2(n10435), .ZN(n10224) );
  NAND2_X1 U11328 ( .A1(n10213), .A2(n10212), .ZN(n10214) );
  NAND2_X1 U11329 ( .A1(n10215), .A2(n10214), .ZN(n10222) );
  NAND2_X1 U11330 ( .A1(n10217), .A2(n10216), .ZN(n10220) );
  NAND2_X1 U11331 ( .A1(n10218), .A2(n8701), .ZN(n10219) );
  NAND2_X1 U11332 ( .A1(n10220), .A2(n10219), .ZN(n10221) );
  AOI21_X1 U11333 ( .B1(n10222), .B2(n10432), .A(n10221), .ZN(n10223) );
  NOR2_X1 U11334 ( .A1(n10237), .A2(n10456), .ZN(n10225) );
  AOI211_X1 U11335 ( .C1(n10228), .C2(n10227), .A(n10226), .B(n10225), .ZN(
        n10229) );
  NAND2_X1 U11336 ( .A1(n10230), .A2(n10229), .ZN(P2_U3283) );
  INV_X1 U11337 ( .A(n10231), .ZN(n10235) );
  OAI21_X1 U11338 ( .B1(n10233), .B2(n10488), .A(n10232), .ZN(n10234) );
  AOI21_X1 U11339 ( .B1(n10235), .B2(n10493), .A(n10234), .ZN(n10236) );
  AOI22_X1 U11340 ( .A1(n10499), .A2(n10240), .B1(n10238), .B2(n10504), .ZN(
        P2_U3533) );
  INV_X1 U11341 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n10239) );
  AOI22_X1 U11342 ( .A1(n10496), .A2(n10240), .B1(n10239), .B2(n10494), .ZN(
        P2_U3490) );
  XNOR2_X1 U11343 ( .A(n10241), .B(n10247), .ZN(n10257) );
  INV_X1 U11344 ( .A(n10257), .ZN(n10274) );
  INV_X1 U11345 ( .A(n10242), .ZN(n10244) );
  OAI21_X1 U11346 ( .B1(n10244), .B2(n10269), .A(n10243), .ZN(n10270) );
  INV_X1 U11347 ( .A(n10270), .ZN(n10245) );
  AOI22_X1 U11348 ( .A1(n10274), .A2(n10344), .B1(n10343), .B2(n10245), .ZN(
        n10263) );
  INV_X1 U11349 ( .A(n10246), .ZN(n10251) );
  NAND3_X1 U11350 ( .A1(n10249), .A2(n10248), .A3(n10247), .ZN(n10250) );
  NAND2_X1 U11351 ( .A1(n10251), .A2(n10250), .ZN(n10256) );
  AOI222_X1 U11352 ( .A1(n10355), .A2(n10256), .B1(n10255), .B2(n10254), .C1(
        n10253), .C2(n10252), .ZN(n10271) );
  OAI21_X1 U11353 ( .B1(n10358), .B2(n10257), .A(n10271), .ZN(n10261) );
  AOI22_X1 U11354 ( .A1(n10362), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n10258), 
        .B2(n10360), .ZN(n10259) );
  OAI21_X1 U11355 ( .B1(n10269), .B2(n10364), .A(n10259), .ZN(n10260) );
  AOI21_X1 U11356 ( .B1(n10261), .B2(n10366), .A(n10260), .ZN(n10262) );
  NAND2_X1 U11357 ( .A1(n10263), .A2(n10262), .ZN(P1_U3278) );
  NOR2_X1 U11358 ( .A1(n10264), .A2(n10388), .ZN(n10265) );
  INV_X1 U11359 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n10268) );
  AOI22_X1 U11360 ( .A1(n4483), .A2(n10288), .B1(n10268), .B2(n10399), .ZN(
        P1_U3553) );
  OAI22_X1 U11361 ( .A1(n10270), .A2(n10388), .B1(n10269), .B2(n10386), .ZN(
        n10273) );
  INV_X1 U11362 ( .A(n10271), .ZN(n10272) );
  AOI211_X1 U11363 ( .C1(n10274), .C2(n10279), .A(n10273), .B(n10272), .ZN(
        n10290) );
  AOI22_X1 U11364 ( .A1(n4483), .A2(n10290), .B1(n6450), .B2(n10399), .ZN(
        P1_U3536) );
  OAI211_X1 U11365 ( .C1(n10277), .C2(n10386), .A(n10276), .B(n10275), .ZN(
        n10278) );
  AOI21_X1 U11366 ( .B1(n10280), .B2(n10279), .A(n10278), .ZN(n10292) );
  AOI22_X1 U11367 ( .A1(n4483), .A2(n10292), .B1(n6235), .B2(n10399), .ZN(
        P1_U3535) );
  OAI22_X1 U11368 ( .A1(n10282), .A2(n10388), .B1(n10281), .B2(n10386), .ZN(
        n10284) );
  AOI211_X1 U11369 ( .C1(n10393), .C2(n10285), .A(n10284), .B(n10283), .ZN(
        n10294) );
  AOI22_X1 U11370 ( .A1(n4483), .A2(n10294), .B1(n10286), .B2(n10399), .ZN(
        P1_U3534) );
  INV_X1 U11371 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n10287) );
  AOI22_X1 U11372 ( .A1(n10396), .A2(n10288), .B1(n10287), .B2(n10394), .ZN(
        P1_U3521) );
  INV_X1 U11373 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n10289) );
  AOI22_X1 U11374 ( .A1(n10396), .A2(n10290), .B1(n10289), .B2(n10394), .ZN(
        P1_U3493) );
  INV_X1 U11375 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n10291) );
  AOI22_X1 U11376 ( .A1(n10396), .A2(n10292), .B1(n10291), .B2(n10394), .ZN(
        P1_U3490) );
  INV_X1 U11377 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n10293) );
  AOI22_X1 U11378 ( .A1(n10396), .A2(n10294), .B1(n10293), .B2(n10394), .ZN(
        P1_U3487) );
  XNOR2_X1 U11379 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  OAI21_X1 U11380 ( .B1(n10297), .B2(n10296), .A(n10295), .ZN(n10298) );
  AOI22_X1 U11381 ( .A1(n10299), .A2(P1_ADDR_REG_8__SCAN_IN), .B1(n10331), 
        .B2(n10298), .ZN(n10307) );
  AND3_X1 U11382 ( .A1(n10332), .A2(P1_REG1_REG_8__SCAN_IN), .A3(n10303), .ZN(
        n10301) );
  OAI21_X1 U11383 ( .B1(n10301), .B2(n10324), .A(n10300), .ZN(n10305) );
  OAI211_X1 U11384 ( .C1(n10303), .C2(n10302), .A(n10332), .B(n10318), .ZN(
        n10304) );
  NAND4_X1 U11385 ( .A1(n10307), .A2(n10306), .A3(n10305), .A4(n10304), .ZN(
        P1_U3249) );
  AOI21_X1 U11386 ( .B1(n10324), .B2(n10309), .A(n10308), .ZN(n10315) );
  AOI21_X1 U11387 ( .B1(n10312), .B2(n10311), .A(n10310), .ZN(n10313) );
  NAND2_X1 U11388 ( .A1(n10331), .A2(n10313), .ZN(n10314) );
  AND2_X1 U11389 ( .A1(n10315), .A2(n10314), .ZN(n10321) );
  OAI21_X1 U11390 ( .B1(n10318), .B2(n10317), .A(n10316), .ZN(n10319) );
  NAND2_X1 U11391 ( .A1(n10319), .A2(n10332), .ZN(n10320) );
  OAI211_X1 U11392 ( .C1(n10537), .C2(n10337), .A(n10321), .B(n10320), .ZN(
        P1_U3250) );
  INV_X1 U11393 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n10336) );
  AOI21_X1 U11394 ( .B1(n10324), .B2(n10323), .A(n10322), .ZN(n10335) );
  OAI21_X1 U11395 ( .B1(n10327), .B2(n10326), .A(n10325), .ZN(n10333) );
  OAI21_X1 U11396 ( .B1(n4560), .B2(n10329), .A(n10328), .ZN(n10330) );
  AOI22_X1 U11397 ( .A1(n10333), .A2(n10332), .B1(n10331), .B2(n10330), .ZN(
        n10334) );
  OAI211_X1 U11398 ( .C1(n10337), .C2(n10336), .A(n10335), .B(n10334), .ZN(
        P1_U3252) );
  XOR2_X1 U11399 ( .A(n10348), .B(n10338), .Z(n10359) );
  INV_X1 U11400 ( .A(n10359), .ZN(n10392) );
  INV_X1 U11401 ( .A(n10339), .ZN(n10341) );
  OAI21_X1 U11402 ( .B1(n10341), .B2(n10387), .A(n10340), .ZN(n10389) );
  INV_X1 U11403 ( .A(n10389), .ZN(n10342) );
  AOI22_X1 U11404 ( .A1(n10392), .A2(n10344), .B1(n10343), .B2(n10342), .ZN(
        n10368) );
  INV_X1 U11405 ( .A(n10345), .ZN(n10346) );
  NOR2_X1 U11406 ( .A1(n10347), .A2(n10346), .ZN(n10349) );
  XNOR2_X1 U11407 ( .A(n10349), .B(n10348), .ZN(n10356) );
  OAI22_X1 U11408 ( .A1(n10353), .A2(n10352), .B1(n10351), .B2(n10350), .ZN(
        n10354) );
  AOI21_X1 U11409 ( .B1(n10356), .B2(n10355), .A(n10354), .ZN(n10357) );
  OAI21_X1 U11410 ( .B1(n10359), .B2(n10358), .A(n10357), .ZN(n10390) );
  AOI22_X1 U11411 ( .A1(n10362), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n10361), 
        .B2(n10360), .ZN(n10363) );
  OAI21_X1 U11412 ( .B1(n10364), .B2(n10387), .A(n10363), .ZN(n10365) );
  AOI21_X1 U11413 ( .B1(n10390), .B2(n10366), .A(n10365), .ZN(n10367) );
  NAND2_X1 U11414 ( .A1(n10368), .A2(n10367), .ZN(P1_U3282) );
  AND2_X1 U11415 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n10371), .ZN(P1_U3292) );
  AND2_X1 U11416 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n10371), .ZN(P1_U3293) );
  AND2_X1 U11417 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n10371), .ZN(P1_U3294) );
  AND2_X1 U11418 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n10371), .ZN(P1_U3295) );
  AND2_X1 U11419 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n10371), .ZN(P1_U3296) );
  AND2_X1 U11420 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n10371), .ZN(P1_U3297) );
  AND2_X1 U11421 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n10371), .ZN(P1_U3298) );
  AND2_X1 U11422 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n10371), .ZN(P1_U3299) );
  AND2_X1 U11423 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n10371), .ZN(P1_U3300) );
  AND2_X1 U11424 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n10371), .ZN(P1_U3301) );
  AND2_X1 U11425 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n10371), .ZN(P1_U3302) );
  AND2_X1 U11426 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n10371), .ZN(P1_U3303) );
  AND2_X1 U11427 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n10371), .ZN(P1_U3304) );
  AND2_X1 U11428 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n10371), .ZN(P1_U3305) );
  AND2_X1 U11429 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n10371), .ZN(P1_U3306) );
  AND2_X1 U11430 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n10371), .ZN(P1_U3307) );
  AND2_X1 U11431 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n10371), .ZN(P1_U3308) );
  AND2_X1 U11432 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n10371), .ZN(P1_U3309) );
  AND2_X1 U11433 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n10371), .ZN(P1_U3310) );
  AND2_X1 U11434 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n10371), .ZN(P1_U3311) );
  AND2_X1 U11435 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n10371), .ZN(P1_U3312) );
  AND2_X1 U11436 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n10371), .ZN(P1_U3313) );
  AND2_X1 U11437 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n10371), .ZN(P1_U3314) );
  AND2_X1 U11438 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n10371), .ZN(P1_U3315) );
  AND2_X1 U11439 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n10371), .ZN(P1_U3316) );
  AND2_X1 U11440 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n10371), .ZN(P1_U3317) );
  AND2_X1 U11441 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n10371), .ZN(P1_U3318) );
  AND2_X1 U11442 ( .A1(n10371), .A2(P1_D_REG_4__SCAN_IN), .ZN(P1_U3319) );
  NOR2_X1 U11443 ( .A1(n10370), .A2(n10369), .ZN(P1_U3320) );
  AND2_X1 U11444 ( .A1(n10371), .A2(P1_D_REG_2__SCAN_IN), .ZN(P1_U3321) );
  NAND2_X1 U11445 ( .A1(n10372), .A2(n6310), .ZN(n10373) );
  OAI211_X1 U11446 ( .C1(n10376), .C2(n10375), .A(n10374), .B(n10373), .ZN(
        n10377) );
  NOR2_X1 U11447 ( .A1(n10378), .A2(n10377), .ZN(n10397) );
  INV_X1 U11448 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n10379) );
  AOI22_X1 U11449 ( .A1(n10396), .A2(n10397), .B1(n10379), .B2(n10394), .ZN(
        P1_U3457) );
  OAI22_X1 U11450 ( .A1(n10381), .A2(n10388), .B1(n10380), .B2(n10386), .ZN(
        n10383) );
  AOI211_X1 U11451 ( .C1(n10393), .C2(n10384), .A(n10383), .B(n10382), .ZN(
        n10398) );
  INV_X1 U11452 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n10385) );
  AOI22_X1 U11453 ( .A1(n10396), .A2(n10398), .B1(n10385), .B2(n10394), .ZN(
        P1_U3463) );
  OAI22_X1 U11454 ( .A1(n10389), .A2(n10388), .B1(n10387), .B2(n10386), .ZN(
        n10391) );
  AOI211_X1 U11455 ( .C1(n10393), .C2(n10392), .A(n10391), .B(n10390), .ZN(
        n10401) );
  INV_X1 U11456 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n10395) );
  AOI22_X1 U11457 ( .A1(n10396), .A2(n10401), .B1(n10395), .B2(n10394), .ZN(
        P1_U3481) );
  AOI22_X1 U11458 ( .A1(n4483), .A2(n10397), .B1(n5952), .B2(n10399), .ZN(
        P1_U3524) );
  AOI22_X1 U11459 ( .A1(n4483), .A2(n10398), .B1(n5958), .B2(n10399), .ZN(
        P1_U3526) );
  INV_X1 U11460 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10400) );
  AOI22_X1 U11461 ( .A1(n4483), .A2(n10401), .B1(n10400), .B2(n10399), .ZN(
        P1_U3532) );
  AOI22_X1 U11462 ( .A1(n10403), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n10402), .ZN(n10412) );
  AOI22_X1 U11463 ( .A1(n10404), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n10411) );
  NOR2_X1 U11464 ( .A1(n10405), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n10409) );
  OAI21_X1 U11465 ( .B1(P2_REG1_REG_0__SCAN_IN), .B2(n10407), .A(n10406), .ZN(
        n10408) );
  OAI21_X1 U11466 ( .B1(n10409), .B2(n10408), .A(n10413), .ZN(n10410) );
  OAI211_X1 U11467 ( .C1(n10413), .C2(n10412), .A(n10411), .B(n10410), .ZN(
        P2_U3245) );
  INV_X1 U11468 ( .A(n10414), .ZN(n10415) );
  AOI21_X1 U11469 ( .B1(n10426), .B2(n10416), .A(n10415), .ZN(n10436) );
  INV_X1 U11470 ( .A(n10436), .ZN(n10492) );
  INV_X1 U11471 ( .A(n10417), .ZN(n10423) );
  OAI211_X1 U11472 ( .C1(n10420), .C2(n10489), .A(n10419), .B(n10418), .ZN(
        n10487) );
  INV_X1 U11473 ( .A(n10487), .ZN(n10421) );
  AOI22_X1 U11474 ( .A1(n10492), .A2(n10423), .B1(n10422), .B2(n10421), .ZN(
        n10442) );
  OAI21_X1 U11475 ( .B1(n10426), .B2(n10425), .A(n10424), .ZN(n10433) );
  OAI22_X1 U11476 ( .A1(n10430), .A2(n10429), .B1(n10428), .B2(n10427), .ZN(
        n10431) );
  AOI21_X1 U11477 ( .B1(n10433), .B2(n10432), .A(n10431), .ZN(n10434) );
  OAI21_X1 U11478 ( .B1(n10436), .B2(n10435), .A(n10434), .ZN(n10490) );
  AOI22_X1 U11479 ( .A1(n10456), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n10437), 
        .B2(n10447), .ZN(n10438) );
  OAI21_X1 U11480 ( .B1(n10489), .B2(n10439), .A(n10438), .ZN(n10440) );
  AOI21_X1 U11481 ( .B1(n10490), .B2(n10211), .A(n10440), .ZN(n10441) );
  NAND2_X1 U11482 ( .A1(n10442), .A2(n10441), .ZN(P2_U3287) );
  INV_X1 U11483 ( .A(n10443), .ZN(n10450) );
  AOI22_X1 U11484 ( .A1(n10447), .A2(n10446), .B1(n10445), .B2(n10444), .ZN(
        n10448) );
  OAI21_X1 U11485 ( .B1(n10450), .B2(n10449), .A(n10448), .ZN(n10451) );
  AOI211_X1 U11486 ( .C1(n10454), .C2(n10453), .A(n10452), .B(n10451), .ZN(
        n10455) );
  AOI22_X1 U11487 ( .A1(n10456), .A2(n5860), .B1(n10455), .B2(n10211), .ZN(
        P2_U3291) );
  AND2_X1 U11488 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n10461), .ZN(P2_U3297) );
  AND2_X1 U11489 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n10461), .ZN(P2_U3298) );
  AND2_X1 U11490 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n10461), .ZN(P2_U3299) );
  AND2_X1 U11491 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n10461), .ZN(P2_U3300) );
  AND2_X1 U11492 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n10461), .ZN(P2_U3301) );
  AND2_X1 U11493 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n10461), .ZN(P2_U3302) );
  AND2_X1 U11494 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n10461), .ZN(P2_U3303) );
  AND2_X1 U11495 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n10461), .ZN(P2_U3304) );
  AND2_X1 U11496 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n10461), .ZN(P2_U3305) );
  AND2_X1 U11497 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n10461), .ZN(P2_U3306) );
  AND2_X1 U11498 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n10461), .ZN(P2_U3307) );
  AND2_X1 U11499 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n10461), .ZN(P2_U3308) );
  AND2_X1 U11500 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n10461), .ZN(P2_U3309) );
  AND2_X1 U11501 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n10461), .ZN(P2_U3310) );
  AND2_X1 U11502 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n10461), .ZN(P2_U3311) );
  AND2_X1 U11503 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n10461), .ZN(P2_U3312) );
  AND2_X1 U11504 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n10461), .ZN(P2_U3313) );
  AND2_X1 U11505 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n10461), .ZN(P2_U3314) );
  AND2_X1 U11506 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n10461), .ZN(P2_U3315) );
  AND2_X1 U11507 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n10461), .ZN(P2_U3316) );
  AND2_X1 U11508 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n10461), .ZN(P2_U3317) );
  AND2_X1 U11509 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n10461), .ZN(P2_U3318) );
  AND2_X1 U11510 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n10461), .ZN(P2_U3319) );
  AND2_X1 U11511 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n10461), .ZN(P2_U3320) );
  AND2_X1 U11512 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n10461), .ZN(P2_U3321) );
  AND2_X1 U11513 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n10461), .ZN(P2_U3322) );
  AND2_X1 U11514 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n10461), .ZN(P2_U3323) );
  AND2_X1 U11515 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n10461), .ZN(P2_U3324) );
  AND2_X1 U11516 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n10461), .ZN(P2_U3325) );
  AND2_X1 U11517 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n10461), .ZN(P2_U3326) );
  AOI22_X1 U11518 ( .A1(n10460), .A2(n10463), .B1(n10459), .B2(n10461), .ZN(
        P2_U3437) );
  AOI22_X1 U11519 ( .A1(n10464), .A2(n10463), .B1(n10462), .B2(n10461), .ZN(
        P2_U3438) );
  OAI22_X1 U11520 ( .A1(n10467), .A2(n10466), .B1(n5212), .B2(n10465), .ZN(
        n10468) );
  NOR2_X1 U11521 ( .A1(n10469), .A2(n10468), .ZN(n10498) );
  INV_X1 U11522 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n10470) );
  AOI22_X1 U11523 ( .A1(n10496), .A2(n10498), .B1(n10470), .B2(n10494), .ZN(
        P2_U3451) );
  OAI22_X1 U11524 ( .A1(n10473), .A2(n10472), .B1(n10471), .B2(n10488), .ZN(
        n10476) );
  INV_X1 U11525 ( .A(n10474), .ZN(n10475) );
  AOI211_X1 U11526 ( .C1(n10493), .C2(n10477), .A(n10476), .B(n10475), .ZN(
        n10501) );
  INV_X1 U11527 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10478) );
  AOI22_X1 U11528 ( .A1(n10496), .A2(n10501), .B1(n10478), .B2(n10494), .ZN(
        P2_U3460) );
  OAI21_X1 U11529 ( .B1(n10480), .B2(n10488), .A(n10479), .ZN(n10483) );
  INV_X1 U11530 ( .A(n10481), .ZN(n10482) );
  AOI211_X1 U11531 ( .C1(n10485), .C2(n10484), .A(n10483), .B(n10482), .ZN(
        n10503) );
  INV_X1 U11532 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10486) );
  AOI22_X1 U11533 ( .A1(n10496), .A2(n10503), .B1(n10486), .B2(n10494), .ZN(
        P2_U3472) );
  OAI21_X1 U11534 ( .B1(n10489), .B2(n10488), .A(n10487), .ZN(n10491) );
  AOI211_X1 U11535 ( .C1(n10493), .C2(n10492), .A(n10491), .B(n10490), .ZN(
        n10506) );
  INV_X1 U11536 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10495) );
  AOI22_X1 U11537 ( .A1(n10496), .A2(n10506), .B1(n10495), .B2(n10494), .ZN(
        P2_U3478) );
  INV_X1 U11538 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10497) );
  AOI22_X1 U11539 ( .A1(n10499), .A2(n10498), .B1(n10497), .B2(n10504), .ZN(
        P2_U3520) );
  INV_X1 U11540 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10500) );
  AOI22_X1 U11541 ( .A1(n10499), .A2(n10501), .B1(n10500), .B2(n10504), .ZN(
        P2_U3523) );
  INV_X1 U11542 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n10502) );
  AOI22_X1 U11543 ( .A1(n10499), .A2(n10503), .B1(n10502), .B2(n10504), .ZN(
        P2_U3527) );
  INV_X1 U11544 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n10505) );
  AOI22_X1 U11545 ( .A1(n10499), .A2(n10506), .B1(n10505), .B2(n10504), .ZN(
        P2_U3529) );
  INV_X1 U11546 ( .A(n10507), .ZN(n10508) );
  NAND2_X1 U11547 ( .A1(n10509), .A2(n10508), .ZN(n10510) );
  XOR2_X1 U11548 ( .A(n10511), .B(n10510), .Z(ADD_1071_U5) );
  XOR2_X1 U11549 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  OAI21_X1 U11550 ( .B1(n10514), .B2(n10513), .A(n10512), .ZN(ADD_1071_U56) );
  OAI21_X1 U11551 ( .B1(n10517), .B2(n10516), .A(n10515), .ZN(ADD_1071_U57) );
  OAI21_X1 U11552 ( .B1(n10520), .B2(n10519), .A(n10518), .ZN(ADD_1071_U58) );
  OAI21_X1 U11553 ( .B1(n10523), .B2(n10522), .A(n10521), .ZN(ADD_1071_U59) );
  OAI21_X1 U11554 ( .B1(n10526), .B2(n10525), .A(n10524), .ZN(ADD_1071_U60) );
  OAI21_X1 U11555 ( .B1(n10529), .B2(n10528), .A(n10527), .ZN(ADD_1071_U61) );
  AOI21_X1 U11556 ( .B1(n10532), .B2(n10531), .A(n10530), .ZN(ADD_1071_U62) );
  AOI21_X1 U11557 ( .B1(n10535), .B2(n10534), .A(n10533), .ZN(ADD_1071_U63) );
  AOI21_X1 U11558 ( .B1(n10538), .B2(n10537), .A(n10536), .ZN(ADD_1071_U47) );
  XOR2_X1 U11559 ( .A(n10539), .B(P2_ADDR_REG_7__SCAN_IN), .Z(ADD_1071_U49) );
  XOR2_X1 U11560 ( .A(n10541), .B(n10540), .Z(ADD_1071_U54) );
  NOR2_X1 U11561 ( .A1(n10543), .A2(n10542), .ZN(n10544) );
  XOR2_X1 U11562 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n10544), .Z(ADD_1071_U51) );
  OAI21_X1 U11563 ( .B1(n9381), .B2(n10546), .A(n10545), .ZN(n10547) );
  XNOR2_X1 U11564 ( .A(n10547), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  XOR2_X1 U11565 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n10548), .Z(ADD_1071_U48) );
  XOR2_X1 U11566 ( .A(P2_ADDR_REG_6__SCAN_IN), .B(n10549), .Z(ADD_1071_U50) );
  XOR2_X1 U11567 ( .A(n10551), .B(n10550), .Z(ADD_1071_U53) );
  XNOR2_X1 U11568 ( .A(n10553), .B(n10552), .ZN(ADD_1071_U52) );
  NAND2_X1 U5521 ( .A1(n7651), .A2(n7650), .ZN(n8818) );
  NAND2_X2 U4999 ( .A1(n5215), .A2(n5214), .ZN(n5263) );
  NOR2_X2 U5018 ( .A1(n8589), .A2(n8818), .ZN(n8574) );
  NOR2_X2 U5021 ( .A1(n8627), .A2(n8828), .ZN(n4880) );
  CLKBUF_X1 U5051 ( .A(n4479), .Z(n5387) );
  CLKBUF_X1 U5181 ( .A(n5589), .Z(n4486) );
  CLKBUF_X1 U6153 ( .A(n9515), .Z(n4485) );
  INV_X2 U6224 ( .A(n10456), .ZN(n10211) );
endmodule

