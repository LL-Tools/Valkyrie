

module b14_C_2inp_gates_syn ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, U3352, U3351, U3350, U3349, 
        U3348, U3347, U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, 
        U3338, U3337, U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, 
        U3328, U3327, U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, 
        U3320, U3319, U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, 
        U3310, U3309, U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, 
        U3300, U3299, U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, 
        U3467, U3469, U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, 
        U3487, U3489, U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, 
        U3506, U3507, U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, 
        U3516, U3517, U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, 
        U3526, U3527, U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, 
        U3536, U3537, U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, 
        U3546, U3547, U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, 
        U3284, U3283, U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, 
        U3274, U3273, U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, 
        U3264, U3263, U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, 
        U3255, U3254, U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, 
        U3245, U3244, U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, 
        U3554, U3555, U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, 
        U3564, U3565, U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, 
        U3574, U3575, U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, 
        U3237, U3236, U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, 
        U3227, U3226, U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, 
        U3217, U3216, U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, 
        U4043, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, 
        keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, 
        keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, 
        keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, 
        keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, 
        keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, 
        keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, 
        keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, 
        keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, 
        keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, 
        keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, 
        keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, 
        keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, 
        keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, 
        keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, 
        keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, 
        keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, 
        keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, 
        keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, 
        keyinput110, keyinput111, keyinput112, keyinput113, keyinput114, 
        keyinput115, keyinput116, keyinput117, keyinput118, keyinput119, 
        keyinput120, keyinput121, keyinput122, keyinput123, keyinput124, 
        keyinput125, keyinput126, keyinput127 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2123, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133,
         n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143,
         n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153,
         n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163,
         n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173,
         n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183,
         n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
         n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
         n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
         n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223,
         n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233,
         n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243,
         n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253,
         n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263,
         n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273,
         n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283,
         n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293,
         n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303,
         n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313,
         n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323,
         n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333,
         n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343,
         n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353,
         n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363,
         n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373,
         n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383,
         n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393,
         n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403,
         n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413,
         n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423,
         n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433,
         n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443,
         n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453,
         n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463,
         n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473,
         n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483,
         n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493,
         n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503,
         n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513,
         n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523,
         n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533,
         n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543,
         n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553,
         n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563,
         n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573,
         n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583,
         n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593,
         n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603,
         n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613,
         n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623,
         n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633,
         n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643,
         n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653,
         n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663,
         n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673,
         n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683,
         n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693,
         n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703,
         n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713,
         n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723,
         n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733,
         n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743,
         n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753,
         n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763,
         n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773,
         n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783,
         n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793,
         n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803,
         n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813,
         n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823,
         n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833,
         n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843,
         n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853,
         n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863,
         n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873,
         n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883,
         n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893,
         n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903,
         n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913,
         n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923,
         n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933,
         n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943,
         n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953,
         n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963,
         n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973,
         n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983,
         n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993,
         n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003,
         n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013,
         n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023,
         n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033,
         n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043,
         n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053,
         n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063,
         n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073,
         n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083,
         n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093,
         n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103,
         n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113,
         n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123,
         n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133,
         n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143,
         n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153,
         n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163,
         n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173,
         n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183,
         n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193,
         n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203,
         n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213,
         n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223,
         n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233,
         n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243,
         n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253,
         n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263,
         n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273,
         n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283,
         n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293,
         n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303,
         n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313,
         n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323,
         n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333,
         n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343,
         n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353,
         n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363,
         n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373,
         n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383,
         n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393,
         n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403,
         n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413,
         n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423,
         n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433,
         n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443,
         n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453,
         n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463,
         n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473,
         n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483,
         n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493,
         n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503,
         n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513,
         n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523,
         n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533,
         n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543,
         n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553,
         n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563,
         n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
         n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583,
         n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593,
         n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603,
         n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613,
         n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
         n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633,
         n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
         n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653,
         n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663,
         n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673,
         n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683,
         n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693,
         n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703,
         n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713,
         n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723,
         n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733,
         n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743,
         n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753,
         n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763,
         n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773,
         n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783,
         n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793,
         n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803,
         n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813,
         n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823,
         n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833,
         n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843,
         n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853,
         n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863,
         n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873,
         n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883,
         n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893,
         n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903,
         n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913,
         n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923,
         n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933,
         n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943,
         n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953,
         n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963,
         n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973,
         n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983,
         n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993,
         n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003,
         n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013,
         n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023,
         n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033,
         n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043,
         n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053,
         n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063,
         n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073,
         n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083,
         n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093,
         n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103,
         n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113,
         n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123,
         n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133,
         n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143,
         n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153,
         n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163,
         n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173,
         n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183,
         n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193,
         n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203,
         n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213,
         n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223,
         n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233,
         n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243,
         n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253,
         n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263,
         n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273,
         n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283,
         n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293,
         n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303,
         n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313,
         n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323,
         n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333,
         n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343,
         n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353,
         n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363,
         n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373,
         n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383,
         n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393,
         n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403,
         n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413,
         n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423,
         n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433,
         n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443,
         n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453,
         n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463,
         n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473,
         n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483,
         n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493,
         n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503,
         n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
         n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
         n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
         n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
         n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
         n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
         n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613,
         n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623,
         n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
         n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643,
         n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653,
         n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663,
         n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673,
         n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683,
         n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693,
         n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703,
         n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713,
         n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723,
         n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733,
         n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743,
         n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753,
         n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763,
         n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773,
         n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783,
         n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793,
         n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803,
         n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813,
         n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823,
         n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833,
         n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843,
         n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853,
         n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863,
         n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873,
         n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883,
         n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893,
         n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903,
         n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913,
         n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923,
         n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933,
         n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943,
         n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953,
         n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963,
         n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973,
         n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983,
         n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993,
         n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003,
         n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013,
         n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023,
         n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033,
         n5034, n5035, n5036;

  INV_X2 U2365 ( .A(n2923), .ZN(n3116) );
  INV_X1 U2366 ( .A(n3117), .ZN(n2930) );
  INV_X2 U2368 ( .A(n2605), .ZN(n2639) );
  NAND3_X1 U2369 ( .A1(n2183), .A2(n2856), .A3(n2136), .ZN(n2888) );
  INV_X1 U2370 ( .A(n4604), .ZN(n2123) );
  INV_X2 U2371 ( .A(n2123), .ZN(U3149) );
  INV_X1 U2372 ( .A(STATE_REG_SCAN_IN), .ZN(n4604) );
  NOR2_X1 U2374 ( .A1(n4698), .A2(n2921), .ZN(n2908) );
  INV_X1 U2375 ( .A(n2908), .ZN(n3051) );
  CLKBUF_X2 U2376 ( .A(n2923), .Z(n3142) );
  OAI21_X1 U2377 ( .B1(n4166), .B2(n2347), .A(n2345), .ZN(n2436) );
  NAND2_X1 U2378 ( .A1(n3214), .A2(n4080), .ZN(n4241) );
  XNOR2_X1 U2379 ( .A(n2444), .B(n3768), .ZN(n3764) );
  CLKBUF_X2 U2380 ( .A(n2501), .Z(n2127) );
  NAND2_X4 U2381 ( .A1(n2488), .A2(n2487), .ZN(n2612) );
  NAND2_X2 U2382 ( .A1(n2816), .A2(n2814), .ZN(n3185) );
  OAI22_X2 U2383 ( .A1(n2242), .A2(n3532), .B1(n2820), .B2(n2240), .ZN(n3382)
         );
  AND2_X4 U2384 ( .A1(n2566), .A2(n4590), .ZN(n2606) );
  INV_X1 U2385 ( .A(n3051), .ZN(n2125) );
  INV_X1 U2386 ( .A(n3051), .ZN(n2126) );
  AND2_X1 U2387 ( .A1(n2181), .A2(n2158), .ZN(n3808) );
  INV_X1 U2388 ( .A(n3440), .ZN(n3924) );
  OR2_X1 U2389 ( .A1(n2986), .A2(n2200), .ZN(n2199) );
  NAND2_X1 U2390 ( .A1(n3400), .A2(n3535), .ZN(n4037) );
  INV_X1 U2391 ( .A(n3535), .ZN(n3367) );
  INV_X2 U2392 ( .A(n3789), .ZN(n2909) );
  CLKBUF_X2 U2393 ( .A(n2639), .Z(n3155) );
  NAND2_X1 U2394 ( .A1(n2606), .A2(REG1_REG_0__SCAN_IN), .ZN(n2584) );
  NAND2_X1 U2395 ( .A1(n2895), .A2(n4094), .ZN(n3140) );
  OR2_X1 U2396 ( .A1(n2189), .A2(n2188), .ZN(n2186) );
  OR2_X1 U2397 ( .A1(n2190), .A2(n2188), .ZN(n2187) );
  OAI21_X1 U2398 ( .B1(n3837), .B2(n2333), .A(n2332), .ZN(n3130) );
  NAND2_X1 U2399 ( .A1(n3837), .A2(n3834), .ZN(n3872) );
  AOI21_X1 U2400 ( .B1(n3202), .B2(n4414), .A(n3201), .ZN(n4486) );
  NOR2_X1 U2401 ( .A1(n3808), .A2(n3814), .ZN(n3049) );
  NAND3_X1 U2402 ( .A1(n2308), .A2(n2307), .A3(n3008), .ZN(n3852) );
  NAND2_X1 U2403 ( .A1(n4438), .A2(n4015), .ZN(n4439) );
  AOI21_X1 U2404 ( .B1(n4425), .B2(n2736), .A(n2735), .ZN(n4404) );
  NAND2_X1 U2405 ( .A1(n2281), .A2(n2280), .ZN(n4425) );
  NAND2_X1 U2406 ( .A1(n2823), .A2(n4052), .ZN(n3650) );
  AND2_X1 U2407 ( .A1(n2199), .A2(n3487), .ZN(n2987) );
  OR2_X1 U2408 ( .A1(n2972), .A2(n2971), .ZN(n2984) );
  OR2_X1 U2409 ( .A1(n3988), .A2(n2710), .ZN(n2712) );
  AND2_X1 U2410 ( .A1(n2954), .A2(n3722), .ZN(n3726) );
  XNOR2_X1 U2411 ( .A(n2423), .B(n4146), .ZN(n4144) );
  NAND2_X1 U2412 ( .A1(n2549), .A2(REG3_REG_19__SCAN_IN), .ZN(n2765) );
  NAND2_X1 U2413 ( .A1(n3278), .A2(n2418), .ZN(n2423) );
  INV_X1 U2414 ( .A(n2750), .ZN(n2549) );
  OR2_X1 U2415 ( .A1(n2962), .A2(n2169), .ZN(n2960) );
  XNOR2_X1 U2416 ( .A(n2407), .B(n3314), .ZN(n3317) );
  NAND2_X1 U2417 ( .A1(n2279), .A2(n2888), .ZN(n2906) );
  AND4_X1 U2418 ( .A1(n2595), .A2(n2594), .A3(n2593), .A4(n2592), .ZN(n3789)
         );
  NAND4_X1 U2419 ( .A1(n2610), .A2(n2609), .A3(n2608), .A4(n2607), .ZN(n3535)
         );
  NAND2_X1 U2420 ( .A1(n2580), .A2(n2579), .ZN(n3455) );
  XNOR2_X1 U2421 ( .A(n2813), .B(n2812), .ZN(n2816) );
  NAND2_X1 U2422 ( .A1(n2811), .A2(n2461), .ZN(n4094) );
  NAND2_X1 U2423 ( .A1(n2811), .A2(IR_REG_31__SCAN_IN), .ZN(n2813) );
  XNOR2_X1 U2424 ( .A(n2485), .B(IR_REG_21__SCAN_IN), .ZN(n2814) );
  OR2_X1 U2425 ( .A1(n2481), .A2(n2360), .ZN(n2482) );
  AND2_X1 U2426 ( .A1(n2484), .A2(n2483), .ZN(n2485) );
  XNOR2_X1 U2427 ( .A(n2470), .B(IR_REG_26__SCAN_IN), .ZN(n2856) );
  OAI21_X1 U2428 ( .B1(n2489), .B2(n2486), .A(n2231), .ZN(n2488) );
  XNOR2_X1 U2429 ( .A(n2563), .B(IR_REG_29__SCAN_IN), .ZN(n4590) );
  NOR2_X1 U2430 ( .A1(n2476), .A2(n2475), .ZN(n2481) );
  NAND2_X1 U2431 ( .A1(n2491), .A2(IR_REG_31__SCAN_IN), .ZN(n2470) );
  NAND2_X1 U2432 ( .A1(n2476), .A2(IR_REG_31__SCAN_IN), .ZN(n2484) );
  OR2_X1 U2433 ( .A1(n2471), .A2(IR_REG_25__SCAN_IN), .ZN(n2491) );
  NAND2_X1 U2434 ( .A1(n2385), .A2(n2182), .ZN(n2476) );
  NAND3_X1 U2435 ( .A1(n2277), .A2(n2276), .A3(n2275), .ZN(n2501) );
  NAND2_X1 U2436 ( .A1(n2555), .A2(IR_REG_27__SCAN_IN), .ZN(n2487) );
  NOR2_X1 U2437 ( .A1(IR_REG_20__SCAN_IN), .A2(IR_REG_21__SCAN_IN), .ZN(n2474)
         );
  INV_X1 U2438 ( .A(IR_REG_28__SCAN_IN), .ZN(n2555) );
  INV_X1 U2439 ( .A(IR_REG_27__SCAN_IN), .ZN(n2486) );
  INV_X1 U2440 ( .A(IR_REG_4__SCAN_IN), .ZN(n2405) );
  INV_X1 U2441 ( .A(IR_REG_3__SCAN_IN), .ZN(n2399) );
  NOR2_X1 U2442 ( .A1(IR_REG_15__SCAN_IN), .A2(IR_REG_6__SCAN_IN), .ZN(n2167)
         );
  NOR2_X1 U2443 ( .A1(IR_REG_12__SCAN_IN), .A2(IR_REG_10__SCAN_IN), .ZN(n2168)
         );
  INV_X1 U2444 ( .A(IR_REG_1__SCAN_IN), .ZN(n2306) );
  INV_X1 U2445 ( .A(IR_REG_0__SCAN_IN), .ZN(n2305) );
  INV_X2 U2446 ( .A(n4265), .ZN(n4306) );
  INV_X4 U2447 ( .A(n2898), .ZN(n2921) );
  INV_X1 U2448 ( .A(n3117), .ZN(n2128) );
  NOR2_X2 U2449 ( .A1(n4429), .A2(n4397), .ZN(n4389) );
  NOR2_X1 U2450 ( .A1(n4698), .A2(n2921), .ZN(n2129) );
  AOI21_X1 U2452 ( .B1(n2263), .B2(n2261), .A(n2260), .ZN(n2259) );
  INV_X1 U2453 ( .A(n4046), .ZN(n2261) );
  INV_X1 U2454 ( .A(n4045), .ZN(n2260) );
  INV_X1 U2455 ( .A(n4603), .ZN(n2507) );
  NOR2_X1 U2456 ( .A1(n4618), .A2(n2528), .ZN(n2530) );
  AND2_X1 U2457 ( .A1(n2322), .A2(n2316), .ZN(n2315) );
  NOR2_X1 U2458 ( .A1(n3177), .A2(n2323), .ZN(n2322) );
  NAND2_X1 U2459 ( .A1(n2319), .A2(n2317), .ZN(n2316) );
  INV_X1 U2460 ( .A(n2324), .ZN(n2323) );
  INV_X1 U2461 ( .A(n2319), .ZN(n2318) );
  NAND2_X1 U2462 ( .A1(n4362), .A2(n2882), .ZN(n2302) );
  NAND2_X1 U2463 ( .A1(n3826), .A2(n4360), .ZN(n2303) );
  AND2_X1 U2464 ( .A1(n2895), .A2(n4591), .ZN(n3125) );
  INV_X1 U2465 ( .A(n3917), .ZN(n2335) );
  AND2_X1 U2466 ( .A1(n2612), .A2(DATAI_25_), .ZN(n3843) );
  NOR2_X1 U2467 ( .A1(n3898), .A2(n2329), .ZN(n2327) );
  OAI21_X1 U2468 ( .B1(n2897), .B2(n2906), .A(n2899), .ZN(n2900) );
  OR2_X1 U2470 ( .A1(n4253), .A2(n2605), .ZN(n2571) );
  INV_X1 U2471 ( .A(n2606), .ZN(n3153) );
  NAND2_X1 U2472 ( .A1(n4182), .A2(n2522), .ZN(n2523) );
  OAI21_X1 U2473 ( .B1(n2442), .B2(IR_REG_14__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2448) );
  NAND2_X1 U2474 ( .A1(n2532), .A2(n4989), .ZN(n2364) );
  INV_X1 U2475 ( .A(n4646), .ZN(n2217) );
  OAI21_X1 U2476 ( .B1(n4279), .B2(n2149), .A(n2799), .ZN(n4259) );
  INV_X1 U2477 ( .A(n2286), .ZN(n2285) );
  INV_X1 U2478 ( .A(n4414), .ZN(n4468) );
  OR2_X1 U2479 ( .A1(n3442), .A2(n2895), .ZN(n4693) );
  INV_X1 U2480 ( .A(n3941), .ZN(n3927) );
  NOR2_X1 U2481 ( .A1(n2212), .A2(n2210), .ZN(n2209) );
  INV_X1 U2482 ( .A(n4160), .ZN(n2212) );
  INV_X1 U2483 ( .A(n4178), .ZN(n2347) );
  INV_X1 U2484 ( .A(n4049), .ZN(n2264) );
  INV_X1 U2485 ( .A(n2961), .ZN(n2169) );
  INV_X1 U2486 ( .A(n3865), .ZN(n2196) );
  OAI21_X1 U2487 ( .B1(n2408), .B2(n2354), .A(n2413), .ZN(n2349) );
  NOR2_X1 U2488 ( .A1(n2821), .A2(n2246), .ZN(n2245) );
  INV_X1 U2489 ( .A(n4034), .ZN(n2246) );
  INV_X1 U2490 ( .A(n3454), .ZN(n4027) );
  AND2_X1 U2491 ( .A1(n4388), .A2(n4369), .ZN(n2221) );
  NAND2_X1 U2492 ( .A1(n2480), .A2(IR_REG_31__SCAN_IN), .ZN(n2857) );
  AND2_X1 U2493 ( .A1(n2168), .A2(n2167), .ZN(n2382) );
  NAND2_X1 U2494 ( .A1(n3002), .A2(n3712), .ZN(n2308) );
  NAND2_X1 U2495 ( .A1(n3004), .A2(n3003), .ZN(n2307) );
  INV_X1 U2496 ( .A(n3908), .ZN(n2191) );
  AND2_X1 U2497 ( .A1(n2130), .A2(n3163), .ZN(n2334) );
  NAND2_X1 U2498 ( .A1(n2612), .A2(DATAI_1_), .ZN(n2579) );
  NAND2_X1 U2499 ( .A1(n2578), .A2(n2127), .ZN(n2580) );
  OR2_X1 U2500 ( .A1(n2765), .A2(n2550), .ZN(n2772) );
  INV_X1 U2501 ( .A(n2612), .ZN(n2728) );
  NAND2_X1 U2502 ( .A1(n2171), .A2(n3486), .ZN(n2176) );
  INV_X1 U2503 ( .A(n3487), .ZN(n2172) );
  INV_X1 U2504 ( .A(n4110), .ZN(n3392) );
  INV_X1 U2505 ( .A(n4107), .ZN(n3554) );
  NAND2_X1 U2506 ( .A1(n2477), .A2(n2859), .ZN(n2183) );
  INV_X1 U2507 ( .A(IR_REG_20__SCAN_IN), .ZN(n2812) );
  AND4_X1 U2508 ( .A1(n2625), .A2(n2624), .A3(n2623), .A4(n2622), .ZN(n2626)
         );
  NAND2_X1 U2509 ( .A1(n4123), .A2(n2403), .ZN(n2407) );
  NAND2_X1 U2510 ( .A1(n2203), .A2(n2509), .ZN(n2510) );
  NAND2_X1 U2511 ( .A1(n4125), .A2(REG1_REG_3__SCAN_IN), .ZN(n2203) );
  INV_X1 U2512 ( .A(n4136), .ZN(n2354) );
  INV_X1 U2513 ( .A(REG2_REG_4__SCAN_IN), .ZN(n2355) );
  OAI21_X1 U2514 ( .B1(n3276), .B2(n3275), .A(n2517), .ZN(n2518) );
  NOR2_X1 U2515 ( .A1(n2518), .A2(n4146), .ZN(n2214) );
  NAND2_X1 U2516 ( .A1(n2339), .A2(n2337), .ZN(n2430) );
  INV_X1 U2517 ( .A(n2338), .ZN(n2337) );
  NAND2_X1 U2518 ( .A1(n4144), .A2(n2342), .ZN(n2339) );
  OAI21_X1 U2519 ( .B1(n2424), .B2(n2343), .A(n2427), .ZN(n2338) );
  NAND2_X1 U2520 ( .A1(n4190), .A2(n2437), .ZN(n2362) );
  OR2_X1 U2521 ( .A1(n2362), .A2(n4595), .ZN(n4200) );
  NAND2_X1 U2522 ( .A1(n2361), .A2(n2138), .ZN(n2444) );
  NAND2_X1 U2523 ( .A1(n4190), .A2(n2134), .ZN(n2361) );
  NOR2_X1 U2524 ( .A1(n4616), .A2(n2451), .ZN(n2455) );
  AND2_X1 U2525 ( .A1(n4622), .A2(REG2_REG_15__SCAN_IN), .ZN(n2451) );
  NAND2_X1 U2526 ( .A1(n4641), .A2(n2164), .ZN(n2459) );
  INV_X1 U2527 ( .A(n4663), .ZN(n2363) );
  INV_X1 U2528 ( .A(n2216), .ZN(n2215) );
  OAI21_X1 U2529 ( .B1(n2531), .B2(n2217), .A(n2165), .ZN(n2216) );
  INV_X1 U2530 ( .A(n4654), .ZN(n2534) );
  NAND2_X1 U2531 ( .A1(n2314), .A2(n2313), .ZN(n3212) );
  AOI21_X1 U2532 ( .B1(n2315), .B2(n2318), .A(n2151), .ZN(n2313) );
  OR2_X1 U2533 ( .A1(n2845), .A2(n3167), .ZN(n3109) );
  NAND2_X1 U2534 ( .A1(n2789), .A2(n2788), .ZN(n4279) );
  NAND2_X1 U2535 ( .A1(n2551), .A2(REG3_REG_22__SCAN_IN), .ZN(n2781) );
  INV_X1 U2536 ( .A(n2772), .ZN(n2551) );
  NAND2_X1 U2537 ( .A1(n2299), .A2(n2302), .ZN(n2294) );
  NAND2_X1 U2538 ( .A1(n2293), .A2(n2302), .ZN(n2292) );
  INV_X1 U2539 ( .A(n2296), .ZN(n2293) );
  AOI21_X1 U2540 ( .B1(n2299), .B2(n2297), .A(n2153), .ZN(n2296) );
  INV_X1 U2541 ( .A(n2289), .ZN(n4319) );
  AOI21_X1 U2542 ( .B1(n4386), .B2(n2292), .A(n2290), .ZN(n2289) );
  NAND2_X1 U2543 ( .A1(n2291), .A2(n4320), .ZN(n2290) );
  NAND2_X1 U2544 ( .A1(n2292), .A2(n2294), .ZN(n2291) );
  INV_X1 U2545 ( .A(n2284), .ZN(n2283) );
  OAI21_X1 U2546 ( .B1(n2143), .B2(n2285), .A(n4450), .ZN(n2284) );
  NAND2_X1 U2547 ( .A1(n2133), .A2(n2144), .ZN(n2286) );
  AND2_X1 U2548 ( .A1(n2691), .A2(n2690), .ZN(n4463) );
  INV_X1 U2549 ( .A(n4470), .ZN(n2831) );
  NAND2_X1 U2550 ( .A1(n3382), .A2(n4039), .ZN(n2822) );
  OAI21_X1 U2551 ( .B1(n2612), .B2(n4602), .A(n2613), .ZN(n3400) );
  NAND2_X1 U2552 ( .A1(n2612), .A2(n2611), .ZN(n2613) );
  AND2_X1 U2553 ( .A1(n4034), .A2(n4032), .ZN(n4004) );
  INV_X1 U2554 ( .A(n3296), .ZN(n3451) );
  NAND2_X1 U2555 ( .A1(n3790), .A2(n3296), .ZN(n3454) );
  NOR3_X1 U2556 ( .A1(n3206), .A2(n4223), .A3(n3970), .ZN(n4221) );
  NAND2_X1 U2557 ( .A1(n4222), .A2(n3207), .ZN(n4490) );
  NAND2_X1 U2558 ( .A1(n3221), .A2(n3220), .ZN(n4227) );
  NOR2_X1 U2559 ( .A1(n3928), .A2(n2224), .ZN(n2223) );
  INV_X1 U2560 ( .A(n2225), .ZN(n2224) );
  OR2_X2 U2561 ( .A1(n4426), .A2(n4427), .ZN(n4429) );
  NAND2_X1 U2562 ( .A1(n4366), .A2(n4693), .ZN(n4545) );
  INV_X1 U2563 ( .A(n4698), .ZN(n4706) );
  AND3_X1 U2564 ( .A1(n2876), .A2(n2875), .A3(n3124), .ZN(n3228) );
  NAND3_X1 U2565 ( .A1(n2856), .A2(n2862), .A3(n2861), .ZN(n3253) );
  XNOR2_X1 U2566 ( .A(n2857), .B(n4840), .ZN(n3136) );
  OR2_X1 U2567 ( .A1(n2432), .A2(n2389), .ZN(n2442) );
  INV_X1 U2568 ( .A(n3163), .ZN(n3164) );
  AOI211_X1 U2569 ( .C1(n3799), .C2(n2131), .A(n2135), .B(n2154), .ZN(n2174)
         );
  MUX2_X1 U2570 ( .A(n4603), .B(DATAI_3_), .S(n2612), .Z(n3507) );
  AND2_X1 U2571 ( .A1(n2802), .A2(n2801), .ZN(n4274) );
  NAND2_X1 U2572 ( .A1(n2612), .A2(n2615), .ZN(n2616) );
  OR2_X1 U2573 ( .A1(n2612), .A2(n2614), .ZN(n2617) );
  INV_X1 U2574 ( .A(n3400), .ZN(n3396) );
  OR3_X1 U2575 ( .A1(n3156), .A2(n4606), .A3(n4097), .ZN(n3920) );
  AND2_X1 U2576 ( .A1(n3148), .A2(n4447), .ZN(n3941) );
  OAI21_X1 U2577 ( .B1(n2127), .B2(n2500), .A(n2278), .ZN(n2503) );
  NAND2_X1 U2578 ( .A1(n2127), .A2(n2500), .ZN(n2278) );
  XNOR2_X1 U2579 ( .A(n2518), .B(n4599), .ZN(n4150) );
  NAND2_X1 U2580 ( .A1(n4150), .A2(REG1_REG_8__SCAN_IN), .ZN(n4149) );
  XNOR2_X1 U2581 ( .A(n2430), .B(n4172), .ZN(n4167) );
  OAI21_X1 U2582 ( .B1(n4171), .B2(n2207), .A(n2204), .ZN(n4182) );
  AOI21_X1 U2583 ( .B1(n2520), .B2(n2206), .A(n2205), .ZN(n2204) );
  INV_X1 U2584 ( .A(REG1_REG_10__SCAN_IN), .ZN(n2206) );
  XNOR2_X1 U2585 ( .A(n2523), .B(n4195), .ZN(n4194) );
  NAND2_X1 U2586 ( .A1(n4194), .A2(REG1_REG_12__SCAN_IN), .ZN(n2202) );
  OAI21_X1 U2587 ( .B1(n2438), .B2(IR_REG_12__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2440) );
  NAND2_X1 U2588 ( .A1(n2325), .A2(n2324), .ZN(n4240) );
  NAND2_X1 U2589 ( .A1(n2321), .A2(n2319), .ZN(n2325) );
  NOR2_X1 U2590 ( .A1(n4237), .A2(n2268), .ZN(n4500) );
  INV_X1 U2591 ( .A(n2269), .ZN(n2268) );
  AOI21_X1 U2592 ( .B1(n4239), .B2(n4418), .A(n4238), .ZN(n2269) );
  XOR2_X1 U2593 ( .A(n4020), .B(n3176), .Z(n4251) );
  NAND2_X1 U2594 ( .A1(n2321), .A2(n2810), .ZN(n3176) );
  OR2_X1 U2595 ( .A1(n4490), .A2(n4706), .ZN(n4495) );
  NOR2_X1 U2596 ( .A1(n3994), .A2(n2235), .ZN(n4003) );
  NAND2_X1 U2597 ( .A1(n2237), .A2(n2236), .ZN(n2235) );
  INV_X1 U2598 ( .A(n3996), .ZN(n2237) );
  INV_X1 U2599 ( .A(n2373), .ZN(n2317) );
  NOR2_X1 U2600 ( .A1(n3188), .A2(n2253), .ZN(n2252) );
  INV_X1 U2601 ( .A(n4075), .ZN(n2253) );
  INV_X1 U2602 ( .A(n3959), .ZN(n2250) );
  NAND2_X1 U2603 ( .A1(n3367), .A2(n3396), .ZN(n4035) );
  NOR2_X1 U2604 ( .A1(IR_REG_16__SCAN_IN), .A2(IR_REG_8__SCAN_IN), .ZN(n2378)
         );
  XNOR2_X1 U2605 ( .A(n2197), .B(n2930), .ZN(n2955) );
  NAND2_X1 U2606 ( .A1(n2945), .A2(n2198), .ZN(n2197) );
  NAND2_X1 U2607 ( .A1(n3490), .A2(n2923), .ZN(n2198) );
  NAND2_X1 U2608 ( .A1(n2984), .A2(n2201), .ZN(n2200) );
  INV_X1 U2609 ( .A(n2985), .ZN(n2201) );
  INV_X1 U2610 ( .A(n3185), .ZN(n2279) );
  NAND2_X1 U2611 ( .A1(n3322), .A2(n2397), .ZN(n2402) );
  NAND2_X1 U2612 ( .A1(n3328), .A2(n2506), .ZN(n2508) );
  NOR2_X1 U2613 ( .A1(n2343), .A2(n2344), .ZN(n2342) );
  NAND2_X1 U2614 ( .A1(n2211), .A2(n2208), .ZN(n2519) );
  AOI21_X1 U2615 ( .B1(n2214), .B2(n4160), .A(n2140), .ZN(n2211) );
  NAND2_X1 U2616 ( .A1(n4150), .A2(n2209), .ZN(n2208) );
  INV_X1 U2617 ( .A(n2346), .ZN(n2345) );
  OAI21_X1 U2618 ( .B1(n2841), .B2(n2251), .A(n2248), .ZN(n4235) );
  INV_X1 U2619 ( .A(n2252), .ZN(n2251) );
  AND2_X1 U2620 ( .A1(n4082), .A2(n2249), .ZN(n2248) );
  NAND2_X1 U2621 ( .A1(n2252), .A2(n2250), .ZN(n2249) );
  NAND2_X1 U2622 ( .A1(n4281), .A2(n4075), .ZN(n4261) );
  NAND2_X1 U2623 ( .A1(n2841), .A2(n3959), .ZN(n4281) );
  INV_X1 U2624 ( .A(n2141), .ZN(n2297) );
  INV_X1 U2625 ( .A(REG3_REG_10__SCAN_IN), .ZN(n2672) );
  INV_X1 U2626 ( .A(n4044), .ZN(n2265) );
  AND2_X1 U2627 ( .A1(n3592), .A2(n2649), .ZN(n2650) );
  AND2_X1 U2628 ( .A1(n3968), .A2(DATAI_29_), .ZN(n3970) );
  NOR2_X1 U2629 ( .A1(n2227), .A2(n3189), .ZN(n3222) );
  NOR2_X1 U2630 ( .A1(n3843), .A2(n2226), .ZN(n2225) );
  INV_X1 U2631 ( .A(n4290), .ZN(n2226) );
  NOR2_X1 U2632 ( .A1(n3431), .A2(n3473), .ZN(n3471) );
  NAND2_X1 U2633 ( .A1(n2257), .A2(n2259), .ZN(n3466) );
  NAND2_X1 U2634 ( .A1(n2258), .A2(n2263), .ZN(n2257) );
  INV_X1 U2635 ( .A(n3576), .ZN(n2258) );
  NAND2_X1 U2636 ( .A1(n4044), .A2(n4046), .ZN(n3592) );
  OR2_X1 U2637 ( .A1(n3253), .A2(n2874), .ZN(n3124) );
  OR2_X1 U2638 ( .A1(n3138), .A2(n3146), .ZN(n3180) );
  INV_X1 U2639 ( .A(IR_REG_22__SCAN_IN), .ZN(n4820) );
  INV_X1 U2640 ( .A(B_REG_SCAN_IN), .ZN(n4976) );
  NAND2_X1 U2641 ( .A1(n2230), .A2(IR_REG_31__SCAN_IN), .ZN(n2489) );
  AND2_X1 U2642 ( .A1(n2560), .A2(n2288), .ZN(n2182) );
  INV_X1 U2643 ( .A(IR_REG_18__SCAN_IN), .ZN(n2288) );
  INV_X1 U2644 ( .A(IR_REG_12__SCAN_IN), .ZN(n4778) );
  INV_X1 U2645 ( .A(IR_REG_10__SCAN_IN), .ZN(n2387) );
  NAND2_X1 U2646 ( .A1(n2305), .A2(n2306), .ZN(n2358) );
  NAND2_X1 U2647 ( .A1(n2178), .A2(n3415), .ZN(n2980) );
  AND2_X1 U2648 ( .A1(n2937), .A2(n2180), .ZN(n2179) );
  INV_X1 U2649 ( .A(n3416), .ZN(n2180) );
  AND2_X1 U2650 ( .A1(n3020), .A2(n3019), .ZN(n3850) );
  AND2_X1 U2651 ( .A1(n3968), .A2(DATAI_23_), .ZN(n3070) );
  INV_X1 U2652 ( .A(n2960), .ZN(n2963) );
  XNOR2_X1 U2653 ( .A(n2956), .B(n2955), .ZN(n2959) );
  INV_X1 U2654 ( .A(n3887), .ZN(n3058) );
  AOI21_X1 U2655 ( .B1(n3837), .B2(n3836), .A(n3835), .ZN(n3874) );
  NAND2_X1 U2656 ( .A1(n3365), .A2(n3366), .ZN(n2304) );
  OR2_X1 U2657 ( .A1(n2693), .A2(n2692), .ZN(n2700) );
  NAND2_X1 U2658 ( .A1(n2330), .A2(n3822), .ZN(n2329) );
  NAND2_X1 U2659 ( .A1(n2162), .A2(n3058), .ZN(n2330) );
  NAND2_X1 U2660 ( .A1(n3811), .A2(n2331), .ZN(n2328) );
  AND2_X1 U2661 ( .A1(n3059), .A2(n2162), .ZN(n2331) );
  NAND2_X1 U2662 ( .A1(n3479), .A2(n2985), .ZN(n2974) );
  INV_X1 U2663 ( .A(n2193), .ZN(n2192) );
  OAI21_X1 U2664 ( .B1(n3025), .B2(n2194), .A(n3864), .ZN(n2193) );
  OR2_X1 U2665 ( .A1(n3026), .A2(n2196), .ZN(n2194) );
  OR2_X1 U2666 ( .A1(n3025), .A2(n2196), .ZN(n2195) );
  INV_X1 U2667 ( .A(REG3_REG_6__SCAN_IN), .ZN(n2640) );
  INV_X1 U2668 ( .A(IR_REG_19__SCAN_IN), .ZN(n2473) );
  AND4_X1 U2669 ( .A1(n2660), .A2(n2659), .A3(n2658), .A4(n2657), .ZN(n3467)
         );
  XNOR2_X1 U2670 ( .A(n2508), .B(n2507), .ZN(n4125) );
  XNOR2_X1 U2671 ( .A(n2402), .B(n2507), .ZN(n4124) );
  NAND2_X1 U2672 ( .A1(n2350), .A2(n2348), .ZN(n2415) );
  NAND2_X1 U2673 ( .A1(n3317), .A2(n2353), .ZN(n2350) );
  NOR2_X1 U2674 ( .A1(n2354), .A2(n2355), .ZN(n2353) );
  INV_X1 U2675 ( .A(IR_REG_7__SCAN_IN), .ZN(n4962) );
  INV_X1 U2676 ( .A(n4155), .ZN(n2343) );
  INV_X1 U2677 ( .A(n4183), .ZN(n2205) );
  NAND2_X1 U2678 ( .A1(n4171), .A2(REG1_REG_10__SCAN_IN), .ZN(n4170) );
  NAND2_X1 U2679 ( .A1(n4206), .A2(n2525), .ZN(n2526) );
  OAI21_X1 U2680 ( .B1(n3764), .B2(n2366), .A(n2365), .ZN(n4616) );
  NAND2_X1 U2681 ( .A1(n2367), .A2(REG2_REG_14__SCAN_IN), .ZN(n2366) );
  INV_X1 U2682 ( .A(n4617), .ZN(n2367) );
  OAI22_X1 U2683 ( .A1(n3766), .A2(n2218), .B1(n2142), .B2(n4619), .ZN(n4618)
         );
  OR2_X1 U2684 ( .A1(n4619), .A2(n4770), .ZN(n2218) );
  OR2_X1 U2685 ( .A1(n3766), .A2(n4770), .ZN(n2219) );
  XNOR2_X1 U2686 ( .A(n2455), .B(n2529), .ZN(n4632) );
  NAND2_X1 U2687 ( .A1(n4632), .A2(n4631), .ZN(n4630) );
  NAND2_X1 U2688 ( .A1(n4633), .A2(n2531), .ZN(n4645) );
  INV_X1 U2689 ( .A(n4606), .ZN(n3307) );
  NAND2_X1 U2690 ( .A1(n4645), .A2(n4646), .ZN(n4644) );
  AND2_X1 U2691 ( .A1(n3192), .A2(n3973), .ZN(n4022) );
  NAND2_X1 U2692 ( .A1(n4234), .A2(n3174), .ZN(n2324) );
  NOR2_X1 U2693 ( .A1(n3175), .A2(n2320), .ZN(n2319) );
  INV_X1 U2694 ( .A(n2810), .ZN(n2320) );
  AND2_X1 U2695 ( .A1(n2798), .A2(n2797), .ZN(n4265) );
  OR2_X1 U2696 ( .A1(n3877), .A2(n2605), .ZN(n2798) );
  AND2_X1 U2697 ( .A1(n2779), .A2(n2778), .ZN(n4341) );
  INV_X1 U2698 ( .A(n2371), .ZN(n2300) );
  NAND2_X1 U2699 ( .A1(n4386), .A2(n2757), .ZN(n2301) );
  AOI21_X1 U2700 ( .B1(n2283), .B2(n2285), .A(n2145), .ZN(n2280) );
  INV_X1 U2701 ( .A(n2720), .ZN(n2547) );
  AND2_X1 U2702 ( .A1(n4457), .A2(n4456), .ZN(n4444) );
  INV_X1 U2703 ( .A(n2239), .ZN(n2238) );
  OAI21_X1 U2704 ( .B1(n4058), .B2(n2829), .A(n3947), .ZN(n2239) );
  AND2_X1 U2705 ( .A1(n2708), .A2(n2707), .ZN(n3638) );
  NAND2_X1 U2706 ( .A1(n2828), .A2(n4058), .ZN(n3948) );
  OR2_X1 U2707 ( .A1(n2673), .A2(n2672), .ZN(n2681) );
  NAND2_X1 U2708 ( .A1(n2544), .A2(REG3_REG_11__SCAN_IN), .ZN(n2693) );
  INV_X1 U2709 ( .A(n2681), .ZN(n2544) );
  AND2_X1 U2710 ( .A1(n3649), .A2(n3647), .ZN(n3988) );
  INV_X1 U2711 ( .A(n3490), .ZN(n3701) );
  INV_X1 U2712 ( .A(n4417), .ZN(n4462) );
  AOI21_X1 U2713 ( .B1(n2132), .B2(n2262), .A(n2256), .ZN(n2255) );
  NAND2_X1 U2714 ( .A1(n3576), .A2(n2132), .ZN(n2254) );
  INV_X1 U2715 ( .A(n4050), .ZN(n2256) );
  OAI21_X1 U2716 ( .B1(n3465), .B2(n2671), .A(n2670), .ZN(n3528) );
  OR2_X1 U2717 ( .A1(n2655), .A2(n4730), .ZN(n2664) );
  OAI21_X1 U2718 ( .B1(n3576), .B2(n2265), .A(n4046), .ZN(n3426) );
  NAND2_X1 U2719 ( .A1(n2247), .A2(n4037), .ZN(n2240) );
  INV_X1 U2720 ( .A(n2243), .ZN(n2242) );
  OAI21_X1 U2721 ( .B1(n2245), .B2(n2244), .A(n4041), .ZN(n2243) );
  NAND2_X1 U2722 ( .A1(n2241), .A2(n4037), .ZN(n3533) );
  NAND2_X1 U2723 ( .A1(n2820), .A2(n2245), .ZN(n2241) );
  NOR2_X1 U2724 ( .A1(n3506), .A2(n3507), .ZN(n3505) );
  NAND2_X1 U2725 ( .A1(n2589), .A2(n2588), .ZN(n3355) );
  NAND2_X1 U2726 ( .A1(n2612), .A2(DATAI_2_), .ZN(n2588) );
  OR2_X1 U2727 ( .A1(n2612), .A2(n2587), .ZN(n2589) );
  NAND2_X1 U2728 ( .A1(n3354), .A2(n3350), .ZN(n3506) );
  INV_X1 U2729 ( .A(n3355), .ZN(n3350) );
  AND2_X1 U2730 ( .A1(n3125), .A2(n3307), .ZN(n4417) );
  NAND2_X1 U2731 ( .A1(n4092), .A2(n2844), .ZN(n4414) );
  OR2_X1 U2732 ( .A1(n2590), .A2(n2573), .ZN(n2575) );
  NAND2_X1 U2733 ( .A1(n2815), .A2(n4094), .ZN(n4366) );
  AND2_X1 U2734 ( .A1(n3124), .A2(n4727), .ZN(n3182) );
  OR2_X1 U2735 ( .A1(n3206), .A2(n3970), .ZN(n4222) );
  AND2_X1 U2736 ( .A1(n3968), .A2(DATAI_30_), .ZN(n4223) );
  AND2_X1 U2737 ( .A1(n3968), .A2(DATAI_28_), .ZN(n3223) );
  NAND2_X1 U2738 ( .A1(n3222), .A2(n3217), .ZN(n3206) );
  NAND2_X1 U2739 ( .A1(n4289), .A2(n2225), .ZN(n4271) );
  NAND2_X1 U2740 ( .A1(n4389), .A2(n2137), .ZN(n4347) );
  INV_X1 U2741 ( .A(n4382), .ZN(n4388) );
  MUX2_X1 U2742 ( .A(n4594), .B(DATAI_14_), .S(n3968), .Z(n3643) );
  NOR2_X1 U2743 ( .A1(n3690), .A2(n3643), .ZN(n4457) );
  NAND2_X1 U2744 ( .A1(n3614), .A2(n2232), .ZN(n3690) );
  NOR2_X1 U2745 ( .A1(n3686), .A2(n3652), .ZN(n2232) );
  AND2_X1 U2746 ( .A1(n3471), .A2(n2881), .ZN(n3613) );
  OR2_X1 U2747 ( .A1(n3399), .A2(n2228), .ZN(n3582) );
  NAND2_X1 U2748 ( .A1(n2880), .A2(n3538), .ZN(n2228) );
  XNOR2_X1 U2749 ( .A(n2472), .B(n2469), .ZN(n2863) );
  XNOR2_X1 U2750 ( .A(n2860), .B(n2859), .ZN(n2878) );
  NAND2_X1 U2751 ( .A1(n2858), .A2(IR_REG_31__SCAN_IN), .ZN(n2860) );
  INV_X1 U2752 ( .A(n2814), .ZN(n4023) );
  INV_X1 U2753 ( .A(IR_REG_17__SCAN_IN), .ZN(n2391) );
  INV_X1 U2754 ( .A(IR_REG_16__SCAN_IN), .ZN(n2453) );
  NAND2_X1 U2755 ( .A1(n2432), .A2(IR_REG_31__SCAN_IN), .ZN(n2434) );
  INV_X1 U2756 ( .A(IR_REG_11__SCAN_IN), .ZN(n4767) );
  NOR2_X1 U2757 ( .A1(n2425), .A2(IR_REG_9__SCAN_IN), .ZN(n2428) );
  OR3_X1 U2758 ( .A1(n2417), .A2(IR_REG_7__SCAN_IN), .A3(IR_REG_8__SCAN_IN), 
        .ZN(n2425) );
  NAND2_X1 U2759 ( .A1(n2357), .A2(n2356), .ZN(n2498) );
  NAND3_X1 U2760 ( .A1(n2358), .A2(n2359), .A3(IR_REG_31__SCAN_IN), .ZN(n2357)
         );
  OAI21_X1 U2761 ( .B1(n2395), .B2(n2360), .A(IR_REG_2__SCAN_IN), .ZN(n2356)
         );
  INV_X1 U2762 ( .A(n2358), .ZN(n2395) );
  INV_X1 U2763 ( .A(n2888), .ZN(n3299) );
  NAND2_X1 U2764 ( .A1(n2612), .A2(n4733), .ZN(n2630) );
  INV_X1 U2765 ( .A(n3070), .ZN(n4313) );
  INV_X1 U2766 ( .A(n3920), .ZN(n3937) );
  AND2_X1 U2767 ( .A1(n2762), .A2(n2761), .ZN(n4385) );
  AOI21_X1 U2768 ( .B1(n2334), .B2(n2173), .A(n2150), .ZN(n2332) );
  INV_X1 U2769 ( .A(n2334), .ZN(n2333) );
  INV_X1 U2770 ( .A(n3455), .ZN(n3798) );
  AND3_X1 U2771 ( .A1(n2704), .A2(n2703), .A3(n2702), .ZN(n3780) );
  NAND2_X1 U2772 ( .A1(n3841), .A2(n3888), .ZN(n2188) );
  INV_X1 U2773 ( .A(n3874), .ZN(n2190) );
  NAND2_X1 U2774 ( .A1(n3872), .A2(n3875), .ZN(n2189) );
  NOR2_X1 U2775 ( .A1(n3841), .A2(n3945), .ZN(n2185) );
  NAND2_X1 U2776 ( .A1(n2612), .A2(DATAI_24_), .ZN(n4290) );
  NAND2_X1 U2777 ( .A1(n2612), .A2(DATAI_0_), .ZN(n2581) );
  INV_X1 U2778 ( .A(n3923), .ZN(n3938) );
  MUX2_X1 U2779 ( .A(n2699), .B(n4209), .S(n2728), .Z(n3717) );
  INV_X1 U2780 ( .A(n3625), .ZN(n2175) );
  NAND2_X1 U2781 ( .A1(n2328), .A2(n2326), .ZN(n3897) );
  INV_X1 U2782 ( .A(n2329), .ZN(n2326) );
  NAND2_X1 U2783 ( .A1(n2974), .A2(n2973), .ZN(n3489) );
  NAND2_X1 U2784 ( .A1(n3837), .A2(n2372), .ZN(n2336) );
  INV_X1 U2785 ( .A(n4474), .ZN(n4456) );
  OR2_X1 U2786 ( .A1(n3144), .A2(n3292), .ZN(n3943) );
  INV_X1 U2787 ( .A(n3200), .ZN(n4239) );
  NAND2_X1 U2788 ( .A1(n2851), .A2(n2850), .ZN(n3440) );
  OR2_X1 U2789 ( .A1(n4246), .A2(n2605), .ZN(n2851) );
  NAND2_X1 U2790 ( .A1(n2808), .A2(n2807), .ZN(n4286) );
  NAND2_X1 U2791 ( .A1(n2787), .A2(n2786), .ZN(n4326) );
  OR2_X1 U2792 ( .A1(n4309), .A2(n2605), .ZN(n2787) );
  INV_X1 U2793 ( .A(n4341), .ZN(n3805) );
  NAND2_X1 U2794 ( .A1(n2771), .A2(n2770), .ZN(n4327) );
  INV_X1 U2795 ( .A(n4385), .ZN(n3826) );
  INV_X1 U2796 ( .A(n4437), .ZN(n3910) );
  INV_X1 U2797 ( .A(n4463), .ZN(n4103) );
  INV_X1 U2798 ( .A(n3780), .ZN(n4104) );
  INV_X1 U2799 ( .A(n3467), .ZN(n3703) );
  NAND4_X1 U2800 ( .A1(n2638), .A2(n2637), .A3(n2636), .A4(n2635), .ZN(n4107)
         );
  INV_X1 U2801 ( .A(n2626), .ZN(n4108) );
  OR2_X1 U2802 ( .A1(n2605), .A2(n2582), .ZN(n2583) );
  NAND2_X1 U2803 ( .A1(n3317), .A2(REG2_REG_4__SCAN_IN), .ZN(n3316) );
  XNOR2_X1 U2804 ( .A(n2510), .B(n3314), .ZN(n3304) );
  NAND2_X1 U2805 ( .A1(n3316), .A2(n2408), .ZN(n4135) );
  OAI21_X1 U2806 ( .B1(n3317), .B2(n2352), .A(n2351), .ZN(n4134) );
  INV_X1 U2807 ( .A(n2408), .ZN(n2352) );
  AOI21_X1 U2808 ( .B1(n2408), .B2(n2355), .A(n2354), .ZN(n2351) );
  OAI21_X1 U2809 ( .B1(n3304), .B2(n2274), .A(n2271), .ZN(n4137) );
  INV_X1 U2810 ( .A(n2511), .ZN(n2274) );
  AOI21_X1 U2811 ( .B1(n2511), .B2(n2273), .A(n2272), .ZN(n2271) );
  INV_X1 U2812 ( .A(n4139), .ZN(n2272) );
  NAND2_X1 U2813 ( .A1(n2270), .A2(n2511), .ZN(n4138) );
  NAND2_X1 U2814 ( .A1(n3304), .A2(REG1_REG_4__SCAN_IN), .ZN(n2270) );
  XNOR2_X1 U2815 ( .A(n2415), .B(n3268), .ZN(n3271) );
  NAND2_X1 U2816 ( .A1(n4144), .A2(REG2_REG_8__SCAN_IN), .ZN(n4143) );
  NAND2_X1 U2817 ( .A1(n4143), .A2(n2424), .ZN(n4156) );
  OAI21_X1 U2818 ( .B1(n4144), .B2(n2341), .A(n2340), .ZN(n4154) );
  INV_X1 U2819 ( .A(n2424), .ZN(n2341) );
  AOI21_X1 U2820 ( .B1(n2424), .B2(n2344), .A(n2343), .ZN(n2340) );
  NAND2_X1 U2821 ( .A1(n4161), .A2(n4160), .ZN(n4159) );
  NAND2_X1 U2822 ( .A1(n4149), .A2(n2213), .ZN(n4161) );
  NAND2_X1 U2823 ( .A1(n4170), .A2(n2520), .ZN(n4184) );
  NAND2_X1 U2824 ( .A1(n4179), .A2(n4178), .ZN(n4177) );
  NAND2_X1 U2825 ( .A1(n4166), .A2(n2431), .ZN(n4179) );
  NAND2_X1 U2826 ( .A1(n2202), .A2(n2524), .ZN(n4208) );
  NAND2_X1 U2827 ( .A1(n2362), .A2(n4595), .ZN(n4201) );
  XNOR2_X1 U2828 ( .A(n2526), .B(n4594), .ZN(n3766) );
  NOR2_X1 U2829 ( .A1(n3764), .A2(n4932), .ZN(n3763) );
  AND2_X1 U2830 ( .A1(n2452), .A2(n2449), .ZN(n4622) );
  AND2_X1 U2831 ( .A1(n2495), .A2(n2494), .ZN(n4657) );
  OR2_X1 U2832 ( .A1(n4614), .A2(n3307), .ZN(n4668) );
  NAND2_X1 U2833 ( .A1(n4641), .A2(n2364), .ZN(n4662) );
  AOI21_X1 U2834 ( .B1(n4655), .B2(n4654), .A(n4653), .ZN(n4660) );
  NAND2_X1 U2835 ( .A1(n4644), .A2(n2533), .ZN(n4655) );
  OAI21_X1 U2836 ( .B1(n4633), .B2(n2217), .A(n2215), .ZN(n4652) );
  OR2_X1 U2837 ( .A1(n4614), .A2(n4096), .ZN(n4615) );
  OAI22_X1 U2838 ( .A1(n2215), .A2(n2166), .B1(n4633), .B2(n2139), .ZN(n2537)
         );
  INV_X1 U2839 ( .A(n4653), .ZN(n4648) );
  INV_X1 U2840 ( .A(n4492), .ZN(n4484) );
  AND2_X1 U2841 ( .A1(n3150), .A2(n3110), .ZN(n4226) );
  NAND2_X1 U2842 ( .A1(n4227), .A2(n4351), .ZN(n4228) );
  AND2_X1 U2843 ( .A1(n2137), .A2(n3069), .ZN(n2220) );
  OAI21_X1 U2844 ( .B1(n4386), .B2(n2294), .A(n2292), .ZN(n4321) );
  INV_X1 U2845 ( .A(n2295), .ZN(n4339) );
  AOI21_X1 U2846 ( .B1(n4386), .B2(n2141), .A(n2298), .ZN(n2295) );
  NAND2_X1 U2847 ( .A1(n2282), .A2(n2286), .ZN(n4451) );
  OAI21_X1 U2848 ( .B1(n2714), .B2(n2285), .A(n2283), .ZN(n4449) );
  NAND2_X1 U2849 ( .A1(n2714), .A2(n2143), .ZN(n2282) );
  OR2_X1 U2850 ( .A1(n4459), .A2(n4593), .ZN(n4409) );
  NAND2_X1 U2851 ( .A1(n2820), .A2(n4034), .ZN(n3391) );
  INV_X1 U2852 ( .A(n4461), .ZN(n4674) );
  OR2_X1 U2853 ( .A1(n4409), .A2(n4706), .ZN(n4461) );
  NOR2_X1 U2854 ( .A1(n4459), .A2(n3404), .ZN(n4672) );
  INV_X1 U2855 ( .A(n4669), .ZN(n4447) );
  OR2_X1 U2856 ( .A1(n4498), .A2(n4706), .ZN(n4499) );
  NAND2_X1 U2857 ( .A1(n4497), .A2(n4545), .ZN(n4501) );
  NAND2_X1 U2858 ( .A1(n3253), .A2(n3252), .ZN(n4678) );
  AND2_X1 U2859 ( .A1(n3136), .A2(STATE_REG_SCAN_IN), .ZN(n4726) );
  INV_X1 U2860 ( .A(n4094), .ZN(n4593) );
  INV_X1 U2861 ( .A(n2535), .ZN(n4679) );
  INV_X1 U2862 ( .A(n2559), .ZN(n2409) );
  AND2_X1 U2863 ( .A1(n2404), .A2(n2401), .ZN(n4603) );
  NAND3_X1 U2864 ( .A1(n2306), .A2(IR_REG_31__SCAN_IN), .A3(IR_REG_0__SCAN_IN), 
        .ZN(n2276) );
  NAND2_X1 U2865 ( .A1(n4685), .A2(IR_REG_1__SCAN_IN), .ZN(n2275) );
  AND2_X1 U2866 ( .A1(n3171), .A2(n3170), .ZN(n3172) );
  NOR2_X1 U2867 ( .A1(n4725), .A2(REG1_REG_29__SCAN_IN), .ZN(n2311) );
  AND3_X1 U2868 ( .A1(n4494), .A2(n4495), .A3(n4725), .ZN(n2309) );
  AND2_X1 U2869 ( .A1(n4551), .A2(n4552), .ZN(n2233) );
  NOR2_X1 U2870 ( .A1(n4717), .A2(REG0_REG_29__SCAN_IN), .ZN(n2312) );
  AND3_X1 U2871 ( .A1(n4494), .A2(n4495), .A3(n4717), .ZN(n2310) );
  NAND2_X1 U2872 ( .A1(n2267), .A2(n2266), .ZN(U3513) );
  OR2_X1 U2873 ( .A1(n4717), .A2(n4807), .ZN(n2266) );
  NAND2_X1 U2874 ( .A1(n4559), .A2(n4717), .ZN(n2267) );
  OR2_X1 U2875 ( .A1(n4505), .A2(n4586), .ZN(n2886) );
  AND2_X1 U2876 ( .A1(n2152), .A2(n3097), .ZN(n2130) );
  AND2_X1 U2877 ( .A1(n2130), .A2(n3079), .ZN(n2131) );
  INV_X4 U2878 ( .A(n2590), .ZN(n2591) );
  AND2_X1 U2879 ( .A1(n2259), .A2(n3464), .ZN(n2132) );
  NAND2_X1 U2880 ( .A1(n4436), .A2(n4456), .ZN(n2133) );
  INV_X1 U2881 ( .A(n3538), .ZN(n3542) );
  NAND2_X1 U2882 ( .A1(n2617), .A2(n2616), .ZN(n3538) );
  INV_X1 U2883 ( .A(n2372), .ZN(n2173) );
  AND2_X1 U2884 ( .A1(n2437), .A2(n2161), .ZN(n2134) );
  NAND2_X1 U2885 ( .A1(n4389), .A2(n2221), .ZN(n2222) );
  AND2_X1 U2886 ( .A1(n2130), .A2(n2173), .ZN(n2135) );
  AND2_X1 U2887 ( .A1(n3234), .A2(n2479), .ZN(n2136) );
  NAND2_X1 U2888 ( .A1(n3614), .A2(n3660), .ZN(n3659) );
  AOI21_X1 U2889 ( .B1(n2265), .B2(n4046), .A(n2264), .ZN(n2263) );
  AND2_X1 U2890 ( .A1(n2221), .A2(n2882), .ZN(n2137) );
  OR2_X1 U2891 ( .A1(n4595), .A2(REG2_REG_13__SCAN_IN), .ZN(n2138) );
  OR2_X1 U2892 ( .A1(n2217), .A2(n2166), .ZN(n2139) );
  AND2_X1 U2893 ( .A1(n4598), .A2(REG1_REG_9__SCAN_IN), .ZN(n2140) );
  NAND2_X1 U2894 ( .A1(n4289), .A2(n4290), .ZN(n4270) );
  AND2_X1 U2895 ( .A1(n2303), .A2(n2757), .ZN(n2141) );
  NAND2_X1 U2896 ( .A1(n2526), .A2(n4594), .ZN(n2142) );
  AND2_X1 U2897 ( .A1(n2133), .A2(n2713), .ZN(n2143) );
  NAND2_X1 U2898 ( .A1(n3581), .A2(n3554), .ZN(n4044) );
  NAND2_X1 U2899 ( .A1(n2328), .A2(n2327), .ZN(n3799) );
  AND2_X1 U2900 ( .A1(n3782), .A2(n4474), .ZN(n2144) );
  AOI21_X1 U2901 ( .B1(n3852), .B2(n3026), .A(n3025), .ZN(n3863) );
  NAND2_X1 U2902 ( .A1(n2181), .A2(n2192), .ZN(n3906) );
  INV_X1 U2903 ( .A(n2829), .ZN(n3989) );
  NAND2_X1 U2904 ( .A1(n3951), .A2(n3947), .ZN(n2829) );
  AND2_X1 U2905 ( .A1(n4416), .A2(n2727), .ZN(n2145) );
  INV_X1 U2906 ( .A(IR_REG_6__SCAN_IN), .ZN(n2386) );
  AOI21_X1 U2907 ( .B1(n3811), .B2(n3059), .A(n3058), .ZN(n3821) );
  INV_X1 U2908 ( .A(n4241), .ZN(n3190) );
  AND3_X1 U2909 ( .A1(n3128), .A2(n3131), .A3(n3888), .ZN(n2146) );
  NOR2_X1 U2910 ( .A1(n3763), .A2(n2446), .ZN(n2147) );
  INV_X1 U2911 ( .A(n4037), .ZN(n2244) );
  AND2_X1 U2912 ( .A1(n4385), .A2(n4369), .ZN(n2148) );
  NAND2_X1 U2913 ( .A1(n4289), .A2(n2223), .ZN(n2227) );
  INV_X1 U2914 ( .A(n3652), .ZN(n3660) );
  MUX2_X1 U2915 ( .A(DATAI_12_), .B(n4596), .S(n2728), .Z(n3652) );
  NOR2_X1 U2916 ( .A1(n4265), .A2(n4290), .ZN(n2149) );
  AND2_X1 U2917 ( .A1(n2154), .A2(n3163), .ZN(n2150) );
  INV_X1 U2918 ( .A(n2263), .ZN(n2262) );
  AND2_X1 U2919 ( .A1(n3440), .A2(n3189), .ZN(n2151) );
  INV_X1 U2920 ( .A(IR_REG_26__SCAN_IN), .ZN(n2556) );
  NAND2_X1 U2921 ( .A1(n3103), .A2(n3102), .ZN(n2152) );
  AND2_X1 U2922 ( .A1(n4327), .A2(n3829), .ZN(n2153) );
  INV_X1 U2923 ( .A(IR_REG_2__SCAN_IN), .ZN(n2359) );
  AND2_X1 U2924 ( .A1(n2152), .A2(n2335), .ZN(n2154) );
  OR2_X1 U2925 ( .A1(n2371), .A2(n2148), .ZN(n2155) );
  INV_X1 U2926 ( .A(n2299), .ZN(n2298) );
  NAND2_X1 U2927 ( .A1(n2155), .A2(n2303), .ZN(n2299) );
  AND2_X1 U2928 ( .A1(n4311), .A2(n4313), .ZN(n4289) );
  INV_X1 U2929 ( .A(n3580), .ZN(n3581) );
  OAI21_X1 U2930 ( .B1(n2612), .B2(n2631), .A(n2630), .ZN(n3580) );
  AND2_X1 U2931 ( .A1(n2301), .A2(n2300), .ZN(n2156) );
  AND2_X1 U2932 ( .A1(n2469), .A2(n2556), .ZN(n2157) );
  AND2_X1 U2933 ( .A1(n2192), .A2(n2191), .ZN(n2158) );
  AND2_X1 U2934 ( .A1(n2219), .A2(n2142), .ZN(n2159) );
  INV_X1 U2935 ( .A(n3532), .ZN(n2247) );
  INV_X1 U2936 ( .A(n3945), .ZN(n3888) );
  AND2_X1 U2937 ( .A1(n2852), .A2(n4023), .ZN(n2885) );
  NAND2_X1 U2938 ( .A1(n2979), .A2(n2980), .ZN(n3479) );
  AND2_X1 U2939 ( .A1(n2604), .A2(n2603), .ZN(n3393) );
  BUF_X1 U2940 ( .A(n2816), .Z(n2884) );
  NAND2_X1 U2941 ( .A1(n2176), .A2(n2989), .ZN(n3623) );
  NAND2_X1 U2942 ( .A1(n2177), .A2(n3624), .ZN(n3710) );
  NAND2_X1 U2943 ( .A1(n2308), .A2(n2307), .ZN(n3776) );
  AND2_X1 U2944 ( .A1(n2714), .A2(n2713), .ZN(n2160) );
  AND2_X1 U2945 ( .A1(n4389), .A2(n2220), .ZN(n4311) );
  NAND2_X1 U2946 ( .A1(n2385), .A2(n2560), .ZN(n2460) );
  OR2_X1 U2947 ( .A1(n4209), .A2(n2441), .ZN(n2161) );
  NAND2_X1 U2948 ( .A1(n3064), .A2(n3065), .ZN(n2162) );
  NAND2_X1 U2949 ( .A1(n4389), .A2(n4388), .ZN(n4368) );
  INV_X1 U2950 ( .A(n4369), .ZN(n4360) );
  NAND2_X1 U2951 ( .A1(n3968), .A2(DATAI_20_), .ZN(n4369) );
  INV_X1 U2952 ( .A(IR_REG_15__SCAN_IN), .ZN(n2447) );
  NOR2_X1 U2953 ( .A1(n3399), .A2(n2229), .ZN(n3430) );
  NAND2_X1 U2954 ( .A1(n3430), .A2(n3557), .ZN(n3431) );
  INV_X1 U2955 ( .A(n3189), .ZN(n4243) );
  NAND2_X1 U2956 ( .A1(n3335), .A2(n2914), .ZN(n3365) );
  AND2_X1 U2957 ( .A1(n3613), .A2(n2977), .ZN(n3614) );
  NAND2_X1 U2958 ( .A1(n2304), .A2(n2920), .ZN(n3372) );
  OR2_X1 U2959 ( .A1(n3399), .A2(n3542), .ZN(n2163) );
  INV_X1 U2960 ( .A(n3174), .ZN(n3928) );
  NAND2_X1 U2961 ( .A1(n3968), .A2(DATAI_26_), .ZN(n3174) );
  AND2_X1 U2962 ( .A1(n2364), .A2(n2363), .ZN(n2164) );
  AND2_X1 U2963 ( .A1(n2533), .A2(n2534), .ZN(n2165) );
  AND2_X1 U2964 ( .A1(n2612), .A2(DATAI_22_), .ZN(n4332) );
  AND2_X1 U2965 ( .A1(n2535), .A2(REG1_REG_18__SCAN_IN), .ZN(n2166) );
  INV_X1 U2966 ( .A(REG1_REG_8__SCAN_IN), .ZN(n2210) );
  INV_X1 U2967 ( .A(REG2_REG_8__SCAN_IN), .ZN(n2344) );
  INV_X1 U2968 ( .A(REG1_REG_4__SCAN_IN), .ZN(n2273) );
  XNOR2_X1 U2969 ( .A(n2953), .B(n3117), .ZN(n2962) );
  NAND2_X2 U2970 ( .A1(n2565), .A2(n4590), .ZN(n2605) );
  XNOR2_X2 U2971 ( .A(n2170), .B(IR_REG_30__SCAN_IN), .ZN(n2565) );
  OR2_X2 U2972 ( .A1(n3772), .A2(n2360), .ZN(n2170) );
  OR2_X2 U2973 ( .A1(n3852), .A2(n2195), .ZN(n2181) );
  NAND2_X2 U2974 ( .A1(n3799), .A2(n3079), .ZN(n3837) );
  NAND3_X1 U2975 ( .A1(n2974), .A2(n2973), .A3(n2172), .ZN(n2171) );
  NAND2_X1 U2976 ( .A1(n2910), .A2(n2911), .ZN(n3335) );
  INV_X1 U2977 ( .A(n2174), .ZN(n3165) );
  NAND3_X1 U2978 ( .A1(n2176), .A2(n2989), .A3(n2175), .ZN(n2177) );
  NAND2_X1 U2979 ( .A1(n3407), .A2(n2179), .ZN(n2178) );
  NAND2_X1 U2980 ( .A1(n3407), .A2(n2937), .ZN(n3418) );
  NAND2_X2 U2981 ( .A1(n3409), .A2(n3408), .ZN(n3407) );
  NAND4_X1 U2982 ( .A1(n2187), .A2(n2186), .A3(n2184), .A4(n3847), .ZN(U3222)
         );
  NAND3_X1 U2983 ( .A1(n2190), .A2(n2189), .A3(n2185), .ZN(n2184) );
  AND2_X1 U2984 ( .A1(n3726), .A2(n3549), .ZN(n2985) );
  NAND3_X1 U2985 ( .A1(n2560), .A2(n2468), .A3(n2559), .ZN(n2471) );
  OAI211_X1 U2986 ( .C1(n4194), .C2(REG1_REG_12__SCAN_IN), .A(n2202), .B(n4648), .ZN(n4197) );
  INV_X1 U2987 ( .A(n2520), .ZN(n2207) );
  INV_X1 U2988 ( .A(n2214), .ZN(n2213) );
  INV_X1 U2989 ( .A(n2219), .ZN(n3765) );
  INV_X1 U2990 ( .A(n2222), .ZN(n4346) );
  INV_X1 U2991 ( .A(n2227), .ZN(n4244) );
  NAND3_X1 U2992 ( .A1(n2880), .A2(n3538), .A3(n3580), .ZN(n2229) );
  NOR2_X2 U2993 ( .A1(n3455), .A2(n3296), .ZN(n3354) );
  NAND4_X1 U2994 ( .A1(n2560), .A2(n2468), .A3(n2157), .A4(n2559), .ZN(n2230)
         );
  NAND2_X1 U2995 ( .A1(n2489), .A2(n2555), .ZN(n2231) );
  XNOR2_X1 U2996 ( .A(n4221), .B(n4216), .ZN(n4553) );
  OAI21_X1 U2997 ( .B1(n4553), .B2(n4586), .A(n2233), .ZN(U3517) );
  NAND2_X1 U2998 ( .A1(n2818), .A2(n2234), .ZN(n3453) );
  INV_X1 U2999 ( .A(n3452), .ZN(n2234) );
  INV_X1 U3000 ( .A(n2817), .ZN(n2818) );
  XNOR2_X1 U3001 ( .A(n2817), .B(n3454), .ZN(n3459) );
  NOR2_X1 U3002 ( .A1(n3995), .A2(n2817), .ZN(n2236) );
  OAI21_X1 U3003 ( .B1(n2828), .B2(n2829), .A(n2238), .ZN(n4470) );
  INV_X1 U3004 ( .A(n4235), .ZN(n3191) );
  NAND2_X1 U3005 ( .A1(n2254), .A2(n2255), .ZN(n3521) );
  NAND3_X1 U3006 ( .A1(n4499), .A2(n4500), .A3(n4501), .ZN(n4559) );
  NAND2_X1 U3007 ( .A1(n2360), .A2(IR_REG_1__SCAN_IN), .ZN(n2277) );
  NAND2_X1 U3008 ( .A1(n2714), .A2(n2283), .ZN(n2281) );
  NAND2_X1 U3009 ( .A1(n2650), .A2(n3381), .ZN(n2653) );
  NAND2_X1 U3010 ( .A1(n2287), .A2(n2629), .ZN(n3381) );
  NAND4_X1 U3011 ( .A1(n2604), .A2(n2628), .A3(n3390), .A4(n2603), .ZN(n2287)
         );
  NAND3_X1 U3012 ( .A1(n2304), .A2(n2920), .A3(n2926), .ZN(n3374) );
  NOR2_X2 U3013 ( .A1(n2398), .A2(n2377), .ZN(n2559) );
  NAND3_X1 U3014 ( .A1(n2306), .A2(n2305), .A3(n2359), .ZN(n2398) );
  AOI21_X1 U3015 ( .B1(n2309), .B2(n4496), .A(n2311), .ZN(U3547) );
  AOI21_X1 U3016 ( .B1(n2310), .B2(n4496), .A(n2312), .ZN(U3515) );
  NAND2_X1 U3017 ( .A1(n2809), .A2(n2315), .ZN(n2314) );
  NAND2_X1 U3018 ( .A1(n2809), .A2(n2373), .ZN(n2321) );
  NAND2_X1 U3019 ( .A1(n2336), .A2(n3097), .ZN(n3916) );
  OAI21_X1 U3020 ( .B1(n2431), .B2(n2347), .A(n2433), .ZN(n2346) );
  XNOR2_X1 U3021 ( .A(n2436), .B(n4195), .ZN(n4191) );
  INV_X1 U3022 ( .A(n2349), .ZN(n2348) );
  INV_X1 U3023 ( .A(IR_REG_31__SCAN_IN), .ZN(n2360) );
  NAND2_X1 U3024 ( .A1(n4642), .A2(n4643), .ZN(n4641) );
  INV_X1 U3025 ( .A(n2459), .ZN(n4661) );
  NAND2_X1 U3026 ( .A1(n2446), .A2(n2367), .ZN(n2365) );
  XNOR2_X1 U3027 ( .A(n2901), .B(n2903), .ZN(n3795) );
  XNOR2_X1 U3028 ( .A(n2900), .B(n2128), .ZN(n2903) );
  NAND2_X1 U3029 ( .A1(n4630), .A2(n2456), .ZN(n4642) );
  NAND2_X1 U3030 ( .A1(n4167), .A2(REG2_REG_10__SCAN_IN), .ZN(n4166) );
  INV_X1 U3031 ( .A(n3710), .ZN(n3004) );
  NAND2_X1 U3032 ( .A1(n4191), .A2(REG2_REG_12__SCAN_IN), .ZN(n4190) );
  INV_X1 U3033 ( .A(n2565), .ZN(n2566) );
  AND2_X2 U3034 ( .A1(n2565), .A2(n2564), .ZN(n2621) );
  OAI22_X2 U3035 ( .A1(n3528), .A2(n2679), .B1(n3701), .B2(n2881), .ZN(n3608)
         );
  AND2_X1 U3036 ( .A1(n3160), .A2(n3159), .ZN(n2368) );
  AND2_X2 U3037 ( .A1(n3228), .A2(n3183), .ZN(n4717) );
  INV_X1 U3038 ( .A(n4725), .ZN(n3232) );
  OR2_X1 U3039 ( .A1(n3971), .A2(n4464), .ZN(n2369) );
  INV_X1 U3040 ( .A(n4600), .ZN(n2631) );
  XOR2_X1 U3041 ( .A(n3179), .B(n4484), .Z(n2370) );
  AND2_X1 U3042 ( .A1(n2833), .A2(n4388), .ZN(n2371) );
  INV_X1 U3043 ( .A(IR_REG_24__SCAN_IN), .ZN(n2859) );
  AND2_X1 U3044 ( .A1(n3838), .A2(n3091), .ZN(n2372) );
  OR2_X1 U3045 ( .A1(n4286), .A2(n3843), .ZN(n2373) );
  AND2_X2 U3046 ( .A1(n3184), .A2(n4447), .ZN(n4459) );
  INV_X1 U3047 ( .A(n4459), .ZN(n4316) );
  NOR2_X1 U3048 ( .A1(n4230), .A2(n4586), .ZN(n2374) );
  NAND2_X1 U3049 ( .A1(n2819), .A2(n4029), .ZN(n3346) );
  NAND2_X1 U3050 ( .A1(n2627), .A2(n3539), .ZN(n2375) );
  AND2_X1 U3051 ( .A1(n2612), .A2(DATAI_21_), .ZN(n3829) );
  INV_X1 U3052 ( .A(n3735), .ZN(n2881) );
  OR2_X1 U3053 ( .A1(n4326), .A2(n3070), .ZN(n2376) );
  XNOR2_X1 U3054 ( .A(n2454), .B(n2453), .ZN(n4682) );
  INV_X1 U3055 ( .A(n4682), .ZN(n2529) );
  XNOR2_X1 U3056 ( .A(n2392), .B(n2391), .ZN(n2729) );
  INV_X1 U3057 ( .A(n3588), .ZN(n2880) );
  AND2_X2 U3058 ( .A1(n3185), .A2(n2888), .ZN(n2898) );
  INV_X1 U3059 ( .A(n2498), .ZN(n2587) );
  INV_X1 U3060 ( .A(n4469), .ZN(n2830) );
  INV_X1 U3061 ( .A(n3711), .ZN(n3003) );
  INV_X1 U3062 ( .A(n3777), .ZN(n3008) );
  AND2_X1 U3063 ( .A1(n4622), .A2(REG1_REG_15__SCAN_IN), .ZN(n2528) );
  INV_X1 U3064 ( .A(n2729), .ZN(n2532) );
  INV_X1 U3065 ( .A(n4435), .ZN(n2727) );
  INV_X1 U3066 ( .A(REG3_REG_12__SCAN_IN), .ZN(n2692) );
  NAND2_X1 U3067 ( .A1(n2831), .A2(n2830), .ZN(n4466) );
  AND2_X1 U3068 ( .A1(n2864), .A2(n3125), .ZN(n3138) );
  INV_X1 U3069 ( .A(IR_REG_25__SCAN_IN), .ZN(n2469) );
  INV_X1 U3070 ( .A(n3223), .ZN(n3217) );
  INV_X1 U3071 ( .A(REG3_REG_8__SCAN_IN), .ZN(n4730) );
  INV_X1 U3072 ( .A(REG3_REG_25__SCAN_IN), .ZN(n4988) );
  AND2_X1 U3073 ( .A1(REG3_REG_15__SCAN_IN), .A2(REG3_REG_14__SCAN_IN), .ZN(
        n2545) );
  NAND2_X1 U3074 ( .A1(n2552), .A2(REG3_REG_24__SCAN_IN), .ZN(n2800) );
  INV_X1 U3075 ( .A(REG3_REG_13__SCAN_IN), .ZN(n4999) );
  AND2_X1 U3076 ( .A1(n2445), .A2(n4594), .ZN(n2446) );
  NAND2_X1 U3077 ( .A1(n2553), .A2(REG3_REG_26__SCAN_IN), .ZN(n2845) );
  AND2_X1 U3078 ( .A1(n3910), .A2(n4427), .ZN(n2735) );
  INV_X1 U3079 ( .A(n4405), .ZN(n4397) );
  INV_X1 U3080 ( .A(n3390), .ZN(n4006) );
  AND2_X1 U3081 ( .A1(n3968), .A2(DATAI_27_), .ZN(n3189) );
  INV_X1 U3082 ( .A(REG3_REG_23__SCAN_IN), .ZN(n4792) );
  NAND2_X1 U3083 ( .A1(n2546), .A2(n2545), .ZN(n2720) );
  OR2_X1 U3084 ( .A1(n3697), .A2(n3696), .ZN(n3727) );
  OR3_X1 U3085 ( .A1(n3156), .A2(n3307), .A3(n4097), .ZN(n3923) );
  OR2_X1 U3086 ( .A1(n3109), .A2(n3149), .ZN(n3150) );
  XNOR2_X1 U3087 ( .A(n2498), .B(n2396), .ZN(n3324) );
  AOI21_X1 U3088 ( .B1(n4657), .B2(ADDR_REG_18__SCAN_IN), .A(n4656), .ZN(n4658) );
  INV_X1 U3089 ( .A(n4327), .ZN(n4362) );
  AND2_X1 U3090 ( .A1(n2734), .A2(n2733), .ZN(n4437) );
  OR2_X1 U3091 ( .A1(n3253), .A2(D_REG_1__SCAN_IN), .ZN(n3181) );
  NOR2_X1 U3092 ( .A1(n4693), .A2(n4591), .ZN(n3147) );
  INV_X1 U3093 ( .A(n4111), .ZN(n3790) );
  OR2_X1 U3094 ( .A1(n3253), .A2(D_REG_0__SCAN_IN), .ZN(n2879) );
  AND2_X1 U3095 ( .A1(n3219), .A2(n2369), .ZN(n3220) );
  INV_X1 U3096 ( .A(n3829), .ZN(n2882) );
  INV_X1 U3097 ( .A(n3717), .ZN(n3686) );
  NAND2_X1 U3098 ( .A1(n2885), .A2(n4592), .ZN(n4422) );
  NAND2_X1 U3099 ( .A1(n3125), .A2(n4606), .ZN(n4464) );
  NAND2_X1 U3100 ( .A1(n2888), .A2(n4726), .ZN(n3146) );
  NAND2_X1 U3101 ( .A1(n2547), .A2(REG3_REG_16__SCAN_IN), .ZN(n2739) );
  NAND2_X1 U3102 ( .A1(n2746), .A2(n2745), .ZN(n4419) );
  XNOR2_X1 U3103 ( .A(n2519), .B(n4172), .ZN(n4171) );
  INV_X1 U3104 ( .A(n4615), .ZN(n4664) );
  INV_X1 U3105 ( .A(n4464), .ZN(n4418) );
  INV_X1 U3106 ( .A(n4422), .ZN(n4473) );
  INV_X1 U3107 ( .A(n4452), .ZN(n4477) );
  AND2_X1 U3108 ( .A1(n3252), .A2(n3147), .ZN(n4669) );
  INV_X1 U3109 ( .A(n4540), .ZN(n4481) );
  AND2_X1 U3110 ( .A1(n2879), .A2(n3254), .ZN(n3227) );
  NOR2_X1 U3111 ( .A1(n4717), .A2(n4810), .ZN(n3225) );
  INV_X1 U3112 ( .A(n4545), .ZN(n4710) );
  INV_X1 U3113 ( .A(n4586), .ZN(n4554) );
  AND2_X2 U3114 ( .A1(n2885), .A2(n2884), .ZN(n4698) );
  INV_X1 U3115 ( .A(n3227), .ZN(n3183) );
  INV_X1 U3116 ( .A(n3146), .ZN(n3252) );
  INV_X1 U3117 ( .A(n2863), .ZN(n3234) );
  INV_X1 U3118 ( .A(n3943), .ZN(n3922) );
  OR2_X1 U3119 ( .A1(n3145), .A2(n3134), .ZN(n3945) );
  INV_X1 U3120 ( .A(U4043), .ZN(n3439) );
  INV_X1 U3121 ( .A(n4234), .ZN(n4267) );
  NAND2_X1 U3122 ( .A1(n2756), .A2(n2755), .ZN(n4398) );
  INV_X1 U3123 ( .A(n3439), .ZN(n4109) );
  OR2_X1 U3124 ( .A1(n4614), .A2(n4611), .ZN(n4653) );
  AOI21_X1 U3125 ( .B1(n4652), .B2(n4660), .A(n4659), .ZN(n4667) );
  INV_X1 U3126 ( .A(n2497), .ZN(n2540) );
  OR2_X1 U3127 ( .A1(n4459), .A2(n3186), .ZN(n4452) );
  AND2_X1 U3128 ( .A1(n4026), .A2(n3454), .ZN(n4007) );
  NAND2_X1 U3129 ( .A1(n4725), .A2(n4698), .ZN(n4540) );
  AND2_X2 U3130 ( .A1(n3228), .A2(n3227), .ZN(n4725) );
  AND2_X1 U3131 ( .A1(n4220), .A2(n4219), .ZN(n4558) );
  NAND2_X1 U3132 ( .A1(n4717), .A2(n4698), .ZN(n4586) );
  INV_X1 U3133 ( .A(n4717), .ZN(n4716) );
  INV_X1 U3134 ( .A(n4678), .ZN(n4729) );
  INV_X1 U3135 ( .A(n4023), .ZN(n4591) );
  AND2_X2 U3136 ( .A1(n3299), .A2(n4726), .ZN(U4043) );
  OAI211_X1 U3137 ( .C1(n2370), .C2(n4452), .A(n3211), .B(n3210), .ZN(U3354)
         );
  OAI21_X1 U3138 ( .B1(n3233), .B2(n3232), .A(n3231), .ZN(U3546) );
  OAI21_X1 U3139 ( .B1(n3233), .B2(n4716), .A(n3226), .ZN(U3514) );
  NAND2_X1 U3140 ( .A1(n2399), .A2(n2405), .ZN(n2377) );
  AND2_X2 U3141 ( .A1(n2559), .A2(n2410), .ZN(n2385) );
  NOR2_X2 U3142 ( .A1(IR_REG_13__SCAN_IN), .A2(IR_REG_11__SCAN_IN), .ZN(n2388)
         );
  AND2_X1 U3143 ( .A1(n2388), .A2(n2378), .ZN(n2383) );
  NOR2_X1 U3144 ( .A1(IR_REG_14__SCAN_IN), .A2(IR_REG_9__SCAN_IN), .ZN(n2380)
         );
  NOR2_X1 U3145 ( .A1(IR_REG_7__SCAN_IN), .A2(IR_REG_17__SCAN_IN), .ZN(n2379)
         );
  AND2_X1 U3146 ( .A1(n2380), .A2(n2379), .ZN(n2381) );
  AND3_X2 U3147 ( .A1(n2383), .A2(n2382), .A3(n2381), .ZN(n2560) );
  NAND2_X1 U31480 ( .A1(n2460), .A2(IR_REG_31__SCAN_IN), .ZN(n2384) );
  XNOR2_X1 U31490 ( .A(n2384), .B(IR_REG_18__SCAN_IN), .ZN(n2535) );
  NAND2_X1 U3150 ( .A1(REG2_REG_18__SCAN_IN), .A2(n2535), .ZN(n2458) );
  OAI21_X1 U3151 ( .B1(REG2_REG_18__SCAN_IN), .B2(n2535), .A(n2458), .ZN(n4663) );
  NAND2_X1 U3152 ( .A1(n2385), .A2(n2386), .ZN(n2417) );
  NAND2_X1 U3153 ( .A1(n2428), .A2(n2387), .ZN(n2432) );
  NAND2_X1 U3154 ( .A1(n2388), .A2(n4778), .ZN(n2389) );
  OAI21_X1 U3155 ( .B1(IR_REG_15__SCAN_IN), .B2(IR_REG_16__SCAN_IN), .A(
        IR_REG_31__SCAN_IN), .ZN(n2390) );
  NAND2_X1 U3156 ( .A1(n2448), .A2(n2390), .ZN(n2392) );
  INV_X1 U3157 ( .A(REG2_REG_1__SCAN_IN), .ZN(n2393) );
  XNOR2_X1 U3158 ( .A(n2501), .B(n2393), .ZN(n4114) );
  INV_X1 U3159 ( .A(IR_REG_0__SCAN_IN), .ZN(n4685) );
  NAND2_X1 U3160 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n3309) );
  INV_X1 U3161 ( .A(n3309), .ZN(n4113) );
  NAND2_X1 U3162 ( .A1(n4114), .A2(n4113), .ZN(n4112) );
  NAND2_X1 U3163 ( .A1(n2127), .A2(REG2_REG_1__SCAN_IN), .ZN(n2394) );
  NAND2_X1 U3164 ( .A1(n4112), .A2(n2394), .ZN(n3323) );
  INV_X1 U3165 ( .A(REG2_REG_2__SCAN_IN), .ZN(n2396) );
  NAND2_X1 U3166 ( .A1(n3323), .A2(n3324), .ZN(n3322) );
  NAND2_X1 U3167 ( .A1(n2498), .A2(REG2_REG_2__SCAN_IN), .ZN(n2397) );
  NAND2_X1 U3168 ( .A1(n2398), .A2(IR_REG_31__SCAN_IN), .ZN(n2400) );
  NAND2_X1 U3169 ( .A1(n2400), .A2(n2399), .ZN(n2404) );
  OR2_X1 U3170 ( .A1(n2400), .A2(n2399), .ZN(n2401) );
  NAND2_X1 U3171 ( .A1(n4124), .A2(REG2_REG_3__SCAN_IN), .ZN(n4123) );
  NAND2_X1 U3172 ( .A1(n2402), .A2(n4603), .ZN(n2403) );
  NAND2_X1 U3173 ( .A1(n2404), .A2(IR_REG_31__SCAN_IN), .ZN(n2406) );
  XNOR2_X1 U3174 ( .A(n2406), .B(n2405), .ZN(n3314) );
  INV_X1 U3175 ( .A(n3314), .ZN(n4602) );
  NAND2_X1 U3176 ( .A1(n2407), .A2(n4602), .ZN(n2408) );
  NAND2_X1 U3177 ( .A1(n2409), .A2(IR_REG_31__SCAN_IN), .ZN(n2411) );
  INV_X1 U3178 ( .A(IR_REG_5__SCAN_IN), .ZN(n2410) );
  XNOR2_X1 U3179 ( .A(n2411), .B(n2410), .ZN(n4131) );
  XNOR2_X1 U3180 ( .A(n4131), .B(REG2_REG_5__SCAN_IN), .ZN(n4136) );
  INV_X1 U3181 ( .A(REG2_REG_5__SCAN_IN), .ZN(n2412) );
  OR2_X1 U3182 ( .A1(n4131), .A2(n2412), .ZN(n2413) );
  OR2_X1 U3183 ( .A1(n2385), .A2(n2360), .ZN(n2414) );
  XNOR2_X1 U3184 ( .A(n2414), .B(IR_REG_6__SCAN_IN), .ZN(n4601) );
  INV_X1 U3185 ( .A(n4601), .ZN(n3268) );
  NAND2_X1 U3186 ( .A1(n3271), .A2(REG2_REG_6__SCAN_IN), .ZN(n3270) );
  NAND2_X1 U3187 ( .A1(n2415), .A2(n4601), .ZN(n2416) );
  NAND2_X1 U3188 ( .A1(n3270), .A2(n2416), .ZN(n3280) );
  INV_X1 U3189 ( .A(REG2_REG_7__SCAN_IN), .ZN(n3587) );
  NAND2_X1 U3190 ( .A1(n2417), .A2(IR_REG_31__SCAN_IN), .ZN(n2419) );
  XNOR2_X1 U3191 ( .A(n2419), .B(n4962), .ZN(n4600) );
  MUX2_X1 U3192 ( .A(n3587), .B(REG2_REG_7__SCAN_IN), .S(n4600), .Z(n3279) );
  NAND2_X1 U3193 ( .A1(n3280), .A2(n3279), .ZN(n3278) );
  OR2_X1 U3194 ( .A1(n4600), .A2(n3587), .ZN(n2418) );
  NAND2_X1 U3195 ( .A1(n2419), .A2(n4962), .ZN(n2420) );
  NAND2_X1 U3196 ( .A1(n2420), .A2(IR_REG_31__SCAN_IN), .ZN(n2422) );
  INV_X1 U3197 ( .A(IR_REG_8__SCAN_IN), .ZN(n2421) );
  XNOR2_X1 U3198 ( .A(n2422), .B(n2421), .ZN(n4146) );
  INV_X1 U3199 ( .A(n4146), .ZN(n4599) );
  NAND2_X1 U3200 ( .A1(n2423), .A2(n4599), .ZN(n2424) );
  INV_X1 U3201 ( .A(REG2_REG_9__SCAN_IN), .ZN(n4931) );
  NAND2_X1 U3202 ( .A1(n2425), .A2(IR_REG_31__SCAN_IN), .ZN(n2426) );
  XNOR2_X1 U3203 ( .A(n2426), .B(IR_REG_9__SCAN_IN), .ZN(n4598) );
  MUX2_X1 U3204 ( .A(REG2_REG_9__SCAN_IN), .B(n4931), .S(n4598), .Z(n4155) );
  NAND2_X1 U3205 ( .A1(n4598), .A2(REG2_REG_9__SCAN_IN), .ZN(n2427) );
  OR2_X1 U3206 ( .A1(n2428), .A2(n2360), .ZN(n2429) );
  XNOR2_X1 U3207 ( .A(n2429), .B(IR_REG_10__SCAN_IN), .ZN(n4597) );
  INV_X1 U3208 ( .A(n4597), .ZN(n4172) );
  NAND2_X1 U3209 ( .A1(n2430), .A2(n4597), .ZN(n2431) );
  XNOR2_X1 U32100 ( .A(n2434), .B(n4767), .ZN(n4185) );
  XNOR2_X1 U32110 ( .A(n4185), .B(REG2_REG_11__SCAN_IN), .ZN(n4178) );
  INV_X1 U32120 ( .A(REG2_REG_11__SCAN_IN), .ZN(n3618) );
  OR2_X1 U32130 ( .A1(n4185), .A2(n3618), .ZN(n2433) );
  NAND2_X1 U32140 ( .A1(n2434), .A2(n4767), .ZN(n2438) );
  NAND2_X1 U32150 ( .A1(n2438), .A2(IR_REG_31__SCAN_IN), .ZN(n2435) );
  XNOR2_X1 U32160 ( .A(n2435), .B(IR_REG_12__SCAN_IN), .ZN(n4596) );
  INV_X1 U32170 ( .A(n4596), .ZN(n4195) );
  NAND2_X1 U32180 ( .A1(n2436), .A2(n4596), .ZN(n2437) );
  INV_X1 U32190 ( .A(IR_REG_13__SCAN_IN), .ZN(n2439) );
  XNOR2_X1 U32200 ( .A(n2440), .B(n2439), .ZN(n4209) );
  INV_X1 U32210 ( .A(n4209), .ZN(n4595) );
  INV_X1 U32220 ( .A(REG2_REG_13__SCAN_IN), .ZN(n2441) );
  NAND2_X1 U32230 ( .A1(n2442), .A2(IR_REG_31__SCAN_IN), .ZN(n2443) );
  XNOR2_X1 U32240 ( .A(n2443), .B(IR_REG_14__SCAN_IN), .ZN(n4594) );
  INV_X1 U32250 ( .A(n4594), .ZN(n3768) );
  INV_X1 U32260 ( .A(REG2_REG_14__SCAN_IN), .ZN(n4932) );
  INV_X1 U32270 ( .A(n2444), .ZN(n2445) );
  NAND2_X1 U32280 ( .A1(n2448), .A2(n2447), .ZN(n2452) );
  OR2_X1 U32290 ( .A1(n2448), .A2(n2447), .ZN(n2449) );
  INV_X1 U32300 ( .A(n4622), .ZN(n4684) );
  INV_X1 U32310 ( .A(REG2_REG_15__SCAN_IN), .ZN(n2450) );
  AOI22_X1 U32320 ( .A1(REG2_REG_15__SCAN_IN), .A2(n4684), .B1(n4622), .B2(
        n2450), .ZN(n4617) );
  NAND2_X1 U32330 ( .A1(n2452), .A2(IR_REG_31__SCAN_IN), .ZN(n2454) );
  INV_X1 U32340 ( .A(REG2_REG_16__SCAN_IN), .ZN(n4631) );
  NAND2_X1 U32350 ( .A1(n2455), .A2(n4682), .ZN(n2456) );
  NOR2_X1 U32360 ( .A1(n2729), .A2(REG2_REG_17__SCAN_IN), .ZN(n2457) );
  AOI21_X1 U32370 ( .B1(REG2_REG_17__SCAN_IN), .B2(n2729), .A(n2457), .ZN(
        n4643) );
  NAND2_X1 U32380 ( .A1(n2459), .A2(n2458), .ZN(n2464) );
  INV_X1 U32390 ( .A(REG2_REG_19__SCAN_IN), .ZN(n2462) );
  NAND2_X1 U32400 ( .A1(n2484), .A2(n2473), .ZN(n2811) );
  OR2_X1 U32410 ( .A1(n2484), .A2(n2473), .ZN(n2461) );
  MUX2_X1 U32420 ( .A(n2462), .B(REG2_REG_19__SCAN_IN), .S(n4094), .Z(n2463)
         );
  XNOR2_X1 U32430 ( .A(n2464), .B(n2463), .ZN(n2541) );
  NOR2_X1 U32440 ( .A1(IR_REG_19__SCAN_IN), .A2(IR_REG_18__SCAN_IN), .ZN(n2467) );
  NOR2_X1 U32450 ( .A1(IR_REG_5__SCAN_IN), .A2(IR_REG_22__SCAN_IN), .ZN(n2466)
         );
  NOR2_X1 U32460 ( .A1(IR_REG_23__SCAN_IN), .A2(IR_REG_24__SCAN_IN), .ZN(n2465) );
  NAND4_X1 U32470 ( .A1(n2474), .A2(n2467), .A3(n2466), .A4(n2465), .ZN(n2558)
         );
  INV_X1 U32480 ( .A(n2558), .ZN(n2468) );
  NAND2_X1 U32490 ( .A1(n2471), .A2(IR_REG_31__SCAN_IN), .ZN(n2472) );
  NAND2_X1 U32500 ( .A1(n2474), .A2(n2473), .ZN(n2475) );
  NAND2_X1 U32510 ( .A1(n2481), .A2(n4820), .ZN(n2480) );
  INV_X1 U32520 ( .A(n2480), .ZN(n2477) );
  NAND2_X1 U32530 ( .A1(IR_REG_24__SCAN_IN), .A2(IR_REG_23__SCAN_IN), .ZN(
        n4761) );
  NAND2_X1 U32540 ( .A1(n4761), .A2(IR_REG_31__SCAN_IN), .ZN(n2478) );
  OAI21_X1 U32550 ( .B1(IR_REG_31__SCAN_IN), .B2(n2859), .A(n2478), .ZN(n2479)
         );
  OR2_X1 U32560 ( .A1(n3136), .A2(U3149), .ZN(n4100) );
  NAND2_X1 U32570 ( .A1(n3146), .A2(n4100), .ZN(n2495) );
  XNOR2_X2 U32580 ( .A(n2482), .B(IR_REG_22__SCAN_IN), .ZN(n2895) );
  OAI21_X1 U32590 ( .B1(IR_REG_19__SCAN_IN), .B2(IR_REG_20__SCAN_IN), .A(
        IR_REG_31__SCAN_IN), .ZN(n2483) );
  AOI21_X1 U32600 ( .B1(n3136), .B2(n3125), .A(n2728), .ZN(n2493) );
  NAND2_X1 U32610 ( .A1(n2495), .A2(n2493), .ZN(n4614) );
  XNOR2_X1 U32620 ( .A(n2489), .B(n2486), .ZN(n3306) );
  NAND2_X1 U32630 ( .A1(n2556), .A2(n2486), .ZN(n2490) );
  OAI21_X1 U32640 ( .B1(n2491), .B2(n2490), .A(IR_REG_31__SCAN_IN), .ZN(n2492)
         );
  XNOR2_X1 U32650 ( .A(n2492), .B(n2555), .ZN(n4606) );
  OR2_X1 U32660 ( .A1(n3306), .A2(n4606), .ZN(n4096) );
  NAND2_X1 U32670 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n3815) );
  INV_X1 U32680 ( .A(n2493), .ZN(n2494) );
  NAND2_X1 U32690 ( .A1(n4657), .A2(ADDR_REG_19__SCAN_IN), .ZN(n2496) );
  OAI211_X1 U32700 ( .C1(n4668), .C2(n4094), .A(n3815), .B(n2496), .ZN(n2497)
         );
  NAND2_X1 U32710 ( .A1(n2498), .A2(n3357), .ZN(n2499) );
  OAI21_X1 U32720 ( .B1(n2498), .B2(n3357), .A(n2499), .ZN(n2505) );
  INV_X1 U32730 ( .A(REG1_REG_1__SCAN_IN), .ZN(n2500) );
  NAND2_X1 U32740 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(
        n2892) );
  INV_X1 U32750 ( .A(n2892), .ZN(n2502) );
  NAND2_X1 U32760 ( .A1(n2503), .A2(n2502), .ZN(n4118) );
  NAND2_X1 U32770 ( .A1(n2127), .A2(REG1_REG_1__SCAN_IN), .ZN(n3325) );
  NAND2_X1 U32780 ( .A1(n4118), .A2(n3325), .ZN(n2504) );
  NAND2_X1 U32790 ( .A1(n2505), .A2(n2504), .ZN(n3328) );
  NAND2_X1 U32800 ( .A1(n2498), .A2(REG1_REG_2__SCAN_IN), .ZN(n2506) );
  NAND2_X1 U32810 ( .A1(n2508), .A2(n4603), .ZN(n2509) );
  NAND2_X1 U32820 ( .A1(n2510), .A2(n4602), .ZN(n2511) );
  INV_X1 U32830 ( .A(REG1_REG_5__SCAN_IN), .ZN(n2512) );
  MUX2_X1 U32840 ( .A(n2512), .B(REG1_REG_5__SCAN_IN), .S(n4131), .Z(n4139) );
  OR2_X1 U32850 ( .A1(n4131), .A2(n2512), .ZN(n2513) );
  NAND2_X1 U32860 ( .A1(n4137), .A2(n2513), .ZN(n2514) );
  XNOR2_X1 U32870 ( .A(n2514), .B(n3268), .ZN(n3266) );
  NAND2_X1 U32880 ( .A1(n3266), .A2(REG1_REG_6__SCAN_IN), .ZN(n2516) );
  NAND2_X1 U32890 ( .A1(n2514), .A2(n4601), .ZN(n2515) );
  NAND2_X1 U32900 ( .A1(n2516), .A2(n2515), .ZN(n3276) );
  INV_X1 U32910 ( .A(REG1_REG_7__SCAN_IN), .ZN(n4723) );
  NOR2_X1 U32920 ( .A1(n4600), .A2(n4723), .ZN(n3275) );
  NAND2_X1 U32930 ( .A1(n4600), .A2(n4723), .ZN(n2517) );
  INV_X1 U32940 ( .A(REG1_REG_9__SCAN_IN), .ZN(n5004) );
  XNOR2_X1 U32950 ( .A(n4598), .B(n5004), .ZN(n4160) );
  NAND2_X1 U32960 ( .A1(n2519), .A2(n4597), .ZN(n2520) );
  XNOR2_X1 U32970 ( .A(n4185), .B(REG1_REG_11__SCAN_IN), .ZN(n4183) );
  INV_X1 U32980 ( .A(REG1_REG_11__SCAN_IN), .ZN(n2521) );
  OR2_X1 U32990 ( .A1(n4185), .A2(n2521), .ZN(n2522) );
  NAND2_X1 U33000 ( .A1(n2523), .A2(n4596), .ZN(n2524) );
  XNOR2_X1 U33010 ( .A(n4209), .B(REG1_REG_13__SCAN_IN), .ZN(n4207) );
  NAND2_X1 U33020 ( .A1(n4208), .A2(n4207), .ZN(n4206) );
  INV_X1 U33030 ( .A(REG1_REG_13__SCAN_IN), .ZN(n5005) );
  OR2_X1 U33040 ( .A1(n4209), .A2(n5005), .ZN(n2525) );
  INV_X1 U33050 ( .A(REG1_REG_14__SCAN_IN), .ZN(n4770) );
  INV_X1 U33060 ( .A(REG1_REG_15__SCAN_IN), .ZN(n2527) );
  AOI22_X1 U33070 ( .A1(REG1_REG_15__SCAN_IN), .A2(n4684), .B1(n4622), .B2(
        n2527), .ZN(n4619) );
  XNOR2_X1 U33080 ( .A(n2530), .B(n2529), .ZN(n4635) );
  INV_X1 U33090 ( .A(REG1_REG_16__SCAN_IN), .ZN(n4634) );
  NAND2_X1 U33100 ( .A1(n4635), .A2(n4634), .ZN(n4633) );
  NAND2_X1 U33110 ( .A1(n2530), .A2(n4682), .ZN(n2531) );
  INV_X1 U33120 ( .A(REG1_REG_17__SCAN_IN), .ZN(n4538) );
  AOI22_X1 U33130 ( .A1(n2729), .A2(REG1_REG_17__SCAN_IN), .B1(n4538), .B2(
        n2532), .ZN(n4646) );
  NAND2_X1 U33140 ( .A1(n2532), .A2(n4538), .ZN(n2533) );
  INV_X1 U33150 ( .A(REG1_REG_18__SCAN_IN), .ZN(n2743) );
  AOI22_X1 U33160 ( .A1(REG1_REG_18__SCAN_IN), .A2(n4679), .B1(n2535), .B2(
        n2743), .ZN(n4654) );
  XNOR2_X1 U33170 ( .A(n4094), .B(REG1_REG_19__SCAN_IN), .ZN(n2536) );
  XNOR2_X1 U33180 ( .A(n2537), .B(n2536), .ZN(n2538) );
  INV_X1 U33190 ( .A(n3306), .ZN(n4611) );
  NAND2_X1 U33200 ( .A1(n2538), .A2(n4648), .ZN(n2539) );
  OAI211_X1 U33210 ( .C1(n2541), .C2(n4615), .A(n2540), .B(n2539), .ZN(U3259)
         );
  INV_X1 U33220 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4795) );
  NAND2_X1 U33230 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .ZN(
        n2619) );
  INV_X1 U33240 ( .A(n2619), .ZN(n2542) );
  NAND2_X1 U33250 ( .A1(n2542), .A2(REG3_REG_5__SCAN_IN), .ZN(n2641) );
  NOR2_X1 U33260 ( .A1(n2641), .A2(n2640), .ZN(n2632) );
  NAND2_X1 U33270 ( .A1(n2632), .A2(REG3_REG_7__SCAN_IN), .ZN(n2655) );
  INV_X1 U33280 ( .A(n2664), .ZN(n2543) );
  NAND2_X1 U33290 ( .A1(n2543), .A2(REG3_REG_9__SCAN_IN), .ZN(n2673) );
  OR2_X2 U33300 ( .A1(n2700), .A2(n4999), .ZN(n2716) );
  INV_X1 U33310 ( .A(n2716), .ZN(n2546) );
  NAND2_X1 U33320 ( .A1(REG3_REG_17__SCAN_IN), .A2(REG3_REG_18__SCAN_IN), .ZN(
        n2548) );
  OR2_X2 U33330 ( .A1(n2739), .A2(n2548), .ZN(n2750) );
  NAND2_X1 U33340 ( .A1(REG3_REG_21__SCAN_IN), .A2(REG3_REG_20__SCAN_IN), .ZN(
        n2550) );
  OR2_X2 U33350 ( .A1(n2781), .A2(n4792), .ZN(n2790) );
  INV_X1 U33360 ( .A(n2790), .ZN(n2552) );
  OR2_X2 U33370 ( .A1(n2800), .A2(n4988), .ZN(n2802) );
  INV_X1 U33380 ( .A(n2802), .ZN(n2553) );
  INV_X1 U33390 ( .A(REG3_REG_26__SCAN_IN), .ZN(n3919) );
  NAND2_X1 U33400 ( .A1(n2802), .A2(n3919), .ZN(n2554) );
  NAND2_X1 U33410 ( .A1(n2845), .A2(n2554), .ZN(n4253) );
  NAND4_X1 U33420 ( .A1(n2556), .A2(n2469), .A3(n2555), .A4(n2486), .ZN(n2557)
         );
  NOR2_X1 U33430 ( .A1(n2558), .A2(n2557), .ZN(n2561) );
  NAND3_X1 U33440 ( .A1(n2561), .A2(n2560), .A3(n2559), .ZN(n2562) );
  NOR2_X2 U33450 ( .A1(n2562), .A2(IR_REG_29__SCAN_IN), .ZN(n3772) );
  NAND2_X1 U33460 ( .A1(n2562), .A2(IR_REG_31__SCAN_IN), .ZN(n2563) );
  OR2_X2 U33470 ( .A1(n2565), .A2(n4590), .ZN(n2590) );
  INV_X1 U33480 ( .A(n2591), .ZN(n2805) );
  INV_X1 U33490 ( .A(n4590), .ZN(n2564) );
  NAND2_X1 U33500 ( .A1(n3964), .A2(REG2_REG_26__SCAN_IN), .ZN(n2568) );
  NAND2_X1 U33510 ( .A1(n2606), .A2(REG1_REG_26__SCAN_IN), .ZN(n2567) );
  OAI211_X1 U33520 ( .C1(n2805), .C2(n4795), .A(n2568), .B(n2567), .ZN(n2569)
         );
  INV_X1 U3353 ( .A(n2569), .ZN(n2570) );
  AND2_X2 U33540 ( .A1(n2571), .A2(n2570), .ZN(n4234) );
  AND2_X1 U3355 ( .A1(n4267), .A2(n3174), .ZN(n3974) );
  INV_X1 U3356 ( .A(n3974), .ZN(n2572) );
  NAND2_X1 U3357 ( .A1(n4234), .A2(n3928), .ZN(n3187) );
  NAND2_X1 U3358 ( .A1(n2572), .A2(n3187), .ZN(n4020) );
  NAND2_X1 U3359 ( .A1(n2621), .A2(REG2_REG_1__SCAN_IN), .ZN(n2577) );
  NAND2_X1 U3360 ( .A1(n2639), .A2(REG3_REG_1__SCAN_IN), .ZN(n2576) );
  INV_X1 U3361 ( .A(REG0_REG_1__SCAN_IN), .ZN(n2573) );
  NAND2_X1 U3362 ( .A1(n2606), .A2(REG1_REG_1__SCAN_IN), .ZN(n2574) );
  AND4_X2 U3363 ( .A1(n2577), .A2(n2576), .A3(n2575), .A4(n2574), .ZN(n2897)
         );
  INV_X1 U3364 ( .A(n2897), .ZN(n2601) );
  INV_X1 U3365 ( .A(n2612), .ZN(n2578) );
  NAND2_X1 U3366 ( .A1(n2601), .A2(n3798), .ZN(n4025) );
  NAND2_X1 U3367 ( .A1(n3455), .A2(n2897), .ZN(n4029) );
  NAND2_X1 U3368 ( .A1(n4025), .A2(n4029), .ZN(n2817) );
  OAI21_X2 U3369 ( .B1(n4685), .B2(n2612), .A(n2581), .ZN(n3296) );
  NAND2_X1 U3370 ( .A1(n2621), .A2(REG2_REG_0__SCAN_IN), .ZN(n2586) );
  NAND2_X1 U3371 ( .A1(n2591), .A2(REG0_REG_0__SCAN_IN), .ZN(n2585) );
  INV_X1 U3372 ( .A(REG3_REG_0__SCAN_IN), .ZN(n2582) );
  NAND4_X2 U3373 ( .A1(n2586), .A2(n2585), .A3(n2584), .A4(n2583), .ZN(n4111)
         );
  AND2_X1 U3374 ( .A1(n3296), .A2(n4111), .ZN(n3452) );
  NAND2_X1 U3375 ( .A1(n2817), .A2(n3452), .ZN(n3343) );
  NAND2_X1 U3376 ( .A1(n2621), .A2(REG2_REG_2__SCAN_IN), .ZN(n2595) );
  NAND2_X1 U3377 ( .A1(n2639), .A2(REG3_REG_2__SCAN_IN), .ZN(n2594) );
  NAND2_X1 U3378 ( .A1(n2591), .A2(REG0_REG_2__SCAN_IN), .ZN(n2593) );
  NAND2_X1 U3379 ( .A1(n2606), .A2(REG1_REG_2__SCAN_IN), .ZN(n2592) );
  NAND2_X1 U3380 ( .A1(n3355), .A2(n3789), .ZN(n4028) );
  NAND2_X1 U3381 ( .A1(n3350), .A2(n2909), .ZN(n4031) );
  NAND2_X1 U3382 ( .A1(n4028), .A2(n4031), .ZN(n3995) );
  INV_X1 U3383 ( .A(REG3_REG_3__SCAN_IN), .ZN(n2596) );
  NAND2_X1 U3384 ( .A1(n2639), .A2(n2596), .ZN(n2600) );
  NAND2_X1 U3385 ( .A1(n2606), .A2(REG1_REG_3__SCAN_IN), .ZN(n2599) );
  NAND2_X1 U3386 ( .A1(n2621), .A2(REG2_REG_3__SCAN_IN), .ZN(n2598) );
  NAND2_X1 U3387 ( .A1(n2591), .A2(REG0_REG_3__SCAN_IN), .ZN(n2597) );
  NAND4_X1 U3388 ( .A1(n2600), .A2(n2599), .A3(n2598), .A4(n2597), .ZN(n4110)
         );
  NAND2_X1 U3389 ( .A1(n3507), .A2(n4110), .ZN(n2602) );
  NAND2_X1 U3390 ( .A1(n3455), .A2(n2601), .ZN(n3344) );
  NAND4_X1 U3391 ( .A1(n3343), .A2(n3995), .A3(n2602), .A4(n3344), .ZN(n2604)
         );
  AND2_X1 U3392 ( .A1(n3350), .A2(n3789), .ZN(n3496) );
  INV_X1 U3393 ( .A(n3507), .ZN(n3501) );
  AOI22_X1 U3394 ( .A1(n3496), .A2(n2602), .B1(n3392), .B2(n3501), .ZN(n2603)
         );
  OAI21_X1 U3395 ( .B1(REG3_REG_3__SCAN_IN), .B2(REG3_REG_4__SCAN_IN), .A(
        n2619), .ZN(n3401) );
  OR2_X1 U3396 ( .A1(n2605), .A2(n3401), .ZN(n2610) );
  NAND2_X1 U3397 ( .A1(n2591), .A2(REG0_REG_4__SCAN_IN), .ZN(n2609) );
  NAND2_X1 U3398 ( .A1(n2606), .A2(REG1_REG_4__SCAN_IN), .ZN(n2608) );
  NAND2_X1 U3399 ( .A1(n2621), .A2(REG2_REG_4__SCAN_IN), .ZN(n2607) );
  INV_X1 U3400 ( .A(DATAI_4_), .ZN(n2611) );
  NAND2_X1 U3401 ( .A1(n4035), .A2(n4037), .ZN(n3390) );
  INV_X1 U3402 ( .A(n4131), .ZN(n2614) );
  INV_X1 U3403 ( .A(DATAI_5_), .ZN(n2615) );
  NAND2_X1 U3404 ( .A1(n2591), .A2(REG0_REG_5__SCAN_IN), .ZN(n2625) );
  NAND2_X1 U3405 ( .A1(n2606), .A2(REG1_REG_5__SCAN_IN), .ZN(n2624) );
  INV_X1 U3406 ( .A(REG3_REG_5__SCAN_IN), .ZN(n2618) );
  NAND2_X1 U3407 ( .A1(n2619), .A2(n2618), .ZN(n2620) );
  AND2_X1 U3408 ( .A1(n2641), .A2(n2620), .ZN(n3544) );
  NAND2_X1 U3409 ( .A1(n2639), .A2(n3544), .ZN(n2623) );
  NAND2_X1 U3410 ( .A1(n2621), .A2(REG2_REG_5__SCAN_IN), .ZN(n2622) );
  NAND2_X1 U3411 ( .A1(n3538), .A2(n2626), .ZN(n2628) );
  NAND2_X1 U3412 ( .A1(n3542), .A2(n4108), .ZN(n2627) );
  NAND2_X1 U3413 ( .A1(n3396), .A2(n3535), .ZN(n3539) );
  NAND2_X1 U3414 ( .A1(n2375), .A2(n2628), .ZN(n2629) );
  INV_X1 U3415 ( .A(DATAI_7_), .ZN(n4733) );
  NAND2_X1 U3416 ( .A1(n2591), .A2(REG0_REG_7__SCAN_IN), .ZN(n2638) );
  NAND2_X1 U3417 ( .A1(n2606), .A2(REG1_REG_7__SCAN_IN), .ZN(n2637) );
  INV_X1 U3418 ( .A(n2632), .ZN(n2643) );
  INV_X1 U3419 ( .A(REG3_REG_7__SCAN_IN), .ZN(n2633) );
  NAND2_X1 U3420 ( .A1(n2643), .A2(n2633), .ZN(n2634) );
  AND2_X1 U3421 ( .A1(n2655), .A2(n2634), .ZN(n3585) );
  NAND2_X1 U3422 ( .A1(n2639), .A2(n3585), .ZN(n2636) );
  NAND2_X1 U3423 ( .A1(n2621), .A2(REG2_REG_7__SCAN_IN), .ZN(n2635) );
  NAND2_X1 U3424 ( .A1(n3580), .A2(n4107), .ZN(n4046) );
  MUX2_X1 U3425 ( .A(n4601), .B(DATAI_6_), .S(n2612), .Z(n3588) );
  NAND2_X1 U3426 ( .A1(n2591), .A2(REG0_REG_6__SCAN_IN), .ZN(n2647) );
  NAND2_X1 U3427 ( .A1(n2606), .A2(REG1_REG_6__SCAN_IN), .ZN(n2646) );
  NAND2_X1 U3428 ( .A1(n2641), .A2(n2640), .ZN(n2642) );
  AND2_X1 U3429 ( .A1(n2643), .A2(n2642), .ZN(n3514) );
  NAND2_X1 U3430 ( .A1(n3155), .A2(n3514), .ZN(n2645) );
  NAND2_X1 U3431 ( .A1(n2621), .A2(REG2_REG_6__SCAN_IN), .ZN(n2644) );
  NAND4_X1 U3432 ( .A1(n2647), .A2(n2646), .A3(n2645), .A4(n2644), .ZN(n3589)
         );
  INV_X1 U3433 ( .A(n3589), .ZN(n2648) );
  NAND2_X1 U3434 ( .A1(n2880), .A2(n2648), .ZN(n2649) );
  AND2_X1 U3435 ( .A1(n3588), .A2(n3589), .ZN(n2651) );
  AOI22_X1 U3436 ( .A1(n3592), .A2(n2651), .B1(n3581), .B2(n4107), .ZN(n2652)
         );
  NAND2_X1 U3437 ( .A1(n2653), .A2(n2652), .ZN(n3425) );
  INV_X1 U3438 ( .A(DATAI_8_), .ZN(n2654) );
  MUX2_X1 U3439 ( .A(n4146), .B(n2654), .S(n3968), .Z(n3557) );
  NAND2_X1 U3440 ( .A1(n2591), .A2(REG0_REG_8__SCAN_IN), .ZN(n2660) );
  NAND2_X1 U3441 ( .A1(n2606), .A2(REG1_REG_8__SCAN_IN), .ZN(n2659) );
  NAND2_X1 U3442 ( .A1(n2655), .A2(n4730), .ZN(n2656) );
  AND2_X1 U3443 ( .A1(n2664), .A2(n2656), .ZN(n3569) );
  NAND2_X1 U3444 ( .A1(n3155), .A2(n3569), .ZN(n2658) );
  NAND2_X1 U3445 ( .A1(n2621), .A2(REG2_REG_8__SCAN_IN), .ZN(n2657) );
  NAND2_X1 U3446 ( .A1(n3557), .A2(n3467), .ZN(n2661) );
  NAND2_X1 U3447 ( .A1(n3425), .A2(n2661), .ZN(n2663) );
  INV_X1 U3448 ( .A(n3557), .ZN(n3434) );
  NAND2_X1 U3449 ( .A1(n3434), .A2(n3703), .ZN(n2662) );
  NAND2_X1 U3450 ( .A1(n2663), .A2(n2662), .ZN(n3465) );
  MUX2_X1 U3451 ( .A(n4598), .B(DATAI_9_), .S(n3968), .Z(n3473) );
  NAND2_X1 U3452 ( .A1(n2591), .A2(REG0_REG_9__SCAN_IN), .ZN(n2669) );
  NAND2_X1 U3453 ( .A1(n2606), .A2(REG1_REG_9__SCAN_IN), .ZN(n2668) );
  INV_X1 U3454 ( .A(REG3_REG_9__SCAN_IN), .ZN(n4913) );
  NAND2_X1 U3455 ( .A1(n2664), .A2(n4913), .ZN(n2665) );
  AND2_X1 U3456 ( .A1(n2673), .A2(n2665), .ZN(n3707) );
  NAND2_X1 U3457 ( .A1(n3155), .A2(n3707), .ZN(n2667) );
  NAND2_X1 U34580 ( .A1(n2621), .A2(REG2_REG_9__SCAN_IN), .ZN(n2666) );
  NAND4_X1 U34590 ( .A1(n2669), .A2(n2668), .A3(n2667), .A4(n2666), .ZN(n4106)
         );
  AND2_X1 U3460 ( .A1(n3473), .A2(n4106), .ZN(n2671) );
  INV_X1 U3461 ( .A(n3473), .ZN(n3705) );
  INV_X1 U3462 ( .A(n4106), .ZN(n2952) );
  NAND2_X1 U3463 ( .A1(n3705), .A2(n2952), .ZN(n2670) );
  MUX2_X1 U3464 ( .A(n4597), .B(DATAI_10_), .S(n2612), .Z(n3735) );
  NAND2_X1 U3465 ( .A1(n2591), .A2(REG0_REG_10__SCAN_IN), .ZN(n2678) );
  NAND2_X1 U3466 ( .A1(n2606), .A2(REG1_REG_10__SCAN_IN), .ZN(n2677) );
  NAND2_X1 U34670 ( .A1(n2673), .A2(n2672), .ZN(n2674) );
  AND2_X1 U3468 ( .A1(n2681), .A2(n2674), .ZN(n3525) );
  NAND2_X1 U34690 ( .A1(n3155), .A2(n3525), .ZN(n2676) );
  NAND2_X1 U3470 ( .A1(n2621), .A2(REG2_REG_10__SCAN_IN), .ZN(n2675) );
  NAND4_X1 U34710 ( .A1(n2678), .A2(n2677), .A3(n2676), .A4(n2675), .ZN(n3490)
         );
  NOR2_X1 U3472 ( .A1(n3735), .A2(n3490), .ZN(n2679) );
  INV_X1 U34730 ( .A(DATAI_11_), .ZN(n3247) );
  MUX2_X1 U3474 ( .A(n4185), .B(n3247), .S(n3968), .Z(n2977) );
  INV_X1 U34750 ( .A(REG3_REG_11__SCAN_IN), .ZN(n2680) );
  NAND2_X1 U3476 ( .A1(n2681), .A2(n2680), .ZN(n2682) );
  NAND2_X1 U34770 ( .A1(n2693), .A2(n2682), .ZN(n3617) );
  OR2_X1 U3478 ( .A1(n3617), .A2(n2605), .ZN(n2686) );
  NAND2_X1 U34790 ( .A1(n2591), .A2(REG0_REG_11__SCAN_IN), .ZN(n2685) );
  NAND2_X1 U3480 ( .A1(n2606), .A2(REG1_REG_11__SCAN_IN), .ZN(n2684) );
  NAND2_X1 U34810 ( .A1(n3964), .A2(REG2_REG_11__SCAN_IN), .ZN(n2683) );
  NAND4_X1 U3482 ( .A1(n2686), .A2(n2685), .A3(n2684), .A4(n2683), .ZN(n4105)
         );
  NAND2_X1 U34830 ( .A1(n2977), .A2(n4105), .ZN(n3649) );
  INV_X1 U3484 ( .A(n2977), .ZN(n3616) );
  INV_X1 U34850 ( .A(n4105), .ZN(n3733) );
  NAND2_X1 U3486 ( .A1(n3616), .A2(n3733), .ZN(n3647) );
  INV_X1 U34870 ( .A(n3643), .ZN(n3784) );
  XNOR2_X1 U3488 ( .A(n2716), .B(REG3_REG_14__SCAN_IN), .ZN(n3786) );
  NAND2_X1 U34890 ( .A1(n3786), .A2(n3155), .ZN(n2691) );
  NAND2_X1 U3490 ( .A1(n2591), .A2(REG0_REG_14__SCAN_IN), .ZN(n2688) );
  NAND2_X1 U34910 ( .A1(n3964), .A2(REG2_REG_14__SCAN_IN), .ZN(n2687) );
  OAI211_X1 U3492 ( .C1(n3153), .C2(n4770), .A(n2688), .B(n2687), .ZN(n2689)
         );
  INV_X1 U34930 ( .A(n2689), .ZN(n2690) );
  NAND2_X1 U3494 ( .A1(n3784), .A2(n4103), .ZN(n3951) );
  NAND2_X1 U34950 ( .A1(n4463), .A2(n3643), .ZN(n3947) );
  INV_X1 U3496 ( .A(n2621), .ZN(n2794) );
  INV_X1 U34970 ( .A(REG2_REG_12__SCAN_IN), .ZN(n3658) );
  NAND2_X1 U3498 ( .A1(n2693), .A2(n2692), .ZN(n2694) );
  NAND2_X1 U34990 ( .A1(n2700), .A2(n2694), .ZN(n3657) );
  OR2_X1 U3500 ( .A1(n3657), .A2(n2605), .ZN(n2698) );
  NAND2_X1 U35010 ( .A1(n2591), .A2(REG0_REG_12__SCAN_IN), .ZN(n2696) );
  NAND2_X1 U3502 ( .A1(n2606), .A2(REG1_REG_12__SCAN_IN), .ZN(n2695) );
  AND2_X1 U35030 ( .A1(n2696), .A2(n2695), .ZN(n2697) );
  OAI211_X1 U3504 ( .C1(n2794), .C2(n3658), .A(n2698), .B(n2697), .ZN(n3256)
         );
  INV_X1 U35050 ( .A(n3256), .ZN(n3714) );
  NAND2_X1 U35060 ( .A1(n3660), .A2(n3714), .ZN(n3681) );
  INV_X1 U35070 ( .A(DATAI_13_), .ZN(n2699) );
  NAND2_X1 U35080 ( .A1(n2700), .A2(n4999), .ZN(n2701) );
  AND2_X1 U35090 ( .A1(n2716), .A2(n2701), .ZN(n3719) );
  NAND2_X1 U35100 ( .A1(n3719), .A2(n3155), .ZN(n2704) );
  AOI22_X1 U35110 ( .A1(n2606), .A2(REG1_REG_13__SCAN_IN), .B1(n2591), .B2(
        REG0_REG_13__SCAN_IN), .ZN(n2703) );
  NAND2_X1 U35120 ( .A1(n2621), .A2(REG2_REG_13__SCAN_IN), .ZN(n2702) );
  NAND2_X1 U35130 ( .A1(n3717), .A2(n3780), .ZN(n2705) );
  AND2_X1 U35140 ( .A1(n3681), .A2(n2705), .ZN(n2709) );
  NAND2_X1 U35150 ( .A1(n3652), .A2(n3256), .ZN(n3679) );
  INV_X1 U35160 ( .A(n3679), .ZN(n2706) );
  NAND2_X1 U35170 ( .A1(n2709), .A2(n2706), .ZN(n2708) );
  NAND2_X1 U35180 ( .A1(n3686), .A2(n4104), .ZN(n2707) );
  NAND2_X1 U35190 ( .A1(n2829), .A2(n3638), .ZN(n2710) );
  NAND2_X1 U35200 ( .A1(n2977), .A2(n3733), .ZN(n3655) );
  AND2_X1 U35210 ( .A1(n3655), .A2(n2709), .ZN(n3637) );
  OR2_X1 U35220 ( .A1(n2710), .A2(n3637), .ZN(n2711) );
  OAI21_X2 U35230 ( .B1(n3608), .B2(n2712), .A(n2711), .ZN(n3641) );
  INV_X1 U35240 ( .A(n3641), .ZN(n2714) );
  NAND2_X1 U35250 ( .A1(n3784), .A2(n4463), .ZN(n2713) );
  INV_X1 U35260 ( .A(REG3_REG_14__SCAN_IN), .ZN(n2715) );
  INV_X1 U35270 ( .A(REG3_REG_15__SCAN_IN), .ZN(n5008) );
  OAI21_X1 U35280 ( .B1(n2716), .B2(n2715), .A(n5008), .ZN(n2717) );
  NAND2_X1 U35290 ( .A1(n2720), .A2(n2717), .ZN(n3936) );
  OR2_X1 U35300 ( .A1(n3936), .A2(n2605), .ZN(n2719) );
  AOI22_X1 U35310 ( .A1(n2606), .A2(REG1_REG_15__SCAN_IN), .B1(n2591), .B2(
        REG0_REG_15__SCAN_IN), .ZN(n2718) );
  OAI211_X1 U35320 ( .C1(n2794), .C2(n2450), .A(n2719), .B(n2718), .ZN(n3782)
         );
  MUX2_X1 U35330 ( .A(n4622), .B(DATAI_15_), .S(n3968), .Z(n4474) );
  INV_X1 U35340 ( .A(n3782), .ZN(n4436) );
  INV_X1 U35350 ( .A(DATAI_16_), .ZN(n4681) );
  MUX2_X1 U35360 ( .A(n4681), .B(n4682), .S(n2728), .Z(n4435) );
  INV_X1 U35370 ( .A(REG3_REG_16__SCAN_IN), .ZN(n4867) );
  NAND2_X1 U35380 ( .A1(n2720), .A2(n4867), .ZN(n2721) );
  NAND2_X1 U35390 ( .A1(n2739), .A2(n2721), .ZN(n4448) );
  OR2_X1 U35400 ( .A1(n4448), .A2(n2605), .ZN(n2726) );
  NAND2_X1 U35410 ( .A1(n2591), .A2(REG0_REG_16__SCAN_IN), .ZN(n2723) );
  NAND2_X1 U35420 ( .A1(n3964), .A2(REG2_REG_16__SCAN_IN), .ZN(n2722) );
  OAI211_X1 U35430 ( .C1(n3153), .C2(n4634), .A(n2723), .B(n2722), .ZN(n2724)
         );
  INV_X1 U35440 ( .A(n2724), .ZN(n2725) );
  NAND2_X1 U35450 ( .A1(n2726), .A2(n2725), .ZN(n4416) );
  OR2_X1 U35460 ( .A1(n4435), .A2(n4416), .ZN(n4065) );
  NAND2_X1 U35470 ( .A1(n4435), .A2(n4416), .ZN(n4412) );
  NAND2_X1 U35480 ( .A1(n4065), .A2(n4412), .ZN(n4450) );
  INV_X1 U35490 ( .A(n4416), .ZN(n4465) );
  MUX2_X1 U35500 ( .A(DATAI_17_), .B(n2729), .S(n2728), .Z(n4427) );
  INV_X1 U35510 ( .A(n4427), .ZN(n4423) );
  XNOR2_X1 U35520 ( .A(n2739), .B(REG3_REG_17__SCAN_IN), .ZN(n4430) );
  NAND2_X1 U35530 ( .A1(n4430), .A2(n3155), .ZN(n2734) );
  INV_X1 U35540 ( .A(REG2_REG_17__SCAN_IN), .ZN(n4989) );
  NAND2_X1 U35550 ( .A1(n2591), .A2(REG0_REG_17__SCAN_IN), .ZN(n2731) );
  NAND2_X1 U35560 ( .A1(n2606), .A2(REG1_REG_17__SCAN_IN), .ZN(n2730) );
  OAI211_X1 U35570 ( .C1(n4989), .C2(n2794), .A(n2731), .B(n2730), .ZN(n2732)
         );
  INV_X1 U35580 ( .A(n2732), .ZN(n2733) );
  NAND2_X1 U35590 ( .A1(n4423), .A2(n4437), .ZN(n2736) );
  INV_X1 U35600 ( .A(REG3_REG_17__SCAN_IN), .ZN(n2738) );
  INV_X1 U35610 ( .A(REG3_REG_18__SCAN_IN), .ZN(n2737) );
  OAI21_X1 U35620 ( .B1(n2739), .B2(n2738), .A(n2737), .ZN(n2740) );
  AND2_X1 U35630 ( .A1(n2740), .A2(n2750), .ZN(n4407) );
  NAND2_X1 U35640 ( .A1(n4407), .A2(n3155), .ZN(n2746) );
  NAND2_X1 U35650 ( .A1(n2591), .A2(REG0_REG_18__SCAN_IN), .ZN(n2742) );
  NAND2_X1 U35660 ( .A1(n3964), .A2(REG2_REG_18__SCAN_IN), .ZN(n2741) );
  OAI211_X1 U35670 ( .C1(n3153), .C2(n2743), .A(n2742), .B(n2741), .ZN(n2744)
         );
  INV_X1 U35680 ( .A(n2744), .ZN(n2745) );
  INV_X1 U35690 ( .A(DATAI_18_), .ZN(n2747) );
  MUX2_X1 U35700 ( .A(n4679), .B(n2747), .S(n3968), .Z(n4405) );
  OR2_X1 U35710 ( .A1(n4419), .A2(n4405), .ZN(n4377) );
  NAND2_X1 U35720 ( .A1(n4419), .A2(n4405), .ZN(n4378) );
  NAND2_X1 U35730 ( .A1(n4377), .A2(n4378), .ZN(n4403) );
  NAND2_X1 U35740 ( .A1(n4404), .A2(n4403), .ZN(n4402) );
  INV_X1 U35750 ( .A(n4419), .ZN(n2748) );
  NAND2_X1 U35760 ( .A1(n2748), .A2(n4405), .ZN(n2749) );
  NAND2_X1 U35770 ( .A1(n4402), .A2(n2749), .ZN(n4386) );
  INV_X1 U35780 ( .A(REG3_REG_19__SCAN_IN), .ZN(n4734) );
  NAND2_X1 U35790 ( .A1(n2750), .A2(n4734), .ZN(n2751) );
  NAND2_X1 U35800 ( .A1(n2765), .A2(n2751), .ZN(n4391) );
  OR2_X1 U35810 ( .A1(n4391), .A2(n2605), .ZN(n2756) );
  INV_X1 U3582 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4947) );
  NAND2_X1 U3583 ( .A1(n3964), .A2(REG2_REG_19__SCAN_IN), .ZN(n2753) );
  NAND2_X1 U3584 ( .A1(n2606), .A2(REG1_REG_19__SCAN_IN), .ZN(n2752) );
  OAI211_X1 U3585 ( .C1(n2805), .C2(n4947), .A(n2753), .B(n2752), .ZN(n2754)
         );
  INV_X1 U3586 ( .A(n2754), .ZN(n2755) );
  MUX2_X1 U3587 ( .A(n4593), .B(DATAI_19_), .S(n3968), .Z(n4382) );
  NAND2_X1 U3588 ( .A1(n4398), .A2(n4382), .ZN(n2757) );
  INV_X1 U3589 ( .A(n4398), .ZN(n2833) );
  XNOR2_X1 U3590 ( .A(n2765), .B(REG3_REG_20__SCAN_IN), .ZN(n4371) );
  NAND2_X1 U3591 ( .A1(n4371), .A2(n3155), .ZN(n2762) );
  INV_X1 U3592 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4946) );
  NAND2_X1 U3593 ( .A1(n2591), .A2(REG0_REG_20__SCAN_IN), .ZN(n2759) );
  NAND2_X1 U3594 ( .A1(n3964), .A2(REG2_REG_20__SCAN_IN), .ZN(n2758) );
  OAI211_X1 U3595 ( .C1(n3153), .C2(n4946), .A(n2759), .B(n2758), .ZN(n2760)
         );
  INV_X1 U3596 ( .A(n2760), .ZN(n2761) );
  INV_X1 U3597 ( .A(REG3_REG_20__SCAN_IN), .ZN(n2764) );
  INV_X1 U3598 ( .A(REG3_REG_21__SCAN_IN), .ZN(n2763) );
  OAI21_X1 U3599 ( .B1(n2765), .B2(n2764), .A(n2763), .ZN(n2766) );
  AND2_X1 U3600 ( .A1(n2766), .A2(n2772), .ZN(n4348) );
  NAND2_X1 U3601 ( .A1(n4348), .A2(n3155), .ZN(n2771) );
  INV_X1 U3602 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4790) );
  NAND2_X1 U3603 ( .A1(n2591), .A2(REG0_REG_21__SCAN_IN), .ZN(n2768) );
  NAND2_X1 U3604 ( .A1(n3964), .A2(REG2_REG_21__SCAN_IN), .ZN(n2767) );
  OAI211_X1 U3605 ( .C1(n3153), .C2(n4790), .A(n2768), .B(n2767), .ZN(n2769)
         );
  INV_X1 U3606 ( .A(n2769), .ZN(n2770) );
  INV_X1 U3607 ( .A(REG3_REG_22__SCAN_IN), .ZN(n4977) );
  NAND2_X1 U3608 ( .A1(n2772), .A2(n4977), .ZN(n2773) );
  NAND2_X1 U3609 ( .A1(n2781), .A2(n2773), .ZN(n3899) );
  OR2_X1 U3610 ( .A1(n3899), .A2(n2605), .ZN(n2779) );
  INV_X1 U3611 ( .A(REG2_REG_22__SCAN_IN), .ZN(n2776) );
  NAND2_X1 U3612 ( .A1(n2591), .A2(REG0_REG_22__SCAN_IN), .ZN(n2775) );
  NAND2_X1 U3613 ( .A1(n2606), .A2(REG1_REG_22__SCAN_IN), .ZN(n2774) );
  OAI211_X1 U3614 ( .C1(n2776), .C2(n2794), .A(n2775), .B(n2774), .ZN(n2777)
         );
  INV_X1 U3615 ( .A(n2777), .ZN(n2778) );
  NAND2_X1 U3616 ( .A1(n4341), .A2(n4332), .ZN(n4302) );
  INV_X1 U3617 ( .A(n4332), .ZN(n3069) );
  NAND2_X1 U3618 ( .A1(n3805), .A2(n3069), .ZN(n2839) );
  NAND2_X1 U3619 ( .A1(n4302), .A2(n2839), .ZN(n4320) );
  NAND2_X1 U3620 ( .A1(n3805), .A2(n4332), .ZN(n2780) );
  NAND2_X1 U3621 ( .A1(n4319), .A2(n2780), .ZN(n4297) );
  NAND2_X1 U3622 ( .A1(n2781), .A2(n4792), .ZN(n2782) );
  NAND2_X1 U3623 ( .A1(n2790), .A2(n2782), .ZN(n4309) );
  INV_X1 U3624 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4793) );
  NAND2_X1 U3625 ( .A1(n3964), .A2(REG2_REG_23__SCAN_IN), .ZN(n2784) );
  NAND2_X1 U3626 ( .A1(n2591), .A2(REG0_REG_23__SCAN_IN), .ZN(n2783) );
  OAI211_X1 U3627 ( .C1(n3153), .C2(n4793), .A(n2784), .B(n2783), .ZN(n2785)
         );
  INV_X1 U3628 ( .A(n2785), .ZN(n2786) );
  NAND2_X1 U3629 ( .A1(n4297), .A2(n2376), .ZN(n2789) );
  NAND2_X1 U3630 ( .A1(n4326), .A2(n3070), .ZN(n2788) );
  INV_X1 U3631 ( .A(REG3_REG_24__SCAN_IN), .ZN(n4991) );
  NAND2_X1 U3632 ( .A1(n2790), .A2(n4991), .ZN(n2791) );
  NAND2_X1 U3633 ( .A1(n2800), .A2(n2791), .ZN(n3877) );
  INV_X1 U3634 ( .A(REG2_REG_24__SCAN_IN), .ZN(n2795) );
  NAND2_X1 U3635 ( .A1(n2591), .A2(REG0_REG_24__SCAN_IN), .ZN(n2793) );
  NAND2_X1 U3636 ( .A1(n2606), .A2(REG1_REG_24__SCAN_IN), .ZN(n2792) );
  OAI211_X1 U3637 ( .C1(n2795), .C2(n2794), .A(n2793), .B(n2792), .ZN(n2796)
         );
  INV_X1 U3638 ( .A(n2796), .ZN(n2797) );
  NAND2_X1 U3639 ( .A1(n4265), .A2(n4290), .ZN(n2799) );
  INV_X1 U3640 ( .A(n4259), .ZN(n2809) );
  NAND2_X1 U3641 ( .A1(n2800), .A2(n4988), .ZN(n2801) );
  NAND2_X1 U3642 ( .A1(n4274), .A2(n3155), .ZN(n2808) );
  INV_X1 U3643 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4796) );
  NAND2_X1 U3644 ( .A1(n2606), .A2(REG1_REG_25__SCAN_IN), .ZN(n2804) );
  NAND2_X1 U3645 ( .A1(n3964), .A2(REG2_REG_25__SCAN_IN), .ZN(n2803) );
  OAI211_X1 U3646 ( .C1(n4796), .C2(n2805), .A(n2804), .B(n2803), .ZN(n2806)
         );
  INV_X1 U3647 ( .A(n2806), .ZN(n2807) );
  NAND2_X1 U3648 ( .A1(n4286), .A2(n3843), .ZN(n2810) );
  XNOR2_X1 U3649 ( .A(n3185), .B(n2895), .ZN(n2815) );
  NAND2_X1 U3650 ( .A1(n2884), .A2(n4593), .ZN(n3442) );
  NAND2_X1 U3651 ( .A1(n2818), .A2(n4027), .ZN(n2819) );
  INV_X1 U3652 ( .A(n3995), .ZN(n3348) );
  NAND2_X1 U3653 ( .A1(n3346), .A2(n3348), .ZN(n3347) );
  NAND2_X1 U3654 ( .A1(n3347), .A2(n4028), .ZN(n3499) );
  NAND2_X1 U3655 ( .A1(n3507), .A2(n3392), .ZN(n4034) );
  NAND2_X1 U3656 ( .A1(n3501), .A2(n4110), .ZN(n4032) );
  NAND2_X1 U3657 ( .A1(n3499), .A2(n4004), .ZN(n2820) );
  INV_X1 U3658 ( .A(n4035), .ZN(n2821) );
  NAND2_X1 U3659 ( .A1(n3542), .A2(n2626), .ZN(n4041) );
  AND2_X1 U3660 ( .A1(n3538), .A2(n4108), .ZN(n3532) );
  NAND2_X1 U3661 ( .A1(n2880), .A2(n3589), .ZN(n4039) );
  NAND2_X1 U3662 ( .A1(n3588), .A2(n2648), .ZN(n4043) );
  NAND2_X1 U3663 ( .A1(n2822), .A2(n4043), .ZN(n3576) );
  NAND2_X1 U3664 ( .A1(n3434), .A2(n3467), .ZN(n4049) );
  NAND2_X1 U3665 ( .A1(n3557), .A2(n3703), .ZN(n4045) );
  AND2_X1 U3666 ( .A1(n3705), .A2(n4106), .ZN(n4053) );
  NAND2_X1 U3667 ( .A1(n3473), .A2(n2952), .ZN(n4050) );
  NAND2_X1 U3668 ( .A1(n2881), .A2(n3490), .ZN(n4055) );
  NAND2_X1 U3669 ( .A1(n3521), .A2(n4055), .ZN(n2823) );
  NAND2_X1 U3670 ( .A1(n3735), .A2(n3701), .ZN(n4052) );
  NAND2_X1 U3671 ( .A1(n3717), .A2(n4104), .ZN(n3677) );
  NAND2_X1 U3672 ( .A1(n3660), .A2(n3256), .ZN(n3672) );
  NAND2_X1 U3673 ( .A1(n3677), .A2(n3672), .ZN(n2826) );
  INV_X1 U3674 ( .A(n3649), .ZN(n2824) );
  NOR2_X1 U3675 ( .A1(n2826), .A2(n2824), .ZN(n4056) );
  NAND2_X1 U3676 ( .A1(n3650), .A2(n4056), .ZN(n2828) );
  NAND2_X1 U3677 ( .A1(n3652), .A2(n3714), .ZN(n3674) );
  AND2_X1 U3678 ( .A1(n3674), .A2(n3647), .ZN(n2825) );
  OR2_X1 U3679 ( .A1(n2826), .A2(n2825), .ZN(n2827) );
  NAND2_X1 U3680 ( .A1(n3686), .A2(n3780), .ZN(n3676) );
  AND2_X1 U3681 ( .A1(n2827), .A2(n3676), .ZN(n4058) );
  NAND2_X1 U3682 ( .A1(n4456), .A2(n3782), .ZN(n3950) );
  NAND2_X1 U3683 ( .A1(n4474), .A2(n4436), .ZN(n3949) );
  NAND2_X1 U3684 ( .A1(n3950), .A2(n3949), .ZN(n4469) );
  NAND2_X1 U3685 ( .A1(n4466), .A2(n3950), .ZN(n4438) );
  INV_X1 U3686 ( .A(n4450), .ZN(n4015) );
  NAND2_X1 U3687 ( .A1(n4423), .A2(n3910), .ZN(n4066) );
  AND2_X1 U3688 ( .A1(n4412), .A2(n4066), .ZN(n3955) );
  NAND2_X1 U3689 ( .A1(n4439), .A2(n3955), .ZN(n4354) );
  NAND2_X1 U3690 ( .A1(n4398), .A2(n4388), .ZN(n3986) );
  AND2_X1 U3691 ( .A1(n3986), .A2(n4378), .ZN(n4356) );
  NAND2_X1 U3692 ( .A1(n4437), .A2(n4427), .ZN(n4376) );
  NAND2_X1 U3693 ( .A1(n4377), .A2(n4376), .ZN(n2832) );
  NAND2_X1 U3694 ( .A1(n4356), .A2(n2832), .ZN(n2834) );
  NAND2_X1 U3695 ( .A1(n2833), .A2(n4382), .ZN(n3987) );
  NAND2_X1 U3696 ( .A1(n2834), .A2(n3987), .ZN(n4355) );
  NOR2_X1 U3697 ( .A1(n3826), .A2(n4369), .ZN(n2835) );
  NOR2_X1 U3698 ( .A1(n4355), .A2(n2835), .ZN(n4070) );
  NAND2_X1 U3699 ( .A1(n4354), .A2(n4070), .ZN(n2838) );
  INV_X1 U3700 ( .A(n4356), .ZN(n2837) );
  AND2_X1 U3701 ( .A1(n3826), .A2(n4369), .ZN(n2836) );
  AOI21_X1 U3702 ( .B1(n4070), .B2(n2837), .A(n2836), .ZN(n3957) );
  NAND2_X1 U3703 ( .A1(n2838), .A2(n3957), .ZN(n4298) );
  NAND2_X1 U3704 ( .A1(n4362), .A2(n3829), .ZN(n4300) );
  AND2_X1 U3705 ( .A1(n4302), .A2(n4300), .ZN(n4072) );
  NAND2_X1 U3706 ( .A1(n4298), .A2(n4072), .ZN(n2841) );
  NAND2_X1 U3707 ( .A1(n4326), .A2(n4313), .ZN(n3993) );
  NAND2_X1 U3708 ( .A1(n3993), .A2(n2839), .ZN(n4077) );
  AND2_X1 U3709 ( .A1(n4327), .A2(n2882), .ZN(n4299) );
  AND2_X1 U3710 ( .A1(n4302), .A2(n4299), .ZN(n2840) );
  NOR2_X1 U3711 ( .A1(n4077), .A2(n2840), .ZN(n3959) );
  OR2_X1 U3712 ( .A1(n4306), .A2(n4290), .ZN(n3992) );
  INV_X1 U3713 ( .A(n4326), .ZN(n4284) );
  NAND2_X1 U3714 ( .A1(n4284), .A2(n3070), .ZN(n4280) );
  AND2_X1 U3715 ( .A1(n3992), .A2(n4280), .ZN(n4075) );
  INV_X1 U3716 ( .A(n4261), .ZN(n2842) );
  INV_X1 U3717 ( .A(n3843), .ZN(n4272) );
  NAND2_X1 U3718 ( .A1(n4286), .A2(n4272), .ZN(n4017) );
  NAND2_X1 U3719 ( .A1(n4306), .A2(n4290), .ZN(n4260) );
  NAND2_X1 U3720 ( .A1(n4017), .A2(n4260), .ZN(n3961) );
  OR2_X1 U3721 ( .A1(n4286), .A2(n4272), .ZN(n4018) );
  OAI21_X1 U3722 ( .B1(n2842), .B2(n3961), .A(n4018), .ZN(n2843) );
  XNOR2_X1 U3723 ( .A(n2843), .B(n4020), .ZN(n2855) );
  INV_X1 U3724 ( .A(n2884), .ZN(n4592) );
  NAND2_X1 U3725 ( .A1(n4592), .A2(n4591), .ZN(n4092) );
  NAND2_X1 U3726 ( .A1(n2895), .A2(n4593), .ZN(n2844) );
  INV_X1 U3727 ( .A(REG3_REG_27__SCAN_IN), .ZN(n3167) );
  NAND2_X1 U3728 ( .A1(n2845), .A2(n3167), .ZN(n2846) );
  NAND2_X1 U3729 ( .A1(n3109), .A2(n2846), .ZN(n4246) );
  INV_X1 U3730 ( .A(REG1_REG_27__SCAN_IN), .ZN(n4798) );
  NAND2_X1 U3731 ( .A1(n3964), .A2(REG2_REG_27__SCAN_IN), .ZN(n2848) );
  NAND2_X1 U3732 ( .A1(n2591), .A2(REG0_REG_27__SCAN_IN), .ZN(n2847) );
  OAI211_X1 U3733 ( .C1(n3153), .C2(n4798), .A(n2848), .B(n2847), .ZN(n2849)
         );
  INV_X1 U3734 ( .A(n2849), .ZN(n2850) );
  INV_X1 U3735 ( .A(n4286), .ZN(n3921) );
  INV_X1 U3736 ( .A(n2895), .ZN(n2852) );
  OAI22_X1 U3737 ( .A1(n3921), .A2(n4462), .B1(n4422), .B2(n3174), .ZN(n2853)
         );
  AOI21_X1 U3738 ( .B1(n4418), .B2(n3440), .A(n2853), .ZN(n2854) );
  OAI21_X1 U3739 ( .B1(n2855), .B2(n4468), .A(n2854), .ZN(n4256) );
  AOI21_X1 U3740 ( .B1(n4251), .B2(n4545), .A(n4256), .ZN(n4502) );
  NAND2_X1 U3741 ( .A1(n2857), .A2(n4840), .ZN(n2858) );
  NAND3_X1 U3742 ( .A1(n2878), .A2(B_REG_SCAN_IN), .A3(n2863), .ZN(n2862) );
  INV_X1 U3743 ( .A(n2878), .ZN(n3249) );
  NAND2_X1 U3744 ( .A1(n3249), .A2(n4976), .ZN(n2861) );
  INV_X1 U3745 ( .A(n2856), .ZN(n2877) );
  NAND2_X1 U3746 ( .A1(n2877), .A2(n2863), .ZN(n4727) );
  NAND2_X1 U3747 ( .A1(n3181), .A2(n4727), .ZN(n2876) );
  NAND2_X1 U3748 ( .A1(n2884), .A2(n4094), .ZN(n2864) );
  NOR2_X1 U3749 ( .A1(n3180), .A2(n3147), .ZN(n2875) );
  INV_X1 U3750 ( .A(D_REG_22__SCAN_IN), .ZN(n4851) );
  INV_X1 U3751 ( .A(D_REG_18__SCAN_IN), .ZN(n4876) );
  INV_X1 U3752 ( .A(D_REG_11__SCAN_IN), .ZN(n4893) );
  INV_X1 U3753 ( .A(D_REG_29__SCAN_IN), .ZN(n4896) );
  NAND4_X1 U3754 ( .A1(n4851), .A2(n4876), .A3(n4893), .A4(n4896), .ZN(n2865)
         );
  NOR4_X1 U3755 ( .A1(D_REG_13__SCAN_IN), .A2(D_REG_7__SCAN_IN), .A3(
        D_REG_8__SCAN_IN), .A4(n2865), .ZN(n4751) );
  NOR4_X1 U3756 ( .A1(D_REG_10__SCAN_IN), .A2(D_REG_17__SCAN_IN), .A3(
        D_REG_3__SCAN_IN), .A4(D_REG_2__SCAN_IN), .ZN(n2867) );
  NOR3_X1 U3757 ( .A1(D_REG_31__SCAN_IN), .A2(D_REG_9__SCAN_IN), .A3(
        D_REG_25__SCAN_IN), .ZN(n2866) );
  NAND3_X1 U3758 ( .A1(n4751), .A2(n2867), .A3(n2866), .ZN(n2873) );
  NOR4_X1 U3759 ( .A1(D_REG_12__SCAN_IN), .A2(D_REG_14__SCAN_IN), .A3(
        D_REG_20__SCAN_IN), .A4(D_REG_16__SCAN_IN), .ZN(n2871) );
  NOR4_X1 U3760 ( .A1(D_REG_6__SCAN_IN), .A2(D_REG_4__SCAN_IN), .A3(
        D_REG_5__SCAN_IN), .A4(D_REG_15__SCAN_IN), .ZN(n2870) );
  NOR4_X1 U3761 ( .A1(D_REG_28__SCAN_IN), .A2(D_REG_26__SCAN_IN), .A3(
        D_REG_27__SCAN_IN), .A4(D_REG_30__SCAN_IN), .ZN(n2869) );
  NOR4_X1 U3762 ( .A1(D_REG_19__SCAN_IN), .A2(D_REG_24__SCAN_IN), .A3(
        D_REG_21__SCAN_IN), .A4(D_REG_23__SCAN_IN), .ZN(n2868) );
  NAND4_X1 U3763 ( .A1(n2871), .A2(n2870), .A3(n2869), .A4(n2868), .ZN(n2872)
         );
  NOR2_X1 U3764 ( .A1(n2873), .A2(n2872), .ZN(n2874) );
  NAND2_X1 U3765 ( .A1(n2878), .A2(n2877), .ZN(n3254) );
  MUX2_X1 U3766 ( .A(n4795), .B(n4502), .S(n4717), .Z(n2887) );
  NAND2_X1 U3767 ( .A1(n3505), .A2(n3400), .ZN(n3399) );
  NAND2_X1 U3768 ( .A1(n4444), .A2(n4435), .ZN(n4426) );
  INV_X1 U3769 ( .A(n4271), .ZN(n2883) );
  OAI21_X1 U3770 ( .B1(n2883), .B2(n3174), .A(n2227), .ZN(n4505) );
  NAND2_X1 U3771 ( .A1(n2887), .A2(n2886), .ZN(U3512) );
  NAND2_X1 U3772 ( .A1(n2129), .A2(n4111), .ZN(n2890) );
  NAND2_X1 U3773 ( .A1(n2923), .A2(n3296), .ZN(n2889) );
  NAND2_X1 U3774 ( .A1(n2890), .A2(n2889), .ZN(n3297) );
  NAND2_X1 U3775 ( .A1(n3296), .A2(n2898), .ZN(n2891) );
  OAI21_X2 U3776 ( .B1(n3790), .B2(n2906), .A(n2891), .ZN(n3298) );
  NAND2_X1 U3777 ( .A1(n3297), .A2(n3298), .ZN(n2894) );
  OR2_X1 U3778 ( .A1(n2888), .A2(n2892), .ZN(n2893) );
  NAND2_X1 U3779 ( .A1(n2894), .A2(n2893), .ZN(n3300) );
  NAND2_X4 U3780 ( .A1(n3185), .A2(n3140), .ZN(n3117) );
  NOR2_X1 U3781 ( .A1(n3298), .A2(n3117), .ZN(n2896) );
  OR2_X2 U3782 ( .A1(n3300), .A2(n2896), .ZN(n3794) );
  AOI22_X1 U3783 ( .A1(n2908), .A2(n2601), .B1(n2923), .B2(n3455), .ZN(n2902)
         );
  INV_X1 U3784 ( .A(n2902), .ZN(n2901) );
  NAND2_X1 U3785 ( .A1(n3455), .A2(n2898), .ZN(n2899) );
  NAND2_X1 U3786 ( .A1(n3794), .A2(n3795), .ZN(n3793) );
  OR2_X1 U3787 ( .A1(n2903), .A2(n2902), .ZN(n2904) );
  NAND2_X1 U3788 ( .A1(n3793), .A2(n2904), .ZN(n3337) );
  INV_X1 U3789 ( .A(n3337), .ZN(n2911) );
  NAND2_X1 U3790 ( .A1(n3355), .A2(n2898), .ZN(n2905) );
  OAI21_X1 U3791 ( .B1(n3789), .B2(n2906), .A(n2905), .ZN(n2907) );
  XNOR2_X1 U3792 ( .A(n2907), .B(n2930), .ZN(n2913) );
  AOI22_X1 U3793 ( .A1(n2908), .A2(n2909), .B1(n2923), .B2(n3355), .ZN(n2912)
         );
  XNOR2_X1 U3794 ( .A(n2913), .B(n2912), .ZN(n3338) );
  INV_X1 U3795 ( .A(n3338), .ZN(n2910) );
  NAND2_X1 U3796 ( .A1(n2913), .A2(n2912), .ZN(n2914) );
  NAND2_X1 U3797 ( .A1(n3507), .A2(n3104), .ZN(n2915) );
  OAI21_X1 U3798 ( .B1(n3392), .B2(n3116), .A(n2915), .ZN(n2916) );
  XNOR2_X1 U3799 ( .A(n2916), .B(n3117), .ZN(n2917) );
  AOI22_X1 U3800 ( .A1(n2125), .A2(n4110), .B1(n3142), .B2(n3507), .ZN(n2918)
         );
  XNOR2_X1 U3801 ( .A(n2917), .B(n2918), .ZN(n3366) );
  INV_X1 U3802 ( .A(n2917), .ZN(n2919) );
  NAND2_X1 U3803 ( .A1(n2919), .A2(n2918), .ZN(n2920) );
  OAI22_X1 U3804 ( .A1(n3400), .A2(n2921), .B1(n3116), .B2(n3367), .ZN(n2922)
         );
  XNOR2_X1 U3805 ( .A(n2922), .B(n3117), .ZN(n2928) );
  NAND2_X1 U3806 ( .A1(n2125), .A2(n3535), .ZN(n2925) );
  NAND2_X1 U3807 ( .A1(n3396), .A2(n3142), .ZN(n2924) );
  NAND2_X1 U3808 ( .A1(n2925), .A2(n2924), .ZN(n2927) );
  XNOR2_X1 U3809 ( .A(n2928), .B(n2927), .ZN(n3373) );
  INV_X1 U3810 ( .A(n3373), .ZN(n2926) );
  NAND2_X1 U3811 ( .A1(n2928), .A2(n2927), .ZN(n2929) );
  NAND2_X1 U3812 ( .A1(n3374), .A2(n2929), .ZN(n3409) );
  OAI22_X1 U3813 ( .A1(n3538), .A2(n2921), .B1(n3116), .B2(n2626), .ZN(n2931)
         );
  XNOR2_X1 U3814 ( .A(n2931), .B(n2930), .ZN(n2934) );
  NAND2_X1 U3815 ( .A1(n2125), .A2(n4108), .ZN(n2933) );
  NAND2_X1 U3816 ( .A1(n3542), .A2(n3142), .ZN(n2932) );
  NAND2_X1 U3817 ( .A1(n2933), .A2(n2932), .ZN(n2935) );
  XNOR2_X1 U3818 ( .A(n2934), .B(n2935), .ZN(n3408) );
  INV_X1 U3819 ( .A(n2934), .ZN(n2936) );
  NAND2_X1 U3820 ( .A1(n2936), .A2(n2935), .ZN(n2937) );
  NAND2_X1 U3821 ( .A1(n2126), .A2(n3589), .ZN(n2939) );
  NAND2_X1 U3822 ( .A1(n3142), .A2(n3588), .ZN(n2938) );
  NAND2_X1 U3823 ( .A1(n2939), .A2(n2938), .ZN(n3416) );
  NAND2_X1 U3824 ( .A1(n3588), .A2(n3104), .ZN(n2940) );
  OAI21_X1 U3825 ( .B1(n2648), .B2(n3116), .A(n2940), .ZN(n2941) );
  XNOR2_X1 U3826 ( .A(n2941), .B(n3117), .ZN(n3415) );
  NAND2_X1 U3827 ( .A1(n3418), .A2(n3416), .ZN(n2979) );
  OAI22_X1 U3828 ( .A1(n3580), .A2(n2921), .B1(n3116), .B2(n3554), .ZN(n2942)
         );
  XNOR2_X1 U3829 ( .A(n2942), .B(n2930), .ZN(n2967) );
  NAND2_X1 U3830 ( .A1(n2126), .A2(n4107), .ZN(n2944) );
  NAND2_X1 U3831 ( .A1(n3581), .A2(n3142), .ZN(n2943) );
  NAND2_X1 U3832 ( .A1(n2944), .A2(n2943), .ZN(n2968) );
  XNOR2_X1 U3833 ( .A(n2967), .B(n2968), .ZN(n3549) );
  NAND2_X1 U3834 ( .A1(n3735), .A2(n3104), .ZN(n2945) );
  AOI22_X1 U3835 ( .A1(n2126), .A2(n3490), .B1(n3142), .B2(n3735), .ZN(n2956)
         );
  INV_X1 U3836 ( .A(n2959), .ZN(n2954) );
  OAI22_X1 U3837 ( .A1(n3557), .A2(n2921), .B1(n3116), .B2(n3467), .ZN(n2946)
         );
  XNOR2_X1 U3838 ( .A(n2946), .B(n3117), .ZN(n2966) );
  INV_X1 U3839 ( .A(n2966), .ZN(n2950) );
  NAND2_X1 U3840 ( .A1(n2126), .A2(n3703), .ZN(n2948) );
  NAND2_X1 U3841 ( .A1(n3434), .A2(n3142), .ZN(n2947) );
  NAND2_X1 U3842 ( .A1(n2948), .A2(n2947), .ZN(n2965) );
  INV_X1 U3843 ( .A(n2965), .ZN(n2949) );
  NAND2_X1 U3844 ( .A1(n2950), .A2(n2949), .ZN(n3698) );
  NAND2_X1 U3845 ( .A1(n3473), .A2(n3104), .ZN(n2951) );
  OAI21_X1 U3846 ( .B1(n2952), .B2(n3116), .A(n2951), .ZN(n2953) );
  AOI22_X1 U3847 ( .A1(n2129), .A2(n4106), .B1(n3142), .B2(n3473), .ZN(n2961)
         );
  AND2_X1 U3848 ( .A1(n3698), .A2(n2960), .ZN(n3722) );
  INV_X1 U3849 ( .A(n2955), .ZN(n2958) );
  INV_X1 U3850 ( .A(n2956), .ZN(n2957) );
  NAND2_X1 U3851 ( .A1(n2958), .A2(n2957), .ZN(n2964) );
  XNOR2_X1 U3852 ( .A(n2962), .B(n2961), .ZN(n3700) );
  OR2_X1 U3853 ( .A1(n2963), .A2(n3700), .ZN(n3723) );
  OR2_X1 U3854 ( .A1(n2959), .A2(n3723), .ZN(n3728) );
  AND2_X1 U3855 ( .A1(n2964), .A2(n3728), .ZN(n2983) );
  INV_X1 U3856 ( .A(n3726), .ZN(n2972) );
  AND2_X1 U3857 ( .A1(n2966), .A2(n2965), .ZN(n3696) );
  INV_X1 U3858 ( .A(n3696), .ZN(n2970) );
  INV_X1 U3859 ( .A(n2967), .ZN(n2969) );
  NAND2_X1 U3860 ( .A1(n2969), .A2(n2968), .ZN(n3550) );
  AND2_X1 U3861 ( .A1(n2970), .A2(n3550), .ZN(n2971) );
  AND2_X1 U3862 ( .A1(n2983), .A2(n2984), .ZN(n2973) );
  NAND2_X1 U3863 ( .A1(n2125), .A2(n4105), .ZN(n2976) );
  NAND2_X1 U3864 ( .A1(n3616), .A2(n3142), .ZN(n2975) );
  NAND2_X1 U3865 ( .A1(n2976), .A2(n2975), .ZN(n3487) );
  OAI22_X1 U3866 ( .A1(n2977), .A2(n2921), .B1(n3116), .B2(n3733), .ZN(n2978)
         );
  XNOR2_X1 U3867 ( .A(n2978), .B(n3117), .ZN(n3486) );
  AND2_X1 U3868 ( .A1(n2979), .A2(n2983), .ZN(n2982) );
  AND2_X1 U3869 ( .A1(n2984), .A2(n2980), .ZN(n2981) );
  NAND2_X1 U3870 ( .A1(n2982), .A2(n2981), .ZN(n2988) );
  INV_X1 U3871 ( .A(n2983), .ZN(n2986) );
  NAND2_X1 U3872 ( .A1(n2988), .A2(n2987), .ZN(n2989) );
  NAND2_X1 U3873 ( .A1(n3652), .A2(n3104), .ZN(n2991) );
  NAND2_X1 U3874 ( .A1(n3142), .A2(n3256), .ZN(n2990) );
  NAND2_X1 U3875 ( .A1(n2991), .A2(n2990), .ZN(n2992) );
  XNOR2_X1 U3876 ( .A(n2992), .B(n3117), .ZN(n2995) );
  NAND2_X1 U3877 ( .A1(n3652), .A2(n3142), .ZN(n2994) );
  NAND2_X1 U3878 ( .A1(n2126), .A2(n3256), .ZN(n2993) );
  NAND2_X1 U3879 ( .A1(n2994), .A2(n2993), .ZN(n2996) );
  AND2_X1 U3880 ( .A1(n2995), .A2(n2996), .ZN(n3625) );
  INV_X1 U3881 ( .A(n2995), .ZN(n2998) );
  INV_X1 U3882 ( .A(n2996), .ZN(n2997) );
  NAND2_X1 U3883 ( .A1(n2998), .A2(n2997), .ZN(n3624) );
  OAI22_X1 U3884 ( .A1(n3717), .A2(n2921), .B1(n3780), .B2(n3116), .ZN(n2999)
         );
  XNOR2_X1 U3885 ( .A(n2999), .B(n2930), .ZN(n3711) );
  NAND2_X1 U3886 ( .A1(n3710), .A2(n3711), .ZN(n3002) );
  OR2_X1 U3887 ( .A1(n3717), .A2(n3116), .ZN(n3001) );
  NAND2_X1 U3888 ( .A1(n4104), .A2(n2126), .ZN(n3000) );
  NAND2_X1 U3889 ( .A1(n3001), .A2(n3000), .ZN(n3712) );
  NAND2_X1 U3890 ( .A1(n3643), .A2(n3104), .ZN(n3005) );
  OAI21_X1 U3891 ( .B1(n4463), .B2(n3116), .A(n3005), .ZN(n3006) );
  XNOR2_X1 U3892 ( .A(n3006), .B(n3117), .ZN(n3017) );
  NAND2_X1 U3893 ( .A1(n3643), .A2(n3142), .ZN(n3007) );
  OAI21_X1 U3894 ( .B1(n4463), .B2(n3051), .A(n3007), .ZN(n3018) );
  AND2_X1 U3895 ( .A1(n3017), .A2(n3018), .ZN(n3777) );
  OAI22_X1 U3896 ( .A1(n4435), .A2(n2921), .B1(n4465), .B2(n3116), .ZN(n3009)
         );
  XNOR2_X1 U3897 ( .A(n3009), .B(n3117), .ZN(n3023) );
  INV_X1 U3898 ( .A(n3023), .ZN(n3013) );
  OR2_X1 U3899 ( .A1(n4435), .A2(n3116), .ZN(n3011) );
  NAND2_X1 U3900 ( .A1(n4416), .A2(n2126), .ZN(n3010) );
  NAND2_X1 U3901 ( .A1(n3011), .A2(n3010), .ZN(n3022) );
  INV_X1 U3902 ( .A(n3022), .ZN(n3012) );
  NAND2_X1 U3903 ( .A1(n3013), .A2(n3012), .ZN(n3849) );
  NAND2_X1 U3904 ( .A1(n4474), .A2(n3104), .ZN(n3015) );
  NAND2_X1 U3905 ( .A1(n3782), .A2(n3142), .ZN(n3014) );
  NAND2_X1 U3906 ( .A1(n3015), .A2(n3014), .ZN(n3016) );
  XNOR2_X1 U3907 ( .A(n3016), .B(n2930), .ZN(n3853) );
  AOI22_X1 U3908 ( .A1(n4474), .A2(n3142), .B1(n2126), .B2(n3782), .ZN(n3934)
         );
  INV_X1 U3909 ( .A(n3017), .ZN(n3020) );
  INV_X1 U3910 ( .A(n3018), .ZN(n3019) );
  AOI21_X1 U3911 ( .B1(n3853), .B2(n3934), .A(n3850), .ZN(n3021) );
  AND2_X1 U3912 ( .A1(n3849), .A2(n3021), .ZN(n3026) );
  NAND2_X1 U3913 ( .A1(n3023), .A2(n3022), .ZN(n3848) );
  OAI21_X1 U3914 ( .B1(n3934), .B2(n3853), .A(n3848), .ZN(n3024) );
  AND2_X1 U3915 ( .A1(n3024), .A2(n3849), .ZN(n3025) );
  NAND2_X1 U3916 ( .A1(n4427), .A2(n3104), .ZN(n3027) );
  OAI21_X1 U3917 ( .B1(n4437), .B2(n3116), .A(n3027), .ZN(n3028) );
  XNOR2_X1 U3918 ( .A(n3028), .B(n3117), .ZN(n3031) );
  OR2_X1 U3919 ( .A1(n4437), .A2(n3051), .ZN(n3030) );
  NAND2_X1 U3920 ( .A1(n4427), .A2(n3142), .ZN(n3029) );
  NAND2_X1 U3921 ( .A1(n3030), .A2(n3029), .ZN(n3032) );
  NAND2_X1 U3922 ( .A1(n3031), .A2(n3032), .ZN(n3865) );
  INV_X1 U3923 ( .A(n3031), .ZN(n3034) );
  INV_X1 U3924 ( .A(n3032), .ZN(n3033) );
  NAND2_X1 U3925 ( .A1(n3034), .A2(n3033), .ZN(n3864) );
  NOR2_X1 U3926 ( .A1(n4405), .A2(n3116), .ZN(n3035) );
  AOI21_X1 U3927 ( .B1(n4419), .B2(n2125), .A(n3035), .ZN(n3908) );
  NAND2_X1 U3928 ( .A1(n4398), .A2(n3142), .ZN(n3037) );
  NAND2_X1 U3929 ( .A1(n4382), .A2(n3104), .ZN(n3036) );
  NAND2_X1 U3930 ( .A1(n3037), .A2(n3036), .ZN(n3038) );
  XNOR2_X1 U3931 ( .A(n3038), .B(n2930), .ZN(n3040) );
  AND2_X1 U3932 ( .A1(n3142), .A2(n4382), .ZN(n3039) );
  AOI21_X1 U3933 ( .B1(n4398), .B2(n2126), .A(n3039), .ZN(n3041) );
  NAND2_X1 U3934 ( .A1(n3040), .A2(n3041), .ZN(n3823) );
  INV_X1 U3935 ( .A(n3040), .ZN(n3043) );
  INV_X1 U3936 ( .A(n3041), .ZN(n3042) );
  NAND2_X1 U3937 ( .A1(n3043), .A2(n3042), .ZN(n3044) );
  NAND2_X1 U3938 ( .A1(n3823), .A2(n3044), .ZN(n3814) );
  NAND2_X1 U3939 ( .A1(n3906), .A2(n3908), .ZN(n3048) );
  NAND2_X1 U3940 ( .A1(n4419), .A2(n3142), .ZN(n3046) );
  NAND2_X1 U3941 ( .A1(n4397), .A2(n3104), .ZN(n3045) );
  NAND2_X1 U3942 ( .A1(n3046), .A2(n3045), .ZN(n3047) );
  XNOR2_X1 U3943 ( .A(n3047), .B(n3117), .ZN(n3907) );
  NAND2_X1 U3944 ( .A1(n3048), .A2(n3907), .ZN(n3810) );
  NAND2_X1 U3945 ( .A1(n3049), .A2(n3810), .ZN(n3811) );
  OAI22_X1 U3946 ( .A1(n4385), .A2(n3116), .B1(n2921), .B2(n4369), .ZN(n3050)
         );
  XNOR2_X1 U3947 ( .A(n3050), .B(n3117), .ZN(n3057) );
  INV_X1 U3948 ( .A(n3057), .ZN(n3055) );
  OR2_X1 U3949 ( .A1(n4385), .A2(n3051), .ZN(n3053) );
  NAND2_X1 U3950 ( .A1(n3142), .A2(n4360), .ZN(n3052) );
  NAND2_X1 U3951 ( .A1(n3053), .A2(n3052), .ZN(n3056) );
  INV_X1 U3952 ( .A(n3056), .ZN(n3054) );
  NAND2_X1 U3953 ( .A1(n3055), .A2(n3054), .ZN(n3886) );
  AND2_X1 U3954 ( .A1(n3823), .A2(n3886), .ZN(n3059) );
  NAND2_X1 U3955 ( .A1(n3057), .A2(n3056), .ZN(n3887) );
  NAND2_X1 U3956 ( .A1(n4327), .A2(n3142), .ZN(n3061) );
  NAND2_X1 U3957 ( .A1(n3104), .A2(n3829), .ZN(n3060) );
  NAND2_X1 U3958 ( .A1(n3061), .A2(n3060), .ZN(n3062) );
  XNOR2_X1 U3959 ( .A(n3062), .B(n2930), .ZN(n3064) );
  NOR2_X1 U3960 ( .A1(n3116), .A2(n2882), .ZN(n3063) );
  AOI21_X1 U3961 ( .B1(n4327), .B2(n2126), .A(n3063), .ZN(n3065) );
  INV_X1 U3962 ( .A(n3064), .ZN(n3067) );
  INV_X1 U3963 ( .A(n3065), .ZN(n3066) );
  NAND2_X1 U3964 ( .A1(n3067), .A2(n3066), .ZN(n3822) );
  OAI22_X1 U3965 ( .A1(n4341), .A2(n3116), .B1(n2921), .B2(n3069), .ZN(n3068)
         );
  XNOR2_X1 U3966 ( .A(n3068), .B(n3117), .ZN(n3075) );
  OAI22_X1 U3967 ( .A1(n4341), .A2(n3051), .B1(n3116), .B2(n3069), .ZN(n3076)
         );
  XNOR2_X1 U3968 ( .A(n3075), .B(n3076), .ZN(n3898) );
  NAND2_X1 U3969 ( .A1(n4326), .A2(n3142), .ZN(n3072) );
  NAND2_X1 U3970 ( .A1(n3104), .A2(n3070), .ZN(n3071) );
  NAND2_X1 U3971 ( .A1(n3072), .A2(n3071), .ZN(n3073) );
  XNOR2_X1 U3972 ( .A(n3073), .B(n3117), .ZN(n3088) );
  NOR2_X1 U3973 ( .A1(n3116), .A2(n4313), .ZN(n3074) );
  AOI21_X1 U3974 ( .B1(n4326), .B2(n2125), .A(n3074), .ZN(n3086) );
  XNOR2_X1 U3975 ( .A(n3088), .B(n3086), .ZN(n3801) );
  INV_X1 U3976 ( .A(n3075), .ZN(n3078) );
  INV_X1 U3977 ( .A(n3076), .ZN(n3077) );
  NAND2_X1 U3978 ( .A1(n3078), .A2(n3077), .ZN(n3800) );
  AND2_X1 U3979 ( .A1(n3801), .A2(n3800), .ZN(n3079) );
  NAND2_X1 U3980 ( .A1(n4286), .A2(n3142), .ZN(n3081) );
  NAND2_X1 U3981 ( .A1(n3104), .A2(n3843), .ZN(n3080) );
  NAND2_X1 U3982 ( .A1(n3081), .A2(n3080), .ZN(n3082) );
  XNOR2_X1 U3983 ( .A(n3082), .B(n3117), .ZN(n3840) );
  NAND2_X1 U3984 ( .A1(n4286), .A2(n2126), .ZN(n3084) );
  NAND2_X1 U3985 ( .A1(n3142), .A2(n3843), .ZN(n3083) );
  NAND2_X1 U3986 ( .A1(n3084), .A2(n3083), .ZN(n3839) );
  NAND2_X1 U3987 ( .A1(n3840), .A2(n3839), .ZN(n3838) );
  OAI22_X1 U3988 ( .A1(n4265), .A2(n3116), .B1(n2921), .B2(n4290), .ZN(n3085)
         );
  XNOR2_X1 U3989 ( .A(n3085), .B(n3117), .ZN(n3875) );
  INV_X1 U3990 ( .A(n3086), .ZN(n3087) );
  NAND2_X1 U3991 ( .A1(n3088), .A2(n3087), .ZN(n3836) );
  INV_X1 U3992 ( .A(n3836), .ZN(n3090) );
  NOR2_X1 U3993 ( .A1(n3116), .A2(n4290), .ZN(n3089) );
  AOI21_X1 U3994 ( .B1(n4306), .B2(n2125), .A(n3089), .ZN(n3835) );
  NAND2_X1 U3995 ( .A1(n3835), .A2(n3836), .ZN(n3833) );
  OAI21_X1 U3996 ( .B1(n3875), .B2(n3090), .A(n3833), .ZN(n3091) );
  INV_X1 U3997 ( .A(n3835), .ZN(n3092) );
  OAI21_X1 U3998 ( .B1(n3875), .B2(n3092), .A(n3839), .ZN(n3096) );
  INV_X1 U3999 ( .A(n3840), .ZN(n3095) );
  INV_X1 U4000 ( .A(n3875), .ZN(n3094) );
  NOR2_X1 U4001 ( .A1(n3839), .A2(n3092), .ZN(n3093) );
  AOI22_X1 U4002 ( .A1(n3096), .A2(n3095), .B1(n3094), .B2(n3093), .ZN(n3097)
         );
  OAI22_X1 U4003 ( .A1(n4234), .A2(n3116), .B1(n2921), .B2(n3174), .ZN(n3098)
         );
  XNOR2_X1 U4004 ( .A(n3098), .B(n2930), .ZN(n3103) );
  INV_X1 U4005 ( .A(n3103), .ZN(n3101) );
  NOR2_X1 U4006 ( .A1(n3116), .A2(n3174), .ZN(n3099) );
  AOI21_X1 U4007 ( .B1(n4267), .B2(n2125), .A(n3099), .ZN(n3102) );
  INV_X1 U4008 ( .A(n3102), .ZN(n3100) );
  NAND2_X1 U4009 ( .A1(n3101), .A2(n3100), .ZN(n3917) );
  NAND2_X1 U4010 ( .A1(n3440), .A2(n3142), .ZN(n3106) );
  NAND2_X1 U4011 ( .A1(n3104), .A2(n3189), .ZN(n3105) );
  NAND2_X1 U4012 ( .A1(n3106), .A2(n3105), .ZN(n3107) );
  XNOR2_X1 U4013 ( .A(n3107), .B(n3117), .ZN(n3123) );
  NOR2_X1 U4014 ( .A1(n3116), .A2(n4243), .ZN(n3108) );
  AOI21_X1 U4015 ( .B1(n3440), .B2(n2126), .A(n3108), .ZN(n3121) );
  XNOR2_X1 U4016 ( .A(n3123), .B(n3121), .ZN(n3163) );
  INV_X1 U4017 ( .A(n3130), .ZN(n3129) );
  INV_X1 U4018 ( .A(REG3_REG_28__SCAN_IN), .ZN(n3149) );
  NAND2_X1 U4019 ( .A1(n3109), .A2(n3149), .ZN(n3110) );
  NAND2_X1 U4020 ( .A1(n4226), .A2(n3155), .ZN(n3115) );
  INV_X1 U4021 ( .A(REG1_REG_28__SCAN_IN), .ZN(n4806) );
  NAND2_X1 U4022 ( .A1(n3964), .A2(REG2_REG_28__SCAN_IN), .ZN(n3112) );
  NAND2_X1 U4023 ( .A1(n2591), .A2(REG0_REG_28__SCAN_IN), .ZN(n3111) );
  OAI211_X1 U4024 ( .C1(n3153), .C2(n4806), .A(n3112), .B(n3111), .ZN(n3113)
         );
  INV_X1 U4025 ( .A(n3113), .ZN(n3114) );
  AND2_X2 U4026 ( .A1(n3115), .A2(n3114), .ZN(n3200) );
  OAI22_X1 U4027 ( .A1(n3200), .A2(n3116), .B1(n2921), .B2(n3217), .ZN(n3118)
         );
  XNOR2_X1 U4028 ( .A(n3118), .B(n3117), .ZN(n3120) );
  OAI22_X1 U4029 ( .A1(n3200), .A2(n3051), .B1(n3116), .B2(n3217), .ZN(n3119)
         );
  XNOR2_X1 U4030 ( .A(n3120), .B(n3119), .ZN(n3133) );
  INV_X1 U4031 ( .A(n3133), .ZN(n3128) );
  INV_X1 U4032 ( .A(n3121), .ZN(n3122) );
  NAND2_X1 U4033 ( .A1(n3123), .A2(n3122), .ZN(n3131) );
  NAND3_X1 U4034 ( .A1(n3182), .A2(n3227), .A3(n3181), .ZN(n3156) );
  OR2_X1 U4035 ( .A1(n3156), .A2(n3146), .ZN(n3145) );
  INV_X1 U4036 ( .A(n3125), .ZN(n3127) );
  NAND2_X1 U4037 ( .A1(n2885), .A2(n4593), .ZN(n3126) );
  NAND3_X1 U4038 ( .A1(n4422), .A2(n3127), .A3(n3126), .ZN(n3134) );
  NAND2_X1 U4039 ( .A1(n3129), .A2(n2146), .ZN(n3162) );
  NAND3_X1 U4040 ( .A1(n3130), .A2(n3888), .A3(n3133), .ZN(n3161) );
  INV_X1 U4041 ( .A(n3131), .ZN(n3132) );
  NAND3_X1 U4042 ( .A1(n3133), .A2(n3888), .A3(n3132), .ZN(n3160) );
  NAND2_X1 U40430 ( .A1(n3134), .A2(n4422), .ZN(n3135) );
  NAND2_X1 U4044 ( .A1(n3156), .A2(n3135), .ZN(n3293) );
  NAND2_X1 U4045 ( .A1(n3136), .A2(n2888), .ZN(n3137) );
  NOR2_X1 U4046 ( .A1(n3138), .A2(n3137), .ZN(n3139) );
  AOI21_X1 U4047 ( .B1(n3293), .B2(n3139), .A(U3149), .ZN(n3144) );
  INV_X1 U4048 ( .A(n3140), .ZN(n3141) );
  NAND3_X1 U4049 ( .A1(n3142), .A2(n4726), .A3(n3141), .ZN(n4097) );
  INV_X1 U4050 ( .A(n4097), .ZN(n3143) );
  AND2_X1 U4051 ( .A1(n3156), .A2(n3143), .ZN(n3292) );
  OR2_X1 U4052 ( .A1(n3145), .A2(n4422), .ZN(n3148) );
  OAI22_X1 U4053 ( .A1(n3941), .A2(n3217), .B1(STATE_REG_SCAN_IN), .B2(n3149), 
        .ZN(n3158) );
  INV_X1 U4054 ( .A(n3150), .ZN(n3203) );
  INV_X1 U4055 ( .A(REG1_REG_29__SCAN_IN), .ZN(n4809) );
  NAND2_X1 U4056 ( .A1(n2591), .A2(REG0_REG_29__SCAN_IN), .ZN(n3152) );
  NAND2_X1 U4057 ( .A1(n3964), .A2(REG2_REG_29__SCAN_IN), .ZN(n3151) );
  OAI211_X1 U4058 ( .C1(n3153), .C2(n4809), .A(n3152), .B(n3151), .ZN(n3154)
         );
  AOI21_X1 U4059 ( .B1(n3203), .B2(n3155), .A(n3154), .ZN(n3971) );
  OAI22_X1 U4060 ( .A1(n3971), .A2(n3923), .B1(n3924), .B2(n3920), .ZN(n3157)
         );
  AOI211_X1 U4061 ( .C1(n4226), .C2(n3943), .A(n3158), .B(n3157), .ZN(n3159)
         );
  NAND3_X1 U4062 ( .A1(n3162), .A2(n3161), .A3(n2368), .ZN(U3217) );
  XNOR2_X1 U4063 ( .A(n3165), .B(n3164), .ZN(n3166) );
  NAND2_X1 U4064 ( .A1(n3166), .A2(n3888), .ZN(n3173) );
  NOR2_X1 U4065 ( .A1(n4246), .A2(n3922), .ZN(n3169) );
  OAI22_X1 U4066 ( .A1(n4234), .A2(n3920), .B1(STATE_REG_SCAN_IN), .B2(n3167), 
        .ZN(n3168) );
  AOI211_X1 U4067 ( .C1(n3189), .C2(n3927), .A(n3169), .B(n3168), .ZN(n3171)
         );
  OR2_X1 U4068 ( .A1(n3200), .A2(n3923), .ZN(n3170) );
  NAND2_X1 U4069 ( .A1(n3173), .A2(n3172), .ZN(U3211) );
  NOR2_X1 U4070 ( .A1(n4234), .A2(n3174), .ZN(n3175) );
  NOR2_X1 U4071 ( .A1(n3440), .A2(n3189), .ZN(n3177) );
  NAND2_X1 U4072 ( .A1(n3200), .A2(n3223), .ZN(n3192) );
  NAND2_X1 U4073 ( .A1(n4239), .A2(n3217), .ZN(n3973) );
  INV_X1 U4074 ( .A(n4022), .ZN(n3178) );
  NAND2_X1 U4075 ( .A1(n3212), .A2(n3178), .ZN(n4493) );
  NAND2_X1 U4076 ( .A1(n4239), .A2(n3223), .ZN(n4491) );
  NAND2_X1 U4077 ( .A1(n4493), .A2(n4491), .ZN(n3179) );
  XNOR2_X1 U4078 ( .A(n3971), .B(n3970), .ZN(n4492) );
  INV_X1 U4079 ( .A(n3180), .ZN(n3294) );
  NAND4_X1 U4080 ( .A1(n3183), .A2(n3182), .A3(n3294), .A4(n3181), .ZN(n3184)
         );
  OR2_X1 U4081 ( .A1(n3185), .A2(n4094), .ZN(n3404) );
  AND2_X1 U4082 ( .A1(n4366), .A2(n3404), .ZN(n3186) );
  NAND2_X1 U4083 ( .A1(n3187), .A2(n4018), .ZN(n3188) );
  INV_X1 U4084 ( .A(n3188), .ZN(n4076) );
  AOI21_X1 U4085 ( .B1(n4076), .B2(n3961), .A(n3974), .ZN(n4082) );
  NAND2_X1 U4086 ( .A1(n3924), .A2(n3189), .ZN(n3214) );
  NAND2_X1 U4087 ( .A1(n3440), .A2(n4243), .ZN(n4080) );
  NAND2_X1 U4088 ( .A1(n3191), .A2(n3190), .ZN(n3213) );
  AND2_X1 U4089 ( .A1(n3192), .A2(n3214), .ZN(n3976) );
  NAND2_X1 U4090 ( .A1(n3213), .A2(n3976), .ZN(n3193) );
  NAND2_X1 U4091 ( .A1(n3193), .A2(n3973), .ZN(n3194) );
  XNOR2_X1 U4092 ( .A(n3194), .B(n4492), .ZN(n3202) );
  NOR2_X1 U4093 ( .A1(n3306), .A2(n4976), .ZN(n3195) );
  NOR2_X1 U4094 ( .A1(n4464), .A2(n3195), .ZN(n4215) );
  NAND2_X1 U4095 ( .A1(n2606), .A2(REG1_REG_30__SCAN_IN), .ZN(n3198) );
  NAND2_X1 U4096 ( .A1(n3964), .A2(REG2_REG_30__SCAN_IN), .ZN(n3197) );
  NAND2_X1 U4097 ( .A1(n2591), .A2(REG0_REG_30__SCAN_IN), .ZN(n3196) );
  NAND3_X1 U4098 ( .A1(n3198), .A2(n3197), .A3(n3196), .ZN(n4102) );
  AOI22_X1 U4099 ( .A1(n4215), .A2(n4102), .B1(n4473), .B2(n3970), .ZN(n3199)
         );
  OAI21_X1 U4100 ( .B1(n3200), .B2(n4462), .A(n3199), .ZN(n3201) );
  NAND2_X1 U4101 ( .A1(n3203), .A2(n4669), .ZN(n3204) );
  AOI21_X1 U4102 ( .B1(n4486), .B2(n3204), .A(n4459), .ZN(n3205) );
  INV_X1 U4103 ( .A(n3205), .ZN(n3211) );
  NAND2_X1 U4104 ( .A1(n3206), .A2(n3970), .ZN(n3207) );
  INV_X1 U4105 ( .A(REG2_REG_29__SCAN_IN), .ZN(n3208) );
  OAI22_X1 U4106 ( .A1(n4490), .A2(n4461), .B1(n3208), .B2(n4351), .ZN(n3209)
         );
  INV_X1 U4107 ( .A(n3209), .ZN(n3210) );
  XNOR2_X1 U4108 ( .A(n3212), .B(n4022), .ZN(n4232) );
  NAND2_X1 U4109 ( .A1(n3213), .A2(n3214), .ZN(n3215) );
  XNOR2_X1 U4110 ( .A(n3215), .B(n4022), .ZN(n3216) );
  NAND2_X1 U4111 ( .A1(n3216), .A2(n4414), .ZN(n3221) );
  NOR2_X1 U4112 ( .A1(n4422), .A2(n3217), .ZN(n3218) );
  AOI21_X1 U4113 ( .B1(n3440), .B2(n4417), .A(n3218), .ZN(n3219) );
  AOI21_X1 U4114 ( .B1(n4232), .B2(n4545), .A(n4227), .ZN(n3233) );
  INV_X1 U4115 ( .A(n3222), .ZN(n4242) );
  NAND2_X1 U4116 ( .A1(n4242), .A2(n3223), .ZN(n3224) );
  NAND2_X1 U4117 ( .A1(n3206), .A2(n3224), .ZN(n4230) );
  INV_X1 U4118 ( .A(REG0_REG_28__SCAN_IN), .ZN(n4810) );
  NOR2_X1 U4119 ( .A1(n2374), .A2(n3225), .ZN(n3226) );
  OR2_X1 U4120 ( .A1(n4725), .A2(n4806), .ZN(n3229) );
  OAI21_X1 U4121 ( .B1(n4230), .B2(n4540), .A(n3229), .ZN(n3230) );
  INV_X1 U4122 ( .A(n3230), .ZN(n3231) );
  INV_X1 U4123 ( .A(DATAI_25_), .ZN(n3236) );
  NAND2_X1 U4124 ( .A1(n3234), .A2(STATE_REG_SCAN_IN), .ZN(n3235) );
  OAI21_X1 U4125 ( .B1(STATE_REG_SCAN_IN), .B2(n3236), .A(n3235), .ZN(U3327)
         );
  INV_X1 U4126 ( .A(DATAI_30_), .ZN(n3238) );
  NAND2_X1 U4127 ( .A1(n2565), .A2(STATE_REG_SCAN_IN), .ZN(n3237) );
  OAI21_X1 U4128 ( .B1(STATE_REG_SCAN_IN), .B2(n3238), .A(n3237), .ZN(U3322)
         );
  INV_X1 U4129 ( .A(DATAI_26_), .ZN(n3240) );
  NAND2_X1 U4130 ( .A1(n2856), .A2(STATE_REG_SCAN_IN), .ZN(n3239) );
  OAI21_X1 U4131 ( .B1(STATE_REG_SCAN_IN), .B2(n3240), .A(n3239), .ZN(U3326)
         );
  INV_X1 U4132 ( .A(DATAI_27_), .ZN(n4865) );
  NAND2_X1 U4133 ( .A1(n4611), .A2(STATE_REG_SCAN_IN), .ZN(n3241) );
  OAI21_X1 U4134 ( .B1(STATE_REG_SCAN_IN), .B2(n4865), .A(n3241), .ZN(U3325)
         );
  INV_X1 U4135 ( .A(DATAI_2_), .ZN(n3242) );
  MUX2_X1 U4136 ( .A(n2587), .B(n3242), .S(U3149), .Z(n3243) );
  INV_X1 U4137 ( .A(n3243), .ZN(U3350) );
  MUX2_X1 U4138 ( .A(n4131), .B(n2615), .S(U3149), .Z(n3244) );
  INV_X1 U4139 ( .A(n3244), .ZN(U3347) );
  INV_X1 U4140 ( .A(DATAI_22_), .ZN(n3246) );
  NAND2_X1 U4141 ( .A1(n2895), .A2(STATE_REG_SCAN_IN), .ZN(n3245) );
  OAI21_X1 U4142 ( .B1(STATE_REG_SCAN_IN), .B2(n3246), .A(n3245), .ZN(U3330)
         );
  MUX2_X1 U4143 ( .A(n3247), .B(n4185), .S(STATE_REG_SCAN_IN), .Z(n3248) );
  INV_X1 U4144 ( .A(n3248), .ZN(U3341) );
  INV_X1 U4145 ( .A(DATAI_24_), .ZN(n3251) );
  NAND2_X1 U4146 ( .A1(n3249), .A2(STATE_REG_SCAN_IN), .ZN(n3250) );
  OAI21_X1 U4147 ( .B1(STATE_REG_SCAN_IN), .B2(n3251), .A(n3250), .ZN(U3328)
         );
  INV_X1 U4148 ( .A(D_REG_0__SCAN_IN), .ZN(n4838) );
  INV_X1 U4149 ( .A(n3254), .ZN(n3255) );
  AOI22_X1 U4150 ( .A1(n4678), .A2(n4838), .B1(n4726), .B2(n3255), .ZN(U3458)
         );
  NOR2_X1 U4151 ( .A1(n4657), .A2(U4043), .ZN(U3148) );
  INV_X1 U4152 ( .A(DATAO_REG_12__SCAN_IN), .ZN(n4853) );
  NAND2_X1 U4153 ( .A1(U4043), .A2(n3256), .ZN(n3257) );
  OAI21_X1 U4154 ( .B1(U4043), .B2(n4853), .A(n3257), .ZN(U3562) );
  INV_X1 U4155 ( .A(DATAO_REG_2__SCAN_IN), .ZN(n4804) );
  NAND2_X1 U4156 ( .A1(U4043), .A2(n2909), .ZN(n3258) );
  OAI21_X1 U4157 ( .B1(U4043), .B2(n4804), .A(n3258), .ZN(U3552) );
  INV_X1 U4158 ( .A(DATAO_REG_6__SCAN_IN), .ZN(n4894) );
  NAND2_X1 U4159 ( .A1(U4043), .A2(n3589), .ZN(n3259) );
  OAI21_X1 U4160 ( .B1(U4043), .B2(n4894), .A(n3259), .ZN(U3556) );
  INV_X1 U4161 ( .A(DATAO_REG_10__SCAN_IN), .ZN(n4862) );
  NAND2_X1 U4162 ( .A1(U4043), .A2(n3490), .ZN(n3260) );
  OAI21_X1 U4163 ( .B1(U4043), .B2(n4862), .A(n3260), .ZN(U3560) );
  INV_X1 U4164 ( .A(DATAO_REG_8__SCAN_IN), .ZN(n4882) );
  NAND2_X1 U4165 ( .A1(U4043), .A2(n3703), .ZN(n3261) );
  OAI21_X1 U4166 ( .B1(U4043), .B2(n4882), .A(n3261), .ZN(U3558) );
  INV_X1 U4167 ( .A(DATAO_REG_15__SCAN_IN), .ZN(n4821) );
  NAND2_X1 U4168 ( .A1(n3782), .A2(U4043), .ZN(n3262) );
  OAI21_X1 U4169 ( .B1(U4043), .B2(n4821), .A(n3262), .ZN(U3565) );
  INV_X1 U4170 ( .A(DATAO_REG_18__SCAN_IN), .ZN(n4881) );
  NAND2_X1 U4171 ( .A1(n4419), .A2(U4043), .ZN(n3263) );
  OAI21_X1 U4172 ( .B1(U4043), .B2(n4881), .A(n3263), .ZN(U3568) );
  INV_X1 U4173 ( .A(DATAO_REG_17__SCAN_IN), .ZN(n4832) );
  NAND2_X1 U4174 ( .A1(n3910), .A2(U4043), .ZN(n3264) );
  OAI21_X1 U4175 ( .B1(U4043), .B2(n4832), .A(n3264), .ZN(U3567) );
  INV_X1 U4176 ( .A(DATAO_REG_4__SCAN_IN), .ZN(n4834) );
  NAND2_X1 U4177 ( .A1(U4043), .A2(n3535), .ZN(n3265) );
  OAI21_X1 U4178 ( .B1(U4043), .B2(n4834), .A(n3265), .ZN(U3554) );
  XNOR2_X1 U4179 ( .A(n3266), .B(REG1_REG_6__SCAN_IN), .ZN(n3274) );
  NAND2_X1 U4180 ( .A1(U3149), .A2(REG3_REG_6__SCAN_IN), .ZN(n3419) );
  NAND2_X1 U4181 ( .A1(n4657), .A2(ADDR_REG_6__SCAN_IN), .ZN(n3267) );
  OAI211_X1 U4182 ( .C1(n4668), .C2(n3268), .A(n3419), .B(n3267), .ZN(n3269)
         );
  INV_X1 U4183 ( .A(n3269), .ZN(n3273) );
  OAI211_X1 U4184 ( .C1(n3271), .C2(REG2_REG_6__SCAN_IN), .A(n3270), .B(n4664), 
        .ZN(n3272) );
  OAI211_X1 U4185 ( .C1(n3274), .C2(n4653), .A(n3273), .B(n3272), .ZN(U3246)
         );
  AOI21_X1 U4186 ( .B1(n4723), .B2(n4600), .A(n3275), .ZN(n3277) );
  XOR2_X1 U4187 ( .A(n3277), .B(n3276), .Z(n3284) );
  OAI211_X1 U4188 ( .C1(n3280), .C2(n3279), .A(n3278), .B(n4664), .ZN(n3282)
         );
  AND2_X1 U4189 ( .A1(U3149), .A2(REG3_REG_7__SCAN_IN), .ZN(n3480) );
  AOI21_X1 U4190 ( .B1(n4657), .B2(ADDR_REG_7__SCAN_IN), .A(n3480), .ZN(n3281)
         );
  OAI211_X1 U4191 ( .C1(n4668), .C2(n4600), .A(n3282), .B(n3281), .ZN(n3283)
         );
  AOI21_X1 U4192 ( .B1(n4648), .B2(n3284), .A(n3283), .ZN(n3285) );
  INV_X1 U4193 ( .A(n3285), .ZN(U3247) );
  INV_X1 U4194 ( .A(DATAO_REG_20__SCAN_IN), .ZN(n4902) );
  NAND2_X1 U4195 ( .A1(n3826), .A2(U4043), .ZN(n3286) );
  OAI21_X1 U4196 ( .B1(U4043), .B2(n4902), .A(n3286), .ZN(U3570) );
  INV_X1 U4197 ( .A(n4693), .ZN(n4702) );
  NAND2_X1 U4198 ( .A1(n3451), .A2(n4111), .ZN(n4026) );
  INV_X1 U4199 ( .A(n4007), .ZN(n3289) );
  NAND2_X1 U4200 ( .A1(n3296), .A2(n2885), .ZN(n3444) );
  INV_X1 U4201 ( .A(n3444), .ZN(n3288) );
  AND2_X1 U4202 ( .A1(n4366), .A2(n4468), .ZN(n3287) );
  OAI22_X1 U4203 ( .A1(n4007), .A2(n3287), .B1(n2897), .B2(n4464), .ZN(n3446)
         );
  AOI211_X1 U4204 ( .C1(n4702), .C2(n3289), .A(n3288), .B(n3446), .ZN(n4687)
         );
  NAND2_X1 U4205 ( .A1(n3232), .A2(REG1_REG_0__SCAN_IN), .ZN(n3290) );
  OAI21_X1 U4206 ( .B1(n4687), .B2(n3232), .A(n3290), .ZN(U3518) );
  INV_X1 U4207 ( .A(DATAO_REG_22__SCAN_IN), .ZN(n4835) );
  NAND2_X1 U4208 ( .A1(n3805), .A2(U4043), .ZN(n3291) );
  OAI21_X1 U4209 ( .B1(n4109), .B2(n4835), .A(n3291), .ZN(U3572) );
  INV_X1 U4210 ( .A(n3292), .ZN(n3295) );
  NAND3_X1 U4211 ( .A1(n3295), .A2(n3294), .A3(n3293), .ZN(n3792) );
  AOI22_X1 U4212 ( .A1(n3927), .A2(n3296), .B1(n3792), .B2(REG3_REG_0__SCAN_IN), .ZN(n3303) );
  INV_X1 U4213 ( .A(REG1_REG_0__SCAN_IN), .ZN(n4116) );
  NAND2_X1 U4214 ( .A1(n4685), .A2(n4116), .ZN(n4610) );
  AOI211_X1 U4215 ( .C1(n3299), .C2(n4610), .A(n3298), .B(n3297), .ZN(n3301)
         );
  NOR2_X1 U4216 ( .A1(n3301), .A2(n3300), .ZN(n3305) );
  AOI22_X1 U4217 ( .A1(n3305), .A2(n3888), .B1(n3938), .B2(n2601), .ZN(n3302)
         );
  NAND2_X1 U4218 ( .A1(n3303), .A2(n3302), .ZN(U3229) );
  XNOR2_X1 U4219 ( .A(n3304), .B(REG1_REG_4__SCAN_IN), .ZN(n3320) );
  NOR3_X1 U4220 ( .A1(n3305), .A2(n4611), .A3(n4606), .ZN(n3311) );
  OR2_X1 U4221 ( .A1(n3306), .A2(REG2_REG_0__SCAN_IN), .ZN(n3308) );
  AND2_X1 U4222 ( .A1(n3308), .A2(n3307), .ZN(n4607) );
  OAI22_X1 U4223 ( .A1(n4607), .A2(IR_REG_0__SCAN_IN), .B1(n3309), .B2(n4096), 
        .ZN(n3310) );
  NOR3_X1 U4224 ( .A1(n3311), .A2(n3439), .A3(n3310), .ZN(n3333) );
  NAND2_X1 U4225 ( .A1(REG3_REG_4__SCAN_IN), .A2(U3149), .ZN(n3376) );
  INV_X1 U4226 ( .A(n3376), .ZN(n3312) );
  AOI21_X1 U4227 ( .B1(n4657), .B2(ADDR_REG_4__SCAN_IN), .A(n3312), .ZN(n3313)
         );
  OAI21_X1 U4228 ( .B1(n4668), .B2(n3314), .A(n3313), .ZN(n3315) );
  NOR2_X1 U4229 ( .A1(n3333), .A2(n3315), .ZN(n3319) );
  OAI211_X1 U4230 ( .C1(REG2_REG_4__SCAN_IN), .C2(n3317), .A(n4664), .B(n3316), 
        .ZN(n3318) );
  OAI211_X1 U4231 ( .C1(n3320), .C2(n4653), .A(n3319), .B(n3318), .ZN(U3244)
         );
  AOI22_X1 U4232 ( .A1(n4657), .A2(ADDR_REG_2__SCAN_IN), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n3321) );
  OAI21_X1 U4233 ( .B1(n2587), .B2(n4668), .A(n3321), .ZN(n3332) );
  OAI211_X1 U4234 ( .C1(n3324), .C2(n3323), .A(n4664), .B(n3322), .ZN(n3330)
         );
  INV_X1 U4235 ( .A(REG1_REG_2__SCAN_IN), .ZN(n3357) );
  MUX2_X1 U4236 ( .A(n3357), .B(REG1_REG_2__SCAN_IN), .S(n2498), .Z(n3326) );
  NAND3_X1 U4237 ( .A1(n3326), .A2(n4118), .A3(n3325), .ZN(n3327) );
  NAND3_X1 U4238 ( .A1(n4648), .A2(n3328), .A3(n3327), .ZN(n3329) );
  NAND2_X1 U4239 ( .A1(n3330), .A2(n3329), .ZN(n3331) );
  OR3_X1 U4240 ( .A1(n3333), .A2(n3332), .A3(n3331), .ZN(U3242) );
  INV_X1 U4241 ( .A(DATAO_REG_23__SCAN_IN), .ZN(n4901) );
  NAND2_X1 U4242 ( .A1(n4326), .A2(U4043), .ZN(n3334) );
  OAI21_X1 U4243 ( .B1(U4043), .B2(n4901), .A(n3334), .ZN(U3573) );
  INV_X1 U4244 ( .A(n3335), .ZN(n3336) );
  AOI21_X1 U4245 ( .B1(n3338), .B2(n3337), .A(n3336), .ZN(n3342) );
  OAI22_X1 U4246 ( .A1(n3392), .A2(n3923), .B1(n3920), .B2(n2897), .ZN(n3340)
         );
  NOR2_X1 U4247 ( .A1(n3941), .A2(n3350), .ZN(n3339) );
  AOI211_X1 U4248 ( .C1(REG3_REG_2__SCAN_IN), .C2(n3792), .A(n3340), .B(n3339), 
        .ZN(n3341) );
  OAI21_X1 U4249 ( .B1(n3342), .B2(n3945), .A(n3341), .ZN(U3234) );
  NAND2_X1 U4250 ( .A1(n3343), .A2(n3344), .ZN(n3345) );
  NOR2_X1 U4251 ( .A1(n3345), .A2(n3348), .ZN(n3497) );
  AOI21_X1 U4252 ( .B1(n3348), .B2(n3345), .A(n3497), .ZN(n4670) );
  OAI21_X1 U4253 ( .B1(n3348), .B2(n3346), .A(n3347), .ZN(n3353) );
  AOI22_X1 U4254 ( .A1(n2601), .A2(n4417), .B1(n4418), .B2(n4110), .ZN(n3349)
         );
  OAI21_X1 U4255 ( .B1(n4422), .B2(n3350), .A(n3349), .ZN(n3352) );
  NOR2_X1 U4256 ( .A1(n4670), .A2(n4366), .ZN(n3351) );
  AOI211_X1 U4257 ( .C1(n4414), .C2(n3353), .A(n3352), .B(n3351), .ZN(n4677)
         );
  OAI21_X1 U4258 ( .B1(n4670), .B2(n4693), .A(n4677), .ZN(n3363) );
  INV_X1 U4259 ( .A(n3354), .ZN(n3450) );
  NAND2_X1 U4260 ( .A1(n3450), .A2(n3355), .ZN(n3356) );
  AND2_X1 U4261 ( .A1(n3356), .A2(n3506), .ZN(n4673) );
  INV_X1 U4262 ( .A(n4673), .ZN(n3361) );
  OAI22_X1 U4263 ( .A1(n4540), .A2(n3361), .B1(n4725), .B2(n3357), .ZN(n3358)
         );
  AOI21_X1 U4264 ( .B1(n3363), .B2(n4725), .A(n3358), .ZN(n3359) );
  INV_X1 U4265 ( .A(n3359), .ZN(U3520) );
  INV_X1 U4266 ( .A(REG0_REG_2__SCAN_IN), .ZN(n3360) );
  OAI22_X1 U4267 ( .A1(n4586), .A2(n3361), .B1(n4717), .B2(n3360), .ZN(n3362)
         );
  AOI21_X1 U4268 ( .B1(n3363), .B2(n4717), .A(n3362), .ZN(n3364) );
  INV_X1 U4269 ( .A(n3364), .ZN(U3471) );
  XOR2_X1 U4270 ( .A(n3366), .B(n3365), .Z(n3371) );
  OAI22_X1 U4271 ( .A1(n3789), .A2(n3920), .B1(n3923), .B2(n3367), .ZN(n3369)
         );
  MUX2_X1 U4272 ( .A(n3943), .B(U3149), .S(REG3_REG_3__SCAN_IN), .Z(n3368) );
  AOI211_X1 U4273 ( .C1(n3507), .C2(n3927), .A(n3369), .B(n3368), .ZN(n3370)
         );
  OAI21_X1 U4274 ( .B1(n3945), .B2(n3371), .A(n3370), .ZN(U3215) );
  AOI21_X1 U4275 ( .B1(n3372), .B2(n3373), .A(n3945), .ZN(n3375) );
  NAND2_X1 U4276 ( .A1(n3375), .A2(n3374), .ZN(n3380) );
  NAND2_X1 U4277 ( .A1(n3938), .A2(n4108), .ZN(n3377) );
  OAI211_X1 U4278 ( .C1(n3392), .C2(n3920), .A(n3377), .B(n3376), .ZN(n3378)
         );
  AOI21_X1 U4279 ( .B1(n3927), .B2(n3396), .A(n3378), .ZN(n3379) );
  OAI211_X1 U4280 ( .C1(n3922), .C2(n3401), .A(n3380), .B(n3379), .ZN(U3227)
         );
  AND2_X1 U4281 ( .A1(n4043), .A2(n4039), .ZN(n4000) );
  XNOR2_X1 U4282 ( .A(n3381), .B(n4000), .ZN(n3518) );
  XNOR2_X1 U4283 ( .A(n3382), .B(n4000), .ZN(n3383) );
  NAND2_X1 U4284 ( .A1(n3383), .A2(n4414), .ZN(n3385) );
  AOI22_X1 U4285 ( .A1(n4108), .A2(n4417), .B1(n4418), .B2(n4107), .ZN(n3384)
         );
  OAI211_X1 U4286 ( .C1(n2880), .C2(n4422), .A(n3385), .B(n3384), .ZN(n3512)
         );
  AOI21_X1 U4287 ( .B1(n3518), .B2(n4545), .A(n3512), .ZN(n3389) );
  INV_X1 U4288 ( .A(n3582), .ZN(n3386) );
  AOI21_X1 U4289 ( .B1(n3588), .B2(n2163), .A(n3386), .ZN(n3513) );
  AOI22_X1 U4290 ( .A1(n3513), .A2(n4481), .B1(REG1_REG_6__SCAN_IN), .B2(n3232), .ZN(n3387) );
  OAI21_X1 U4291 ( .B1(n3389), .B2(n3232), .A(n3387), .ZN(U3524) );
  AOI22_X1 U4292 ( .A1(n3513), .A2(n4554), .B1(REG0_REG_6__SCAN_IN), .B2(n4716), .ZN(n3388) );
  OAI21_X1 U4293 ( .B1(n3389), .B2(n4716), .A(n3388), .ZN(U3479) );
  XOR2_X1 U4294 ( .A(n4006), .B(n3391), .Z(n3398) );
  OAI22_X1 U4295 ( .A1(n4462), .A2(n3392), .B1(n2626), .B2(n4464), .ZN(n3395)
         );
  NAND2_X1 U4296 ( .A1(n3393), .A2(n3390), .ZN(n3540) );
  OAI21_X1 U4297 ( .B1(n3393), .B2(n3390), .A(n3540), .ZN(n3403) );
  NOR2_X1 U4298 ( .A1(n3403), .A2(n4366), .ZN(n3394) );
  AOI211_X1 U4299 ( .C1(n3396), .C2(n4473), .A(n3395), .B(n3394), .ZN(n3397)
         );
  OAI21_X1 U4300 ( .B1(n4468), .B2(n3398), .A(n3397), .ZN(n4700) );
  OAI211_X1 U4301 ( .C1(n3505), .C2(n3400), .A(n3399), .B(n4698), .ZN(n4699)
         );
  OAI22_X1 U4302 ( .A1(n4699), .A2(n4593), .B1(n4447), .B2(n3401), .ZN(n3402)
         );
  OAI21_X1 U4303 ( .B1(n4700), .B2(n3402), .A(n4351), .ZN(n3406) );
  INV_X1 U4304 ( .A(n3403), .ZN(n4703) );
  AOI22_X1 U4305 ( .A1(n4703), .A2(n4672), .B1(REG2_REG_4__SCAN_IN), .B2(n4459), .ZN(n3405) );
  NAND2_X1 U4306 ( .A1(n3406), .A2(n3405), .ZN(U3286) );
  OAI211_X1 U4307 ( .C1(n3409), .C2(n3408), .A(n3407), .B(n3888), .ZN(n3414)
         );
  AND2_X1 U4308 ( .A1(U3149), .A2(REG3_REG_5__SCAN_IN), .ZN(n4133) );
  AOI21_X1 U4309 ( .B1(n3937), .B2(n3535), .A(n4133), .ZN(n3411) );
  NAND2_X1 U4310 ( .A1(n3938), .A2(n3589), .ZN(n3410) );
  OAI211_X1 U4311 ( .C1(n3941), .C2(n3538), .A(n3411), .B(n3410), .ZN(n3412)
         );
  AOI21_X1 U4312 ( .B1(n3544), .B2(n3943), .A(n3412), .ZN(n3413) );
  NAND2_X1 U4313 ( .A1(n3414), .A2(n3413), .ZN(U3224) );
  XOR2_X1 U4314 ( .A(n3416), .B(n3415), .Z(n3417) );
  XNOR2_X1 U4315 ( .A(n3418), .B(n3417), .ZN(n3424) );
  OAI21_X1 U4316 ( .B1(n3923), .B2(n3554), .A(n3419), .ZN(n3420) );
  AOI21_X1 U4317 ( .B1(n3937), .B2(n4108), .A(n3420), .ZN(n3421) );
  OAI21_X1 U4318 ( .B1(n3941), .B2(n2880), .A(n3421), .ZN(n3422) );
  AOI21_X1 U4319 ( .B1(n3514), .B2(n3943), .A(n3422), .ZN(n3423) );
  OAI21_X1 U4320 ( .B1(n3424), .B2(n3945), .A(n3423), .ZN(U3236) );
  AND2_X1 U4321 ( .A1(n4045), .A2(n4049), .ZN(n4001) );
  XNOR2_X1 U4322 ( .A(n3425), .B(n4001), .ZN(n3573) );
  XNOR2_X1 U4323 ( .A(n3426), .B(n4001), .ZN(n3429) );
  AOI22_X1 U4324 ( .A1(n4418), .A2(n4106), .B1(n4417), .B2(n4107), .ZN(n3428)
         );
  NAND2_X1 U4325 ( .A1(n3434), .A2(n4473), .ZN(n3427) );
  OAI211_X1 U4326 ( .C1(n3429), .C2(n4468), .A(n3428), .B(n3427), .ZN(n3567)
         );
  AOI21_X1 U4327 ( .B1(n3573), .B2(n4545), .A(n3567), .ZN(n3437) );
  INV_X1 U4328 ( .A(n3430), .ZN(n3433) );
  INV_X1 U4329 ( .A(n3431), .ZN(n3432) );
  AOI21_X1 U4330 ( .B1(n3434), .B2(n3433), .A(n3432), .ZN(n3568) );
  AOI22_X1 U4331 ( .A1(n3568), .A2(n4554), .B1(REG0_REG_8__SCAN_IN), .B2(n4716), .ZN(n3435) );
  OAI21_X1 U4332 ( .B1(n3437), .B2(n4716), .A(n3435), .ZN(U3483) );
  AOI22_X1 U4333 ( .A1(n3568), .A2(n4481), .B1(REG1_REG_8__SCAN_IN), .B2(n3232), .ZN(n3436) );
  OAI21_X1 U4334 ( .B1(n3437), .B2(n3232), .A(n3436), .ZN(U3526) );
  NAND2_X1 U4335 ( .A1(n3439), .A2(DATAO_REG_29__SCAN_IN), .ZN(n3438) );
  OAI21_X1 U4336 ( .B1(n3971), .B2(n3439), .A(n3438), .ZN(U3579) );
  INV_X1 U4337 ( .A(DATAO_REG_27__SCAN_IN), .ZN(n4880) );
  NAND2_X1 U4338 ( .A1(n3440), .A2(U4043), .ZN(n3441) );
  OAI21_X1 U4339 ( .B1(n4109), .B2(n4880), .A(n3441), .ZN(U3577) );
  INV_X1 U4340 ( .A(n4672), .ZN(n3622) );
  INV_X1 U4341 ( .A(n3442), .ZN(n3443) );
  NOR2_X1 U4342 ( .A1(n3444), .A2(n3443), .ZN(n3445) );
  NOR2_X1 U4343 ( .A1(n3446), .A2(n3445), .ZN(n3447) );
  OAI22_X1 U4344 ( .A1(n4459), .A2(n3447), .B1(n2582), .B2(n4447), .ZN(n3448)
         );
  AOI21_X1 U4345 ( .B1(REG2_REG_0__SCAN_IN), .B2(n4459), .A(n3448), .ZN(n3449)
         );
  OAI21_X1 U4346 ( .B1(n3622), .B2(n4007), .A(n3449), .ZN(U3290) );
  OAI21_X1 U4347 ( .B1(n3451), .B2(n3798), .A(n3450), .ZN(n4689) );
  NAND2_X1 U4348 ( .A1(n3343), .A2(n3453), .ZN(n4690) );
  INV_X1 U4349 ( .A(n4690), .ZN(n3462) );
  AOI22_X1 U4350 ( .A1(n2909), .A2(n4418), .B1(n4417), .B2(n4111), .ZN(n3457)
         );
  NAND2_X1 U4351 ( .A1(n3455), .A2(n4473), .ZN(n3456) );
  OAI211_X1 U4352 ( .C1(n4690), .C2(n4366), .A(n3457), .B(n3456), .ZN(n3458)
         );
  AOI21_X1 U4353 ( .B1(n4414), .B2(n3459), .A(n3458), .ZN(n4688) );
  AOI22_X1 U4354 ( .A1(n4459), .A2(REG2_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(n4669), .ZN(n3460) );
  OAI21_X1 U4355 ( .B1(n4688), .B2(n4459), .A(n3460), .ZN(n3461) );
  AOI21_X1 U4356 ( .B1(n4672), .B2(n3462), .A(n3461), .ZN(n3463) );
  OAI21_X1 U4357 ( .B1(n4461), .B2(n4689), .A(n3463), .ZN(U3289) );
  INV_X1 U4358 ( .A(n4053), .ZN(n3464) );
  NAND2_X1 U4359 ( .A1(n3464), .A2(n4050), .ZN(n3999) );
  XOR2_X1 U4360 ( .A(n3999), .B(n3465), .Z(n3600) );
  XOR2_X1 U4361 ( .A(n3999), .B(n3466), .Z(n3470) );
  OAI22_X1 U4362 ( .A1(n4462), .A2(n3467), .B1(n3701), .B2(n4464), .ZN(n3468)
         );
  AOI21_X1 U4363 ( .B1(n4473), .B2(n3473), .A(n3468), .ZN(n3469) );
  OAI21_X1 U4364 ( .B1(n3470), .B2(n4468), .A(n3469), .ZN(n3601) );
  AOI21_X1 U4365 ( .B1(n3600), .B2(n4545), .A(n3601), .ZN(n3478) );
  INV_X1 U4366 ( .A(n3471), .ZN(n3472) );
  NAND2_X1 U4367 ( .A1(n3431), .A2(n3473), .ZN(n3474) );
  AND2_X1 U4368 ( .A1(n3472), .A2(n3474), .ZN(n3603) );
  NOR2_X1 U4369 ( .A1(n4725), .A2(n5004), .ZN(n3475) );
  AOI21_X1 U4370 ( .B1(n3603), .B2(n4481), .A(n3475), .ZN(n3476) );
  OAI21_X1 U4371 ( .B1(n3478), .B2(n3232), .A(n3476), .ZN(U3527) );
  AOI22_X1 U4372 ( .A1(n3603), .A2(n4554), .B1(REG0_REG_9__SCAN_IN), .B2(n4716), .ZN(n3477) );
  OAI21_X1 U4373 ( .B1(n3478), .B2(n4716), .A(n3477), .ZN(U3485) );
  XNOR2_X1 U4374 ( .A(n3479), .B(n3549), .ZN(n3485) );
  AOI21_X1 U4375 ( .B1(n3937), .B2(n3589), .A(n3480), .ZN(n3482) );
  NAND2_X1 U4376 ( .A1(n3938), .A2(n3703), .ZN(n3481) );
  OAI211_X1 U4377 ( .C1(n3941), .C2(n3580), .A(n3482), .B(n3481), .ZN(n3483)
         );
  AOI21_X1 U4378 ( .B1(n3585), .B2(n3943), .A(n3483), .ZN(n3484) );
  OAI21_X1 U4379 ( .B1(n3485), .B2(n3945), .A(n3484), .ZN(U3210) );
  XOR2_X1 U4380 ( .A(n3487), .B(n3486), .Z(n3488) );
  XNOR2_X1 U4381 ( .A(n3489), .B(n3488), .ZN(n3495) );
  NAND2_X1 U4382 ( .A1(n3937), .A2(n3490), .ZN(n3491) );
  NAND2_X1 U4383 ( .A1(U3149), .A2(REG3_REG_11__SCAN_IN), .ZN(n4180) );
  OAI211_X1 U4384 ( .C1(n3714), .C2(n3923), .A(n3491), .B(n4180), .ZN(n3493)
         );
  NOR2_X1 U4385 ( .A1(n3922), .A2(n3617), .ZN(n3492) );
  AOI211_X1 U4386 ( .C1(n3616), .C2(n3927), .A(n3493), .B(n3492), .ZN(n3494)
         );
  OAI21_X1 U4387 ( .B1(n3495), .B2(n3945), .A(n3494), .ZN(U3233) );
  NOR2_X1 U4388 ( .A1(n3497), .A2(n3496), .ZN(n3498) );
  XOR2_X1 U4389 ( .A(n4004), .B(n3498), .Z(n4694) );
  XNOR2_X1 U4390 ( .A(n3499), .B(n4004), .ZN(n3503) );
  AOI22_X1 U4391 ( .A1(n2909), .A2(n4417), .B1(n4418), .B2(n3535), .ZN(n3500)
         );
  OAI21_X1 U4392 ( .B1(n4422), .B2(n3501), .A(n3500), .ZN(n3502) );
  AOI21_X1 U4393 ( .B1(n3503), .B2(n4414), .A(n3502), .ZN(n3504) );
  OAI21_X1 U4394 ( .B1(n4694), .B2(n4366), .A(n3504), .ZN(n4695) );
  NAND2_X1 U4395 ( .A1(n4695), .A2(n4351), .ZN(n3511) );
  AOI21_X1 U4396 ( .B1(n3507), .B2(n3506), .A(n3505), .ZN(n4697) );
  INV_X1 U4397 ( .A(REG2_REG_3__SCAN_IN), .ZN(n3508) );
  OAI22_X1 U4398 ( .A1(n4351), .A2(n3508), .B1(REG3_REG_3__SCAN_IN), .B2(n4447), .ZN(n3509) );
  AOI21_X1 U4399 ( .B1(n4674), .B2(n4697), .A(n3509), .ZN(n3510) );
  OAI211_X1 U4400 ( .C1(n4694), .C2(n3622), .A(n3511), .B(n3510), .ZN(U3287)
         );
  INV_X1 U4401 ( .A(n3512), .ZN(n3520) );
  INV_X1 U4402 ( .A(n3513), .ZN(n3516) );
  AOI22_X1 U4403 ( .A1(n4459), .A2(REG2_REG_6__SCAN_IN), .B1(n3514), .B2(n4669), .ZN(n3515) );
  OAI21_X1 U4404 ( .B1(n3516), .B2(n4461), .A(n3515), .ZN(n3517) );
  AOI21_X1 U4405 ( .B1(n3518), .B2(n4477), .A(n3517), .ZN(n3519) );
  OAI21_X1 U4406 ( .B1(n3520), .B2(n4459), .A(n3519), .ZN(U3284) );
  NAND2_X1 U4407 ( .A1(n4052), .A2(n4055), .ZN(n3994) );
  XNOR2_X1 U4408 ( .A(n3521), .B(n3994), .ZN(n3524) );
  AOI22_X1 U4409 ( .A1(n4418), .A2(n4105), .B1(n4417), .B2(n4106), .ZN(n3523)
         );
  NAND2_X1 U4410 ( .A1(n3735), .A2(n4473), .ZN(n3522) );
  OAI211_X1 U4411 ( .C1(n3524), .C2(n4468), .A(n3523), .B(n3522), .ZN(n3561)
         );
  INV_X1 U4412 ( .A(n3561), .ZN(n3531) );
  AOI21_X1 U4413 ( .B1(n3735), .B2(n3472), .A(n3613), .ZN(n3564) );
  INV_X1 U4414 ( .A(REG2_REG_10__SCAN_IN), .ZN(n3526) );
  INV_X1 U4415 ( .A(n3525), .ZN(n3738) );
  OAI22_X1 U4416 ( .A1(n4351), .A2(n3526), .B1(n3738), .B2(n4447), .ZN(n3527)
         );
  AOI21_X1 U4417 ( .B1(n3564), .B2(n4674), .A(n3527), .ZN(n3530) );
  XNOR2_X1 U4418 ( .A(n3528), .B(n3994), .ZN(n3562) );
  NAND2_X1 U4419 ( .A1(n3562), .A2(n4477), .ZN(n3529) );
  OAI211_X1 U4420 ( .C1(n3531), .C2(n4459), .A(n3530), .B(n3529), .ZN(U3280)
         );
  NAND2_X1 U4421 ( .A1(n2247), .A2(n4041), .ZN(n3996) );
  XNOR2_X1 U4422 ( .A(n3533), .B(n3996), .ZN(n3534) );
  NAND2_X1 U4423 ( .A1(n3534), .A2(n4414), .ZN(n3537) );
  AOI22_X1 U4424 ( .A1(n4418), .A2(n3589), .B1(n4417), .B2(n3535), .ZN(n3536)
         );
  OAI211_X1 U4425 ( .C1(n3538), .C2(n4422), .A(n3537), .B(n3536), .ZN(n4709)
         );
  INV_X1 U4426 ( .A(n4459), .ZN(n4351) );
  NAND2_X1 U4427 ( .A1(n3540), .A2(n3539), .ZN(n3541) );
  XNOR2_X1 U4428 ( .A(n3541), .B(n3996), .ZN(n4707) );
  NOR2_X1 U4429 ( .A1(n4707), .A2(n4452), .ZN(n3547) );
  NAND2_X1 U4430 ( .A1(n3399), .A2(n3542), .ZN(n3543) );
  NAND2_X1 U4431 ( .A1(n2163), .A2(n3543), .ZN(n4705) );
  AOI22_X1 U4432 ( .A1(n4459), .A2(REG2_REG_5__SCAN_IN), .B1(n3544), .B2(n4669), .ZN(n3545) );
  OAI21_X1 U4433 ( .B1(n4461), .B2(n4705), .A(n3545), .ZN(n3546) );
  AOI211_X1 U4434 ( .C1(n4709), .C2(n4351), .A(n3547), .B(n3546), .ZN(n3548)
         );
  INV_X1 U4435 ( .A(n3548), .ZN(U3285) );
  NAND2_X1 U4436 ( .A1(n3479), .A2(n3549), .ZN(n3551) );
  NAND2_X1 U4437 ( .A1(n3551), .A2(n3550), .ZN(n3697) );
  INV_X1 U4438 ( .A(n3698), .ZN(n3552) );
  NOR2_X1 U4439 ( .A1(n3552), .A2(n3696), .ZN(n3553) );
  XNOR2_X1 U4440 ( .A(n3697), .B(n3553), .ZN(n3560) );
  NAND2_X1 U4441 ( .A1(U3149), .A2(REG3_REG_8__SCAN_IN), .ZN(n4145) );
  OAI21_X1 U4442 ( .B1(n3920), .B2(n3554), .A(n4145), .ZN(n3555) );
  AOI21_X1 U4443 ( .B1(n3938), .B2(n4106), .A(n3555), .ZN(n3556) );
  OAI21_X1 U4444 ( .B1(n3941), .B2(n3557), .A(n3556), .ZN(n3558) );
  AOI21_X1 U4445 ( .B1(n3569), .B2(n3943), .A(n3558), .ZN(n3559) );
  OAI21_X1 U4446 ( .B1(n3560), .B2(n3945), .A(n3559), .ZN(U3218) );
  AOI21_X1 U4447 ( .B1(n4545), .B2(n3562), .A(n3561), .ZN(n3566) );
  AOI22_X1 U4448 ( .A1(n3564), .A2(n4554), .B1(REG0_REG_10__SCAN_IN), .B2(
        n4716), .ZN(n3563) );
  OAI21_X1 U4449 ( .B1(n3566), .B2(n4716), .A(n3563), .ZN(U3487) );
  AOI22_X1 U4450 ( .A1(n3564), .A2(n4481), .B1(REG1_REG_10__SCAN_IN), .B2(
        n3232), .ZN(n3565) );
  OAI21_X1 U4451 ( .B1(n3566), .B2(n3232), .A(n3565), .ZN(U3528) );
  INV_X1 U4452 ( .A(n3567), .ZN(n3575) );
  INV_X1 U4453 ( .A(n3568), .ZN(n3571) );
  AOI22_X1 U4454 ( .A1(n4459), .A2(REG2_REG_8__SCAN_IN), .B1(n3569), .B2(n4669), .ZN(n3570) );
  OAI21_X1 U4455 ( .B1(n3571), .B2(n4461), .A(n3570), .ZN(n3572) );
  AOI21_X1 U4456 ( .B1(n3573), .B2(n4477), .A(n3572), .ZN(n3574) );
  OAI21_X1 U4457 ( .B1(n3575), .B2(n4459), .A(n3574), .ZN(U3282) );
  INV_X1 U4458 ( .A(n3592), .ZN(n4005) );
  XNOR2_X1 U4459 ( .A(n3576), .B(n4005), .ZN(n3577) );
  NAND2_X1 U4460 ( .A1(n3577), .A2(n4414), .ZN(n3579) );
  AOI22_X1 U4461 ( .A1(n3703), .A2(n4418), .B1(n4417), .B2(n3589), .ZN(n3578)
         );
  OAI211_X1 U4462 ( .C1(n3580), .C2(n4422), .A(n3579), .B(n3578), .ZN(n4714)
         );
  INV_X1 U4463 ( .A(n4714), .ZN(n3599) );
  INV_X1 U4464 ( .A(n4409), .ZN(n3597) );
  NAND2_X1 U4465 ( .A1(n3582), .A2(n3581), .ZN(n3583) );
  NAND2_X1 U4466 ( .A1(n3583), .A2(n4698), .ZN(n3584) );
  NOR2_X1 U4467 ( .A1(n3430), .A2(n3584), .ZN(n4713) );
  INV_X1 U4468 ( .A(n3585), .ZN(n3586) );
  OAI22_X1 U4469 ( .A1(n4351), .A2(n3587), .B1(n3586), .B2(n4447), .ZN(n3596)
         );
  INV_X1 U4470 ( .A(n3381), .ZN(n3591) );
  AOI21_X1 U4471 ( .B1(n3381), .B2(n3589), .A(n3588), .ZN(n3590) );
  AOI21_X1 U4472 ( .B1(n3591), .B2(n2648), .A(n3590), .ZN(n3593) );
  NOR2_X1 U4473 ( .A1(n3593), .A2(n3592), .ZN(n4712) );
  INV_X1 U4474 ( .A(n3593), .ZN(n3594) );
  NOR2_X1 U4475 ( .A1(n3594), .A2(n4005), .ZN(n4711) );
  NOR3_X1 U4476 ( .A1(n4712), .A2(n4711), .A3(n4452), .ZN(n3595) );
  AOI211_X1 U4477 ( .C1(n3597), .C2(n4713), .A(n3596), .B(n3595), .ZN(n3598)
         );
  OAI21_X1 U4478 ( .B1(n4459), .B2(n3599), .A(n3598), .ZN(U3283) );
  INV_X1 U4479 ( .A(n3600), .ZN(n3606) );
  INV_X1 U4480 ( .A(n3601), .ZN(n3602) );
  MUX2_X1 U4481 ( .A(n4931), .B(n3602), .S(n4351), .Z(n3605) );
  AOI22_X1 U4482 ( .A1(n3603), .A2(n4674), .B1(n3707), .B2(n4669), .ZN(n3604)
         );
  OAI211_X1 U4483 ( .C1(n4452), .C2(n3606), .A(n3605), .B(n3604), .ZN(U3281)
         );
  OR2_X1 U4484 ( .A1(n3608), .A2(n3988), .ZN(n3656) );
  INV_X1 U4485 ( .A(n3656), .ZN(n3607) );
  AOI21_X1 U4486 ( .B1(n3988), .B2(n3608), .A(n3607), .ZN(n3665) );
  XOR2_X1 U4487 ( .A(n3988), .B(n3650), .Z(n3612) );
  OAI22_X1 U4488 ( .A1(n3701), .A2(n4462), .B1(n3714), .B2(n4464), .ZN(n3610)
         );
  NOR2_X1 U4489 ( .A1(n3665), .A2(n4366), .ZN(n3609) );
  AOI211_X1 U4490 ( .C1(n3616), .C2(n4473), .A(n3610), .B(n3609), .ZN(n3611)
         );
  OAI21_X1 U4491 ( .B1(n4468), .B2(n3612), .A(n3611), .ZN(n3666) );
  NAND2_X1 U4492 ( .A1(n3666), .A2(n4351), .ZN(n3621) );
  INV_X1 U4493 ( .A(n3613), .ZN(n3615) );
  AOI21_X1 U4494 ( .B1(n3616), .B2(n3615), .A(n3614), .ZN(n3669) );
  OAI22_X1 U4495 ( .A1(n4351), .A2(n3618), .B1(n3617), .B2(n4447), .ZN(n3619)
         );
  AOI21_X1 U4496 ( .B1(n3669), .B2(n4674), .A(n3619), .ZN(n3620) );
  OAI211_X1 U4497 ( .C1(n3665), .C2(n3622), .A(n3621), .B(n3620), .ZN(U3279)
         );
  INV_X1 U4498 ( .A(n3624), .ZN(n3626) );
  NOR2_X1 U4499 ( .A1(n3626), .A2(n3625), .ZN(n3627) );
  XNOR2_X1 U4500 ( .A(n3623), .B(n3627), .ZN(n3632) );
  NAND2_X1 U4501 ( .A1(n3937), .A2(n4105), .ZN(n3628) );
  NAND2_X1 U4502 ( .A1(U3149), .A2(REG3_REG_12__SCAN_IN), .ZN(n4192) );
  OAI211_X1 U4503 ( .C1(n3780), .C2(n3923), .A(n3628), .B(n4192), .ZN(n3630)
         );
  NOR2_X1 U4504 ( .A1(n3922), .A2(n3657), .ZN(n3629) );
  AOI211_X1 U4505 ( .C1(n3652), .C2(n3927), .A(n3630), .B(n3629), .ZN(n3631)
         );
  OAI21_X1 U4506 ( .B1(n3632), .B2(n3945), .A(n3631), .ZN(U3221) );
  XNOR2_X1 U4507 ( .A(n3948), .B(n3989), .ZN(n3636) );
  NAND2_X1 U4508 ( .A1(n3782), .A2(n4418), .ZN(n3634) );
  NAND2_X1 U4509 ( .A1(n3643), .A2(n4473), .ZN(n3633) );
  OAI211_X1 U4510 ( .C1(n3780), .C2(n4462), .A(n3634), .B(n3633), .ZN(n3635)
         );
  AOI21_X1 U4511 ( .B1(n3636), .B2(n4414), .A(n3635), .ZN(n3748) );
  NAND2_X1 U4512 ( .A1(n3656), .A2(n3637), .ZN(n3639) );
  NAND2_X1 U4513 ( .A1(n3639), .A2(n3638), .ZN(n3640) );
  AND2_X1 U4514 ( .A1(n3640), .A2(n3989), .ZN(n3642) );
  OR2_X1 U4515 ( .A1(n3642), .A2(n3641), .ZN(n3747) );
  AOI21_X1 U4516 ( .B1(n3643), .B2(n3690), .A(n4457), .ZN(n3761) );
  INV_X1 U4517 ( .A(n3761), .ZN(n3752) );
  AOI22_X1 U4518 ( .A1(n4459), .A2(REG2_REG_14__SCAN_IN), .B1(n3786), .B2(
        n4669), .ZN(n3644) );
  OAI21_X1 U4519 ( .B1(n3752), .B2(n4461), .A(n3644), .ZN(n3645) );
  AOI21_X1 U4520 ( .B1(n3747), .B2(n4477), .A(n3645), .ZN(n3646) );
  OAI21_X1 U4521 ( .B1(n4459), .B2(n3748), .A(n3646), .ZN(U3276) );
  NAND2_X1 U4522 ( .A1(n3672), .A2(n3674), .ZN(n4011) );
  INV_X1 U4523 ( .A(n3647), .ZN(n3648) );
  AOI21_X1 U4524 ( .B1(n3650), .B2(n3649), .A(n3648), .ZN(n3675) );
  XOR2_X1 U4525 ( .A(n4011), .B(n3675), .Z(n3654) );
  OAI22_X1 U4526 ( .A1(n3780), .A2(n4464), .B1(n3733), .B2(n4462), .ZN(n3651)
         );
  AOI21_X1 U4527 ( .B1(n4473), .B2(n3652), .A(n3651), .ZN(n3653) );
  OAI21_X1 U4528 ( .B1(n3654), .B2(n4468), .A(n3653), .ZN(n3739) );
  INV_X1 U4529 ( .A(n3739), .ZN(n3664) );
  NAND2_X1 U4530 ( .A1(n3656), .A2(n3655), .ZN(n3680) );
  XNOR2_X1 U4531 ( .A(n3680), .B(n4011), .ZN(n3740) );
  OAI22_X1 U4532 ( .A1(n4351), .A2(n3658), .B1(n3657), .B2(n4447), .ZN(n3662)
         );
  OAI21_X1 U4533 ( .B1(n3614), .B2(n3660), .A(n3659), .ZN(n3746) );
  NOR2_X1 U4534 ( .A1(n3746), .A2(n4461), .ZN(n3661) );
  AOI211_X1 U4535 ( .C1(n3740), .C2(n4477), .A(n3662), .B(n3661), .ZN(n3663)
         );
  OAI21_X1 U4536 ( .B1(n3664), .B2(n4459), .A(n3663), .ZN(U3278) );
  INV_X1 U4537 ( .A(n3665), .ZN(n3667) );
  AOI21_X1 U4538 ( .B1(n4702), .B2(n3667), .A(n3666), .ZN(n3671) );
  AOI22_X1 U4539 ( .A1(n3669), .A2(n4481), .B1(REG1_REG_11__SCAN_IN), .B2(
        n3232), .ZN(n3668) );
  OAI21_X1 U4540 ( .B1(n3671), .B2(n3232), .A(n3668), .ZN(U3529) );
  AOI22_X1 U4541 ( .A1(n3669), .A2(n4554), .B1(REG0_REG_11__SCAN_IN), .B2(
        n4716), .ZN(n3670) );
  OAI21_X1 U4542 ( .B1(n3671), .B2(n4716), .A(n3670), .ZN(U3489) );
  INV_X1 U4543 ( .A(n3672), .ZN(n3673) );
  AOI21_X1 U4544 ( .B1(n3675), .B2(n3674), .A(n3673), .ZN(n3678) );
  NAND2_X1 U4545 ( .A1(n3677), .A2(n3676), .ZN(n4012) );
  XNOR2_X1 U4546 ( .A(n3678), .B(n4012), .ZN(n3688) );
  OAI22_X1 U4547 ( .A1(n4463), .A2(n4464), .B1(n3714), .B2(n4462), .ZN(n3685)
         );
  NAND2_X1 U4548 ( .A1(n3680), .A2(n3679), .ZN(n3682) );
  NAND2_X1 U4549 ( .A1(n3682), .A2(n3681), .ZN(n3683) );
  XOR2_X1 U4550 ( .A(n4012), .B(n3683), .Z(n3689) );
  NOR2_X1 U4551 ( .A1(n3689), .A2(n4366), .ZN(n3684) );
  AOI211_X1 U4552 ( .C1(n3686), .C2(n4473), .A(n3685), .B(n3684), .ZN(n3687)
         );
  OAI21_X1 U4553 ( .B1(n4468), .B2(n3688), .A(n3687), .ZN(n3753) );
  INV_X1 U4554 ( .A(n3753), .ZN(n3695) );
  INV_X1 U4555 ( .A(n3689), .ZN(n3754) );
  INV_X1 U4556 ( .A(n3659), .ZN(n3691) );
  OAI21_X1 U4557 ( .B1(n3691), .B2(n3717), .A(n3690), .ZN(n3758) );
  AOI22_X1 U4558 ( .A1(n4459), .A2(REG2_REG_13__SCAN_IN), .B1(n3719), .B2(
        n4669), .ZN(n3692) );
  OAI21_X1 U4559 ( .B1(n3758), .B2(n4461), .A(n3692), .ZN(n3693) );
  AOI21_X1 U4560 ( .B1(n3754), .B2(n4672), .A(n3693), .ZN(n3694) );
  OAI21_X1 U4561 ( .B1(n3695), .B2(n4459), .A(n3694), .ZN(U3277) );
  NAND2_X1 U4562 ( .A1(n3727), .A2(n3698), .ZN(n3699) );
  XOR2_X1 U4563 ( .A(n3700), .B(n3699), .Z(n3709) );
  NAND2_X1 U4564 ( .A1(U3149), .A2(REG3_REG_9__SCAN_IN), .ZN(n4157) );
  OAI21_X1 U4565 ( .B1(n3923), .B2(n3701), .A(n4157), .ZN(n3702) );
  AOI21_X1 U4566 ( .B1(n3937), .B2(n3703), .A(n3702), .ZN(n3704) );
  OAI21_X1 U4567 ( .B1(n3941), .B2(n3705), .A(n3704), .ZN(n3706) );
  AOI21_X1 U4568 ( .B1(n3707), .B2(n3943), .A(n3706), .ZN(n3708) );
  OAI21_X1 U4569 ( .B1(n3709), .B2(n3945), .A(n3708), .ZN(U3228) );
  XOR2_X1 U4570 ( .A(n3712), .B(n3711), .Z(n3713) );
  XNOR2_X1 U4571 ( .A(n3710), .B(n3713), .ZN(n3721) );
  NAND2_X1 U4572 ( .A1(U3149), .A2(REG3_REG_13__SCAN_IN), .ZN(n4204) );
  OAI21_X1 U4573 ( .B1(n3920), .B2(n3714), .A(n4204), .ZN(n3715) );
  AOI21_X1 U4574 ( .B1(n3938), .B2(n4103), .A(n3715), .ZN(n3716) );
  OAI21_X1 U4575 ( .B1(n3941), .B2(n3717), .A(n3716), .ZN(n3718) );
  AOI21_X1 U4576 ( .B1(n3719), .B2(n3943), .A(n3718), .ZN(n3720) );
  OAI21_X1 U4577 ( .B1(n3721), .B2(n3945), .A(n3720), .ZN(U3231) );
  NAND2_X1 U4578 ( .A1(n3727), .A2(n3722), .ZN(n3724) );
  AND2_X1 U4579 ( .A1(n3724), .A2(n3723), .ZN(n3725) );
  AOI21_X1 U4580 ( .B1(n3725), .B2(n2959), .A(n3945), .ZN(n3731) );
  NAND2_X1 U4581 ( .A1(n3727), .A2(n3726), .ZN(n3729) );
  AND2_X1 U4582 ( .A1(n3729), .A2(n3728), .ZN(n3730) );
  NAND2_X1 U4583 ( .A1(n3731), .A2(n3730), .ZN(n3737) );
  NAND2_X1 U4584 ( .A1(n3937), .A2(n4106), .ZN(n3732) );
  NAND2_X1 U4585 ( .A1(U3149), .A2(REG3_REG_10__SCAN_IN), .ZN(n4168) );
  OAI211_X1 U4586 ( .C1(n3733), .C2(n3923), .A(n3732), .B(n4168), .ZN(n3734)
         );
  AOI21_X1 U4587 ( .B1(n3927), .B2(n3735), .A(n3734), .ZN(n3736) );
  OAI211_X1 U4588 ( .C1(n3922), .C2(n3738), .A(n3737), .B(n3736), .ZN(U3214)
         );
  INV_X1 U4589 ( .A(REG0_REG_12__SCAN_IN), .ZN(n3741) );
  AOI21_X1 U4590 ( .B1(n4545), .B2(n3740), .A(n3739), .ZN(n3743) );
  MUX2_X1 U4591 ( .A(n3741), .B(n3743), .S(n4717), .Z(n3742) );
  OAI21_X1 U4592 ( .B1(n3746), .B2(n4586), .A(n3742), .ZN(U3491) );
  INV_X1 U4593 ( .A(REG1_REG_12__SCAN_IN), .ZN(n3744) );
  MUX2_X1 U4594 ( .A(n3744), .B(n3743), .S(n4725), .Z(n3745) );
  OAI21_X1 U4595 ( .B1(n4540), .B2(n3746), .A(n3745), .ZN(U3530) );
  NAND2_X1 U4596 ( .A1(n3747), .A2(n4545), .ZN(n3749) );
  NAND2_X1 U4597 ( .A1(n3749), .A2(n3748), .ZN(n3759) );
  INV_X1 U4598 ( .A(n3759), .ZN(n3750) );
  MUX2_X1 U4599 ( .A(n3750), .B(n4770), .S(n3232), .Z(n3751) );
  OAI21_X1 U4600 ( .B1(n4540), .B2(n3752), .A(n3751), .ZN(U3532) );
  AOI21_X1 U4601 ( .B1(n4702), .B2(n3754), .A(n3753), .ZN(n3756) );
  MUX2_X1 U4602 ( .A(n5005), .B(n3756), .S(n4725), .Z(n3755) );
  OAI21_X1 U4603 ( .B1(n4540), .B2(n3758), .A(n3755), .ZN(U3531) );
  INV_X1 U4604 ( .A(REG0_REG_13__SCAN_IN), .ZN(n4956) );
  MUX2_X1 U4605 ( .A(n4956), .B(n3756), .S(n4717), .Z(n3757) );
  OAI21_X1 U4606 ( .B1(n3758), .B2(n4586), .A(n3757), .ZN(U3493) );
  MUX2_X1 U4607 ( .A(REG0_REG_14__SCAN_IN), .B(n3759), .S(n4717), .Z(n3760) );
  AOI21_X1 U4608 ( .B1(n3761), .B2(n4554), .A(n3760), .ZN(n3762) );
  INV_X1 U4609 ( .A(n3762), .ZN(U3495) );
  AOI211_X1 U4610 ( .C1(n4932), .C2(n3764), .A(n4615), .B(n3763), .ZN(n3771)
         );
  AOI211_X1 U4611 ( .C1(n3766), .C2(n4770), .A(n4653), .B(n3765), .ZN(n3770)
         );
  NAND2_X1 U4612 ( .A1(U3149), .A2(REG3_REG_14__SCAN_IN), .ZN(n3779) );
  NAND2_X1 U4613 ( .A1(n4657), .A2(ADDR_REG_14__SCAN_IN), .ZN(n3767) );
  OAI211_X1 U4614 ( .C1(n4668), .C2(n3768), .A(n3779), .B(n3767), .ZN(n3769)
         );
  OR3_X1 U4615 ( .A1(n3771), .A2(n3770), .A3(n3769), .ZN(U3254) );
  INV_X1 U4616 ( .A(n3772), .ZN(n3775) );
  INV_X1 U4617 ( .A(IR_REG_30__SCAN_IN), .ZN(n4868) );
  NAND3_X1 U4618 ( .A1(IR_REG_31__SCAN_IN), .A2(STATE_REG_SCAN_IN), .A3(n4868), 
        .ZN(n3774) );
  INV_X1 U4619 ( .A(DATAI_31_), .ZN(n3773) );
  OAI22_X1 U4620 ( .A1(n3775), .A2(n3774), .B1(STATE_REG_SCAN_IN), .B2(n3773), 
        .ZN(U3321) );
  NOR2_X1 U4621 ( .A1(n3850), .A2(n3777), .ZN(n3778) );
  XNOR2_X1 U4622 ( .A(n3776), .B(n3778), .ZN(n3788) );
  OAI21_X1 U4623 ( .B1(n3920), .B2(n3780), .A(n3779), .ZN(n3781) );
  AOI21_X1 U4624 ( .B1(n3938), .B2(n3782), .A(n3781), .ZN(n3783) );
  OAI21_X1 U4625 ( .B1(n3941), .B2(n3784), .A(n3783), .ZN(n3785) );
  AOI21_X1 U4626 ( .B1(n3786), .B2(n3943), .A(n3785), .ZN(n3787) );
  OAI21_X1 U4627 ( .B1(n3788), .B2(n3945), .A(n3787), .ZN(U3212) );
  OAI22_X1 U4628 ( .A1(n3790), .A2(n3920), .B1(n3923), .B2(n3789), .ZN(n3791)
         );
  AOI21_X1 U4629 ( .B1(n3792), .B2(REG3_REG_1__SCAN_IN), .A(n3791), .ZN(n3797)
         );
  OAI211_X1 U4630 ( .C1(n3795), .C2(n3794), .A(n3888), .B(n3793), .ZN(n3796)
         );
  OAI211_X1 U4631 ( .C1(n3941), .C2(n3798), .A(n3797), .B(n3796), .ZN(U3219)
         );
  AND2_X1 U4632 ( .A1(n3799), .A2(n3800), .ZN(n3802) );
  OAI211_X1 U4633 ( .C1(n3802), .C2(n3801), .A(n3888), .B(n3837), .ZN(n3807)
         );
  NOR2_X1 U4634 ( .A1(n3941), .A2(n4313), .ZN(n3804) );
  OAI22_X1 U4635 ( .A1(n4265), .A2(n3923), .B1(STATE_REG_SCAN_IN), .B2(n4792), 
        .ZN(n3803) );
  AOI211_X1 U4636 ( .C1(n3937), .C2(n3805), .A(n3804), .B(n3803), .ZN(n3806)
         );
  OAI211_X1 U4637 ( .C1(n3922), .C2(n4309), .A(n3807), .B(n3806), .ZN(U3213)
         );
  INV_X1 U4638 ( .A(n3808), .ZN(n3809) );
  NAND2_X1 U4639 ( .A1(n3810), .A2(n3809), .ZN(n3813) );
  INV_X1 U4640 ( .A(n3811), .ZN(n3812) );
  AOI21_X1 U4641 ( .B1(n3814), .B2(n3813), .A(n3812), .ZN(n3820) );
  NAND2_X1 U4642 ( .A1(n3937), .A2(n4419), .ZN(n3816) );
  OAI211_X1 U4643 ( .C1(n4385), .C2(n3923), .A(n3816), .B(n3815), .ZN(n3818)
         );
  NOR2_X1 U4644 ( .A1(n3922), .A2(n4391), .ZN(n3817) );
  AOI211_X1 U4645 ( .C1(n4382), .C2(n3927), .A(n3818), .B(n3817), .ZN(n3819)
         );
  OAI21_X1 U4646 ( .B1(n3820), .B2(n3945), .A(n3819), .ZN(U3216) );
  INV_X1 U4647 ( .A(n4348), .ZN(n3832) );
  NAND2_X1 U4648 ( .A1(n2162), .A2(n3822), .ZN(n3825) );
  NAND2_X1 U4649 ( .A1(n3811), .A2(n3823), .ZN(n3885) );
  INV_X1 U4650 ( .A(n3886), .ZN(n3883) );
  OAI211_X1 U4651 ( .C1(n3885), .C2(n3883), .A(n3887), .B(n3825), .ZN(n3824)
         );
  OAI211_X1 U4652 ( .C1(n3821), .C2(n3825), .A(n3888), .B(n3824), .ZN(n3831)
         );
  AOI22_X1 U4653 ( .A1(n3826), .A2(n3937), .B1(REG3_REG_21__SCAN_IN), .B2(
        U3149), .ZN(n3827) );
  OAI21_X1 U4654 ( .B1(n4341), .B2(n3923), .A(n3827), .ZN(n3828) );
  AOI21_X1 U4655 ( .B1(n3829), .B2(n3927), .A(n3828), .ZN(n3830) );
  OAI211_X1 U4656 ( .C1(n3922), .C2(n3832), .A(n3831), .B(n3830), .ZN(U3220)
         );
  INV_X1 U4657 ( .A(n3833), .ZN(n3834) );
  OAI21_X1 U4658 ( .B1(n3840), .B2(n3839), .A(n3838), .ZN(n3841) );
  OAI22_X1 U4659 ( .A1(n4265), .A2(n3920), .B1(STATE_REG_SCAN_IN), .B2(n4988), 
        .ZN(n3842) );
  INV_X1 U4660 ( .A(n3842), .ZN(n3845) );
  NAND2_X1 U4661 ( .A1(n3927), .A2(n3843), .ZN(n3844) );
  OAI211_X1 U4662 ( .C1(n4234), .C2(n3923), .A(n3845), .B(n3844), .ZN(n3846)
         );
  AOI21_X1 U4663 ( .B1(n4274), .B2(n3943), .A(n3846), .ZN(n3847) );
  NAND2_X1 U4664 ( .A1(n3849), .A2(n3848), .ZN(n3857) );
  INV_X1 U4665 ( .A(n3850), .ZN(n3851) );
  NAND2_X1 U4666 ( .A1(n3852), .A2(n3851), .ZN(n3854) );
  NOR2_X1 U4667 ( .A1(n3854), .A2(n3853), .ZN(n3931) );
  INV_X1 U4668 ( .A(n3934), .ZN(n3855) );
  NAND2_X1 U4669 ( .A1(n3854), .A2(n3853), .ZN(n3932) );
  OAI21_X1 U4670 ( .B1(n3931), .B2(n3855), .A(n3932), .ZN(n3856) );
  XOR2_X1 U4671 ( .A(n3857), .B(n3856), .Z(n3858) );
  NAND2_X1 U4672 ( .A1(n3858), .A2(n3888), .ZN(n3862) );
  NAND2_X1 U4673 ( .A1(U3149), .A2(REG3_REG_16__SCAN_IN), .ZN(n4628) );
  OAI21_X1 U4674 ( .B1(n3920), .B2(n4436), .A(n4628), .ZN(n3860) );
  NOR2_X1 U4675 ( .A1(n3941), .A2(n4435), .ZN(n3859) );
  AOI211_X1 U4676 ( .C1(n3938), .C2(n3910), .A(n3860), .B(n3859), .ZN(n3861)
         );
  OAI211_X1 U4677 ( .C1(n3922), .C2(n4448), .A(n3862), .B(n3861), .ZN(U3223)
         );
  NAND2_X1 U4678 ( .A1(n3865), .A2(n3864), .ZN(n3866) );
  XNOR2_X1 U4679 ( .A(n3863), .B(n3866), .ZN(n3871) );
  AND2_X1 U4680 ( .A1(U3149), .A2(REG3_REG_17__SCAN_IN), .ZN(n4640) );
  AOI21_X1 U4681 ( .B1(n3937), .B2(n4416), .A(n4640), .ZN(n3868) );
  NAND2_X1 U4682 ( .A1(n3938), .A2(n4419), .ZN(n3867) );
  OAI211_X1 U4683 ( .C1(n3941), .C2(n4423), .A(n3868), .B(n3867), .ZN(n3869)
         );
  AOI21_X1 U4684 ( .B1(n4430), .B2(n3943), .A(n3869), .ZN(n3870) );
  OAI21_X1 U4685 ( .B1(n3871), .B2(n3945), .A(n3870), .ZN(U3225) );
  INV_X1 U4686 ( .A(n3872), .ZN(n3873) );
  NOR2_X1 U4687 ( .A1(n3874), .A2(n3873), .ZN(n3876) );
  XNOR2_X1 U4688 ( .A(n3876), .B(n3875), .ZN(n3882) );
  INV_X1 U4689 ( .A(n3877), .ZN(n4292) );
  NAND2_X1 U4690 ( .A1(n4286), .A2(n3938), .ZN(n3879) );
  AOI22_X1 U4691 ( .A1(n4326), .A2(n3937), .B1(REG3_REG_24__SCAN_IN), .B2(
        U3149), .ZN(n3878) );
  OAI211_X1 U4692 ( .C1(n3941), .C2(n4290), .A(n3879), .B(n3878), .ZN(n3880)
         );
  AOI21_X1 U4693 ( .B1(n4292), .B2(n3943), .A(n3880), .ZN(n3881) );
  OAI21_X1 U4694 ( .B1(n3882), .B2(n3945), .A(n3881), .ZN(U3226) );
  INV_X1 U4695 ( .A(n4371), .ZN(n3895) );
  NAND2_X1 U4696 ( .A1(n3885), .A2(n3887), .ZN(n3884) );
  NOR2_X1 U4697 ( .A1(n3884), .A2(n3883), .ZN(n3890) );
  AOI21_X1 U4698 ( .B1(n3887), .B2(n3886), .A(n3885), .ZN(n3889) );
  OAI21_X1 U4699 ( .B1(n3890), .B2(n3889), .A(n3888), .ZN(n3894) );
  AOI22_X1 U4700 ( .A1(n3937), .A2(n4398), .B1(REG3_REG_20__SCAN_IN), .B2(
        U3149), .ZN(n3891) );
  OAI21_X1 U4701 ( .B1(n4362), .B2(n3923), .A(n3891), .ZN(n3892) );
  AOI21_X1 U4702 ( .B1(n4360), .B2(n3927), .A(n3892), .ZN(n3893) );
  OAI211_X1 U4703 ( .C1(n3922), .C2(n3895), .A(n3894), .B(n3893), .ZN(U3230)
         );
  INV_X1 U4704 ( .A(n3799), .ZN(n3896) );
  AOI21_X1 U4705 ( .B1(n3898), .B2(n3897), .A(n3896), .ZN(n3905) );
  AOI22_X1 U4706 ( .A1(n4326), .A2(n3938), .B1(REG3_REG_22__SCAN_IN), .B2(
        U3149), .ZN(n3903) );
  INV_X1 U4707 ( .A(n3899), .ZN(n4333) );
  NAND2_X1 U4708 ( .A1(n3943), .A2(n4333), .ZN(n3902) );
  NAND2_X1 U4709 ( .A1(n3927), .A2(n4332), .ZN(n3901) );
  NAND2_X1 U4710 ( .A1(n3937), .A2(n4327), .ZN(n3900) );
  AND4_X1 U4711 ( .A1(n3903), .A2(n3902), .A3(n3901), .A4(n3900), .ZN(n3904)
         );
  OAI21_X1 U4712 ( .B1(n3905), .B2(n3945), .A(n3904), .ZN(U3232) );
  XOR2_X1 U4713 ( .A(n3908), .B(n3907), .Z(n3909) );
  XNOR2_X1 U4714 ( .A(n3906), .B(n3909), .ZN(n3915) );
  AND2_X1 U4715 ( .A1(U3149), .A2(REG3_REG_18__SCAN_IN), .ZN(n4656) );
  AOI21_X1 U4716 ( .B1(n3937), .B2(n3910), .A(n4656), .ZN(n3912) );
  NAND2_X1 U4717 ( .A1(n3938), .A2(n4398), .ZN(n3911) );
  OAI211_X1 U4718 ( .C1(n3941), .C2(n4405), .A(n3912), .B(n3911), .ZN(n3913)
         );
  AOI21_X1 U4719 ( .B1(n4407), .B2(n3943), .A(n3913), .ZN(n3914) );
  OAI21_X1 U4720 ( .B1(n3915), .B2(n3945), .A(n3914), .ZN(U3235) );
  NAND2_X1 U4721 ( .A1(n2152), .A2(n3917), .ZN(n3918) );
  XNOR2_X1 U4722 ( .A(n3916), .B(n3918), .ZN(n3930) );
  OAI22_X1 U4723 ( .A1(n3921), .A2(n3920), .B1(STATE_REG_SCAN_IN), .B2(n3919), 
        .ZN(n3926) );
  OAI22_X1 U4724 ( .A1(n3924), .A2(n3923), .B1(n3922), .B2(n4253), .ZN(n3925)
         );
  AOI211_X1 U4725 ( .C1(n3928), .C2(n3927), .A(n3926), .B(n3925), .ZN(n3929)
         );
  OAI21_X1 U4726 ( .B1(n3930), .B2(n3945), .A(n3929), .ZN(U3237) );
  INV_X1 U4727 ( .A(n3931), .ZN(n3933) );
  NAND2_X1 U4728 ( .A1(n3933), .A2(n3932), .ZN(n3935) );
  XNOR2_X1 U4729 ( .A(n3935), .B(n3934), .ZN(n3946) );
  INV_X1 U4730 ( .A(n3936), .ZN(n4458) );
  AND2_X1 U4731 ( .A1(U3149), .A2(REG3_REG_15__SCAN_IN), .ZN(n4624) );
  AOI21_X1 U4732 ( .B1(n3937), .B2(n4103), .A(n4624), .ZN(n3940) );
  NAND2_X1 U4733 ( .A1(n3938), .A2(n4416), .ZN(n3939) );
  OAI211_X1 U4734 ( .C1(n3941), .C2(n4456), .A(n3940), .B(n3939), .ZN(n3942)
         );
  AOI21_X1 U4735 ( .B1(n4458), .B2(n3943), .A(n3942), .ZN(n3944) );
  OAI21_X1 U4736 ( .B1(n3946), .B2(n3945), .A(n3944), .ZN(U3238) );
  NAND2_X1 U4737 ( .A1(n3949), .A2(n3947), .ZN(n4059) );
  NOR2_X1 U4738 ( .A1(n3948), .A2(n4059), .ZN(n3953) );
  INV_X1 U4739 ( .A(n3949), .ZN(n3952) );
  OAI21_X1 U4740 ( .B1(n3952), .B2(n3951), .A(n3950), .ZN(n4061) );
  OAI21_X1 U4741 ( .B1(n3953), .B2(n4061), .A(n4065), .ZN(n3956) );
  INV_X1 U4742 ( .A(n4070), .ZN(n3954) );
  AOI21_X1 U4743 ( .B1(n3956), .B2(n3955), .A(n3954), .ZN(n3958) );
  INV_X1 U4744 ( .A(n3957), .ZN(n4069) );
  OAI21_X1 U4745 ( .B1(n3958), .B2(n4069), .A(n4072), .ZN(n3960) );
  NAND2_X1 U4746 ( .A1(n3960), .A2(n3959), .ZN(n3962) );
  AOI21_X1 U4747 ( .B1(n3962), .B2(n4075), .A(n3961), .ZN(n3979) );
  INV_X1 U4748 ( .A(n4102), .ZN(n3963) );
  NAND2_X1 U4749 ( .A1(n3963), .A2(n4223), .ZN(n3969) );
  NAND2_X1 U4750 ( .A1(n2606), .A2(REG1_REG_31__SCAN_IN), .ZN(n3967) );
  NAND2_X1 U4751 ( .A1(n3964), .A2(REG2_REG_31__SCAN_IN), .ZN(n3966) );
  NAND2_X1 U4752 ( .A1(n2591), .A2(REG0_REG_31__SCAN_IN), .ZN(n3965) );
  NAND3_X1 U4753 ( .A1(n3967), .A2(n3966), .A3(n3965), .ZN(n4214) );
  NAND2_X1 U4754 ( .A1(n3968), .A2(DATAI_31_), .ZN(n4216) );
  NAND2_X1 U4755 ( .A1(n4214), .A2(n4216), .ZN(n4086) );
  NAND2_X1 U4756 ( .A1(n3969), .A2(n4086), .ZN(n3998) );
  AOI21_X1 U4757 ( .B1(n3971), .B2(n3970), .A(n3998), .ZN(n3975) );
  NAND3_X1 U4758 ( .A1(n3976), .A2(n4076), .A3(n3975), .ZN(n3978) );
  OR2_X1 U4759 ( .A1(n3971), .A2(n3970), .ZN(n3972) );
  NAND2_X1 U4760 ( .A1(n3973), .A2(n3972), .ZN(n4079) );
  NOR3_X1 U4761 ( .A1(n4079), .A2(n4241), .A3(n3974), .ZN(n3977) );
  OAI21_X1 U4762 ( .B1(n3976), .B2(n4079), .A(n3975), .ZN(n4084) );
  OAI22_X1 U4763 ( .A1(n3979), .A2(n3978), .B1(n3977), .B2(n4084), .ZN(n3984)
         );
  INV_X1 U4764 ( .A(n4214), .ZN(n3980) );
  NAND2_X1 U4765 ( .A1(n3980), .A2(n4223), .ZN(n3983) );
  INV_X1 U4766 ( .A(n4223), .ZN(n3981) );
  NAND2_X1 U4767 ( .A1(n3981), .A2(n4102), .ZN(n3997) );
  AOI21_X1 U4768 ( .B1(n3997), .B2(n4214), .A(n4216), .ZN(n3982) );
  AOI21_X1 U4769 ( .B1(n3984), .B2(n3983), .A(n3982), .ZN(n4093) );
  INV_X1 U4770 ( .A(n4299), .ZN(n3985) );
  NAND2_X1 U4771 ( .A1(n3985), .A2(n4300), .ZN(n4340) );
  NAND2_X1 U4772 ( .A1(n3987), .A2(n3986), .ZN(n4387) );
  INV_X1 U4773 ( .A(n4387), .ZN(n3990) );
  NAND3_X1 U4774 ( .A1(n3990), .A2(n3989), .A3(n3988), .ZN(n3991) );
  NAND2_X1 U4775 ( .A1(n4376), .A2(n4066), .ZN(n4424) );
  NOR4_X1 U4776 ( .A1(n4340), .A2(n4320), .A3(n3991), .A4(n4424), .ZN(n4016)
         );
  NAND2_X1 U4777 ( .A1(n3992), .A2(n4260), .ZN(n4282) );
  INV_X1 U4778 ( .A(n4282), .ZN(n4014) );
  NAND2_X1 U4779 ( .A1(n4280), .A2(n3993), .ZN(n4303) );
  OAI21_X1 U4780 ( .B1(n4214), .B2(n4216), .A(n3997), .ZN(n4085) );
  NOR3_X1 U4781 ( .A1(n3999), .A2(n3998), .A3(n4085), .ZN(n4002) );
  NAND4_X1 U4782 ( .A1(n4003), .A2(n4002), .A3(n4001), .A4(n4000), .ZN(n4009)
         );
  NAND4_X1 U4783 ( .A1(n4007), .A2(n4006), .A3(n4005), .A4(n4004), .ZN(n4008)
         );
  OR4_X1 U4784 ( .A1(n4403), .A2(n4469), .A3(n4009), .A4(n4008), .ZN(n4010) );
  NOR4_X1 U4785 ( .A1(n4303), .A2(n4012), .A3(n4011), .A4(n4010), .ZN(n4013)
         );
  NAND4_X1 U4786 ( .A1(n4016), .A2(n4015), .A3(n4014), .A4(n4013), .ZN(n4019)
         );
  NAND2_X1 U4787 ( .A1(n4018), .A2(n4017), .ZN(n4262) );
  XNOR2_X1 U4788 ( .A(n4385), .B(n4360), .ZN(n4358) );
  NOR4_X1 U4789 ( .A1(n4020), .A2(n4019), .A3(n4262), .A4(n4358), .ZN(n4021)
         );
  NAND4_X1 U4790 ( .A1(n4022), .A2(n4484), .A3(n3190), .A4(n4021), .ZN(n4024)
         );
  NAND2_X1 U4791 ( .A1(n4024), .A2(n4023), .ZN(n4090) );
  OAI211_X1 U4792 ( .C1(n4027), .C2(n4591), .A(n4025), .B(n4026), .ZN(n4030)
         );
  NAND3_X1 U4793 ( .A1(n4030), .A2(n4029), .A3(n4028), .ZN(n4033) );
  NAND3_X1 U4794 ( .A1(n4033), .A2(n4031), .A3(n4032), .ZN(n4036) );
  NAND3_X1 U4795 ( .A1(n4036), .A2(n4035), .A3(n4034), .ZN(n4038) );
  NAND3_X1 U4796 ( .A1(n4038), .A2(n4037), .A3(n2247), .ZN(n4042) );
  INV_X1 U4797 ( .A(n4039), .ZN(n4040) );
  AOI21_X1 U4798 ( .B1(n4042), .B2(n4041), .A(n4040), .ZN(n4048) );
  NAND2_X1 U4799 ( .A1(n4044), .A2(n4043), .ZN(n4047) );
  OAI211_X1 U4800 ( .C1(n4048), .C2(n4047), .A(n4046), .B(n4045), .ZN(n4051)
         );
  AND3_X1 U4801 ( .A1(n4051), .A2(n4050), .A3(n4049), .ZN(n4054) );
  OAI21_X1 U4802 ( .B1(n4054), .B2(n4053), .A(n4052), .ZN(n4057) );
  NAND3_X1 U4803 ( .A1(n4057), .A2(n4056), .A3(n4055), .ZN(n4064) );
  INV_X1 U4804 ( .A(n4058), .ZN(n4060) );
  NOR2_X1 U4805 ( .A1(n4060), .A2(n4059), .ZN(n4063) );
  INV_X1 U4806 ( .A(n4412), .ZN(n4062) );
  AOI211_X1 U4807 ( .C1(n4064), .C2(n4063), .A(n4062), .B(n4061), .ZN(n4068)
         );
  INV_X1 U4808 ( .A(n4065), .ZN(n4067) );
  OAI21_X1 U4809 ( .B1(n4068), .B2(n4067), .A(n4066), .ZN(n4071) );
  AOI211_X1 U4810 ( .C1(n4071), .C2(n4070), .A(n4299), .B(n4069), .ZN(n4074)
         );
  INV_X1 U4811 ( .A(n4072), .ZN(n4073) );
  NOR2_X1 U4812 ( .A1(n4074), .A2(n4073), .ZN(n4078) );
  OAI211_X1 U4813 ( .C1(n4078), .C2(n4077), .A(n4076), .B(n4075), .ZN(n4083)
         );
  INV_X1 U4814 ( .A(n4079), .ZN(n4081) );
  NAND4_X1 U4815 ( .A1(n4083), .A2(n4082), .A3(n4081), .A4(n4080), .ZN(n4088)
         );
  INV_X1 U4816 ( .A(n4084), .ZN(n4087) );
  AOI22_X1 U4817 ( .A1(n4088), .A2(n4087), .B1(n4086), .B2(n4085), .ZN(n4089)
         );
  MUX2_X1 U4818 ( .A(n4090), .B(n4089), .S(n2816), .Z(n4091) );
  OAI21_X1 U4819 ( .B1(n4093), .B2(n4092), .A(n4091), .ZN(n4095) );
  XNOR2_X1 U4820 ( .A(n4095), .B(n4094), .ZN(n4101) );
  NOR2_X1 U4821 ( .A1(n4097), .A2(n4096), .ZN(n4099) );
  OAI21_X1 U4822 ( .B1(n4100), .B2(n2895), .A(B_REG_SCAN_IN), .ZN(n4098) );
  OAI22_X1 U4823 ( .A1(n4101), .A2(n4100), .B1(n4099), .B2(n4098), .ZN(U3239)
         );
  MUX2_X1 U4824 ( .A(DATAO_REG_31__SCAN_IN), .B(n4214), .S(n4109), .Z(U3581)
         );
  MUX2_X1 U4825 ( .A(DATAO_REG_30__SCAN_IN), .B(n4102), .S(n4109), .Z(U3580)
         );
  MUX2_X1 U4826 ( .A(DATAO_REG_28__SCAN_IN), .B(n4239), .S(n4109), .Z(U3578)
         );
  MUX2_X1 U4827 ( .A(DATAO_REG_26__SCAN_IN), .B(n4267), .S(n4109), .Z(U3576)
         );
  MUX2_X1 U4828 ( .A(DATAO_REG_25__SCAN_IN), .B(n4286), .S(n4109), .Z(U3575)
         );
  MUX2_X1 U4829 ( .A(DATAO_REG_24__SCAN_IN), .B(n4306), .S(n4109), .Z(U3574)
         );
  MUX2_X1 U4830 ( .A(DATAO_REG_21__SCAN_IN), .B(n4327), .S(n4109), .Z(U3571)
         );
  MUX2_X1 U4831 ( .A(n4398), .B(DATAO_REG_19__SCAN_IN), .S(n3439), .Z(U3569)
         );
  MUX2_X1 U4832 ( .A(DATAO_REG_16__SCAN_IN), .B(n4416), .S(n4109), .Z(U3566)
         );
  MUX2_X1 U4833 ( .A(DATAO_REG_14__SCAN_IN), .B(n4103), .S(n4109), .Z(U3564)
         );
  MUX2_X1 U4834 ( .A(DATAO_REG_13__SCAN_IN), .B(n4104), .S(n4109), .Z(U3563)
         );
  MUX2_X1 U4835 ( .A(DATAO_REG_11__SCAN_IN), .B(n4105), .S(n4109), .Z(U3561)
         );
  MUX2_X1 U4836 ( .A(DATAO_REG_9__SCAN_IN), .B(n4106), .S(n4109), .Z(U3559) );
  MUX2_X1 U4837 ( .A(DATAO_REG_7__SCAN_IN), .B(n4107), .S(n4109), .Z(U3557) );
  MUX2_X1 U4838 ( .A(DATAO_REG_5__SCAN_IN), .B(n4108), .S(n4109), .Z(U3555) );
  MUX2_X1 U4839 ( .A(DATAO_REG_3__SCAN_IN), .B(n4110), .S(n4109), .Z(U3553) );
  MUX2_X1 U4840 ( .A(DATAO_REG_1__SCAN_IN), .B(n2601), .S(U4043), .Z(U3551) );
  MUX2_X1 U4841 ( .A(DATAO_REG_0__SCAN_IN), .B(n4111), .S(U4043), .Z(U3550) );
  OAI211_X1 U4842 ( .C1(n4114), .C2(n4113), .A(n4664), .B(n4112), .ZN(n4122)
         );
  MUX2_X1 U4843 ( .A(n2500), .B(REG1_REG_1__SCAN_IN), .S(n2127), .Z(n4115) );
  OAI21_X1 U4844 ( .B1(n4685), .B2(n4116), .A(n4115), .ZN(n4117) );
  NAND3_X1 U4845 ( .A1(n4648), .A2(n4118), .A3(n4117), .ZN(n4121) );
  INV_X1 U4846 ( .A(n4668), .ZN(n4623) );
  NAND2_X1 U4847 ( .A1(n4623), .A2(n2127), .ZN(n4120) );
  AOI22_X1 U4848 ( .A1(n4657), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n4119) );
  NAND4_X1 U4849 ( .A1(n4122), .A2(n4121), .A3(n4120), .A4(n4119), .ZN(U3241)
         );
  OAI211_X1 U4850 ( .C1(REG2_REG_3__SCAN_IN), .C2(n4124), .A(n4664), .B(n4123), 
        .ZN(n4130) );
  NAND2_X1 U4851 ( .A1(n4623), .A2(n4603), .ZN(n4129) );
  XOR2_X1 U4852 ( .A(n4125), .B(REG1_REG_3__SCAN_IN), .Z(n4126) );
  NAND2_X1 U4853 ( .A1(n4648), .A2(n4126), .ZN(n4128) );
  AOI22_X1 U4854 ( .A1(n4657), .A2(ADDR_REG_3__SCAN_IN), .B1(
        REG3_REG_3__SCAN_IN), .B2(U3149), .ZN(n4127) );
  NAND4_X1 U4855 ( .A1(n4130), .A2(n4129), .A3(n4128), .A4(n4127), .ZN(U3243)
         );
  NOR2_X1 U4856 ( .A1(n4668), .A2(n4131), .ZN(n4132) );
  AOI211_X1 U4857 ( .C1(n4657), .C2(ADDR_REG_5__SCAN_IN), .A(n4133), .B(n4132), 
        .ZN(n4142) );
  OAI211_X1 U4858 ( .C1(n4136), .C2(n4135), .A(n4664), .B(n4134), .ZN(n4141)
         );
  OAI211_X1 U4859 ( .C1(n4139), .C2(n4138), .A(n4648), .B(n4137), .ZN(n4140)
         );
  NAND3_X1 U4860 ( .A1(n4142), .A2(n4141), .A3(n4140), .ZN(U3245) );
  OAI211_X1 U4861 ( .C1(n4144), .C2(REG2_REG_8__SCAN_IN), .A(n4143), .B(n4664), 
        .ZN(n4153) );
  INV_X1 U4862 ( .A(n4145), .ZN(n4148) );
  NOR2_X1 U4863 ( .A1(n4668), .A2(n4146), .ZN(n4147) );
  AOI211_X1 U4864 ( .C1(n4657), .C2(ADDR_REG_8__SCAN_IN), .A(n4148), .B(n4147), 
        .ZN(n4152) );
  OAI211_X1 U4865 ( .C1(n4150), .C2(REG1_REG_8__SCAN_IN), .A(n4149), .B(n4648), 
        .ZN(n4151) );
  NAND3_X1 U4866 ( .A1(n4153), .A2(n4152), .A3(n4151), .ZN(U3248) );
  OAI211_X1 U4867 ( .C1(n4156), .C2(n4155), .A(n4154), .B(n4664), .ZN(n4165)
         );
  INV_X1 U4868 ( .A(n4157), .ZN(n4158) );
  AOI21_X1 U4869 ( .B1(n4657), .B2(ADDR_REG_9__SCAN_IN), .A(n4158), .ZN(n4164)
         );
  OAI211_X1 U4870 ( .C1(n4161), .C2(n4160), .A(n4159), .B(n4648), .ZN(n4163)
         );
  NAND2_X1 U4871 ( .A1(n4623), .A2(n4598), .ZN(n4162) );
  NAND4_X1 U4872 ( .A1(n4165), .A2(n4164), .A3(n4163), .A4(n4162), .ZN(U3249)
         );
  OAI211_X1 U4873 ( .C1(n4167), .C2(REG2_REG_10__SCAN_IN), .A(n4166), .B(n4664), .ZN(n4176) );
  INV_X1 U4874 ( .A(n4168), .ZN(n4169) );
  AOI21_X1 U4875 ( .B1(n4657), .B2(ADDR_REG_10__SCAN_IN), .A(n4169), .ZN(n4175) );
  OAI211_X1 U4876 ( .C1(n4171), .C2(REG1_REG_10__SCAN_IN), .A(n4170), .B(n4648), .ZN(n4174) );
  OR2_X1 U4877 ( .A1(n4668), .A2(n4172), .ZN(n4173) );
  NAND4_X1 U4878 ( .A1(n4176), .A2(n4175), .A3(n4174), .A4(n4173), .ZN(U3250)
         );
  OAI211_X1 U4879 ( .C1(n4179), .C2(n4178), .A(n4177), .B(n4664), .ZN(n4189)
         );
  INV_X1 U4880 ( .A(n4180), .ZN(n4181) );
  AOI21_X1 U4881 ( .B1(n4657), .B2(ADDR_REG_11__SCAN_IN), .A(n4181), .ZN(n4188) );
  OAI211_X1 U4882 ( .C1(n4184), .C2(n4183), .A(n4182), .B(n4648), .ZN(n4187)
         );
  OR2_X1 U4883 ( .A1(n4668), .A2(n4185), .ZN(n4186) );
  NAND4_X1 U4884 ( .A1(n4189), .A2(n4188), .A3(n4187), .A4(n4186), .ZN(U3251)
         );
  OAI211_X1 U4885 ( .C1(n4191), .C2(REG2_REG_12__SCAN_IN), .A(n4190), .B(n4664), .ZN(n4199) );
  INV_X1 U4886 ( .A(n4192), .ZN(n4193) );
  AOI21_X1 U4887 ( .B1(n4657), .B2(ADDR_REG_12__SCAN_IN), .A(n4193), .ZN(n4198) );
  OR2_X1 U4888 ( .A1(n4668), .A2(n4195), .ZN(n4196) );
  NAND4_X1 U4889 ( .A1(n4199), .A2(n4198), .A3(n4197), .A4(n4196), .ZN(U3252)
         );
  AND2_X1 U4890 ( .A1(n4201), .A2(n4200), .ZN(n4203) );
  AOI21_X1 U4891 ( .B1(REG2_REG_13__SCAN_IN), .B2(n4203), .A(n4615), .ZN(n4202) );
  OAI21_X1 U4892 ( .B1(n4203), .B2(REG2_REG_13__SCAN_IN), .A(n4202), .ZN(n4213) );
  INV_X1 U4893 ( .A(n4204), .ZN(n4205) );
  AOI21_X1 U4894 ( .B1(n4657), .B2(ADDR_REG_13__SCAN_IN), .A(n4205), .ZN(n4212) );
  OAI211_X1 U4895 ( .C1(n4208), .C2(n4207), .A(n4206), .B(n4648), .ZN(n4211)
         );
  OR2_X1 U4896 ( .A1(n4668), .A2(n4209), .ZN(n4210) );
  NAND4_X1 U4897 ( .A1(n4213), .A2(n4212), .A3(n4211), .A4(n4210), .ZN(U3253)
         );
  NAND2_X1 U4898 ( .A1(n4215), .A2(n4214), .ZN(n4220) );
  OAI21_X1 U4899 ( .B1(n4216), .B2(n4422), .A(n4220), .ZN(n4550) );
  NAND2_X1 U4900 ( .A1(n4351), .A2(n4550), .ZN(n4218) );
  NAND2_X1 U4901 ( .A1(n4459), .A2(REG2_REG_31__SCAN_IN), .ZN(n4217) );
  OAI211_X1 U4902 ( .C1(n4553), .C2(n4461), .A(n4218), .B(n4217), .ZN(U3260)
         );
  NAND2_X1 U4903 ( .A1(n4473), .A2(n4223), .ZN(n4219) );
  AOI21_X1 U4904 ( .B1(n4223), .B2(n4222), .A(n4221), .ZN(n4555) );
  NAND2_X1 U4905 ( .A1(n4555), .A2(n4674), .ZN(n4225) );
  NAND2_X1 U4906 ( .A1(n4459), .A2(REG2_REG_30__SCAN_IN), .ZN(n4224) );
  OAI211_X1 U4907 ( .C1(n4459), .C2(n4558), .A(n4225), .B(n4224), .ZN(U3261)
         );
  AOI22_X1 U4908 ( .A1(n4226), .A2(n4669), .B1(REG2_REG_28__SCAN_IN), .B2(
        n4459), .ZN(n4229) );
  OAI211_X1 U4909 ( .C1(n4230), .C2(n4461), .A(n4229), .B(n4228), .ZN(n4231)
         );
  AOI21_X1 U4910 ( .B1(n4232), .B2(n4477), .A(n4231), .ZN(n4233) );
  INV_X1 U4911 ( .A(n4233), .ZN(U3262) );
  OAI22_X1 U4912 ( .A1(n4234), .A2(n4462), .B1(n4422), .B2(n4243), .ZN(n4238)
         );
  NAND2_X1 U4913 ( .A1(n4235), .A2(n4241), .ZN(n4236) );
  AOI21_X1 U4914 ( .B1(n3213), .B2(n4236), .A(n4468), .ZN(n4237) );
  XNOR2_X1 U4915 ( .A(n4240), .B(n4241), .ZN(n4497) );
  NAND2_X1 U4916 ( .A1(n4497), .A2(n4477), .ZN(n4250) );
  OAI21_X1 U4917 ( .B1(n4244), .B2(n4243), .A(n4242), .ZN(n4498) );
  INV_X1 U4918 ( .A(n4498), .ZN(n4248) );
  INV_X1 U4919 ( .A(REG2_REG_27__SCAN_IN), .ZN(n4245) );
  OAI22_X1 U4920 ( .A1(n4246), .A2(n4447), .B1(n4245), .B2(n4351), .ZN(n4247)
         );
  AOI21_X1 U4921 ( .B1(n4248), .B2(n4674), .A(n4247), .ZN(n4249) );
  OAI211_X1 U4922 ( .C1(n4500), .C2(n4459), .A(n4250), .B(n4249), .ZN(U3263)
         );
  INV_X1 U4923 ( .A(n4251), .ZN(n4258) );
  INV_X1 U4924 ( .A(REG2_REG_26__SCAN_IN), .ZN(n4252) );
  OAI22_X1 U4925 ( .A1(n4253), .A2(n4447), .B1(n4252), .B2(n4351), .ZN(n4255)
         );
  NOR2_X1 U4926 ( .A1(n4505), .A2(n4461), .ZN(n4254) );
  AOI211_X1 U4927 ( .C1(n4256), .C2(n4351), .A(n4255), .B(n4254), .ZN(n4257)
         );
  OAI21_X1 U4928 ( .B1(n4258), .B2(n4452), .A(n4257), .ZN(U3264) );
  XNOR2_X1 U4929 ( .A(n4259), .B(n4262), .ZN(n4507) );
  INV_X1 U4930 ( .A(n4507), .ZN(n4278) );
  NAND2_X1 U4931 ( .A1(n4261), .A2(n4260), .ZN(n4263) );
  XNOR2_X1 U4932 ( .A(n4263), .B(n4262), .ZN(n4264) );
  NAND2_X1 U4933 ( .A1(n4264), .A2(n4414), .ZN(n4269) );
  OAI22_X1 U4934 ( .A1(n4265), .A2(n4462), .B1(n4422), .B2(n4272), .ZN(n4266)
         );
  AOI21_X1 U4935 ( .B1(n4267), .B2(n4418), .A(n4266), .ZN(n4268) );
  NAND2_X1 U4936 ( .A1(n4269), .A2(n4268), .ZN(n4506) );
  INV_X1 U4937 ( .A(n4270), .ZN(n4273) );
  OAI21_X1 U4938 ( .B1(n4273), .B2(n4272), .A(n4271), .ZN(n4562) );
  AOI22_X1 U4939 ( .A1(n4274), .A2(n4669), .B1(REG2_REG_25__SCAN_IN), .B2(
        n4459), .ZN(n4275) );
  OAI21_X1 U4940 ( .B1(n4562), .B2(n4461), .A(n4275), .ZN(n4276) );
  AOI21_X1 U4941 ( .B1(n4316), .B2(n4506), .A(n4276), .ZN(n4277) );
  OAI21_X1 U4942 ( .B1(n4278), .B2(n4452), .A(n4277), .ZN(U3265) );
  XOR2_X1 U4943 ( .A(n4282), .B(n4279), .Z(n4511) );
  INV_X1 U4944 ( .A(n4511), .ZN(n4296) );
  NAND2_X1 U4945 ( .A1(n4281), .A2(n4280), .ZN(n4283) );
  XNOR2_X1 U4946 ( .A(n4283), .B(n4282), .ZN(n4288) );
  OAI22_X1 U4947 ( .A1(n4284), .A2(n4462), .B1(n4422), .B2(n4290), .ZN(n4285)
         );
  AOI21_X1 U4948 ( .B1(n4286), .B2(n4418), .A(n4285), .ZN(n4287) );
  OAI21_X1 U4949 ( .B1(n4288), .B2(n4468), .A(n4287), .ZN(n4510) );
  OR2_X1 U4950 ( .A1(n4289), .A2(n4290), .ZN(n4291) );
  NAND2_X1 U4951 ( .A1(n4270), .A2(n4291), .ZN(n4566) );
  AOI22_X1 U4952 ( .A1(n4292), .A2(n4669), .B1(REG2_REG_24__SCAN_IN), .B2(
        n4459), .ZN(n4293) );
  OAI21_X1 U4953 ( .B1(n4566), .B2(n4461), .A(n4293), .ZN(n4294) );
  AOI21_X1 U4954 ( .B1(n4316), .B2(n4510), .A(n4294), .ZN(n4295) );
  OAI21_X1 U4955 ( .B1(n4296), .B2(n4452), .A(n4295), .ZN(U3266) );
  XOR2_X1 U4956 ( .A(n4303), .B(n4297), .Z(n4515) );
  INV_X1 U4957 ( .A(n4515), .ZN(n4318) );
  OR2_X1 U4958 ( .A1(n4298), .A2(n4299), .ZN(n4301) );
  NAND2_X1 U4959 ( .A1(n4301), .A2(n4300), .ZN(n4323) );
  INV_X1 U4960 ( .A(n4320), .ZN(n4322) );
  NAND2_X1 U4961 ( .A1(n4323), .A2(n4322), .ZN(n4325) );
  NAND2_X1 U4962 ( .A1(n4325), .A2(n4302), .ZN(n4304) );
  XNOR2_X1 U4963 ( .A(n4304), .B(n4303), .ZN(n4308) );
  OAI22_X1 U4964 ( .A1(n4341), .A2(n4462), .B1(n4422), .B2(n4313), .ZN(n4305)
         );
  AOI21_X1 U4965 ( .B1(n4306), .B2(n4418), .A(n4305), .ZN(n4307) );
  OAI21_X1 U4966 ( .B1(n4308), .B2(n4468), .A(n4307), .ZN(n4514) );
  INV_X1 U4967 ( .A(REG2_REG_23__SCAN_IN), .ZN(n4310) );
  OAI22_X1 U4968 ( .A1(n4351), .A2(n4310), .B1(n4309), .B2(n4447), .ZN(n4315)
         );
  INV_X1 U4969 ( .A(n4289), .ZN(n4312) );
  OAI21_X1 U4970 ( .B1(n4311), .B2(n4313), .A(n4312), .ZN(n4570) );
  NOR2_X1 U4971 ( .A1(n4570), .A2(n4461), .ZN(n4314) );
  AOI211_X1 U4972 ( .C1(n4316), .C2(n4514), .A(n4315), .B(n4314), .ZN(n4317)
         );
  OAI21_X1 U4973 ( .B1(n4318), .B2(n4452), .A(n4317), .ZN(U3267) );
  OAI21_X1 U4974 ( .B1(n4321), .B2(n4320), .A(n4319), .ZN(n4521) );
  OR2_X1 U4975 ( .A1(n4323), .A2(n4322), .ZN(n4324) );
  NAND2_X1 U4976 ( .A1(n4325), .A2(n4324), .ZN(n4331) );
  NAND2_X1 U4977 ( .A1(n4326), .A2(n4418), .ZN(n4329) );
  AOI22_X1 U4978 ( .A1(n4327), .A2(n4417), .B1(n4473), .B2(n4332), .ZN(n4328)
         );
  NAND2_X1 U4979 ( .A1(n4329), .A2(n4328), .ZN(n4330) );
  AOI21_X1 U4980 ( .B1(n4331), .B2(n4414), .A(n4330), .ZN(n4520) );
  INV_X1 U4981 ( .A(n4520), .ZN(n4337) );
  NAND2_X1 U4982 ( .A1(n4347), .A2(n4332), .ZN(n4517) );
  NAND2_X1 U4983 ( .A1(n4517), .A2(n4674), .ZN(n4335) );
  AOI22_X1 U4984 ( .A1(REG2_REG_22__SCAN_IN), .A2(n4459), .B1(n4333), .B2(
        n4669), .ZN(n4334) );
  OAI21_X1 U4985 ( .B1(n4311), .B2(n4335), .A(n4334), .ZN(n4336) );
  AOI21_X1 U4986 ( .B1(n4337), .B2(n4351), .A(n4336), .ZN(n4338) );
  OAI21_X1 U4987 ( .B1(n4521), .B2(n4452), .A(n4338), .ZN(U3268) );
  XNOR2_X1 U4988 ( .A(n4339), .B(n4340), .ZN(n4523) );
  INV_X1 U4989 ( .A(n4523), .ZN(n4353) );
  XNOR2_X1 U4990 ( .A(n4298), .B(n4340), .ZN(n4344) );
  NOR2_X1 U4991 ( .A1(n4385), .A2(n4462), .ZN(n4343) );
  OAI22_X1 U4992 ( .A1(n4341), .A2(n4464), .B1(n4422), .B2(n2882), .ZN(n4342)
         );
  AOI211_X1 U4993 ( .C1(n4344), .C2(n4414), .A(n4343), .B(n4342), .ZN(n4345)
         );
  INV_X1 U4994 ( .A(n4345), .ZN(n4522) );
  OAI21_X1 U4995 ( .B1(n4346), .B2(n2882), .A(n4347), .ZN(n4575) );
  AOI22_X1 U4996 ( .A1(n4459), .A2(REG2_REG_21__SCAN_IN), .B1(n4348), .B2(
        n4669), .ZN(n4349) );
  OAI21_X1 U4997 ( .B1(n4575), .B2(n4461), .A(n4349), .ZN(n4350) );
  AOI21_X1 U4998 ( .B1(n4522), .B2(n4351), .A(n4350), .ZN(n4352) );
  OAI21_X1 U4999 ( .B1(n4353), .B2(n4452), .A(n4352), .ZN(U3269) );
  XNOR2_X1 U5000 ( .A(n2156), .B(n4358), .ZN(n4367) );
  INV_X1 U5001 ( .A(n4354), .ZN(n4357) );
  AOI21_X1 U5002 ( .B1(n4357), .B2(n4356), .A(n4355), .ZN(n4359) );
  XNOR2_X1 U5003 ( .A(n4359), .B(n4358), .ZN(n4364) );
  AOI22_X1 U5004 ( .A1(n4398), .A2(n4417), .B1(n4473), .B2(n4360), .ZN(n4361)
         );
  OAI21_X1 U5005 ( .B1(n4362), .B2(n4464), .A(n4361), .ZN(n4363) );
  AOI21_X1 U5006 ( .B1(n4364), .B2(n4414), .A(n4363), .ZN(n4365) );
  OAI21_X1 U5007 ( .B1(n4367), .B2(n4366), .A(n4365), .ZN(n4525) );
  INV_X1 U5008 ( .A(n4525), .ZN(n4375) );
  INV_X1 U5009 ( .A(n4367), .ZN(n4526) );
  INV_X1 U5010 ( .A(n4368), .ZN(n4370) );
  OAI21_X1 U5011 ( .B1(n4370), .B2(n4369), .A(n2222), .ZN(n4579) );
  AOI22_X1 U5012 ( .A1(n4459), .A2(REG2_REG_20__SCAN_IN), .B1(n4371), .B2(
        n4669), .ZN(n4372) );
  OAI21_X1 U5013 ( .B1(n4579), .B2(n4461), .A(n4372), .ZN(n4373) );
  AOI21_X1 U5014 ( .B1(n4526), .B2(n4672), .A(n4373), .ZN(n4374) );
  OAI21_X1 U5015 ( .B1(n4375), .B2(n4459), .A(n4374), .ZN(U3270) );
  NAND2_X1 U5016 ( .A1(n4354), .A2(n4376), .ZN(n4396) );
  INV_X1 U5017 ( .A(n4377), .ZN(n4379) );
  OAI21_X1 U5018 ( .B1(n4396), .B2(n4379), .A(n4378), .ZN(n4380) );
  XNOR2_X1 U5019 ( .A(n4380), .B(n4387), .ZN(n4381) );
  NAND2_X1 U5020 ( .A1(n4381), .A2(n4414), .ZN(n4384) );
  AOI22_X1 U5021 ( .A1(n4419), .A2(n4417), .B1(n4473), .B2(n4382), .ZN(n4383)
         );
  OAI211_X1 U5022 ( .C1(n4385), .C2(n4464), .A(n4384), .B(n4383), .ZN(n4528)
         );
  INV_X1 U5023 ( .A(n4528), .ZN(n4395) );
  XNOR2_X1 U5024 ( .A(n4386), .B(n4387), .ZN(n4529) );
  OR2_X1 U5025 ( .A1(n4389), .A2(n4388), .ZN(n4390) );
  NAND2_X1 U5026 ( .A1(n4368), .A2(n4390), .ZN(n4582) );
  NOR2_X1 U5027 ( .A1(n4582), .A2(n4461), .ZN(n4393) );
  OAI22_X1 U5028 ( .A1(n4351), .A2(n2462), .B1(n4391), .B2(n4447), .ZN(n4392)
         );
  AOI211_X1 U5029 ( .C1(n4529), .C2(n4477), .A(n4393), .B(n4392), .ZN(n4394)
         );
  OAI21_X1 U5030 ( .B1(n4459), .B2(n4395), .A(n4394), .ZN(U3271) );
  XOR2_X1 U5031 ( .A(n4403), .B(n4396), .Z(n4401) );
  AOI22_X1 U5032 ( .A1(n4398), .A2(n4418), .B1(n4473), .B2(n4397), .ZN(n4399)
         );
  OAI21_X1 U5033 ( .B1(n4437), .B2(n4462), .A(n4399), .ZN(n4400) );
  AOI21_X1 U5034 ( .B1(n4401), .B2(n4414), .A(n4400), .ZN(n4534) );
  OAI21_X1 U5035 ( .B1(n4404), .B2(n4403), .A(n4402), .ZN(n4532) );
  XNOR2_X1 U5036 ( .A(n4429), .B(n4405), .ZN(n4406) );
  NAND2_X1 U5037 ( .A1(n4406), .A2(n4698), .ZN(n4533) );
  AOI22_X1 U5038 ( .A1(n4459), .A2(REG2_REG_18__SCAN_IN), .B1(n4407), .B2(
        n4669), .ZN(n4408) );
  OAI21_X1 U5039 ( .B1(n4533), .B2(n4409), .A(n4408), .ZN(n4410) );
  AOI21_X1 U5040 ( .B1(n4532), .B2(n4477), .A(n4410), .ZN(n4411) );
  OAI21_X1 U5041 ( .B1(n4459), .B2(n4534), .A(n4411), .ZN(U3272) );
  NAND2_X1 U5042 ( .A1(n4439), .A2(n4412), .ZN(n4413) );
  XNOR2_X1 U5043 ( .A(n4413), .B(n4424), .ZN(n4415) );
  NAND2_X1 U5044 ( .A1(n4415), .A2(n4414), .ZN(n4421) );
  AOI22_X1 U5045 ( .A1(n4419), .A2(n4418), .B1(n4417), .B2(n4416), .ZN(n4420)
         );
  OAI211_X1 U5046 ( .C1(n4423), .C2(n4422), .A(n4421), .B(n4420), .ZN(n4536)
         );
  INV_X1 U5047 ( .A(n4536), .ZN(n4434) );
  XOR2_X1 U5048 ( .A(n4425), .B(n4424), .Z(n4537) );
  NAND2_X1 U5049 ( .A1(n4426), .A2(n4427), .ZN(n4428) );
  NAND2_X1 U5050 ( .A1(n4429), .A2(n4428), .ZN(n4587) );
  AOI22_X1 U5051 ( .A1(n4459), .A2(REG2_REG_17__SCAN_IN), .B1(n4430), .B2(
        n4669), .ZN(n4431) );
  OAI21_X1 U5052 ( .B1(n4587), .B2(n4461), .A(n4431), .ZN(n4432) );
  AOI21_X1 U5053 ( .B1(n4537), .B2(n4477), .A(n4432), .ZN(n4433) );
  OAI21_X1 U5054 ( .B1(n4459), .B2(n4434), .A(n4433), .ZN(U3273) );
  OAI22_X1 U5055 ( .A1(n4437), .A2(n4464), .B1(n4436), .B2(n4462), .ZN(n4443)
         );
  INV_X1 U5056 ( .A(n4438), .ZN(n4441) );
  INV_X1 U5057 ( .A(n4439), .ZN(n4440) );
  AOI211_X1 U5058 ( .C1(n4441), .C2(n4450), .A(n4468), .B(n4440), .ZN(n4442)
         );
  AOI211_X1 U5059 ( .C1(n2727), .C2(n4473), .A(n4443), .B(n4442), .ZN(n4543)
         );
  INV_X1 U5060 ( .A(n4444), .ZN(n4446) );
  INV_X1 U5061 ( .A(n4426), .ZN(n4445) );
  AOI21_X1 U5062 ( .B1(n2727), .B2(n4446), .A(n4445), .ZN(n4541) );
  OAI22_X1 U5063 ( .A1(n4351), .A2(n4631), .B1(n4448), .B2(n4447), .ZN(n4454)
         );
  OAI21_X1 U5064 ( .B1(n4451), .B2(n4450), .A(n4449), .ZN(n4544) );
  NOR2_X1 U5065 ( .A1(n4544), .A2(n4452), .ZN(n4453) );
  AOI211_X1 U5066 ( .C1(n4541), .C2(n4674), .A(n4454), .B(n4453), .ZN(n4455)
         );
  OAI21_X1 U5067 ( .B1(n4459), .B2(n4543), .A(n4455), .ZN(U3274) );
  XOR2_X1 U5068 ( .A(n2160), .B(n4469), .Z(n4546) );
  XNOR2_X1 U5069 ( .A(n4457), .B(n4456), .ZN(n4549) );
  AOI22_X1 U5070 ( .A1(n4459), .A2(REG2_REG_15__SCAN_IN), .B1(n4458), .B2(
        n4669), .ZN(n4460) );
  OAI21_X1 U5071 ( .B1(n4549), .B2(n4461), .A(n4460), .ZN(n4476) );
  OAI22_X1 U5072 ( .A1(n4465), .A2(n4464), .B1(n4463), .B2(n4462), .ZN(n4472)
         );
  INV_X1 U5073 ( .A(n4466), .ZN(n4467) );
  AOI211_X1 U5074 ( .C1(n4470), .C2(n4469), .A(n4468), .B(n4467), .ZN(n4471)
         );
  AOI211_X1 U5075 ( .C1(n4474), .C2(n4473), .A(n4472), .B(n4471), .ZN(n4548)
         );
  NOR2_X1 U5076 ( .A1(n4548), .A2(n4459), .ZN(n4475) );
  AOI211_X1 U5077 ( .C1(n4477), .C2(n4546), .A(n4476), .B(n4475), .ZN(n4478)
         );
  INV_X1 U5078 ( .A(n4478), .ZN(U3275) );
  NAND2_X1 U5079 ( .A1(n4725), .A2(n4550), .ZN(n4480) );
  NAND2_X1 U5080 ( .A1(n3232), .A2(REG1_REG_31__SCAN_IN), .ZN(n4479) );
  OAI211_X1 U5081 ( .C1(n4553), .C2(n4540), .A(n4480), .B(n4479), .ZN(U3549)
         );
  NAND2_X1 U5082 ( .A1(n4555), .A2(n4481), .ZN(n4483) );
  NAND2_X1 U5083 ( .A1(n3232), .A2(REG1_REG_30__SCAN_IN), .ZN(n4482) );
  OAI211_X1 U5084 ( .C1(n4558), .C2(n3232), .A(n4483), .B(n4482), .ZN(U3548)
         );
  NAND2_X1 U5085 ( .A1(n4484), .A2(n4545), .ZN(n4488) );
  INV_X1 U5086 ( .A(n4491), .ZN(n4485) );
  NAND3_X1 U5087 ( .A1(n4485), .A2(n4484), .A3(n4545), .ZN(n4487) );
  OAI211_X1 U5088 ( .C1(n4493), .C2(n4488), .A(n4487), .B(n4486), .ZN(n4489)
         );
  INV_X1 U5089 ( .A(n4489), .ZN(n4496) );
  NAND4_X1 U5090 ( .A1(n4493), .A2(n4545), .A3(n4492), .A4(n4491), .ZN(n4494)
         );
  MUX2_X1 U5091 ( .A(REG1_REG_27__SCAN_IN), .B(n4559), .S(n4725), .Z(U3545) );
  INV_X1 U5092 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4503) );
  MUX2_X1 U5093 ( .A(n4503), .B(n4502), .S(n4725), .Z(n4504) );
  OAI21_X1 U5094 ( .B1(n4540), .B2(n4505), .A(n4504), .ZN(U3544) );
  INV_X1 U5095 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4508) );
  AOI21_X1 U5096 ( .B1(n4507), .B2(n4545), .A(n4506), .ZN(n4560) );
  MUX2_X1 U5097 ( .A(n4508), .B(n4560), .S(n4725), .Z(n4509) );
  OAI21_X1 U5098 ( .B1(n4540), .B2(n4562), .A(n4509), .ZN(U3543) );
  INV_X1 U5099 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4512) );
  AOI21_X1 U5100 ( .B1(n4511), .B2(n4545), .A(n4510), .ZN(n4563) );
  MUX2_X1 U5101 ( .A(n4512), .B(n4563), .S(n4725), .Z(n4513) );
  OAI21_X1 U5102 ( .B1(n4540), .B2(n4566), .A(n4513), .ZN(U3542) );
  AOI21_X1 U5103 ( .B1(n4515), .B2(n4545), .A(n4514), .ZN(n4567) );
  MUX2_X1 U5104 ( .A(n4793), .B(n4567), .S(n4725), .Z(n4516) );
  OAI21_X1 U5105 ( .B1(n4540), .B2(n4570), .A(n4516), .ZN(U3541) );
  INV_X1 U5106 ( .A(n4311), .ZN(n4518) );
  NAND3_X1 U5107 ( .A1(n4518), .A2(n4698), .A3(n4517), .ZN(n4519) );
  OAI211_X1 U5108 ( .C1(n4521), .C2(n4710), .A(n4520), .B(n4519), .ZN(n4571)
         );
  MUX2_X1 U5109 ( .A(REG1_REG_22__SCAN_IN), .B(n4571), .S(n4725), .Z(U3540) );
  AOI21_X1 U5110 ( .B1(n4523), .B2(n4545), .A(n4522), .ZN(n4572) );
  MUX2_X1 U5111 ( .A(n4790), .B(n4572), .S(n4725), .Z(n4524) );
  OAI21_X1 U5112 ( .B1(n4540), .B2(n4575), .A(n4524), .ZN(U3539) );
  AOI21_X1 U5113 ( .B1(n4702), .B2(n4526), .A(n4525), .ZN(n4576) );
  MUX2_X1 U5114 ( .A(n4946), .B(n4576), .S(n4725), .Z(n4527) );
  OAI21_X1 U5115 ( .B1(n4540), .B2(n4579), .A(n4527), .ZN(U3538) );
  INV_X1 U5116 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4530) );
  AOI21_X1 U5117 ( .B1(n4529), .B2(n4545), .A(n4528), .ZN(n4580) );
  MUX2_X1 U5118 ( .A(n4530), .B(n4580), .S(n4725), .Z(n4531) );
  OAI21_X1 U5119 ( .B1(n4540), .B2(n4582), .A(n4531), .ZN(U3537) );
  INV_X1 U5120 ( .A(n4532), .ZN(n4535) );
  OAI211_X1 U5121 ( .C1(n4535), .C2(n4710), .A(n4534), .B(n4533), .ZN(n4583)
         );
  MUX2_X1 U5122 ( .A(REG1_REG_18__SCAN_IN), .B(n4583), .S(n4725), .Z(U3536) );
  AOI21_X1 U5123 ( .B1(n4537), .B2(n4545), .A(n4536), .ZN(n4584) );
  MUX2_X1 U5124 ( .A(n4538), .B(n4584), .S(n4725), .Z(n4539) );
  OAI21_X1 U5125 ( .B1(n4540), .B2(n4587), .A(n4539), .ZN(U3535) );
  NAND2_X1 U5126 ( .A1(n4541), .A2(n4698), .ZN(n4542) );
  OAI211_X1 U5127 ( .C1(n4710), .C2(n4544), .A(n4543), .B(n4542), .ZN(n4588)
         );
  MUX2_X1 U5128 ( .A(REG1_REG_16__SCAN_IN), .B(n4588), .S(n4725), .Z(U3534) );
  NAND2_X1 U5129 ( .A1(n4546), .A2(n4545), .ZN(n4547) );
  OAI211_X1 U5130 ( .C1(n4549), .C2(n4706), .A(n4548), .B(n4547), .ZN(n4589)
         );
  MUX2_X1 U5131 ( .A(REG1_REG_15__SCAN_IN), .B(n4589), .S(n4725), .Z(U3533) );
  NAND2_X1 U5132 ( .A1(n4717), .A2(n4550), .ZN(n4552) );
  NAND2_X1 U5133 ( .A1(n4716), .A2(REG0_REG_31__SCAN_IN), .ZN(n4551) );
  NAND2_X1 U5134 ( .A1(n4555), .A2(n4554), .ZN(n4557) );
  NAND2_X1 U5135 ( .A1(n4716), .A2(REG0_REG_30__SCAN_IN), .ZN(n4556) );
  OAI211_X1 U5136 ( .C1(n4558), .C2(n4716), .A(n4557), .B(n4556), .ZN(U3516)
         );
  MUX2_X1 U5137 ( .A(n4796), .B(n4560), .S(n4717), .Z(n4561) );
  OAI21_X1 U5138 ( .B1(n4562), .B2(n4586), .A(n4561), .ZN(U3511) );
  INV_X1 U5139 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4564) );
  MUX2_X1 U5140 ( .A(n4564), .B(n4563), .S(n4717), .Z(n4565) );
  OAI21_X1 U5141 ( .B1(n4566), .B2(n4586), .A(n4565), .ZN(U3510) );
  INV_X1 U5142 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4568) );
  MUX2_X1 U5143 ( .A(n4568), .B(n4567), .S(n4717), .Z(n4569) );
  OAI21_X1 U5144 ( .B1(n4570), .B2(n4586), .A(n4569), .ZN(U3509) );
  MUX2_X1 U5145 ( .A(REG0_REG_22__SCAN_IN), .B(n4571), .S(n4717), .Z(U3508) );
  INV_X1 U5146 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4573) );
  MUX2_X1 U5147 ( .A(n4573), .B(n4572), .S(n4717), .Z(n4574) );
  OAI21_X1 U5148 ( .B1(n4575), .B2(n4586), .A(n4574), .ZN(U3507) );
  INV_X1 U5149 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4577) );
  MUX2_X1 U5150 ( .A(n4577), .B(n4576), .S(n4717), .Z(n4578) );
  OAI21_X1 U5151 ( .B1(n4579), .B2(n4586), .A(n4578), .ZN(U3506) );
  MUX2_X1 U5152 ( .A(n4947), .B(n4580), .S(n4717), .Z(n4581) );
  OAI21_X1 U5153 ( .B1(n4582), .B2(n4586), .A(n4581), .ZN(U3505) );
  MUX2_X1 U5154 ( .A(REG0_REG_18__SCAN_IN), .B(n4583), .S(n4717), .Z(U3503) );
  INV_X1 U5155 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4949) );
  MUX2_X1 U5156 ( .A(n4949), .B(n4584), .S(n4717), .Z(n4585) );
  OAI21_X1 U5157 ( .B1(n4587), .B2(n4586), .A(n4585), .ZN(U3501) );
  MUX2_X1 U5158 ( .A(REG0_REG_16__SCAN_IN), .B(n4588), .S(n4717), .Z(U3499) );
  MUX2_X1 U5159 ( .A(REG0_REG_15__SCAN_IN), .B(n4589), .S(n4717), .Z(U3497) );
  MUX2_X1 U5160 ( .A(n4590), .B(DATAI_29_), .S(U3149), .Z(U3323) );
  MUX2_X1 U5161 ( .A(n4591), .B(DATAI_21_), .S(U3149), .Z(U3331) );
  MUX2_X1 U5162 ( .A(DATAI_20_), .B(n4592), .S(STATE_REG_SCAN_IN), .Z(U3332)
         );
  MUX2_X1 U5163 ( .A(n4593), .B(DATAI_19_), .S(U3149), .Z(U3333) );
  MUX2_X1 U5164 ( .A(n4594), .B(DATAI_14_), .S(U3149), .Z(U3338) );
  MUX2_X1 U5165 ( .A(DATAI_13_), .B(n4595), .S(STATE_REG_SCAN_IN), .Z(U3339)
         );
  MUX2_X1 U5166 ( .A(DATAI_12_), .B(n4596), .S(STATE_REG_SCAN_IN), .Z(U3340)
         );
  MUX2_X1 U5167 ( .A(n4597), .B(DATAI_10_), .S(U3149), .Z(U3342) );
  MUX2_X1 U5168 ( .A(n4598), .B(DATAI_9_), .S(U3149), .Z(U3343) );
  MUX2_X1 U5169 ( .A(DATAI_8_), .B(n4599), .S(STATE_REG_SCAN_IN), .Z(U3344) );
  MUX2_X1 U5170 ( .A(DATAI_7_), .B(n2631), .S(STATE_REG_SCAN_IN), .Z(U3345) );
  MUX2_X1 U5171 ( .A(n4601), .B(DATAI_6_), .S(U3149), .Z(U3346) );
  MUX2_X1 U5172 ( .A(DATAI_4_), .B(n4602), .S(STATE_REG_SCAN_IN), .Z(U3348) );
  MUX2_X1 U5173 ( .A(n4603), .B(DATAI_3_), .S(U3149), .Z(U3349) );
  MUX2_X1 U5174 ( .A(n2127), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  INV_X1 U5175 ( .A(DATAI_28_), .ZN(n4605) );
  AOI22_X1 U5176 ( .A1(STATE_REG_SCAN_IN), .A2(n4606), .B1(n4605), .B2(U3149), 
        .ZN(U3324) );
  OAI21_X1 U5177 ( .B1(REG1_REG_0__SCAN_IN), .B2(n4611), .A(n4607), .ZN(n4608)
         );
  MUX2_X1 U5178 ( .A(n4608), .B(n4607), .S(n4685), .Z(n4609) );
  OAI21_X1 U5179 ( .B1(n4611), .B2(n4610), .A(n4609), .ZN(n4613) );
  AOI22_X1 U5180 ( .A1(ADDR_REG_0__SCAN_IN), .A2(n4657), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n4612) );
  OAI21_X1 U5181 ( .B1(n4614), .B2(n4613), .A(n4612), .ZN(U3240) );
  INV_X1 U5182 ( .A(n4657), .ZN(n4627) );
  INV_X1 U5183 ( .A(ADDR_REG_15__SCAN_IN), .ZN(n4877) );
  AOI211_X1 U5184 ( .C1(n2147), .C2(n4617), .A(n4616), .B(n4615), .ZN(n4621)
         );
  AOI211_X1 U5185 ( .C1(n2159), .C2(n4619), .A(n4618), .B(n4653), .ZN(n4620)
         );
  AOI211_X1 U5186 ( .C1(n4623), .C2(n4622), .A(n4621), .B(n4620), .ZN(n4626)
         );
  INV_X1 U5187 ( .A(n4624), .ZN(n4625) );
  OAI211_X1 U5188 ( .C1(n4627), .C2(n4877), .A(n4626), .B(n4625), .ZN(U3255)
         );
  INV_X1 U5189 ( .A(n4628), .ZN(n4629) );
  AOI21_X1 U5190 ( .B1(n4657), .B2(ADDR_REG_16__SCAN_IN), .A(n4629), .ZN(n4639) );
  OAI21_X1 U5191 ( .B1(n4632), .B2(n4631), .A(n4630), .ZN(n4637) );
  OAI21_X1 U5192 ( .B1(n4635), .B2(n4634), .A(n4633), .ZN(n4636) );
  AOI22_X1 U5193 ( .A1(n4664), .A2(n4637), .B1(n4648), .B2(n4636), .ZN(n4638)
         );
  OAI211_X1 U5194 ( .C1(n4682), .C2(n4668), .A(n4639), .B(n4638), .ZN(U3256)
         );
  AOI21_X1 U5195 ( .B1(n4657), .B2(ADDR_REG_17__SCAN_IN), .A(n4640), .ZN(n4651) );
  OAI21_X1 U5196 ( .B1(n4643), .B2(n4642), .A(n4641), .ZN(n4649) );
  OAI21_X1 U5197 ( .B1(n4646), .B2(n4645), .A(n4644), .ZN(n4647) );
  AOI22_X1 U5198 ( .A1(n4664), .A2(n4649), .B1(n4648), .B2(n4647), .ZN(n4650)
         );
  OAI211_X1 U5199 ( .C1(n2532), .C2(n4668), .A(n4651), .B(n4650), .ZN(U3257)
         );
  INV_X1 U5200 ( .A(n4658), .ZN(n4659) );
  AOI21_X1 U5201 ( .B1(n4663), .B2(n4662), .A(n4661), .ZN(n4665) );
  NAND2_X1 U5202 ( .A1(n4665), .A2(n4664), .ZN(n4666) );
  OAI211_X1 U5203 ( .C1(n4668), .C2(n4679), .A(n4667), .B(n4666), .ZN(U3258)
         );
  AOI22_X1 U5204 ( .A1(REG3_REG_2__SCAN_IN), .A2(n4669), .B1(
        REG2_REG_2__SCAN_IN), .B2(n4459), .ZN(n4676) );
  INV_X1 U5205 ( .A(n4670), .ZN(n4671) );
  AOI22_X1 U5206 ( .A1(n4674), .A2(n4673), .B1(n4672), .B2(n4671), .ZN(n4675)
         );
  OAI211_X1 U5207 ( .C1(n4459), .C2(n4677), .A(n4676), .B(n4675), .ZN(U3288)
         );
  AND2_X1 U5208 ( .A1(D_REG_31__SCAN_IN), .A2(n4678), .ZN(U3291) );
  AND2_X1 U5209 ( .A1(D_REG_30__SCAN_IN), .A2(n4678), .ZN(U3292) );
  NOR2_X1 U5210 ( .A1(n4729), .A2(n4896), .ZN(U3293) );
  AND2_X1 U5211 ( .A1(D_REG_28__SCAN_IN), .A2(n4678), .ZN(U3294) );
  AND2_X1 U5212 ( .A1(D_REG_27__SCAN_IN), .A2(n4678), .ZN(U3295) );
  AND2_X1 U5213 ( .A1(D_REG_26__SCAN_IN), .A2(n4678), .ZN(U3296) );
  INV_X1 U5214 ( .A(D_REG_25__SCAN_IN), .ZN(n4943) );
  NOR2_X1 U5215 ( .A1(n4729), .A2(n4943), .ZN(U3297) );
  AND2_X1 U5216 ( .A1(D_REG_24__SCAN_IN), .A2(n4678), .ZN(U3298) );
  AND2_X1 U5217 ( .A1(D_REG_23__SCAN_IN), .A2(n4678), .ZN(U3299) );
  NOR2_X1 U5218 ( .A1(n4729), .A2(n4851), .ZN(U3300) );
  AND2_X1 U5219 ( .A1(D_REG_21__SCAN_IN), .A2(n4678), .ZN(U3301) );
  AND2_X1 U5220 ( .A1(D_REG_20__SCAN_IN), .A2(n4678), .ZN(U3302) );
  AND2_X1 U5221 ( .A1(D_REG_19__SCAN_IN), .A2(n4678), .ZN(U3303) );
  NOR2_X1 U5222 ( .A1(n4729), .A2(n4876), .ZN(U3304) );
  INV_X1 U5223 ( .A(D_REG_17__SCAN_IN), .ZN(n4940) );
  NOR2_X1 U5224 ( .A1(n4729), .A2(n4940), .ZN(U3305) );
  AND2_X1 U5225 ( .A1(D_REG_16__SCAN_IN), .A2(n4678), .ZN(U3306) );
  AND2_X1 U5226 ( .A1(D_REG_15__SCAN_IN), .A2(n4678), .ZN(U3307) );
  AND2_X1 U5227 ( .A1(D_REG_14__SCAN_IN), .A2(n4678), .ZN(U3308) );
  INV_X1 U5228 ( .A(D_REG_13__SCAN_IN), .ZN(n4899) );
  NOR2_X1 U5229 ( .A1(n4729), .A2(n4899), .ZN(U3309) );
  AND2_X1 U5230 ( .A1(D_REG_12__SCAN_IN), .A2(n4678), .ZN(U3310) );
  NOR2_X1 U5231 ( .A1(n4729), .A2(n4893), .ZN(U3311) );
  INV_X1 U5232 ( .A(D_REG_10__SCAN_IN), .ZN(n4941) );
  NOR2_X1 U5233 ( .A1(n4729), .A2(n4941), .ZN(U3312) );
  INV_X1 U5234 ( .A(D_REG_9__SCAN_IN), .ZN(n4944) );
  NOR2_X1 U5235 ( .A1(n4729), .A2(n4944), .ZN(U3313) );
  INV_X1 U5236 ( .A(D_REG_8__SCAN_IN), .ZN(n4818) );
  NOR2_X1 U5237 ( .A1(n4729), .A2(n4818), .ZN(U3314) );
  INV_X1 U5238 ( .A(D_REG_7__SCAN_IN), .ZN(n4819) );
  NOR2_X1 U5239 ( .A1(n4729), .A2(n4819), .ZN(U3315) );
  AND2_X1 U5240 ( .A1(D_REG_6__SCAN_IN), .A2(n4678), .ZN(U3316) );
  AND2_X1 U5241 ( .A1(D_REG_5__SCAN_IN), .A2(n4678), .ZN(U3317) );
  AND2_X1 U5242 ( .A1(D_REG_4__SCAN_IN), .A2(n4678), .ZN(U3318) );
  AND2_X1 U5243 ( .A1(D_REG_3__SCAN_IN), .A2(n4678), .ZN(U3319) );
  AND2_X1 U5244 ( .A1(D_REG_2__SCAN_IN), .A2(n4678), .ZN(U3320) );
  INV_X1 U5245 ( .A(DATAI_23_), .ZN(n4831) );
  AOI21_X1 U5246 ( .B1(U3149), .B2(n4831), .A(n4726), .ZN(U3329) );
  AOI22_X1 U5247 ( .A1(STATE_REG_SCAN_IN), .A2(n4679), .B1(n2747), .B2(U3149), 
        .ZN(U3334) );
  INV_X1 U5248 ( .A(DATAI_17_), .ZN(n4680) );
  AOI22_X1 U5249 ( .A1(STATE_REG_SCAN_IN), .A2(n2532), .B1(n4680), .B2(U3149), 
        .ZN(U3335) );
  AOI22_X1 U5250 ( .A1(STATE_REG_SCAN_IN), .A2(n4682), .B1(n4681), .B2(U3149), 
        .ZN(U3336) );
  INV_X1 U5251 ( .A(DATAI_15_), .ZN(n4683) );
  AOI22_X1 U5252 ( .A1(STATE_REG_SCAN_IN), .A2(n4684), .B1(n4683), .B2(U3149), 
        .ZN(U3337) );
  INV_X1 U5253 ( .A(DATAI_0_), .ZN(n4837) );
  AOI22_X1 U5254 ( .A1(STATE_REG_SCAN_IN), .A2(n4685), .B1(n4837), .B2(U3149), 
        .ZN(U3352) );
  INV_X1 U5255 ( .A(REG0_REG_0__SCAN_IN), .ZN(n4686) );
  AOI22_X1 U5256 ( .A1(n4717), .A2(n4687), .B1(n4686), .B2(n4716), .ZN(U3467)
         );
  INV_X1 U5257 ( .A(n4688), .ZN(n4692) );
  OAI22_X1 U5258 ( .A1(n4690), .A2(n4693), .B1(n4689), .B2(n4706), .ZN(n4691)
         );
  NOR2_X1 U5259 ( .A1(n4692), .A2(n4691), .ZN(n4718) );
  AOI22_X1 U5260 ( .A1(n4717), .A2(n4718), .B1(n2573), .B2(n4716), .ZN(U3469)
         );
  NOR2_X1 U5261 ( .A1(n4694), .A2(n4693), .ZN(n4696) );
  AOI211_X1 U5262 ( .C1(n4698), .C2(n4697), .A(n4696), .B(n4695), .ZN(n4720)
         );
  INV_X1 U5263 ( .A(REG0_REG_3__SCAN_IN), .ZN(n4927) );
  AOI22_X1 U5264 ( .A1(n4717), .A2(n4720), .B1(n4927), .B2(n4716), .ZN(U3473)
         );
  INV_X1 U5265 ( .A(n4699), .ZN(n4701) );
  AOI211_X1 U5266 ( .C1(n4703), .C2(n4702), .A(n4701), .B(n4700), .ZN(n4721)
         );
  INV_X1 U5267 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4704) );
  AOI22_X1 U5268 ( .A1(n4717), .A2(n4721), .B1(n4704), .B2(n4716), .ZN(U3475)
         );
  OAI22_X1 U5269 ( .A1(n4707), .A2(n4710), .B1(n4706), .B2(n4705), .ZN(n4708)
         );
  NOR2_X1 U5270 ( .A1(n4709), .A2(n4708), .ZN(n4722) );
  INV_X1 U5271 ( .A(REG0_REG_5__SCAN_IN), .ZN(n4919) );
  AOI22_X1 U5272 ( .A1(n4717), .A2(n4722), .B1(n4919), .B2(n4716), .ZN(U3477)
         );
  NOR3_X1 U5273 ( .A1(n4712), .A2(n4711), .A3(n4710), .ZN(n4715) );
  NOR3_X1 U5274 ( .A1(n4715), .A2(n4714), .A3(n4713), .ZN(n4724) );
  INV_X1 U5275 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4916) );
  AOI22_X1 U5276 ( .A1(n4717), .A2(n4724), .B1(n4916), .B2(n4716), .ZN(U3481)
         );
  AOI22_X1 U5277 ( .A1(n4725), .A2(n4718), .B1(n2500), .B2(n3232), .ZN(U3519)
         );
  INV_X1 U5278 ( .A(REG1_REG_3__SCAN_IN), .ZN(n4719) );
  AOI22_X1 U5279 ( .A1(n4725), .A2(n4720), .B1(n4719), .B2(n3232), .ZN(U3521)
         );
  AOI22_X1 U5280 ( .A1(n4725), .A2(n4721), .B1(n2273), .B2(n3232), .ZN(U3522)
         );
  AOI22_X1 U5281 ( .A1(n4725), .A2(n4722), .B1(n2512), .B2(n3232), .ZN(U3523)
         );
  AOI22_X1 U5282 ( .A1(n4725), .A2(n4724), .B1(n4723), .B2(n3232), .ZN(U3525)
         );
  INV_X1 U5283 ( .A(n4726), .ZN(n4728) );
  OAI22_X1 U5284 ( .A1(n4729), .A2(D_REG_1__SCAN_IN), .B1(n4728), .B2(n4727), 
        .ZN(n5036) );
  INV_X1 U5285 ( .A(DATAI_14_), .ZN(n4731) );
  NAND4_X1 U5286 ( .A1(n4731), .A2(n4730), .A3(REG3_REG_6__SCAN_IN), .A4(
        DATAI_0_), .ZN(n4732) );
  OR3_X1 U5287 ( .A1(n4732), .A2(REG3_REG_10__SCAN_IN), .A3(n4838), .ZN(n4745)
         );
  NAND4_X1 U5288 ( .A1(n4868), .A2(n4734), .A3(n4733), .A4(DATAI_27_), .ZN(
        n4735) );
  NOR3_X1 U5289 ( .A1(DATAO_REG_10__SCAN_IN), .A2(DATAO_REG_8__SCAN_IN), .A3(
        n4735), .ZN(n4743) );
  NAND4_X1 U5290 ( .A1(DATAO_REG_4__SCAN_IN), .A2(DATAI_23_), .A3(
        DATAO_REG_17__SCAN_IN), .A4(n4835), .ZN(n4741) );
  NAND4_X1 U5291 ( .A1(ADDR_REG_13__SCAN_IN), .A2(n2654), .A3(n4902), .A4(
        n4901), .ZN(n4736) );
  NOR2_X1 U5292 ( .A1(IR_REG_28__SCAN_IN), .A2(n4736), .ZN(n4738) );
  INV_X1 U5293 ( .A(DATAI_20_), .ZN(n4737) );
  NAND4_X1 U5294 ( .A1(n4738), .A2(DATAO_REG_2__SCAN_IN), .A3(n4737), .A4(
        DATAO_REG_15__SCAN_IN), .ZN(n4740) );
  NAND4_X1 U5295 ( .A1(ADDR_REG_15__SCAN_IN), .A2(DATAO_REG_27__SCAN_IN), .A3(
        DATAO_REG_6__SCAN_IN), .A4(DATAO_REG_18__SCAN_IN), .ZN(n4739) );
  NOR3_X1 U5296 ( .A1(n4741), .A2(n4740), .A3(n4739), .ZN(n4742) );
  NAND4_X1 U5297 ( .A1(REG3_REG_16__SCAN_IN), .A2(DATAI_4_), .A3(n4743), .A4(
        n4742), .ZN(n4744) );
  NOR4_X1 U5298 ( .A1(IR_REG_29__SCAN_IN), .A2(n4853), .A3(n4745), .A4(n4744), 
        .ZN(n4788) );
  NAND2_X1 U5299 ( .A1(IR_REG_10__SCAN_IN), .A2(IR_REG_31__SCAN_IN), .ZN(n4747) );
  NAND4_X1 U5300 ( .A1(STATE_REG_SCAN_IN), .A2(IR_REG_22__SCAN_IN), .A3(
        IR_REG_14__SCAN_IN), .A4(IR_REG_9__SCAN_IN), .ZN(n4746) );
  NOR4_X1 U5301 ( .A1(IR_REG_8__SCAN_IN), .A2(IR_REG_7__SCAN_IN), .A3(n4747), 
        .A4(n4746), .ZN(n4750) );
  INV_X1 U5302 ( .A(REG2_REG_18__SCAN_IN), .ZN(n4993) );
  NOR4_X1 U5303 ( .A1(REG3_REG_24__SCAN_IN), .A2(n4977), .A3(n2582), .A4(n4993), .ZN(n4749) );
  NOR4_X1 U5304 ( .A1(REG2_REG_17__SCAN_IN), .A2(ADDR_REG_19__SCAN_IN), .A3(
        n4988), .A4(n4976), .ZN(n4748) );
  AND4_X1 U5305 ( .A1(n4751), .A2(n4750), .A3(n4749), .A4(n4748), .ZN(n4786)
         );
  NAND4_X1 U5306 ( .A1(REG1_REG_13__SCAN_IN), .A2(REG1_REG_9__SCAN_IN), .A3(
        REG2_REG_0__SCAN_IN), .A4(n2441), .ZN(n4755) );
  NAND4_X1 U5307 ( .A1(REG3_REG_15__SCAN_IN), .A2(REG3_REG_13__SCAN_IN), .A3(
        ADDR_REG_16__SCAN_IN), .A4(ADDR_REG_12__SCAN_IN), .ZN(n4754) );
  NAND4_X1 U5308 ( .A1(REG0_REG_7__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .A3(
        REG0_REG_5__SCAN_IN), .A4(n4927), .ZN(n4753) );
  NAND4_X1 U5309 ( .A1(REG2_REG_14__SCAN_IN), .A2(REG2_REG_9__SCAN_IN), .A3(
        REG0_REG_1__SCAN_IN), .A4(n3618), .ZN(n4752) );
  NOR4_X1 U5310 ( .A1(n4755), .A2(n4754), .A3(n4753), .A4(n4752), .ZN(n4785)
         );
  NAND4_X1 U5311 ( .A1(REG0_REG_25__SCAN_IN), .A2(REG1_REG_23__SCAN_IN), .A3(
        REG2_REG_23__SCAN_IN), .A4(n4792), .ZN(n4760) );
  NAND4_X1 U5312 ( .A1(REG1_REG_20__SCAN_IN), .A2(REG0_REG_17__SCAN_IN), .A3(
        n4790), .A4(n4947), .ZN(n4759) );
  INV_X1 U5313 ( .A(REG0_REG_29__SCAN_IN), .ZN(n4756) );
  NAND4_X1 U5314 ( .A1(REG1_REG_29__SCAN_IN), .A2(REG0_REG_28__SCAN_IN), .A3(
        REG1_REG_28__SCAN_IN), .A4(n4756), .ZN(n4758) );
  INV_X1 U5315 ( .A(REG0_REG_27__SCAN_IN), .ZN(n4807) );
  NAND4_X1 U5316 ( .A1(REG1_REG_27__SCAN_IN), .A2(REG0_REG_26__SCAN_IN), .A3(
        REG2_REG_26__SCAN_IN), .A4(n4807), .ZN(n4757) );
  NOR4_X1 U5317 ( .A1(n4760), .A2(n4759), .A3(n4758), .A4(n4757), .ZN(n4784)
         );
  INV_X1 U5318 ( .A(n4761), .ZN(n4763) );
  INV_X1 U5319 ( .A(REG3_REG_1__SCAN_IN), .ZN(n4762) );
  AND4_X1 U5320 ( .A1(n4763), .A2(REG3_REG_2__SCAN_IN), .A3(D_REG_9__SCAN_IN), 
        .A4(n4762), .ZN(n4782) );
  INV_X1 U5321 ( .A(REG0_REG_16__SCAN_IN), .ZN(n4950) );
  NAND4_X1 U5322 ( .A1(D_REG_10__SCAN_IN), .A2(D_REG_25__SCAN_IN), .A3(
        D_REG_17__SCAN_IN), .A4(n4950), .ZN(n4766) );
  INV_X1 U5323 ( .A(DATAI_3_), .ZN(n4764) );
  NAND4_X1 U5324 ( .A1(n4764), .A2(DATAI_13_), .A3(REG3_REG_11__SCAN_IN), .A4(
        DATAI_9_), .ZN(n4765) );
  NOR2_X1 U5325 ( .A1(n4766), .A2(n4765), .ZN(n4781) );
  NAND2_X1 U5326 ( .A1(n4767), .A2(IR_REG_16__SCAN_IN), .ZN(n4777) );
  INV_X1 U5327 ( .A(ADDR_REG_0__SCAN_IN), .ZN(n5020) );
  NAND4_X1 U5328 ( .A1(REG1_REG_0__SCAN_IN), .A2(REG2_REG_6__SCAN_IN), .A3(
        ADDR_REG_1__SCAN_IN), .A4(n5020), .ZN(n4769) );
  INV_X1 U5329 ( .A(ADDR_REG_10__SCAN_IN), .ZN(n5002) );
  NAND4_X1 U5330 ( .A1(REG2_REG_10__SCAN_IN), .A2(REG2_REG_12__SCAN_IN), .A3(
        REG2_REG_8__SCAN_IN), .A4(n5002), .ZN(n4768) );
  NOR2_X1 U5331 ( .A1(n4769), .A2(n4768), .ZN(n4775) );
  INV_X1 U5332 ( .A(DATAI_21_), .ZN(n4973) );
  NAND4_X1 U5333 ( .A1(REG2_REG_27__SCAN_IN), .A2(REG2_REG_20__SCAN_IN), .A3(
        REG2_REG_24__SCAN_IN), .A4(n4973), .ZN(n4773) );
  INV_X1 U5334 ( .A(REG0_REG_9__SCAN_IN), .ZN(n4918) );
  NAND4_X1 U5335 ( .A1(REG3_REG_9__SCAN_IN), .A2(REG1_REG_8__SCAN_IN), .A3(
        REG0_REG_8__SCAN_IN), .A4(n4918), .ZN(n4772) );
  INV_X1 U5336 ( .A(REG0_REG_11__SCAN_IN), .ZN(n4957) );
  INV_X1 U5337 ( .A(REG0_REG_10__SCAN_IN), .ZN(n4912) );
  NAND4_X1 U5338 ( .A1(n4770), .A2(n4956), .A3(n4957), .A4(n4912), .ZN(n4771)
         );
  NOR3_X1 U5339 ( .A1(n4773), .A2(n4772), .A3(n4771), .ZN(n4774) );
  NAND3_X1 U5340 ( .A1(IR_REG_5__SCAN_IN), .A2(n4775), .A3(n4774), .ZN(n4776)
         );
  NOR2_X1 U5341 ( .A1(n4777), .A2(n4776), .ZN(n4780) );
  AND4_X1 U5342 ( .A1(n4778), .A2(n2469), .A3(IR_REG_26__SCAN_IN), .A4(
        DATAI_19_), .ZN(n4779) );
  AND4_X1 U5343 ( .A1(n4782), .A2(n4781), .A3(n4780), .A4(n4779), .ZN(n4783)
         );
  AND4_X1 U5344 ( .A1(n4786), .A2(n4785), .A3(n4784), .A4(n4783), .ZN(n4787)
         );
  AOI21_X1 U5345 ( .B1(n4788), .B2(n4787), .A(IR_REG_18__SCAN_IN), .ZN(n5034)
         );
  AOI22_X1 U5346 ( .A1(n4790), .A2(keyinput78), .B1(n4310), .B2(keyinput114), 
        .ZN(n4789) );
  OAI221_X1 U5347 ( .B1(n4790), .B2(keyinput78), .C1(n4310), .C2(keyinput114), 
        .A(n4789), .ZN(n4802) );
  AOI22_X1 U5348 ( .A1(n4793), .A2(keyinput11), .B1(n4792), .B2(keyinput33), 
        .ZN(n4791) );
  OAI221_X1 U5349 ( .B1(n4793), .B2(keyinput11), .C1(n4792), .C2(keyinput33), 
        .A(n4791), .ZN(n4801) );
  AOI22_X1 U5350 ( .A1(n4796), .A2(keyinput56), .B1(n4795), .B2(keyinput20), 
        .ZN(n4794) );
  OAI221_X1 U5351 ( .B1(n4796), .B2(keyinput56), .C1(n4795), .C2(keyinput20), 
        .A(n4794), .ZN(n4800) );
  AOI22_X1 U5352 ( .A1(n4252), .A2(keyinput21), .B1(n4798), .B2(keyinput30), 
        .ZN(n4797) );
  OAI221_X1 U5353 ( .B1(n4252), .B2(keyinput21), .C1(n4798), .C2(keyinput30), 
        .A(n4797), .ZN(n4799) );
  NOR4_X1 U5354 ( .A1(n4802), .A2(n4801), .A3(n4800), .A4(n4799), .ZN(n4849)
         );
  AOI22_X1 U5355 ( .A1(n2556), .A2(keyinput67), .B1(keyinput47), .B2(n4804), 
        .ZN(n4803) );
  OAI221_X1 U5356 ( .B1(n2556), .B2(keyinput67), .C1(n4804), .C2(keyinput47), 
        .A(n4803), .ZN(n4816) );
  AOI22_X1 U5357 ( .A1(n4807), .A2(keyinput70), .B1(n4806), .B2(keyinput18), 
        .ZN(n4805) );
  OAI221_X1 U5358 ( .B1(n4807), .B2(keyinput70), .C1(n4806), .C2(keyinput18), 
        .A(n4805), .ZN(n4815) );
  AOI22_X1 U5359 ( .A1(n4810), .A2(keyinput103), .B1(n4809), .B2(keyinput25), 
        .ZN(n4808) );
  OAI221_X1 U5360 ( .B1(n4810), .B2(keyinput103), .C1(n4809), .C2(keyinput25), 
        .A(n4808), .ZN(n4814) );
  XNOR2_X1 U5361 ( .A(REG0_REG_29__SCAN_IN), .B(keyinput83), .ZN(n4812) );
  XNOR2_X1 U5362 ( .A(IR_REG_28__SCAN_IN), .B(keyinput69), .ZN(n4811) );
  NAND2_X1 U5363 ( .A1(n4812), .A2(n4811), .ZN(n4813) );
  NOR4_X1 U5364 ( .A1(n4816), .A2(n4815), .A3(n4814), .A4(n4813), .ZN(n4848)
         );
  AOI22_X1 U5365 ( .A1(n4819), .A2(keyinput15), .B1(keyinput87), .B2(n4818), 
        .ZN(n4817) );
  OAI221_X1 U5366 ( .B1(n4819), .B2(keyinput15), .C1(n4818), .C2(keyinput87), 
        .A(n4817), .ZN(n4829) );
  XNOR2_X1 U5367 ( .A(n4820), .B(keyinput99), .ZN(n4828) );
  XNOR2_X1 U5368 ( .A(keyinput3), .B(n4821), .ZN(n4827) );
  XNOR2_X1 U5369 ( .A(IR_REG_14__SCAN_IN), .B(keyinput43), .ZN(n4825) );
  XNOR2_X1 U5370 ( .A(DATAI_20_), .B(keyinput27), .ZN(n4824) );
  XNOR2_X1 U5371 ( .A(IR_REG_8__SCAN_IN), .B(keyinput63), .ZN(n4823) );
  XNOR2_X1 U5372 ( .A(IR_REG_5__SCAN_IN), .B(keyinput127), .ZN(n4822) );
  NAND4_X1 U5373 ( .A1(n4825), .A2(n4824), .A3(n4823), .A4(n4822), .ZN(n4826)
         );
  NOR4_X1 U5374 ( .A1(n4829), .A2(n4828), .A3(n4827), .A4(n4826), .ZN(n4847)
         );
  AOI22_X1 U5375 ( .A1(n4832), .A2(keyinput111), .B1(n4831), .B2(keyinput119), 
        .ZN(n4830) );
  OAI221_X1 U5376 ( .B1(n4832), .B2(keyinput111), .C1(n4831), .C2(keyinput119), 
        .A(n4830), .ZN(n4845) );
  AOI22_X1 U5377 ( .A1(n4835), .A2(keyinput107), .B1(n4834), .B2(keyinput115), 
        .ZN(n4833) );
  OAI221_X1 U5378 ( .B1(n4835), .B2(keyinput107), .C1(n4834), .C2(keyinput115), 
        .A(n4833), .ZN(n4844) );
  AOI22_X1 U5379 ( .A1(n4838), .A2(keyinput51), .B1(keyinput75), .B2(n4837), 
        .ZN(n4836) );
  OAI221_X1 U5380 ( .B1(n4838), .B2(keyinput51), .C1(n4837), .C2(keyinput75), 
        .A(n4836), .ZN(n4843) );
  INV_X1 U5381 ( .A(IR_REG_29__SCAN_IN), .ZN(n4841) );
  INV_X1 U5382 ( .A(IR_REG_23__SCAN_IN), .ZN(n4840) );
  AOI22_X1 U5383 ( .A1(n4841), .A2(keyinput28), .B1(n4840), .B2(keyinput24), 
        .ZN(n4839) );
  OAI221_X1 U5384 ( .B1(n4841), .B2(keyinput28), .C1(n4840), .C2(keyinput24), 
        .A(n4839), .ZN(n4842) );
  NOR4_X1 U5385 ( .A1(n4845), .A2(n4844), .A3(n4843), .A4(n4842), .ZN(n4846)
         );
  NAND4_X1 U5386 ( .A1(n4849), .A2(n4848), .A3(n4847), .A4(n4846), .ZN(n5032)
         );
  AOI22_X1 U5387 ( .A1(n2859), .A2(keyinput40), .B1(keyinput32), .B2(n4851), 
        .ZN(n4850) );
  OAI221_X1 U5388 ( .B1(n2859), .B2(keyinput40), .C1(n4851), .C2(keyinput32), 
        .A(n4850), .ZN(n4860) );
  AOI22_X1 U5389 ( .A1(n4853), .A2(keyinput36), .B1(n4731), .B2(keyinput41), 
        .ZN(n4852) );
  OAI221_X1 U5390 ( .B1(n4853), .B2(keyinput36), .C1(n4731), .C2(keyinput41), 
        .A(n4852), .ZN(n4859) );
  XNOR2_X1 U5391 ( .A(REG3_REG_10__SCAN_IN), .B(keyinput6), .ZN(n4857) );
  XNOR2_X1 U5392 ( .A(REG3_REG_8__SCAN_IN), .B(keyinput4), .ZN(n4856) );
  XNOR2_X1 U5393 ( .A(REG3_REG_6__SCAN_IN), .B(keyinput9), .ZN(n4855) );
  XNOR2_X1 U5394 ( .A(REG3_REG_19__SCAN_IN), .B(keyinput0), .ZN(n4854) );
  NAND4_X1 U5395 ( .A1(n4857), .A2(n4856), .A3(n4855), .A4(n4854), .ZN(n4858)
         );
  NOR3_X1 U5396 ( .A1(n4860), .A2(n4859), .A3(n4858), .ZN(n4910) );
  INV_X1 U5397 ( .A(IR_REG_9__SCAN_IN), .ZN(n4863) );
  AOI22_X1 U5398 ( .A1(n4863), .A2(keyinput120), .B1(keyinput117), .B2(n4862), 
        .ZN(n4861) );
  OAI221_X1 U5399 ( .B1(n4863), .B2(keyinput120), .C1(n4862), .C2(keyinput117), 
        .A(n4861), .ZN(n4874) );
  AOI22_X1 U5400 ( .A1(n4865), .A2(keyinput122), .B1(n2453), .B2(keyinput125), 
        .ZN(n4864) );
  OAI221_X1 U5401 ( .B1(n4865), .B2(keyinput122), .C1(n2453), .C2(keyinput125), 
        .A(n4864), .ZN(n4873) );
  AOI22_X1 U5402 ( .A1(n4868), .A2(keyinput17), .B1(keyinput10), .B2(n4867), 
        .ZN(n4866) );
  OAI221_X1 U5403 ( .B1(n4868), .B2(keyinput17), .C1(n4867), .C2(keyinput10), 
        .A(n4866), .ZN(n4872) );
  XNOR2_X1 U5404 ( .A(IR_REG_12__SCAN_IN), .B(keyinput126), .ZN(n4870) );
  XNOR2_X1 U5405 ( .A(DATAI_4_), .B(keyinput12), .ZN(n4869) );
  NAND2_X1 U5406 ( .A1(n4870), .A2(n4869), .ZN(n4871) );
  NOR4_X1 U5407 ( .A1(n4874), .A2(n4873), .A3(n4872), .A4(n4871), .ZN(n4909)
         );
  AOI22_X1 U5408 ( .A1(n4877), .A2(keyinput97), .B1(n4876), .B2(keyinput72), 
        .ZN(n4875) );
  OAI221_X1 U5409 ( .B1(n4877), .B2(keyinput97), .C1(n4876), .C2(keyinput72), 
        .A(n4875), .ZN(n4878) );
  INV_X1 U5410 ( .A(n4878), .ZN(n4891) );
  INV_X1 U5411 ( .A(keyinput100), .ZN(n4879) );
  XNOR2_X1 U5412 ( .A(n4880), .B(n4879), .ZN(n4890) );
  XNOR2_X1 U5413 ( .A(n4881), .B(keyinput64), .ZN(n4884) );
  XNOR2_X1 U5414 ( .A(n4882), .B(keyinput106), .ZN(n4883) );
  NOR2_X1 U5415 ( .A1(n4884), .A2(n4883), .ZN(n4889) );
  XNOR2_X1 U5416 ( .A(IR_REG_10__SCAN_IN), .B(keyinput65), .ZN(n4887) );
  XNOR2_X1 U5417 ( .A(IR_REG_25__SCAN_IN), .B(keyinput104), .ZN(n4886) );
  XNOR2_X1 U5418 ( .A(DATAI_7_), .B(keyinput105), .ZN(n4885) );
  AND3_X1 U5419 ( .A1(n4887), .A2(n4886), .A3(n4885), .ZN(n4888) );
  AND4_X1 U5420 ( .A1(n4891), .A2(n4890), .A3(n4889), .A4(n4888), .ZN(n4908)
         );
  AOI22_X1 U5421 ( .A1(n4894), .A2(keyinput62), .B1(n4893), .B2(keyinput57), 
        .ZN(n4892) );
  OAI221_X1 U5422 ( .B1(n4894), .B2(keyinput62), .C1(n4893), .C2(keyinput57), 
        .A(n4892), .ZN(n4906) );
  AOI22_X1 U5423 ( .A1(n2654), .A2(keyinput54), .B1(n4896), .B2(keyinput50), 
        .ZN(n4895) );
  OAI221_X1 U5424 ( .B1(n2654), .B2(keyinput54), .C1(n4896), .C2(keyinput50), 
        .A(n4895), .ZN(n4905) );
  INV_X1 U5425 ( .A(ADDR_REG_13__SCAN_IN), .ZN(n4898) );
  AOI22_X1 U5426 ( .A1(n4899), .A2(keyinput53), .B1(keyinput46), .B2(n4898), 
        .ZN(n4897) );
  OAI221_X1 U5427 ( .B1(n4899), .B2(keyinput53), .C1(n4898), .C2(keyinput46), 
        .A(n4897), .ZN(n4904) );
  AOI22_X1 U5428 ( .A1(n4902), .A2(keyinput42), .B1(keyinput45), .B2(n4901), 
        .ZN(n4900) );
  OAI221_X1 U5429 ( .B1(n4902), .B2(keyinput42), .C1(n4901), .C2(keyinput45), 
        .A(n4900), .ZN(n4903) );
  NOR4_X1 U5430 ( .A1(n4906), .A2(n4905), .A3(n4904), .A4(n4903), .ZN(n4907)
         );
  NAND4_X1 U5431 ( .A1(n4910), .A2(n4909), .A3(n4908), .A4(n4907), .ZN(n5031)
         );
  AOI22_X1 U5432 ( .A1(n4913), .A2(keyinput52), .B1(keyinput118), .B2(n4912), 
        .ZN(n4911) );
  OAI221_X1 U5433 ( .B1(n4913), .B2(keyinput52), .C1(n4912), .C2(keyinput118), 
        .A(n4911), .ZN(n4925) );
  INV_X1 U5434 ( .A(REG0_REG_8__SCAN_IN), .ZN(n4915) );
  AOI22_X1 U5435 ( .A1(n4916), .A2(keyinput19), .B1(n4915), .B2(keyinput77), 
        .ZN(n4914) );
  OAI221_X1 U5436 ( .B1(n4916), .B2(keyinput19), .C1(n4915), .C2(keyinput77), 
        .A(n4914), .ZN(n4924) );
  AOI22_X1 U5437 ( .A1(n2210), .A2(keyinput93), .B1(n4918), .B2(keyinput60), 
        .ZN(n4917) );
  OAI221_X1 U5438 ( .B1(n2210), .B2(keyinput93), .C1(n4918), .C2(keyinput60), 
        .A(n4917), .ZN(n4923) );
  XOR2_X1 U5439 ( .A(n4919), .B(keyinput121), .Z(n4921) );
  XNOR2_X1 U5440 ( .A(REG3_REG_4__SCAN_IN), .B(keyinput80), .ZN(n4920) );
  NAND2_X1 U5441 ( .A1(n4921), .A2(n4920), .ZN(n4922) );
  NOR4_X1 U5442 ( .A1(n4925), .A2(n4924), .A3(n4923), .A4(n4922), .ZN(n4970)
         );
  AOI22_X1 U5443 ( .A1(n2573), .A2(keyinput59), .B1(n4927), .B2(keyinput7), 
        .ZN(n4926) );
  OAI221_X1 U5444 ( .B1(n2573), .B2(keyinput59), .C1(n4927), .C2(keyinput7), 
        .A(n4926), .ZN(n4938) );
  INV_X1 U5445 ( .A(REG2_REG_0__SCAN_IN), .ZN(n4929) );
  AOI22_X1 U5446 ( .A1(n2441), .A2(keyinput94), .B1(keyinput37), .B2(n4929), 
        .ZN(n4928) );
  OAI221_X1 U5447 ( .B1(n2441), .B2(keyinput94), .C1(n4929), .C2(keyinput37), 
        .A(n4928), .ZN(n4937) );
  AOI22_X1 U5448 ( .A1(n4931), .A2(keyinput13), .B1(n3618), .B2(keyinput81), 
        .ZN(n4930) );
  OAI221_X1 U5449 ( .B1(n4931), .B2(keyinput13), .C1(n3618), .C2(keyinput81), 
        .A(n4930), .ZN(n4936) );
  XOR2_X1 U5450 ( .A(n4932), .B(keyinput85), .Z(n4934) );
  XNOR2_X1 U5451 ( .A(IR_REG_31__SCAN_IN), .B(keyinput2), .ZN(n4933) );
  NAND2_X1 U5452 ( .A1(n4934), .A2(n4933), .ZN(n4935) );
  NOR4_X1 U5453 ( .A1(n4938), .A2(n4937), .A3(n4936), .A4(n4935), .ZN(n4969)
         );
  AOI22_X1 U5454 ( .A1(n4941), .A2(keyinput26), .B1(keyinput16), .B2(n4940), 
        .ZN(n4939) );
  OAI221_X1 U5455 ( .B1(n4941), .B2(keyinput26), .C1(n4940), .C2(keyinput16), 
        .A(n4939), .ZN(n4954) );
  AOI22_X1 U5456 ( .A1(n4944), .A2(keyinput76), .B1(keyinput116), .B2(n4943), 
        .ZN(n4942) );
  OAI221_X1 U5457 ( .B1(n4944), .B2(keyinput76), .C1(n4943), .C2(keyinput116), 
        .A(n4942), .ZN(n4953) );
  AOI22_X1 U5458 ( .A1(n4947), .A2(keyinput22), .B1(n4946), .B2(keyinput95), 
        .ZN(n4945) );
  OAI221_X1 U5459 ( .B1(n4947), .B2(keyinput22), .C1(n4946), .C2(keyinput95), 
        .A(n4945), .ZN(n4952) );
  AOI22_X1 U5460 ( .A1(n4950), .A2(keyinput88), .B1(n4949), .B2(keyinput29), 
        .ZN(n4948) );
  OAI221_X1 U5461 ( .B1(n4950), .B2(keyinput88), .C1(n4949), .C2(keyinput29), 
        .A(n4948), .ZN(n4951) );
  NOR4_X1 U5462 ( .A1(n4954), .A2(n4953), .A3(n4952), .A4(n4951), .ZN(n4968)
         );
  AOI22_X1 U5463 ( .A1(n4957), .A2(keyinput68), .B1(n4956), .B2(keyinput108), 
        .ZN(n4955) );
  OAI221_X1 U5464 ( .B1(n4957), .B2(keyinput68), .C1(n4956), .C2(keyinput108), 
        .A(n4955), .ZN(n4966) );
  XNOR2_X1 U5465 ( .A(REG1_REG_14__SCAN_IN), .B(keyinput124), .ZN(n4961) );
  XNOR2_X1 U5466 ( .A(DATAI_3_), .B(keyinput5), .ZN(n4960) );
  XNOR2_X1 U5467 ( .A(DATAI_9_), .B(keyinput109), .ZN(n4959) );
  XNOR2_X1 U5468 ( .A(IR_REG_11__SCAN_IN), .B(keyinput112), .ZN(n4958) );
  NAND4_X1 U5469 ( .A1(n4961), .A2(n4960), .A3(n4959), .A4(n4958), .ZN(n4965)
         );
  XNOR2_X1 U5470 ( .A(n4962), .B(keyinput61), .ZN(n4964) );
  XNOR2_X1 U5471 ( .A(keyinput90), .B(n2699), .ZN(n4963) );
  NOR4_X1 U5472 ( .A1(n4966), .A2(n4965), .A3(n4964), .A4(n4963), .ZN(n4967)
         );
  NAND4_X1 U5473 ( .A1(n4970), .A2(n4969), .A3(n4968), .A4(n4967), .ZN(n5030)
         );
  AOI22_X1 U5474 ( .A1(n4245), .A2(keyinput86), .B1(keyinput92), .B2(n2795), 
        .ZN(n4971) );
  OAI221_X1 U5475 ( .B1(n4245), .B2(keyinput86), .C1(n2795), .C2(keyinput92), 
        .A(n4971), .ZN(n4983) );
  INV_X1 U5476 ( .A(REG2_REG_20__SCAN_IN), .ZN(n4974) );
  AOI22_X1 U5477 ( .A1(n4974), .A2(keyinput110), .B1(n4973), .B2(keyinput55), 
        .ZN(n4972) );
  OAI221_X1 U5478 ( .B1(n4974), .B2(keyinput110), .C1(n4973), .C2(keyinput55), 
        .A(n4972), .ZN(n4982) );
  AOI22_X1 U5479 ( .A1(n4977), .A2(keyinput31), .B1(n4976), .B2(keyinput82), 
        .ZN(n4975) );
  OAI221_X1 U5480 ( .B1(n4977), .B2(keyinput31), .C1(n4976), .C2(keyinput82), 
        .A(n4975), .ZN(n4981) );
  XNOR2_X1 U5481 ( .A(REG3_REG_1__SCAN_IN), .B(keyinput96), .ZN(n4979) );
  XNOR2_X1 U5482 ( .A(DATAI_19_), .B(keyinput71), .ZN(n4978) );
  NAND2_X1 U5483 ( .A1(n4979), .A2(n4978), .ZN(n4980) );
  NOR4_X1 U5484 ( .A1(n4983), .A2(n4982), .A3(n4981), .A4(n4980), .ZN(n5028)
         );
  INV_X1 U5485 ( .A(keyinput39), .ZN(n4986) );
  INV_X1 U5486 ( .A(ADDR_REG_19__SCAN_IN), .ZN(n4984) );
  XOR2_X1 U5487 ( .A(n4984), .B(keyinput74), .Z(n4985) );
  OAI21_X1 U5488 ( .B1(IR_REG_18__SCAN_IN), .B2(n4986), .A(n4985), .ZN(n4997)
         );
  AOI22_X1 U5489 ( .A1(n4989), .A2(keyinput84), .B1(n4988), .B2(keyinput123), 
        .ZN(n4987) );
  OAI221_X1 U5490 ( .B1(n4989), .B2(keyinput84), .C1(n4988), .C2(keyinput123), 
        .A(n4987), .ZN(n4996) );
  AOI22_X1 U5491 ( .A1(n2582), .A2(keyinput101), .B1(n4991), .B2(keyinput102), 
        .ZN(n4990) );
  OAI221_X1 U5492 ( .B1(n2582), .B2(keyinput101), .C1(n4991), .C2(keyinput102), 
        .A(n4990), .ZN(n4995) );
  AOI22_X1 U5493 ( .A1(n4993), .A2(keyinput49), .B1(U3149), .B2(keyinput73), 
        .ZN(n4992) );
  OAI221_X1 U5494 ( .B1(n4993), .B2(keyinput49), .C1(U3149), .C2(keyinput73), 
        .A(n4992), .ZN(n4994) );
  NOR4_X1 U5495 ( .A1(n4997), .A2(n4996), .A3(n4995), .A4(n4994), .ZN(n5027)
         );
  INV_X1 U5496 ( .A(ADDR_REG_12__SCAN_IN), .ZN(n5000) );
  AOI22_X1 U5497 ( .A1(n5000), .A2(keyinput44), .B1(n4999), .B2(keyinput98), 
        .ZN(n4998) );
  OAI221_X1 U5498 ( .B1(n5000), .B2(keyinput44), .C1(n4999), .C2(keyinput98), 
        .A(n4998), .ZN(n5012) );
  AOI22_X1 U5499 ( .A1(n5002), .A2(keyinput48), .B1(n3658), .B2(keyinput113), 
        .ZN(n5001) );
  OAI221_X1 U5500 ( .B1(n5002), .B2(keyinput48), .C1(n3658), .C2(keyinput113), 
        .A(n5001), .ZN(n5011) );
  AOI22_X1 U5501 ( .A1(n5005), .A2(keyinput1), .B1(keyinput34), .B2(n5004), 
        .ZN(n5003) );
  OAI221_X1 U5502 ( .B1(n5005), .B2(keyinput1), .C1(n5004), .C2(keyinput34), 
        .A(n5003), .ZN(n5010) );
  INV_X1 U5503 ( .A(ADDR_REG_16__SCAN_IN), .ZN(n5007) );
  AOI22_X1 U5504 ( .A1(n5008), .A2(keyinput66), .B1(keyinput91), .B2(n5007), 
        .ZN(n5006) );
  OAI221_X1 U5505 ( .B1(n5008), .B2(keyinput66), .C1(n5007), .C2(keyinput91), 
        .A(n5006), .ZN(n5009) );
  NOR4_X1 U5506 ( .A1(n5012), .A2(n5011), .A3(n5010), .A4(n5009), .ZN(n5026)
         );
  INV_X1 U5507 ( .A(ADDR_REG_1__SCAN_IN), .ZN(n5015) );
  INV_X1 U5508 ( .A(REG2_REG_6__SCAN_IN), .ZN(n5014) );
  AOI22_X1 U5509 ( .A1(n5015), .A2(keyinput8), .B1(n5014), .B2(keyinput38), 
        .ZN(n5013) );
  OAI221_X1 U5510 ( .B1(n5015), .B2(keyinput8), .C1(n5014), .C2(keyinput38), 
        .A(n5013), .ZN(n5024) );
  AOI22_X1 U5511 ( .A1(n2344), .A2(keyinput58), .B1(n3526), .B2(keyinput89), 
        .ZN(n5016) );
  OAI221_X1 U5512 ( .B1(n2344), .B2(keyinput58), .C1(n3526), .C2(keyinput89), 
        .A(n5016), .ZN(n5023) );
  XNOR2_X1 U5513 ( .A(REG3_REG_11__SCAN_IN), .B(keyinput35), .ZN(n5019) );
  XNOR2_X1 U5514 ( .A(REG1_REG_0__SCAN_IN), .B(keyinput79), .ZN(n5018) );
  XNOR2_X1 U5515 ( .A(REG3_REG_2__SCAN_IN), .B(keyinput14), .ZN(n5017) );
  NAND3_X1 U5516 ( .A1(n5019), .A2(n5018), .A3(n5017), .ZN(n5022) );
  XNOR2_X1 U5517 ( .A(n5020), .B(keyinput23), .ZN(n5021) );
  NOR4_X1 U5518 ( .A1(n5024), .A2(n5023), .A3(n5022), .A4(n5021), .ZN(n5025)
         );
  NAND4_X1 U5519 ( .A1(n5028), .A2(n5027), .A3(n5026), .A4(n5025), .ZN(n5029)
         );
  NOR4_X1 U5520 ( .A1(n5032), .A2(n5031), .A3(n5030), .A4(n5029), .ZN(n5033)
         );
  OAI21_X1 U5521 ( .B1(keyinput39), .B2(n5034), .A(n5033), .ZN(n5035) );
  XOR2_X1 U5522 ( .A(n5036), .B(n5035), .Z(U3459) );
  CLKBUF_X1 U2367 ( .A(n2898), .Z(n3104) );
  INV_X1 U2373 ( .A(n2906), .ZN(n2923) );
  CLKBUF_X1 U2451 ( .A(n2621), .Z(n3964) );
  CLKBUF_X1 U2469 ( .A(n2612), .Z(n3968) );
endmodule

