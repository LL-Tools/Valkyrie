

module b21_C_AntiSAT_k_128_1 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3, 
        keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, 
        keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, 
        keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, 
        keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, 
        keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, 
        keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, 
        keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, 
        keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, 
        keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, 
        keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, 
        keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, 
        keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, 
        keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, 
        keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, 
        keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, 
        keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, 
        keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, 
        keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, 
        keyinput110, keyinput111, keyinput112, keyinput113, keyinput114, 
        keyinput115, keyinput116, keyinput117, keyinput118, keyinput119, 
        keyinput120, keyinput121, keyinput122, keyinput123, keyinput124, 
        keyinput125, keyinput126, keyinput127, ADD_1071_U4, ADD_1071_U55, 
        ADD_1071_U56, ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, 
        ADD_1071_U61, ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, 
        ADD_1071_U49, ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, 
        ADD_1071_U54, ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, 
        P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, 
        P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, 
        P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, 
        P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, 
        P1_U3324, P1_U3323, P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, 
        P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, 
        P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, 
        P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, 
        P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, 
        P1_U3454, P1_U3457, P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, 
        P1_U3475, P1_U3478, P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, 
        P1_U3496, P1_U3499, P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, 
        P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, 
        P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, 
        P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, 
        P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, 
        P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, 
        P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, 
        P1_U3554, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, 
        P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, 
        P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, 
        P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, 
        P1_U3264, P1_U3263, P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, 
        P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, 
        P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, 
        P1_U3244, P1_U3243, P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, 
        P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, 
        P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, 
        P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, 
        P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, 
        P1_U3586, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, 
        P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, 
        P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, 
        P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, 
        P1_U3213, P1_U3212, P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, 
        P2_U3357, P2_U3356, P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, 
        P2_U3350, P2_U3349, P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, 
        P2_U3343, P2_U3342, P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, 
        P2_U3336, P2_U3335, P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, 
        P2_U3329, P2_U3328, P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, 
        P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, 
        P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, 
        P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, 
        P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, 
        P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, 
        P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, 
        P2_U3493, P2_U3496, P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, 
        P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, 
        P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, 
        P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, 
        P2_U3530, P2_U3531, P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, 
        P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, 
        P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, 
        P2_U3551, P2_U3296, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, 
        P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, 
        P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, 
        P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, 
        P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, 
        P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, 
        P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, 
        P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, 
        P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, 
        P2_U3562, P2_U3563, P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, 
        P2_U3569, P2_U3570, P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, 
        P2_U3576, P2_U3577, P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, 
        P2_U3583, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, 
        P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, 
        P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, 
        P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, 
        P2_U3217, P2_U3216, P2_U3215, P2_U3152, P2_U3151, P2_U3966 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298,
         n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308,
         n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318,
         n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328,
         n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338,
         n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348,
         n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
         n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368,
         n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378,
         n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
         n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
         n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
         n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
         n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
         n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
         n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
         n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
         n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
         n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
         n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
         n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
         n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
         n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
         n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
         n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
         n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
         n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
         n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
         n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
         n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
         n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
         n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
         n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
         n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
         n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
         n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
         n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
         n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
         n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
         n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
         n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
         n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718,
         n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728,
         n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738,
         n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748,
         n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758,
         n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768,
         n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778,
         n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788,
         n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798,
         n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808,
         n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818,
         n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828,
         n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838,
         n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848,
         n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858,
         n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868,
         n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878,
         n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888,
         n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898,
         n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908,
         n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918,
         n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928,
         n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938,
         n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948,
         n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958,
         n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968,
         n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978,
         n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988,
         n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998,
         n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008,
         n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018,
         n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028,
         n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038,
         n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048,
         n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058,
         n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068,
         n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078,
         n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088,
         n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098,
         n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108,
         n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118,
         n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128,
         n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138,
         n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148,
         n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158,
         n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168,
         n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178,
         n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188,
         n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198,
         n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208,
         n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218,
         n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228,
         n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238,
         n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248,
         n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258,
         n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268,
         n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278,
         n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288,
         n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298,
         n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308,
         n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318,
         n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328,
         n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338,
         n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348,
         n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358,
         n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368,
         n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378,
         n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388,
         n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398,
         n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408,
         n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418,
         n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428,
         n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438,
         n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448,
         n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458,
         n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468,
         n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478,
         n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488,
         n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498,
         n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508,
         n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518,
         n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528,
         n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538,
         n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548,
         n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558,
         n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568,
         n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578,
         n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588,
         n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598,
         n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608,
         n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618,
         n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628,
         n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638,
         n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648,
         n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658,
         n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668,
         n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678,
         n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688,
         n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698,
         n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708,
         n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718,
         n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728,
         n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738,
         n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748,
         n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758,
         n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768,
         n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778,
         n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788,
         n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798,
         n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808,
         n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818,
         n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828,
         n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838,
         n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848,
         n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858,
         n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868,
         n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878,
         n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888,
         n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898,
         n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908,
         n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918,
         n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928,
         n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938,
         n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948,
         n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958,
         n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968,
         n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978,
         n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988,
         n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998,
         n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008,
         n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018,
         n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028,
         n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038,
         n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048,
         n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058,
         n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068,
         n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078,
         n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088,
         n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098,
         n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108,
         n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118,
         n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128,
         n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138,
         n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148,
         n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158,
         n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168,
         n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178,
         n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188,
         n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198,
         n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208,
         n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218,
         n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228,
         n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238,
         n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248,
         n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258,
         n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268,
         n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278,
         n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288,
         n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298,
         n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308,
         n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318,
         n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328,
         n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338,
         n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348,
         n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358,
         n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368,
         n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378,
         n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388,
         n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398,
         n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408,
         n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418,
         n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428,
         n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438,
         n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448,
         n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458,
         n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468,
         n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478,
         n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488,
         n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498,
         n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508,
         n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518,
         n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528,
         n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538,
         n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548,
         n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558,
         n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568,
         n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578,
         n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588,
         n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598,
         n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608,
         n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618,
         n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628,
         n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638,
         n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648,
         n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658,
         n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668,
         n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678,
         n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688,
         n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698,
         n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708,
         n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718,
         n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728,
         n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738,
         n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748,
         n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758,
         n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768,
         n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778,
         n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788,
         n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798,
         n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808,
         n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818,
         n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828,
         n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838,
         n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848,
         n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858,
         n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868,
         n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878,
         n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888,
         n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898,
         n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908,
         n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918,
         n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928,
         n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938,
         n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948,
         n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958,
         n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968,
         n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978,
         n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988,
         n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998,
         n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008,
         n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018,
         n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028,
         n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038,
         n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048,
         n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058,
         n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068,
         n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078,
         n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088,
         n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098,
         n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108,
         n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118,
         n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128,
         n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138,
         n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148,
         n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158,
         n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168,
         n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178,
         n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188,
         n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198,
         n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208,
         n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218,
         n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228,
         n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238,
         n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248,
         n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258,
         n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268,
         n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278,
         n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288,
         n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298,
         n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308,
         n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318,
         n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328,
         n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338,
         n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348,
         n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358,
         n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368,
         n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378,
         n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388,
         n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398,
         n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408,
         n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418,
         n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428,
         n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438,
         n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448,
         n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458,
         n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468,
         n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478,
         n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488,
         n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498,
         n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508,
         n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518,
         n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528,
         n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538,
         n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548,
         n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558,
         n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568,
         n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578,
         n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588,
         n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598,
         n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608,
         n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618,
         n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628,
         n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638,
         n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648,
         n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658,
         n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668,
         n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678,
         n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688,
         n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698,
         n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708,
         n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718,
         n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728,
         n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738,
         n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748,
         n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758,
         n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768,
         n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778,
         n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788,
         n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798,
         n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808,
         n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818,
         n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828,
         n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838,
         n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848,
         n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858,
         n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868,
         n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878,
         n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888,
         n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898,
         n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908,
         n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918,
         n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928,
         n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938,
         n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948,
         n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958,
         n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968,
         n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978,
         n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988,
         n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998,
         n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008,
         n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018,
         n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028,
         n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038,
         n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048,
         n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058,
         n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068,
         n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078,
         n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088,
         n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098,
         n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108,
         n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118,
         n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128,
         n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138,
         n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148,
         n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158,
         n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168,
         n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178,
         n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188,
         n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198,
         n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208,
         n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218,
         n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228,
         n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238,
         n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248,
         n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258,
         n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268,
         n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278,
         n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288,
         n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298,
         n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308,
         n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318,
         n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328,
         n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338,
         n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348,
         n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358,
         n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368,
         n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378,
         n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388,
         n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398,
         n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408,
         n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418,
         n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428,
         n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438,
         n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448,
         n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458,
         n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468,
         n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478,
         n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488,
         n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498,
         n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508,
         n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518,
         n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528,
         n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538,
         n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548,
         n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558,
         n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568,
         n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578,
         n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588,
         n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598,
         n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608,
         n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618,
         n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628,
         n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638,
         n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648,
         n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658,
         n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668,
         n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678,
         n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688,
         n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698,
         n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708,
         n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718,
         n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728,
         n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738,
         n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748,
         n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758,
         n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768,
         n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778,
         n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788,
         n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798,
         n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808,
         n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818,
         n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828,
         n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838,
         n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848,
         n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858,
         n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868,
         n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878,
         n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888,
         n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898,
         n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908,
         n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918,
         n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928,
         n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938,
         n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948,
         n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958,
         n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968,
         n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978,
         n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988,
         n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998,
         n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008,
         n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018,
         n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028,
         n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038,
         n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048,
         n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058,
         n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068,
         n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078,
         n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088,
         n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098,
         n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108,
         n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118,
         n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128,
         n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138,
         n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148,
         n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158,
         n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168,
         n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178,
         n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188,
         n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198,
         n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208,
         n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218,
         n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228,
         n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238,
         n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248,
         n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258,
         n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268,
         n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278,
         n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288,
         n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298,
         n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308,
         n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318,
         n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328,
         n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338,
         n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348,
         n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358,
         n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368,
         n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378,
         n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388,
         n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398,
         n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408,
         n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418,
         n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428,
         n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438,
         n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448,
         n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458,
         n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468,
         n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478,
         n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488,
         n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498,
         n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508,
         n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518,
         n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528,
         n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538,
         n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548,
         n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558,
         n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568,
         n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578,
         n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588,
         n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598,
         n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608,
         n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618,
         n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628,
         n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638,
         n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648,
         n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659,
         n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669,
         n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679,
         n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689,
         n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699,
         n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709,
         n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719,
         n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729,
         n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739,
         n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749,
         n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759,
         n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769,
         n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779,
         n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789,
         n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799,
         n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809,
         n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819,
         n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829,
         n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839,
         n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849,
         n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859,
         n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869,
         n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879,
         n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889,
         n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899,
         n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909,
         n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919,
         n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929,
         n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939,
         n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949,
         n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959,
         n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969,
         n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979,
         n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989,
         n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999,
         n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198;

  OAI22_X1 U4794 ( .A1(n6890), .A2(n6889), .B1(n6888), .B2(n6887), .ZN(n6977)
         );
  CLKBUF_X1 U4795 ( .A(n6686), .Z(n7321) );
  AND2_X1 U4797 ( .A1(n8842), .A2(n5005), .ZN(n4292) );
  AND2_X2 U4798 ( .A1(n5006), .A2(n5005), .ZN(n4293) );
  CLKBUF_X2 U4799 ( .A(n5806), .Z(n6262) );
  INV_X1 U4801 ( .A(n7482), .ZN(n7452) );
  INV_X1 U4802 ( .A(n6682), .ZN(n6686) );
  INV_X1 U4803 ( .A(n9897), .ZN(n7859) );
  INV_X2 U4805 ( .A(n5665), .ZN(n5581) );
  OAI21_X2 U4806 ( .B1(n4318), .B2(P2_IR_REG_21__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5475) );
  INV_X1 U4807 ( .A(n5600), .ZN(n5696) );
  NAND2_X1 U4808 ( .A1(n5699), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5706) );
  XNOR2_X1 U4809 ( .A(n5475), .B(n5474), .ZN(n7833) );
  INV_X1 U4810 ( .A(n9660), .ZN(n7199) );
  XOR2_X1 U4811 ( .A(n7996), .B(n8682), .Z(n4289) );
  NAND2_X1 U4812 ( .A1(n5711), .A2(n7686), .ZN(n4290) );
  NAND2_X1 U4813 ( .A1(n5711), .A2(n7686), .ZN(n8084) );
  INV_X1 U4814 ( .A(n8084), .ZN(n5862) );
  AND2_X1 U4815 ( .A1(n8842), .A2(n5005), .ZN(n4291) );
  AND2_X1 U4816 ( .A1(n8842), .A2(n5005), .ZN(n5347) );
  OAI21_X2 U4817 ( .B1(n5174), .B2(n4907), .A(n4906), .ZN(n5204) );
  AND2_X1 U4818 ( .A1(n5006), .A2(n5005), .ZN(n4294) );
  INV_X1 U4819 ( .A(n4294), .ZN(n4295) );
  AND2_X2 U4820 ( .A1(n5006), .A2(n5005), .ZN(n5078) );
  INV_X2 U4821 ( .A(n7153), .ZN(n4297) );
  INV_X1 U4822 ( .A(n9667), .ZN(n7285) );
  NAND2_X1 U4823 ( .A1(n7041), .A2(n6286), .ZN(n4320) );
  BUF_X4 U4824 ( .A(n7764), .Z(n4296) );
  INV_X2 U4825 ( .A(n5826), .ZN(n5803) );
  INV_X2 U4826 ( .A(n5050), .ZN(n5305) );
  XNOR2_X1 U4827 ( .A(n5706), .B(n5707), .ZN(n8201) );
  NAND2_X1 U4828 ( .A1(n4982), .A2(n4981), .ZN(n5459) );
  INV_X2 U4829 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  OAI21_X1 U4830 ( .B1(n6281), .B2(n4785), .A(n8901), .ZN(n4784) );
  CLKBUF_X1 U4831 ( .A(n6245), .Z(n8871) );
  NOR2_X1 U4832 ( .A1(n7754), .A2(n7753), .ZN(n8379) );
  XNOR2_X1 U4833 ( .A(n7745), .B(n4357), .ZN(n8400) );
  AOI22_X1 U4834 ( .A1(n7735), .A2(n7734), .B1(n7733), .B2(n7732), .ZN(n8351)
         );
  OR2_X1 U4835 ( .A1(n7654), .A2(n8125), .ZN(n7690) );
  AND2_X1 U4836 ( .A1(n5861), .A2(n7025), .ZN(n7016) );
  NAND2_X1 U4837 ( .A1(n5212), .A2(n5211), .ZN(n8796) );
  NAND2_X1 U4838 ( .A1(n5629), .A2(n5628), .ZN(n9460) );
  AND2_X2 U4839 ( .A1(n6915), .A2(n5502), .ZN(n9944) );
  NAND2_X1 U4840 ( .A1(n5620), .A2(n5619), .ZN(n7645) );
  CLKBUF_X1 U4841 ( .A(n9226), .Z(n9615) );
  NAND2_X1 U4842 ( .A1(n7042), .A2(n6222), .ZN(n7153) );
  NAND2_X1 U4843 ( .A1(n5780), .A2(n8985), .ZN(n7042) );
  INV_X1 U4844 ( .A(n7280), .ZN(n8957) );
  OAI211_X1 U4845 ( .C1(n5029), .C2(n6333), .A(n5113), .B(n5112), .ZN(n9897)
         );
  AND3_X1 U4846 ( .A1(n4343), .A2(n5805), .A3(n5804), .ZN(n7280) );
  INV_X4 U4847 ( .A(n4320), .ZN(n6261) );
  NAND4_X1 U4848 ( .A1(n5832), .A2(n5831), .A3(n5830), .A4(n5829), .ZN(n9668)
         );
  OAI211_X1 U4849 ( .C1(n6340), .C2(n5600), .A(n5580), .B(n5579), .ZN(n9667)
         );
  CLKBUF_X2 U4850 ( .A(n5717), .Z(n4299) );
  AND4_X1 U4851 ( .A1(n5074), .A2(n5073), .A3(n5072), .A4(n5071), .ZN(n6865)
         );
  AND2_X1 U4852 ( .A1(n6222), .A2(n6286), .ZN(n5806) );
  NAND2_X1 U4853 ( .A1(n6675), .A2(n7831), .ZN(n6676) );
  CLKBUF_X1 U4854 ( .A(n5777), .Z(n8206) );
  NAND2_X1 U4855 ( .A1(n5702), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5704) );
  NAND2_X1 U4856 ( .A1(n5777), .A2(n8201), .ZN(n6222) );
  INV_X1 U4857 ( .A(n5770), .ZN(n7686) );
  INV_X2 U4858 ( .A(n5029), .ZN(n7792) );
  INV_X1 U4859 ( .A(n7675), .ZN(n5005) );
  NAND2_X1 U4860 ( .A1(n5004), .A2(n5003), .ZN(n7675) );
  XNOR2_X1 U4861 ( .A(n4998), .B(P2_IR_REG_30__SCAN_IN), .ZN(n8842) );
  NAND2_X1 U4862 ( .A1(n4414), .A2(n4411), .ZN(n8002) );
  OR2_X1 U4863 ( .A1(n9383), .A2(n9385), .ZN(n5710) );
  INV_X2 U4864 ( .A(n8253), .ZN(n8844) );
  INV_X1 U4865 ( .A(n5729), .ZN(n5555) );
  NAND2_X1 U4866 ( .A1(n4976), .A2(n4835), .ZN(n5302) );
  NAND2_X2 U4867 ( .A1(n4749), .A2(n4439), .ZN(n5563) );
  NOR2_X1 U4868 ( .A1(n5551), .A2(n5550), .ZN(n5658) );
  AND2_X1 U4869 ( .A1(n5051), .A2(n4972), .ZN(n5094) );
  AND4_X1 U4870 ( .A1(n5141), .A2(n4970), .A3(n4969), .A4(n4968), .ZN(n4974)
         );
  AND4_X1 U4871 ( .A1(n4971), .A2(n5164), .A3(n10080), .A4(n5257), .ZN(n4973)
         );
  NOR2_X1 U4872 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5051) );
  INV_X1 U4873 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5622) );
  NOR2_X1 U4874 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n5546) );
  INV_X1 U4875 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5634) );
  INV_X1 U4876 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n10080) );
  INV_X4 U4877 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  INV_X1 U4878 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5257) );
  NOR2_X1 U4879 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n4446) );
  NOR2_X1 U4880 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n4970) );
  NOR2_X1 U4881 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n4445) );
  NOR2_X1 U4882 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n4969) );
  NOR2_X1 U4883 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n4968) );
  INV_X1 U4884 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5164) );
  NOR2_X1 U4885 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n5141) );
  NOR2_X1 U4886 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n4971) );
  NAND2_X1 U4887 ( .A1(n6676), .A2(n6926), .ZN(n7764) );
  XNOR2_X1 U4888 ( .A(n5704), .B(n5703), .ZN(n5717) );
  AOI21_X2 U4889 ( .B1(n7552), .B2(n7551), .A(n7550), .ZN(n7553) );
  AOI21_X1 U4890 ( .B1(n5329), .B2(n4960), .A(n4728), .ZN(n4727) );
  INV_X1 U4891 ( .A(n5337), .ZN(n4728) );
  OR2_X1 U4892 ( .A1(n7799), .A2(n7988), .ZN(n7982) );
  AND2_X1 U4893 ( .A1(n4746), .A2(n4745), .ZN(n8241) );
  NOR2_X1 U4894 ( .A1(n5239), .A2(n4720), .ZN(n4719) );
  INV_X1 U4895 ( .A(n4921), .ZN(n4720) );
  NOR2_X1 U4896 ( .A1(n5528), .A2(n8476), .ZN(n8466) );
  NAND2_X1 U4897 ( .A1(n5050), .A2(n5563), .ZN(n5029) );
  NAND2_X1 U4898 ( .A1(n4501), .A2(n4500), .ZN(n4504) );
  AOI21_X1 U4899 ( .B1(n7930), .B2(n8565), .A(n7981), .ZN(n4500) );
  NAND2_X1 U4900 ( .A1(n7931), .A2(n8565), .ZN(n4501) );
  AND2_X1 U4901 ( .A1(n5223), .A2(n5225), .ZN(n4918) );
  INV_X1 U4902 ( .A(n5207), .ZN(n4917) );
  AOI21_X1 U4903 ( .B1(n4304), .B2(n4603), .A(n4520), .ZN(n4602) );
  NOR2_X1 U4904 ( .A1(n4606), .A2(n7970), .ZN(n4603) );
  INV_X1 U4905 ( .A(n8842), .ZN(n5006) );
  NAND2_X1 U4906 ( .A1(n4640), .A2(n4641), .ZN(n4639) );
  INV_X1 U4907 ( .A(n4642), .ZN(n4640) );
  OR2_X1 U4908 ( .A1(n8791), .A2(n7411), .ZN(n8697) );
  OR2_X1 U4909 ( .A1(n9809), .A2(n7412), .ZN(n7895) );
  OR2_X1 U4910 ( .A1(n6687), .A2(n9887), .ZN(n7854) );
  NAND2_X1 U4911 ( .A1(n6673), .A2(n6903), .ZN(n7842) );
  OR2_X1 U4912 ( .A1(n5408), .A2(n8501), .ZN(n5409) );
  AOI21_X1 U4913 ( .B1(n5697), .B2(n5600), .A(n8097), .ZN(n4744) );
  NOR2_X1 U4914 ( .A1(n8140), .A2(n8091), .ZN(n4468) );
  INV_X1 U4915 ( .A(n4693), .ZN(n4692) );
  OAI21_X1 U4916 ( .B1(n8270), .B2(n4694), .A(n8273), .ZN(n4693) );
  INV_X1 U4917 ( .A(n4678), .ZN(n4677) );
  OAI21_X1 U4918 ( .B1(n8264), .B2(n4679), .A(n8267), .ZN(n4678) );
  AND2_X1 U4919 ( .A1(n4355), .A2(n4684), .ZN(n4682) );
  NOR2_X1 U4920 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(n5557), .ZN(n4695) );
  NOR2_X1 U4921 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), .ZN(
        n4791) );
  NAND2_X1 U4922 ( .A1(n4739), .A2(n4738), .ZN(n5540) );
  AOI21_X1 U4923 ( .B1(n4741), .B2(n4743), .A(n4383), .ZN(n4738) );
  NAND2_X1 U4924 ( .A1(n5415), .A2(n4741), .ZN(n4739) );
  NAND2_X1 U4925 ( .A1(n5560), .A2(n4791), .ZN(n5709) );
  INV_X1 U4926 ( .A(n4696), .ZN(n5560) );
  NAND2_X1 U4927 ( .A1(n4722), .A2(n4721), .ZN(n5375) );
  AOI21_X1 U4928 ( .B1(n4724), .B2(n4726), .A(n4384), .ZN(n4721) );
  NAND2_X1 U4929 ( .A1(n5330), .A2(n4724), .ZN(n4722) );
  NAND2_X1 U4930 ( .A1(n4723), .A2(n4727), .ZN(n5340) );
  NAND2_X1 U4931 ( .A1(n5013), .A2(n5012), .ZN(n4730) );
  OAI21_X1 U4932 ( .B1(n5274), .B2(n4938), .A(n4937), .ZN(n5287) );
  NAND2_X1 U4933 ( .A1(n4927), .A2(n4926), .ZN(n5239) );
  NAND2_X1 U4934 ( .A1(n4905), .A2(SI_11_), .ZN(n4906) );
  INV_X1 U4935 ( .A(n5173), .ZN(n4907) );
  OAI21_X1 U4936 ( .B1(n5139), .B2(n5138), .A(n4893), .ZN(n5148) );
  INV_X1 U4937 ( .A(n5347), .ZN(n5423) );
  NAND2_X1 U4938 ( .A1(n4558), .A2(n4557), .ZN(n4556) );
  NOR2_X1 U4939 ( .A1(n7772), .A2(n8731), .ZN(n4557) );
  NOR2_X1 U4940 ( .A1(n8511), .A2(n5451), .ZN(n8502) );
  OR2_X1 U4941 ( .A1(n8731), .A2(n8413), .ZN(n8510) );
  AND2_X1 U4942 ( .A1(n8834), .A2(n8431), .ZN(n5272) );
  AOI21_X1 U4943 ( .B1(n7407), .B2(n4328), .A(n4651), .ZN(n7503) );
  NAND2_X1 U4944 ( .A1(n4652), .A2(n4333), .ZN(n4651) );
  NAND2_X1 U4945 ( .A1(n7794), .A2(n7793), .ZN(n7799) );
  AND2_X1 U4947 ( .A1(n4613), .A2(n4978), .ZN(n4612) );
  NOR2_X1 U4948 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(P2_IR_REG_26__SCAN_IN), .ZN(
        n4613) );
  NAND2_X1 U4949 ( .A1(n4648), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n4749) );
  NAND2_X1 U4950 ( .A1(n4440), .A2(n4750), .ZN(n4439) );
  INV_X1 U4951 ( .A(n4857), .ZN(n4440) );
  AOI21_X1 U4952 ( .B1(n8200), .B2(n9127), .A(n8201), .ZN(n4731) );
  NAND2_X1 U4953 ( .A1(n4735), .A2(n4734), .ZN(n4733) );
  INV_X1 U4954 ( .A(n9345), .ZN(n8999) );
  NOR2_X1 U4955 ( .A1(n9013), .A2(n9248), .ZN(n8996) );
  NAND2_X1 U4956 ( .A1(n8194), .A2(n8237), .ZN(n8322) );
  NOR2_X1 U4957 ( .A1(n9027), .A2(n8073), .ZN(n4687) );
  NAND2_X1 U4958 ( .A1(n4689), .A2(n4688), .ZN(n9004) );
  AND2_X1 U4959 ( .A1(n8287), .A2(n8286), .ZN(n4688) );
  AOI21_X1 U4960 ( .B1(n7450), .B2(n4668), .A(n4666), .ZN(n4665) );
  NAND2_X1 U4961 ( .A1(n4667), .A2(n7649), .ZN(n4666) );
  INV_X1 U4962 ( .A(n7448), .ZN(n4673) );
  OR2_X1 U4963 ( .A1(n9633), .A2(n7047), .ZN(n9236) );
  OR2_X1 U4964 ( .A1(n7057), .A2(n7056), .ZN(n7170) );
  NAND2_X1 U4965 ( .A1(n4418), .A2(n4862), .ZN(n5049) );
  NAND2_X1 U4966 ( .A1(n5028), .A2(n5027), .ZN(n4418) );
  XNOR2_X1 U4967 ( .A(n7752), .B(n7753), .ZN(n8381) );
  NAND2_X1 U4968 ( .A1(n5531), .A2(n9959), .ZN(n4392) );
  AOI21_X1 U4969 ( .B1(n7791), .B2(n5696), .A(n4747), .ZN(n8995) );
  NAND2_X1 U4970 ( .A1(n4513), .A2(n4511), .ZN(n4510) );
  NOR2_X1 U4971 ( .A1(n7879), .A2(n4512), .ZN(n4511) );
  OAI21_X1 U4972 ( .B1(n7871), .B2(n4514), .A(n4331), .ZN(n4513) );
  INV_X1 U4973 ( .A(n7881), .ZN(n4512) );
  NOR2_X1 U4974 ( .A1(n7889), .A2(n4509), .ZN(n4508) );
  INV_X1 U4975 ( .A(n7885), .ZN(n4509) );
  NAND2_X1 U4976 ( .A1(n7901), .A2(n7900), .ZN(n7908) );
  AOI21_X1 U4977 ( .B1(n7893), .B2(n7978), .A(n7892), .ZN(n7901) );
  NAND2_X1 U4978 ( .A1(n8699), .A2(n7911), .ZN(n4518) );
  AND2_X1 U4979 ( .A1(n7923), .A2(n7922), .ZN(n7934) );
  NAND2_X1 U4980 ( .A1(n4515), .A2(n7917), .ZN(n7923) );
  NOR2_X1 U4981 ( .A1(n7950), .A2(n4506), .ZN(n4505) );
  AND2_X1 U4982 ( .A1(n7932), .A2(n7981), .ZN(n4506) );
  NAND2_X1 U4983 ( .A1(n4490), .A2(n4488), .ZN(n4487) );
  NOR2_X1 U4984 ( .A1(n8051), .A2(n4489), .ZN(n4488) );
  NAND2_X1 U4985 ( .A1(n8045), .A2(n4366), .ZN(n4490) );
  NAND2_X1 U4986 ( .A1(n4358), .A2(n8093), .ZN(n4489) );
  OAI21_X1 U4987 ( .B1(n8032), .B2(n4485), .A(n4482), .ZN(n4481) );
  NAND2_X1 U4988 ( .A1(n4486), .A2(n8034), .ZN(n4485) );
  NOR2_X1 U4989 ( .A1(n8170), .A2(n4483), .ZN(n4482) );
  NAND2_X1 U4990 ( .A1(n8493), .A2(n4309), .ZN(n4525) );
  NOR2_X1 U4991 ( .A1(n7965), .A2(n7966), .ZN(n4524) );
  AND2_X1 U4992 ( .A1(n8306), .A2(n4457), .ZN(n4456) );
  NAND2_X1 U4993 ( .A1(n4375), .A2(n8305), .ZN(n4457) );
  AOI21_X1 U4994 ( .B1(n4456), .B2(n4535), .A(n4455), .ZN(n4454) );
  INV_X1 U4995 ( .A(n8308), .ZN(n4455) );
  INV_X1 U4996 ( .A(n8301), .ZN(n4536) );
  INV_X1 U4997 ( .A(n4927), .ZN(n4718) );
  NOR2_X1 U4998 ( .A1(n5127), .A2(n4709), .ZN(n4708) );
  INV_X1 U4999 ( .A(n5108), .ZN(n4709) );
  INV_X1 U5000 ( .A(n4886), .ZN(n4711) );
  OAI21_X1 U5001 ( .B1(n5563), .B2(n4438), .A(n4437), .ZN(n4888) );
  NAND2_X1 U5002 ( .A1(n7359), .A2(n7352), .ZN(n7358) );
  INV_X1 U5003 ( .A(n8333), .ZN(n4819) );
  NAND2_X1 U5004 ( .A1(n4521), .A2(n4519), .ZN(n7973) );
  NAND2_X1 U5005 ( .A1(n8519), .A2(n8338), .ZN(n7956) );
  NOR2_X1 U5006 ( .A1(n4637), .A2(n4394), .ZN(n4393) );
  NAND2_X1 U5007 ( .A1(n4641), .A2(n4644), .ZN(n4637) );
  INV_X1 U5008 ( .A(n4395), .ZN(n4394) );
  OAI211_X1 U5009 ( .C1(n4610), .C2(n8631), .A(n5447), .B(n4608), .ZN(n8564)
         );
  NAND2_X1 U5010 ( .A1(n4611), .A2(n4609), .ZN(n4608) );
  INV_X1 U5011 ( .A(n4611), .ZN(n4610) );
  NAND2_X1 U5012 ( .A1(n4436), .A2(n4338), .ZN(n8565) );
  INV_X1 U5013 ( .A(n8363), .ZN(n4435) );
  NOR2_X1 U5014 ( .A1(n8769), .A2(n8668), .ZN(n4548) );
  INV_X1 U5015 ( .A(n5285), .ZN(n4402) );
  OR2_X1 U5016 ( .A1(n8668), .A2(n8654), .ZN(n7920) );
  OR2_X1 U5017 ( .A1(n5231), .A2(n10091), .ZN(n5247) );
  NAND2_X1 U5018 ( .A1(n9915), .A2(n4563), .ZN(n4562) );
  NOR2_X1 U5019 ( .A1(n6768), .A2(n6960), .ZN(n4552) );
  OR2_X1 U5020 ( .A1(n6673), .A2(n6903), .ZN(n7853) );
  OR2_X1 U5021 ( .A1(n5412), .A2(n5411), .ZN(n5508) );
  NAND2_X1 U5022 ( .A1(n4975), .A2(n4838), .ZN(n4837) );
  INV_X1 U5023 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n4838) );
  NAND2_X1 U5024 ( .A1(n4441), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n4648) );
  INV_X1 U5025 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4441) );
  NOR2_X1 U5026 ( .A1(P1_RD_REG_SCAN_IN), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(
        n4857) );
  NAND2_X1 U5027 ( .A1(n4780), .A2(n4779), .ZN(n4778) );
  INV_X1 U5028 ( .A(n7238), .ZN(n4779) );
  INV_X1 U5029 ( .A(n4777), .ZN(n4776) );
  OAI21_X1 U5030 ( .B1(n4781), .B2(n4778), .A(n7237), .ZN(n4777) );
  NAND2_X1 U5031 ( .A1(n5903), .A2(n8957), .ZN(n5807) );
  NOR2_X1 U5032 ( .A1(n8093), .A2(n4466), .ZN(n4465) );
  INV_X1 U5033 ( .A(n8320), .ZN(n4466) );
  AND2_X1 U5034 ( .A1(n8319), .A2(n8093), .ZN(n4469) );
  NAND2_X1 U5035 ( .A1(n4470), .A2(n4543), .ZN(n4467) );
  NAND2_X1 U5036 ( .A1(n8968), .A2(n8969), .ZN(n8971) );
  OR2_X1 U5037 ( .A1(n9015), .A2(n8288), .ZN(n8319) );
  AND2_X1 U5038 ( .A1(n9027), .A2(n8316), .ZN(n4544) );
  AND2_X1 U5039 ( .A1(n8144), .A2(n9043), .ZN(n8315) );
  OR2_X1 U5040 ( .A1(n9096), .A2(n9289), .ZN(n8312) );
  NOR2_X1 U5041 ( .A1(n9141), .A2(n9157), .ZN(n4581) );
  NOR2_X1 U5042 ( .A1(n9154), .A2(n4539), .ZN(n4538) );
  INV_X1 U5043 ( .A(n8304), .ZN(n4539) );
  INV_X1 U5044 ( .A(n9174), .ZN(n8264) );
  OR2_X1 U5045 ( .A1(n9325), .A2(n9331), .ZN(n8299) );
  OR2_X1 U5046 ( .A1(n7695), .A2(n7694), .ZN(n7717) );
  OR2_X1 U5047 ( .A1(n7500), .A2(n7444), .ZN(n8041) );
  NOR2_X1 U5048 ( .A1(n7168), .A2(n7174), .ZN(n7169) );
  NAND3_X1 U5049 ( .A1(n4588), .A2(n4589), .A3(n7257), .ZN(n7168) );
  NOR2_X1 U5050 ( .A1(n9694), .A2(n9623), .ZN(n4589) );
  INV_X1 U5051 ( .A(n5771), .ZN(n5711) );
  XNOR2_X1 U5052 ( .A(n7040), .B(n8204), .ZN(n8114) );
  NAND2_X1 U5053 ( .A1(n5563), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4567) );
  OR2_X1 U5054 ( .A1(n6344), .A2(n5563), .ZN(n4573) );
  NOR2_X1 U5055 ( .A1(n4317), .A2(n9096), .ZN(n9095) );
  NAND2_X1 U5056 ( .A1(n7450), .A2(n7449), .ZN(n4674) );
  INV_X1 U5057 ( .A(n7038), .ZN(n8204) );
  NOR2_X1 U5058 ( .A1(n7038), .A2(n9640), .ZN(n7200) );
  OAI21_X1 U5059 ( .B1(n5540), .B2(n5539), .A(n5538), .ZN(n5691) );
  NAND2_X1 U5060 ( .A1(n5395), .A2(n5394), .ZN(n5415) );
  NAND2_X1 U5061 ( .A1(n4955), .A2(n4954), .ZN(n5330) );
  NAND2_X1 U5062 ( .A1(n4730), .A2(n4359), .ZN(n4955) );
  NAND2_X1 U5063 ( .A1(n4912), .A2(SI_13_), .ZN(n5207) );
  AOI21_X1 U5064 ( .B1(n5148), .B2(n4701), .A(n4699), .ZN(n4698) );
  NAND2_X1 U5065 ( .A1(n4700), .A2(n4903), .ZN(n4699) );
  NAND2_X1 U5066 ( .A1(n4701), .A2(n4703), .ZN(n4700) );
  INV_X1 U5067 ( .A(n4867), .ZN(n4705) );
  AND2_X1 U5068 ( .A1(n4821), .A2(n8370), .ZN(n4820) );
  INV_X1 U5069 ( .A(n8409), .ZN(n4821) );
  NAND2_X1 U5070 ( .A1(n4826), .A2(n4825), .ZN(n4824) );
  OR2_X1 U5071 ( .A1(n8409), .A2(n4827), .ZN(n4822) );
  INV_X1 U5072 ( .A(n7760), .ZN(n4826) );
  AND2_X1 U5073 ( .A1(n7350), .A2(n7349), .ZN(n7359) );
  NAND2_X1 U5074 ( .A1(n7358), .A2(n7362), .ZN(n4808) );
  OR2_X1 U5075 ( .A1(n5116), .A2(n5115), .ZN(n5132) );
  XNOR2_X1 U5076 ( .A(n6690), .B(n6903), .ZN(n6678) );
  NAND2_X1 U5077 ( .A1(n4801), .A2(n4803), .ZN(n7625) );
  OR2_X1 U5078 ( .A1(n6701), .A2(n9879), .ZN(n6969) );
  NAND2_X1 U5079 ( .A1(n4995), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5344) );
  NAND2_X1 U5080 ( .A1(n7757), .A2(n7758), .ZN(n4827) );
  AND2_X1 U5081 ( .A1(n5428), .A2(n5427), .ZN(n8336) );
  OR2_X1 U5082 ( .A1(n8484), .A2(n5423), .ZN(n5428) );
  OR2_X1 U5083 ( .A1(n5402), .A2(n8335), .ZN(n5421) );
  INV_X1 U5084 ( .A(n4558), .ZN(n4555) );
  NAND2_X1 U5085 ( .A1(n7958), .A2(n7956), .ZN(n8515) );
  NOR2_X1 U5086 ( .A1(n8553), .A2(n8731), .ZN(n8536) );
  OR2_X1 U5087 ( .A1(n8735), .A2(n8372), .ZN(n8529) );
  AOI21_X1 U5088 ( .B1(n8563), .B2(n8566), .A(n4643), .ZN(n8552) );
  AND2_X1 U5089 ( .A1(n8346), .A2(n8546), .ZN(n4643) );
  OR2_X1 U5090 ( .A1(n8572), .A2(n8735), .ZN(n8553) );
  NOR2_X1 U5091 ( .A1(n5328), .A2(n4646), .ZN(n4642) );
  NAND2_X1 U5092 ( .A1(n7929), .A2(n8565), .ZN(n8590) );
  NAND2_X1 U5093 ( .A1(n8631), .A2(n7926), .ZN(n8612) );
  XNOR2_X1 U5094 ( .A(n8751), .B(n8617), .ZN(n8597) );
  NOR2_X1 U5095 ( .A1(n5315), .A2(n4396), .ZN(n4395) );
  NAND2_X1 U5096 ( .A1(n5317), .A2(n5316), .ZN(n4397) );
  INV_X1 U5097 ( .A(n8630), .ZN(n5317) );
  AND2_X1 U5098 ( .A1(n8665), .A2(n4546), .ZN(n8622) );
  AND2_X1 U5099 ( .A1(n4301), .A2(n8626), .ZN(n4546) );
  AND3_X1 U5100 ( .A1(n5021), .A2(n5020), .A3(n5019), .ZN(n8638) );
  NOR2_X1 U5101 ( .A1(n8689), .A2(n8834), .ZN(n8665) );
  NAND2_X1 U5102 ( .A1(n4403), .A2(n4404), .ZN(n8676) );
  NOR2_X1 U5103 ( .A1(n5272), .A2(n8671), .ZN(n4404) );
  AND2_X1 U5104 ( .A1(n7503), .A2(n7918), .ZN(n7505) );
  NAND2_X1 U5105 ( .A1(n4991), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5266) );
  INV_X1 U5106 ( .A(n5247), .ZN(n4991) );
  NOR2_X1 U5107 ( .A1(n8690), .A2(n8786), .ZN(n5436) );
  OAI21_X1 U5108 ( .B1(n7179), .B2(n5198), .A(n4416), .ZN(n7407) );
  AND2_X1 U5109 ( .A1(n5221), .A2(n5202), .ZN(n4416) );
  NAND2_X1 U5110 ( .A1(n7407), .A2(n4323), .ZN(n7596) );
  NAND2_X1 U5111 ( .A1(n4990), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5231) );
  INV_X1 U5112 ( .A(n5214), .ZN(n4990) );
  AOI21_X1 U5113 ( .B1(n5441), .B2(n4300), .A(n4310), .ZN(n9799) );
  OR2_X1 U5114 ( .A1(n9810), .A2(n9809), .ZN(n9811) );
  OR2_X1 U5115 ( .A1(n5192), .A2(n10078), .ZN(n5214) );
  NAND2_X1 U5116 ( .A1(n7425), .A2(n7814), .ZN(n4659) );
  NAND2_X1 U5117 ( .A1(n4661), .A2(n4660), .ZN(n7425) );
  INV_X1 U5118 ( .A(n5200), .ZN(n4660) );
  NAND2_X1 U5119 ( .A1(n9816), .A2(n9824), .ZN(n4661) );
  NOR2_X1 U5120 ( .A1(n9897), .A2(n8440), .ZN(n4408) );
  OAI211_X1 U5121 ( .C1(n7845), .C2(n4595), .A(n7848), .B(n4594), .ZN(n6772)
         );
  NAND2_X1 U5122 ( .A1(n5372), .A2(n5371), .ZN(n8516) );
  NAND2_X1 U5123 ( .A1(n5370), .A2(n8413), .ZN(n5371) );
  NOR2_X1 U5124 ( .A1(n4983), .A2(P2_IR_REG_28__SCAN_IN), .ZN(n5000) );
  NAND2_X1 U5125 ( .A1(n4356), .A2(n4766), .ZN(n4757) );
  NAND2_X1 U5126 ( .A1(n4316), .A2(n4766), .ZN(n4758) );
  OR2_X1 U5127 ( .A1(n6151), .A2(n4765), .ZN(n4759) );
  AND2_X1 U5128 ( .A1(n6154), .A2(n4764), .ZN(n4763) );
  AND2_X1 U5129 ( .A1(n6216), .A2(n6215), .ZN(n6217) );
  NAND2_X1 U5130 ( .A1(n7111), .A2(n7112), .ZN(n4780) );
  NAND2_X1 U5131 ( .A1(n8863), .A2(n8864), .ZN(n8862) );
  OR2_X1 U5132 ( .A1(n5964), .A2(n5944), .ZN(n5946) );
  NAND2_X1 U5133 ( .A1(n4794), .A2(n4793), .ZN(n8881) );
  AND2_X1 U5134 ( .A1(n6046), .A2(n4795), .ZN(n4793) );
  INV_X1 U5135 ( .A(n4780), .ZN(n4775) );
  INV_X1 U5136 ( .A(n4774), .ZN(n4773) );
  OAI21_X1 U5137 ( .B1(n4781), .B2(n4775), .A(n7238), .ZN(n4774) );
  OR2_X1 U5138 ( .A1(n4776), .A2(n4773), .ZN(n4771) );
  NAND2_X1 U5139 ( .A1(n4776), .A2(n4778), .ZN(n4769) );
  NAND3_X1 U5140 ( .A1(n4792), .A2(n6095), .A3(n8933), .ZN(n8916) );
  INV_X1 U5141 ( .A(n8856), .ZN(n6095) );
  OR2_X1 U5142 ( .A1(n7460), .A2(n7462), .ZN(n7582) );
  INV_X1 U5143 ( .A(n5799), .ZN(n6202) );
  OR2_X1 U5144 ( .A1(n5826), .A2(n5815), .ZN(n5819) );
  AND2_X1 U5145 ( .A1(n5771), .A2(n5770), .ZN(n5845) );
  NAND2_X1 U5146 ( .A1(n4624), .A2(n4623), .ZN(n4622) );
  NAND2_X1 U5147 ( .A1(n9492), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n4623) );
  NAND2_X1 U5148 ( .A1(n4622), .A2(n4621), .ZN(n4620) );
  INV_X1 U5149 ( .A(n9428), .ZN(n4621) );
  XNOR2_X1 U5150 ( .A(n8971), .B(n8970), .ZN(n9552) );
  NOR2_X1 U5151 ( .A1(n9552), .A2(n9551), .ZN(n9550) );
  NOR2_X1 U5152 ( .A1(n9576), .A2(n4616), .ZN(n9593) );
  AND2_X1 U5153 ( .A1(n8975), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n4616) );
  NAND2_X1 U5154 ( .A1(n9080), .A2(n4574), .ZN(n9013) );
  NOR2_X1 U5155 ( .A1(n9015), .A2(n4575), .ZN(n4574) );
  INV_X1 U5156 ( .A(n4576), .ZN(n4575) );
  OR2_X1 U5157 ( .A1(n9021), .A2(n9047), .ZN(n8286) );
  AND2_X1 U5158 ( .A1(n8282), .A2(n9035), .ZN(n8283) );
  OR2_X1 U5159 ( .A1(n9065), .A2(n8060), .ZN(n9043) );
  INV_X1 U5160 ( .A(n4531), .ZN(n4530) );
  OAI21_X1 U5161 ( .B1(n8312), .B2(n4532), .A(n9070), .ZN(n4531) );
  NAND2_X1 U5162 ( .A1(n9043), .A2(n8314), .ZN(n9058) );
  AOI21_X1 U5163 ( .B1(n4692), .B2(n4694), .A(n4363), .ZN(n4691) );
  AND2_X1 U5164 ( .A1(n8102), .A2(n8309), .ZN(n9106) );
  INV_X1 U5165 ( .A(n9117), .ZN(n8270) );
  AOI21_X1 U5166 ( .B1(n4677), .B2(n4679), .A(n4364), .ZN(n4676) );
  NAND2_X1 U5167 ( .A1(n4540), .A2(n4538), .ZN(n9149) );
  NAND2_X1 U5168 ( .A1(n9197), .A2(n8301), .ZN(n4540) );
  OR2_X1 U5169 ( .A1(n9179), .A2(n9313), .ZN(n9180) );
  NOR2_X1 U5170 ( .A1(n9180), .A2(n9157), .ZN(n9156) );
  NAND2_X1 U5171 ( .A1(n8265), .A2(n8264), .ZN(n9171) );
  INV_X1 U5172 ( .A(n6050), .ZN(n6048) );
  OR2_X1 U5173 ( .A1(n6002), .A2(n10161), .ZN(n6030) );
  NOR2_X1 U5174 ( .A1(n9237), .A2(n9325), .ZN(n9203) );
  AOI21_X1 U5175 ( .B1(n7691), .B2(n4685), .A(n4339), .ZN(n4684) );
  INV_X1 U5176 ( .A(n7689), .ZN(n4685) );
  INV_X1 U5177 ( .A(n7691), .ZN(n4686) );
  NAND2_X1 U5178 ( .A1(n7718), .A2(n8008), .ZN(n7701) );
  AND2_X1 U5179 ( .A1(n8034), .A2(n8165), .ZN(n8125) );
  AOI21_X1 U5180 ( .B1(n4671), .B2(n4669), .A(n4341), .ZN(n4668) );
  INV_X1 U5181 ( .A(n7449), .ZN(n4669) );
  OR2_X1 U5182 ( .A1(n7481), .A2(n7500), .ZN(n7482) );
  NAND2_X1 U5183 ( .A1(n4664), .A2(n4662), .ZN(n7292) );
  NOR2_X1 U5184 ( .A1(n8118), .A2(n4663), .ZN(n4662) );
  INV_X1 U5185 ( .A(n7270), .ZN(n4663) );
  OAI21_X1 U5186 ( .B1(n7306), .B2(n8117), .A(n7152), .ZN(n7268) );
  NAND2_X1 U5187 ( .A1(n7195), .A2(n7196), .ZN(n7141) );
  NAND2_X1 U5188 ( .A1(n8209), .A2(n8213), .ZN(n8108) );
  INV_X1 U5189 ( .A(n6792), .ZN(n7142) );
  INV_X1 U5190 ( .A(n4573), .ZN(n4570) );
  INV_X1 U5191 ( .A(n5719), .ZN(n4571) );
  AND2_X1 U5192 ( .A1(n9639), .A2(n8242), .ZN(n7037) );
  NAND2_X1 U5193 ( .A1(n5688), .A2(n5687), .ZN(n9248) );
  NAND2_X1 U5194 ( .A1(n8327), .A2(n8326), .ZN(n8328) );
  NAND2_X1 U5195 ( .A1(n5682), .A2(n5681), .ZN(n9265) );
  NAND2_X1 U5196 ( .A1(n5653), .A2(n5652), .ZN(n9320) );
  INV_X1 U5197 ( .A(n8952), .ZN(n7444) );
  AND2_X1 U5198 ( .A1(n5739), .A2(n5738), .ZN(n7054) );
  XNOR2_X1 U5199 ( .A(n5691), .B(n5690), .ZN(n5689) );
  XNOR2_X1 U5200 ( .A(n4545), .B(P1_IR_REG_29__SCAN_IN), .ZN(n5770) );
  NAND2_X1 U5201 ( .A1(n5709), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4545) );
  MUX2_X1 U5202 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5558), .S(
        P1_IR_REG_28__SCAN_IN), .Z(n5559) );
  XNOR2_X1 U5203 ( .A(n5562), .B(n5561), .ZN(n5719) );
  NAND2_X1 U5204 ( .A1(n4696), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5562) );
  AND2_X1 U5205 ( .A1(n4787), .A2(n5732), .ZN(n4526) );
  NAND2_X1 U5206 ( .A1(n5340), .A2(n4967), .ZN(n5357) );
  NAND2_X1 U5207 ( .A1(n4730), .A2(n4951), .ZN(n5319) );
  NAND2_X1 U5208 ( .A1(n5663), .A2(n5662), .ZN(n5699) );
  INV_X1 U5209 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5662) );
  INV_X1 U5210 ( .A(n5661), .ZN(n5663) );
  NAND2_X1 U5211 ( .A1(n4430), .A2(n4941), .ZN(n5301) );
  NAND2_X1 U5212 ( .A1(n5287), .A2(n4939), .ZN(n4430) );
  OR3_X1 U5213 ( .A1(n5644), .A2(P1_IR_REG_15__SCAN_IN), .A3(
        P1_IR_REG_14__SCAN_IN), .ZN(n5648) );
  NAND2_X1 U5214 ( .A1(n4715), .A2(n4927), .ZN(n5255) );
  NAND2_X1 U5215 ( .A1(n4922), .A2(n4719), .ZN(n4715) );
  NAND2_X1 U5216 ( .A1(n4922), .A2(n4921), .ZN(n5240) );
  XNOR2_X1 U5217 ( .A(n5204), .B(n5203), .ZN(n6422) );
  NAND2_X1 U5218 ( .A1(n4647), .A2(n4898), .ZN(n5160) );
  NAND2_X1 U5219 ( .A1(n5148), .A2(n4850), .ZN(n4647) );
  AND2_X1 U5220 ( .A1(n5608), .A2(n5607), .ZN(n6610) );
  XNOR2_X1 U5221 ( .A(n4884), .B(SI_6_), .ZN(n5108) );
  NAND2_X1 U5222 ( .A1(n4883), .A2(n4882), .ZN(n4417) );
  NOR2_X1 U5223 ( .A1(n4881), .A2(n4853), .ZN(n4882) );
  NOR2_X1 U5224 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5541) );
  NOR2_X1 U5225 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n5542) );
  XNOR2_X1 U5226 ( .A(n4861), .B(n4860), .ZN(n5028) );
  NAND2_X1 U5227 ( .A1(n5230), .A2(n5229), .ZN(n8791) );
  INV_X1 U5228 ( .A(n8429), .ZN(n8675) );
  NAND2_X1 U5229 ( .A1(n5419), .A2(n5418), .ZN(n7772) );
  INV_X1 U5230 ( .A(n6903), .ZN(n7102) );
  AOI21_X1 U5231 ( .B1(n8381), .B2(n7751), .A(n7750), .ZN(n7756) );
  INV_X1 U5232 ( .A(n7747), .ZN(n7751) );
  AND4_X1 U5233 ( .A1(n5271), .A2(n5270), .A3(n5269), .A4(n5268), .ZN(n8674)
         );
  INV_X1 U5234 ( .A(n6743), .ZN(n6739) );
  NAND2_X1 U5235 ( .A1(n4443), .A2(n4499), .ZN(n4442) );
  NAND2_X1 U5236 ( .A1(n4498), .A2(n4497), .ZN(n4499) );
  NAND2_X1 U5237 ( .A1(n7999), .A2(n8000), .ZN(n4443) );
  NOR2_X1 U5238 ( .A1(n7998), .A2(n7829), .ZN(n4497) );
  NAND2_X1 U5239 ( .A1(n5518), .A2(n5517), .ZN(n8476) );
  NAND2_X1 U5240 ( .A1(n4604), .A2(n4605), .ZN(n5520) );
  NOR2_X1 U5241 ( .A1(n8487), .A2(n8480), .ZN(n4626) );
  OAI211_X1 U5242 ( .C1(n5413), .C2(n4607), .A(n4633), .B(n4631), .ZN(n8481)
         );
  NAND2_X1 U5243 ( .A1(n4634), .A2(n7824), .ZN(n4633) );
  NAND2_X1 U5244 ( .A1(n5413), .A2(n4632), .ZN(n4631) );
  NAND2_X1 U5245 ( .A1(n8516), .A2(n5506), .ZN(n5413) );
  INV_X1 U5246 ( .A(n4628), .ZN(n4627) );
  OAI21_X1 U5247 ( .B1(n8487), .B2(n4625), .A(n4636), .ZN(n4628) );
  OR2_X1 U5248 ( .A1(n9959), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n4636) );
  OR2_X1 U5249 ( .A1(n8480), .A2(n4629), .ZN(n4625) );
  AOI21_X1 U5250 ( .B1(n8470), .B2(n9941), .A(n4349), .ZN(n5531) );
  INV_X1 U5251 ( .A(n6828), .ZN(n7212) );
  AND3_X1 U5252 ( .A1(n5066), .A2(n5065), .A3(n5064), .ZN(n7225) );
  AND2_X1 U5253 ( .A1(n4980), .A2(n5001), .ZN(n4839) );
  OAI21_X1 U5254 ( .B1(n5471), .B2(P2_IR_REG_26__SCAN_IN), .A(n4347), .ZN(
        n4414) );
  NOR2_X1 U5255 ( .A1(n4413), .A2(n4412), .ZN(n4411) );
  INV_X1 U5256 ( .A(n5567), .ZN(n6288) );
  NAND2_X1 U5257 ( .A1(n5876), .A2(n7027), .ZN(n7114) );
  OR2_X1 U5258 ( .A1(n7525), .A2(n7524), .ZN(n5999) );
  AND2_X1 U5259 ( .A1(n6239), .A2(n4568), .ZN(n8938) );
  NOR2_X1 U5260 ( .A1(n4303), .A2(n8251), .ZN(n4472) );
  OR2_X1 U5261 ( .A1(n8095), .A2(n8096), .ZN(n4737) );
  NAND2_X1 U5262 ( .A1(n4348), .A2(n4475), .ZN(n4474) );
  NAND2_X1 U5263 ( .A1(n4478), .A2(n4479), .ZN(n4475) );
  NOR2_X1 U5264 ( .A1(n8098), .A2(n8985), .ZN(n4479) );
  NOR2_X1 U5265 ( .A1(n5708), .A2(n9236), .ZN(n8991) );
  XNOR2_X1 U5266 ( .A(n8289), .B(n8322), .ZN(n9251) );
  MUX2_X1 U5267 ( .A(n7837), .B(n7836), .S(n7978), .Z(n7862) );
  OR2_X1 U5268 ( .A1(n7870), .A2(n7869), .ZN(n4514) );
  NAND2_X1 U5269 ( .A1(n4507), .A2(n7888), .ZN(n7896) );
  NAND2_X1 U5270 ( .A1(n4510), .A2(n4508), .ZN(n4507) );
  MUX2_X1 U5271 ( .A(n8011), .B(n8010), .S(n8093), .Z(n8019) );
  OAI21_X1 U5272 ( .B1(n4517), .B2(n7914), .A(n4516), .ZN(n4515) );
  INV_X1 U5273 ( .A(n7918), .ZN(n4516) );
  AOI21_X1 U5274 ( .B1(n7908), .B2(n7907), .A(n4518), .ZN(n4517) );
  MUX2_X1 U5275 ( .A(n8028), .B(n8027), .S(n8093), .Z(n8035) );
  AOI211_X1 U5276 ( .C1(n7927), .C2(n7926), .A(n4444), .B(n7939), .ZN(n7931)
         );
  NOR2_X1 U5277 ( .A1(n8046), .A2(n4492), .ZN(n4491) );
  INV_X1 U5278 ( .A(n8044), .ZN(n4492) );
  NAND2_X1 U5279 ( .A1(n4484), .A2(n8014), .ZN(n4483) );
  NAND2_X1 U5280 ( .A1(n8033), .A2(n8034), .ZN(n4484) );
  NOR2_X1 U5281 ( .A1(n8123), .A2(n8167), .ZN(n4486) );
  INV_X1 U5282 ( .A(n7948), .ZN(n7949) );
  NAND2_X1 U5283 ( .A1(n4480), .A2(n4368), .ZN(n8056) );
  NAND2_X1 U5284 ( .A1(n4523), .A2(n4522), .ZN(n4521) );
  INV_X1 U5285 ( .A(n7969), .ZN(n4522) );
  OAI21_X1 U5286 ( .B1(n7960), .B2(n4525), .A(n4524), .ZN(n4523) );
  NOR2_X1 U5287 ( .A1(n7970), .A2(n4520), .ZN(n4519) );
  INV_X1 U5288 ( .A(n7926), .ZN(n4609) );
  INV_X1 U5289 ( .A(n8847), .ZN(n4761) );
  OAI21_X1 U5290 ( .B1(n4373), .B2(n8310), .A(n4449), .ZN(n4448) );
  NAND2_X1 U5291 ( .A1(n4454), .A2(n4452), .ZN(n4451) );
  INV_X1 U5292 ( .A(n4456), .ZN(n4452) );
  NOR2_X1 U5293 ( .A1(n4453), .A2(n8310), .ZN(n4450) );
  INV_X1 U5294 ( .A(n4454), .ZN(n4453) );
  NAND2_X1 U5295 ( .A1(n4581), .A2(n9125), .ZN(n4580) );
  INV_X1 U5296 ( .A(n4742), .ZN(n4741) );
  OAI21_X1 U5297 ( .B1(n5414), .B2(n4743), .A(n5512), .ZN(n4742) );
  INV_X1 U5298 ( .A(n5416), .ZN(n4743) );
  AOI21_X1 U5299 ( .B1(n4727), .B2(n4725), .A(n4374), .ZN(n4724) );
  INV_X1 U5300 ( .A(n4960), .ZN(n4725) );
  INV_X1 U5301 ( .A(n4967), .ZN(n4729) );
  INV_X1 U5302 ( .A(n4727), .ZN(n4726) );
  INV_X1 U5303 ( .A(n5300), .ZN(n4434) );
  AND2_X1 U5304 ( .A1(n4716), .A2(n4427), .ZN(n4426) );
  NAND2_X1 U5305 ( .A1(n4918), .A2(n4913), .ZN(n4427) );
  INV_X1 U5306 ( .A(n4717), .ZN(n4716) );
  OAI21_X1 U5307 ( .B1(n4719), .B2(n4718), .A(n5254), .ZN(n4717) );
  INV_X1 U5308 ( .A(n4933), .ZN(n4714) );
  NAND2_X1 U5309 ( .A1(n4426), .A2(n4424), .ZN(n4423) );
  INV_X1 U5310 ( .A(n4918), .ZN(n4424) );
  OR2_X1 U5311 ( .A1(n5203), .A2(n4917), .ZN(n4913) );
  INV_X1 U5312 ( .A(n4702), .ZN(n4701) );
  OAI21_X1 U5313 ( .B1(n4850), .B2(n4703), .A(n4851), .ZN(n4702) );
  NAND2_X1 U5314 ( .A1(n4890), .A2(n4889), .ZN(n4893) );
  INV_X1 U5315 ( .A(n7759), .ZN(n4825) );
  INV_X1 U5316 ( .A(n7764), .ZN(n6690) );
  AND2_X1 U5317 ( .A1(n8493), .A2(n4607), .ZN(n4606) );
  NOR2_X1 U5318 ( .A1(n8719), .A2(n8519), .ZN(n4558) );
  NOR2_X1 U5319 ( .A1(n8597), .A2(n4444), .ZN(n4611) );
  NAND2_X1 U5320 ( .A1(n7909), .A2(n4653), .ZN(n4652) );
  INV_X1 U5321 ( .A(n5238), .ZN(n4653) );
  AND2_X1 U5322 ( .A1(n9799), .A2(n7895), .ZN(n7410) );
  NAND2_X1 U5323 ( .A1(n4659), .A2(n4658), .ZN(n7404) );
  INV_X1 U5324 ( .A(n5201), .ZN(n4658) );
  NOR2_X1 U5325 ( .A1(n9823), .A2(n4562), .ZN(n4561) );
  AND3_X1 U5326 ( .A1(n7859), .A2(n4552), .A3(n7212), .ZN(n4549) );
  INV_X1 U5327 ( .A(n6919), .ZN(n4550) );
  INV_X1 U5328 ( .A(n6948), .ZN(n4593) );
  OR2_X1 U5329 ( .A1(n8443), .A2(n7225), .ZN(n7838) );
  NAND2_X1 U5330 ( .A1(n7854), .A2(n7856), .ZN(n4596) );
  NAND2_X1 U5331 ( .A1(n8665), .A2(n4548), .ZN(n8656) );
  OR2_X1 U5332 ( .A1(n6919), .A2(n6768), .ZN(n6954) );
  NOR2_X1 U5333 ( .A1(n4837), .A2(P2_IR_REG_19__SCAN_IN), .ZN(n4836) );
  OR2_X1 U5334 ( .A1(n4765), .A2(n4761), .ZN(n4760) );
  NOR2_X1 U5335 ( .A1(n4763), .A2(n4761), .ZN(n4754) );
  INV_X1 U5336 ( .A(n4757), .ZN(n4755) );
  NAND2_X1 U5337 ( .A1(n4465), .A2(n4370), .ZN(n4464) );
  NAND2_X1 U5338 ( .A1(n8199), .A2(n8198), .ZN(n4735) );
  NOR2_X1 U5339 ( .A1(n8239), .A2(n8197), .ZN(n4734) );
  INV_X1 U5340 ( .A(n8200), .ZN(n4736) );
  AND2_X1 U5341 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_REG3_REG_7__SCAN_IN), 
        .ZN(n5881) );
  OR2_X1 U5342 ( .A1(n9248), .A2(n8080), .ZN(n8194) );
  AND2_X1 U5343 ( .A1(n4578), .A2(n4577), .ZN(n4576) );
  NOR2_X1 U5344 ( .A1(n9265), .A2(n9065), .ZN(n4578) );
  INV_X1 U5345 ( .A(n8272), .ZN(n4694) );
  INV_X1 U5346 ( .A(n8266), .ZN(n4679) );
  NOR2_X1 U5347 ( .A1(n7723), .A2(n9460), .ZN(n4585) );
  NAND2_X1 U5348 ( .A1(n4668), .A2(n4672), .ZN(n4667) );
  NAND2_X1 U5349 ( .A1(n5845), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5801) );
  NAND2_X1 U5350 ( .A1(n7142), .A2(n9667), .ZN(n8213) );
  INV_X1 U5351 ( .A(n4542), .ZN(n4541) );
  OAI21_X1 U5352 ( .B1(n4544), .B2(n4306), .A(n8320), .ZN(n4542) );
  AND2_X1 U5353 ( .A1(n9095), .A2(n9085), .ZN(n9080) );
  AOI21_X1 U5354 ( .B1(n4538), .B2(n4536), .A(n4535), .ZN(n4534) );
  INV_X1 U5355 ( .A(n4538), .ZN(n4537) );
  AND2_X1 U5356 ( .A1(n8201), .A2(n8985), .ZN(n8243) );
  AND2_X1 U5357 ( .A1(n4695), .A2(n5561), .ZN(n4587) );
  OAI21_X1 U5358 ( .B1(n5375), .B2(n5374), .A(n5373), .ZN(n5393) );
  INV_X1 U5359 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5732) );
  AND2_X1 U5360 ( .A1(n4967), .A2(n4966), .ZN(n5337) );
  OAI21_X1 U5361 ( .B1(n5287), .B2(n4433), .A(n4431), .ZN(n5013) );
  INV_X1 U5362 ( .A(n4432), .ZN(n4431) );
  OAI21_X1 U5363 ( .B1(n4433), .B2(n4939), .A(n4946), .ZN(n4432) );
  NAND2_X1 U5364 ( .A1(n4434), .A2(n4941), .ZN(n4433) );
  AND2_X1 U5365 ( .A1(n4951), .A2(n4950), .ZN(n5012) );
  OAI21_X1 U5366 ( .B1(n5204), .B2(n4425), .A(n4422), .ZN(n5274) );
  INV_X1 U5367 ( .A(n4426), .ZN(n4425) );
  AND2_X1 U5368 ( .A1(n4423), .A2(n4713), .ZN(n4422) );
  AOI21_X1 U5369 ( .B1(n4716), .B2(n4718), .A(n4714), .ZN(n4713) );
  XNOR2_X1 U5370 ( .A(n4935), .B(SI_17_), .ZN(n5273) );
  NAND2_X1 U5371 ( .A1(n4924), .A2(n4923), .ZN(n4927) );
  NAND2_X1 U5372 ( .A1(n4920), .A2(SI_14_), .ZN(n4921) );
  NAND2_X1 U5373 ( .A1(n5224), .A2(n4918), .ZN(n4922) );
  OR2_X1 U5374 ( .A1(n4917), .A2(n4916), .ZN(n5223) );
  NAND2_X1 U5375 ( .A1(n4429), .A2(n4428), .ZN(n5224) );
  INV_X1 U5376 ( .A(n4913), .ZN(n4428) );
  INV_X1 U5377 ( .A(n5204), .ZN(n4429) );
  XNOR2_X1 U5378 ( .A(n4904), .B(SI_11_), .ZN(n5173) );
  NAND2_X1 U5379 ( .A1(n4707), .A2(n4710), .ZN(n5139) );
  AOI21_X1 U5380 ( .B1(n4887), .B2(n4711), .A(n4340), .ZN(n4710) );
  AND2_X1 U5381 ( .A1(n5086), .A2(n5090), .ZN(n4875) );
  AND2_X1 U5382 ( .A1(n5090), .A2(n4878), .ZN(n4881) );
  NAND2_X1 U5383 ( .A1(n5039), .A2(n5570), .ZN(n4861) );
  NAND2_X1 U5384 ( .A1(n4748), .A2(n4649), .ZN(n4873) );
  NAND2_X1 U5385 ( .A1(n4650), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n4649) );
  INV_X1 U5386 ( .A(n4648), .ZN(n4650) );
  NAND2_X1 U5387 ( .A1(n4987), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5116) );
  NOR2_X1 U5388 ( .A1(n4818), .A2(n4345), .ZN(n4816) );
  NOR2_X1 U5389 ( .A1(n4322), .A2(n4819), .ZN(n4818) );
  INV_X1 U5390 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n5131) );
  OR2_X1 U5391 ( .A1(n5132), .A2(n5131), .ZN(n5154) );
  INV_X1 U5392 ( .A(n7998), .ZN(n6675) );
  OAI21_X1 U5393 ( .B1(n8383), .B2(n8425), .A(n8380), .ZN(n7747) );
  AND2_X1 U5394 ( .A1(n6660), .A2(n6659), .ZN(n6670) );
  OR2_X1 U5395 ( .A1(n5308), .A2(n8354), .ZN(n5310) );
  OR2_X1 U5396 ( .A1(n5310), .A2(n8393), .ZN(n5323) );
  NAND2_X1 U5397 ( .A1(n4994), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n5332) );
  INV_X1 U5398 ( .A(n5323), .ZN(n4994) );
  NAND2_X1 U5399 ( .A1(n4834), .A2(n4833), .ZN(n4829) );
  NAND2_X1 U5400 ( .A1(n4831), .A2(n4833), .ZN(n4828) );
  OR2_X1 U5401 ( .A1(n5364), .A2(n10142), .ZN(n5384) );
  OR2_X1 U5402 ( .A1(n7985), .A2(n7984), .ZN(n4498) );
  AOI21_X1 U5403 ( .B1(n7991), .B2(n7990), .A(n4387), .ZN(n4419) );
  AND2_X1 U5404 ( .A1(n5011), .A2(n5010), .ZN(n8372) );
  AND4_X1 U5405 ( .A1(n5187), .A2(n5186), .A3(n5185), .A4(n5184), .ZN(n5199)
         );
  NOR2_X1 U5406 ( .A1(n4842), .A2(n5509), .ZN(n5510) );
  NAND2_X1 U5407 ( .A1(n8516), .A2(n5507), .ZN(n5511) );
  NAND2_X1 U5408 ( .A1(n4607), .A2(n7964), .ZN(n4605) );
  AND2_X1 U5409 ( .A1(n5421), .A2(n5403), .ZN(n8498) );
  NOR3_X1 U5410 ( .A1(n8509), .A2(n5450), .A3(n8515), .ZN(n8511) );
  AND2_X1 U5411 ( .A1(n8536), .A2(n8814), .ZN(n8517) );
  NAND2_X1 U5412 ( .A1(n8510), .A2(n7954), .ZN(n8530) );
  OR2_X1 U5413 ( .A1(n5344), .A2(n5343), .ZN(n5346) );
  NAND2_X1 U5414 ( .A1(n4996), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5364) );
  INV_X1 U5415 ( .A(n5346), .ZN(n4996) );
  NAND2_X1 U5416 ( .A1(n8529), .A2(n7951), .ZN(n8551) );
  AOI21_X1 U5417 ( .B1(n8564), .B2(n5449), .A(n5448), .ZN(n8544) );
  NAND2_X1 U5418 ( .A1(n4399), .A2(n4398), .ZN(n8563) );
  NAND2_X1 U5419 ( .A1(n4312), .A2(n4644), .ZN(n4398) );
  NAND2_X1 U5420 ( .A1(n4397), .A2(n4393), .ZN(n4399) );
  NAND2_X1 U5421 ( .A1(n8612), .A2(n4611), .ZN(n8603) );
  AND2_X1 U5422 ( .A1(n8622), .A2(n8602), .ZN(n8599) );
  NAND2_X1 U5423 ( .A1(n4405), .A2(n4367), .ZN(n8630) );
  NAND2_X1 U5424 ( .A1(n8676), .A2(n4401), .ZN(n4405) );
  NOR2_X1 U5425 ( .A1(n5299), .A2(n4402), .ZN(n4401) );
  NAND2_X1 U5426 ( .A1(n8634), .A2(n5446), .ZN(n8631) );
  NAND2_X1 U5427 ( .A1(n4993), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5308) );
  INV_X1 U5428 ( .A(n5293), .ZN(n4993) );
  NAND2_X1 U5429 ( .A1(n4600), .A2(n4599), .ZN(n8650) );
  NOR2_X1 U5430 ( .A1(n4848), .A2(n4342), .ZN(n4599) );
  AND2_X1 U5431 ( .A1(n8665), .A2(n8830), .ZN(n8666) );
  OR2_X1 U5432 ( .A1(n5266), .A2(n7558), .ZN(n5279) );
  AND4_X1 U5433 ( .A1(n5253), .A2(n5252), .A3(n5251), .A4(n5250), .ZN(n7607)
         );
  NAND2_X1 U5434 ( .A1(n7409), .A2(n7903), .ZN(n7605) );
  NOR2_X1 U5435 ( .A1(n9811), .A2(n8796), .ZN(n7599) );
  AND4_X1 U5436 ( .A1(n5237), .A2(n5236), .A3(n5235), .A4(n5234), .ZN(n7411)
         );
  AND2_X1 U5437 ( .A1(n7895), .A2(n7897), .ZN(n9800) );
  NAND2_X1 U5438 ( .A1(n4656), .A2(n4654), .ZN(n7885) );
  AND2_X1 U5439 ( .A1(n4655), .A2(n5167), .ZN(n4654) );
  AOI21_X1 U5440 ( .B1(n9841), .B2(n7875), .A(n7883), .ZN(n4598) );
  INV_X1 U5441 ( .A(n9826), .ZN(n9816) );
  NAND2_X1 U5442 ( .A1(n4560), .A2(n4561), .ZN(n9830) );
  NAND2_X1 U5443 ( .A1(n6362), .A2(n7792), .ZN(n4656) );
  OR2_X1 U5444 ( .A1(n5154), .A2(n5153), .ZN(n5181) );
  AND2_X1 U5445 ( .A1(n7884), .A2(n7885), .ZN(n9826) );
  NOR2_X1 U5446 ( .A1(n9858), .A2(n4562), .ZN(n9831) );
  AND2_X1 U5447 ( .A1(n7880), .A2(n7881), .ZN(n7811) );
  OR2_X1 U5448 ( .A1(n9842), .A2(n9841), .ZN(n9845) );
  NOR2_X1 U5449 ( .A1(n9858), .A2(n9857), .ZN(n9859) );
  OAI21_X1 U5450 ( .B1(n7775), .B2(n4409), .A(n4407), .ZN(n9839) );
  NAND2_X1 U5451 ( .A1(n7869), .A2(n4410), .ZN(n4409) );
  AOI21_X1 U5452 ( .B1(n7869), .B2(n4408), .A(n4371), .ZN(n4407) );
  INV_X1 U5453 ( .A(n5114), .ZN(n4410) );
  OR2_X1 U5454 ( .A1(n9839), .A2(n9840), .ZN(n9837) );
  NAND2_X1 U5455 ( .A1(n7782), .A2(n5438), .ZN(n7130) );
  NAND2_X1 U5456 ( .A1(n4592), .A2(n4590), .ZN(n7782) );
  INV_X1 U5457 ( .A(n4591), .ZN(n4590) );
  NAND2_X1 U5458 ( .A1(n4593), .A2(n4335), .ZN(n4592) );
  OAI21_X1 U5459 ( .B1(n6848), .B2(n7840), .A(n7810), .ZN(n4591) );
  NAND2_X1 U5460 ( .A1(n8442), .A2(n9891), .ZN(n7835) );
  NAND2_X1 U5461 ( .A1(n4552), .A2(n7212), .ZN(n4551) );
  NOR2_X1 U5462 ( .A1(n6919), .A2(n4553), .ZN(n6955) );
  INV_X1 U5463 ( .A(n4552), .ZN(n4553) );
  NAND2_X1 U5464 ( .A1(n7839), .A2(n7835), .ZN(n7807) );
  NAND2_X1 U5465 ( .A1(n7838), .A2(n7858), .ZN(n6770) );
  OAI22_X1 U5466 ( .A1(n6925), .A2(n7805), .B1(n6924), .B2(n6687), .ZN(n6765)
         );
  AND2_X1 U5467 ( .A1(n5437), .A2(n7842), .ZN(n7845) );
  INV_X1 U5468 ( .A(n9846), .ZN(n8545) );
  INV_X1 U5469 ( .A(n4596), .ZN(n7805) );
  NOR2_X1 U5470 ( .A1(n7102), .A2(n6972), .ZN(n6920) );
  NAND2_X1 U5471 ( .A1(n7853), .A2(n7842), .ZN(n7803) );
  INV_X1 U5472 ( .A(n9848), .ZN(n8547) );
  AND2_X1 U5473 ( .A1(n8515), .A2(n5409), .ZN(n5506) );
  AND2_X1 U5474 ( .A1(n5508), .A2(n4607), .ZN(n4632) );
  INV_X1 U5475 ( .A(n5508), .ZN(n4634) );
  NAND2_X1 U5476 ( .A1(n9959), .A2(n9932), .ZN(n4629) );
  INV_X1 U5477 ( .A(n8466), .ZN(n5529) );
  AND2_X1 U5478 ( .A1(n5152), .A2(n5151), .ZN(n9915) );
  OAI211_X1 U5479 ( .C1(n5029), .C2(n6343), .A(n5096), .B(n5095), .ZN(n6828)
         );
  AND3_X1 U5480 ( .A1(n5055), .A2(n5054), .A3(n5053), .ZN(n9887) );
  OR2_X1 U5481 ( .A1(n5029), .A2(n6338), .ZN(n5054) );
  INV_X1 U5482 ( .A(n9937), .ZN(n9927) );
  NOR2_X1 U5483 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n4412) );
  INV_X1 U5484 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5474) );
  INV_X1 U5485 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5429) );
  INV_X1 U5486 ( .A(n4837), .ZN(n4835) );
  NAND2_X1 U5487 ( .A1(n8932), .A2(n8935), .ZN(n4792) );
  NAND2_X1 U5488 ( .A1(n4783), .A2(n4782), .ZN(n4781) );
  INV_X1 U5489 ( .A(n7112), .ZN(n4782) );
  INV_X1 U5490 ( .A(n7111), .ZN(n4783) );
  AND2_X1 U5491 ( .A1(n5975), .A2(n7534), .ZN(n7535) );
  NAND2_X1 U5492 ( .A1(n7664), .A2(n7665), .ZN(n4795) );
  OR2_X1 U5493 ( .A1(n7664), .A2(n7665), .ZN(n4796) );
  INV_X1 U5494 ( .A(n4752), .ZN(n8899) );
  OAI21_X1 U5495 ( .B1(n6151), .B2(n4751), .A(n4753), .ZN(n4752) );
  NOR2_X1 U5496 ( .A1(n4755), .A2(n4754), .ZN(n4753) );
  AND2_X1 U5497 ( .A1(n4760), .A2(n4758), .ZN(n4751) );
  OR2_X1 U5498 ( .A1(n5910), .A2(n5909), .ZN(n5962) );
  AND2_X1 U5499 ( .A1(n6114), .A2(n6112), .ZN(n8913) );
  OR2_X1 U5500 ( .A1(n6080), .A2(n6079), .ZN(n6098) );
  NAND2_X1 U5501 ( .A1(n6130), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n6158) );
  INV_X1 U5502 ( .A(n6132), .ZN(n6130) );
  NAND2_X1 U5503 ( .A1(n6076), .A2(n6075), .ZN(n8933) );
  INV_X1 U5504 ( .A(n6074), .ZN(n6075) );
  AND2_X1 U5505 ( .A1(n5858), .A2(n5843), .ZN(n4797) );
  CLKBUF_X1 U5506 ( .A(n7015), .Z(n7026) );
  NAND2_X1 U5507 ( .A1(n4468), .A2(n4336), .ZN(n4461) );
  OAI21_X1 U5508 ( .B1(n8077), .B2(n8076), .A(n8075), .ZN(n8079) );
  NAND2_X1 U5509 ( .A1(n4468), .A2(n4460), .ZN(n4459) );
  INV_X1 U5510 ( .A(n4462), .ZN(n4460) );
  AOI21_X1 U5511 ( .B1(n4307), .B2(n8143), .A(n4463), .ZN(n4462) );
  NAND2_X1 U5512 ( .A1(n4464), .A2(n8323), .ZN(n4463) );
  NAND2_X1 U5513 ( .A1(n9425), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n4619) );
  NOR2_X2 U5514 ( .A1(n5605), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n5659) );
  NOR2_X1 U5515 ( .A1(n6609), .A2(n4369), .ZN(n6613) );
  NOR2_X1 U5516 ( .A1(n6613), .A2(n6612), .ZN(n6804) );
  NOR2_X1 U5517 ( .A1(n6804), .A2(n4617), .ZN(n9542) );
  AND2_X1 U5518 ( .A1(n6805), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4617) );
  NAND2_X1 U5519 ( .A1(n9542), .A2(n9543), .ZN(n9541) );
  NOR2_X1 U5520 ( .A1(n5624), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n5635) );
  NOR2_X1 U5521 ( .A1(n6935), .A2(n4362), .ZN(n6939) );
  NOR2_X1 U5522 ( .A1(n6939), .A2(n6938), .ZN(n7083) );
  NOR2_X1 U5523 ( .A1(n7083), .A2(n4618), .ZN(n8967) );
  AND2_X1 U5524 ( .A1(n7084), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4618) );
  NOR2_X1 U5525 ( .A1(n9550), .A2(n8972), .ZN(n9563) );
  NOR2_X1 U5526 ( .A1(n9593), .A2(n9594), .ZN(n9592) );
  OR2_X1 U5527 ( .A1(n6200), .A2(n6199), .ZN(n8290) );
  NAND2_X1 U5528 ( .A1(n9026), .A2(n8318), .ZN(n9008) );
  AOI21_X1 U5529 ( .B1(n4530), .B2(n4532), .A(n4529), .ZN(n4528) );
  INV_X1 U5530 ( .A(n8314), .ZN(n4529) );
  NAND2_X1 U5531 ( .A1(n9080), .A2(n9354), .ZN(n9062) );
  NAND2_X1 U5532 ( .A1(n9080), .A2(n4578), .ZN(n9038) );
  OR2_X1 U5533 ( .A1(n8278), .A2(n8073), .ZN(n9046) );
  AND2_X1 U5534 ( .A1(n8281), .A2(n8280), .ZN(n9035) );
  OR2_X1 U5535 ( .A1(n8279), .A2(n9056), .ZN(n8281) );
  NAND2_X1 U5536 ( .A1(n9089), .A2(n8312), .ZN(n9074) );
  NAND2_X1 U5537 ( .A1(n9074), .A2(n8313), .ZN(n9072) );
  OAI21_X1 U5538 ( .B1(n9122), .B2(n8270), .A(n8308), .ZN(n9103) );
  AND2_X1 U5539 ( .A1(n8104), .A2(n8308), .ZN(n9117) );
  OAI21_X1 U5540 ( .B1(n9138), .B2(n8269), .A(n8268), .ZN(n9118) );
  AND2_X1 U5541 ( .A1(n8306), .A2(n8105), .ZN(n9137) );
  NOR2_X1 U5542 ( .A1(n9180), .A2(n4579), .ZN(n9139) );
  INV_X1 U5543 ( .A(n4581), .ZN(n4579) );
  AND2_X1 U5544 ( .A1(n8107), .A2(n8302), .ZN(n9174) );
  NAND2_X1 U5545 ( .A1(n6027), .A2(n6026), .ZN(n6050) );
  AND2_X1 U5546 ( .A1(n8296), .A2(n8295), .ZN(n9224) );
  NAND2_X1 U5547 ( .A1(n7658), .A2(n4582), .ZN(n9237) );
  AND2_X1 U5548 ( .A1(n4302), .A2(n4583), .ZN(n4582) );
  AOI21_X1 U5549 ( .B1(n4682), .B2(n4686), .A(n4344), .ZN(n4680) );
  NAND2_X1 U5550 ( .A1(n7658), .A2(n4302), .ZN(n4852) );
  INV_X1 U5551 ( .A(n5946), .ZN(n5930) );
  NAND2_X1 U5552 ( .A1(n7699), .A2(n8127), .ZN(n7718) );
  AND2_X1 U5553 ( .A1(n7642), .A2(n8007), .ZN(n8164) );
  NOR2_X1 U5554 ( .A1(n7482), .A2(n7645), .ZN(n7658) );
  NAND2_X1 U5555 ( .A1(n7264), .A2(n8148), .ZN(n7293) );
  INV_X1 U5556 ( .A(n8955), .ZN(n7294) );
  OAI211_X1 U5557 ( .C1(n6348), .C2(n5600), .A(n5599), .B(n5598), .ZN(n7174)
         );
  NAND2_X1 U5558 ( .A1(n7163), .A2(n7162), .ZN(n7264) );
  INV_X1 U5559 ( .A(n7165), .ZN(n7163) );
  NAND2_X1 U5560 ( .A1(n9625), .A2(n7257), .ZN(n7312) );
  AND2_X1 U5561 ( .A1(n8155), .A2(n8012), .ZN(n8112) );
  OAI21_X1 U5562 ( .B1(n7197), .B2(n4495), .A(n4493), .ZN(n9613) );
  INV_X1 U5563 ( .A(n4494), .ZN(n4493) );
  OAI21_X1 U5564 ( .B1(n7158), .B2(n4495), .A(n8213), .ZN(n4494) );
  INV_X1 U5565 ( .A(n8209), .ZN(n4495) );
  NOR2_X1 U5566 ( .A1(n9624), .A2(n9623), .ZN(n9625) );
  INV_X1 U5567 ( .A(n9236), .ZN(n9626) );
  NAND2_X1 U5568 ( .A1(n7197), .A2(n7158), .ZN(n8154) );
  INV_X1 U5569 ( .A(n7196), .ZN(n8111) );
  NAND2_X1 U5570 ( .A1(n8210), .A2(n7158), .ZN(n7196) );
  NAND2_X1 U5571 ( .A1(n7137), .A2(n8114), .ZN(n7139) );
  NOR2_X1 U5572 ( .A1(n6638), .A2(n8109), .ZN(n8110) );
  AND2_X1 U5573 ( .A1(n8201), .A2(n9127), .ZN(n8242) );
  NAND2_X1 U5574 ( .A1(n5678), .A2(n5677), .ZN(n9278) );
  INV_X1 U5575 ( .A(n8948), .ZN(n9331) );
  NAND2_X1 U5576 ( .A1(n4674), .A2(n4671), .ZN(n7471) );
  NOR2_X1 U5577 ( .A1(n4670), .A2(n7448), .ZN(n7472) );
  INV_X1 U5578 ( .A(n4674), .ZN(n4670) );
  OR2_X1 U5579 ( .A1(n9633), .A2(n8243), .ZN(n9678) );
  OAI211_X1 U5580 ( .C1(n6338), .C2(n5600), .A(n5575), .B(n5574), .ZN(n9660)
         );
  INV_X1 U5581 ( .A(n9678), .ZN(n9695) );
  OAI21_X1 U5582 ( .B1(n5567), .B2(n5573), .A(n5572), .ZN(n9640) );
  NAND2_X1 U5583 ( .A1(n5567), .A2(n9393), .ZN(n5572) );
  INV_X1 U5584 ( .A(SI_30_), .ZN(n4697) );
  AND2_X1 U5585 ( .A1(n4789), .A2(n4695), .ZN(n4496) );
  AND2_X1 U5586 ( .A1(n4791), .A2(n4790), .ZN(n4789) );
  INV_X1 U5587 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n4790) );
  XNOR2_X1 U5588 ( .A(n5540), .B(n5516), .ZN(n7673) );
  XNOR2_X1 U5589 ( .A(n5513), .B(n5512), .ZN(n7545) );
  NAND2_X1 U5590 ( .A1(n4740), .A2(n5416), .ZN(n5513) );
  XNOR2_X1 U5591 ( .A(n5415), .B(n5414), .ZN(n7519) );
  XNOR2_X1 U5592 ( .A(n5210), .B(n5209), .ZN(n6485) );
  OR2_X1 U5593 ( .A1(n5204), .A2(n5203), .ZN(n5206) );
  NAND2_X1 U5594 ( .A1(n4712), .A2(n4886), .ZN(n5128) );
  INV_X1 U5595 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n4788) );
  NAND2_X1 U5596 ( .A1(n4704), .A2(n4657), .ZN(n5087) );
  AOI21_X1 U5597 ( .B1(n4705), .B2(n5061), .A(n4346), .ZN(n4704) );
  OAI21_X1 U5598 ( .B1(P1_IR_REG_1__SCAN_IN), .B2(P1_IR_REG_0__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5576) );
  NAND2_X1 U5599 ( .A1(n4817), .A2(n4322), .ZN(n8334) );
  AND4_X1 U5600 ( .A1(n5220), .A2(n5219), .A3(n5218), .A4(n5217), .ZN(n7606)
         );
  AOI21_X1 U5601 ( .B1(n7364), .B2(n7363), .A(n4807), .ZN(n7365) );
  NOR2_X1 U5602 ( .A1(n7361), .A2(n4808), .ZN(n4807) );
  NAND2_X1 U5603 ( .A1(n7070), .A2(n4805), .ZN(n7364) );
  NOR2_X1 U5604 ( .A1(n7077), .A2(n4806), .ZN(n4805) );
  NAND2_X1 U5605 ( .A1(n7070), .A2(n7069), .ZN(n7076) );
  AND2_X1 U5606 ( .A1(n4325), .A2(n4823), .ZN(n4811) );
  OAI21_X1 U5607 ( .B1(n4823), .B2(n4816), .A(n4813), .ZN(n4812) );
  NAND2_X1 U5608 ( .A1(n4816), .A2(n4814), .ZN(n4813) );
  OR2_X1 U5609 ( .A1(n4325), .A2(n4823), .ZN(n4814) );
  NAND2_X1 U5610 ( .A1(n4816), .A2(n7767), .ZN(n4815) );
  OAI22_X1 U5611 ( .A1(n6700), .A2(n6686), .B1(n6972), .B2(n4296), .ZN(n6717)
         );
  NAND2_X1 U5612 ( .A1(n4830), .A2(n4834), .ZN(n8362) );
  NAND2_X1 U5613 ( .A1(n8349), .A2(n4305), .ZN(n4830) );
  NAND2_X1 U5614 ( .A1(n7625), .A2(n7624), .ZN(n7679) );
  NAND2_X1 U5615 ( .A1(n4985), .A2(n4984), .ZN(n8735) );
  NAND2_X1 U5616 ( .A1(n8349), .A2(n7739), .ZN(n8392) );
  AND4_X1 U5617 ( .A1(n5197), .A2(n5196), .A3(n5195), .A4(n5194), .ZN(n7412)
         );
  NAND2_X1 U5618 ( .A1(n4436), .A2(n5331), .ZN(n8745) );
  AND4_X1 U5619 ( .A1(n5122), .A2(n5121), .A3(n5120), .A4(n5119), .ZN(n9847)
         );
  INV_X1 U5620 ( .A(n8441), .ZN(n6951) );
  INV_X1 U5621 ( .A(n4827), .ZN(n4810) );
  NAND2_X1 U5622 ( .A1(n5245), .A2(n5244), .ZN(n8786) );
  NAND2_X1 U5623 ( .A1(n6662), .A2(n8556), .ZN(n8420) );
  OR2_X1 U5624 ( .A1(n8521), .A2(n5423), .ZN(n5391) );
  AND3_X1 U5625 ( .A1(n5336), .A2(n5335), .A3(n5334), .ZN(n8363) );
  INV_X1 U5626 ( .A(n6865), .ZN(n8442) );
  AND2_X1 U5627 ( .A1(n5023), .A2(n5022), .ZN(n5026) );
  NAND4_X1 U5628 ( .A1(n5036), .A2(n5035), .A3(n5034), .A4(n5033), .ZN(n6701)
         );
  OAI211_X1 U5629 ( .C1(n5511), .C2(n7826), .A(n4389), .B(n4388), .ZN(n8470)
         );
  NAND2_X1 U5630 ( .A1(n4390), .A2(n5521), .ZN(n4389) );
  NAND2_X1 U5631 ( .A1(n5511), .A2(n4308), .ZN(n4388) );
  INV_X1 U5632 ( .A(n5510), .ZN(n4390) );
  NAND2_X1 U5633 ( .A1(n5363), .A2(n5362), .ZN(n8731) );
  INV_X1 U5634 ( .A(n8745), .ZN(n8586) );
  NAND2_X1 U5635 ( .A1(n4638), .A2(n4641), .ZN(n8582) );
  NAND2_X1 U5636 ( .A1(n8755), .A2(n4642), .ZN(n4638) );
  NAND2_X1 U5637 ( .A1(n8755), .A2(n4645), .ZN(n8598) );
  NAND2_X1 U5638 ( .A1(n4397), .A2(n4395), .ZN(n8755) );
  AND2_X1 U5639 ( .A1(n4397), .A2(n4400), .ZN(n8621) );
  NAND2_X1 U5640 ( .A1(n8665), .A2(n4301), .ZN(n8623) );
  NAND2_X1 U5641 ( .A1(n8676), .A2(n5285), .ZN(n8648) );
  AND2_X1 U5642 ( .A1(n4600), .A2(n4601), .ZN(n8670) );
  NOR2_X1 U5643 ( .A1(n7505), .A2(n5272), .ZN(n8678) );
  NAND2_X1 U5644 ( .A1(n7596), .A2(n5238), .ZN(n8688) );
  AND2_X1 U5645 ( .A1(n7407), .A2(n5222), .ZN(n7597) );
  NAND2_X1 U5646 ( .A1(n5191), .A2(n5190), .ZN(n9809) );
  INV_X1 U5647 ( .A(n4659), .ZN(n7426) );
  OAI21_X1 U5648 ( .B1(n7775), .B2(n5114), .A(n4406), .ZN(n7123) );
  INV_X1 U5649 ( .A(n4408), .ZN(n4406) );
  INV_X1 U5650 ( .A(n9856), .ZN(n8693) );
  NOR2_X1 U5651 ( .A1(n9866), .A2(n6927), .ZN(n9834) );
  OR2_X1 U5652 ( .A1(n9868), .A2(n6663), .ZN(n8556) );
  AND2_X1 U5653 ( .A1(n7790), .A2(n7789), .ZN(n8810) );
  AND2_X1 U5654 ( .A1(n8716), .A2(n8715), .ZN(n8807) );
  AOI21_X1 U5655 ( .B1(n8481), .B2(n9941), .A(n4635), .ZN(n5503) );
  INV_X1 U5656 ( .A(n4626), .ZN(n4635) );
  AND2_X1 U5657 ( .A1(n5342), .A2(n5341), .ZN(n8819) );
  NAND2_X1 U5658 ( .A1(n5265), .A2(n5264), .ZN(n8834) );
  OAI21_X1 U5659 ( .B1(n6344), .B2(n5029), .A(n5032), .ZN(n4415) );
  INV_X1 U5660 ( .A(n9944), .ZN(n9942) );
  NAND2_X1 U5661 ( .A1(n5003), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4998) );
  MUX2_X1 U5662 ( .A(n5002), .B(P2_IR_REG_31__SCAN_IN), .S(n5001), .Z(n5004)
         );
  OR2_X1 U5663 ( .A1(n5000), .A2(n4999), .ZN(n5002) );
  MUX2_X1 U5664 ( .A(P2_IR_REG_31__SCAN_IN), .B(n4979), .S(
        P2_IR_REG_28__SCAN_IN), .Z(n4982) );
  XNOR2_X1 U5665 ( .A(n5478), .B(n5477), .ZN(n9870) );
  AND2_X1 U5666 ( .A1(n5175), .A2(n5166), .ZN(n9770) );
  AOI21_X1 U5667 ( .B1(n6248), .B2(n6220), .A(n6219), .ZN(n4785) );
  NAND2_X1 U5668 ( .A1(n4756), .A2(n4757), .ZN(n8846) );
  OR2_X1 U5669 ( .A1(n6151), .A2(n4758), .ZN(n4756) );
  NAND2_X1 U5670 ( .A1(n5676), .A2(n5675), .ZN(n9096) );
  NAND2_X1 U5671 ( .A1(n4792), .A2(n8933), .ZN(n8855) );
  NAND2_X1 U5672 ( .A1(n5668), .A2(n5667), .ZN(n9157) );
  AND2_X1 U5673 ( .A1(n6248), .A2(n4376), .ZN(n6281) );
  NAND2_X1 U5674 ( .A1(n4772), .A2(n4780), .ZN(n7240) );
  NAND2_X1 U5675 ( .A1(n7114), .A2(n4781), .ZN(n4772) );
  NAND2_X1 U5676 ( .A1(n4794), .A2(n4795), .ZN(n8884) );
  NAND2_X1 U5677 ( .A1(n5647), .A2(n5646), .ZN(n9325) );
  INV_X1 U5678 ( .A(n9687), .ZN(n7166) );
  AND2_X1 U5679 ( .A1(n4769), .A2(n4768), .ZN(n4767) );
  NAND2_X1 U5680 ( .A1(n7114), .A2(n4771), .ZN(n4770) );
  NAND2_X1 U5681 ( .A1(n4773), .A2(n4775), .ZN(n4768) );
  OR2_X1 U5682 ( .A1(n6151), .A2(n6152), .ZN(n8928) );
  OAI211_X1 U5683 ( .C1(n6333), .C2(n5600), .A(n5594), .B(n5593), .ZN(n9694)
         );
  NAND2_X1 U5684 ( .A1(n6245), .A2(n4786), .ZN(n6248) );
  AND2_X1 U5685 ( .A1(n6246), .A2(n6247), .ZN(n4786) );
  OAI21_X1 U5686 ( .B1(n9042), .B2(n8910), .A(n6252), .ZN(n6253) );
  INV_X1 U5687 ( .A(n8910), .ZN(n8942) );
  NAND4_X1 U5688 ( .A1(n5968), .A2(n5967), .A3(n5966), .A4(n5965), .ZN(n8952)
         );
  NAND4_X1 U5689 ( .A1(n5854), .A2(n5853), .A3(n5852), .A4(n5851), .ZN(n9614)
         );
  OR2_X1 U5690 ( .A1(n8082), .A2(n6303), .ZN(n5853) );
  NAND2_X1 U5691 ( .A1(n4319), .A2(n5820), .ZN(n6792) );
  AND2_X1 U5692 ( .A1(n5788), .A2(n5787), .ZN(n5789) );
  INV_X1 U5693 ( .A(n4622), .ZN(n9427) );
  INV_X1 U5694 ( .A(n4620), .ZN(n9426) );
  AND2_X1 U5695 ( .A1(n5542), .A2(n5541), .ZN(n5582) );
  XNOR2_X1 U5696 ( .A(n8967), .B(n7088), .ZN(n7085) );
  XNOR2_X1 U5697 ( .A(n4614), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n8984) );
  OR2_X1 U5698 ( .A1(n9592), .A2(n4615), .ZN(n4614) );
  AND2_X1 U5699 ( .A1(n8979), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n4615) );
  AOI211_X1 U5700 ( .C1(n9000), .C2(n8999), .A(n9236), .B(n8998), .ZN(n9245)
         );
  NAND2_X1 U5701 ( .A1(n4689), .A2(n8286), .ZN(n9005) );
  NAND2_X1 U5702 ( .A1(n8285), .A2(n8284), .ZN(n9020) );
  OAI21_X1 U5703 ( .B1(n9089), .B2(n4532), .A(n4530), .ZN(n9052) );
  INV_X1 U5704 ( .A(n9075), .ZN(n9289) );
  NAND2_X1 U5705 ( .A1(n9116), .A2(n8272), .ZN(n9107) );
  NAND2_X1 U5706 ( .A1(n5674), .A2(n5673), .ZN(n9286) );
  NAND2_X1 U5707 ( .A1(n8271), .A2(n8270), .ZN(n9116) );
  NAND2_X1 U5708 ( .A1(n5672), .A2(n5671), .ZN(n9296) );
  NAND2_X1 U5709 ( .A1(n9171), .A2(n8266), .ZN(n9155) );
  NAND2_X1 U5710 ( .A1(n4540), .A2(n8304), .ZN(n9151) );
  NAND2_X1 U5711 ( .A1(n5657), .A2(n5656), .ZN(n9313) );
  NAND2_X1 U5712 ( .A1(n4683), .A2(n4684), .ZN(n8258) );
  OR2_X1 U5713 ( .A1(n7690), .A2(n4686), .ZN(n4683) );
  NAND2_X1 U5714 ( .A1(n7690), .A2(n7689), .ZN(n7715) );
  OAI21_X1 U5715 ( .B1(n7450), .B2(n4672), .A(n4668), .ZN(n7650) );
  NAND2_X1 U5716 ( .A1(n5615), .A2(n5614), .ZN(n7500) );
  NAND2_X1 U5717 ( .A1(n5611), .A2(n5610), .ZN(n7468) );
  INV_X1 U5718 ( .A(n9622), .ZN(n9204) );
  INV_X1 U5719 ( .A(n9646), .ZN(n9206) );
  INV_X1 U5720 ( .A(n9222), .ZN(n9231) );
  OR2_X1 U5721 ( .A1(n5826), .A2(n5825), .ZN(n5831) );
  NAND2_X1 U5722 ( .A1(n4571), .A2(n4570), .ZN(n4569) );
  NAND2_X1 U5723 ( .A1(n5718), .A2(n4329), .ZN(n4572) );
  AOI21_X1 U5724 ( .B1(n4568), .B2(n4566), .A(n4565), .ZN(n4564) );
  AND2_X1 U5725 ( .A1(n5565), .A2(n5564), .ZN(n9345) );
  INV_X1 U5726 ( .A(n9096), .ZN(n9358) );
  OR2_X1 U5727 ( .A1(n6234), .A2(n5764), .ZN(n9718) );
  AND2_X1 U5728 ( .A1(n6235), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9654) );
  OAI21_X1 U5729 ( .B1(n5689), .B2(n4697), .A(n5692), .ZN(n5695) );
  CLKBUF_X1 U5730 ( .A(n5719), .Z(n9479) );
  XNOR2_X1 U5731 ( .A(n5724), .B(P1_IR_REG_26__SCAN_IN), .ZN(n7385) );
  INV_X1 U5732 ( .A(n8206), .ZN(n8197) );
  AND2_X1 U5733 ( .A1(n5654), .A2(n5651), .ZN(n8975) );
  INV_X1 U5734 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6363) );
  INV_X1 U5735 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6361) );
  INV_X1 U5736 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6330) );
  NAND2_X1 U5737 ( .A1(n4706), .A2(n4867), .ZN(n5062) );
  NAND2_X1 U5738 ( .A1(n5049), .A2(n5048), .ZN(n4706) );
  XNOR2_X1 U5739 ( .A(n5566), .B(P1_IR_REG_1__SCAN_IN), .ZN(n6630) );
  INV_X1 U5740 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n9394) );
  NAND2_X1 U5741 ( .A1(n6827), .A2(n6826), .ZN(n6862) );
  AOI21_X1 U5742 ( .B1(n4289), .B2(n4385), .A(n4442), .ZN(n8006) );
  NAND2_X1 U5743 ( .A1(n4392), .A2(n4391), .ZN(n5530) );
  OR2_X1 U5744 ( .A1(n9959), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n4391) );
  OAI21_X1 U5745 ( .B1(n8481), .B2(n4630), .A(n4627), .ZN(n5499) );
  OR2_X1 U5746 ( .A1(n8250), .A2(n8249), .ZN(n4476) );
  NAND2_X1 U5747 ( .A1(n4474), .A2(n4477), .ZN(n4473) );
  OR2_X1 U5748 ( .A1(n9251), .A2(n9222), .ZN(n4533) );
  MUX2_X1 U5749 ( .A(n5755), .B(n5765), .S(n9733), .Z(n5758) );
  MUX2_X1 U5750 ( .A(n5712), .B(n5765), .S(n9720), .Z(n5768) );
  NOR2_X1 U5751 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n4787) );
  NOR2_X1 U5752 ( .A1(n9796), .A2(n9807), .ZN(n4300) );
  AND2_X1 U5753 ( .A1(n4548), .A2(n4547), .ZN(n4301) );
  AND2_X1 U5754 ( .A1(n4585), .A2(n4584), .ZN(n4302) );
  AND2_X1 U5755 ( .A1(n4348), .A2(n4311), .ZN(n4303) );
  XNOR2_X1 U5757 ( .A(n5710), .B(P1_IR_REG_30__SCAN_IN), .ZN(n5771) );
  INV_X1 U5758 ( .A(n7831), .ZN(n7989) );
  AND2_X1 U5759 ( .A1(n4605), .A2(n5519), .ZN(n4304) );
  NOR2_X1 U5760 ( .A1(n8391), .A2(n7738), .ZN(n4305) );
  OR2_X1 U5761 ( .A1(n8321), .A2(n4543), .ZN(n4306) );
  AND2_X1 U5762 ( .A1(n4467), .A2(n4469), .ZN(n4307) );
  NAND2_X1 U5763 ( .A1(n5519), .A2(n7967), .ZN(n7824) );
  INV_X1 U5764 ( .A(n7824), .ZN(n4607) );
  NAND2_X1 U5765 ( .A1(n5277), .A2(n5276), .ZN(n8668) );
  NAND2_X1 U5766 ( .A1(n5633), .A2(n5632), .ZN(n7723) );
  NAND2_X1 U5767 ( .A1(n4976), .A2(n4836), .ZN(n5431) );
  AND2_X1 U5768 ( .A1(n5510), .A2(n7826), .ZN(n4308) );
  NAND2_X1 U5769 ( .A1(n7959), .A2(n7978), .ZN(n4309) );
  INV_X1 U5770 ( .A(n8719), .ZN(n8500) );
  NAND2_X1 U5771 ( .A1(n5401), .A2(n5400), .ZN(n8719) );
  NOR2_X1 U5772 ( .A1(n9807), .A2(n9797), .ZN(n4310) );
  NAND2_X1 U5773 ( .A1(n4478), .A2(n4386), .ZN(n4311) );
  INV_X1 U5774 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5544) );
  NAND2_X1 U5775 ( .A1(n8602), .A2(n8617), .ZN(n4641) );
  INV_X1 U5776 ( .A(n4800), .ZN(n4799) );
  OR2_X1 U5777 ( .A1(n7678), .A2(n7623), .ZN(n4800) );
  NAND2_X1 U5778 ( .A1(n4639), .A2(n8590), .ZN(n4312) );
  AND2_X1 U5779 ( .A1(n4561), .A2(n4559), .ZN(n4313) );
  AND2_X1 U5780 ( .A1(n4836), .A2(n4327), .ZN(n4314) );
  NAND2_X1 U5781 ( .A1(n7658), .A2(n7659), .ZN(n4315) );
  NOR2_X1 U5782 ( .A1(n8639), .A2(n8428), .ZN(n5315) );
  OR2_X1 U5783 ( .A1(n4762), .A2(n8926), .ZN(n4316) );
  INV_X1 U5784 ( .A(n8189), .ZN(n4449) );
  INV_X1 U5785 ( .A(n8305), .ZN(n4535) );
  INV_X1 U5786 ( .A(n8639), .ZN(n4547) );
  NAND2_X1 U5787 ( .A1(n5637), .A2(n5636), .ZN(n8257) );
  INV_X1 U5788 ( .A(n8257), .ZN(n4584) );
  AND2_X1 U5789 ( .A1(n5433), .A2(n4318), .ZN(n7829) );
  OR3_X1 U5790 ( .A1(n9180), .A2(n9286), .A3(n4580), .ZN(n4317) );
  OR2_X1 U5791 ( .A1(n5431), .A2(P2_IR_REG_20__SCAN_IN), .ZN(n4318) );
  NAND2_X1 U5792 ( .A1(n7280), .A2(n9660), .ZN(n7158) );
  INV_X1 U5793 ( .A(n5092), .ZN(n5109) );
  INV_X2 U5794 ( .A(n5109), .ZN(n7788) );
  AND3_X1 U5795 ( .A1(n5819), .A2(n5818), .A3(n5817), .ZN(n4319) );
  XNOR2_X1 U5796 ( .A(n5695), .B(n5694), .ZN(n7791) );
  INV_X1 U5797 ( .A(n5845), .ZN(n5827) );
  NAND3_X1 U5798 ( .A1(n5791), .A2(n5790), .A3(n5789), .ZN(n7040) );
  OAI211_X1 U5799 ( .C1(n5776), .C2(n5826), .A(n5775), .B(n5774), .ZN(n6638)
         );
  NAND4_X1 U5800 ( .A1(n5047), .A2(n5046), .A3(n5045), .A4(n5044), .ZN(n6687)
         );
  AND2_X1 U5801 ( .A1(n9080), .A2(n4576), .ZN(n4321) );
  AND2_X1 U5802 ( .A1(n4822), .A2(n4824), .ZN(n4322) );
  NOR2_X1 U5803 ( .A1(n8553), .A2(n4556), .ZN(n4554) );
  INV_X1 U5804 ( .A(n4672), .ZN(n4671) );
  NAND2_X1 U5805 ( .A1(n8120), .A2(n4673), .ZN(n4672) );
  AND2_X1 U5806 ( .A1(n7902), .A2(n5222), .ZN(n4323) );
  NAND2_X1 U5807 ( .A1(n5872), .A2(n5873), .ZN(n4324) );
  NAND2_X1 U5808 ( .A1(n5770), .A2(n5711), .ZN(n5799) );
  AND2_X1 U5809 ( .A1(n8333), .A2(n4820), .ZN(n4325) );
  INV_X1 U5810 ( .A(n7987), .ZN(n4520) );
  AND2_X1 U5811 ( .A1(n8925), .A2(n8926), .ZN(n4326) );
  AND4_X1 U5812 ( .A1(n4977), .A2(n9995), .A3(n5474), .A4(n5429), .ZN(n4327)
         );
  AND2_X1 U5813 ( .A1(n4323), .A2(n7909), .ZN(n4328) );
  AND2_X1 U5814 ( .A1(n5719), .A2(n6630), .ZN(n4329) );
  NAND2_X1 U5815 ( .A1(n6151), .A2(n6152), .ZN(n8925) );
  AND3_X1 U5816 ( .A1(n5658), .A2(n5553), .A3(n5552), .ZN(n4330) );
  OR2_X1 U5817 ( .A1(n8757), .A2(n8638), .ZN(n8615) );
  INV_X1 U5818 ( .A(n8615), .ZN(n4444) );
  AND2_X1 U5819 ( .A1(n7874), .A2(n9840), .ZN(n4331) );
  AND2_X1 U5820 ( .A1(n4759), .A2(n4763), .ZN(n4332) );
  NAND2_X1 U5821 ( .A1(n5555), .A2(n5554), .ZN(n5722) );
  NAND2_X1 U5822 ( .A1(n5291), .A2(n5290), .ZN(n8769) );
  OR2_X1 U5823 ( .A1(n8786), .A2(n8432), .ZN(n4333) );
  AND2_X1 U5824 ( .A1(n4620), .A2(n4619), .ZN(n4334) );
  NAND2_X1 U5825 ( .A1(n5771), .A2(n7686), .ZN(n5826) );
  NOR2_X1 U5826 ( .A1(n7807), .A2(n7840), .ZN(n4335) );
  NAND2_X1 U5827 ( .A1(n4656), .A2(n5167), .ZN(n9823) );
  INV_X1 U5828 ( .A(n5127), .ZN(n4887) );
  XNOR2_X1 U5829 ( .A(n4888), .B(SI_7_), .ZN(n5127) );
  OR2_X1 U5830 ( .A1(n4307), .A2(n4465), .ZN(n4336) );
  AND2_X1 U5831 ( .A1(n5092), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n4337) );
  INV_X1 U5832 ( .A(n8251), .ZN(n4477) );
  AND2_X1 U5833 ( .A1(n4435), .A2(n5331), .ZN(n4338) );
  OR2_X1 U5834 ( .A1(n7772), .A2(n8336), .ZN(n5519) );
  AND2_X1 U5835 ( .A1(n7723), .A2(n9459), .ZN(n4339) );
  AND2_X1 U5836 ( .A1(n4888), .A2(SI_7_), .ZN(n4340) );
  INV_X1 U5837 ( .A(n4898), .ZN(n4703) );
  NAND2_X1 U5838 ( .A1(n4895), .A2(n4894), .ZN(n4898) );
  AND2_X1 U5839 ( .A1(n8149), .A2(n8029), .ZN(n8118) );
  NOR2_X1 U5840 ( .A1(n7500), .A2(n8952), .ZN(n4341) );
  INV_X1 U5841 ( .A(n8814), .ZN(n8519) );
  NAND2_X1 U5842 ( .A1(n8669), .A2(n7920), .ZN(n4342) );
  INV_X1 U5843 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9385) );
  NAND2_X1 U5844 ( .A1(n7961), .A2(n7962), .ZN(n8501) );
  XNOR2_X1 U5845 ( .A(n5835), .B(n4298), .ZN(n5840) );
  INV_X1 U5846 ( .A(n4646), .ZN(n4645) );
  NOR2_X1 U5847 ( .A1(n8626), .A2(n8638), .ZN(n4646) );
  AND2_X1 U5848 ( .A1(n5801), .A2(n5800), .ZN(n4343) );
  NOR2_X1 U5849 ( .A1(n8257), .A2(n9225), .ZN(n4344) );
  AND2_X1 U5850 ( .A1(n7763), .A2(n7762), .ZN(n4345) );
  INV_X1 U5851 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5303) );
  AND2_X1 U5852 ( .A1(n4871), .A2(SI_3_), .ZN(n4346) );
  AND2_X1 U5853 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n4347) );
  AND2_X1 U5854 ( .A1(n4732), .A2(n4731), .ZN(n4348) );
  NAND2_X1 U5855 ( .A1(n8479), .A2(n8473), .ZN(n4349) );
  OAI21_X1 U5856 ( .B1(n4305), .B2(n4832), .A(n8361), .ZN(n4831) );
  OR2_X1 U5857 ( .A1(n8476), .A2(n6784), .ZN(n7986) );
  NAND2_X1 U5858 ( .A1(n5700), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5705) );
  OR2_X1 U5859 ( .A1(n8719), .A2(n8412), .ZN(n7961) );
  AND2_X1 U5860 ( .A1(n4604), .A2(n4304), .ZN(n4350) );
  AND4_X1 U5861 ( .A1(n5172), .A2(n5171), .A3(n5170), .A4(n5169), .ZN(n7232)
         );
  INV_X1 U5862 ( .A(n7232), .ZN(n4655) );
  NAND2_X1 U5863 ( .A1(n5479), .A2(n4612), .ZN(n4983) );
  INV_X1 U5864 ( .A(n4983), .ZN(n4413) );
  AND2_X1 U5865 ( .A1(n6826), .A2(n6829), .ZN(n4351) );
  AND2_X1 U5866 ( .A1(n8118), .A2(n8148), .ZN(n4352) );
  AND2_X1 U5867 ( .A1(n4849), .A2(n7903), .ZN(n4353) );
  AND2_X1 U5868 ( .A1(n7700), .A2(n8008), .ZN(n4354) );
  NAND2_X1 U5869 ( .A1(n8257), .A2(n9225), .ZN(n4355) );
  AND2_X1 U5870 ( .A1(n8318), .A2(n8100), .ZN(n9027) );
  NAND2_X1 U5871 ( .A1(n4770), .A2(n4767), .ZN(n7460) );
  NAND2_X1 U5872 ( .A1(n5479), .A2(n4978), .ZN(n5471) );
  OR2_X1 U5873 ( .A1(n9021), .A2(n8078), .ZN(n8318) );
  INV_X1 U5874 ( .A(n8318), .ZN(n4543) );
  AND2_X1 U5875 ( .A1(n8926), .A2(n4762), .ZN(n4356) );
  NAND2_X1 U5876 ( .A1(n4681), .A2(n4680), .ZN(n9229) );
  OAI21_X1 U5877 ( .B1(n7460), .B2(n5986), .A(n5985), .ZN(n7523) );
  NAND2_X1 U5878 ( .A1(n5680), .A2(n5679), .ZN(n9065) );
  INV_X1 U5879 ( .A(n7833), .ZN(n5453) );
  XOR2_X1 U5880 ( .A(n8745), .B(n4296), .Z(n4357) );
  INV_X1 U5881 ( .A(n8313), .ZN(n4532) );
  OR2_X1 U5882 ( .A1(n8047), .A2(n8046), .ZN(n4358) );
  INV_X1 U5883 ( .A(n8620), .ZN(n4396) );
  AND2_X1 U5884 ( .A1(n4314), .A2(n4976), .ZN(n5479) );
  NAND2_X1 U5885 ( .A1(n7410), .A2(n7817), .ZN(n7409) );
  AND2_X1 U5886 ( .A1(n5318), .A2(n4951), .ZN(n4359) );
  NAND2_X1 U5887 ( .A1(n7717), .A2(n7716), .ZN(n4360) );
  OR2_X1 U5888 ( .A1(n9180), .A2(n4580), .ZN(n4361) );
  NAND2_X1 U5889 ( .A1(n5307), .A2(n5306), .ZN(n8639) );
  NAND2_X1 U5890 ( .A1(n5670), .A2(n5669), .ZN(n9141) );
  INV_X1 U5891 ( .A(n7767), .ZN(n4823) );
  NAND2_X1 U5892 ( .A1(n5596), .A2(n5544), .ZN(n5601) );
  AND2_X1 U5893 ( .A1(n8319), .A2(n8320), .ZN(n9007) );
  AND2_X1 U5894 ( .A1(n6936), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n4362) );
  AND2_X1 U5895 ( .A1(n9286), .A2(n9295), .ZN(n4363) );
  AND2_X1 U5896 ( .A1(n9157), .A2(n9312), .ZN(n4364) );
  INV_X1 U5897 ( .A(n9015), .ZN(n9254) );
  NAND2_X1 U5898 ( .A1(n5686), .A2(n5685), .ZN(n9015) );
  AND2_X1 U5899 ( .A1(n8612), .A2(n8615), .ZN(n4365) );
  AND2_X1 U5900 ( .A1(n8043), .A2(n4491), .ZN(n4366) );
  OR2_X1 U5901 ( .A1(n8662), .A2(n8675), .ZN(n4367) );
  AND2_X1 U5902 ( .A1(n8131), .A2(n8054), .ZN(n4368) );
  AND2_X1 U5903 ( .A1(n6610), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n4369) );
  OR2_X1 U5904 ( .A1(n9460), .A2(n7641), .ZN(n8034) );
  INV_X1 U5905 ( .A(n6152), .ZN(n4762) );
  NAND2_X1 U5906 ( .A1(n8319), .A2(n8318), .ZN(n4370) );
  NAND2_X1 U5907 ( .A1(n8586), .A2(n8363), .ZN(n4644) );
  AND2_X1 U5908 ( .A1(n9847), .A2(n9904), .ZN(n4371) );
  INV_X1 U5909 ( .A(n8602), .ZN(n8751) );
  AND2_X1 U5910 ( .A1(n5321), .A2(n5320), .ZN(n8602) );
  NAND2_X1 U5911 ( .A1(n7676), .A2(n7677), .ZN(n4372) );
  AND2_X1 U5912 ( .A1(n4451), .A2(n8062), .ZN(n4373) );
  OR2_X1 U5913 ( .A1(n5356), .A2(n4729), .ZN(n4374) );
  INV_X1 U5914 ( .A(n4834), .ZN(n4832) );
  NAND2_X1 U5915 ( .A1(n7740), .A2(n7741), .ZN(n4834) );
  NAND2_X1 U5916 ( .A1(n8106), .A2(n8107), .ZN(n4375) );
  NAND2_X1 U5917 ( .A1(n5015), .A2(n5014), .ZN(n8757) );
  NAND2_X1 U5918 ( .A1(n5684), .A2(n5683), .ZN(n9021) );
  INV_X1 U5919 ( .A(n9021), .ZN(n4577) );
  NOR2_X1 U5920 ( .A1(n6218), .A2(n6217), .ZN(n4376) );
  NOR2_X1 U5921 ( .A1(n7553), .A2(n4804), .ZN(n4377) );
  NAND2_X1 U5922 ( .A1(n9320), .A2(n9169), .ZN(n4378) );
  AND2_X1 U5923 ( .A1(n8053), .A2(n9223), .ZN(n4379) );
  AND2_X1 U5924 ( .A1(n5382), .A2(n5381), .ZN(n8814) );
  INV_X1 U5925 ( .A(n5315), .ZN(n4400) );
  INV_X1 U5926 ( .A(n4848), .ZN(n4601) );
  NAND2_X1 U5927 ( .A1(n5643), .A2(n5642), .ZN(n9328) );
  INV_X1 U5928 ( .A(n9328), .ZN(n4583) );
  AND2_X1 U5929 ( .A1(n7169), .A2(n7302), .ZN(n7274) );
  NAND2_X1 U5930 ( .A1(n5453), .A2(n8539), .ZN(n6674) );
  OR2_X1 U5931 ( .A1(n4551), .A2(n6919), .ZN(n4380) );
  AND2_X1 U5932 ( .A1(n7658), .A2(n4585), .ZN(n4381) );
  NAND2_X1 U5933 ( .A1(n9845), .A2(n7875), .ZN(n7181) );
  NAND3_X1 U5934 ( .A1(n4330), .A2(n4787), .A3(n5596), .ZN(n4382) );
  NAND2_X1 U5935 ( .A1(n4664), .A2(n7270), .ZN(n7290) );
  NAND2_X1 U5936 ( .A1(n4976), .A2(n4975), .ZN(n5288) );
  OR2_X1 U5937 ( .A1(n7124), .A2(n7126), .ZN(n9858) );
  INV_X1 U5938 ( .A(n9858), .ZN(n4560) );
  AND2_X1 U5939 ( .A1(n5515), .A2(n5514), .ZN(n4383) );
  AND2_X1 U5940 ( .A1(n5355), .A2(SI_24_), .ZN(n4384) );
  INV_X1 U5941 ( .A(n9926), .ZN(n4559) );
  NAND2_X1 U5942 ( .A1(n5146), .A2(n5145), .ZN(n9857) );
  INV_X1 U5943 ( .A(n9857), .ZN(n4563) );
  INV_X1 U5944 ( .A(n7069), .ZN(n4806) );
  NAND2_X1 U5945 ( .A1(n6682), .A2(n7997), .ZN(n4385) );
  AND2_X1 U5946 ( .A1(n4299), .A2(n8206), .ZN(n4386) );
  OR2_X1 U5947 ( .A1(n7282), .A2(n9667), .ZN(n9624) );
  INV_X1 U5948 ( .A(n9624), .ZN(n4588) );
  AND2_X1 U5949 ( .A1(n7988), .A2(n7989), .ZN(n4387) );
  INV_X1 U5950 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n5573) );
  AND2_X1 U5951 ( .A1(n5555), .A2(n4496), .ZN(n9383) );
  NAND2_X1 U5952 ( .A1(n9477), .A2(n9478), .ZN(n4624) );
  INV_X1 U5953 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n4438) );
  INV_X1 U5954 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4750) );
  AOI21_X1 U5955 ( .B1(n8329), .B2(n9227), .A(n8328), .ZN(n9250) );
  INV_X1 U5956 ( .A(n7505), .ZN(n4403) );
  NOR2_X2 U5957 ( .A1(n4337), .A2(n4415), .ZN(n6903) );
  NAND2_X1 U5958 ( .A1(n4708), .A2(n4417), .ZN(n4707) );
  NAND2_X1 U5959 ( .A1(n4417), .A2(n5108), .ZN(n4712) );
  XNOR2_X1 U5960 ( .A(n4417), .B(n5108), .ZN(n6333) );
  AOI21_X1 U5961 ( .B1(n7992), .B2(n8810), .A(n4419), .ZN(n7995) );
  NAND2_X1 U5962 ( .A1(n4602), .A2(n4420), .ZN(n7991) );
  NAND3_X1 U5963 ( .A1(n4304), .A2(n4421), .A3(n7986), .ZN(n4420) );
  INV_X1 U5964 ( .A(n8502), .ZN(n4421) );
  NAND2_X1 U5965 ( .A1(n6992), .A2(n7792), .ZN(n4436) );
  INV_X2 U5966 ( .A(n5563), .ZN(n6327) );
  NAND2_X1 U5967 ( .A1(n5563), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n4437) );
  NAND4_X1 U5968 ( .A1(n4788), .A2(n5543), .A3(n4446), .A4(n4445), .ZN(n5586)
         );
  INV_X1 U5969 ( .A(n8063), .ZN(n4447) );
  AOI21_X1 U5970 ( .B1(n4447), .B2(n4450), .A(n4448), .ZN(n8061) );
  OR2_X1 U5971 ( .A1(n8079), .A2(n4461), .ZN(n4458) );
  NAND2_X1 U5972 ( .A1(n4458), .A2(n4459), .ZN(n8096) );
  INV_X1 U5973 ( .A(n8143), .ZN(n4470) );
  NAND2_X1 U5974 ( .A1(n4737), .A2(n4472), .ZN(n4471) );
  OAI211_X1 U5975 ( .C1(n4737), .C2(n4473), .A(n4476), .B(n4471), .ZN(P1_U3240) );
  INV_X1 U5976 ( .A(n8239), .ZN(n4478) );
  NAND3_X1 U5977 ( .A1(n4487), .A2(n4481), .A3(n4379), .ZN(n4480) );
  NAND2_X1 U5978 ( .A1(n5555), .A2(n4695), .ZN(n4696) );
  NAND2_X1 U5979 ( .A1(n4498), .A2(n7983), .ZN(n7999) );
  NAND2_X1 U5980 ( .A1(n4502), .A2(n4843), .ZN(n7953) );
  NAND2_X1 U5981 ( .A1(n4503), .A2(n7949), .ZN(n4502) );
  NAND2_X1 U5982 ( .A1(n4505), .A2(n4504), .ZN(n4503) );
  NAND3_X1 U5983 ( .A1(n4330), .A2(n4526), .A3(n5596), .ZN(n5729) );
  NOR2_X2 U5984 ( .A1(n5586), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n5596) );
  NAND2_X1 U5985 ( .A1(n9089), .A2(n4530), .ZN(n4527) );
  NAND2_X1 U5986 ( .A1(n4527), .A2(n4528), .ZN(n9044) );
  NAND2_X1 U5987 ( .A1(n8332), .A2(n4533), .ZN(P1_U3355) );
  AOI22_X1 U5988 ( .A1(n6261), .A2(n9660), .B1(n6257), .B2(n8957), .ZN(n5811)
         );
  OAI21_X1 U5989 ( .B1(n9197), .B2(n4537), .A(n4534), .ZN(n8307) );
  NAND2_X1 U5990 ( .A1(n7718), .A2(n4354), .ZN(n8296) );
  NAND2_X1 U5991 ( .A1(n7264), .A2(n4352), .ZN(n7265) );
  NAND2_X1 U5992 ( .A1(n8317), .A2(n4544), .ZN(n9026) );
  OAI21_X1 U5993 ( .B1(n8317), .B2(n4306), .A(n4541), .ZN(n8324) );
  AND2_X1 U5994 ( .A1(n8317), .A2(n8316), .ZN(n4854) );
  AND2_X2 U5995 ( .A1(n5050), .A2(n6327), .ZN(n5092) );
  NAND2_X1 U5996 ( .A1(n4550), .A2(n4549), .ZN(n7124) );
  OR3_X1 U5997 ( .A1(n8553), .A2(n4555), .A3(n8731), .ZN(n8495) );
  INV_X1 U5998 ( .A(n4554), .ZN(n5528) );
  NAND2_X1 U5999 ( .A1(n4560), .A2(n4313), .ZN(n9810) );
  NOR2_X1 U6000 ( .A1(n5719), .A2(n4567), .ZN(n4565) );
  NAND2_X1 U6001 ( .A1(n4573), .A2(n4567), .ZN(n4566) );
  INV_X1 U6002 ( .A(n5718), .ZN(n4568) );
  NAND2_X2 U6003 ( .A1(n5567), .A2(n5563), .ZN(n5665) );
  NAND2_X2 U6004 ( .A1(n5718), .A2(n5719), .ZN(n5567) );
  NAND3_X1 U6005 ( .A1(n4572), .A2(n4564), .A3(n4569), .ZN(n7038) );
  NAND2_X2 U6006 ( .A1(n5567), .A2(n6327), .ZN(n5600) );
  NAND2_X1 U6007 ( .A1(n5555), .A2(n4587), .ZN(n4586) );
  NAND2_X1 U6008 ( .A1(n4586), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5558) );
  NAND2_X1 U6009 ( .A1(n7845), .A2(n7805), .ZN(n6907) );
  NAND2_X1 U6010 ( .A1(n4596), .A2(n7854), .ZN(n4594) );
  INV_X1 U6011 ( .A(n7854), .ZN(n4595) );
  NAND2_X1 U6012 ( .A1(n4597), .A2(n4598), .ZN(n5439) );
  NAND2_X1 U6013 ( .A1(n9842), .A2(n7875), .ZN(n4597) );
  NAND2_X1 U6014 ( .A1(n7409), .A2(n4353), .ZN(n4600) );
  NAND2_X1 U6015 ( .A1(n8502), .A2(n4606), .ZN(n4604) );
  NAND2_X1 U6016 ( .A1(n8502), .A2(n8493), .ZN(n5452) );
  NOR2_X1 U6017 ( .A1(n9613), .A2(n7251), .ZN(n8011) );
  AOI21_X1 U6018 ( .B1(n8531), .B2(n8529), .A(n8530), .ZN(n8509) );
  NAND2_X1 U6019 ( .A1(n8544), .A2(n7822), .ZN(n8531) );
  INV_X2 U6020 ( .A(n6366), .ZN(n5070) );
  INV_X1 U6021 ( .A(n8710), .ZN(n8712) );
  NAND2_X1 U6022 ( .A1(n4626), .A2(n9959), .ZN(n4630) );
  NAND3_X1 U6023 ( .A1(n5049), .A2(n5061), .A3(n5048), .ZN(n4657) );
  NAND2_X1 U6024 ( .A1(n7268), .A2(n8116), .ZN(n4664) );
  INV_X1 U6025 ( .A(n4665), .ZN(n7652) );
  NAND2_X1 U6026 ( .A1(n8265), .A2(n4677), .ZN(n4675) );
  NAND2_X1 U6027 ( .A1(n4675), .A2(n4676), .ZN(n9138) );
  NAND2_X1 U6028 ( .A1(n7690), .A2(n4682), .ZN(n4681) );
  NAND2_X1 U6029 ( .A1(n8285), .A2(n4687), .ZN(n4689) );
  NAND2_X1 U6030 ( .A1(n8271), .A2(n4692), .ZN(n4690) );
  NAND2_X1 U6031 ( .A1(n4690), .A2(n4691), .ZN(n9088) );
  INV_X1 U6032 ( .A(n4698), .ZN(n5174) );
  NAND2_X1 U6033 ( .A1(n5330), .A2(n4960), .ZN(n4723) );
  OAI21_X1 U6034 ( .B1(n5330), .B2(n5329), .A(n4960), .ZN(n5338) );
  NAND3_X1 U6035 ( .A1(n4736), .A2(n8985), .A3(n4733), .ZN(n4732) );
  NAND2_X1 U6036 ( .A1(n5415), .A2(n5414), .ZN(n4740) );
  NAND2_X1 U6037 ( .A1(n9345), .A2(n8946), .ZN(n4745) );
  OAI21_X1 U6038 ( .B1(n7791), .B2(n4747), .A(n4744), .ZN(n4746) );
  INV_X1 U6039 ( .A(n4746), .ZN(n8092) );
  INV_X1 U6040 ( .A(n5697), .ZN(n4747) );
  NAND2_X1 U6041 ( .A1(n4857), .A2(n4750), .ZN(n4748) );
  NAND2_X1 U6042 ( .A1(n8926), .A2(n4762), .ZN(n4764) );
  NOR2_X1 U6043 ( .A1(n8926), .A2(n4762), .ZN(n4765) );
  INV_X1 U6044 ( .A(n6154), .ZN(n4766) );
  NAND3_X1 U6045 ( .A1(n4784), .A2(n4844), .A3(n6244), .ZN(P1_U3212) );
  NAND2_X1 U6046 ( .A1(n5596), .A2(n4787), .ZN(n5605) );
  NAND3_X1 U6047 ( .A1(n5542), .A2(n5541), .A3(n5543), .ZN(n5587) );
  NAND2_X1 U6048 ( .A1(n7667), .A2(n4796), .ZN(n4794) );
  NAND2_X1 U6049 ( .A1(n6788), .A2(n4797), .ZN(n7025) );
  NAND2_X1 U6050 ( .A1(n6788), .A2(n5843), .ZN(n5860) );
  OAI211_X2 U6051 ( .C1(n4801), .C2(n4800), .A(n4372), .B(n4798), .ZN(n7735)
         );
  NAND2_X1 U6052 ( .A1(n7553), .A2(n4799), .ZN(n4798) );
  NOR2_X2 U6053 ( .A1(n4804), .A2(n4802), .ZN(n4801) );
  AND2_X2 U6054 ( .A1(n7555), .A2(n7554), .ZN(n4804) );
  INV_X1 U6055 ( .A(n7556), .ZN(n4802) );
  INV_X1 U6056 ( .A(n7553), .ZN(n4803) );
  NAND2_X1 U6057 ( .A1(n8371), .A2(n4811), .ZN(n4809) );
  OAI211_X1 U6058 ( .C1(n8371), .C2(n4815), .A(n4812), .B(n4809), .ZN(n7774)
         );
  NAND2_X1 U6059 ( .A1(n8371), .A2(n4820), .ZN(n4817) );
  AOI21_X1 U6060 ( .B1(n8371), .B2(n8370), .A(n4810), .ZN(n8410) );
  OAI21_X2 U6061 ( .B1(n8349), .B2(n4829), .A(n4828), .ZN(n7745) );
  NAND2_X1 U6062 ( .A1(n7743), .A2(n7744), .ZN(n4833) );
  NAND2_X1 U6063 ( .A1(n6827), .A2(n4351), .ZN(n6836) );
  NAND2_X1 U6064 ( .A1(n6740), .A2(n6739), .ZN(n6827) );
  NAND2_X1 U6065 ( .A1(n4413), .A2(n4839), .ZN(n5003) );
  XNOR2_X1 U6066 ( .A(n5357), .B(n5353), .ZN(n7218) );
  NAND2_X1 U6067 ( .A1(n7274), .A2(n7393), .ZN(n7481) );
  XNOR2_X1 U6068 ( .A(n5689), .B(SI_30_), .ZN(n8840) );
  OAI21_X1 U6069 ( .B1(n7995), .B2(n7994), .A(n7993), .ZN(n7996) );
  OR2_X1 U6070 ( .A1(n5665), .A2(n4863), .ZN(n5575) );
  NAND2_X1 U6071 ( .A1(n5393), .A2(n5392), .ZN(n5395) );
  XNOR2_X1 U6072 ( .A(n5393), .B(n5392), .ZN(n7384) );
  INV_X1 U6073 ( .A(n6073), .ZN(n6076) );
  OR2_X1 U6074 ( .A1(n4290), .A2(n5802), .ZN(n5805) );
  OR2_X1 U6075 ( .A1(n4290), .A2(n5769), .ZN(n5775) );
  NAND2_X1 U6076 ( .A1(n5068), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5022) );
  NAND2_X1 U6077 ( .A1(n5068), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5044) );
  CLKBUF_X1 U6078 ( .A(n6977), .Z(n6891) );
  NAND2_X1 U6079 ( .A1(n6366), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5025) );
  INV_X2 U6080 ( .A(n5563), .ZN(n6326) );
  XNOR2_X1 U6081 ( .A(n5375), .B(n5374), .ZN(n7397) );
  AND2_X4 U6082 ( .A1(n5006), .A2(n7675), .ZN(n5068) );
  CLKBUF_X1 U6083 ( .A(n6733), .Z(n6691) );
  AND2_X1 U6084 ( .A1(n7745), .A2(n4357), .ZN(n7746) );
  OR3_X1 U6085 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .A3(
        P2_IR_REG_0__SCAN_IN), .ZN(n4840) );
  INV_X1 U6086 ( .A(n8428), .ZN(n8655) );
  INV_X1 U6087 ( .A(n8901), .ZN(n8944) );
  OR2_X1 U6088 ( .A1(n5533), .A2(n8777), .ZN(n4841) );
  NOR2_X1 U6089 ( .A1(n4607), .A2(n5508), .ZN(n4842) );
  AND2_X1 U6090 ( .A1(n8527), .A2(n7952), .ZN(n4843) );
  OR2_X1 U6091 ( .A1(n4577), .A2(n8910), .ZN(n4844) );
  OR2_X1 U6092 ( .A1(n8482), .A2(n8831), .ZN(n4845) );
  OR2_X1 U6093 ( .A1(n8482), .A2(n8777), .ZN(n4846) );
  OR2_X1 U6094 ( .A1(n5533), .A2(n8831), .ZN(n4847) );
  NOR2_X1 U6095 ( .A1(n5443), .A2(n7507), .ZN(n4848) );
  NOR2_X1 U6096 ( .A1(n7506), .A2(n5443), .ZN(n4849) );
  AND2_X1 U6097 ( .A1(n4898), .A2(n4897), .ZN(n4850) );
  AND2_X1 U6098 ( .A1(n4903), .A2(n4902), .ZN(n4851) );
  INV_X1 U6099 ( .A(n9342), .ZN(n5756) );
  INV_X1 U6100 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n4975) );
  NAND2_X1 U6101 ( .A1(n5796), .A2(n5795), .ZN(n6635) );
  AND2_X1 U6102 ( .A1(n4880), .A2(SI_5_), .ZN(n4853) );
  NAND2_X1 U6103 ( .A1(n9088), .A2(n8274), .ZN(n9054) );
  AND2_X1 U6104 ( .A1(n9250), .A2(n9249), .ZN(n4855) );
  OR2_X1 U6105 ( .A1(n7987), .A2(n7978), .ZN(n4856) );
  INV_X1 U6106 ( .A(n8322), .ZN(n8323) );
  INV_X1 U6107 ( .A(n7986), .ZN(n7970) );
  NAND2_X1 U6108 ( .A1(n7899), .A2(n7981), .ZN(n7900) );
  AND2_X1 U6109 ( .A1(n7906), .A2(n7905), .ZN(n7907) );
  AND2_X1 U6110 ( .A1(n8671), .A2(n7916), .ZN(n7917) );
  AOI21_X1 U6111 ( .B1(n7942), .B2(n7941), .A(n8566), .ZN(n7943) );
  OAI21_X1 U6112 ( .B1(n7986), .B2(n7981), .A(n4856), .ZN(n7971) );
  INV_X1 U6113 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5543) );
  INV_X1 U6114 ( .A(n7351), .ZN(n7352) );
  INV_X1 U6115 ( .A(n7971), .ZN(n7972) );
  INV_X1 U6116 ( .A(n5841), .ZN(n5842) );
  INV_X1 U6117 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5554) );
  INV_X1 U6118 ( .A(n5279), .ZN(n4992) );
  NAND2_X1 U6120 ( .A1(n5840), .A2(n5842), .ZN(n5843) );
  INV_X1 U6121 ( .A(n8116), .ZN(n7162) );
  INV_X1 U6122 ( .A(n5332), .ZN(n4995) );
  NOR2_X1 U6123 ( .A1(n7772), .A2(n8503), .ZN(n5509) );
  INV_X1 U6124 ( .A(n8731), .ZN(n5370) );
  NAND2_X1 U6125 ( .A1(n4992), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n5293) );
  INV_X1 U6126 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n9995) );
  NOR2_X1 U6127 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n4972) );
  NOR2_X1 U6128 ( .A1(n5976), .A2(n7535), .ZN(n5984) );
  NOR2_X1 U6129 ( .A1(n8241), .A2(n8995), .ZN(n8140) );
  NAND2_X1 U6130 ( .A1(n5845), .A2(n5816), .ZN(n5818) );
  NAND2_X1 U6131 ( .A1(n8325), .A2(n8946), .ZN(n8326) );
  INV_X1 U6132 ( .A(n6098), .ZN(n6096) );
  INV_X1 U6133 ( .A(n6030), .ZN(n6027) );
  INV_X1 U6134 ( .A(n5962), .ZN(n5929) );
  INV_X1 U6135 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5638) );
  OR2_X1 U6136 ( .A1(n5621), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n5624) );
  INV_X1 U6137 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5115) );
  NOR2_X1 U6138 ( .A1(n7749), .A2(n7748), .ZN(n7750) );
  OAI22_X1 U6139 ( .A1(n6722), .A2(n6721), .B1(n6689), .B2(n6688), .ZN(n6733)
         );
  INV_X1 U6140 ( .A(n5181), .ZN(n4989) );
  NAND2_X1 U6141 ( .A1(n6673), .A2(n6682), .ZN(n6680) );
  NAND2_X1 U6142 ( .A1(n8639), .A2(n8428), .ZN(n5316) );
  NAND2_X1 U6143 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5080) );
  OR2_X1 U6144 ( .A1(n5050), .A2(n5031), .ZN(n5032) );
  OR4_X1 U6145 ( .A1(n5188), .A2(P2_IR_REG_11__SCAN_IN), .A3(
        P2_IR_REG_10__SCAN_IN), .A4(P2_IR_REG_9__SCAN_IN), .ZN(n5260) );
  XNOR2_X1 U6146 ( .A(n5971), .B(n4298), .ZN(n5977) );
  INV_X1 U6147 ( .A(n8883), .ZN(n6046) );
  OR2_X1 U6148 ( .A1(n6158), .A2(n6157), .ZN(n6176) );
  NAND2_X1 U6149 ( .A1(n5930), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5988) );
  OR2_X1 U6150 ( .A1(n5799), .A2(n6305), .ZN(n5787) );
  INV_X1 U6151 ( .A(n8995), .ZN(n5698) );
  OR2_X1 U6152 ( .A1(n6115), .A2(n8866), .ZN(n6132) );
  OR2_X1 U6153 ( .A1(n9141), .A2(n9123), .ZN(n8268) );
  NAND2_X1 U6154 ( .A1(n6048), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n6080) );
  OR2_X1 U6155 ( .A1(n5988), .A2(n5987), .ZN(n6002) );
  INV_X1 U6156 ( .A(n8112), .ZN(n7149) );
  INV_X1 U6157 ( .A(n5273), .ZN(n4938) );
  NAND2_X1 U6158 ( .A1(n4900), .A2(n4899), .ZN(n4903) );
  INV_X1 U6159 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n4868) );
  NAND2_X1 U6160 ( .A1(n4989), .A2(n4988), .ZN(n5192) );
  AND2_X1 U6161 ( .A1(n6426), .A2(n6407), .ZN(n6535) );
  NAND2_X1 U6162 ( .A1(n7944), .A2(n7945), .ZN(n8566) );
  OR2_X1 U6163 ( .A1(n8668), .A2(n8430), .ZN(n5285) );
  OR2_X1 U6164 ( .A1(n6682), .A2(n8682), .ZN(n6663) );
  INV_X1 U6165 ( .A(n8715), .ZN(n8711) );
  AND2_X1 U6166 ( .A1(n6789), .A2(n6787), .ZN(n5839) );
  INV_X1 U6167 ( .A(n8907), .ZN(n8940) );
  AND2_X1 U6168 ( .A1(n8995), .A2(n8097), .ZN(n8239) );
  NAND2_X1 U6169 ( .A1(n5803), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5804) );
  OR2_X1 U6170 ( .A1(n9580), .A2(n9579), .ZN(n9582) );
  XNOR2_X1 U6171 ( .A(n8997), .B(n5698), .ZN(n5708) );
  INV_X1 U6172 ( .A(n8311), .ZN(n9090) );
  AND2_X1 U6173 ( .A1(n8156), .A2(n8016), .ZN(n8117) );
  INV_X1 U6174 ( .A(n9629), .ZN(n9239) );
  AND2_X1 U6175 ( .A1(n5753), .A2(n9382), .ZN(n6232) );
  NAND2_X1 U6176 ( .A1(n7652), .A2(n7651), .ZN(n7654) );
  INV_X1 U6177 ( .A(n7468), .ZN(n7393) );
  INV_X1 U6178 ( .A(n9686), .ZN(n9705) );
  AND2_X1 U6179 ( .A1(n7045), .A2(n7044), .ZN(n9610) );
  AND2_X1 U6180 ( .A1(n4933), .A2(n4932), .ZN(n5254) );
  NAND2_X1 U6181 ( .A1(n4893), .A2(n4892), .ZN(n5138) );
  OR3_X1 U6182 ( .A1(n9870), .A2(n9869), .A3(n7400), .ZN(n6665) );
  INV_X1 U6183 ( .A(n8819), .ZN(n8346) );
  AND2_X1 U6184 ( .A1(n5384), .A2(n5365), .ZN(n8537) );
  INV_X1 U6185 ( .A(n8417), .ZN(n8364) );
  AND3_X1 U6186 ( .A1(n5327), .A2(n5326), .A3(n5325), .ZN(n8617) );
  AND4_X1 U6187 ( .A1(n5284), .A2(n5283), .A3(n5282), .A4(n5281), .ZN(n8654)
         );
  AND2_X1 U6188 ( .A1(n6395), .A2(n6394), .ZN(n9783) );
  INV_X1 U6189 ( .A(n8501), .ZN(n8493) );
  AND2_X1 U6190 ( .A1(n8633), .A2(n7924), .ZN(n8651) );
  INV_X1 U6191 ( .A(n8556), .ZN(n9854) );
  INV_X1 U6192 ( .A(n9866), .ZN(n8579) );
  AOI21_X1 U6193 ( .B1(n8712), .B2(n7321), .A(n8711), .ZN(n8804) );
  INV_X1 U6194 ( .A(n5489), .ZN(n9867) );
  NAND2_X1 U6195 ( .A1(n6665), .A2(n5495), .ZN(n9868) );
  INV_X1 U6196 ( .A(n9599), .ZN(n9567) );
  AND2_X1 U6197 ( .A1(n8049), .A2(n8008), .ZN(n8127) );
  AND2_X1 U6198 ( .A1(n7037), .A2(n9654), .ZN(n9646) );
  INV_X1 U6199 ( .A(n9379), .ZN(n5766) );
  OR2_X1 U6200 ( .A1(n9252), .A2(n9699), .ZN(n9258) );
  AND2_X1 U6201 ( .A1(n9610), .A2(n9712), .ZN(n9699) );
  INV_X1 U6202 ( .A(n9699), .ZN(n9710) );
  OR2_X1 U6203 ( .A1(n7056), .A2(n7037), .ZN(n6234) );
  AND2_X1 U6204 ( .A1(n5626), .A2(n5625), .ZN(n6936) );
  XNOR2_X1 U6205 ( .A(n4879), .B(SI_5_), .ZN(n5090) );
  INV_X1 U6206 ( .A(n8464), .ZN(n9781) );
  INV_X1 U6207 ( .A(n8420), .ZN(n8360) );
  NAND2_X1 U6208 ( .A1(n6694), .A2(n6693), .ZN(n8422) );
  AOI21_X1 U6209 ( .B1(n8498), .B2(n5347), .A(n5407), .ZN(n8412) );
  INV_X1 U6210 ( .A(n7607), .ZN(n8432) );
  INV_X1 U6211 ( .A(n8579), .ZN(n9855) );
  INV_X1 U6212 ( .A(n9834), .ZN(n8709) );
  INV_X1 U6213 ( .A(n9959), .ZN(n9956) );
  INV_X1 U6214 ( .A(n9874), .ZN(n9989) );
  INV_X1 U6215 ( .A(n7829), .ZN(n7983) );
  INV_X1 U6216 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n10004) );
  INV_X1 U6217 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6324) );
  OR2_X1 U6218 ( .A1(n6281), .A2(n6280), .ZN(n6282) );
  INV_X1 U6219 ( .A(n6253), .ZN(n6254) );
  OR2_X1 U6220 ( .A1(n6316), .A2(n6315), .ZN(n9605) );
  OR2_X1 U6221 ( .A1(P1_U3083), .A2(n6320), .ZN(n9609) );
  OR2_X1 U6224 ( .A1(n6234), .A2(n5754), .ZN(n9731) );
  INV_X1 U6225 ( .A(n9065), .ZN(n9354) );
  AND4_X1 U6226 ( .A1(n9692), .A2(n9691), .A3(n9690), .A4(n9689), .ZN(n9728)
         );
  INV_X1 U6227 ( .A(n9650), .ZN(n9651) );
  INV_X1 U6228 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6372) );
  AND2_X1 U6229 ( .A1(n6377), .A2(n9871), .ZN(P2_U3966) );
  AND2_X1 U6230 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n4858) );
  NAND2_X1 U6231 ( .A1(n4873), .A2(n4858), .ZN(n5570) );
  AND2_X1 U6232 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n4859) );
  NAND2_X1 U6233 ( .A1(n5563), .A2(n4859), .ZN(n5039) );
  INV_X1 U6234 ( .A(SI_1_), .ZN(n4860) );
  MUX2_X1 U6235 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n4873), .Z(n5027) );
  NAND2_X1 U6236 ( .A1(n4861), .A2(SI_1_), .ZN(n4862) );
  INV_X1 U6237 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n4864) );
  INV_X1 U6238 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n4863) );
  MUX2_X1 U6239 ( .A(n4864), .B(n4863), .S(n4873), .Z(n4865) );
  XNOR2_X1 U6240 ( .A(n4865), .B(SI_2_), .ZN(n5048) );
  INV_X1 U6241 ( .A(n4865), .ZN(n4866) );
  NAND2_X1 U6242 ( .A1(n4866), .A2(SI_2_), .ZN(n4867) );
  INV_X1 U6243 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n4869) );
  MUX2_X1 U6244 ( .A(n4869), .B(n4868), .S(n4873), .Z(n4870) );
  XNOR2_X1 U6245 ( .A(n4870), .B(SI_3_), .ZN(n5061) );
  INV_X1 U6246 ( .A(n4870), .ZN(n4871) );
  INV_X1 U6247 ( .A(n5563), .ZN(n4872) );
  MUX2_X1 U6248 ( .A(n6324), .B(n6330), .S(n4872), .Z(n4876) );
  XNOR2_X1 U6249 ( .A(n4876), .B(SI_4_), .ZN(n5086) );
  INV_X1 U6250 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6325) );
  INV_X1 U6251 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n4874) );
  MUX2_X1 U6252 ( .A(n6325), .B(n4874), .S(n4873), .Z(n4879) );
  NAND2_X1 U6253 ( .A1(n5087), .A2(n4875), .ZN(n4883) );
  INV_X1 U6254 ( .A(n4876), .ZN(n4877) );
  NAND2_X1 U6255 ( .A1(n4877), .A2(SI_4_), .ZN(n5088) );
  INV_X1 U6256 ( .A(n5088), .ZN(n4878) );
  INV_X1 U6257 ( .A(n4879), .ZN(n4880) );
  INV_X1 U6258 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6334) );
  INV_X1 U6259 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6332) );
  MUX2_X1 U6260 ( .A(n6334), .B(n6332), .S(n6326), .Z(n4884) );
  INV_X1 U6261 ( .A(n4884), .ZN(n4885) );
  NAND2_X1 U6262 ( .A1(n4885), .A2(SI_6_), .ZN(n4886) );
  INV_X1 U6263 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6351) );
  INV_X1 U6264 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6354) );
  MUX2_X1 U6265 ( .A(n6351), .B(n6354), .S(n6327), .Z(n4890) );
  INV_X1 U6266 ( .A(SI_8_), .ZN(n4889) );
  INV_X1 U6267 ( .A(n4890), .ZN(n4891) );
  NAND2_X1 U6268 ( .A1(n4891), .A2(SI_8_), .ZN(n4892) );
  INV_X1 U6269 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6358) );
  MUX2_X1 U6270 ( .A(n6358), .B(n6361), .S(n6327), .Z(n4895) );
  INV_X1 U6271 ( .A(SI_9_), .ZN(n4894) );
  INV_X1 U6272 ( .A(n4895), .ZN(n4896) );
  NAND2_X1 U6273 ( .A1(n4896), .A2(SI_9_), .ZN(n4897) );
  MUX2_X1 U6274 ( .A(n10004), .B(n6363), .S(n6327), .Z(n4900) );
  INV_X1 U6275 ( .A(SI_10_), .ZN(n4899) );
  INV_X1 U6276 ( .A(n4900), .ZN(n4901) );
  NAND2_X1 U6277 ( .A1(n4901), .A2(SI_10_), .ZN(n4902) );
  INV_X1 U6278 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6374) );
  MUX2_X1 U6279 ( .A(n6374), .B(n6372), .S(n6327), .Z(n4904) );
  INV_X1 U6280 ( .A(n4904), .ZN(n4905) );
  INV_X1 U6281 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6425) );
  INV_X1 U6282 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6423) );
  MUX2_X1 U6283 ( .A(n6425), .B(n6423), .S(n6327), .Z(n4909) );
  INV_X1 U6284 ( .A(SI_12_), .ZN(n4908) );
  NAND2_X1 U6285 ( .A1(n4909), .A2(n4908), .ZN(n5205) );
  INV_X1 U6286 ( .A(n4909), .ZN(n4910) );
  NAND2_X1 U6287 ( .A1(n4910), .A2(SI_12_), .ZN(n4911) );
  NAND2_X1 U6288 ( .A1(n5205), .A2(n4911), .ZN(n5203) );
  INV_X1 U6289 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6488) );
  INV_X1 U6290 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n6486) );
  MUX2_X1 U6291 ( .A(n6488), .B(n6486), .S(n6327), .Z(n4915) );
  INV_X1 U6292 ( .A(n4915), .ZN(n4912) );
  INV_X1 U6293 ( .A(SI_13_), .ZN(n4914) );
  NAND2_X1 U6294 ( .A1(n4915), .A2(n4914), .ZN(n5208) );
  AND2_X1 U6295 ( .A1(n5205), .A2(n5208), .ZN(n4916) );
  INV_X1 U6296 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6482) );
  INV_X1 U6297 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n6484) );
  MUX2_X1 U6298 ( .A(n6482), .B(n6484), .S(n6326), .Z(n4919) );
  XNOR2_X1 U6299 ( .A(n4919), .B(SI_14_), .ZN(n5225) );
  INV_X1 U6300 ( .A(n4919), .ZN(n4920) );
  INV_X1 U6301 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6554) );
  INV_X1 U6302 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6556) );
  MUX2_X1 U6303 ( .A(n6554), .B(n6556), .S(n6327), .Z(n4924) );
  INV_X1 U6304 ( .A(SI_15_), .ZN(n4923) );
  INV_X1 U6305 ( .A(n4924), .ZN(n4925) );
  NAND2_X1 U6306 ( .A1(n4925), .A2(SI_15_), .ZN(n4926) );
  INV_X1 U6307 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n6600) );
  INV_X1 U6308 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n4928) );
  MUX2_X1 U6309 ( .A(n6600), .B(n4928), .S(n6326), .Z(n4930) );
  INV_X1 U6310 ( .A(SI_16_), .ZN(n4929) );
  NAND2_X1 U6311 ( .A1(n4930), .A2(n4929), .ZN(n4933) );
  INV_X1 U6312 ( .A(n4930), .ZN(n4931) );
  NAND2_X1 U6313 ( .A1(n4931), .A2(SI_16_), .ZN(n4932) );
  INV_X1 U6314 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n6632) );
  INV_X1 U6315 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n4934) );
  MUX2_X1 U6316 ( .A(n6632), .B(n4934), .S(n6326), .Z(n4935) );
  INV_X1 U6317 ( .A(n4935), .ZN(n4936) );
  NAND2_X1 U6318 ( .A1(n4936), .A2(SI_17_), .ZN(n4937) );
  MUX2_X1 U6319 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n6327), .Z(n4940) );
  XNOR2_X1 U6320 ( .A(n4940), .B(SI_18_), .ZN(n5286) );
  INV_X1 U6321 ( .A(n5286), .ZN(n4939) );
  NAND2_X1 U6322 ( .A1(n4940), .A2(SI_18_), .ZN(n4941) );
  INV_X1 U6323 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n6780) );
  INV_X1 U6324 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n6782) );
  MUX2_X1 U6325 ( .A(n6780), .B(n6782), .S(n6326), .Z(n4943) );
  INV_X1 U6326 ( .A(SI_19_), .ZN(n4942) );
  NAND2_X1 U6327 ( .A1(n4943), .A2(n4942), .ZN(n4946) );
  INV_X1 U6328 ( .A(n4943), .ZN(n4944) );
  NAND2_X1 U6329 ( .A1(n4944), .A2(SI_19_), .ZN(n4945) );
  NAND2_X1 U6330 ( .A1(n4946), .A2(n4945), .ZN(n5300) );
  INV_X1 U6331 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n6873) );
  INV_X1 U6332 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n6871) );
  MUX2_X1 U6333 ( .A(n6873), .B(n6871), .S(n6326), .Z(n4948) );
  INV_X1 U6334 ( .A(SI_20_), .ZN(n4947) );
  NAND2_X1 U6335 ( .A1(n4948), .A2(n4947), .ZN(n4951) );
  INV_X1 U6336 ( .A(n4948), .ZN(n4949) );
  NAND2_X1 U6337 ( .A1(n4949), .A2(SI_20_), .ZN(n4950) );
  INV_X1 U6338 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n10082) );
  INV_X1 U6339 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n6945) );
  MUX2_X1 U6340 ( .A(n10082), .B(n6945), .S(n6327), .Z(n4952) );
  XNOR2_X1 U6341 ( .A(n4952), .B(SI_21_), .ZN(n5318) );
  INV_X1 U6342 ( .A(n4952), .ZN(n4953) );
  NAND2_X1 U6343 ( .A1(n4953), .A2(SI_21_), .ZN(n4954) );
  INV_X1 U6344 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n6995) );
  INV_X1 U6345 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n6993) );
  MUX2_X1 U6346 ( .A(n6995), .B(n6993), .S(n6326), .Z(n4957) );
  INV_X1 U6347 ( .A(SI_22_), .ZN(n4956) );
  NAND2_X1 U6348 ( .A1(n4957), .A2(n4956), .ZN(n4960) );
  INV_X1 U6349 ( .A(n4957), .ZN(n4958) );
  NAND2_X1 U6350 ( .A1(n4958), .A2(SI_22_), .ZN(n4959) );
  NAND2_X1 U6351 ( .A1(n4960), .A2(n4959), .ZN(n5329) );
  INV_X1 U6352 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n4962) );
  INV_X1 U6353 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n4961) );
  MUX2_X1 U6354 ( .A(n4962), .B(n4961), .S(n6326), .Z(n4964) );
  INV_X1 U6355 ( .A(SI_23_), .ZN(n4963) );
  NAND2_X1 U6356 ( .A1(n4964), .A2(n4963), .ZN(n4967) );
  INV_X1 U6357 ( .A(n4964), .ZN(n4965) );
  NAND2_X1 U6358 ( .A1(n4965), .A2(SI_23_), .ZN(n4966) );
  INV_X1 U6359 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7219) );
  INV_X1 U6360 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7220) );
  MUX2_X1 U6361 ( .A(n7219), .B(n7220), .S(n6327), .Z(n5354) );
  XNOR2_X1 U6362 ( .A(n5354), .B(SI_24_), .ZN(n5353) );
  NAND3_X1 U6363 ( .A1(n4974), .A2(n4973), .A3(n5094), .ZN(n5262) );
  INV_X1 U6364 ( .A(n5262), .ZN(n4976) );
  NOR2_X1 U6365 ( .A1(P2_IR_REG_24__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .ZN(
        n4977) );
  INV_X1 U6366 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n4978) );
  NAND2_X1 U6367 ( .A1(n4983), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4979) );
  INV_X1 U6368 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n4980) );
  INV_X1 U6369 ( .A(n5000), .ZN(n4981) );
  NAND2_X1 U6370 ( .A1(n7218), .A2(n7792), .ZN(n4985) );
  NAND2_X1 U6371 ( .A1(n5092), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n4984) );
  INV_X1 U6372 ( .A(n5080), .ZN(n4986) );
  NAND2_X1 U6373 ( .A1(n4986), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5102) );
  INV_X1 U6374 ( .A(n5102), .ZN(n4987) );
  INV_X1 U6375 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5153) );
  AND2_X1 U6376 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_REG3_REG_11__SCAN_IN), 
        .ZN(n4988) );
  INV_X1 U6377 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n10078) );
  INV_X1 U6378 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n10091) );
  INV_X1 U6379 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n7558) );
  INV_X1 U6380 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n8354) );
  INV_X1 U6381 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n8393) );
  INV_X1 U6382 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n5343) );
  INV_X1 U6383 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n8386) );
  NAND2_X1 U6384 ( .A1(n5346), .A2(n8386), .ZN(n4997) );
  NAND2_X1 U6385 ( .A1(n5364), .A2(n4997), .ZN(n8557) );
  INV_X1 U6386 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5001) );
  INV_X1 U6387 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n4999) );
  OR2_X1 U6388 ( .A1(n8557), .A2(n5423), .ZN(n5011) );
  INV_X1 U6389 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n8558) );
  AND2_X4 U6390 ( .A1(n8842), .A2(n7675), .ZN(n6366) );
  NAND2_X1 U6391 ( .A1(n5068), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n5008) );
  NAND2_X1 U6392 ( .A1(n5078), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n5007) );
  OAI211_X1 U6393 ( .C1(n8558), .C2(n5070), .A(n5008), .B(n5007), .ZN(n5009)
         );
  INV_X1 U6394 ( .A(n5009), .ZN(n5010) );
  INV_X1 U6395 ( .A(n8372), .ZN(n8425) );
  XNOR2_X1 U6396 ( .A(n5013), .B(n5012), .ZN(n6870) );
  NAND2_X1 U6397 ( .A1(n6870), .A2(n7792), .ZN(n5015) );
  NAND2_X1 U6398 ( .A1(n5092), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n5014) );
  INV_X1 U6399 ( .A(n8757), .ZN(n8626) );
  NAND2_X1 U6400 ( .A1(n5310), .A2(n8393), .ZN(n5016) );
  NAND2_X1 U6401 ( .A1(n5323), .A2(n5016), .ZN(n8394) );
  INV_X1 U6402 ( .A(n8394), .ZN(n8624) );
  NAND2_X1 U6403 ( .A1(n8624), .A2(n5347), .ZN(n5021) );
  NAND2_X1 U6404 ( .A1(n5068), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n5018) );
  NAND2_X1 U6405 ( .A1(n5078), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n5017) );
  AND2_X1 U6406 ( .A1(n5018), .A2(n5017), .ZN(n5020) );
  NAND2_X1 U6407 ( .A1(n6366), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n5019) );
  NAND2_X1 U6408 ( .A1(n4294), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5023) );
  NAND2_X1 U6409 ( .A1(n4291), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n5024) );
  NAND3_X2 U6410 ( .A1(n5026), .A2(n5025), .A3(n5024), .ZN(n6673) );
  XNOR2_X1 U6411 ( .A(n5028), .B(n5027), .ZN(n6344) );
  NAND2_X1 U6412 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5030) );
  XNOR2_X1 U6413 ( .A(n5030), .B(P2_IR_REG_1__SCAN_IN), .ZN(n6443) );
  INV_X1 U6414 ( .A(n6443), .ZN(n5031) );
  NAND2_X1 U6415 ( .A1(n6366), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5036) );
  NAND2_X1 U6416 ( .A1(n4292), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n5035) );
  NAND2_X1 U6417 ( .A1(n5068), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5034) );
  NAND2_X1 U6418 ( .A1(n5078), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5033) );
  NAND2_X1 U6419 ( .A1(n5563), .A2(SI_0_), .ZN(n5038) );
  INV_X1 U6420 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5037) );
  NAND2_X1 U6421 ( .A1(n5038), .A2(n5037), .ZN(n5040) );
  AND2_X1 U6422 ( .A1(n5040), .A2(n5039), .ZN(n8845) );
  MUX2_X1 U6423 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8845), .S(n5050), .Z(n6972) );
  NAND2_X1 U6424 ( .A1(n6701), .A2(n6972), .ZN(n6700) );
  NAND2_X1 U6425 ( .A1(n7803), .A2(n6700), .ZN(n6699) );
  NAND2_X1 U6426 ( .A1(n6699), .A2(n7102), .ZN(n5043) );
  INV_X1 U6427 ( .A(n6700), .ZN(n5041) );
  NAND2_X1 U6428 ( .A1(n5041), .A2(n6673), .ZN(n5042) );
  NAND2_X1 U6429 ( .A1(n5043), .A2(n5042), .ZN(n6925) );
  NAND2_X1 U6430 ( .A1(n5078), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5047) );
  NAND2_X1 U6431 ( .A1(n4292), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n5046) );
  NAND2_X1 U6432 ( .A1(n6366), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5045) );
  NAND2_X1 U6433 ( .A1(n5092), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n5055) );
  XNOR2_X1 U6434 ( .A(n5049), .B(n5048), .ZN(n6338) );
  OR2_X1 U6435 ( .A1(n5051), .A2(n4999), .ZN(n5052) );
  XNOR2_X1 U6436 ( .A(n5052), .B(P2_IR_REG_2__SCAN_IN), .ZN(n9437) );
  NAND2_X1 U6437 ( .A1(n5305), .A2(n9437), .ZN(n5053) );
  NAND2_X1 U6438 ( .A1(n6687), .A2(n9887), .ZN(n7856) );
  INV_X1 U6439 ( .A(n9887), .ZN(n6924) );
  NAND2_X1 U6440 ( .A1(n5078), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5060) );
  INV_X1 U6441 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n5056) );
  NAND2_X1 U6442 ( .A1(n4292), .A2(n5056), .ZN(n5059) );
  NAND2_X1 U6443 ( .A1(n6366), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5058) );
  NAND2_X1 U6444 ( .A1(n5068), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5057) );
  NAND4_X1 U6445 ( .A1(n5060), .A2(n5059), .A3(n5058), .A4(n5057), .ZN(n8443)
         );
  NAND2_X1 U6446 ( .A1(n5092), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n5066) );
  XNOR2_X1 U6447 ( .A(n5062), .B(n5061), .ZN(n6340) );
  OR2_X1 U6448 ( .A1(n5029), .A2(n6340), .ZN(n5065) );
  NAND2_X1 U6449 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n4840), .ZN(n5063) );
  XNOR2_X1 U6450 ( .A(n5063), .B(P2_IR_REG_3__SCAN_IN), .ZN(n9744) );
  NAND2_X1 U6451 ( .A1(n5305), .A2(n9744), .ZN(n5064) );
  NAND2_X1 U6452 ( .A1(n8443), .A2(n7225), .ZN(n7858) );
  NAND2_X1 U6453 ( .A1(n6765), .A2(n6770), .ZN(n6767) );
  INV_X1 U6454 ( .A(n8443), .ZN(n6950) );
  NAND2_X1 U6455 ( .A1(n6950), .A2(n7225), .ZN(n5067) );
  NAND2_X1 U6456 ( .A1(n6767), .A2(n5067), .ZN(n6947) );
  NAND2_X1 U6457 ( .A1(n5068), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5074) );
  NAND2_X1 U6458 ( .A1(n4293), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5073) );
  OAI21_X1 U6459 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(P2_REG3_REG_4__SCAN_IN), 
        .A(n5080), .ZN(n6958) );
  INV_X1 U6460 ( .A(n6958), .ZN(n5069) );
  NAND2_X1 U6461 ( .A1(n4291), .A2(n5069), .ZN(n5072) );
  INV_X1 U6462 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6953) );
  OR2_X1 U6463 ( .A1(n5070), .A2(n6953), .ZN(n5071) );
  OR2_X1 U6464 ( .A1(n5094), .A2(n4999), .ZN(n5075) );
  XNOR2_X1 U6465 ( .A(n5075), .B(P2_IR_REG_4__SCAN_IN), .ZN(n6427) );
  NAND2_X1 U6466 ( .A1(n5305), .A2(n6427), .ZN(n5077) );
  XNOR2_X1 U6467 ( .A(n5087), .B(n5086), .ZN(n6329) );
  OR2_X1 U6468 ( .A1(n5029), .A2(n6329), .ZN(n5076) );
  OAI211_X2 U6469 ( .C1(n5109), .C2(n6324), .A(n5077), .B(n5076), .ZN(n6960)
         );
  NAND2_X1 U6470 ( .A1(n6865), .A2(n6960), .ZN(n7839) );
  INV_X1 U6471 ( .A(n6960), .ZN(n9891) );
  NAND2_X1 U6472 ( .A1(n6947), .A2(n7807), .ZN(n6946) );
  NAND2_X1 U6473 ( .A1(n6865), .A2(n9891), .ZN(n6846) );
  NAND2_X1 U6474 ( .A1(n5068), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5085) );
  NAND2_X1 U6475 ( .A1(n5078), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5084) );
  INV_X1 U6476 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5079) );
  NAND2_X1 U6477 ( .A1(n5080), .A2(n5079), .ZN(n5081) );
  AND2_X1 U6478 ( .A1(n5102), .A2(n5081), .ZN(n7210) );
  NAND2_X1 U6479 ( .A1(n4292), .A2(n7210), .ZN(n5083) );
  NAND2_X1 U6480 ( .A1(n6366), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5082) );
  NAND4_X1 U6481 ( .A1(n5085), .A2(n5084), .A3(n5083), .A4(n5082), .ZN(n8441)
         );
  NAND2_X1 U6482 ( .A1(n5087), .A2(n5086), .ZN(n5089) );
  NAND2_X1 U6483 ( .A1(n5089), .A2(n5088), .ZN(n5091) );
  XNOR2_X1 U6484 ( .A(n5091), .B(n5090), .ZN(n6343) );
  NAND2_X1 U6485 ( .A1(n5092), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n5096) );
  INV_X1 U6486 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5093) );
  NAND2_X1 U6487 ( .A1(n5094), .A2(n5093), .ZN(n5143) );
  NAND2_X1 U6488 ( .A1(n5143), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5110) );
  XNOR2_X1 U6489 ( .A(n5110), .B(P2_IR_REG_5__SCAN_IN), .ZN(n6551) );
  NAND2_X1 U6490 ( .A1(n5305), .A2(n6551), .ZN(n5095) );
  OR2_X1 U6491 ( .A1(n8441), .A2(n6828), .ZN(n5097) );
  AND2_X1 U6492 ( .A1(n6846), .A2(n5097), .ZN(n5098) );
  NAND2_X1 U6493 ( .A1(n6946), .A2(n5098), .ZN(n5100) );
  NAND2_X1 U6494 ( .A1(n6951), .A2(n6828), .ZN(n7834) );
  NAND2_X1 U6495 ( .A1(n8441), .A2(n7212), .ZN(n7860) );
  NAND2_X1 U6496 ( .A1(n7834), .A2(n7860), .ZN(n7808) );
  OR2_X1 U6497 ( .A1(n7808), .A2(n7212), .ZN(n5099) );
  NAND2_X1 U6498 ( .A1(n5100), .A2(n5099), .ZN(n7775) );
  NAND2_X1 U6499 ( .A1(n5078), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5107) );
  NAND2_X1 U6500 ( .A1(n6366), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5106) );
  INV_X1 U6501 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n5101) );
  NAND2_X1 U6502 ( .A1(n5102), .A2(n5101), .ZN(n5103) );
  AND2_X1 U6503 ( .A1(n5116), .A2(n5103), .ZN(n6839) );
  NAND2_X1 U6504 ( .A1(n4291), .A2(n6839), .ZN(n5105) );
  NAND2_X1 U6505 ( .A1(n5068), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5104) );
  NAND4_X1 U6506 ( .A1(n5107), .A2(n5106), .A3(n5105), .A4(n5104), .ZN(n8440)
         );
  NAND2_X1 U6507 ( .A1(n7788), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n5113) );
  INV_X1 U6508 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5140) );
  NAND2_X1 U6509 ( .A1(n5110), .A2(n5140), .ZN(n5111) );
  NAND2_X1 U6510 ( .A1(n5111), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5124) );
  XNOR2_X1 U6511 ( .A(n5124), .B(P2_IR_REG_6__SCAN_IN), .ZN(n6413) );
  NAND2_X1 U6512 ( .A1(n5305), .A2(n6413), .ZN(n5112) );
  AND2_X1 U6513 ( .A1(n8440), .A2(n9897), .ZN(n5114) );
  NAND2_X1 U6514 ( .A1(n5068), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5122) );
  NAND2_X1 U6515 ( .A1(n4293), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5121) );
  NAND2_X1 U6516 ( .A1(n5116), .A2(n5115), .ZN(n5117) );
  AND2_X1 U6517 ( .A1(n5132), .A2(n5117), .ZN(n7125) );
  NAND2_X1 U6518 ( .A1(n4292), .A2(n7125), .ZN(n5120) );
  INV_X1 U6519 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n5118) );
  OR2_X1 U6520 ( .A1(n5070), .A2(n5118), .ZN(n5119) );
  INV_X1 U6521 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5123) );
  NAND2_X1 U6522 ( .A1(n5124), .A2(n5123), .ZN(n5125) );
  NAND2_X1 U6523 ( .A1(n5125), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5126) );
  XNOR2_X1 U6524 ( .A(n5126), .B(P2_IR_REG_7__SCAN_IN), .ZN(n9757) );
  INV_X1 U6525 ( .A(n9757), .ZN(n6347) );
  XNOR2_X1 U6526 ( .A(n5128), .B(n5127), .ZN(n5595) );
  NAND2_X1 U6527 ( .A1(n5595), .A2(n7792), .ZN(n5130) );
  NAND2_X1 U6528 ( .A1(n7788), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n5129) );
  OAI211_X1 U6529 ( .C1(n5050), .C2(n6347), .A(n5130), .B(n5129), .ZN(n7126)
         );
  NAND2_X1 U6530 ( .A1(n9847), .A2(n7126), .ZN(n7872) );
  INV_X1 U6531 ( .A(n9847), .ZN(n8439) );
  INV_X1 U6532 ( .A(n7126), .ZN(n9904) );
  NAND2_X1 U6533 ( .A1(n8439), .A2(n9904), .ZN(n7873) );
  NAND2_X1 U6534 ( .A1(n7872), .A2(n7873), .ZN(n7869) );
  NAND2_X1 U6535 ( .A1(n5068), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5137) );
  NAND2_X1 U6536 ( .A1(n4293), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5136) );
  NAND2_X1 U6537 ( .A1(n5132), .A2(n5131), .ZN(n5133) );
  NAND2_X1 U6538 ( .A1(n5154), .A2(n5133), .ZN(n6893) );
  INV_X1 U6539 ( .A(n6893), .ZN(n9853) );
  NAND2_X1 U6540 ( .A1(n4292), .A2(n9853), .ZN(n5135) );
  NAND2_X1 U6541 ( .A1(n6366), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5134) );
  NAND4_X1 U6542 ( .A1(n5137), .A2(n5136), .A3(n5135), .A4(n5134), .ZN(n8438)
         );
  XNOR2_X1 U6543 ( .A(n5139), .B(n5138), .ZN(n6350) );
  NAND2_X1 U6544 ( .A1(n6350), .A2(n7792), .ZN(n5146) );
  NAND2_X1 U6545 ( .A1(n5141), .A2(n5140), .ZN(n5142) );
  NOR2_X1 U6546 ( .A1(n5143), .A2(n5142), .ZN(n5150) );
  OR2_X1 U6547 ( .A1(n5150), .A2(n4999), .ZN(n5144) );
  XNOR2_X1 U6548 ( .A(n5144), .B(P2_IR_REG_8__SCAN_IN), .ZN(n6495) );
  AOI22_X1 U6549 ( .A1(n7788), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n5305), .B2(
        n6495), .ZN(n5145) );
  XNOR2_X1 U6550 ( .A(n8438), .B(n9857), .ZN(n9840) );
  NAND2_X1 U6551 ( .A1(n8438), .A2(n9857), .ZN(n5147) );
  NAND2_X1 U6552 ( .A1(n9837), .A2(n5147), .ZN(n7179) );
  XNOR2_X1 U6553 ( .A(n5148), .B(n4850), .ZN(n6357) );
  NAND2_X1 U6554 ( .A1(n6357), .A2(n7792), .ZN(n5152) );
  INV_X1 U6555 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5149) );
  NAND2_X1 U6556 ( .A1(n5150), .A2(n5149), .ZN(n5188) );
  NAND2_X1 U6557 ( .A1(n5188), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5162) );
  XNOR2_X1 U6558 ( .A(n5162), .B(P2_IR_REG_9__SCAN_IN), .ZN(n6507) );
  AOI22_X1 U6559 ( .A1(n7788), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n5305), .B2(
        n6507), .ZN(n5151) );
  NAND2_X1 U6560 ( .A1(n5068), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5159) );
  NAND2_X1 U6561 ( .A1(n4293), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5158) );
  NAND2_X1 U6562 ( .A1(n5154), .A2(n5153), .ZN(n5155) );
  AND2_X1 U6563 ( .A1(n5181), .A2(n5155), .ZN(n7188) );
  NAND2_X1 U6564 ( .A1(n4292), .A2(n7188), .ZN(n5157) );
  NAND2_X1 U6565 ( .A1(n6366), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5156) );
  NAND4_X1 U6566 ( .A1(n5159), .A2(n5158), .A3(n5157), .A4(n5156), .ZN(n8437)
         );
  NAND2_X1 U6567 ( .A1(n9915), .A2(n8437), .ZN(n7880) );
  INV_X1 U6568 ( .A(n9915), .ZN(n7189) );
  INV_X1 U6569 ( .A(n8437), .ZN(n9849) );
  NAND2_X1 U6570 ( .A1(n7189), .A2(n9849), .ZN(n7881) );
  XNOR2_X1 U6571 ( .A(n5160), .B(n4851), .ZN(n6362) );
  INV_X1 U6572 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5161) );
  NAND2_X1 U6573 ( .A1(n5162), .A2(n5161), .ZN(n5163) );
  NAND2_X1 U6574 ( .A1(n5163), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5165) );
  NAND2_X1 U6575 ( .A1(n5165), .A2(n5164), .ZN(n5175) );
  OR2_X1 U6576 ( .A1(n5165), .A2(n5164), .ZN(n5166) );
  AOI22_X1 U6577 ( .A1(n7788), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n5305), .B2(
        n9770), .ZN(n5167) );
  NAND2_X1 U6578 ( .A1(n5078), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5172) );
  XNOR2_X1 U6579 ( .A(n5181), .B(P2_REG3_REG_10__SCAN_IN), .ZN(n9822) );
  NAND2_X1 U6580 ( .A1(n4291), .A2(n9822), .ZN(n5171) );
  NAND2_X1 U6581 ( .A1(n6366), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5170) );
  INV_X1 U6582 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n5168) );
  OR2_X1 U6583 ( .A1(n5388), .A2(n5168), .ZN(n5169) );
  AND2_X1 U6584 ( .A1(n9823), .A2(n4655), .ZN(n5200) );
  OR2_X1 U6585 ( .A1(n7811), .A2(n5200), .ZN(n7424) );
  XNOR2_X1 U6586 ( .A(n5174), .B(n5173), .ZN(n6371) );
  NAND2_X1 U6587 ( .A1(n6371), .A2(n7792), .ZN(n5178) );
  NAND2_X1 U6588 ( .A1(n5175), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5176) );
  XNOR2_X1 U6589 ( .A(n5176), .B(P2_IR_REG_11__SCAN_IN), .ZN(n6524) );
  AOI22_X1 U6590 ( .A1(n7788), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n5305), .B2(
        n6524), .ZN(n5177) );
  NAND2_X1 U6591 ( .A1(n5178), .A2(n5177), .ZN(n9926) );
  NAND2_X1 U6592 ( .A1(n5078), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5187) );
  INV_X1 U6593 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n5180) );
  INV_X1 U6594 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n5179) );
  OAI21_X1 U6595 ( .B1(n5181), .B2(n5180), .A(n5179), .ZN(n5182) );
  AND2_X1 U6596 ( .A1(n5182), .A2(n5192), .ZN(n7431) );
  NAND2_X1 U6597 ( .A1(n4291), .A2(n7431), .ZN(n5186) );
  NAND2_X1 U6598 ( .A1(n5068), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5185) );
  INV_X1 U6599 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n5183) );
  OR2_X1 U6600 ( .A1(n5070), .A2(n5183), .ZN(n5184) );
  INV_X1 U6601 ( .A(n5199), .ZN(n8436) );
  AND2_X1 U6602 ( .A1(n9926), .A2(n8436), .ZN(n5201) );
  OR2_X1 U6603 ( .A1(n7424), .A2(n5201), .ZN(n7403) );
  NAND2_X1 U6604 ( .A1(n6422), .A2(n7792), .ZN(n5191) );
  NAND2_X1 U6605 ( .A1(n5260), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5189) );
  XNOR2_X1 U6606 ( .A(n5189), .B(P2_IR_REG_12__SCAN_IN), .ZN(n6574) );
  AOI22_X1 U6607 ( .A1(n7788), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n5305), .B2(
        n6574), .ZN(n5190) );
  NAND2_X1 U6608 ( .A1(n4293), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5197) );
  NAND2_X1 U6609 ( .A1(n5192), .A2(n10078), .ZN(n5193) );
  AND2_X1 U6610 ( .A1(n5214), .A2(n5193), .ZN(n9804) );
  NAND2_X1 U6611 ( .A1(n4291), .A2(n9804), .ZN(n5196) );
  NAND2_X1 U6612 ( .A1(n6366), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5195) );
  NAND2_X1 U6613 ( .A1(n5068), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5194) );
  NAND2_X1 U6614 ( .A1(n9809), .A2(n7412), .ZN(n7897) );
  OR2_X1 U6615 ( .A1(n7403), .A2(n9800), .ZN(n5198) );
  OR2_X1 U6616 ( .A1(n9926), .A2(n5199), .ZN(n7894) );
  NAND2_X1 U6617 ( .A1(n9926), .A2(n5199), .ZN(n7890) );
  NAND2_X1 U6618 ( .A1(n7894), .A2(n7890), .ZN(n7814) );
  NAND2_X1 U6619 ( .A1(n9823), .A2(n7232), .ZN(n7884) );
  OR2_X1 U6620 ( .A1(n7189), .A2(n8437), .ZN(n9824) );
  OR2_X1 U6621 ( .A1(n9800), .A2(n7404), .ZN(n5202) );
  NAND2_X1 U6622 ( .A1(n5206), .A2(n5205), .ZN(n5210) );
  AND2_X1 U6623 ( .A1(n5208), .A2(n5207), .ZN(n5209) );
  NAND2_X1 U6624 ( .A1(n6485), .A2(n7792), .ZN(n5212) );
  OAI21_X1 U6625 ( .B1(n5260), .B2(P2_IR_REG_12__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5227) );
  XNOR2_X1 U6626 ( .A(n5227), .B(P2_IR_REG_13__SCAN_IN), .ZN(n6577) );
  AOI22_X1 U6627 ( .A1(n7788), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n5305), .B2(
        n6577), .ZN(n5211) );
  NAND2_X1 U6628 ( .A1(n5078), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n5220) );
  NAND2_X1 U6629 ( .A1(n5068), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5219) );
  INV_X1 U6630 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5213) );
  NAND2_X1 U6631 ( .A1(n5214), .A2(n5213), .ZN(n5215) );
  AND2_X1 U6632 ( .A1(n5231), .A2(n5215), .ZN(n7419) );
  NAND2_X1 U6633 ( .A1(n4292), .A2(n7419), .ZN(n5218) );
  INV_X1 U6634 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n5216) );
  OR2_X1 U6635 ( .A1(n5070), .A2(n5216), .ZN(n5217) );
  OR2_X1 U6636 ( .A1(n8796), .A2(n7606), .ZN(n7904) );
  NAND2_X1 U6637 ( .A1(n8796), .A2(n7606), .ZN(n7903) );
  NAND2_X1 U6638 ( .A1(n7904), .A2(n7903), .ZN(n7892) );
  INV_X1 U6639 ( .A(n7412), .ZN(n8435) );
  OR2_X1 U6640 ( .A1(n9809), .A2(n8435), .ZN(n7406) );
  AND2_X1 U6641 ( .A1(n7892), .A2(n7406), .ZN(n5221) );
  INV_X1 U6642 ( .A(n7606), .ZN(n8434) );
  NAND2_X1 U6643 ( .A1(n8796), .A2(n8434), .ZN(n5222) );
  NAND2_X1 U6644 ( .A1(n5224), .A2(n5223), .ZN(n5226) );
  XNOR2_X1 U6645 ( .A(n5226), .B(n5225), .ZN(n6481) );
  NAND2_X1 U6646 ( .A1(n6481), .A2(n7792), .ZN(n5230) );
  NAND2_X1 U6647 ( .A1(n5227), .A2(n5257), .ZN(n5228) );
  NAND2_X1 U6648 ( .A1(n5228), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5241) );
  XNOR2_X1 U6649 ( .A(n5241), .B(P2_IR_REG_14__SCAN_IN), .ZN(n6649) );
  AOI22_X1 U6650 ( .A1(n7788), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n5305), .B2(
        n6649), .ZN(n5229) );
  NAND2_X1 U6651 ( .A1(n4293), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n5237) );
  NAND2_X1 U6652 ( .A1(n5231), .A2(n10091), .ZN(n5232) );
  AND2_X1 U6653 ( .A1(n5247), .A2(n5232), .ZN(n7602) );
  NAND2_X1 U6654 ( .A1(n4291), .A2(n7602), .ZN(n5236) );
  NAND2_X1 U6655 ( .A1(n5068), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5235) );
  INV_X1 U6656 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n5233) );
  OR2_X1 U6657 ( .A1(n5070), .A2(n5233), .ZN(n5234) );
  NAND2_X1 U6658 ( .A1(n8791), .A2(n7411), .ZN(n7910) );
  NAND2_X1 U6659 ( .A1(n8697), .A2(n7910), .ZN(n7902) );
  INV_X1 U6660 ( .A(n7411), .ZN(n8433) );
  OR2_X1 U6661 ( .A1(n8791), .A2(n8433), .ZN(n5238) );
  XNOR2_X1 U6662 ( .A(n5240), .B(n5239), .ZN(n6553) );
  NAND2_X1 U6663 ( .A1(n6553), .A2(n7792), .ZN(n5245) );
  INV_X1 U6664 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5258) );
  NAND2_X1 U6665 ( .A1(n5241), .A2(n5258), .ZN(n5242) );
  NAND2_X1 U6666 ( .A1(n5242), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5243) );
  XNOR2_X1 U6667 ( .A(n5243), .B(P2_IR_REG_15__SCAN_IN), .ZN(n7004) );
  AOI22_X1 U6668 ( .A1(n7788), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n5305), .B2(
        n7004), .ZN(n5244) );
  NAND2_X1 U6669 ( .A1(n5068), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5253) );
  NAND2_X1 U6670 ( .A1(n5078), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n5252) );
  INV_X1 U6671 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n5246) );
  NAND2_X1 U6672 ( .A1(n5247), .A2(n5246), .ZN(n5248) );
  AND2_X1 U6673 ( .A1(n5266), .A2(n5248), .ZN(n8691) );
  NAND2_X1 U6674 ( .A1(n5347), .A2(n8691), .ZN(n5251) );
  INV_X1 U6675 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n5249) );
  OR2_X1 U6676 ( .A1(n5070), .A2(n5249), .ZN(n5250) );
  XNOR2_X1 U6677 ( .A(n8786), .B(n7607), .ZN(n7909) );
  XNOR2_X1 U6678 ( .A(n5255), .B(n5254), .ZN(n6513) );
  NAND2_X1 U6679 ( .A1(n6513), .A2(n7792), .ZN(n5265) );
  INV_X1 U6680 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5256) );
  NAND4_X1 U6681 ( .A1(n5258), .A2(n10080), .A3(n5257), .A4(n5256), .ZN(n5259)
         );
  OAI21_X1 U6682 ( .B1(n5260), .B2(n5259), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n5261) );
  MUX2_X1 U6683 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5261), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n5263) );
  NAND2_X1 U6684 ( .A1(n5263), .A2(n5262), .ZN(n7571) );
  INV_X1 U6685 ( .A(n7571), .ZN(n7008) );
  AOI22_X1 U6686 ( .A1(n7788), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n5305), .B2(
        n7008), .ZN(n5264) );
  NAND2_X1 U6687 ( .A1(n5068), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5271) );
  NAND2_X1 U6688 ( .A1(n4293), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n5270) );
  NAND2_X1 U6689 ( .A1(n5266), .A2(n7558), .ZN(n5267) );
  AND2_X1 U6690 ( .A1(n5279), .A2(n5267), .ZN(n7561) );
  NAND2_X1 U6691 ( .A1(n5347), .A2(n7561), .ZN(n5269) );
  INV_X1 U6692 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n7566) );
  OR2_X1 U6693 ( .A1(n5070), .A2(n7566), .ZN(n5268) );
  OR2_X1 U6694 ( .A1(n8834), .A2(n8674), .ZN(n8669) );
  NAND2_X1 U6695 ( .A1(n8834), .A2(n8674), .ZN(n7915) );
  NAND2_X1 U6696 ( .A1(n8669), .A2(n7915), .ZN(n7918) );
  INV_X1 U6697 ( .A(n8674), .ZN(n8431) );
  XNOR2_X1 U6698 ( .A(n5274), .B(n5273), .ZN(n6601) );
  NAND2_X1 U6699 ( .A1(n6601), .A2(n7792), .ZN(n5277) );
  NAND2_X1 U6700 ( .A1(n5262), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5275) );
  XNOR2_X1 U6701 ( .A(n5275), .B(n4975), .ZN(n7572) );
  INV_X1 U6702 ( .A(n7572), .ZN(n9790) );
  AOI22_X1 U6703 ( .A1(n7788), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n5305), .B2(
        n9790), .ZN(n5276) );
  NAND2_X1 U6704 ( .A1(n5068), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5284) );
  NAND2_X1 U6705 ( .A1(n5078), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n5283) );
  INV_X1 U6706 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n5278) );
  NAND2_X1 U6707 ( .A1(n5279), .A2(n5278), .ZN(n5280) );
  AND2_X1 U6708 ( .A1(n5293), .A2(n5280), .ZN(n8683) );
  NAND2_X1 U6709 ( .A1(n5347), .A2(n8683), .ZN(n5282) );
  INV_X1 U6710 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n7567) );
  OR2_X1 U6711 ( .A1(n5070), .A2(n7567), .ZN(n5281) );
  NAND2_X1 U6712 ( .A1(n8668), .A2(n8654), .ZN(n7919) );
  NAND2_X1 U6713 ( .A1(n7920), .A2(n7919), .ZN(n8677) );
  INV_X1 U6714 ( .A(n8654), .ZN(n8430) );
  XNOR2_X1 U6715 ( .A(n5287), .B(n5286), .ZN(n6749) );
  NAND2_X1 U6716 ( .A1(n6749), .A2(n7792), .ZN(n5291) );
  NAND2_X1 U6717 ( .A1(n5288), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5289) );
  XNOR2_X1 U6718 ( .A(n5289), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8446) );
  AOI22_X1 U6719 ( .A1(n5092), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n5305), .B2(
        n8446), .ZN(n5290) );
  NAND2_X1 U6720 ( .A1(n4293), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n5298) );
  NAND2_X1 U6721 ( .A1(n6366), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n5297) );
  INV_X1 U6722 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n5292) );
  NAND2_X1 U6723 ( .A1(n5293), .A2(n5292), .ZN(n5294) );
  AND2_X1 U6724 ( .A1(n5308), .A2(n5294), .ZN(n8659) );
  NAND2_X1 U6725 ( .A1(n5347), .A2(n8659), .ZN(n5296) );
  NAND2_X1 U6726 ( .A1(n5068), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n5295) );
  NAND4_X1 U6727 ( .A1(n5298), .A2(n5297), .A3(n5296), .A4(n5295), .ZN(n8429)
         );
  NOR2_X1 U6728 ( .A1(n8769), .A2(n8429), .ZN(n5299) );
  INV_X1 U6729 ( .A(n8769), .ZN(n8662) );
  XNOR2_X1 U6730 ( .A(n5301), .B(n5300), .ZN(n6779) );
  NAND2_X1 U6731 ( .A1(n6779), .A2(n7792), .ZN(n5307) );
  NAND2_X1 U6732 ( .A1(n5302), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5304) );
  XNOR2_X2 U6733 ( .A(n5304), .B(n5303), .ZN(n8682) );
  INV_X1 U6734 ( .A(n8682), .ZN(n8539) );
  AOI22_X1 U6735 ( .A1(n7788), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n5305), .B2(
        n8539), .ZN(n5306) );
  NAND2_X1 U6736 ( .A1(n5068), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n5314) );
  NAND2_X1 U6737 ( .A1(n4293), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n5313) );
  NAND2_X1 U6738 ( .A1(n5308), .A2(n8354), .ZN(n5309) );
  AND2_X1 U6739 ( .A1(n5310), .A2(n5309), .ZN(n8642) );
  NAND2_X1 U6740 ( .A1(n5347), .A2(n8642), .ZN(n5312) );
  NAND2_X1 U6741 ( .A1(n6366), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n5311) );
  NAND4_X1 U6742 ( .A1(n5314), .A2(n5313), .A3(n5312), .A4(n5311), .ZN(n8428)
         );
  NAND2_X1 U6743 ( .A1(n8757), .A2(n8638), .ZN(n7937) );
  NAND2_X1 U6744 ( .A1(n8615), .A2(n7937), .ZN(n8620) );
  XNOR2_X1 U6745 ( .A(n5319), .B(n5318), .ZN(n6944) );
  NAND2_X1 U6746 ( .A1(n6944), .A2(n7792), .ZN(n5321) );
  NAND2_X1 U6747 ( .A1(n5092), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n5320) );
  INV_X1 U6748 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n5322) );
  NAND2_X1 U6749 ( .A1(n5323), .A2(n5322), .ZN(n5324) );
  AND2_X1 U6750 ( .A1(n5332), .A2(n5324), .ZN(n8607) );
  NAND2_X1 U6751 ( .A1(n8607), .A2(n5347), .ZN(n5327) );
  AOI22_X1 U6752 ( .A1(n5068), .A2(P2_REG0_REG_21__SCAN_IN), .B1(n4293), .B2(
        P2_REG1_REG_21__SCAN_IN), .ZN(n5326) );
  NAND2_X1 U6753 ( .A1(n6366), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n5325) );
  NOR2_X1 U6754 ( .A1(n8602), .A2(n8617), .ZN(n5328) );
  INV_X1 U6755 ( .A(n8617), .ZN(n8426) );
  XNOR2_X1 U6756 ( .A(n5330), .B(n5329), .ZN(n6992) );
  NAND2_X1 U6757 ( .A1(n5092), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n5331) );
  INV_X1 U6758 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n8402) );
  NAND2_X1 U6759 ( .A1(n5332), .A2(n8402), .ZN(n5333) );
  NAND2_X1 U6760 ( .A1(n5344), .A2(n5333), .ZN(n8583) );
  OR2_X1 U6761 ( .A1(n8583), .A2(n5423), .ZN(n5336) );
  AOI22_X1 U6762 ( .A1(n5068), .A2(P2_REG0_REG_22__SCAN_IN), .B1(n4293), .B2(
        P2_REG1_REG_22__SCAN_IN), .ZN(n5335) );
  NAND2_X1 U6763 ( .A1(n6366), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n5334) );
  NAND2_X1 U6764 ( .A1(n8745), .A2(n8363), .ZN(n7929) );
  OR2_X1 U6765 ( .A1(n5338), .A2(n5337), .ZN(n5339) );
  NAND2_X1 U6766 ( .A1(n5340), .A2(n5339), .ZN(n7097) );
  NAND2_X1 U6767 ( .A1(n7097), .A2(n7792), .ZN(n5342) );
  NAND2_X1 U6768 ( .A1(n5092), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n5341) );
  NAND2_X1 U6769 ( .A1(n5344), .A2(n5343), .ZN(n5345) );
  AND2_X1 U6770 ( .A1(n5346), .A2(n5345), .ZN(n8575) );
  NAND2_X1 U6771 ( .A1(n8575), .A2(n5347), .ZN(n5352) );
  INV_X1 U6772 ( .A(n5068), .ZN(n5388) );
  INV_X1 U6773 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n10075) );
  NAND2_X1 U6774 ( .A1(n6366), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n5349) );
  NAND2_X1 U6775 ( .A1(n4293), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n5348) );
  OAI211_X1 U6776 ( .C1(n5388), .C2(n10075), .A(n5349), .B(n5348), .ZN(n5350)
         );
  INV_X1 U6777 ( .A(n5350), .ZN(n5351) );
  NAND2_X1 U6778 ( .A1(n5352), .A2(n5351), .ZN(n8546) );
  NAND2_X1 U6779 ( .A1(n8819), .A2(n8546), .ZN(n7944) );
  INV_X1 U6780 ( .A(n8546), .ZN(n8591) );
  NAND2_X1 U6781 ( .A1(n8346), .A2(n8591), .ZN(n7945) );
  NAND2_X1 U6782 ( .A1(n8735), .A2(n8372), .ZN(n7951) );
  NAND2_X1 U6783 ( .A1(n8552), .A2(n8551), .ZN(n8550) );
  OAI21_X1 U6784 ( .B1(n8735), .B2(n8425), .A(n8550), .ZN(n8528) );
  INV_X1 U6785 ( .A(n5353), .ZN(n5356) );
  INV_X1 U6786 ( .A(n5354), .ZN(n5355) );
  INV_X1 U6787 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7402) );
  INV_X1 U6788 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n10121) );
  MUX2_X1 U6789 ( .A(n7402), .B(n10121), .S(n6326), .Z(n5359) );
  INV_X1 U6790 ( .A(SI_25_), .ZN(n5358) );
  NAND2_X1 U6791 ( .A1(n5359), .A2(n5358), .ZN(n5373) );
  INV_X1 U6792 ( .A(n5359), .ZN(n5360) );
  NAND2_X1 U6793 ( .A1(n5360), .A2(SI_25_), .ZN(n5361) );
  NAND2_X1 U6794 ( .A1(n5373), .A2(n5361), .ZN(n5374) );
  NAND2_X1 U6795 ( .A1(n7397), .A2(n7792), .ZN(n5363) );
  NAND2_X1 U6796 ( .A1(n5092), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n5362) );
  INV_X1 U6797 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n10142) );
  NAND2_X1 U6798 ( .A1(n5364), .A2(n10142), .ZN(n5365) );
  INV_X1 U6799 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n5368) );
  NAND2_X1 U6800 ( .A1(n5068), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n5367) );
  NAND2_X1 U6801 ( .A1(n4293), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n5366) );
  OAI211_X1 U6802 ( .C1(n5368), .C2(n5070), .A(n5367), .B(n5366), .ZN(n5369)
         );
  AOI21_X1 U6803 ( .B1(n8537), .B2(n5347), .A(n5369), .ZN(n8413) );
  NAND2_X1 U6804 ( .A1(n8731), .A2(n8413), .ZN(n7954) );
  NAND2_X1 U6805 ( .A1(n8528), .A2(n8530), .ZN(n5372) );
  INV_X1 U6806 ( .A(n8413), .ZN(n8548) );
  INV_X1 U6807 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7442) );
  INV_X1 U6808 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n5376) );
  MUX2_X1 U6809 ( .A(n7442), .B(n5376), .S(n6326), .Z(n5378) );
  INV_X1 U6810 ( .A(SI_26_), .ZN(n5377) );
  NAND2_X1 U6811 ( .A1(n5378), .A2(n5377), .ZN(n5394) );
  INV_X1 U6812 ( .A(n5378), .ZN(n5379) );
  NAND2_X1 U6813 ( .A1(n5379), .A2(SI_26_), .ZN(n5380) );
  AND2_X1 U6814 ( .A1(n5394), .A2(n5380), .ZN(n5392) );
  NAND2_X1 U6815 ( .A1(n7384), .A2(n7792), .ZN(n5382) );
  NAND2_X1 U6816 ( .A1(n7788), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n5381) );
  INV_X1 U6817 ( .A(n5384), .ZN(n5383) );
  NAND2_X1 U6818 ( .A1(n5383), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5402) );
  INV_X1 U6819 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8416) );
  NAND2_X1 U6820 ( .A1(n5384), .A2(n8416), .ZN(n5385) );
  NAND2_X1 U6821 ( .A1(n5402), .A2(n5385), .ZN(n8521) );
  INV_X1 U6822 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n10077) );
  NAND2_X1 U6823 ( .A1(n6366), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n5387) );
  NAND2_X1 U6824 ( .A1(n4293), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n5386) );
  OAI211_X1 U6825 ( .C1(n5388), .C2(n10077), .A(n5387), .B(n5386), .ZN(n5389)
         );
  INV_X1 U6826 ( .A(n5389), .ZN(n5390) );
  NAND2_X1 U6827 ( .A1(n5391), .A2(n5390), .ZN(n8504) );
  NAND2_X1 U6828 ( .A1(n8814), .A2(n8504), .ZN(n7958) );
  INV_X1 U6829 ( .A(n8504), .ZN(n8338) );
  INV_X1 U6830 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n7522) );
  INV_X1 U6831 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n7520) );
  MUX2_X1 U6832 ( .A(n7522), .B(n7520), .S(n6327), .Z(n5397) );
  INV_X1 U6833 ( .A(SI_27_), .ZN(n5396) );
  NAND2_X1 U6834 ( .A1(n5397), .A2(n5396), .ZN(n5416) );
  INV_X1 U6835 ( .A(n5397), .ZN(n5398) );
  NAND2_X1 U6836 ( .A1(n5398), .A2(SI_27_), .ZN(n5399) );
  AND2_X1 U6837 ( .A1(n5416), .A2(n5399), .ZN(n5414) );
  NAND2_X1 U6838 ( .A1(n7519), .A2(n7792), .ZN(n5401) );
  NAND2_X1 U6839 ( .A1(n5092), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n5400) );
  INV_X1 U6840 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n8335) );
  NAND2_X1 U6841 ( .A1(n5402), .A2(n8335), .ZN(n5403) );
  INV_X1 U6842 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n5406) );
  NAND2_X1 U6843 ( .A1(n5068), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n5405) );
  NAND2_X1 U6844 ( .A1(n4294), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n5404) );
  OAI211_X1 U6845 ( .C1(n5406), .C2(n5070), .A(n5405), .B(n5404), .ZN(n5407)
         );
  NAND2_X1 U6846 ( .A1(n8500), .A2(n8412), .ZN(n5410) );
  INV_X1 U6847 ( .A(n5410), .ZN(n5408) );
  NAND2_X1 U6848 ( .A1(n8719), .A2(n8412), .ZN(n7962) );
  INV_X1 U6849 ( .A(n5409), .ZN(n5412) );
  NAND2_X1 U6850 ( .A1(n8814), .A2(n8338), .ZN(n8491) );
  AND2_X1 U6851 ( .A1(n8491), .A2(n5410), .ZN(n5411) );
  INV_X1 U6852 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n7713) );
  INV_X1 U6853 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n5417) );
  MUX2_X1 U6854 ( .A(n7713), .B(n5417), .S(n6326), .Z(n5515) );
  XNOR2_X1 U6855 ( .A(n5515), .B(SI_28_), .ZN(n5512) );
  NAND2_X1 U6856 ( .A1(n7545), .A2(n7792), .ZN(n5419) );
  NAND2_X1 U6857 ( .A1(n5092), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n5418) );
  INV_X1 U6858 ( .A(n5421), .ZN(n5420) );
  NAND2_X1 U6859 ( .A1(n5420), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n8472) );
  INV_X1 U6860 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n7768) );
  NAND2_X1 U6861 ( .A1(n5421), .A2(n7768), .ZN(n5422) );
  NAND2_X1 U6862 ( .A1(n8472), .A2(n5422), .ZN(n8484) );
  INV_X1 U6863 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n8483) );
  NAND2_X1 U6864 ( .A1(n5068), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n5425) );
  NAND2_X1 U6865 ( .A1(n4293), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n5424) );
  OAI211_X1 U6866 ( .C1(n8483), .C2(n5070), .A(n5425), .B(n5424), .ZN(n5426)
         );
  INV_X1 U6867 ( .A(n5426), .ZN(n5427) );
  NAND2_X1 U6868 ( .A1(n7772), .A2(n8336), .ZN(n7967) );
  NAND2_X1 U6869 ( .A1(n4318), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5430) );
  XNOR2_X1 U6870 ( .A(n5430), .B(n5429), .ZN(n7831) );
  NAND2_X1 U6871 ( .A1(n5431), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5432) );
  MUX2_X1 U6872 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5432), .S(
        P2_IR_REG_20__SCAN_IN), .Z(n5433) );
  NAND2_X1 U6873 ( .A1(n7989), .A2(n7983), .ZN(n6926) );
  XNOR2_X1 U6874 ( .A(n5453), .B(n6926), .ZN(n5434) );
  NAND2_X1 U6875 ( .A1(n5434), .A2(n8682), .ZN(n8679) );
  AND2_X1 U6876 ( .A1(n7983), .A2(n8539), .ZN(n5435) );
  NAND2_X1 U6877 ( .A1(n7833), .A2(n5435), .ZN(n6764) );
  NAND2_X1 U6878 ( .A1(n8679), .A2(n6764), .ZN(n9941) );
  NAND2_X1 U6879 ( .A1(n6920), .A2(n9887), .ZN(n6919) );
  INV_X1 U6880 ( .A(n7225), .ZN(n6768) );
  INV_X1 U6881 ( .A(n9823), .ZN(n9923) );
  INV_X1 U6882 ( .A(n8791), .ZN(n7604) );
  NAND2_X1 U6883 ( .A1(n7599), .A2(n7604), .ZN(n8690) );
  INV_X1 U6884 ( .A(n5436), .ZN(n8689) );
  INV_X1 U6885 ( .A(n8668), .ZN(n8830) );
  NAND3_X1 U6886 ( .A1(n8599), .A2(n8586), .A3(n8819), .ZN(n8572) );
  NAND2_X1 U6887 ( .A1(n7833), .A2(n7831), .ZN(n9880) );
  OR2_X2 U6888 ( .A1(n9880), .A2(n7829), .ZN(n6682) );
  AOI211_X1 U6889 ( .C1(n7772), .C2(n8495), .A(n6682), .B(n4554), .ZN(n8487)
         );
  INV_X1 U6890 ( .A(n6972), .ZN(n9879) );
  NAND2_X1 U6891 ( .A1(n6969), .A2(n7853), .ZN(n5437) );
  INV_X1 U6892 ( .A(n6770), .ZN(n7848) );
  NAND2_X1 U6893 ( .A1(n6772), .A2(n7838), .ZN(n6948) );
  INV_X1 U6894 ( .A(n7834), .ZN(n7840) );
  INV_X1 U6895 ( .A(n7808), .ZN(n6851) );
  AND2_X1 U6896 ( .A1(n6851), .A2(n7835), .ZN(n6848) );
  XNOR2_X1 U6897 ( .A(n8440), .B(n9897), .ZN(n7810) );
  NOR2_X1 U6898 ( .A1(n8440), .A2(n7859), .ZN(n7868) );
  NOR2_X1 U6899 ( .A1(n7869), .A2(n7868), .ZN(n5438) );
  NAND2_X1 U6900 ( .A1(n7130), .A2(n7873), .ZN(n9842) );
  INV_X1 U6901 ( .A(n9840), .ZN(n9841) );
  INV_X1 U6902 ( .A(n8438), .ZN(n7876) );
  NAND2_X1 U6903 ( .A1(n7876), .A2(n9857), .ZN(n7875) );
  NAND2_X1 U6904 ( .A1(n5439), .A2(n7881), .ZN(n7433) );
  INV_X1 U6905 ( .A(n7433), .ZN(n5441) );
  INV_X1 U6906 ( .A(n7890), .ZN(n5440) );
  OR2_X1 U6907 ( .A1(n9816), .A2(n5440), .ZN(n9796) );
  INV_X1 U6908 ( .A(n9800), .ZN(n9807) );
  INV_X1 U6909 ( .A(n7814), .ZN(n7437) );
  AND2_X1 U6910 ( .A1(n7437), .A2(n7885), .ZN(n7434) );
  OR2_X1 U6911 ( .A1(n5440), .A2(n7434), .ZN(n9797) );
  INV_X1 U6912 ( .A(n7892), .ZN(n7817) );
  OR2_X1 U6913 ( .A1(n7902), .A2(n7909), .ZN(n7506) );
  INV_X1 U6914 ( .A(n7915), .ZN(n5443) );
  OR2_X1 U6915 ( .A1(n7909), .A2(n8697), .ZN(n8695) );
  INV_X1 U6916 ( .A(n8786), .ZN(n8694) );
  NAND2_X1 U6917 ( .A1(n8694), .A2(n8432), .ZN(n5442) );
  AND2_X1 U6918 ( .A1(n8695), .A2(n5442), .ZN(n7507) );
  OR2_X1 U6919 ( .A1(n8769), .A2(n8675), .ZN(n8633) );
  NAND2_X1 U6920 ( .A1(n8769), .A2(n8675), .ZN(n7924) );
  INV_X1 U6921 ( .A(n7920), .ZN(n5444) );
  INV_X1 U6922 ( .A(n8677), .ZN(n8671) );
  OR2_X1 U6923 ( .A1(n5444), .A2(n8671), .ZN(n8649) );
  AND2_X1 U6924 ( .A1(n8651), .A2(n8649), .ZN(n5445) );
  NAND2_X1 U6925 ( .A1(n8650), .A2(n5445), .ZN(n8634) );
  OR2_X1 U6926 ( .A1(n8639), .A2(n8655), .ZN(n7935) );
  NAND2_X1 U6927 ( .A1(n8639), .A2(n8655), .ZN(n8613) );
  NAND2_X1 U6928 ( .A1(n7935), .A2(n8613), .ZN(n7802) );
  INV_X1 U6929 ( .A(n8633), .ZN(n7933) );
  NOR2_X1 U6930 ( .A1(n7802), .A2(n7933), .ZN(n5446) );
  AND2_X1 U6931 ( .A1(n7937), .A2(n8613), .ZN(n7926) );
  AND2_X1 U6932 ( .A1(n8751), .A2(n8617), .ZN(n7928) );
  NOR2_X1 U6933 ( .A1(n8590), .A2(n7928), .ZN(n5447) );
  INV_X1 U6934 ( .A(n8565), .ZN(n7940) );
  NOR2_X1 U6935 ( .A1(n8566), .A2(n7940), .ZN(n5449) );
  INV_X1 U6936 ( .A(n7945), .ZN(n5448) );
  INV_X1 U6937 ( .A(n8551), .ZN(n7822) );
  INV_X1 U6938 ( .A(n8510), .ZN(n5450) );
  INV_X1 U6939 ( .A(n7956), .ZN(n5451) );
  NAND3_X1 U6940 ( .A1(n5452), .A2(n7824), .A3(n7961), .ZN(n5454) );
  NAND2_X1 U6941 ( .A1(n7989), .A2(n7829), .ZN(n7997) );
  NAND2_X1 U6942 ( .A1(n6674), .A2(n7997), .ZN(n9818) );
  NAND2_X1 U6943 ( .A1(n5454), .A2(n9818), .ZN(n5462) );
  INV_X1 U6944 ( .A(n8472), .ZN(n5458) );
  INV_X1 U6945 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n10006) );
  NAND2_X1 U6946 ( .A1(n5068), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n5456) );
  NAND2_X1 U6947 ( .A1(n6366), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n5455) );
  OAI211_X1 U6948 ( .C1(n4295), .C2(n10006), .A(n5456), .B(n5455), .ZN(n5457)
         );
  AOI21_X1 U6949 ( .B1(n5458), .B2(n5347), .A(n5457), .ZN(n6784) );
  NAND2_X1 U6950 ( .A1(n5453), .A2(n7989), .ZN(n6692) );
  INV_X1 U6951 ( .A(n6692), .ZN(n6379) );
  NAND2_X1 U6952 ( .A1(n5459), .A2(n6379), .ZN(n9848) );
  OR2_X1 U6953 ( .A1(n6784), .A2(n9848), .ZN(n5461) );
  INV_X1 U6954 ( .A(n5459), .ZN(n6394) );
  NAND2_X1 U6955 ( .A1(n6394), .A2(n6379), .ZN(n9846) );
  OR2_X1 U6956 ( .A1(n8412), .A2(n9846), .ZN(n5460) );
  AND2_X1 U6957 ( .A1(n5461), .A2(n5460), .ZN(n7769) );
  OAI21_X1 U6958 ( .B1(n5520), .B2(n5462), .A(n7769), .ZN(n8480) );
  NOR4_X1 U6959 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_17__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_19__SCAN_IN), .ZN(n5466) );
  NOR4_X1 U6960 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_12__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_15__SCAN_IN), .ZN(n5465) );
  NOR4_X1 U6961 ( .A1(P2_D_REG_25__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n5464) );
  NOR4_X1 U6962 ( .A1(P2_D_REG_20__SCAN_IN), .A2(P2_D_REG_21__SCAN_IN), .A3(
        P2_D_REG_23__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n5463) );
  NAND4_X1 U6963 ( .A1(n5466), .A2(n5465), .A3(n5464), .A4(n5463), .ZN(n5488)
         );
  NOR2_X1 U6964 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .ZN(
        n5470) );
  NOR4_X1 U6965 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_2__SCAN_IN), .A4(P2_D_REG_3__SCAN_IN), .ZN(n5469) );
  NOR4_X1 U6966 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), .A3(
        P2_D_REG_10__SCAN_IN), .A4(P2_D_REG_11__SCAN_IN), .ZN(n5468) );
  NOR4_X1 U6967 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_5__SCAN_IN), .A3(
        P2_D_REG_6__SCAN_IN), .A4(P2_D_REG_7__SCAN_IN), .ZN(n5467) );
  NAND4_X1 U6968 ( .A1(n5470), .A2(n5469), .A3(n5468), .A4(n5467), .ZN(n5487)
         );
  NAND2_X1 U6969 ( .A1(n5471), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5473) );
  INV_X1 U6970 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5472) );
  XNOR2_X1 U6971 ( .A(n5473), .B(n5472), .ZN(n9869) );
  INV_X1 U6972 ( .A(n9869), .ZN(n5486) );
  INV_X1 U6973 ( .A(P2_B_REG_SCAN_IN), .ZN(n5484) );
  NAND2_X1 U6974 ( .A1(n5475), .A2(n5474), .ZN(n5476) );
  NAND2_X1 U6975 ( .A1(n5476), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5492) );
  INV_X1 U6976 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5491) );
  NAND2_X1 U6977 ( .A1(n5492), .A2(n5491), .ZN(n5494) );
  NAND2_X1 U6978 ( .A1(n5494), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5478) );
  INV_X1 U6979 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5477) );
  NOR2_X1 U6980 ( .A1(n5479), .A2(n4999), .ZN(n5480) );
  MUX2_X1 U6981 ( .A(n4999), .B(n5480), .S(P2_IR_REG_25__SCAN_IN), .Z(n5481)
         );
  INV_X1 U6982 ( .A(n5481), .ZN(n5482) );
  NAND2_X1 U6983 ( .A1(n5482), .A2(n5471), .ZN(n7400) );
  NAND2_X1 U6984 ( .A1(n9870), .A2(n5484), .ZN(n5483) );
  OAI211_X1 U6985 ( .C1(n5484), .C2(n9870), .A(n7400), .B(n5483), .ZN(n5485)
         );
  NAND2_X1 U6986 ( .A1(n5486), .A2(n5485), .ZN(n5489) );
  OAI21_X1 U6987 ( .B1(n5488), .B2(n5487), .A(n9867), .ZN(n6915) );
  NOR2_X1 U6988 ( .A1(P2_D_REG_0__SCAN_IN), .A2(n5489), .ZN(n5490) );
  AOI21_X1 U6989 ( .B1(n9870), .B2(n9869), .A(n5490), .ZN(n6912) );
  AND2_X1 U6990 ( .A1(n6915), .A2(n6912), .ZN(n6660) );
  OR2_X1 U6991 ( .A1(n5492), .A2(n5491), .ZN(n5493) );
  NAND2_X1 U6992 ( .A1(n5494), .A2(n5493), .ZN(n9871) );
  AND2_X1 U6993 ( .A1(n9871), .A2(P2_STATE_REG_SCAN_IN), .ZN(n5495) );
  NAND2_X1 U6994 ( .A1(n7400), .A2(n9869), .ZN(n9876) );
  INV_X1 U6995 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n5496) );
  NAND2_X1 U6996 ( .A1(n5496), .A2(n9867), .ZN(n5497) );
  NAND2_X1 U6997 ( .A1(n9876), .A2(n5497), .ZN(n6910) );
  AND2_X1 U6998 ( .A1(n7983), .A2(n8682), .ZN(n6668) );
  OR2_X1 U6999 ( .A1(n6692), .A2(n6668), .ZN(n6909) );
  NAND3_X1 U7000 ( .A1(n6663), .A2(n6910), .A3(n6909), .ZN(n5498) );
  NOR2_X1 U7001 ( .A1(n9868), .A2(n5498), .ZN(n5501) );
  AND2_X2 U7002 ( .A1(n6660), .A2(n5501), .ZN(n9959) );
  INV_X1 U7003 ( .A(n7772), .ZN(n8482) );
  OR2_X1 U7004 ( .A1(n9880), .A2(n6668), .ZN(n9937) );
  NAND2_X1 U7005 ( .A1(n9959), .A2(n9927), .ZN(n8777) );
  NAND2_X1 U7006 ( .A1(n5499), .A2(n4846), .ZN(P2_U3548) );
  INV_X1 U7007 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n5504) );
  INV_X1 U7008 ( .A(n6912), .ZN(n5500) );
  AND2_X1 U7009 ( .A1(n5501), .A2(n5500), .ZN(n5502) );
  MUX2_X1 U7010 ( .A(n5504), .B(n5503), .S(n9944), .Z(n5505) );
  NAND2_X1 U7011 ( .A1(n9944), .A2(n9927), .ZN(n8831) );
  NAND2_X1 U7012 ( .A1(n5505), .A2(n4845), .ZN(P2_U3516) );
  AND2_X1 U7013 ( .A1(n5506), .A2(n7824), .ZN(n5507) );
  INV_X1 U7014 ( .A(n8336), .ZN(n8503) );
  INV_X1 U7015 ( .A(SI_28_), .ZN(n5514) );
  INV_X1 U7016 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n7674) );
  INV_X1 U7017 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n10089) );
  MUX2_X1 U7018 ( .A(n7674), .B(n10089), .S(n6327), .Z(n5536) );
  XNOR2_X1 U7019 ( .A(n5536), .B(SI_29_), .ZN(n5516) );
  NAND2_X1 U7020 ( .A1(n7673), .A2(n7792), .ZN(n5518) );
  NAND2_X1 U7021 ( .A1(n5092), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n5517) );
  NAND2_X1 U7022 ( .A1(n8476), .A2(n6784), .ZN(n7987) );
  NAND2_X1 U7023 ( .A1(n7986), .A2(n7987), .ZN(n5521) );
  INV_X1 U7024 ( .A(n5519), .ZN(n7966) );
  INV_X1 U7025 ( .A(n5521), .ZN(n7826) );
  XNOR2_X1 U7026 ( .A(n4350), .B(n7826), .ZN(n5527) );
  NAND2_X1 U7027 ( .A1(n4293), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n5524) );
  NAND2_X1 U7028 ( .A1(n6366), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n5523) );
  NAND2_X1 U7029 ( .A1(n5068), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n5522) );
  AND3_X1 U7030 ( .A1(n5524), .A2(n5523), .A3(n5522), .ZN(n7800) );
  NOR2_X1 U7031 ( .A1(n8002), .A2(n5484), .ZN(n5525) );
  OR2_X1 U7032 ( .A1(n5525), .A2(n9848), .ZN(n7795) );
  OAI22_X1 U7033 ( .A1(n8336), .A2(n9846), .B1(n7800), .B2(n7795), .ZN(n5526)
         );
  AOI21_X1 U7034 ( .B1(n5527), .B2(n9818), .A(n5526), .ZN(n8479) );
  INV_X1 U7035 ( .A(n8476), .ZN(n5533) );
  OAI211_X1 U7036 ( .C1(n5533), .C2(n4554), .A(n5529), .B(n7321), .ZN(n8473)
         );
  NAND2_X1 U7037 ( .A1(n5530), .A2(n4841), .ZN(P2_U3549) );
  INV_X1 U7038 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n5532) );
  MUX2_X1 U7039 ( .A(n5532), .B(n5531), .S(n9944), .Z(n5534) );
  NAND2_X1 U7040 ( .A1(n5534), .A2(n4847), .ZN(P2_U3517) );
  INV_X1 U7041 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n5755) );
  INV_X1 U7042 ( .A(SI_29_), .ZN(n5535) );
  AND2_X1 U7043 ( .A1(n5536), .A2(n5535), .ZN(n5539) );
  INV_X1 U7044 ( .A(n5536), .ZN(n5537) );
  NAND2_X1 U7045 ( .A1(n5537), .A2(SI_29_), .ZN(n5538) );
  MUX2_X1 U7046 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .S(n6326), .Z(n5690) );
  INV_X1 U7047 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5545) );
  NAND4_X1 U7048 ( .A1(n5546), .A2(n5638), .A3(n5634), .A4(n5545), .ZN(n5551)
         );
  INV_X1 U7049 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n5549) );
  INV_X1 U7050 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5548) );
  INV_X1 U7051 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5547) );
  NAND4_X1 U7052 ( .A1(n5622), .A2(n5549), .A3(n5548), .A4(n5547), .ZN(n5550)
         );
  NOR2_X1 U7053 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n5553) );
  NOR3_X1 U7054 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .A3(
        P1_IR_REG_9__SCAN_IN), .ZN(n5552) );
  INV_X1 U7055 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5723) );
  INV_X1 U7056 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5556) );
  NAND2_X1 U7057 ( .A1(n5723), .A2(n5556), .ZN(n5557) );
  INV_X1 U7058 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5561) );
  NAND2_X2 U7059 ( .A1(n5709), .A2(n5559), .ZN(n5718) );
  NAND2_X1 U7060 ( .A1(n8840), .A2(n5696), .ZN(n5565) );
  NAND2_X1 U7061 ( .A1(n5581), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n5564) );
  NAND2_X1 U7062 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5566) );
  NAND2_X1 U7063 ( .A1(n6327), .A2(SI_0_), .ZN(n5569) );
  INV_X1 U7064 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5568) );
  NAND2_X1 U7065 ( .A1(n5569), .A2(n5568), .ZN(n5571) );
  AND2_X1 U7066 ( .A1(n5571), .A2(n5570), .ZN(n9393) );
  XNOR2_X1 U7067 ( .A(n5576), .B(P1_IR_REG_2__SCAN_IN), .ZN(n9492) );
  NAND2_X1 U7068 ( .A1(n6288), .A2(n9492), .ZN(n5574) );
  NAND2_X1 U7069 ( .A1(n7200), .A2(n7199), .ZN(n7282) );
  NAND2_X1 U7070 ( .A1(n5581), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n5580) );
  INV_X1 U7071 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n10156) );
  NAND2_X1 U7072 ( .A1(n5576), .A2(n10156), .ZN(n5577) );
  NAND2_X1 U7073 ( .A1(n5577), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5578) );
  XNOR2_X1 U7074 ( .A(n5578), .B(P1_IR_REG_3__SCAN_IN), .ZN(n9425) );
  NAND2_X1 U7075 ( .A1(n6288), .A2(n9425), .ZN(n5579) );
  NAND2_X1 U7076 ( .A1(n5581), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n5585) );
  OR2_X1 U7077 ( .A1(n5582), .A2(n9385), .ZN(n5583) );
  XNOR2_X1 U7078 ( .A(n5583), .B(P1_IR_REG_4__SCAN_IN), .ZN(n9501) );
  NAND2_X1 U7079 ( .A1(n6288), .A2(n9501), .ZN(n5584) );
  OAI211_X1 U7080 ( .C1(n6329), .C2(n5600), .A(n5585), .B(n5584), .ZN(n9623)
         );
  NAND2_X1 U7081 ( .A1(n5581), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n5591) );
  NAND2_X1 U7082 ( .A1(n5587), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5588) );
  MUX2_X1 U7083 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5588), .S(
        P1_IR_REG_5__SCAN_IN), .Z(n5589) );
  AND2_X1 U7084 ( .A1(n5586), .A2(n5589), .ZN(n9511) );
  NAND2_X1 U7085 ( .A1(n6288), .A2(n9511), .ZN(n5590) );
  OAI211_X1 U7086 ( .C1(n6343), .C2(n5600), .A(n5591), .B(n5590), .ZN(n9685)
         );
  INV_X1 U7087 ( .A(n9685), .ZN(n7257) );
  NAND2_X1 U7088 ( .A1(n5581), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n5594) );
  NAND2_X1 U7089 ( .A1(n5586), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5592) );
  XNOR2_X1 U7090 ( .A(n5592), .B(P1_IR_REG_6__SCAN_IN), .ZN(n6597) );
  NAND2_X1 U7091 ( .A1(n6288), .A2(n6597), .ZN(n5593) );
  INV_X1 U7092 ( .A(n5595), .ZN(n6348) );
  NAND2_X1 U7093 ( .A1(n5581), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n5599) );
  OR2_X1 U7094 ( .A1(n5596), .A2(n9385), .ZN(n5597) );
  XNOR2_X1 U7095 ( .A(n5597), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6564) );
  NAND2_X1 U7096 ( .A1(n6288), .A2(n6564), .ZN(n5598) );
  NAND2_X1 U7097 ( .A1(n5601), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5602) );
  XNOR2_X1 U7098 ( .A(n5602), .B(P1_IR_REG_8__SCAN_IN), .ZN(n9523) );
  INV_X1 U7099 ( .A(n9523), .ZN(n6352) );
  NAND2_X1 U7100 ( .A1(n6350), .A2(n5696), .ZN(n5604) );
  NAND2_X1 U7101 ( .A1(n5581), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n5603) );
  OAI211_X1 U7102 ( .C1(n5567), .C2(n6352), .A(n5604), .B(n5603), .ZN(n7299)
         );
  INV_X1 U7103 ( .A(n7299), .ZN(n7302) );
  NAND2_X1 U7104 ( .A1(n6357), .A2(n5696), .ZN(n5611) );
  NAND2_X1 U7105 ( .A1(n5605), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5606) );
  MUX2_X1 U7106 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5606), .S(
        P1_IR_REG_9__SCAN_IN), .Z(n5608) );
  INV_X1 U7107 ( .A(n5659), .ZN(n5607) );
  INV_X1 U7108 ( .A(n6610), .ZN(n6359) );
  OAI22_X1 U7109 ( .A1(n5665), .A2(n6361), .B1(n5567), .B2(n6359), .ZN(n5609)
         );
  INV_X1 U7110 ( .A(n5609), .ZN(n5610) );
  NAND2_X1 U7111 ( .A1(n6362), .A2(n5696), .ZN(n5615) );
  OR2_X1 U7112 ( .A1(n5659), .A2(n9385), .ZN(n5612) );
  XNOR2_X1 U7113 ( .A(n5612), .B(P1_IR_REG_10__SCAN_IN), .ZN(n6805) );
  INV_X1 U7114 ( .A(n6805), .ZN(n6605) );
  OAI22_X1 U7115 ( .A1(n5665), .A2(n6363), .B1(n5567), .B2(n6605), .ZN(n5613)
         );
  INV_X1 U7116 ( .A(n5613), .ZN(n5614) );
  NAND2_X1 U7117 ( .A1(n6371), .A2(n5696), .ZN(n5620) );
  INV_X1 U7118 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5616) );
  NAND2_X1 U7119 ( .A1(n5659), .A2(n5616), .ZN(n5621) );
  NAND2_X1 U7120 ( .A1(n5621), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5617) );
  XNOR2_X1 U7121 ( .A(n5617), .B(P1_IR_REG_11__SCAN_IN), .ZN(n9536) );
  INV_X1 U7122 ( .A(n9536), .ZN(n6803) );
  OAI22_X1 U7123 ( .A1(n5665), .A2(n6372), .B1(n5567), .B2(n6803), .ZN(n5618)
         );
  INV_X1 U7124 ( .A(n5618), .ZN(n5619) );
  NAND2_X1 U7125 ( .A1(n6422), .A2(n5696), .ZN(n5629) );
  NAND2_X1 U7126 ( .A1(n5624), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5623) );
  MUX2_X1 U7127 ( .A(n5623), .B(P1_IR_REG_31__SCAN_IN), .S(n5622), .Z(n5626)
         );
  INV_X1 U7128 ( .A(n5635), .ZN(n5625) );
  INV_X1 U7129 ( .A(n6936), .ZN(n6931) );
  OAI22_X1 U7130 ( .A1(n5665), .A2(n6423), .B1(n5567), .B2(n6931), .ZN(n5627)
         );
  INV_X1 U7131 ( .A(n5627), .ZN(n5628) );
  INV_X1 U7132 ( .A(n9460), .ZN(n7659) );
  NAND2_X1 U7133 ( .A1(n6485), .A2(n5696), .ZN(n5633) );
  OR2_X1 U7134 ( .A1(n5635), .A2(n9385), .ZN(n5630) );
  XNOR2_X1 U7135 ( .A(n5630), .B(P1_IR_REG_13__SCAN_IN), .ZN(n7084) );
  INV_X1 U7136 ( .A(n7084), .ZN(n7087) );
  OAI22_X1 U7137 ( .A1(n5665), .A2(n6486), .B1(n5567), .B2(n7087), .ZN(n5631)
         );
  INV_X1 U7138 ( .A(n5631), .ZN(n5632) );
  INV_X1 U7139 ( .A(n7723), .ZN(n9380) );
  NAND2_X1 U7140 ( .A1(n6481), .A2(n5696), .ZN(n5637) );
  NAND2_X1 U7141 ( .A1(n5635), .A2(n5634), .ZN(n5644) );
  NAND2_X1 U7142 ( .A1(n5644), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5639) );
  XNOR2_X1 U7143 ( .A(n5639), .B(P1_IR_REG_14__SCAN_IN), .ZN(n7088) );
  AOI22_X1 U7144 ( .A1(n5581), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n6288), .B2(
        n7088), .ZN(n5636) );
  NAND2_X1 U7145 ( .A1(n6553), .A2(n5696), .ZN(n5643) );
  NAND2_X1 U7146 ( .A1(n5639), .A2(n5638), .ZN(n5640) );
  NAND2_X1 U7147 ( .A1(n5640), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5641) );
  XNOR2_X1 U7148 ( .A(n5641), .B(P1_IR_REG_15__SCAN_IN), .ZN(n9555) );
  AOI22_X1 U7149 ( .A1(n5581), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n6288), .B2(
        n9555), .ZN(n5642) );
  NAND2_X1 U7150 ( .A1(n6513), .A2(n5696), .ZN(n5647) );
  NAND2_X1 U7151 ( .A1(n5648), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5645) );
  XNOR2_X1 U7152 ( .A(n5645), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9566) );
  AOI22_X1 U7153 ( .A1(n5581), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n6288), .B2(
        n9566), .ZN(n5646) );
  NAND2_X1 U7154 ( .A1(n6601), .A2(n5696), .ZN(n5653) );
  OAI21_X1 U7155 ( .B1(n5648), .B2(P1_IR_REG_16__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5650) );
  INV_X1 U7156 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5649) );
  NAND2_X1 U7157 ( .A1(n5650), .A2(n5649), .ZN(n5654) );
  OR2_X1 U7158 ( .A1(n5650), .A2(n5649), .ZN(n5651) );
  AOI22_X1 U7159 ( .A1(n5581), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n8975), .B2(
        n6288), .ZN(n5652) );
  INV_X1 U7160 ( .A(n9320), .ZN(n9191) );
  NAND2_X1 U7161 ( .A1(n9203), .A2(n9191), .ZN(n9179) );
  NAND2_X1 U7162 ( .A1(n6749), .A2(n5696), .ZN(n5657) );
  NAND2_X1 U7163 ( .A1(n5654), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5655) );
  XNOR2_X1 U7164 ( .A(n5655), .B(P1_IR_REG_18__SCAN_IN), .ZN(n8979) );
  AOI22_X1 U7165 ( .A1(n8979), .A2(n6288), .B1(n5581), .B2(
        P2_DATAO_REG_18__SCAN_IN), .ZN(n5656) );
  NAND2_X1 U7166 ( .A1(n6779), .A2(n5696), .ZN(n5668) );
  NAND2_X1 U7167 ( .A1(n5659), .A2(n5658), .ZN(n5661) );
  NAND2_X1 U7168 ( .A1(n5661), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5660) );
  MUX2_X1 U7169 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5660), .S(
        P1_IR_REG_19__SCAN_IN), .Z(n5664) );
  NAND2_X1 U7170 ( .A1(n5664), .A2(n5699), .ZN(n8985) );
  OAI22_X1 U7171 ( .A1(n5665), .A2(n6782), .B1(n8985), .B2(n5567), .ZN(n5666)
         );
  INV_X1 U7172 ( .A(n5666), .ZN(n5667) );
  NAND2_X1 U7173 ( .A1(n6870), .A2(n5696), .ZN(n5670) );
  NAND2_X1 U7174 ( .A1(n5581), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n5669) );
  INV_X1 U7175 ( .A(n9141), .ZN(n9367) );
  NAND2_X1 U7176 ( .A1(n6944), .A2(n5696), .ZN(n5672) );
  NAND2_X1 U7177 ( .A1(n5581), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n5671) );
  INV_X1 U7178 ( .A(n9296), .ZN(n9125) );
  NAND2_X1 U7179 ( .A1(n6992), .A2(n5696), .ZN(n5674) );
  NAND2_X1 U7180 ( .A1(n5581), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n5673) );
  NAND2_X1 U7181 ( .A1(n7097), .A2(n5696), .ZN(n5676) );
  NAND2_X1 U7182 ( .A1(n5581), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n5675) );
  NAND2_X1 U7183 ( .A1(n7218), .A2(n5696), .ZN(n5678) );
  NAND2_X1 U7184 ( .A1(n5581), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n5677) );
  INV_X1 U7185 ( .A(n9278), .ZN(n9085) );
  NAND2_X1 U7186 ( .A1(n7397), .A2(n5696), .ZN(n5680) );
  NAND2_X1 U7187 ( .A1(n5581), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n5679) );
  NAND2_X1 U7188 ( .A1(n7384), .A2(n5696), .ZN(n5682) );
  NAND2_X1 U7189 ( .A1(n5581), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n5681) );
  NAND2_X1 U7190 ( .A1(n7519), .A2(n5696), .ZN(n5684) );
  NAND2_X1 U7191 ( .A1(n5581), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n5683) );
  NAND2_X1 U7192 ( .A1(n7545), .A2(n5696), .ZN(n5686) );
  NAND2_X1 U7193 ( .A1(n5581), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n5685) );
  NAND2_X1 U7194 ( .A1(n7673), .A2(n5696), .ZN(n5688) );
  NAND2_X1 U7195 ( .A1(n5581), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n5687) );
  NAND2_X1 U7196 ( .A1(n9345), .A2(n8996), .ZN(n8997) );
  NAND2_X1 U7197 ( .A1(n5691), .A2(n5690), .ZN(n5692) );
  MUX2_X1 U7198 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n6327), .Z(n5693) );
  XNOR2_X1 U7199 ( .A(n5693), .B(SI_31_), .ZN(n5694) );
  NAND2_X1 U7200 ( .A1(n5581), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n5697) );
  INV_X1 U7201 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5707) );
  NAND2_X1 U7202 ( .A1(n5706), .A2(n5707), .ZN(n5700) );
  INV_X1 U7203 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5701) );
  NAND2_X1 U7204 ( .A1(n5705), .A2(n5701), .ZN(n5702) );
  INV_X1 U7205 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5703) );
  XNOR2_X1 U7206 ( .A(n5705), .B(P1_IR_REG_21__SCAN_IN), .ZN(n5777) );
  NAND2_X1 U7207 ( .A1(n4299), .A2(n8197), .ZN(n9633) );
  INV_X1 U7208 ( .A(n8201), .ZN(n7047) );
  NOR2_X1 U7209 ( .A1(n8082), .A2(n5755), .ZN(n5716) );
  INV_X1 U7210 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n5712) );
  NOR2_X1 U7211 ( .A1(n8084), .A2(n5712), .ZN(n5715) );
  INV_X1 U7212 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n5713) );
  NOR2_X1 U7213 ( .A1(n8088), .A2(n5713), .ZN(n5714) );
  OR3_X1 U7214 ( .A1(n5716), .A2(n5715), .A3(n5714), .ZN(n8097) );
  INV_X1 U7215 ( .A(n5717), .ZN(n5780) );
  NAND2_X1 U7216 ( .A1(n5780), .A2(n8206), .ZN(n8098) );
  NOR2_X2 U7217 ( .A1(n8098), .A2(n4568), .ZN(n9686) );
  INV_X1 U7218 ( .A(P1_B_REG_SCAN_IN), .ZN(n5720) );
  OR2_X1 U7219 ( .A1(n9479), .A2(n5720), .ZN(n5721) );
  AND2_X1 U7220 ( .A1(n9686), .A2(n5721), .ZN(n8325) );
  AND2_X1 U7221 ( .A1(n8097), .A2(n8325), .ZN(n9244) );
  NOR2_X1 U7222 ( .A1(n8991), .A2(n9244), .ZN(n5765) );
  NAND2_X1 U7223 ( .A1(n5722), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5725) );
  NAND2_X1 U7224 ( .A1(n5725), .A2(n5723), .ZN(n5727) );
  NAND2_X1 U7225 ( .A1(n5727), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5724) );
  INV_X1 U7226 ( .A(n5725), .ZN(n5726) );
  NAND2_X1 U7227 ( .A1(n5726), .A2(P1_IR_REG_25__SCAN_IN), .ZN(n5728) );
  NAND2_X1 U7228 ( .A1(n5728), .A2(n5727), .ZN(n7398) );
  NAND2_X1 U7229 ( .A1(n5729), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5730) );
  XNOR2_X1 U7230 ( .A(n5730), .B(n5554), .ZN(n7222) );
  NOR2_X1 U7231 ( .A1(n7398), .A2(n7222), .ZN(n5731) );
  NAND2_X1 U7232 ( .A1(n7385), .A2(n5731), .ZN(n6286) );
  NAND2_X1 U7233 ( .A1(n4382), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5733) );
  XNOR2_X1 U7234 ( .A(n5733), .B(n5732), .ZN(n7098) );
  AND2_X1 U7235 ( .A1(n6286), .A2(n7098), .ZN(n6235) );
  OR2_X1 U7236 ( .A1(n8098), .A2(n8243), .ZN(n6236) );
  NAND2_X1 U7237 ( .A1(n9654), .A2(n6236), .ZN(n7056) );
  INV_X1 U7238 ( .A(n9633), .ZN(n9639) );
  INV_X1 U7239 ( .A(n8985), .ZN(n9127) );
  NAND3_X1 U7240 ( .A1(n7398), .A2(P1_B_REG_SCAN_IN), .A3(n7222), .ZN(n5735)
         );
  OR2_X1 U7241 ( .A1(n7222), .A2(P1_B_REG_SCAN_IN), .ZN(n5734) );
  AND2_X1 U7242 ( .A1(n5735), .A2(n5734), .ZN(n5736) );
  NAND2_X1 U7243 ( .A1(n5736), .A2(n7385), .ZN(n9381) );
  OR2_X1 U7244 ( .A1(n9381), .A2(P1_D_REG_1__SCAN_IN), .ZN(n5739) );
  INV_X1 U7245 ( .A(n7398), .ZN(n5737) );
  OR2_X1 U7246 ( .A1(n7385), .A2(n5737), .ZN(n5738) );
  INV_X1 U7247 ( .A(n7054), .ZN(n5763) );
  NOR4_X1 U7248 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n5743) );
  NOR4_X1 U7249 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n5742) );
  NOR4_X1 U7250 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5741) );
  NOR4_X1 U7251 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n5740) );
  AND4_X1 U7252 ( .A1(n5743), .A2(n5742), .A3(n5741), .A4(n5740), .ZN(n5749)
         );
  NOR2_X1 U7253 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .ZN(
        n5747) );
  NOR4_X1 U7254 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_11__SCAN_IN), .A4(P1_D_REG_14__SCAN_IN), .ZN(n5746) );
  NOR4_X1 U7255 ( .A1(P1_D_REG_5__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n5745) );
  NOR4_X1 U7256 ( .A1(P1_D_REG_13__SCAN_IN), .A2(P1_D_REG_2__SCAN_IN), .A3(
        P1_D_REG_3__SCAN_IN), .A4(P1_D_REG_4__SCAN_IN), .ZN(n5744) );
  AND4_X1 U7257 ( .A1(n5747), .A2(n5746), .A3(n5745), .A4(n5744), .ZN(n5748)
         );
  NAND2_X1 U7258 ( .A1(n5749), .A2(n5748), .ZN(n5759) );
  INV_X1 U7259 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n5750) );
  NOR2_X1 U7260 ( .A1(n5759), .A2(n5750), .ZN(n5751) );
  OR2_X1 U7261 ( .A1(n9381), .A2(n5751), .ZN(n5753) );
  INV_X1 U7262 ( .A(n7222), .ZN(n5752) );
  OR2_X1 U7263 ( .A1(n7385), .A2(n5752), .ZN(n9382) );
  NAND2_X1 U7264 ( .A1(n5763), .A2(n6232), .ZN(n5754) );
  INV_X2 U7265 ( .A(n9731), .ZN(n9733) );
  NAND2_X1 U7266 ( .A1(n9733), .A2(n9695), .ZN(n9342) );
  NAND2_X1 U7267 ( .A1(n5698), .A2(n5756), .ZN(n5757) );
  NAND2_X1 U7268 ( .A1(n5758), .A2(n5757), .ZN(P1_U3554) );
  OAI21_X1 U7269 ( .B1(n9381), .B2(P1_D_REG_0__SCAN_IN), .A(n9382), .ZN(n5762)
         );
  INV_X1 U7270 ( .A(n5759), .ZN(n5760) );
  OR2_X1 U7271 ( .A1(n9381), .A2(n5760), .ZN(n5761) );
  AND2_X1 U7272 ( .A1(n5762), .A2(n5761), .ZN(n7055) );
  NAND2_X1 U7273 ( .A1(n5763), .A2(n7055), .ZN(n5764) );
  INV_X2 U7274 ( .A(n9718), .ZN(n9720) );
  NAND2_X1 U7275 ( .A1(n9720), .A2(n9695), .ZN(n9379) );
  NAND2_X1 U7276 ( .A1(n5698), .A2(n5766), .ZN(n5767) );
  NAND2_X1 U7277 ( .A1(n5768), .A2(n5767), .ZN(P1_U3522) );
  INV_X1 U7278 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n5776) );
  INV_X1 U7279 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n5769) );
  INV_X1 U7280 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9721) );
  OR2_X1 U7281 ( .A1(n5799), .A2(n9721), .ZN(n5773) );
  NAND2_X1 U7282 ( .A1(n5845), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5772) );
  AND2_X1 U7283 ( .A1(n5773), .A2(n5772), .ZN(n5774) );
  INV_X1 U7284 ( .A(n6222), .ZN(n7041) );
  INV_X2 U7285 ( .A(n4320), .ZN(n5903) );
  NAND2_X1 U7286 ( .A1(n6638), .A2(n5903), .ZN(n5779) );
  INV_X1 U7287 ( .A(n6286), .ZN(n5782) );
  AOI22_X1 U7288 ( .A1(n9640), .A2(n6262), .B1(P1_REG1_REG_0__SCAN_IN), .B2(
        n5782), .ZN(n5778) );
  NAND2_X1 U7289 ( .A1(n5779), .A2(n5778), .ZN(n6515) );
  INV_X1 U7290 ( .A(n6515), .ZN(n5781) );
  NAND2_X1 U7291 ( .A1(n5781), .A2(n4298), .ZN(n5785) );
  NAND2_X1 U7292 ( .A1(n4299), .A2(n8243), .ZN(n7043) );
  AND2_X4 U7293 ( .A1(n5806), .A2(n7043), .ZN(n6257) );
  NAND2_X1 U7294 ( .A1(n6638), .A2(n6257), .ZN(n5784) );
  AOI22_X1 U7295 ( .A1(n9640), .A2(n5903), .B1(P1_IR_REG_0__SCAN_IN), .B2(
        n5782), .ZN(n5783) );
  AND2_X1 U7296 ( .A1(n5784), .A2(n5783), .ZN(n6517) );
  NAND2_X1 U7297 ( .A1(n6517), .A2(n6515), .ZN(n6516) );
  NAND2_X1 U7298 ( .A1(n5785), .A2(n6516), .ZN(n5798) );
  INV_X1 U7299 ( .A(n5798), .ZN(n5796) );
  NAND2_X1 U7300 ( .A1(n5803), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5791) );
  INV_X1 U7301 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n5786) );
  OR2_X1 U7302 ( .A1(n4290), .A2(n5786), .ZN(n5790) );
  NAND2_X1 U7303 ( .A1(n5845), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5788) );
  INV_X1 U7304 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6305) );
  NAND2_X1 U7305 ( .A1(n7040), .A2(n5903), .ZN(n5793) );
  NAND2_X1 U7306 ( .A1(n7038), .A2(n6262), .ZN(n5792) );
  NAND2_X1 U7307 ( .A1(n5793), .A2(n5792), .ZN(n5794) );
  XNOR2_X1 U7308 ( .A(n5794), .B(n4297), .ZN(n5797) );
  INV_X1 U7309 ( .A(n5797), .ZN(n5795) );
  AOI22_X1 U7310 ( .A1(n7040), .A2(n6257), .B1(n6261), .B2(n7038), .ZN(n6636)
         );
  NAND2_X1 U7311 ( .A1(n6635), .A2(n6636), .ZN(n6634) );
  NAND2_X1 U7312 ( .A1(n5798), .A2(n5797), .ZN(n6753) );
  NAND2_X1 U7313 ( .A1(n6634), .A2(n6753), .ZN(n5813) );
  INV_X1 U7314 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n9724) );
  OR2_X1 U7315 ( .A1(n5799), .A2(n9724), .ZN(n5800) );
  INV_X1 U7316 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n5802) );
  NAND2_X1 U7317 ( .A1(n9660), .A2(n6139), .ZN(n5808) );
  NAND2_X1 U7318 ( .A1(n5808), .A2(n5807), .ZN(n5809) );
  XNOR2_X1 U7319 ( .A(n5809), .B(n4297), .ZN(n5810) );
  NAND2_X1 U7320 ( .A1(n5810), .A2(n5811), .ZN(n5814) );
  OAI21_X1 U7321 ( .B1(n5811), .B2(n5810), .A(n5814), .ZN(n5812) );
  INV_X1 U7322 ( .A(n5812), .ZN(n6755) );
  NAND2_X1 U7323 ( .A1(n5813), .A2(n6755), .ZN(n6757) );
  NAND2_X1 U7324 ( .A1(n6757), .A2(n5814), .ZN(n6813) );
  INV_X1 U7325 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n5815) );
  INV_X1 U7326 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n5816) );
  INV_X1 U7327 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6304) );
  OR2_X1 U7328 ( .A1(n5799), .A2(n6304), .ZN(n5817) );
  NAND2_X1 U7329 ( .A1(n5862), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5820) );
  NAND2_X1 U7330 ( .A1(n6792), .A2(n5903), .ZN(n5822) );
  NAND2_X1 U7331 ( .A1(n9667), .A2(n6262), .ZN(n5821) );
  NAND2_X1 U7332 ( .A1(n5822), .A2(n5821), .ZN(n5823) );
  XNOR2_X1 U7333 ( .A(n5823), .B(n4298), .ZN(n5836) );
  AOI22_X1 U7334 ( .A1(n6792), .A2(n6257), .B1(n6261), .B2(n9667), .ZN(n5837)
         );
  XNOR2_X1 U7335 ( .A(n5836), .B(n5837), .ZN(n6814) );
  NAND2_X1 U7336 ( .A1(n6813), .A2(n6814), .ZN(n6786) );
  INV_X1 U7337 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n5824) );
  OR2_X1 U7338 ( .A1(n5799), .A2(n5824), .ZN(n5832) );
  INV_X1 U7339 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n5825) );
  NAND2_X1 U7340 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5848) );
  OAI21_X1 U7341 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(n5848), .ZN(n6791) );
  OR2_X1 U7342 ( .A1(n5827), .A2(n6791), .ZN(n5830) );
  INV_X1 U7343 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n5828) );
  OR2_X1 U7344 ( .A1(n4290), .A2(n5828), .ZN(n5829) );
  NAND2_X1 U7345 ( .A1(n9668), .A2(n5903), .ZN(n5834) );
  NAND2_X1 U7346 ( .A1(n9623), .A2(n6262), .ZN(n5833) );
  NAND2_X1 U7347 ( .A1(n5834), .A2(n5833), .ZN(n5835) );
  AOI22_X1 U7348 ( .A1(n9668), .A2(n6257), .B1(n6261), .B2(n9623), .ZN(n5841)
         );
  XNOR2_X1 U7349 ( .A(n5840), .B(n5841), .ZN(n6789) );
  INV_X1 U7350 ( .A(n5836), .ZN(n5838) );
  NAND2_X1 U7351 ( .A1(n5838), .A2(n5837), .ZN(n6787) );
  NAND2_X1 U7352 ( .A1(n6786), .A2(n5839), .ZN(n6788) );
  INV_X1 U7353 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n5844) );
  OR2_X1 U7354 ( .A1(n4290), .A2(n5844), .ZN(n5854) );
  INV_X1 U7355 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6303) );
  INV_X1 U7356 ( .A(n5848), .ZN(n5846) );
  NAND2_X1 U7357 ( .A1(n5846), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5880) );
  INV_X1 U7358 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5847) );
  NAND2_X1 U7359 ( .A1(n5848), .A2(n5847), .ZN(n5849) );
  NAND2_X1 U7360 ( .A1(n5880), .A2(n5849), .ZN(n7019) );
  OR2_X1 U7361 ( .A1(n5827), .A2(n7019), .ZN(n5852) );
  INV_X1 U7362 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n5850) );
  OR2_X1 U7363 ( .A1(n8088), .A2(n5850), .ZN(n5851) );
  NAND2_X1 U7364 ( .A1(n9614), .A2(n5903), .ZN(n5856) );
  NAND2_X1 U7365 ( .A1(n9685), .A2(n6139), .ZN(n5855) );
  NAND2_X1 U7366 ( .A1(n5856), .A2(n5855), .ZN(n5857) );
  XNOR2_X1 U7367 ( .A(n5857), .B(n4298), .ZN(n5859) );
  INV_X1 U7368 ( .A(n5859), .ZN(n5858) );
  NAND2_X1 U7369 ( .A1(n5860), .A2(n5859), .ZN(n5861) );
  AOI22_X1 U7370 ( .A1(n9614), .A2(n6257), .B1(n6261), .B2(n9685), .ZN(n7017)
         );
  NAND2_X1 U7371 ( .A1(n7016), .A2(n7017), .ZN(n7015) );
  NAND2_X1 U7372 ( .A1(n5862), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5867) );
  INV_X1 U7373 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n5863) );
  OR2_X1 U7374 ( .A1(n8082), .A2(n5863), .ZN(n5866) );
  INV_X1 U7375 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n5879) );
  XNOR2_X1 U7376 ( .A(n5880), .B(n5879), .ZN(n7313) );
  OR2_X1 U7377 ( .A1(n5827), .A2(n7313), .ZN(n5865) );
  INV_X1 U7378 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n7310) );
  OR2_X1 U7379 ( .A1(n8088), .A2(n7310), .ZN(n5864) );
  NAND4_X1 U7380 ( .A1(n5867), .A2(n5866), .A3(n5865), .A4(n5864), .ZN(n9687)
         );
  NAND2_X1 U7381 ( .A1(n9687), .A2(n5903), .ZN(n5869) );
  NAND2_X1 U7382 ( .A1(n9694), .A2(n6139), .ZN(n5868) );
  NAND2_X1 U7383 ( .A1(n5869), .A2(n5868), .ZN(n5870) );
  XNOR2_X1 U7384 ( .A(n5870), .B(n4297), .ZN(n5872) );
  AOI22_X1 U7385 ( .A1(n9687), .A2(n6257), .B1(n6261), .B2(n9694), .ZN(n5873)
         );
  AND2_X1 U7386 ( .A1(n4324), .A2(n7025), .ZN(n5871) );
  NAND2_X1 U7387 ( .A1(n7015), .A2(n5871), .ZN(n5876) );
  INV_X1 U7388 ( .A(n5872), .ZN(n5875) );
  INV_X1 U7389 ( .A(n5873), .ZN(n5874) );
  NAND2_X1 U7390 ( .A1(n5875), .A2(n5874), .ZN(n7027) );
  NAND2_X1 U7391 ( .A1(n5862), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5888) );
  INV_X1 U7392 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n5877) );
  OR2_X1 U7393 ( .A1(n8082), .A2(n5877), .ZN(n5887) );
  INV_X1 U7394 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5878) );
  OAI21_X1 U7395 ( .B1(n5880), .B2(n5879), .A(n5878), .ZN(n5883) );
  INV_X1 U7396 ( .A(n5880), .ZN(n5882) );
  NAND2_X1 U7397 ( .A1(n5882), .A2(n5881), .ZN(n5896) );
  NAND2_X1 U7398 ( .A1(n5883), .A2(n5896), .ZN(n7115) );
  OR2_X1 U7399 ( .A1(n5827), .A2(n7115), .ZN(n5886) );
  INV_X1 U7400 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n5884) );
  OR2_X1 U7401 ( .A1(n8088), .A2(n5884), .ZN(n5885) );
  NAND4_X1 U7402 ( .A1(n5888), .A2(n5887), .A3(n5886), .A4(n5885), .ZN(n8955)
         );
  NAND2_X1 U7403 ( .A1(n8955), .A2(n6257), .ZN(n5890) );
  NAND2_X1 U7404 ( .A1(n7174), .A2(n5903), .ZN(n5889) );
  NAND2_X1 U7405 ( .A1(n5890), .A2(n5889), .ZN(n7112) );
  NAND2_X1 U7406 ( .A1(n8955), .A2(n6261), .ZN(n5892) );
  NAND2_X1 U7407 ( .A1(n7174), .A2(n6139), .ZN(n5891) );
  NAND2_X1 U7408 ( .A1(n5892), .A2(n5891), .ZN(n5893) );
  XNOR2_X1 U7409 ( .A(n5893), .B(n4298), .ZN(n7111) );
  NAND2_X1 U7410 ( .A1(n5862), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5902) );
  INV_X1 U7411 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6302) );
  OR2_X1 U7412 ( .A1(n8082), .A2(n6302), .ZN(n5901) );
  INV_X1 U7413 ( .A(n5896), .ZN(n5894) );
  NAND2_X1 U7414 ( .A1(n5894), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5910) );
  INV_X1 U7415 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n5895) );
  NAND2_X1 U7416 ( .A1(n5896), .A2(n5895), .ZN(n5897) );
  NAND2_X1 U7417 ( .A1(n5910), .A2(n5897), .ZN(n7243) );
  OR2_X1 U7418 ( .A1(n5827), .A2(n7243), .ZN(n5900) );
  INV_X1 U7419 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n5898) );
  OR2_X1 U7420 ( .A1(n8088), .A2(n5898), .ZN(n5899) );
  NAND4_X1 U7421 ( .A1(n5902), .A2(n5901), .A3(n5900), .A4(n5899), .ZN(n8954)
         );
  NAND2_X1 U7422 ( .A1(n8954), .A2(n6257), .ZN(n5905) );
  NAND2_X1 U7423 ( .A1(n7299), .A2(n5903), .ZN(n5904) );
  NAND2_X1 U7424 ( .A1(n5905), .A2(n5904), .ZN(n7238) );
  NAND2_X1 U7425 ( .A1(n8954), .A2(n6261), .ZN(n5907) );
  NAND2_X1 U7426 ( .A1(n7299), .A2(n6139), .ZN(n5906) );
  NAND2_X1 U7427 ( .A1(n5907), .A2(n5906), .ZN(n5908) );
  XNOR2_X1 U7428 ( .A(n5908), .B(n4298), .ZN(n7237) );
  NAND2_X1 U7429 ( .A1(n7468), .A2(n6139), .ZN(n5919) );
  NAND2_X1 U7430 ( .A1(n5803), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5917) );
  INV_X1 U7431 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5909) );
  NAND2_X1 U7432 ( .A1(n5910), .A2(n5909), .ZN(n5911) );
  NAND2_X1 U7433 ( .A1(n5962), .A2(n5911), .ZN(n7466) );
  OR2_X1 U7434 ( .A1(n5827), .A2(n7466), .ZN(n5916) );
  INV_X1 U7435 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n5912) );
  OR2_X1 U7436 ( .A1(n8082), .A2(n5912), .ZN(n5915) );
  INV_X1 U7437 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n5913) );
  OR2_X1 U7438 ( .A1(n4290), .A2(n5913), .ZN(n5914) );
  NAND4_X1 U7439 ( .A1(n5917), .A2(n5916), .A3(n5915), .A4(n5914), .ZN(n8953)
         );
  NAND2_X1 U7440 ( .A1(n8953), .A2(n6261), .ZN(n5918) );
  NAND2_X1 U7441 ( .A1(n5919), .A2(n5918), .ZN(n5920) );
  XNOR2_X1 U7442 ( .A(n5920), .B(n4297), .ZN(n5923) );
  NAND2_X1 U7443 ( .A1(n7468), .A2(n6261), .ZN(n5922) );
  NAND2_X1 U7444 ( .A1(n8953), .A2(n6257), .ZN(n5921) );
  AND2_X1 U7445 ( .A1(n5922), .A2(n5921), .ZN(n5924) );
  NAND2_X1 U7446 ( .A1(n5923), .A2(n5924), .ZN(n7489) );
  INV_X1 U7447 ( .A(n5923), .ZN(n5926) );
  INV_X1 U7448 ( .A(n5924), .ZN(n5925) );
  NAND2_X1 U7449 ( .A1(n5926), .A2(n5925), .ZN(n5927) );
  NAND2_X1 U7450 ( .A1(n7489), .A2(n5927), .ZN(n7462) );
  NAND2_X1 U7451 ( .A1(n9460), .A2(n6139), .ZN(n5939) );
  NAND2_X1 U7452 ( .A1(n5803), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5937) );
  INV_X1 U7453 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n5928) );
  OR2_X1 U7454 ( .A1(n8082), .A2(n5928), .ZN(n5936) );
  NAND2_X1 U7455 ( .A1(n5929), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5964) );
  INV_X1 U7456 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5944) );
  INV_X1 U7457 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5931) );
  NAND2_X1 U7458 ( .A1(n5946), .A2(n5931), .ZN(n5932) );
  NAND2_X1 U7459 ( .A1(n5988), .A2(n5932), .ZN(n7655) );
  OR2_X1 U7460 ( .A1(n5827), .A2(n7655), .ZN(n5935) );
  INV_X1 U7461 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n5933) );
  OR2_X1 U7462 ( .A1(n4290), .A2(n5933), .ZN(n5934) );
  NAND4_X1 U7463 ( .A1(n5937), .A2(n5936), .A3(n5935), .A4(n5934), .ZN(n8950)
         );
  NAND2_X1 U7464 ( .A1(n8950), .A2(n6261), .ZN(n5938) );
  NAND2_X1 U7465 ( .A1(n5939), .A2(n5938), .ZN(n5940) );
  XNOR2_X1 U7466 ( .A(n5940), .B(n4297), .ZN(n5943) );
  AND2_X1 U7467 ( .A1(n8950), .A2(n6257), .ZN(n5941) );
  AOI21_X1 U7468 ( .B1(n9460), .B2(n6261), .A(n5941), .ZN(n5942) );
  NAND2_X1 U7469 ( .A1(n5943), .A2(n5942), .ZN(n5982) );
  INV_X1 U7470 ( .A(n5982), .ZN(n5976) );
  XNOR2_X1 U7471 ( .A(n5943), .B(n5942), .ZN(n7538) );
  INV_X1 U7472 ( .A(n7538), .ZN(n5975) );
  NAND2_X1 U7473 ( .A1(n7645), .A2(n6139), .ZN(n5953) );
  NAND2_X1 U7474 ( .A1(n5862), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5951) );
  INV_X1 U7475 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n6799) );
  OR2_X1 U7476 ( .A1(n8082), .A2(n6799), .ZN(n5950) );
  NAND2_X1 U7477 ( .A1(n5964), .A2(n5944), .ZN(n5945) );
  NAND2_X1 U7478 ( .A1(n5946), .A2(n5945), .ZN(n7591) );
  OR2_X1 U7479 ( .A1(n5827), .A2(n7591), .ZN(n5949) );
  INV_X1 U7480 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n5947) );
  OR2_X1 U7481 ( .A1(n8088), .A2(n5947), .ZN(n5948) );
  NAND4_X1 U7482 ( .A1(n5951), .A2(n5950), .A3(n5949), .A4(n5948), .ZN(n8951)
         );
  NAND2_X1 U7483 ( .A1(n8951), .A2(n6261), .ZN(n5952) );
  NAND2_X1 U7484 ( .A1(n5953), .A2(n5952), .ZN(n5954) );
  XNOR2_X1 U7485 ( .A(n5954), .B(n4297), .ZN(n5959) );
  INV_X1 U7486 ( .A(n5959), .ZN(n5957) );
  AND2_X1 U7487 ( .A1(n8951), .A2(n6257), .ZN(n5955) );
  AOI21_X1 U7488 ( .B1(n7645), .B2(n6261), .A(n5955), .ZN(n5958) );
  INV_X1 U7489 ( .A(n5958), .ZN(n5956) );
  NAND2_X1 U7490 ( .A1(n5957), .A2(n5956), .ZN(n5974) );
  XNOR2_X1 U7491 ( .A(n5959), .B(n5958), .ZN(n7585) );
  NAND2_X1 U7492 ( .A1(n7500), .A2(n6139), .ZN(n5970) );
  NAND2_X1 U7493 ( .A1(n6202), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5968) );
  INV_X1 U7494 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n5960) );
  OR2_X1 U7495 ( .A1(n4290), .A2(n5960), .ZN(n5967) );
  INV_X1 U7496 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n5961) );
  NAND2_X1 U7497 ( .A1(n5962), .A2(n5961), .ZN(n5963) );
  NAND2_X1 U7498 ( .A1(n5964), .A2(n5963), .ZN(n7498) );
  OR2_X1 U7499 ( .A1(n5827), .A2(n7498), .ZN(n5966) );
  INV_X1 U7500 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7480) );
  OR2_X1 U7501 ( .A1(n8088), .A2(n7480), .ZN(n5965) );
  NAND2_X1 U7502 ( .A1(n8952), .A2(n6261), .ZN(n5969) );
  NAND2_X1 U7503 ( .A1(n5970), .A2(n5969), .ZN(n5971) );
  NAND2_X1 U7504 ( .A1(n7500), .A2(n6261), .ZN(n5973) );
  NAND2_X1 U7505 ( .A1(n8952), .A2(n6257), .ZN(n5972) );
  NAND2_X1 U7506 ( .A1(n5973), .A2(n5972), .ZN(n5978) );
  NAND2_X1 U7507 ( .A1(n5977), .A2(n5978), .ZN(n7583) );
  OR2_X1 U7508 ( .A1(n7585), .A2(n7583), .ZN(n7587) );
  AND2_X1 U7509 ( .A1(n5974), .A2(n7587), .ZN(n7534) );
  OR2_X1 U7510 ( .A1(n7462), .A2(n5984), .ZN(n5986) );
  INV_X1 U7511 ( .A(n5977), .ZN(n5980) );
  INV_X1 U7512 ( .A(n5978), .ZN(n5979) );
  NAND2_X1 U7513 ( .A1(n5980), .A2(n5979), .ZN(n7490) );
  AND2_X1 U7514 ( .A1(n7489), .A2(n7490), .ZN(n7581) );
  INV_X1 U7515 ( .A(n7585), .ZN(n5981) );
  AND2_X1 U7516 ( .A1(n7581), .A2(n5981), .ZN(n7533) );
  AND2_X1 U7517 ( .A1(n7533), .A2(n5982), .ZN(n5983) );
  OR2_X1 U7518 ( .A1(n5984), .A2(n5983), .ZN(n5985) );
  NAND2_X1 U7519 ( .A1(n7723), .A2(n6139), .ZN(n5996) );
  NAND2_X1 U7520 ( .A1(n6202), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5994) );
  INV_X1 U7521 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7725) );
  OR2_X1 U7522 ( .A1(n8088), .A2(n7725), .ZN(n5993) );
  INV_X1 U7523 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5987) );
  NAND2_X1 U7524 ( .A1(n5988), .A2(n5987), .ZN(n5989) );
  NAND2_X1 U7525 ( .A1(n6002), .A2(n5989), .ZN(n7724) );
  OR2_X1 U7526 ( .A1(n5827), .A2(n7724), .ZN(n5992) );
  INV_X1 U7527 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n5990) );
  OR2_X1 U7528 ( .A1(n4290), .A2(n5990), .ZN(n5991) );
  NAND4_X1 U7529 ( .A1(n5994), .A2(n5993), .A3(n5992), .A4(n5991), .ZN(n9459)
         );
  NAND2_X1 U7530 ( .A1(n9459), .A2(n6261), .ZN(n5995) );
  NAND2_X1 U7531 ( .A1(n5996), .A2(n5995), .ZN(n5997) );
  XNOR2_X1 U7532 ( .A(n5997), .B(n4297), .ZN(n7525) );
  AND2_X1 U7533 ( .A1(n9459), .A2(n6257), .ZN(n5998) );
  AOI21_X1 U7534 ( .B1(n7723), .B2(n6261), .A(n5998), .ZN(n7524) );
  AND2_X1 U7535 ( .A1(n7525), .A2(n7524), .ZN(n6000) );
  OAI21_X1 U7536 ( .B1(n7523), .B2(n6000), .A(n5999), .ZN(n7613) );
  NAND2_X1 U7537 ( .A1(n8257), .A2(n6139), .ZN(n6009) );
  NAND2_X1 U7538 ( .A1(n5862), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n6007) );
  INV_X1 U7539 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n6001) );
  OR2_X1 U7540 ( .A1(n8082), .A2(n6001), .ZN(n6006) );
  INV_X1 U7541 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n10161) );
  NAND2_X1 U7542 ( .A1(n6002), .A2(n10161), .ZN(n6003) );
  NAND2_X1 U7543 ( .A1(n6030), .A2(n6003), .ZN(n7705) );
  OR2_X1 U7544 ( .A1(n5827), .A2(n7705), .ZN(n6005) );
  INV_X1 U7545 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7706) );
  OR2_X1 U7546 ( .A1(n8088), .A2(n7706), .ZN(n6004) );
  NAND4_X1 U7547 ( .A1(n6007), .A2(n6006), .A3(n6005), .A4(n6004), .ZN(n9225)
         );
  NAND2_X1 U7548 ( .A1(n9225), .A2(n6261), .ZN(n6008) );
  NAND2_X1 U7549 ( .A1(n6009), .A2(n6008), .ZN(n6010) );
  XNOR2_X1 U7550 ( .A(n6010), .B(n4297), .ZN(n7615) );
  AND2_X1 U7551 ( .A1(n9225), .A2(n6257), .ZN(n6011) );
  AOI21_X1 U7552 ( .B1(n8257), .B2(n5903), .A(n6011), .ZN(n6013) );
  NAND2_X1 U7553 ( .A1(n7615), .A2(n6013), .ZN(n6012) );
  NAND2_X1 U7554 ( .A1(n7613), .A2(n6012), .ZN(n6016) );
  INV_X1 U7555 ( .A(n7615), .ZN(n6014) );
  INV_X1 U7556 ( .A(n6013), .ZN(n7614) );
  NAND2_X1 U7557 ( .A1(n6014), .A2(n7614), .ZN(n6015) );
  NAND2_X1 U7558 ( .A1(n6016), .A2(n6015), .ZN(n7667) );
  NAND2_X1 U7559 ( .A1(n9328), .A2(n6261), .ZN(n6022) );
  NAND2_X1 U7560 ( .A1(n5803), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n6020) );
  INV_X1 U7561 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n10062) );
  OR2_X1 U7562 ( .A1(n4290), .A2(n10062), .ZN(n6019) );
  INV_X1 U7563 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9334) );
  OR2_X1 U7564 ( .A1(n8082), .A2(n9334), .ZN(n6018) );
  INV_X1 U7565 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n6029) );
  XNOR2_X1 U7566 ( .A(n6030), .B(n6029), .ZN(n9232) );
  OR2_X1 U7567 ( .A1(n5827), .A2(n9232), .ZN(n6017) );
  NAND4_X1 U7568 ( .A1(n6020), .A2(n6019), .A3(n6018), .A4(n6017), .ZN(n8949)
         );
  NAND2_X1 U7569 ( .A1(n8949), .A2(n6257), .ZN(n6021) );
  NAND2_X1 U7570 ( .A1(n6022), .A2(n6021), .ZN(n7665) );
  NAND2_X1 U7571 ( .A1(n9328), .A2(n6262), .ZN(n6024) );
  NAND2_X1 U7572 ( .A1(n8949), .A2(n6261), .ZN(n6023) );
  NAND2_X1 U7573 ( .A1(n6024), .A2(n6023), .ZN(n6025) );
  XNOR2_X1 U7574 ( .A(n6025), .B(n4298), .ZN(n7664) );
  NAND2_X1 U7575 ( .A1(n9325), .A2(n6262), .ZN(n6038) );
  NAND2_X1 U7576 ( .A1(n6202), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n6036) );
  INV_X1 U7577 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n9208) );
  OR2_X1 U7578 ( .A1(n8088), .A2(n9208), .ZN(n6035) );
  AND2_X1 U7579 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_REG3_REG_16__SCAN_IN), 
        .ZN(n6026) );
  INV_X1 U7580 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n6028) );
  OAI21_X1 U7581 ( .B1(n6030), .B2(n6029), .A(n6028), .ZN(n6031) );
  NAND2_X1 U7582 ( .A1(n6050), .A2(n6031), .ZN(n9207) );
  OR2_X1 U7583 ( .A1(n5827), .A2(n9207), .ZN(n6034) );
  INV_X1 U7584 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n6032) );
  OR2_X1 U7585 ( .A1(n8084), .A2(n6032), .ZN(n6033) );
  NAND4_X1 U7586 ( .A1(n6036), .A2(n6035), .A3(n6034), .A4(n6033), .ZN(n8948)
         );
  NAND2_X1 U7587 ( .A1(n8948), .A2(n6261), .ZN(n6037) );
  NAND2_X1 U7588 ( .A1(n6038), .A2(n6037), .ZN(n6039) );
  XNOR2_X1 U7589 ( .A(n6039), .B(n4297), .ZN(n6041) );
  AND2_X1 U7590 ( .A1(n8948), .A2(n6257), .ZN(n6040) );
  AOI21_X1 U7591 ( .B1(n9325), .B2(n6261), .A(n6040), .ZN(n6042) );
  NAND2_X1 U7592 ( .A1(n6041), .A2(n6042), .ZN(n6047) );
  INV_X1 U7593 ( .A(n6041), .ZN(n6044) );
  INV_X1 U7594 ( .A(n6042), .ZN(n6043) );
  NAND2_X1 U7595 ( .A1(n6044), .A2(n6043), .ZN(n6045) );
  NAND2_X1 U7596 ( .A1(n6047), .A2(n6045), .ZN(n8883) );
  NAND2_X1 U7597 ( .A1(n8881), .A2(n6047), .ZN(n8890) );
  NAND2_X1 U7598 ( .A1(n9320), .A2(n6262), .ZN(n6057) );
  NAND2_X1 U7599 ( .A1(n5862), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n6055) );
  INV_X1 U7600 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n8963) );
  OR2_X1 U7601 ( .A1(n8082), .A2(n8963), .ZN(n6054) );
  INV_X1 U7602 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n6049) );
  NAND2_X1 U7603 ( .A1(n6050), .A2(n6049), .ZN(n6051) );
  NAND2_X1 U7604 ( .A1(n6080), .A2(n6051), .ZN(n9192) );
  OR2_X1 U7605 ( .A1(n5827), .A2(n9192), .ZN(n6053) );
  INV_X1 U7606 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n9193) );
  OR2_X1 U7607 ( .A1(n8088), .A2(n9193), .ZN(n6052) );
  NAND4_X1 U7608 ( .A1(n6055), .A2(n6054), .A3(n6053), .A4(n6052), .ZN(n9169)
         );
  NAND2_X1 U7609 ( .A1(n9169), .A2(n6261), .ZN(n6056) );
  NAND2_X1 U7610 ( .A1(n6057), .A2(n6056), .ZN(n6058) );
  XNOR2_X1 U7611 ( .A(n6058), .B(n4298), .ZN(n6060) );
  AND2_X1 U7612 ( .A1(n9169), .A2(n6257), .ZN(n6059) );
  AOI21_X1 U7613 ( .B1(n9320), .B2(n6261), .A(n6059), .ZN(n6061) );
  XNOR2_X1 U7614 ( .A(n6060), .B(n6061), .ZN(n8892) );
  NAND2_X1 U7615 ( .A1(n8890), .A2(n8892), .ZN(n8891) );
  INV_X1 U7616 ( .A(n6060), .ZN(n6062) );
  NAND2_X1 U7617 ( .A1(n6062), .A2(n6061), .ZN(n6063) );
  NAND2_X1 U7618 ( .A1(n8891), .A2(n6063), .ZN(n6073) );
  NAND2_X1 U7619 ( .A1(n9313), .A2(n6262), .ZN(n6069) );
  NAND2_X1 U7620 ( .A1(n5862), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n6067) );
  INV_X1 U7621 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n8964) );
  OR2_X1 U7622 ( .A1(n8082), .A2(n8964), .ZN(n6066) );
  INV_X1 U7623 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n6078) );
  XNOR2_X1 U7624 ( .A(n6080), .B(n6078), .ZN(n9175) );
  OR2_X1 U7625 ( .A1(n5827), .A2(n9175), .ZN(n6065) );
  INV_X1 U7626 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n8976) );
  OR2_X1 U7627 ( .A1(n8088), .A2(n8976), .ZN(n6064) );
  NAND4_X1 U7628 ( .A1(n6067), .A2(n6066), .A3(n6065), .A4(n6064), .ZN(n8947)
         );
  NAND2_X1 U7629 ( .A1(n8947), .A2(n6261), .ZN(n6068) );
  NAND2_X1 U7630 ( .A1(n6069), .A2(n6068), .ZN(n6070) );
  XNOR2_X1 U7631 ( .A(n6070), .B(n4297), .ZN(n6074) );
  NAND2_X1 U7632 ( .A1(n6073), .A2(n6074), .ZN(n8932) );
  NAND2_X1 U7633 ( .A1(n9313), .A2(n6261), .ZN(n6072) );
  NAND2_X1 U7634 ( .A1(n8947), .A2(n6257), .ZN(n6071) );
  NAND2_X1 U7635 ( .A1(n6072), .A2(n6071), .ZN(n8935) );
  NAND2_X1 U7636 ( .A1(n9157), .A2(n6262), .ZN(n6087) );
  NAND2_X1 U7637 ( .A1(n5862), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n6085) );
  INV_X1 U7638 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9309) );
  OR2_X1 U7639 ( .A1(n8082), .A2(n9309), .ZN(n6084) );
  INV_X1 U7640 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n6077) );
  OAI21_X1 U7641 ( .B1(n6080), .B2(n6078), .A(n6077), .ZN(n6081) );
  NAND2_X1 U7642 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_REG3_REG_19__SCAN_IN), 
        .ZN(n6079) );
  NAND2_X1 U7643 ( .A1(n6081), .A2(n6098), .ZN(n9158) );
  OR2_X1 U7644 ( .A1(n5827), .A2(n9158), .ZN(n6083) );
  INV_X1 U7645 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n9159) );
  OR2_X1 U7646 ( .A1(n8088), .A2(n9159), .ZN(n6082) );
  NAND4_X1 U7647 ( .A1(n6085), .A2(n6084), .A3(n6083), .A4(n6082), .ZN(n9312)
         );
  NAND2_X1 U7648 ( .A1(n9312), .A2(n6261), .ZN(n6086) );
  NAND2_X1 U7649 ( .A1(n6087), .A2(n6086), .ZN(n6088) );
  XNOR2_X1 U7650 ( .A(n6088), .B(n4297), .ZN(n6090) );
  AND2_X1 U7651 ( .A1(n9312), .A2(n6257), .ZN(n6089) );
  AOI21_X1 U7652 ( .B1(n9157), .B2(n6261), .A(n6089), .ZN(n6091) );
  NAND2_X1 U7653 ( .A1(n6090), .A2(n6091), .ZN(n8915) );
  INV_X1 U7654 ( .A(n6090), .ZN(n6093) );
  INV_X1 U7655 ( .A(n6091), .ZN(n6092) );
  NAND2_X1 U7656 ( .A1(n6093), .A2(n6092), .ZN(n6094) );
  NAND2_X1 U7657 ( .A1(n8915), .A2(n6094), .ZN(n8856) );
  NAND2_X1 U7658 ( .A1(n8916), .A2(n8915), .ZN(n6113) );
  NAND2_X1 U7659 ( .A1(n9141), .A2(n6262), .ZN(n6105) );
  NAND2_X1 U7660 ( .A1(n5862), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n6103) );
  INV_X1 U7661 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n9304) );
  OR2_X1 U7662 ( .A1(n8082), .A2(n9304), .ZN(n6102) );
  NAND2_X1 U7663 ( .A1(n6096), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n6115) );
  INV_X1 U7664 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n6097) );
  NAND2_X1 U7665 ( .A1(n6098), .A2(n6097), .ZN(n6099) );
  NAND2_X1 U7666 ( .A1(n6115), .A2(n6099), .ZN(n9142) );
  OR2_X1 U7667 ( .A1(n5827), .A2(n9142), .ZN(n6101) );
  INV_X1 U7668 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n9143) );
  OR2_X1 U7669 ( .A1(n8088), .A2(n9143), .ZN(n6100) );
  NAND4_X1 U7670 ( .A1(n6103), .A2(n6102), .A3(n6101), .A4(n6100), .ZN(n9123)
         );
  NAND2_X1 U7671 ( .A1(n9123), .A2(n5903), .ZN(n6104) );
  NAND2_X1 U7672 ( .A1(n6105), .A2(n6104), .ZN(n6106) );
  XNOR2_X1 U7673 ( .A(n6106), .B(n4297), .ZN(n6108) );
  AND2_X1 U7674 ( .A1(n9123), .A2(n6257), .ZN(n6107) );
  AOI21_X1 U7675 ( .B1(n9141), .B2(n6261), .A(n6107), .ZN(n6109) );
  NAND2_X1 U7676 ( .A1(n6108), .A2(n6109), .ZN(n6114) );
  INV_X1 U7677 ( .A(n6108), .ZN(n6111) );
  INV_X1 U7678 ( .A(n6109), .ZN(n6110) );
  NAND2_X1 U7679 ( .A1(n6111), .A2(n6110), .ZN(n6112) );
  NAND2_X1 U7680 ( .A1(n6113), .A2(n8913), .ZN(n8918) );
  NAND2_X1 U7681 ( .A1(n8918), .A2(n6114), .ZN(n8863) );
  NAND2_X1 U7682 ( .A1(n9296), .A2(n6262), .ZN(n6123) );
  NAND2_X1 U7683 ( .A1(n5862), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n6121) );
  INV_X1 U7684 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n8866) );
  NAND2_X1 U7685 ( .A1(n6115), .A2(n8866), .ZN(n6116) );
  NAND2_X1 U7686 ( .A1(n6132), .A2(n6116), .ZN(n9126) );
  OR2_X1 U7687 ( .A1(n9126), .A2(n5827), .ZN(n6120) );
  INV_X1 U7688 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n6117) );
  OR2_X1 U7689 ( .A1(n8082), .A2(n6117), .ZN(n6119) );
  INV_X1 U7690 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n9119) );
  OR2_X1 U7691 ( .A1(n8088), .A2(n9119), .ZN(n6118) );
  NAND4_X1 U7692 ( .A1(n6121), .A2(n6120), .A3(n6119), .A4(n6118), .ZN(n9104)
         );
  NAND2_X1 U7693 ( .A1(n9104), .A2(n6261), .ZN(n6122) );
  NAND2_X1 U7694 ( .A1(n6123), .A2(n6122), .ZN(n6124) );
  XNOR2_X1 U7695 ( .A(n6124), .B(n4298), .ZN(n6126) );
  AND2_X1 U7696 ( .A1(n9104), .A2(n6257), .ZN(n6125) );
  AOI21_X1 U7697 ( .B1(n9296), .B2(n6261), .A(n6125), .ZN(n6127) );
  XNOR2_X1 U7698 ( .A(n6126), .B(n6127), .ZN(n8864) );
  INV_X1 U7699 ( .A(n6126), .ZN(n6128) );
  NAND2_X1 U7700 ( .A1(n6128), .A2(n6127), .ZN(n6129) );
  NAND2_X1 U7701 ( .A1(n8862), .A2(n6129), .ZN(n6151) );
  INV_X1 U7702 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n6131) );
  NAND2_X1 U7703 ( .A1(n6132), .A2(n6131), .ZN(n6133) );
  NAND2_X1 U7704 ( .A1(n6158), .A2(n6133), .ZN(n9108) );
  OR2_X1 U7705 ( .A1(n9108), .A2(n5827), .ZN(n6137) );
  NAND2_X1 U7706 ( .A1(n6202), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n6136) );
  NAND2_X1 U7707 ( .A1(n5803), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n6135) );
  NAND2_X1 U7708 ( .A1(n5862), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n6134) );
  NAND4_X1 U7709 ( .A1(n6137), .A2(n6136), .A3(n6135), .A4(n6134), .ZN(n9295)
         );
  AND2_X1 U7710 ( .A1(n9295), .A2(n6257), .ZN(n6138) );
  AOI21_X1 U7711 ( .B1(n9286), .B2(n6261), .A(n6138), .ZN(n6152) );
  NAND2_X1 U7712 ( .A1(n9286), .A2(n6139), .ZN(n6141) );
  NAND2_X1 U7713 ( .A1(n9295), .A2(n6261), .ZN(n6140) );
  NAND2_X1 U7714 ( .A1(n6141), .A2(n6140), .ZN(n6142) );
  XNOR2_X1 U7715 ( .A(n6142), .B(n4298), .ZN(n8926) );
  NAND2_X1 U7716 ( .A1(n9096), .A2(n6262), .ZN(n6149) );
  INV_X1 U7717 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n10066) );
  NAND2_X1 U7718 ( .A1(n6202), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n6144) );
  NAND2_X1 U7719 ( .A1(n5803), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n6143) );
  OAI211_X1 U7720 ( .C1(n10066), .C2(n8084), .A(n6144), .B(n6143), .ZN(n6145)
         );
  INV_X1 U7721 ( .A(n6145), .ZN(n6147) );
  XNOR2_X1 U7722 ( .A(n6158), .B(P1_REG3_REG_23__SCAN_IN), .ZN(n9097) );
  NAND2_X1 U7723 ( .A1(n9097), .A2(n5845), .ZN(n6146) );
  NAND2_X1 U7724 ( .A1(n6147), .A2(n6146), .ZN(n9075) );
  NAND2_X1 U7725 ( .A1(n9075), .A2(n6261), .ZN(n6148) );
  NAND2_X1 U7726 ( .A1(n6149), .A2(n6148), .ZN(n6150) );
  XNOR2_X1 U7727 ( .A(n6150), .B(n4297), .ZN(n6154) );
  INV_X1 U7728 ( .A(n6257), .ZN(n6153) );
  OAI22_X1 U7729 ( .A1(n9358), .A2(n4320), .B1(n9289), .B2(n6153), .ZN(n8847)
         );
  NAND2_X1 U7730 ( .A1(n9278), .A2(n5806), .ZN(n6166) );
  INV_X1 U7731 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n6164) );
  INV_X1 U7732 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n6156) );
  INV_X1 U7733 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n6155) );
  OAI21_X1 U7734 ( .B1(n6158), .B2(n6156), .A(n6155), .ZN(n6159) );
  NAND2_X1 U7735 ( .A1(P1_REG3_REG_24__SCAN_IN), .A2(P1_REG3_REG_23__SCAN_IN), 
        .ZN(n6157) );
  NAND2_X1 U7736 ( .A1(n6159), .A2(n6176), .ZN(n8903) );
  OR2_X1 U7737 ( .A1(n8903), .A2(n5827), .ZN(n6163) );
  NAND2_X1 U7738 ( .A1(n6202), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n6161) );
  NAND2_X1 U7739 ( .A1(n5803), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n6160) );
  AND2_X1 U7740 ( .A1(n6161), .A2(n6160), .ZN(n6162) );
  OAI211_X1 U7741 ( .C1(n8084), .C2(n6164), .A(n6163), .B(n6162), .ZN(n9092)
         );
  NAND2_X1 U7742 ( .A1(n9092), .A2(n6261), .ZN(n6165) );
  NAND2_X1 U7743 ( .A1(n6166), .A2(n6165), .ZN(n6167) );
  XNOR2_X1 U7744 ( .A(n6167), .B(n4298), .ZN(n6171) );
  NAND2_X1 U7745 ( .A1(n9278), .A2(n5903), .ZN(n6169) );
  NAND2_X1 U7746 ( .A1(n9092), .A2(n6257), .ZN(n6168) );
  NAND2_X1 U7747 ( .A1(n6169), .A2(n6168), .ZN(n6170) );
  NOR2_X1 U7748 ( .A1(n6171), .A2(n6170), .ZN(n6172) );
  AOI21_X1 U7749 ( .B1(n6171), .B2(n6170), .A(n6172), .ZN(n8900) );
  NAND2_X1 U7750 ( .A1(n8899), .A2(n8900), .ZN(n8898) );
  INV_X1 U7751 ( .A(n6172), .ZN(n6173) );
  NAND2_X1 U7752 ( .A1(n8898), .A2(n6173), .ZN(n8872) );
  NAND2_X1 U7753 ( .A1(n9065), .A2(n6262), .ZN(n6181) );
  INV_X1 U7754 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n10158) );
  INV_X1 U7755 ( .A(n6176), .ZN(n6174) );
  NAND2_X1 U7756 ( .A1(n6174), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n6185) );
  INV_X1 U7757 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n6175) );
  NAND2_X1 U7758 ( .A1(n6176), .A2(n6175), .ZN(n6177) );
  NAND2_X1 U7759 ( .A1(n6185), .A2(n6177), .ZN(n8875) );
  OR2_X1 U7760 ( .A1(n8875), .A2(n5827), .ZN(n6179) );
  AOI22_X1 U7761 ( .A1(n5803), .A2(P1_REG2_REG_25__SCAN_IN), .B1(n6202), .B2(
        P1_REG1_REG_25__SCAN_IN), .ZN(n6178) );
  OAI211_X1 U7762 ( .C1(n8084), .C2(n10158), .A(n6179), .B(n6178), .ZN(n9076)
         );
  NAND2_X1 U7763 ( .A1(n9076), .A2(n6261), .ZN(n6180) );
  NAND2_X1 U7764 ( .A1(n6181), .A2(n6180), .ZN(n6182) );
  XNOR2_X1 U7765 ( .A(n6182), .B(n4298), .ZN(n6196) );
  AOI22_X1 U7766 ( .A1(n9065), .A2(n6261), .B1(n6257), .B2(n9076), .ZN(n6197)
         );
  XNOR2_X1 U7767 ( .A(n6196), .B(n6197), .ZN(n8873) );
  NAND2_X1 U7768 ( .A1(n8872), .A2(n8873), .ZN(n6245) );
  NAND2_X1 U7769 ( .A1(n9265), .A2(n5806), .ZN(n6193) );
  INV_X1 U7770 ( .A(n6185), .ZN(n6183) );
  NAND2_X1 U7771 ( .A1(n6183), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n6200) );
  INV_X1 U7772 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n6184) );
  NAND2_X1 U7773 ( .A1(n6185), .A2(n6184), .ZN(n6186) );
  NAND2_X1 U7774 ( .A1(n6200), .A2(n6186), .ZN(n6249) );
  OR2_X1 U7775 ( .A1(n6249), .A2(n5827), .ZN(n6191) );
  INV_X1 U7776 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n10163) );
  NAND2_X1 U7777 ( .A1(n5803), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n6188) );
  INV_X1 U7778 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n10123) );
  OR2_X1 U7779 ( .A1(n8084), .A2(n10123), .ZN(n6187) );
  OAI211_X1 U7780 ( .C1(n8082), .C2(n10163), .A(n6188), .B(n6187), .ZN(n6189)
         );
  INV_X1 U7781 ( .A(n6189), .ZN(n6190) );
  NAND2_X1 U7782 ( .A1(n6191), .A2(n6190), .ZN(n9028) );
  NAND2_X1 U7783 ( .A1(n9028), .A2(n6261), .ZN(n6192) );
  NAND2_X1 U7784 ( .A1(n6193), .A2(n6192), .ZN(n6194) );
  XNOR2_X1 U7785 ( .A(n6194), .B(n4298), .ZN(n6216) );
  AND2_X1 U7786 ( .A1(n9028), .A2(n6257), .ZN(n6195) );
  AOI21_X1 U7787 ( .B1(n9265), .B2(n6261), .A(n6195), .ZN(n6214) );
  XNOR2_X1 U7788 ( .A(n6216), .B(n6214), .ZN(n6246) );
  INV_X1 U7789 ( .A(n6196), .ZN(n6198) );
  NAND2_X1 U7790 ( .A1(n6198), .A2(n6197), .ZN(n6247) );
  NAND2_X1 U7791 ( .A1(n9021), .A2(n6262), .ZN(n6209) );
  INV_X1 U7792 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n6199) );
  NAND2_X1 U7793 ( .A1(n6200), .A2(n6199), .ZN(n6201) );
  NAND2_X1 U7794 ( .A1(n8290), .A2(n6201), .ZN(n9023) );
  OR2_X1 U7795 ( .A1(n9023), .A2(n5827), .ZN(n6207) );
  INV_X1 U7796 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n9022) );
  NAND2_X1 U7797 ( .A1(n5862), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n6204) );
  NAND2_X1 U7798 ( .A1(n6202), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n6203) );
  OAI211_X1 U7799 ( .C1(n9022), .C2(n8088), .A(n6204), .B(n6203), .ZN(n6205)
         );
  INV_X1 U7800 ( .A(n6205), .ZN(n6206) );
  NAND2_X1 U7801 ( .A1(n6207), .A2(n6206), .ZN(n9047) );
  NAND2_X1 U7802 ( .A1(n9047), .A2(n6261), .ZN(n6208) );
  NAND2_X1 U7803 ( .A1(n6209), .A2(n6208), .ZN(n6210) );
  XNOR2_X1 U7804 ( .A(n6210), .B(n4297), .ZN(n6213) );
  AND2_X1 U7805 ( .A1(n9047), .A2(n6257), .ZN(n6211) );
  AOI21_X1 U7806 ( .B1(n9021), .B2(n6261), .A(n6211), .ZN(n6212) );
  NAND2_X1 U7807 ( .A1(n6213), .A2(n6212), .ZN(n6278) );
  OAI21_X1 U7808 ( .B1(n6213), .B2(n6212), .A(n6278), .ZN(n6218) );
  INV_X1 U7809 ( .A(n6214), .ZN(n6215) );
  INV_X1 U7810 ( .A(n6217), .ZN(n6220) );
  INV_X1 U7811 ( .A(n6218), .ZN(n6219) );
  NAND2_X1 U7812 ( .A1(n9654), .A2(n7054), .ZN(n9652) );
  NAND3_X1 U7813 ( .A1(n9678), .A2(n6232), .A3(n8098), .ZN(n6221) );
  NOR2_X2 U7814 ( .A1(n9652), .A2(n6221), .ZN(n8901) );
  INV_X1 U7815 ( .A(n6232), .ZN(n6223) );
  OR2_X1 U7816 ( .A1(n7042), .A2(n6222), .ZN(n9634) );
  OR2_X1 U7817 ( .A1(n6223), .A2(n9634), .ZN(n6224) );
  NOR2_X1 U7818 ( .A1(n9652), .A2(n6224), .ZN(n6239) );
  AND2_X1 U7819 ( .A1(n6239), .A2(n5718), .ZN(n8922) );
  XNOR2_X1 U7820 ( .A(n8290), .B(P1_REG3_REG_28__SCAN_IN), .ZN(n9014) );
  NAND2_X1 U7821 ( .A1(n9014), .A2(n5845), .ZN(n6231) );
  INV_X1 U7822 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n6228) );
  NAND2_X1 U7823 ( .A1(n5803), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n6227) );
  INV_X1 U7824 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n6225) );
  OR2_X1 U7825 ( .A1(n8084), .A2(n6225), .ZN(n6226) );
  OAI211_X1 U7826 ( .C1(n8082), .C2(n6228), .A(n6227), .B(n6226), .ZN(n6229)
         );
  INV_X1 U7827 ( .A(n6229), .ZN(n6230) );
  NAND2_X1 U7828 ( .A1(n6231), .A2(n6230), .ZN(n9029) );
  AND2_X1 U7829 ( .A1(n6232), .A2(n7054), .ZN(n6233) );
  OR2_X1 U7830 ( .A1(n6234), .A2(n6233), .ZN(n6243) );
  NAND2_X1 U7831 ( .A1(n6236), .A2(n6235), .ZN(n6237) );
  NAND2_X1 U7832 ( .A1(n6237), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6238) );
  NAND2_X1 U7833 ( .A1(n6243), .A2(n6238), .ZN(n8907) );
  AOI22_X1 U7834 ( .A1(n9028), .A2(n8938), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3084), .ZN(n6240) );
  OAI21_X1 U7835 ( .B1(n8940), .B2(n9023), .A(n6240), .ZN(n6241) );
  AOI21_X1 U7836 ( .B1(n8922), .B2(n9029), .A(n6241), .ZN(n6244) );
  INV_X1 U7837 ( .A(n7056), .ZN(n6242) );
  NAND2_X1 U7838 ( .A1(n6243), .A2(n6242), .ZN(n6761) );
  INV_X1 U7839 ( .A(n6761), .ZN(n7241) );
  NAND2_X1 U7840 ( .A1(n7241), .A2(n9695), .ZN(n8910) );
  AOI21_X1 U7841 ( .B1(n8871), .B2(n6247), .A(n6246), .ZN(n6256) );
  NAND2_X1 U7842 ( .A1(n6248), .A2(n8901), .ZN(n6255) );
  INV_X1 U7843 ( .A(n9265), .ZN(n9042) );
  INV_X1 U7844 ( .A(n6249), .ZN(n9040) );
  INV_X1 U7845 ( .A(n9047), .ZN(n8078) );
  INV_X1 U7846 ( .A(n8922), .ZN(n8936) );
  AOI22_X1 U7847 ( .A1(n9076), .A2(n8938), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3084), .ZN(n6250) );
  OAI21_X1 U7848 ( .B1(n8078), .B2(n8936), .A(n6250), .ZN(n6251) );
  AOI21_X1 U7849 ( .B1(n9040), .B2(n8907), .A(n6251), .ZN(n6252) );
  OAI21_X1 U7850 ( .B1(n6256), .B2(n6255), .A(n6254), .ZN(P1_U3238) );
  NAND2_X1 U7851 ( .A1(n9015), .A2(n5903), .ZN(n6259) );
  NAND2_X1 U7852 ( .A1(n9029), .A2(n6257), .ZN(n6258) );
  NAND2_X1 U7853 ( .A1(n6259), .A2(n6258), .ZN(n6260) );
  XNOR2_X1 U7854 ( .A(n6260), .B(n4298), .ZN(n6264) );
  AOI22_X1 U7855 ( .A1(n9015), .A2(n6262), .B1(n6261), .B2(n9029), .ZN(n6263)
         );
  XNOR2_X1 U7856 ( .A(n6264), .B(n6263), .ZN(n6275) );
  NAND3_X1 U7857 ( .A1(n6281), .A2(n8901), .A3(n6275), .ZN(n6284) );
  INV_X1 U7858 ( .A(n8938), .ZN(n8905) );
  NAND2_X1 U7859 ( .A1(n5845), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n6265) );
  OR2_X1 U7860 ( .A1(n8290), .A2(n6265), .ZN(n6272) );
  INV_X1 U7861 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n6269) );
  INV_X1 U7862 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n8294) );
  OR2_X1 U7863 ( .A1(n8088), .A2(n8294), .ZN(n6268) );
  INV_X1 U7864 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n6266) );
  OR2_X1 U7865 ( .A1(n8084), .A2(n6266), .ZN(n6267) );
  OAI211_X1 U7866 ( .C1(n8082), .C2(n6269), .A(n6268), .B(n6267), .ZN(n6270)
         );
  INV_X1 U7867 ( .A(n6270), .ZN(n6271) );
  NAND2_X1 U7868 ( .A1(n6272), .A2(n6271), .ZN(n9010) );
  AOI22_X1 U7869 ( .A1(n9010), .A2(n8922), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n6274) );
  NAND2_X1 U7870 ( .A1(n9014), .A2(n8907), .ZN(n6273) );
  OAI211_X1 U7871 ( .C1(n8078), .C2(n8905), .A(n6274), .B(n6273), .ZN(n6277)
         );
  INV_X1 U7872 ( .A(n6275), .ZN(n6279) );
  NOR3_X1 U7873 ( .A1(n6279), .A2(n8944), .A3(n6278), .ZN(n6276) );
  AOI211_X1 U7874 ( .C1(n8942), .C2(n9015), .A(n6277), .B(n6276), .ZN(n6283)
         );
  NAND3_X1 U7875 ( .A1(n6279), .A2(n8901), .A3(n6278), .ZN(n6280) );
  NAND3_X1 U7876 ( .A1(n6284), .A2(n6283), .A3(n6282), .ZN(P1_U3218) );
  INV_X1 U7877 ( .A(n7098), .ZN(n6285) );
  OR2_X1 U7878 ( .A1(n8098), .A2(n6285), .ZN(n6287) );
  OR2_X1 U7879 ( .A1(n6286), .A2(n6285), .ZN(n6319) );
  NAND2_X1 U7880 ( .A1(n6287), .A2(n6319), .ZN(n6315) );
  OAI21_X1 U7881 ( .B1(n6315), .B2(n6288), .A(P1_STATE_REG_SCAN_IN), .ZN(
        P1_U3083) );
  OR2_X2 U7882 ( .A1(n6319), .A2(P1_U3084), .ZN(n8956) );
  INV_X1 U7883 ( .A(n8956), .ZN(P1_U4006) );
  NOR2_X1 U7884 ( .A1(n6665), .A2(P2_U3152), .ZN(n6377) );
  AND2_X1 U7885 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7464) );
  NOR2_X1 U7886 ( .A1(n9523), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6289) );
  AOI21_X1 U7887 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n9523), .A(n6289), .ZN(
        n9525) );
  NOR2_X1 U7888 ( .A1(P1_REG2_REG_7__SCAN_IN), .A2(n6564), .ZN(n6290) );
  AOI21_X1 U7889 ( .B1(n6564), .B2(P1_REG2_REG_7__SCAN_IN), .A(n6290), .ZN(
        n6562) );
  NOR2_X1 U7890 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(n9511), .ZN(n6291) );
  AOI21_X1 U7891 ( .B1(n9511), .B2(P1_REG2_REG_5__SCAN_IN), .A(n6291), .ZN(
        n9513) );
  INV_X1 U7892 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6292) );
  MUX2_X1 U7893 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n6292), .S(n6630), .Z(n6620)
         );
  AND2_X1 U7894 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n6619) );
  NAND2_X1 U7895 ( .A1(n6620), .A2(n6619), .ZN(n6618) );
  NAND2_X1 U7896 ( .A1(n6630), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6293) );
  NAND2_X1 U7897 ( .A1(n6618), .A2(n6293), .ZN(n9477) );
  OR2_X1 U7898 ( .A1(n9492), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6295) );
  NAND2_X1 U7899 ( .A1(n9492), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6294) );
  AND2_X1 U7900 ( .A1(n6295), .A2(n6294), .ZN(n9478) );
  NAND2_X1 U7901 ( .A1(n9425), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6296) );
  OAI21_X1 U7902 ( .B1(n9425), .B2(P1_REG2_REG_3__SCAN_IN), .A(n6296), .ZN(
        n9428) );
  NOR2_X1 U7903 ( .A1(n9501), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6297) );
  AOI21_X1 U7904 ( .B1(P1_REG2_REG_4__SCAN_IN), .B2(n9501), .A(n6297), .ZN(
        n9499) );
  NAND2_X1 U7905 ( .A1(n4334), .A2(n9499), .ZN(n9498) );
  OAI21_X1 U7906 ( .B1(n9501), .B2(P1_REG2_REG_4__SCAN_IN), .A(n9498), .ZN(
        n9514) );
  NAND2_X1 U7907 ( .A1(n9513), .A2(n9514), .ZN(n9512) );
  OAI21_X1 U7908 ( .B1(P1_REG2_REG_5__SCAN_IN), .B2(n9511), .A(n9512), .ZN(
        n6594) );
  MUX2_X1 U7909 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n7310), .S(n6597), .Z(n6298)
         );
  INV_X1 U7910 ( .A(n6298), .ZN(n6593) );
  NOR2_X1 U7911 ( .A1(n6594), .A2(n6593), .ZN(n6592) );
  AOI21_X1 U7912 ( .B1(P1_REG2_REG_6__SCAN_IN), .B2(n6597), .A(n6592), .ZN(
        n6561) );
  NAND2_X1 U7913 ( .A1(n6562), .A2(n6561), .ZN(n6560) );
  OAI21_X1 U7914 ( .B1(P1_REG2_REG_7__SCAN_IN), .B2(n6564), .A(n6560), .ZN(
        n9526) );
  NAND2_X1 U7915 ( .A1(n9525), .A2(n9526), .ZN(n9524) );
  OAI21_X1 U7916 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n9523), .A(n9524), .ZN(
        n6301) );
  NAND2_X1 U7917 ( .A1(n6610), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6299) );
  OAI21_X1 U7918 ( .B1(n6610), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6299), .ZN(
        n6300) );
  NOR2_X1 U7919 ( .A1(n6301), .A2(n6300), .ZN(n6609) );
  OR2_X1 U7920 ( .A1(n6315), .A2(P1_U3084), .ZN(n9471) );
  NOR2_X1 U7921 ( .A1(n9471), .A2(n9479), .ZN(n8980) );
  INV_X1 U7922 ( .A(n8980), .ZN(n6318) );
  OR2_X1 U7923 ( .A1(n6318), .A2(n5718), .ZN(n9580) );
  AOI211_X1 U7924 ( .C1(n6301), .C2(n6300), .A(n6609), .B(n9580), .ZN(n6323)
         );
  NAND2_X1 U7925 ( .A1(n9523), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6312) );
  MUX2_X1 U7926 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n6302), .S(n9523), .Z(n9529)
         );
  NOR2_X1 U7927 ( .A1(P1_REG1_REG_7__SCAN_IN), .A2(n6564), .ZN(n6311) );
  INV_X1 U7928 ( .A(n6597), .ZN(n6331) );
  NAND2_X1 U7929 ( .A1(P1_REG1_REG_5__SCAN_IN), .A2(n9511), .ZN(n6310) );
  MUX2_X1 U7930 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n6303), .S(n9511), .Z(n9517)
         );
  NOR2_X1 U7931 ( .A1(n9501), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6309) );
  INV_X1 U7932 ( .A(n9501), .ZN(n6328) );
  AOI22_X1 U7933 ( .A1(n9501), .A2(n5824), .B1(P1_REG1_REG_4__SCAN_IN), .B2(
        n6328), .ZN(n9504) );
  NAND2_X1 U7934 ( .A1(n9425), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6308) );
  MUX2_X1 U7935 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n6304), .S(n9425), .Z(n9431)
         );
  MUX2_X1 U7936 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n6305), .S(n6630), .Z(n6624)
         );
  AND2_X1 U7937 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n6625) );
  NAND2_X1 U7938 ( .A1(n6624), .A2(n6625), .ZN(n6623) );
  NAND2_X1 U7939 ( .A1(n6630), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6306) );
  NAND2_X1 U7940 ( .A1(n6623), .A2(n6306), .ZN(n9488) );
  XNOR2_X1 U7941 ( .A(n9492), .B(n9724), .ZN(n9487) );
  AOI22_X1 U7942 ( .A1(n9488), .A2(n9487), .B1(P1_REG1_REG_2__SCAN_IN), .B2(
        n9492), .ZN(n6307) );
  INV_X1 U7943 ( .A(n6307), .ZN(n9432) );
  NAND2_X1 U7944 ( .A1(n9431), .A2(n9432), .ZN(n9430) );
  NAND2_X1 U7945 ( .A1(n6308), .A2(n9430), .ZN(n9503) );
  NOR2_X1 U7946 ( .A1(n9504), .A2(n9503), .ZN(n9502) );
  NOR2_X1 U7947 ( .A1(n6309), .A2(n9502), .ZN(n9518) );
  NAND2_X1 U7948 ( .A1(n9517), .A2(n9518), .ZN(n9516) );
  NAND2_X1 U7949 ( .A1(n6310), .A2(n9516), .ZN(n6589) );
  AOI22_X1 U7950 ( .A1(n6597), .A2(n5863), .B1(P1_REG1_REG_6__SCAN_IN), .B2(
        n6331), .ZN(n6588) );
  NOR2_X1 U7951 ( .A1(n6589), .A2(n6588), .ZN(n6587) );
  AOI21_X1 U7952 ( .B1(n6331), .B2(n5863), .A(n6587), .ZN(n6559) );
  INV_X1 U7953 ( .A(n6564), .ZN(n6346) );
  AOI22_X1 U7954 ( .A1(P1_REG1_REG_7__SCAN_IN), .A2(n6346), .B1(n6564), .B2(
        n5877), .ZN(n6558) );
  NOR2_X1 U7955 ( .A1(n6559), .A2(n6558), .ZN(n6557) );
  NOR2_X1 U7956 ( .A1(n6311), .A2(n6557), .ZN(n9530) );
  NAND2_X1 U7957 ( .A1(n9529), .A2(n9530), .ZN(n9528) );
  NAND2_X1 U7958 ( .A1(n6312), .A2(n9528), .ZN(n6314) );
  AOI22_X1 U7959 ( .A1(n6610), .A2(n5912), .B1(P1_REG1_REG_9__SCAN_IN), .B2(
        n6359), .ZN(n6313) );
  NOR2_X1 U7960 ( .A1(n6314), .A2(n6313), .ZN(n6603) );
  AOI21_X1 U7961 ( .B1(n6314), .B2(n6313), .A(n6603), .ZN(n6317) );
  NOR2_X1 U7962 ( .A1(n5718), .A2(P1_U3084), .ZN(n7546) );
  NAND2_X1 U7963 ( .A1(n7546), .A2(n9479), .ZN(n6316) );
  NOR2_X1 U7964 ( .A1(n6317), .A2(n9605), .ZN(n6322) );
  OR2_X1 U7965 ( .A1(n6318), .A2(n4568), .ZN(n9599) );
  INV_X1 U7966 ( .A(n6319), .ZN(n6320) );
  INV_X1 U7967 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10192) );
  OAI22_X1 U7968 ( .A1(n9599), .A2(n6359), .B1(n9609), .B2(n10192), .ZN(n6321)
         );
  OR4_X1 U7969 ( .A1(n7464), .A2(n6323), .A3(n6322), .A4(n6321), .ZN(P1_U3250)
         );
  AND2_X1 U7970 ( .A1(n6327), .A2(P2_U3152), .ZN(n8841) );
  INV_X1 U7971 ( .A(n8841), .ZN(n7714) );
  NOR2_X1 U7972 ( .A1(n6326), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8253) );
  INV_X1 U7973 ( .A(n6427), .ZN(n6436) );
  OAI222_X1 U7974 ( .A1(n7714), .A2(n6324), .B1(n8844), .B2(n6329), .C1(
        P2_U3152), .C2(n6436), .ZN(P2_U3354) );
  INV_X1 U7975 ( .A(n6551), .ZN(n6389) );
  OAI222_X1 U7976 ( .A1(n7714), .A2(n6325), .B1(n8844), .B2(n6343), .C1(
        P2_U3152), .C2(n6389), .ZN(P2_U3353) );
  NOR2_X1 U7977 ( .A1(n6326), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9389) );
  INV_X1 U7978 ( .A(n9389), .ZN(n7688) );
  NAND2_X1 U7979 ( .A1(n6327), .A2(P1_U3084), .ZN(n7399) );
  OAI222_X1 U7980 ( .A1(n7688), .A2(n6330), .B1(n7399), .B2(n6329), .C1(
        P1_U3084), .C2(n6328), .ZN(P1_U3349) );
  OAI222_X1 U7981 ( .A1(n7688), .A2(n6332), .B1(n7399), .B2(n6333), .C1(
        P1_U3084), .C2(n6331), .ZN(P1_U3347) );
  INV_X1 U7982 ( .A(n6413), .ZN(n6466) );
  OAI222_X1 U7983 ( .A1(n7714), .A2(n6334), .B1(n8844), .B2(n6333), .C1(
        P2_U3152), .C2(n6466), .ZN(P2_U3352) );
  AOI22_X1 U7984 ( .A1(n8841), .A2(P1_DATAO_REG_3__SCAN_IN), .B1(n9744), .B2(
        P2_STATE_REG_SCAN_IN), .ZN(n6335) );
  OAI21_X1 U7985 ( .B1(n6340), .B2(n8844), .A(n6335), .ZN(P2_U3355) );
  AOI22_X1 U7986 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(n8841), .B1(n9437), .B2(
        P2_STATE_REG_SCAN_IN), .ZN(n6336) );
  OAI21_X1 U7987 ( .B1(n6338), .B2(n8844), .A(n6336), .ZN(P2_U3356) );
  CLKBUF_X1 U7988 ( .A(n7399), .Z(n9391) );
  AOI22_X1 U7989 ( .A1(n9389), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(n9492), .B2(
        P1_STATE_REG_SCAN_IN), .ZN(n6337) );
  OAI21_X1 U7990 ( .B1(n6338), .B2(n9391), .A(n6337), .ZN(P1_U3351) );
  AOI22_X1 U7991 ( .A1(P2_DATAO_REG_3__SCAN_IN), .A2(n9389), .B1(n9425), .B2(
        P1_STATE_REG_SCAN_IN), .ZN(n6339) );
  OAI21_X1 U7992 ( .B1(n6340), .B2(n9391), .A(n6339), .ZN(P1_U3350) );
  AOI22_X1 U7993 ( .A1(n9389), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(n6630), .B2(
        P1_STATE_REG_SCAN_IN), .ZN(n6341) );
  OAI21_X1 U7994 ( .B1(n6344), .B2(n9391), .A(n6341), .ZN(P1_U3352) );
  AOI22_X1 U7995 ( .A1(n9511), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n9389), .ZN(n6342) );
  OAI21_X1 U7996 ( .B1(n6343), .B2(n9391), .A(n6342), .ZN(P1_U3348) );
  INV_X1 U7997 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6345) );
  OAI222_X1 U7998 ( .A1(n7714), .A2(n6345), .B1(n8844), .B2(n6344), .C1(
        P2_U3152), .C2(n5031), .ZN(P2_U3357) );
  OAI222_X1 U7999 ( .A1(n7688), .A2(n4438), .B1(n7399), .B2(n6348), .C1(
        P1_U3084), .C2(n6346), .ZN(P1_U3346) );
  INV_X1 U8000 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6349) );
  OAI222_X1 U8001 ( .A1(n7714), .A2(n6349), .B1(n8844), .B2(n6348), .C1(
        P2_U3152), .C2(n6347), .ZN(P2_U3351) );
  INV_X1 U8002 ( .A(n6350), .ZN(n6353) );
  INV_X1 U8003 ( .A(n6495), .ZN(n6468) );
  OAI222_X1 U8004 ( .A1(n7714), .A2(n6351), .B1(n8844), .B2(n6353), .C1(
        P2_U3152), .C2(n6468), .ZN(P2_U3350) );
  OAI222_X1 U8005 ( .A1(n7688), .A2(n6354), .B1(n7399), .B2(n6353), .C1(
        P1_U3084), .C2(n6352), .ZN(P1_U3345) );
  OAI21_X1 U8006 ( .B1(n9868), .B2(n6692), .A(n5050), .ZN(n6356) );
  OR2_X1 U8007 ( .A1(n9871), .A2(P2_U3152), .ZN(n8005) );
  NAND2_X1 U8008 ( .A1(n9868), .A2(n8005), .ZN(n6355) );
  NAND2_X1 U8009 ( .A1(n6356), .A2(n6355), .ZN(n8464) );
  NOR2_X1 U8010 ( .A1(n9781), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U8011 ( .A(n6357), .ZN(n6360) );
  INV_X1 U8012 ( .A(n6507), .ZN(n6469) );
  OAI222_X1 U8013 ( .A1(n7714), .A2(n6358), .B1(n8844), .B2(n6360), .C1(n6469), 
        .C2(P2_U3152), .ZN(P2_U3349) );
  OAI222_X1 U8014 ( .A1(n7688), .A2(n6361), .B1(n7399), .B2(n6360), .C1(n6359), 
        .C2(P1_U3084), .ZN(P1_U3344) );
  INV_X1 U8015 ( .A(n6362), .ZN(n6365) );
  OAI222_X1 U8016 ( .A1(n7688), .A2(n6363), .B1(n7399), .B2(n6365), .C1(n6605), 
        .C2(P1_U3084), .ZN(P1_U3343) );
  INV_X1 U8017 ( .A(n9770), .ZN(n6364) );
  OAI222_X1 U8018 ( .A1(n7714), .A2(n10004), .B1(n8844), .B2(n6365), .C1(n6364), .C2(P2_U3152), .ZN(P2_U3348) );
  NAND2_X1 U8019 ( .A1(n5078), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n6369) );
  NAND2_X1 U8020 ( .A1(n6366), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n6368) );
  NAND2_X1 U8021 ( .A1(n5068), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n6367) );
  AND3_X1 U8022 ( .A1(n6369), .A2(n6368), .A3(n6367), .ZN(n7988) );
  INV_X2 U8023 ( .A(P2_U3966), .ZN(n8444) );
  NAND2_X1 U8024 ( .A1(n8444), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n6370) );
  OAI21_X1 U8025 ( .B1(n7988), .B2(n8444), .A(n6370), .ZN(P2_U3583) );
  INV_X1 U8026 ( .A(n6371), .ZN(n6373) );
  OAI222_X1 U8027 ( .A1(n7688), .A2(n6372), .B1(n7399), .B2(n6373), .C1(n6803), 
        .C2(P1_U3084), .ZN(P1_U3342) );
  INV_X1 U8028 ( .A(n6524), .ZN(n6521) );
  OAI222_X1 U8029 ( .A1(n7714), .A2(n6374), .B1(n8844), .B2(n6373), .C1(n6521), 
        .C2(P2_U3152), .ZN(P2_U3347) );
  INV_X1 U8030 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6376) );
  NAND2_X1 U8031 ( .A1(n8097), .A2(P1_U4006), .ZN(n6375) );
  OAI21_X1 U8032 ( .B1(P1_U4006), .B2(n6376), .A(n6375), .ZN(P1_U3586) );
  INV_X1 U8033 ( .A(n6377), .ZN(n6378) );
  OAI211_X1 U8034 ( .C1(n6379), .C2(n9868), .A(n6378), .B(n8005), .ZN(n6380)
         );
  AND2_X1 U8035 ( .A1(n6380), .A2(n5050), .ZN(n6399) );
  INV_X1 U8036 ( .A(n6399), .ZN(n6381) );
  NAND2_X1 U8037 ( .A1(n6381), .A2(n8444), .ZN(n6393) );
  NAND2_X1 U8038 ( .A1(n6393), .A2(n5459), .ZN(n9734) );
  NAND2_X1 U8039 ( .A1(P2_REG2_REG_3__SCAN_IN), .A2(n9744), .ZN(n6387) );
  INV_X1 U8040 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6382) );
  MUX2_X1 U8041 ( .A(n6382), .B(P2_REG2_REG_3__SCAN_IN), .S(n9744), .Z(n6383)
         );
  INV_X1 U8042 ( .A(n6383), .ZN(n9749) );
  INV_X1 U8043 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6384) );
  MUX2_X1 U8044 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n6384), .S(n9437), .Z(n9442)
         );
  INV_X1 U8045 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n7107) );
  MUX2_X1 U8046 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n7107), .S(n6443), .Z(n6385)
         );
  NAND3_X1 U8047 ( .A1(n6385), .A2(P2_REG2_REG_0__SCAN_IN), .A3(
        P2_IR_REG_0__SCAN_IN), .ZN(n6445) );
  OAI21_X1 U8048 ( .B1(n7107), .B2(n5031), .A(n6445), .ZN(n9443) );
  NAND2_X1 U8049 ( .A1(n9442), .A2(n9443), .ZN(n9441) );
  NAND2_X1 U8050 ( .A1(P2_REG2_REG_2__SCAN_IN), .A2(n9437), .ZN(n6386) );
  NAND2_X1 U8051 ( .A1(n9441), .A2(n6386), .ZN(n9750) );
  NAND2_X1 U8052 ( .A1(n9749), .A2(n9750), .ZN(n9748) );
  NAND2_X1 U8053 ( .A1(n6387), .A2(n9748), .ZN(n6433) );
  MUX2_X1 U8054 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n6953), .S(n6427), .Z(n6432)
         );
  NAND2_X1 U8055 ( .A1(n6433), .A2(n6432), .ZN(n6546) );
  NAND2_X1 U8056 ( .A1(n6427), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6545) );
  INV_X1 U8057 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n6388) );
  MUX2_X1 U8058 ( .A(n6388), .B(P2_REG2_REG_5__SCAN_IN), .S(n6551), .Z(n6544)
         );
  AOI21_X1 U8059 ( .B1(n6546), .B2(n6545), .A(n6544), .ZN(n6548) );
  INV_X1 U8060 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6456) );
  MUX2_X1 U8061 ( .A(n6456), .B(P2_REG2_REG_6__SCAN_IN), .S(n6413), .Z(n6391)
         );
  NOR2_X1 U8062 ( .A1(n6389), .A2(n6388), .ZN(n6397) );
  INV_X1 U8063 ( .A(n6397), .ZN(n6390) );
  NAND2_X1 U8064 ( .A1(n6391), .A2(n6390), .ZN(n6398) );
  INV_X1 U8065 ( .A(n8002), .ZN(n6392) );
  NAND2_X1 U8066 ( .A1(n6393), .A2(n6392), .ZN(n9736) );
  INV_X1 U8067 ( .A(n9736), .ZN(n6395) );
  MUX2_X1 U8068 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n6456), .S(n6413), .Z(n6396)
         );
  OAI21_X1 U8069 ( .B1(n6548), .B2(n6397), .A(n6396), .ZN(n6455) );
  OAI211_X1 U8070 ( .C1(n6548), .C2(n6398), .A(n9783), .B(n6455), .ZN(n6421)
         );
  AND2_X1 U8071 ( .A1(n6399), .A2(n8002), .ZN(n9786) );
  NAND2_X1 U8072 ( .A1(P2_REG1_REG_3__SCAN_IN), .A2(n9744), .ZN(n6405) );
  INV_X1 U8073 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6400) );
  MUX2_X1 U8074 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n6400), .S(n9744), .Z(n9746)
         );
  INV_X1 U8075 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6704) );
  MUX2_X1 U8076 ( .A(n6704), .B(P2_REG1_REG_1__SCAN_IN), .S(n6443), .Z(n6439)
         );
  INV_X1 U8077 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n6401) );
  INV_X1 U8078 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n6437) );
  NOR3_X1 U8079 ( .A1(n6439), .A2(n6401), .A3(n6437), .ZN(n6438) );
  INV_X1 U8080 ( .A(n6438), .ZN(n6402) );
  OAI21_X1 U8081 ( .B1(n6704), .B2(n5031), .A(n6402), .ZN(n9440) );
  INV_X1 U8082 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6403) );
  MUX2_X1 U8083 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n6403), .S(n9437), .Z(n9439)
         );
  NAND2_X1 U8084 ( .A1(n9440), .A2(n9439), .ZN(n9438) );
  NAND2_X1 U8085 ( .A1(P2_REG1_REG_2__SCAN_IN), .A2(n9437), .ZN(n6404) );
  NAND2_X1 U8086 ( .A1(n9438), .A2(n6404), .ZN(n9747) );
  NAND2_X1 U8087 ( .A1(n9746), .A2(n9747), .ZN(n9745) );
  NAND2_X1 U8088 ( .A1(n6405), .A2(n9745), .ZN(n6426) );
  INV_X1 U8089 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6406) );
  MUX2_X1 U8090 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n6406), .S(n6427), .Z(n6407)
         );
  AND2_X1 U8091 ( .A1(n6427), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6536) );
  INV_X1 U8092 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6408) );
  MUX2_X1 U8093 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n6408), .S(n6551), .Z(n6409)
         );
  OAI21_X1 U8094 ( .B1(n6535), .B2(n6536), .A(n6409), .ZN(n6541) );
  NAND2_X1 U8095 ( .A1(n6551), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6415) );
  NAND2_X1 U8096 ( .A1(n6541), .A2(n6415), .ZN(n6412) );
  INV_X1 U8097 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6410) );
  MUX2_X1 U8098 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n6410), .S(n6413), .Z(n6411)
         );
  NAND2_X1 U8099 ( .A1(n6412), .A2(n6411), .ZN(n6465) );
  MUX2_X1 U8100 ( .A(n6410), .B(P2_REG1_REG_6__SCAN_IN), .S(n6413), .Z(n6414)
         );
  NAND3_X1 U8101 ( .A1(n6541), .A2(n6415), .A3(n6414), .ZN(n6416) );
  AND2_X1 U8102 ( .A1(n6465), .A2(n6416), .ZN(n6419) );
  INV_X1 U8103 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n6417) );
  NAND2_X1 U8104 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3152), .ZN(n6840) );
  OAI21_X1 U8105 ( .B1(n8464), .B2(n6417), .A(n6840), .ZN(n6418) );
  AOI21_X1 U8106 ( .B1(n9786), .B2(n6419), .A(n6418), .ZN(n6420) );
  OAI211_X1 U8107 ( .C1(n9734), .C2(n6466), .A(n6421), .B(n6420), .ZN(P2_U3251) );
  INV_X1 U8108 ( .A(n6422), .ZN(n6424) );
  OAI222_X1 U8109 ( .A1(n7688), .A2(n6423), .B1(n7399), .B2(n6424), .C1(
        P1_U3084), .C2(n6931), .ZN(P1_U3341) );
  INV_X1 U8110 ( .A(n6574), .ZN(n6571) );
  OAI222_X1 U8111 ( .A1(n7714), .A2(n6425), .B1(n8844), .B2(n6424), .C1(
        P2_U3152), .C2(n6571), .ZN(P2_U3346) );
  NAND2_X1 U8112 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3152), .ZN(n6744) );
  INV_X1 U8113 ( .A(n6744), .ZN(n6431) );
  INV_X1 U8114 ( .A(n6426), .ZN(n6429) );
  MUX2_X1 U8115 ( .A(n6406), .B(P2_REG1_REG_4__SCAN_IN), .S(n6427), .Z(n6428)
         );
  INV_X1 U8116 ( .A(n9786), .ZN(n9735) );
  AOI211_X1 U8117 ( .C1(n6429), .C2(n6428), .A(n6535), .B(n9735), .ZN(n6430)
         );
  AOI211_X1 U8118 ( .C1(n9781), .C2(P2_ADDR_REG_4__SCAN_IN), .A(n6431), .B(
        n6430), .ZN(n6435) );
  OAI211_X1 U8119 ( .C1(n6433), .C2(n6432), .A(n9783), .B(n6546), .ZN(n6434)
         );
  OAI211_X1 U8120 ( .C1(n9734), .C2(n6436), .A(n6435), .B(n6434), .ZN(P2_U3249) );
  INV_X1 U8121 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n9964) );
  NOR2_X1 U8122 ( .A1(n8464), .A2(n9964), .ZN(n6442) );
  OR2_X1 U8123 ( .A1(n6437), .A2(n6401), .ZN(n6440) );
  AOI211_X1 U8124 ( .C1(n6440), .C2(n6439), .A(n6438), .B(n9735), .ZN(n6441)
         );
  AOI211_X1 U8125 ( .C1(P2_REG3_REG_1__SCAN_IN), .C2(P2_U3152), .A(n6442), .B(
        n6441), .ZN(n6449) );
  AND2_X1 U8126 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(
        n6447) );
  MUX2_X1 U8127 ( .A(n7107), .B(P2_REG2_REG_1__SCAN_IN), .S(n6443), .Z(n6444)
         );
  INV_X1 U8128 ( .A(n6444), .ZN(n6446) );
  OAI211_X1 U8129 ( .C1(n6447), .C2(n6446), .A(n9783), .B(n6445), .ZN(n6448)
         );
  OAI211_X1 U8130 ( .C1(n9734), .C2(n5031), .A(n6449), .B(n6448), .ZN(P2_U3246) );
  AOI22_X1 U8131 ( .A1(P2_REG2_REG_11__SCAN_IN), .A2(n6521), .B1(n6524), .B2(
        n5183), .ZN(n6462) );
  NAND2_X1 U8132 ( .A1(P2_REG2_REG_10__SCAN_IN), .A2(n9770), .ZN(n6460) );
  INV_X1 U8133 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n6450) );
  MUX2_X1 U8134 ( .A(n6450), .B(P2_REG2_REG_10__SCAN_IN), .S(n9770), .Z(n6451)
         );
  INV_X1 U8135 ( .A(n6451), .ZN(n9775) );
  NAND2_X1 U8136 ( .A1(P2_REG2_REG_9__SCAN_IN), .A2(n6507), .ZN(n6459) );
  INV_X1 U8137 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n6452) );
  MUX2_X1 U8138 ( .A(n6452), .B(P2_REG2_REG_9__SCAN_IN), .S(n6507), .Z(n6453)
         );
  INV_X1 U8139 ( .A(n6453), .ZN(n6509) );
  INV_X1 U8140 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n6458) );
  MUX2_X1 U8141 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n6458), .S(n6495), .Z(n6497)
         );
  NAND2_X1 U8142 ( .A1(n9757), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6457) );
  MUX2_X1 U8143 ( .A(n5118), .B(P2_REG2_REG_7__SCAN_IN), .S(n9757), .Z(n6454)
         );
  INV_X1 U8144 ( .A(n6454), .ZN(n9762) );
  OAI21_X1 U8145 ( .B1(n6456), .B2(n6466), .A(n6455), .ZN(n9763) );
  NAND2_X1 U8146 ( .A1(n9762), .A2(n9763), .ZN(n9761) );
  NAND2_X1 U8147 ( .A1(n6457), .A2(n9761), .ZN(n6498) );
  NAND2_X1 U8148 ( .A1(n6497), .A2(n6498), .ZN(n6496) );
  OAI21_X1 U8149 ( .B1(n6468), .B2(n6458), .A(n6496), .ZN(n6510) );
  NAND2_X1 U8150 ( .A1(n6509), .A2(n6510), .ZN(n6508) );
  NAND2_X1 U8151 ( .A1(n6459), .A2(n6508), .ZN(n9776) );
  NAND2_X1 U8152 ( .A1(n9775), .A2(n9776), .ZN(n9774) );
  NAND2_X1 U8153 ( .A1(n6460), .A2(n9774), .ZN(n6461) );
  NOR2_X1 U8154 ( .A1(n6461), .A2(n6462), .ZN(n6526) );
  AOI21_X1 U8155 ( .B1(n6462), .B2(n6461), .A(n6526), .ZN(n6479) );
  INV_X1 U8156 ( .A(n9783), .ZN(n7579) );
  NAND2_X1 U8157 ( .A1(n9770), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n6470) );
  INV_X1 U8158 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n6463) );
  MUX2_X1 U8159 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n6463), .S(n9770), .Z(n9772)
         );
  INV_X1 U8160 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n9952) );
  MUX2_X1 U8161 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n9952), .S(n6507), .Z(n6502)
         );
  INV_X1 U8162 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n9950) );
  MUX2_X1 U8163 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n9950), .S(n6495), .Z(n6490)
         );
  NAND2_X1 U8164 ( .A1(n9757), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6467) );
  INV_X1 U8165 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6464) );
  MUX2_X1 U8166 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n6464), .S(n9757), .Z(n9759)
         );
  OAI21_X1 U8167 ( .B1(n6410), .B2(n6466), .A(n6465), .ZN(n9760) );
  NAND2_X1 U8168 ( .A1(n9759), .A2(n9760), .ZN(n9758) );
  NAND2_X1 U8169 ( .A1(n6467), .A2(n9758), .ZN(n6491) );
  NAND2_X1 U8170 ( .A1(n6490), .A2(n6491), .ZN(n6489) );
  OAI21_X1 U8171 ( .B1(n6468), .B2(n9950), .A(n6489), .ZN(n6503) );
  NAND2_X1 U8172 ( .A1(n6502), .A2(n6503), .ZN(n6501) );
  OAI21_X1 U8173 ( .B1(n6469), .B2(n9952), .A(n6501), .ZN(n9773) );
  NAND2_X1 U8174 ( .A1(n9772), .A2(n9773), .ZN(n9771) );
  NAND2_X1 U8175 ( .A1(n6470), .A2(n9771), .ZN(n6473) );
  INV_X1 U8176 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n6471) );
  MUX2_X1 U8177 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n6471), .S(n6524), .Z(n6472)
         );
  NAND2_X1 U8178 ( .A1(n6472), .A2(n6473), .ZN(n6520) );
  OAI211_X1 U8179 ( .C1(n6473), .C2(n6472), .A(n9786), .B(n6520), .ZN(n6476)
         );
  NOR2_X1 U8180 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5179), .ZN(n6474) );
  AOI21_X1 U8181 ( .B1(n9781), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n6474), .ZN(
        n6475) );
  OAI211_X1 U8182 ( .C1(n9734), .C2(n6521), .A(n6476), .B(n6475), .ZN(n6477)
         );
  INV_X1 U8183 ( .A(n6477), .ZN(n6478) );
  OAI21_X1 U8184 ( .B1(n6479), .B2(n7579), .A(n6478), .ZN(P2_U3256) );
  NAND2_X1 U8185 ( .A1(n8444), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n6480) );
  OAI21_X1 U8186 ( .B1(n8363), .B2(n8444), .A(n6480), .ZN(P2_U3574) );
  INV_X1 U8187 ( .A(n6481), .ZN(n6483) );
  INV_X1 U8188 ( .A(n6649), .ZN(n6877) );
  OAI222_X1 U8189 ( .A1(n7714), .A2(n6482), .B1(n8844), .B2(n6483), .C1(n6877), 
        .C2(P2_U3152), .ZN(P2_U3344) );
  INV_X1 U8190 ( .A(n7088), .ZN(n8966) );
  OAI222_X1 U8191 ( .A1(n7688), .A2(n6484), .B1(n9391), .B2(n6483), .C1(n8966), 
        .C2(P1_U3084), .ZN(P1_U3339) );
  INV_X1 U8192 ( .A(n6485), .ZN(n6487) );
  OAI222_X1 U8193 ( .A1(n7688), .A2(n6486), .B1(n7399), .B2(n6487), .C1(n7087), 
        .C2(P1_U3084), .ZN(P1_U3340) );
  INV_X1 U8194 ( .A(n6577), .ZN(n6648) );
  OAI222_X1 U8195 ( .A1(n7714), .A2(n6488), .B1(n8844), .B2(n6487), .C1(n6648), 
        .C2(P2_U3152), .ZN(P2_U3345) );
  INV_X1 U8196 ( .A(n9734), .ZN(n9791) );
  INV_X1 U8197 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n6493) );
  OAI211_X1 U8198 ( .C1(n6491), .C2(n6490), .A(n9786), .B(n6489), .ZN(n6492)
         );
  NAND2_X1 U8199 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3152), .ZN(n6892) );
  OAI211_X1 U8200 ( .C1(n8464), .C2(n6493), .A(n6492), .B(n6892), .ZN(n6494)
         );
  AOI21_X1 U8201 ( .B1(n6495), .B2(n9791), .A(n6494), .ZN(n6500) );
  OAI211_X1 U8202 ( .C1(n6498), .C2(n6497), .A(n9783), .B(n6496), .ZN(n6499)
         );
  NAND2_X1 U8203 ( .A1(n6500), .A2(n6499), .ZN(P2_U3253) );
  INV_X1 U8204 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n6505) );
  OAI211_X1 U8205 ( .C1(n6503), .C2(n6502), .A(n9786), .B(n6501), .ZN(n6504)
         );
  NAND2_X1 U8206 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3152), .ZN(n6987) );
  OAI211_X1 U8207 ( .C1(n8464), .C2(n6505), .A(n6504), .B(n6987), .ZN(n6506)
         );
  AOI21_X1 U8208 ( .B1(n6507), .B2(n9791), .A(n6506), .ZN(n6512) );
  OAI211_X1 U8209 ( .C1(n6510), .C2(n6509), .A(n9783), .B(n6508), .ZN(n6511)
         );
  NAND2_X1 U8210 ( .A1(n6512), .A2(n6511), .ZN(P2_U3254) );
  INV_X1 U8211 ( .A(n6513), .ZN(n6599) );
  AOI22_X1 U8212 ( .A1(n9566), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n9389), .ZN(n6514) );
  OAI21_X1 U8213 ( .B1(n6599), .B2(n9391), .A(n6514), .ZN(P1_U3337) );
  INV_X1 U8214 ( .A(n9640), .ZN(n8109) );
  OAI21_X1 U8215 ( .B1(n6517), .B2(n6515), .A(n6516), .ZN(n9480) );
  NAND2_X1 U8216 ( .A1(n9480), .A2(n8901), .ZN(n6519) );
  AOI22_X1 U8217 ( .A1(n8922), .A2(n7040), .B1(n6761), .B2(
        P1_REG3_REG_0__SCAN_IN), .ZN(n6518) );
  OAI211_X1 U8218 ( .C1(n8910), .C2(n8109), .A(n6519), .B(n6518), .ZN(P1_U3230) );
  OAI21_X1 U8219 ( .B1(n6521), .B2(n6471), .A(n6520), .ZN(n6523) );
  INV_X1 U8220 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n9957) );
  AOI22_X1 U8221 ( .A1(P2_REG1_REG_12__SCAN_IN), .A2(n6571), .B1(n6574), .B2(
        n9957), .ZN(n6522) );
  NOR2_X1 U8222 ( .A1(n6523), .A2(n6522), .ZN(n6570) );
  AOI21_X1 U8223 ( .B1(n6523), .B2(n6522), .A(n6570), .ZN(n6534) );
  NOR2_X1 U8224 ( .A1(n6524), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n6525) );
  NOR2_X1 U8225 ( .A1(n6526), .A2(n6525), .ZN(n6529) );
  INV_X1 U8226 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n6527) );
  MUX2_X1 U8227 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n6527), .S(n6574), .Z(n6528)
         );
  NAND2_X1 U8228 ( .A1(n6528), .A2(n6529), .ZN(n6575) );
  OAI211_X1 U8229 ( .C1(n6529), .C2(n6528), .A(n9783), .B(n6575), .ZN(n6533)
         );
  NOR2_X1 U8230 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10078), .ZN(n6531) );
  NOR2_X1 U8231 ( .A1(n9734), .A2(n6571), .ZN(n6530) );
  AOI211_X1 U8232 ( .C1(n9781), .C2(P2_ADDR_REG_12__SCAN_IN), .A(n6531), .B(
        n6530), .ZN(n6532) );
  OAI211_X1 U8233 ( .C1(n6534), .C2(n9735), .A(n6533), .B(n6532), .ZN(P2_U3257) );
  INV_X1 U8234 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n6543) );
  INV_X1 U8235 ( .A(n6535), .ZN(n6539) );
  INV_X1 U8236 ( .A(n6536), .ZN(n6538) );
  MUX2_X1 U8237 ( .A(n6408), .B(P2_REG1_REG_5__SCAN_IN), .S(n6551), .Z(n6537)
         );
  NAND3_X1 U8238 ( .A1(n6539), .A2(n6538), .A3(n6537), .ZN(n6540) );
  NAND3_X1 U8239 ( .A1(n9786), .A2(n6541), .A3(n6540), .ZN(n6542) );
  NAND2_X1 U8240 ( .A1(P2_U3152), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n6863) );
  OAI211_X1 U8241 ( .C1(n6543), .C2(n8464), .A(n6542), .B(n6863), .ZN(n6550)
         );
  AND3_X1 U8242 ( .A1(n6546), .A2(n6545), .A3(n6544), .ZN(n6547) );
  NOR3_X1 U8243 ( .A1(n7579), .A2(n6548), .A3(n6547), .ZN(n6549) );
  AOI211_X1 U8244 ( .C1(n9791), .C2(n6551), .A(n6550), .B(n6549), .ZN(n6552)
         );
  INV_X1 U8245 ( .A(n6552), .ZN(P2_U3250) );
  INV_X1 U8246 ( .A(n6553), .ZN(n6555) );
  INV_X1 U8247 ( .A(n7004), .ZN(n6882) );
  OAI222_X1 U8248 ( .A1(n7714), .A2(n6554), .B1(n8844), .B2(n6555), .C1(
        P2_U3152), .C2(n6882), .ZN(P2_U3343) );
  INV_X1 U8249 ( .A(n9555), .ZN(n8970) );
  OAI222_X1 U8250 ( .A1(n7688), .A2(n6556), .B1(n9391), .B2(n6555), .C1(
        P1_U3084), .C2(n8970), .ZN(P1_U3338) );
  AOI21_X1 U8251 ( .B1(n6559), .B2(n6558), .A(n6557), .ZN(n6569) );
  INV_X1 U8252 ( .A(n9580), .ZN(n9595) );
  OAI21_X1 U8253 ( .B1(n6562), .B2(n6561), .A(n6560), .ZN(n6563) );
  AOI22_X1 U8254 ( .A1(n6564), .A2(n9567), .B1(n9595), .B2(n6563), .ZN(n6568)
         );
  INV_X1 U8255 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n6565) );
  NAND2_X1 U8256 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3084), .ZN(n7117) );
  OAI21_X1 U8257 ( .B1(n9609), .B2(n6565), .A(n7117), .ZN(n6566) );
  INV_X1 U8258 ( .A(n6566), .ZN(n6567) );
  OAI211_X1 U8259 ( .C1(n6569), .C2(n9605), .A(n6568), .B(n6567), .ZN(P1_U3248) );
  AOI21_X1 U8260 ( .B1(n9957), .B2(n6571), .A(n6570), .ZN(n6573) );
  INV_X1 U8261 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n6644) );
  AOI22_X1 U8262 ( .A1(P2_REG1_REG_13__SCAN_IN), .A2(n6648), .B1(n6577), .B2(
        n6644), .ZN(n6572) );
  NOR2_X1 U8263 ( .A1(n6573), .A2(n6572), .ZN(n6643) );
  AOI21_X1 U8264 ( .B1(n6573), .B2(n6572), .A(n6643), .ZN(n6586) );
  NAND2_X1 U8265 ( .A1(P2_REG2_REG_12__SCAN_IN), .A2(n6574), .ZN(n6576) );
  NAND2_X1 U8266 ( .A1(n6576), .A2(n6575), .ZN(n6579) );
  AOI22_X1 U8267 ( .A1(P2_REG2_REG_13__SCAN_IN), .A2(n6648), .B1(n6577), .B2(
        n5216), .ZN(n6578) );
  NOR2_X1 U8268 ( .A1(n6579), .A2(n6578), .ZN(n6647) );
  AOI21_X1 U8269 ( .B1(n6579), .B2(n6578), .A(n6647), .ZN(n6580) );
  NOR2_X1 U8270 ( .A1(n6580), .A2(n7579), .ZN(n6584) );
  NOR2_X1 U8271 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5213), .ZN(n6581) );
  AOI21_X1 U8272 ( .B1(n9781), .B2(P2_ADDR_REG_13__SCAN_IN), .A(n6581), .ZN(
        n6582) );
  OAI21_X1 U8273 ( .B1(n9734), .B2(n6648), .A(n6582), .ZN(n6583) );
  NOR2_X1 U8274 ( .A1(n6584), .A2(n6583), .ZN(n6585) );
  OAI21_X1 U8275 ( .B1(n6586), .B2(n9735), .A(n6585), .ZN(P2_U3258) );
  AOI21_X1 U8276 ( .B1(n6589), .B2(n6588), .A(n6587), .ZN(n6591) );
  INV_X1 U8277 ( .A(n9609), .ZN(n9535) );
  NAND2_X1 U8278 ( .A1(n9535), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n6590) );
  NAND2_X1 U8279 ( .A1(P1_U3084), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n7030) );
  OAI211_X1 U8280 ( .C1(n6591), .C2(n9605), .A(n6590), .B(n7030), .ZN(n6596)
         );
  AOI211_X1 U8281 ( .C1(n6594), .C2(n6593), .A(n6592), .B(n9580), .ZN(n6595)
         );
  AOI211_X1 U8282 ( .C1(n9567), .C2(n6597), .A(n6596), .B(n6595), .ZN(n6598)
         );
  INV_X1 U8283 ( .A(n6598), .ZN(P1_U3247) );
  OAI222_X1 U8284 ( .A1(n7714), .A2(n6600), .B1(n8844), .B2(n6599), .C1(n7571), 
        .C2(P2_U3152), .ZN(P2_U3342) );
  INV_X1 U8285 ( .A(n6601), .ZN(n6633) );
  AOI22_X1 U8286 ( .A1(n8975), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n9389), .ZN(n6602) );
  OAI21_X1 U8287 ( .B1(n6633), .B2(n9391), .A(n6602), .ZN(P1_U3336) );
  NOR2_X1 U8288 ( .A1(n6610), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6604) );
  NOR2_X1 U8289 ( .A1(n6604), .A2(n6603), .ZN(n6607) );
  INV_X1 U8290 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n9453) );
  AOI22_X1 U8291 ( .A1(n6805), .A2(n9453), .B1(P1_REG1_REG_10__SCAN_IN), .B2(
        n6605), .ZN(n6606) );
  NOR2_X1 U8292 ( .A1(n6607), .A2(n6606), .ZN(n6798) );
  AOI21_X1 U8293 ( .B1(n6607), .B2(n6606), .A(n6798), .ZN(n6617) );
  INV_X1 U8294 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n6608) );
  NAND2_X1 U8295 ( .A1(P1_U3084), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n7493) );
  OAI21_X1 U8296 ( .B1(n9609), .B2(n6608), .A(n7493), .ZN(n6615) );
  NAND2_X1 U8297 ( .A1(n6805), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6611) );
  OAI21_X1 U8298 ( .B1(n6805), .B2(P1_REG2_REG_10__SCAN_IN), .A(n6611), .ZN(
        n6612) );
  AOI211_X1 U8299 ( .C1(n6613), .C2(n6612), .A(n6804), .B(n9580), .ZN(n6614)
         );
  AOI211_X1 U8300 ( .C1(n9567), .C2(n6805), .A(n6615), .B(n6614), .ZN(n6616)
         );
  OAI21_X1 U8301 ( .B1(n6617), .B2(n9605), .A(n6616), .ZN(P1_U3251) );
  INV_X1 U8302 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n6622) );
  OAI211_X1 U8303 ( .C1(n6620), .C2(n6619), .A(n9595), .B(n6618), .ZN(n6621)
         );
  OAI21_X1 U8304 ( .B1(n6622), .B2(n9609), .A(n6621), .ZN(n6629) );
  INV_X1 U8305 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n6627) );
  INV_X1 U8306 ( .A(n9605), .ZN(n9585) );
  OAI211_X1 U8307 ( .C1(n6625), .C2(n6624), .A(n9585), .B(n6623), .ZN(n6626)
         );
  OAI21_X1 U8308 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n6627), .A(n6626), .ZN(n6628) );
  AOI211_X1 U8309 ( .C1(n9567), .C2(n6630), .A(n6629), .B(n6628), .ZN(n6631)
         );
  INV_X1 U8310 ( .A(n6631), .ZN(P1_U3242) );
  OAI222_X1 U8311 ( .A1(P2_U3152), .A2(n7572), .B1(n8844), .B2(n6633), .C1(
        n6632), .C2(n7714), .ZN(P2_U3341) );
  INV_X1 U8312 ( .A(n6634), .ZN(n6756) );
  AOI21_X1 U8313 ( .B1(n6635), .B2(n6753), .A(n6636), .ZN(n6637) );
  AOI21_X1 U8314 ( .B1(n6756), .B2(n6753), .A(n6637), .ZN(n6642) );
  NAND2_X1 U8315 ( .A1(n7038), .A2(n9695), .ZN(n9655) );
  AOI22_X1 U8316 ( .A1(n8938), .A2(n6638), .B1(n8922), .B2(n8957), .ZN(n6639)
         );
  OAI21_X1 U8317 ( .B1(n6761), .B2(n9655), .A(n6639), .ZN(n6640) );
  AOI21_X1 U8318 ( .B1(P1_REG3_REG_1__SCAN_IN), .B2(n6761), .A(n6640), .ZN(
        n6641) );
  OAI21_X1 U8319 ( .B1(n6642), .B2(n8944), .A(n6641), .ZN(P1_U3220) );
  AOI21_X1 U8320 ( .B1(n6644), .B2(n6648), .A(n6643), .ZN(n6646) );
  INV_X1 U8321 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n6878) );
  AOI22_X1 U8322 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n6877), .B1(n6649), .B2(
        n6878), .ZN(n6645) );
  NOR2_X1 U8323 ( .A1(n6646), .A2(n6645), .ZN(n6876) );
  AOI21_X1 U8324 ( .B1(n6646), .B2(n6645), .A(n6876), .ZN(n6658) );
  AOI21_X1 U8325 ( .B1(n5216), .B2(n6648), .A(n6647), .ZN(n6651) );
  AOI22_X1 U8326 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n6877), .B1(n6649), .B2(
        n5233), .ZN(n6650) );
  NOR2_X1 U8327 ( .A1(n6651), .A2(n6650), .ZN(n6874) );
  AOI21_X1 U8328 ( .B1(n6651), .B2(n6650), .A(n6874), .ZN(n6652) );
  NOR2_X1 U8329 ( .A1(n6652), .A2(n7579), .ZN(n6656) );
  NOR2_X1 U8330 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10091), .ZN(n6653) );
  AOI21_X1 U8331 ( .B1(n9781), .B2(P2_ADDR_REG_14__SCAN_IN), .A(n6653), .ZN(
        n6654) );
  OAI21_X1 U8332 ( .B1(n9734), .B2(n6877), .A(n6654), .ZN(n6655) );
  NOR2_X1 U8333 ( .A1(n6656), .A2(n6655), .ZN(n6657) );
  OAI21_X1 U8334 ( .B1(n6658), .B2(n9735), .A(n6657), .ZN(P2_U3259) );
  INV_X1 U8335 ( .A(n6910), .ZN(n6659) );
  INV_X1 U8336 ( .A(n6670), .ZN(n6664) );
  NOR2_X1 U8337 ( .A1(n6664), .A2(n9868), .ZN(n6694) );
  OR2_X1 U8338 ( .A1(n9880), .A2(n7983), .ZN(n6916) );
  INV_X1 U8339 ( .A(n6916), .ZN(n6661) );
  NAND2_X1 U8340 ( .A1(n6694), .A2(n6661), .ZN(n6662) );
  NAND2_X1 U8341 ( .A1(n6664), .A2(n6663), .ZN(n6667) );
  AND3_X1 U8342 ( .A1(n6665), .A2(n9871), .A3(n6909), .ZN(n6666) );
  NAND2_X1 U8343 ( .A1(n6667), .A2(n6666), .ZN(n6707) );
  NAND2_X1 U8344 ( .A1(n6707), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8411) );
  NAND2_X1 U8345 ( .A1(P2_U3152), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n9742) );
  INV_X1 U8346 ( .A(n6668), .ZN(n8001) );
  NOR2_X1 U8347 ( .A1(n9868), .A2(n8001), .ZN(n6669) );
  NAND2_X1 U8348 ( .A1(n6670), .A2(n6669), .ZN(n8417) );
  NAND2_X1 U8349 ( .A1(n6687), .A2(n8545), .ZN(n6671) );
  OAI21_X1 U8350 ( .B1(n6865), .B2(n9848), .A(n6671), .ZN(n6773) );
  NAND2_X1 U8351 ( .A1(n8364), .A2(n6773), .ZN(n6672) );
  OAI211_X1 U8352 ( .C1(n8411), .C2(P2_REG3_REG_3__SCAN_IN), .A(n9742), .B(
        n6672), .ZN(n6697) );
  INV_X1 U8353 ( .A(n6680), .ZN(n6677) );
  NAND2_X1 U8354 ( .A1(n9880), .A2(n6674), .ZN(n7998) );
  NAND2_X1 U8355 ( .A1(n6677), .A2(n6678), .ZN(n6681) );
  INV_X1 U8356 ( .A(n6678), .ZN(n6679) );
  NAND2_X1 U8357 ( .A1(n6680), .A2(n6679), .ZN(n6685) );
  NAND2_X1 U8358 ( .A1(n6681), .A2(n6685), .ZN(n6714) );
  INV_X1 U8359 ( .A(n6714), .ZN(n6684) );
  INV_X1 U8360 ( .A(n6717), .ZN(n6683) );
  NAND2_X1 U8361 ( .A1(n6684), .A2(n6683), .ZN(n6715) );
  NAND2_X1 U8362 ( .A1(n6715), .A2(n6685), .ZN(n6722) );
  XNOR2_X1 U8363 ( .A(n9887), .B(n4296), .ZN(n6689) );
  NAND2_X1 U8364 ( .A1(n6687), .A2(n6682), .ZN(n6688) );
  XNOR2_X1 U8365 ( .A(n6689), .B(n6688), .ZN(n6721) );
  XNOR2_X1 U8366 ( .A(n7225), .B(n7375), .ZN(n6735) );
  NAND2_X1 U8367 ( .A1(n8443), .A2(n6682), .ZN(n6734) );
  XNOR2_X1 U8368 ( .A(n6735), .B(n6734), .ZN(n6732) );
  XNOR2_X1 U8369 ( .A(n6691), .B(n6732), .ZN(n6695) );
  AND2_X1 U8370 ( .A1(n9937), .A2(n6692), .ZN(n6693) );
  NOR2_X1 U8371 ( .A1(n6695), .A2(n8422), .ZN(n6696) );
  AOI211_X1 U8372 ( .C1(n6768), .C2(n8420), .A(n6697), .B(n6696), .ZN(n6698)
         );
  INV_X1 U8373 ( .A(n6698), .ZN(P2_U3220) );
  OAI21_X1 U8374 ( .B1(n7803), .B2(n6700), .A(n6699), .ZN(n7103) );
  AOI211_X1 U8375 ( .C1(n6972), .C2(n7102), .A(n6682), .B(n6920), .ZN(n7104)
         );
  INV_X1 U8376 ( .A(n6687), .ZN(n6703) );
  INV_X1 U8377 ( .A(n6701), .ZN(n6708) );
  INV_X1 U8378 ( .A(n9818), .ZN(n9843) );
  INV_X1 U8379 ( .A(n6969), .ZN(n6710) );
  XNOR2_X1 U8380 ( .A(n7803), .B(n6710), .ZN(n6702) );
  OAI222_X1 U8381 ( .A1(n9848), .A2(n6703), .B1(n9846), .B2(n6708), .C1(n9843), 
        .C2(n6702), .ZN(n7109) );
  AOI211_X1 U8382 ( .C1(n9941), .C2(n7103), .A(n7104), .B(n7109), .ZN(n6906)
         );
  OAI22_X1 U8383 ( .A1(n8777), .A2(n6903), .B1(n9959), .B2(n6704), .ZN(n6705)
         );
  INV_X1 U8384 ( .A(n6705), .ZN(n6706) );
  OAI21_X1 U8385 ( .B1(n6906), .B2(n9956), .A(n6706), .ZN(P2_U3521) );
  INV_X1 U8386 ( .A(n6673), .ZN(n6713) );
  NAND2_X1 U8387 ( .A1(n8364), .A2(n8547), .ZN(n8403) );
  OR2_X1 U8388 ( .A1(n6707), .A2(P2_U3152), .ZN(n6723) );
  AOI22_X1 U8389 ( .A1(n8420), .A2(n6972), .B1(P2_REG3_REG_0__SCAN_IN), .B2(
        n6723), .ZN(n6712) );
  NOR2_X1 U8390 ( .A1(n6708), .A2(n6972), .ZN(n7844) );
  MUX2_X1 U8391 ( .A(n6972), .B(n7844), .S(n6682), .Z(n6709) );
  INV_X1 U8392 ( .A(n8422), .ZN(n8352) );
  OAI21_X1 U8393 ( .B1(n6710), .B2(n6709), .A(n8352), .ZN(n6711) );
  OAI211_X1 U8394 ( .C1(n6713), .C2(n8403), .A(n6712), .B(n6711), .ZN(P2_U3234) );
  INV_X1 U8395 ( .A(n6715), .ZN(n6716) );
  AOI21_X1 U8396 ( .B1(n6714), .B2(n6717), .A(n6716), .ZN(n6720) );
  NAND2_X1 U8397 ( .A1(n8364), .A2(n8545), .ZN(n8404) );
  INV_X1 U8398 ( .A(n8404), .ZN(n7680) );
  INV_X1 U8399 ( .A(n8403), .ZN(n8357) );
  AOI22_X1 U8400 ( .A1(n7680), .A2(n6701), .B1(n8357), .B2(n6687), .ZN(n6719)
         );
  AOI22_X1 U8401 ( .A1(n8420), .A2(n7102), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n6723), .ZN(n6718) );
  OAI211_X1 U8402 ( .C1(n6720), .C2(n8422), .A(n6719), .B(n6718), .ZN(P2_U3224) );
  XNOR2_X1 U8403 ( .A(n6722), .B(n6721), .ZN(n6726) );
  AOI22_X1 U8404 ( .A1(n7680), .A2(n6673), .B1(n8357), .B2(n8443), .ZN(n6725)
         );
  AOI22_X1 U8405 ( .A1(n8420), .A2(n6924), .B1(P2_REG3_REG_2__SCAN_IN), .B2(
        n6723), .ZN(n6724) );
  OAI211_X1 U8406 ( .C1(n6726), .C2(n8422), .A(n6725), .B(n6724), .ZN(P2_U3239) );
  NAND2_X1 U8407 ( .A1(n8442), .A2(n6682), .ZN(n6727) );
  XNOR2_X1 U8408 ( .A(n6960), .B(n7375), .ZN(n6728) );
  NAND2_X1 U8409 ( .A1(n6727), .A2(n6728), .ZN(n6826) );
  INV_X1 U8410 ( .A(n6727), .ZN(n6730) );
  INV_X1 U8411 ( .A(n6728), .ZN(n6729) );
  NAND2_X1 U8412 ( .A1(n6730), .A2(n6729), .ZN(n6731) );
  NAND2_X1 U8413 ( .A1(n6826), .A2(n6731), .ZN(n6743) );
  NAND2_X1 U8414 ( .A1(n6733), .A2(n6732), .ZN(n6738) );
  INV_X1 U8415 ( .A(n6734), .ZN(n6736) );
  NAND2_X1 U8416 ( .A1(n6736), .A2(n6735), .ZN(n6737) );
  NAND2_X1 U8417 ( .A1(n6738), .A2(n6737), .ZN(n6742) );
  INV_X1 U8418 ( .A(n6742), .ZN(n6740) );
  INV_X1 U8419 ( .A(n6827), .ZN(n6741) );
  AOI21_X1 U8420 ( .B1(n6743), .B2(n6742), .A(n6741), .ZN(n6748) );
  OAI21_X1 U8421 ( .B1(n8403), .B2(n6951), .A(n6744), .ZN(n6746) );
  OAI22_X1 U8422 ( .A1(n8404), .A2(n6950), .B1(n8411), .B2(n6958), .ZN(n6745)
         );
  AOI211_X1 U8423 ( .C1(n6960), .C2(n8420), .A(n6746), .B(n6745), .ZN(n6747)
         );
  OAI21_X1 U8424 ( .B1(n6748), .B2(n8422), .A(n6747), .ZN(P2_U3232) );
  INV_X1 U8425 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n6750) );
  INV_X1 U8426 ( .A(n6749), .ZN(n6751) );
  INV_X1 U8427 ( .A(n8446), .ZN(n8451) );
  OAI222_X1 U8428 ( .A1(n7714), .A2(n6750), .B1(n8844), .B2(n6751), .C1(
        P2_U3152), .C2(n8451), .ZN(P2_U3340) );
  INV_X1 U8429 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n6752) );
  INV_X1 U8430 ( .A(n8979), .ZN(n9600) );
  OAI222_X1 U8431 ( .A1(n7688), .A2(n6752), .B1(n9391), .B2(n6751), .C1(
        P1_U3084), .C2(n9600), .ZN(P1_U3335) );
  INV_X1 U8432 ( .A(n6753), .ZN(n6754) );
  NOR3_X1 U8433 ( .A1(n6756), .A2(n6755), .A3(n6754), .ZN(n6759) );
  INV_X1 U8434 ( .A(n6757), .ZN(n6758) );
  OAI21_X1 U8435 ( .B1(n6759), .B2(n6758), .A(n8901), .ZN(n6763) );
  INV_X1 U8436 ( .A(n7040), .ZN(n7155) );
  OAI22_X1 U8437 ( .A1(n7142), .A2(n8936), .B1(n8905), .B2(n7155), .ZN(n6760)
         );
  AOI21_X1 U8438 ( .B1(P1_REG3_REG_2__SCAN_IN), .B2(n6761), .A(n6760), .ZN(
        n6762) );
  OAI211_X1 U8439 ( .C1(n7199), .C2(n8910), .A(n6763), .B(n6762), .ZN(P1_U3235) );
  INV_X1 U8440 ( .A(n6764), .ZN(n9920) );
  OR2_X1 U8441 ( .A1(n6765), .A2(n6770), .ZN(n6766) );
  NAND2_X1 U8442 ( .A1(n6767), .A2(n6766), .ZN(n7229) );
  AOI21_X1 U8443 ( .B1(n6919), .B2(n6768), .A(n6682), .ZN(n6769) );
  AND2_X1 U8444 ( .A1(n6769), .A2(n6954), .ZN(n7223) );
  INV_X1 U8445 ( .A(n8679), .ZN(n9852) );
  NAND2_X1 U8446 ( .A1(n7229), .A2(n9852), .ZN(n6776) );
  NAND3_X1 U8447 ( .A1(n6907), .A2(n6770), .A3(n7854), .ZN(n6771) );
  NAND2_X1 U8448 ( .A1(n6772), .A2(n6771), .ZN(n6774) );
  AOI21_X1 U8449 ( .B1(n6774), .B2(n9818), .A(n6773), .ZN(n6775) );
  NAND2_X1 U8450 ( .A1(n6776), .A2(n6775), .ZN(n7226) );
  AOI211_X1 U8451 ( .C1(n9920), .C2(n7229), .A(n7223), .B(n7226), .ZN(n6901)
         );
  OAI22_X1 U8452 ( .A1(n8777), .A2(n7225), .B1(n9959), .B2(n6400), .ZN(n6777)
         );
  INV_X1 U8453 ( .A(n6777), .ZN(n6778) );
  OAI21_X1 U8454 ( .B1(n6901), .B2(n9956), .A(n6778), .ZN(P2_U3523) );
  INV_X1 U8455 ( .A(n6779), .ZN(n6781) );
  OAI222_X1 U8456 ( .A1(n7714), .A2(n6780), .B1(n8844), .B2(n6781), .C1(n8682), 
        .C2(P2_U3152), .ZN(P2_U3339) );
  OAI222_X1 U8457 ( .A1(n7688), .A2(n6782), .B1(n9391), .B2(n6781), .C1(
        P1_U3084), .C2(n8985), .ZN(P1_U3334) );
  NAND2_X1 U8458 ( .A1(n8444), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n6783) );
  OAI21_X1 U8459 ( .B1(n6784), .B2(n8444), .A(n6783), .ZN(P2_U3581) );
  NAND2_X1 U8460 ( .A1(n8444), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n6785) );
  OAI21_X1 U8461 ( .B1(n8412), .B2(n8444), .A(n6785), .ZN(P2_U3579) );
  INV_X1 U8462 ( .A(n9623), .ZN(n9679) );
  AND2_X1 U8463 ( .A1(n6786), .A2(n6787), .ZN(n6790) );
  OAI211_X1 U8464 ( .C1(n6790), .C2(n6789), .A(n8901), .B(n6788), .ZN(n6796)
         );
  INV_X1 U8465 ( .A(n6791), .ZN(n9621) );
  INV_X1 U8466 ( .A(n9614), .ZN(n7148) );
  AND2_X1 U8467 ( .A1(P1_U3084), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n9507) );
  AOI21_X1 U8468 ( .B1(n8938), .B2(n6792), .A(n9507), .ZN(n6793) );
  OAI21_X1 U8469 ( .B1(n8936), .B2(n7148), .A(n6793), .ZN(n6794) );
  AOI21_X1 U8470 ( .B1(n9621), .B2(n8907), .A(n6794), .ZN(n6795) );
  OAI211_X1 U8471 ( .C1(n9679), .C2(n8910), .A(n6796), .B(n6795), .ZN(P1_U3228) );
  NOR2_X1 U8472 ( .A1(n6805), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6797) );
  NOR2_X1 U8473 ( .A1(n6798), .A2(n6797), .ZN(n9539) );
  MUX2_X1 U8474 ( .A(n6799), .B(P1_REG1_REG_11__SCAN_IN), .S(n9536), .Z(n9538)
         );
  NOR2_X1 U8475 ( .A1(n9539), .A2(n9538), .ZN(n9537) );
  AOI21_X1 U8476 ( .B1(n6799), .B2(n6803), .A(n9537), .ZN(n6801) );
  AOI22_X1 U8477 ( .A1(P1_REG1_REG_12__SCAN_IN), .A2(n6931), .B1(n6936), .B2(
        n5928), .ZN(n6800) );
  NOR2_X1 U8478 ( .A1(n6801), .A2(n6800), .ZN(n6930) );
  AOI21_X1 U8479 ( .B1(n6801), .B2(n6800), .A(n6930), .ZN(n6812) );
  INV_X1 U8480 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n6802) );
  NAND2_X1 U8481 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_U3084), .ZN(n7539) );
  OAI21_X1 U8482 ( .B1(n9609), .B2(n6802), .A(n7539), .ZN(n6810) );
  AOI22_X1 U8483 ( .A1(P1_REG2_REG_11__SCAN_IN), .A2(n9536), .B1(n6803), .B2(
        n5947), .ZN(n9543) );
  OAI21_X1 U8484 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n9536), .A(n9541), .ZN(
        n6808) );
  NAND2_X1 U8485 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n6936), .ZN(n6806) );
  OAI21_X1 U8486 ( .B1(n6936), .B2(P1_REG2_REG_12__SCAN_IN), .A(n6806), .ZN(
        n6807) );
  NOR2_X1 U8487 ( .A1(n6807), .A2(n6808), .ZN(n6935) );
  AOI211_X1 U8488 ( .C1(n6808), .C2(n6807), .A(n6935), .B(n9580), .ZN(n6809)
         );
  AOI211_X1 U8489 ( .C1(n9567), .C2(n6936), .A(n6810), .B(n6809), .ZN(n6811)
         );
  OAI21_X1 U8490 ( .B1(n6812), .B2(n9605), .A(n6811), .ZN(P1_U3253) );
  OAI21_X1 U8491 ( .B1(n6814), .B2(n6813), .A(n6786), .ZN(n6815) );
  NAND2_X1 U8492 ( .A1(n6815), .A2(n8901), .ZN(n6820) );
  INV_X1 U8493 ( .A(n9668), .ZN(n7145) );
  NAND2_X1 U8494 ( .A1(P1_U3084), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9435) );
  INV_X1 U8495 ( .A(n9435), .ZN(n6816) );
  AOI21_X1 U8496 ( .B1(n8938), .B2(n8957), .A(n6816), .ZN(n6817) );
  OAI21_X1 U8497 ( .B1(n8936), .B2(n7145), .A(n6817), .ZN(n6818) );
  AOI21_X1 U8498 ( .B1(n5816), .B2(n8907), .A(n6818), .ZN(n6819) );
  OAI211_X1 U8499 ( .C1(n7285), .C2(n8910), .A(n6820), .B(n6819), .ZN(P1_U3216) );
  AND2_X1 U8500 ( .A1(n8440), .A2(n6682), .ZN(n6821) );
  XNOR2_X1 U8501 ( .A(n9897), .B(n4296), .ZN(n6822) );
  NAND2_X1 U8502 ( .A1(n6821), .A2(n6822), .ZN(n6825) );
  INV_X1 U8503 ( .A(n6821), .ZN(n6824) );
  INV_X1 U8504 ( .A(n6822), .ZN(n6823) );
  NAND2_X1 U8505 ( .A1(n6824), .A2(n6823), .ZN(n6855) );
  AND2_X1 U8506 ( .A1(n6825), .A2(n6855), .ZN(n6838) );
  NAND2_X1 U8507 ( .A1(n8441), .A2(n6682), .ZN(n6830) );
  XNOR2_X1 U8508 ( .A(n6828), .B(n7375), .ZN(n6831) );
  XNOR2_X1 U8509 ( .A(n6830), .B(n6831), .ZN(n6861) );
  INV_X1 U8510 ( .A(n6861), .ZN(n6829) );
  INV_X1 U8511 ( .A(n6830), .ZN(n6833) );
  INV_X1 U8512 ( .A(n6831), .ZN(n6832) );
  NAND2_X1 U8513 ( .A1(n6833), .A2(n6832), .ZN(n6834) );
  AND2_X1 U8514 ( .A1(n6836), .A2(n6834), .ZN(n6837) );
  AND2_X1 U8515 ( .A1(n6838), .A2(n6834), .ZN(n6835) );
  NAND2_X1 U8516 ( .A1(n6836), .A2(n6835), .ZN(n6856) );
  OAI21_X1 U8517 ( .B1(n6838), .B2(n6837), .A(n6856), .ZN(n6844) );
  INV_X1 U8518 ( .A(n6839), .ZN(n7777) );
  OAI22_X1 U8519 ( .A1(n8404), .A2(n6951), .B1(n8411), .B2(n7777), .ZN(n6843)
         );
  NAND2_X1 U8520 ( .A1(n8420), .A2(n9897), .ZN(n6841) );
  OAI211_X1 U8521 ( .C1(n8403), .C2(n9847), .A(n6841), .B(n6840), .ZN(n6842)
         );
  AOI211_X1 U8522 ( .C1(n6844), .C2(n8352), .A(n6843), .B(n6842), .ZN(n6845)
         );
  INV_X1 U8523 ( .A(n6845), .ZN(P2_U3241) );
  INV_X1 U8524 ( .A(n9941), .ZN(n9932) );
  NAND2_X1 U8525 ( .A1(n6946), .A2(n6846), .ZN(n6847) );
  XNOR2_X1 U8526 ( .A(n6847), .B(n6851), .ZN(n7217) );
  OR2_X1 U8527 ( .A1(n6948), .A2(n7807), .ZN(n6849) );
  AND2_X1 U8528 ( .A1(n6849), .A2(n7835), .ZN(n6850) );
  NAND2_X1 U8529 ( .A1(n6849), .A2(n6848), .ZN(n7780) );
  OAI21_X1 U8530 ( .B1(n6851), .B2(n6850), .A(n7780), .ZN(n6852) );
  AOI222_X1 U8531 ( .A1(n9818), .A2(n6852), .B1(n8440), .B2(n8547), .C1(n8442), 
        .C2(n8545), .ZN(n7208) );
  OAI211_X1 U8532 ( .C1(n7212), .C2(n6955), .A(n4380), .B(n7321), .ZN(n7209)
         );
  OAI211_X1 U8533 ( .C1(n9932), .C2(n7217), .A(n7208), .B(n7209), .ZN(n6966)
         );
  OAI22_X1 U8534 ( .A1(n8777), .A2(n7212), .B1(n9959), .B2(n6408), .ZN(n6853)
         );
  AOI21_X1 U8535 ( .B1(n6966), .B2(n9959), .A(n6853), .ZN(n6854) );
  INV_X1 U8536 ( .A(n6854), .ZN(P2_U3525) );
  NAND2_X1 U8537 ( .A1(n6856), .A2(n6855), .ZN(n6890) );
  NAND2_X1 U8538 ( .A1(n8439), .A2(n6682), .ZN(n6887) );
  XNOR2_X1 U8539 ( .A(n7126), .B(n7375), .ZN(n6888) );
  XNOR2_X1 U8540 ( .A(n6887), .B(n6888), .ZN(n6889) );
  XNOR2_X1 U8541 ( .A(n6890), .B(n6889), .ZN(n6860) );
  INV_X1 U8542 ( .A(n8411), .ZN(n8375) );
  NAND2_X1 U8543 ( .A1(P2_U3152), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n9755) );
  OAI21_X1 U8544 ( .B1(n8403), .B2(n7876), .A(n9755), .ZN(n6858) );
  INV_X1 U8545 ( .A(n8440), .ZN(n6864) );
  OAI22_X1 U8546 ( .A1(n8360), .A2(n9904), .B1(n6864), .B2(n8404), .ZN(n6857)
         );
  AOI211_X1 U8547 ( .C1(n7125), .C2(n8375), .A(n6858), .B(n6857), .ZN(n6859)
         );
  OAI21_X1 U8548 ( .B1(n6860), .B2(n8422), .A(n6859), .ZN(P2_U3215) );
  XNOR2_X1 U8549 ( .A(n6862), .B(n6861), .ZN(n6869) );
  OAI21_X1 U8550 ( .B1(n8403), .B2(n6864), .A(n6863), .ZN(n6867) );
  OAI22_X1 U8551 ( .A1(n8360), .A2(n7212), .B1(n6865), .B2(n8404), .ZN(n6866)
         );
  AOI211_X1 U8552 ( .C1(n7210), .C2(n8375), .A(n6867), .B(n6866), .ZN(n6868)
         );
  OAI21_X1 U8553 ( .B1(n6869), .B2(n8422), .A(n6868), .ZN(P2_U3229) );
  INV_X1 U8554 ( .A(n6870), .ZN(n6872) );
  OAI222_X1 U8555 ( .A1(n7688), .A2(n6871), .B1(n9391), .B2(n6872), .C1(n8201), 
        .C2(P1_U3084), .ZN(P1_U3333) );
  OAI222_X1 U8556 ( .A1(n7714), .A2(n6873), .B1(P2_U3152), .B2(n7983), .C1(
        n8844), .C2(n6872), .ZN(P2_U3338) );
  AOI21_X1 U8557 ( .B1(n5233), .B2(n6877), .A(n6874), .ZN(n7003) );
  XNOR2_X1 U8558 ( .A(n7004), .B(n7003), .ZN(n6875) );
  NOR2_X1 U8559 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n6875), .ZN(n7005) );
  AOI21_X1 U8560 ( .B1(P2_REG2_REG_15__SCAN_IN), .B2(n6875), .A(n7005), .ZN(
        n6886) );
  AOI21_X1 U8561 ( .B1(n6878), .B2(n6877), .A(n6876), .ZN(n6996) );
  XOR2_X1 U8562 ( .A(n7004), .B(n6996), .Z(n6879) );
  NAND2_X1 U8563 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n6879), .ZN(n6997) );
  OAI211_X1 U8564 ( .C1(n6879), .C2(P2_REG1_REG_15__SCAN_IN), .A(n9786), .B(
        n6997), .ZN(n6885) );
  AND2_X1 U8565 ( .A1(P2_U3152), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6880) );
  AOI21_X1 U8566 ( .B1(n9781), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n6880), .ZN(
        n6881) );
  OAI21_X1 U8567 ( .B1(n9734), .B2(n6882), .A(n6881), .ZN(n6883) );
  INV_X1 U8568 ( .A(n6883), .ZN(n6884) );
  OAI211_X1 U8569 ( .C1(n6886), .C2(n7579), .A(n6885), .B(n6884), .ZN(P2_U3260) );
  XNOR2_X1 U8570 ( .A(n9857), .B(n4296), .ZN(n6980) );
  NAND2_X1 U8571 ( .A1(n8438), .A2(n6682), .ZN(n6978) );
  XNOR2_X1 U8572 ( .A(n6980), .B(n6978), .ZN(n6976) );
  XNOR2_X1 U8573 ( .A(n6891), .B(n6976), .ZN(n6897) );
  OAI21_X1 U8574 ( .B1(n8403), .B2(n9849), .A(n6892), .ZN(n6895) );
  OAI22_X1 U8575 ( .A1(n8404), .A2(n9847), .B1(n8411), .B2(n6893), .ZN(n6894)
         );
  AOI211_X1 U8576 ( .C1(n9857), .C2(n8420), .A(n6895), .B(n6894), .ZN(n6896)
         );
  OAI21_X1 U8577 ( .B1(n6897), .B2(n8422), .A(n6896), .ZN(P2_U3223) );
  INV_X1 U8578 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n6898) );
  OAI22_X1 U8579 ( .A1(n8831), .A2(n7225), .B1(n9944), .B2(n6898), .ZN(n6899)
         );
  INV_X1 U8580 ( .A(n6899), .ZN(n6900) );
  OAI21_X1 U8581 ( .B1(n6901), .B2(n9942), .A(n6900), .ZN(P2_U3460) );
  INV_X1 U8582 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n6902) );
  OAI22_X1 U8583 ( .A1(n8831), .A2(n6903), .B1(n9944), .B2(n6902), .ZN(n6904)
         );
  INV_X1 U8584 ( .A(n6904), .ZN(n6905) );
  OAI21_X1 U8585 ( .B1(n6906), .B2(n9942), .A(n6905), .ZN(P2_U3454) );
  OAI21_X1 U8586 ( .B1(n7805), .B2(n7845), .A(n6907), .ZN(n6908) );
  AOI222_X1 U8587 ( .A1(n9818), .A2(n6908), .B1(n8443), .B2(n8547), .C1(n6673), 
        .C2(n8545), .ZN(n9886) );
  INV_X1 U8588 ( .A(n6909), .ZN(n6911) );
  OR3_X1 U8589 ( .A1(n6912), .A2(n6911), .A3(n6910), .ZN(n6913) );
  NOR2_X1 U8590 ( .A1(n6913), .A2(n9868), .ZN(n6914) );
  NAND2_X1 U8591 ( .A1(n6915), .A2(n6914), .ZN(n6917) );
  AND2_X2 U8592 ( .A1(n6917), .A2(n8556), .ZN(n9866) );
  NOR2_X2 U8593 ( .A1(n9855), .A2(n6916), .ZN(n9856) );
  INV_X1 U8594 ( .A(n6917), .ZN(n6918) );
  NAND2_X1 U8595 ( .A1(n6918), .A2(n8682), .ZN(n9832) );
  OAI211_X1 U8596 ( .C1(n6920), .C2(n9887), .A(n7321), .B(n6919), .ZN(n9885)
         );
  NAND2_X1 U8597 ( .A1(n9866), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6922) );
  NAND2_X1 U8598 ( .A1(n9854), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n6921) );
  OAI211_X1 U8599 ( .C1(n9832), .C2(n9885), .A(n6922), .B(n6921), .ZN(n6923)
         );
  AOI21_X1 U8600 ( .B1(n9856), .B2(n6924), .A(n6923), .ZN(n6929) );
  XNOR2_X1 U8601 ( .A(n6925), .B(n7805), .ZN(n9889) );
  OR2_X1 U8602 ( .A1(n6926), .A2(n8682), .ZN(n7186) );
  AND2_X1 U8603 ( .A1(n8679), .A2(n7186), .ZN(n6927) );
  NAND2_X1 U8604 ( .A1(n9889), .A2(n9834), .ZN(n6928) );
  OAI211_X1 U8605 ( .C1(n9886), .C2(n9855), .A(n6929), .B(n6928), .ZN(P2_U3294) );
  AOI21_X1 U8606 ( .B1(n5928), .B2(n6931), .A(n6930), .ZN(n6933) );
  INV_X1 U8607 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n9340) );
  AOI22_X1 U8608 ( .A1(P1_REG1_REG_13__SCAN_IN), .A2(n7087), .B1(n7084), .B2(
        n9340), .ZN(n6932) );
  NOR2_X1 U8609 ( .A1(n6933), .A2(n6932), .ZN(n7086) );
  AOI21_X1 U8610 ( .B1(n6933), .B2(n6932), .A(n7086), .ZN(n6943) );
  INV_X1 U8611 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n6934) );
  NAND2_X1 U8612 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3084), .ZN(n7527) );
  OAI21_X1 U8613 ( .B1(n9609), .B2(n6934), .A(n7527), .ZN(n6941) );
  NAND2_X1 U8614 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n7084), .ZN(n6937) );
  OAI21_X1 U8615 ( .B1(n7084), .B2(P1_REG2_REG_13__SCAN_IN), .A(n6937), .ZN(
        n6938) );
  AOI211_X1 U8616 ( .C1(n6939), .C2(n6938), .A(n7083), .B(n9580), .ZN(n6940)
         );
  AOI211_X1 U8617 ( .C1(n9567), .C2(n7084), .A(n6941), .B(n6940), .ZN(n6942)
         );
  OAI21_X1 U8618 ( .B1(n6943), .B2(n9605), .A(n6942), .ZN(P1_U3254) );
  INV_X1 U8619 ( .A(n6944), .ZN(n6975) );
  OAI222_X1 U8620 ( .A1(n7688), .A2(n6945), .B1(n7399), .B2(n6975), .C1(n8197), 
        .C2(P1_U3084), .ZN(P1_U3332) );
  OAI21_X1 U8621 ( .B1(n6947), .B2(n7807), .A(n6946), .ZN(n9894) );
  INV_X1 U8622 ( .A(n9894), .ZN(n6963) );
  XNOR2_X1 U8623 ( .A(n6948), .B(n7807), .ZN(n6949) );
  OAI222_X1 U8624 ( .A1(n9848), .A2(n6951), .B1(n9846), .B2(n6950), .C1(n6949), 
        .C2(n9843), .ZN(n9892) );
  INV_X1 U8625 ( .A(n9892), .ZN(n6952) );
  MUX2_X1 U8626 ( .A(n6953), .B(n6952), .S(n8579), .Z(n6962) );
  INV_X1 U8627 ( .A(n6954), .ZN(n6957) );
  INV_X1 U8628 ( .A(n6955), .ZN(n6956) );
  OAI211_X1 U8629 ( .C1(n9891), .C2(n6957), .A(n6956), .B(n7321), .ZN(n9890)
         );
  OAI22_X1 U8630 ( .A1(n9890), .A2(n9832), .B1(n6958), .B2(n8556), .ZN(n6959)
         );
  AOI21_X1 U8631 ( .B1(n9856), .B2(n6960), .A(n6959), .ZN(n6961) );
  OAI211_X1 U8632 ( .C1(n6963), .C2(n8709), .A(n6962), .B(n6961), .ZN(P2_U3292) );
  INV_X1 U8633 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n6964) );
  OAI22_X1 U8634 ( .A1(n8831), .A2(n7212), .B1(n9944), .B2(n6964), .ZN(n6965)
         );
  AOI21_X1 U8635 ( .B1(n6966), .B2(n9944), .A(n6965), .ZN(n6967) );
  INV_X1 U8636 ( .A(n6967), .ZN(P2_U3466) );
  INV_X1 U8637 ( .A(n7844), .ZN(n6968) );
  NAND2_X1 U8638 ( .A1(n6969), .A2(n6968), .ZN(n7806) );
  INV_X1 U8639 ( .A(n7806), .ZN(n9881) );
  AOI22_X1 U8640 ( .A1(n7806), .A2(n9818), .B1(n8547), .B2(n6673), .ZN(n9878)
         );
  INV_X1 U8641 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n6970) );
  OAI22_X1 U8642 ( .A1(n9878), .A2(n9866), .B1(n6970), .B2(n8556), .ZN(n6971)
         );
  AOI21_X1 U8643 ( .B1(P2_REG2_REG_0__SCAN_IN), .B2(n9855), .A(n6971), .ZN(
        n6974) );
  OR2_X1 U8644 ( .A1(n9832), .A2(n6682), .ZN(n7798) );
  INV_X1 U8645 ( .A(n7798), .ZN(n8707) );
  OAI21_X1 U8646 ( .B1(n8707), .B2(n9856), .A(n6972), .ZN(n6973) );
  OAI211_X1 U8647 ( .C1(n9881), .C2(n8709), .A(n6974), .B(n6973), .ZN(P2_U3296) );
  OAI222_X1 U8648 ( .A1(n7714), .A2(n10082), .B1(P2_U3152), .B2(n7831), .C1(
        n8844), .C2(n6975), .ZN(P2_U3337) );
  NAND2_X1 U8649 ( .A1(n6977), .A2(n6976), .ZN(n7068) );
  INV_X1 U8650 ( .A(n6978), .ZN(n6979) );
  NAND2_X1 U8651 ( .A1(n6980), .A2(n6979), .ZN(n7066) );
  NAND2_X1 U8652 ( .A1(n7068), .A2(n7066), .ZN(n6986) );
  XNOR2_X1 U8653 ( .A(n9915), .B(n7375), .ZN(n6984) );
  INV_X1 U8654 ( .A(n6984), .ZN(n6982) );
  AND2_X1 U8655 ( .A1(n8437), .A2(n6682), .ZN(n6983) );
  INV_X1 U8656 ( .A(n6983), .ZN(n6981) );
  NAND2_X1 U8657 ( .A1(n6982), .A2(n6981), .ZN(n7069) );
  AND2_X1 U8658 ( .A1(n6984), .A2(n6983), .ZN(n7064) );
  NOR2_X1 U8659 ( .A1(n4806), .A2(n7064), .ZN(n6985) );
  XNOR2_X1 U8660 ( .A(n6986), .B(n6985), .ZN(n6991) );
  AOI22_X1 U8661 ( .A1(n7680), .A2(n8438), .B1(n8375), .B2(n7188), .ZN(n6988)
         );
  OAI211_X1 U8662 ( .C1(n7232), .C2(n8403), .A(n6988), .B(n6987), .ZN(n6989)
         );
  AOI21_X1 U8663 ( .B1(n7189), .B2(n8420), .A(n6989), .ZN(n6990) );
  OAI21_X1 U8664 ( .B1(n6991), .B2(n8422), .A(n6990), .ZN(P2_U3233) );
  INV_X1 U8665 ( .A(n6992), .ZN(n6994) );
  OAI222_X1 U8666 ( .A1(n7688), .A2(n6993), .B1(n9391), .B2(n6994), .C1(
        P1_U3084), .C2(n4299), .ZN(P1_U3331) );
  OAI222_X1 U8667 ( .A1(n7714), .A2(n6995), .B1(n8844), .B2(n6994), .C1(n7833), 
        .C2(P2_U3152), .ZN(P2_U3336) );
  NAND2_X1 U8668 ( .A1(n7004), .A2(n6996), .ZN(n6998) );
  NAND2_X1 U8669 ( .A1(n6998), .A2(n6997), .ZN(n7000) );
  XNOR2_X1 U8670 ( .A(n7008), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n6999) );
  NOR2_X1 U8671 ( .A1(n7000), .A2(n6999), .ZN(n7569) );
  AOI21_X1 U8672 ( .B1(n7000), .B2(n6999), .A(n7569), .ZN(n7014) );
  NOR2_X1 U8673 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7558), .ZN(n7002) );
  NOR2_X1 U8674 ( .A1(n9734), .A2(n7571), .ZN(n7001) );
  AOI211_X1 U8675 ( .C1(n9781), .C2(P2_ADDR_REG_16__SCAN_IN), .A(n7002), .B(
        n7001), .ZN(n7013) );
  NOR2_X1 U8676 ( .A1(n7004), .A2(n7003), .ZN(n7006) );
  NOR2_X1 U8677 ( .A1(n7006), .A2(n7005), .ZN(n7011) );
  NAND2_X1 U8678 ( .A1(n7008), .A2(n7566), .ZN(n7007) );
  OAI21_X1 U8679 ( .B1(n7008), .B2(n7566), .A(n7007), .ZN(n7010) );
  NAND2_X1 U8680 ( .A1(n7571), .A2(n7566), .ZN(n7009) );
  OAI211_X1 U8681 ( .C1(n7566), .C2(n7571), .A(n7011), .B(n7009), .ZN(n7565)
         );
  OAI211_X1 U8682 ( .C1(n7011), .C2(n7010), .A(n7565), .B(n9783), .ZN(n7012)
         );
  OAI211_X1 U8683 ( .C1(n7014), .C2(n9735), .A(n7013), .B(n7012), .ZN(P2_U3261) );
  OAI21_X1 U8684 ( .B1(n7017), .B2(n7016), .A(n7026), .ZN(n7018) );
  NAND2_X1 U8685 ( .A1(n7018), .A2(n8901), .ZN(n7024) );
  INV_X1 U8686 ( .A(n7019), .ZN(n7255) );
  NAND2_X1 U8687 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n9521) );
  INV_X1 U8688 ( .A(n9521), .ZN(n7020) );
  AOI21_X1 U8689 ( .B1(n8938), .B2(n9668), .A(n7020), .ZN(n7021) );
  OAI21_X1 U8690 ( .B1(n8936), .B2(n7166), .A(n7021), .ZN(n7022) );
  AOI21_X1 U8691 ( .B1(n7255), .B2(n8907), .A(n7022), .ZN(n7023) );
  OAI211_X1 U8692 ( .C1(n7257), .C2(n8910), .A(n7024), .B(n7023), .ZN(P1_U3225) );
  NAND2_X1 U8693 ( .A1(n7026), .A2(n7025), .ZN(n7029) );
  NAND2_X1 U8694 ( .A1(n4324), .A2(n7027), .ZN(n7028) );
  XNOR2_X1 U8695 ( .A(n7029), .B(n7028), .ZN(n7036) );
  INV_X1 U8696 ( .A(n7030), .ZN(n7032) );
  NOR2_X1 U8697 ( .A1(n8905), .A2(n7148), .ZN(n7031) );
  AOI211_X1 U8698 ( .C1(n8922), .C2(n8955), .A(n7032), .B(n7031), .ZN(n7033)
         );
  OAI21_X1 U8699 ( .B1(n8940), .B2(n7313), .A(n7033), .ZN(n7034) );
  AOI21_X1 U8700 ( .B1(n8942), .B2(n9694), .A(n7034), .ZN(n7035) );
  OAI21_X1 U8701 ( .B1(n7036), .B2(n8944), .A(n7035), .ZN(P1_U3237) );
  INV_X1 U8702 ( .A(n7200), .ZN(n7039) );
  OAI211_X1 U8703 ( .C1(n8204), .C2(n8109), .A(n7039), .B(n9626), .ZN(n9656)
         );
  NOR2_X1 U8704 ( .A1(n9656), .A2(n9127), .ZN(n7053) );
  INV_X1 U8705 ( .A(n8114), .ZN(n7046) );
  NAND2_X1 U8706 ( .A1(n6638), .A2(n9640), .ZN(n7137) );
  XNOR2_X1 U8707 ( .A(n7046), .B(n7137), .ZN(n9657) );
  OR2_X1 U8708 ( .A1(n7042), .A2(n7041), .ZN(n7045) );
  OR2_X1 U8709 ( .A1(n7043), .A2(n8197), .ZN(n7044) );
  NOR2_X1 U8710 ( .A1(n8098), .A2(n5718), .ZN(n9226) );
  AOI22_X1 U8711 ( .A1(n9226), .A2(n6638), .B1(n8957), .B2(n9686), .ZN(n7052)
         );
  NAND2_X1 U8712 ( .A1(n7046), .A2(n8110), .ZN(n7157) );
  OAI21_X1 U8713 ( .B1(n7046), .B2(n8110), .A(n7157), .ZN(n7050) );
  OR2_X1 U8714 ( .A1(n4299), .A2(n8985), .ZN(n7049) );
  NAND2_X1 U8715 ( .A1(n8206), .A2(n7047), .ZN(n7048) );
  NAND2_X1 U8716 ( .A1(n7049), .A2(n7048), .ZN(n9227) );
  NAND2_X1 U8717 ( .A1(n7050), .A2(n9227), .ZN(n7051) );
  OAI211_X1 U8718 ( .C1(n9657), .C2(n9610), .A(n7052), .B(n7051), .ZN(n9659)
         );
  AOI211_X1 U8719 ( .C1(n9646), .C2(P1_REG3_REG_1__SCAN_IN), .A(n7053), .B(
        n9659), .ZN(n7058) );
  NAND2_X1 U8720 ( .A1(n7055), .A2(n7054), .ZN(n7057) );
  NAND2_X2 U8721 ( .A1(n9206), .A2(n7170), .ZN(n9219) );
  MUX2_X1 U8722 ( .A(n6292), .B(n7058), .S(n9219), .Z(n7063) );
  INV_X1 U8723 ( .A(n9657), .ZN(n7061) );
  AND2_X1 U8724 ( .A1(n8206), .A2(n8242), .ZN(n7059) );
  NAND2_X1 U8725 ( .A1(n9219), .A2(n7059), .ZN(n7730) );
  INV_X1 U8726 ( .A(n7730), .ZN(n9630) );
  OR2_X1 U8727 ( .A1(n9633), .A2(n8201), .ZN(n7060) );
  NOR2_X2 U8728 ( .A1(n9620), .A2(n7060), .ZN(n9622) );
  AOI22_X1 U8729 ( .A1(n7061), .A2(n9630), .B1(n9622), .B2(n7038), .ZN(n7062)
         );
  NAND2_X1 U8730 ( .A1(n7063), .A2(n7062), .ZN(P1_U3290) );
  INV_X1 U8731 ( .A(n7064), .ZN(n7065) );
  AND2_X1 U8732 ( .A1(n7066), .A2(n7065), .ZN(n7067) );
  NAND2_X1 U8733 ( .A1(n7068), .A2(n7067), .ZN(n7070) );
  XNOR2_X1 U8734 ( .A(n9823), .B(n4296), .ZN(n7071) );
  NOR2_X1 U8735 ( .A1(n7232), .A2(n7321), .ZN(n7072) );
  NAND2_X1 U8736 ( .A1(n7071), .A2(n7072), .ZN(n7353) );
  INV_X1 U8737 ( .A(n7071), .ZN(n7074) );
  INV_X1 U8738 ( .A(n7072), .ZN(n7073) );
  NAND2_X1 U8739 ( .A1(n7074), .A2(n7073), .ZN(n7075) );
  NAND2_X1 U8740 ( .A1(n7353), .A2(n7075), .ZN(n7077) );
  AOI21_X1 U8741 ( .B1(n7076), .B2(n7077), .A(n8422), .ZN(n7078) );
  NAND2_X1 U8742 ( .A1(n7078), .A2(n7364), .ZN(n7082) );
  AND2_X1 U8743 ( .A1(n8437), .A2(n8545), .ZN(n7079) );
  AOI21_X1 U8744 ( .B1(n8436), .B2(n8547), .A(n7079), .ZN(n9820) );
  NAND2_X1 U8745 ( .A1(P2_U3152), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n9768) );
  OAI21_X1 U8746 ( .B1(n8417), .B2(n9820), .A(n9768), .ZN(n7080) );
  AOI21_X1 U8747 ( .B1(n9822), .B2(n8375), .A(n7080), .ZN(n7081) );
  OAI211_X1 U8748 ( .C1(n9923), .C2(n8360), .A(n7082), .B(n7081), .ZN(P2_U3219) );
  NAND2_X1 U8749 ( .A1(n7085), .A2(n7706), .ZN(n8968) );
  OAI21_X1 U8750 ( .B1(n7085), .B2(n7706), .A(n8968), .ZN(n7095) );
  AOI21_X1 U8751 ( .B1(n9340), .B2(n7087), .A(n7086), .ZN(n7090) );
  AOI22_X1 U8752 ( .A1(n7088), .A2(n6001), .B1(P1_REG1_REG_14__SCAN_IN), .B2(
        n8966), .ZN(n7089) );
  NOR2_X1 U8753 ( .A1(n7090), .A2(n7089), .ZN(n8958) );
  AOI21_X1 U8754 ( .B1(n7090), .B2(n7089), .A(n8958), .ZN(n7091) );
  OR2_X1 U8755 ( .A1(n7091), .A2(n9605), .ZN(n7093) );
  NOR2_X1 U8756 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n10161), .ZN(n7618) );
  AOI21_X1 U8757 ( .B1(n9535), .B2(P1_ADDR_REG_14__SCAN_IN), .A(n7618), .ZN(
        n7092) );
  OAI211_X1 U8758 ( .C1(n9599), .C2(n8966), .A(n7093), .B(n7092), .ZN(n7094)
         );
  AOI21_X1 U8759 ( .B1(n9595), .B2(n7095), .A(n7094), .ZN(n7096) );
  INV_X1 U8760 ( .A(n7096), .ZN(P1_U3255) );
  INV_X1 U8761 ( .A(n7097), .ZN(n7101) );
  NOR2_X1 U8762 ( .A1(n7098), .A2(P1_U3084), .ZN(n8247) );
  AOI21_X1 U8763 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(n9389), .A(n8247), .ZN(
        n7099) );
  OAI21_X1 U8764 ( .B1(n7101), .B2(n9391), .A(n7099), .ZN(P1_U3330) );
  NAND2_X1 U8765 ( .A1(n8841), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n7100) );
  OAI211_X1 U8766 ( .C1(n7101), .C2(n8844), .A(n7100), .B(n8005), .ZN(P2_U3335) );
  AOI22_X1 U8767 ( .A1(n9834), .A2(n7103), .B1(n9856), .B2(n7102), .ZN(n7106)
         );
  INV_X1 U8768 ( .A(n9832), .ZN(n9862) );
  AOI22_X1 U8769 ( .A1(n7104), .A2(n9862), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n9854), .ZN(n7105) );
  OAI211_X1 U8770 ( .C1(n7107), .C2(n8579), .A(n7106), .B(n7105), .ZN(n7108)
         );
  AOI21_X1 U8771 ( .B1(n8579), .B2(n7109), .A(n7108), .ZN(n7110) );
  INV_X1 U8772 ( .A(n7110), .ZN(P2_U3295) );
  XOR2_X1 U8773 ( .A(n7112), .B(n7111), .Z(n7113) );
  XNOR2_X1 U8774 ( .A(n7114), .B(n7113), .ZN(n7122) );
  INV_X1 U8775 ( .A(n7174), .ZN(n7269) );
  NOR2_X1 U8776 ( .A1(n7269), .A2(n9678), .ZN(n9702) );
  NAND2_X1 U8777 ( .A1(n8938), .A2(n9687), .ZN(n7119) );
  NAND2_X1 U8778 ( .A1(n8922), .A2(n8954), .ZN(n7118) );
  INV_X1 U8779 ( .A(n7115), .ZN(n7171) );
  NAND2_X1 U8780 ( .A1(n8907), .A2(n7171), .ZN(n7116) );
  NAND4_X1 U8781 ( .A1(n7119), .A2(n7118), .A3(n7117), .A4(n7116), .ZN(n7120)
         );
  AOI21_X1 U8782 ( .B1(n7241), .B2(n9702), .A(n7120), .ZN(n7121) );
  OAI21_X1 U8783 ( .B1(n7122), .B2(n8944), .A(n7121), .ZN(P1_U3211) );
  XNOR2_X1 U8784 ( .A(n7123), .B(n7869), .ZN(n9907) );
  INV_X1 U8785 ( .A(n7124), .ZN(n7776) );
  OAI211_X1 U8786 ( .C1(n7776), .C2(n9904), .A(n7321), .B(n9858), .ZN(n9903)
         );
  AOI22_X1 U8787 ( .A1(n9856), .A2(n7126), .B1(n9854), .B2(n7125), .ZN(n7127)
         );
  OAI21_X1 U8788 ( .B1(n9903), .B2(n9832), .A(n7127), .ZN(n7135) );
  INV_X1 U8789 ( .A(n7868), .ZN(n7128) );
  NAND2_X1 U8790 ( .A1(n7782), .A2(n7128), .ZN(n7129) );
  NAND2_X1 U8791 ( .A1(n7129), .A2(n7869), .ZN(n7131) );
  NAND3_X1 U8792 ( .A1(n7131), .A2(n9818), .A3(n7130), .ZN(n7133) );
  AOI22_X1 U8793 ( .A1(n8545), .A2(n8440), .B1(n8438), .B2(n8547), .ZN(n7132)
         );
  NAND2_X1 U8794 ( .A1(n7133), .A2(n7132), .ZN(n9905) );
  MUX2_X1 U8795 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n9905), .S(n8579), .Z(n7134)
         );
  AOI211_X1 U8796 ( .C1(n9834), .C2(n9907), .A(n7135), .B(n7134), .ZN(n7136)
         );
  INV_X1 U8797 ( .A(n7136), .ZN(P2_U3289) );
  NAND2_X1 U8798 ( .A1(n7155), .A2(n8204), .ZN(n7138) );
  NAND2_X1 U8799 ( .A1(n7139), .A2(n7138), .ZN(n7195) );
  NAND2_X1 U8800 ( .A1(n8957), .A2(n7199), .ZN(n8210) );
  NAND2_X1 U8801 ( .A1(n7280), .A2(n7199), .ZN(n7140) );
  NAND2_X1 U8802 ( .A1(n7141), .A2(n7140), .ZN(n7279) );
  NAND2_X1 U8803 ( .A1(n6792), .A2(n7285), .ZN(n8209) );
  NAND2_X1 U8804 ( .A1(n7279), .A2(n8108), .ZN(n7144) );
  NAND2_X1 U8805 ( .A1(n7142), .A2(n7285), .ZN(n7143) );
  NAND2_X1 U8806 ( .A1(n7144), .A2(n7143), .ZN(n9611) );
  NAND2_X1 U8807 ( .A1(n7145), .A2(n9623), .ZN(n7250) );
  NAND2_X1 U8808 ( .A1(n9668), .A2(n9679), .ZN(n8215) );
  NAND2_X1 U8809 ( .A1(n7250), .A2(n8215), .ZN(n9612) );
  NAND2_X1 U8810 ( .A1(n9611), .A2(n9612), .ZN(n7147) );
  NAND2_X1 U8811 ( .A1(n7145), .A2(n9679), .ZN(n7146) );
  NAND2_X1 U8812 ( .A1(n7147), .A2(n7146), .ZN(n7261) );
  INV_X1 U8813 ( .A(n7261), .ZN(n7150) );
  NAND2_X1 U8814 ( .A1(n7148), .A2(n9685), .ZN(n8155) );
  NAND2_X1 U8815 ( .A1(n9614), .A2(n7257), .ZN(n8012) );
  NAND2_X1 U8816 ( .A1(n7150), .A2(n7149), .ZN(n7260) );
  NAND2_X1 U8817 ( .A1(n9614), .A2(n9685), .ZN(n7151) );
  NAND2_X1 U8818 ( .A1(n7260), .A2(n7151), .ZN(n7306) );
  NAND2_X1 U8819 ( .A1(n7166), .A2(n9694), .ZN(n8156) );
  INV_X1 U8820 ( .A(n9694), .ZN(n7314) );
  NAND2_X1 U8821 ( .A1(n9687), .A2(n7314), .ZN(n8016) );
  NAND2_X1 U8822 ( .A1(n7166), .A2(n7314), .ZN(n7152) );
  NAND2_X1 U8823 ( .A1(n7294), .A2(n7174), .ZN(n8148) );
  NAND2_X1 U8824 ( .A1(n8955), .A2(n7269), .ZN(n8024) );
  NAND2_X1 U8825 ( .A1(n8148), .A2(n8024), .ZN(n8116) );
  XNOR2_X1 U8826 ( .A(n7268), .B(n8116), .ZN(n9709) );
  INV_X1 U8827 ( .A(n9709), .ZN(n7178) );
  AND2_X1 U8828 ( .A1(n9634), .A2(n4298), .ZN(n7154) );
  NAND2_X1 U8829 ( .A1(n9219), .A2(n7154), .ZN(n9222) );
  NAND2_X1 U8830 ( .A1(n7155), .A2(n7038), .ZN(n7156) );
  NAND2_X1 U8831 ( .A1(n7157), .A2(n7156), .ZN(n8212) );
  NAND2_X1 U8832 ( .A1(n8212), .A2(n8111), .ZN(n7197) );
  NAND2_X1 U8833 ( .A1(n9613), .A2(n8215), .ZN(n8009) );
  AND3_X1 U8834 ( .A1(n8156), .A2(n8155), .A3(n7250), .ZN(n8219) );
  NAND2_X1 U8835 ( .A1(n8009), .A2(n8219), .ZN(n7161) );
  INV_X1 U8836 ( .A(n8012), .ZN(n7159) );
  NAND2_X1 U8837 ( .A1(n8156), .A2(n7159), .ZN(n8153) );
  AND2_X1 U8838 ( .A1(n8153), .A2(n8016), .ZN(n7160) );
  NAND2_X1 U8839 ( .A1(n7161), .A2(n7160), .ZN(n7165) );
  INV_X1 U8840 ( .A(n7264), .ZN(n7164) );
  AOI21_X1 U8841 ( .B1(n8116), .B2(n7165), .A(n7164), .ZN(n7167) );
  INV_X1 U8842 ( .A(n9227), .ZN(n9617) );
  INV_X1 U8843 ( .A(n9226), .ZN(n9217) );
  OAI22_X1 U8844 ( .A1(n7167), .A2(n9617), .B1(n7166), .B2(n9217), .ZN(n9707)
         );
  INV_X1 U8845 ( .A(n7168), .ZN(n7311) );
  INV_X1 U8846 ( .A(n7169), .ZN(n7298) );
  OAI211_X1 U8847 ( .C1(n7269), .C2(n7311), .A(n7298), .B(n9626), .ZN(n9704)
         );
  NOR2_X2 U8848 ( .A1(n7170), .A2(n9127), .ZN(n9629) );
  NAND2_X1 U8849 ( .A1(n9219), .A2(n9686), .ZN(n9235) );
  INV_X1 U8850 ( .A(n8954), .ZN(n9706) );
  AOI22_X1 U8851 ( .A1(n9620), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n7171), .B2(
        n9646), .ZN(n7172) );
  OAI21_X1 U8852 ( .B1(n9235), .B2(n9706), .A(n7172), .ZN(n7173) );
  AOI21_X1 U8853 ( .B1(n9622), .B2(n7174), .A(n7173), .ZN(n7175) );
  OAI21_X1 U8854 ( .B1(n9704), .B2(n9239), .A(n7175), .ZN(n7176) );
  AOI21_X1 U8855 ( .B1(n9707), .B2(n9219), .A(n7176), .ZN(n7177) );
  OAI21_X1 U8856 ( .B1(n7178), .B2(n9222), .A(n7177), .ZN(P1_U3284) );
  OR2_X1 U8857 ( .A1(n7179), .A2(n7811), .ZN(n9825) );
  INV_X1 U8858 ( .A(n9825), .ZN(n7180) );
  AOI21_X1 U8859 ( .B1(n7811), .B2(n7179), .A(n7180), .ZN(n7185) );
  XNOR2_X1 U8860 ( .A(n7181), .B(n7811), .ZN(n7183) );
  OAI22_X1 U8861 ( .A1(n7876), .A2(n9846), .B1(n7232), .B2(n9848), .ZN(n7182)
         );
  AOI21_X1 U8862 ( .B1(n7183), .B2(n9818), .A(n7182), .ZN(n7184) );
  OAI21_X1 U8863 ( .B1(n7185), .B2(n8679), .A(n7184), .ZN(n9917) );
  INV_X1 U8864 ( .A(n9917), .ZN(n7194) );
  INV_X1 U8865 ( .A(n7185), .ZN(n9919) );
  NOR2_X1 U8866 ( .A1(n9866), .A2(n7186), .ZN(n9863) );
  NOR2_X1 U8867 ( .A1(n9859), .A2(n9915), .ZN(n7187) );
  OR2_X1 U8868 ( .A1(n9831), .A2(n7187), .ZN(n9916) );
  AOI22_X1 U8869 ( .A1(n9866), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n7188), .B2(
        n9854), .ZN(n7191) );
  NAND2_X1 U8870 ( .A1(n9856), .A2(n7189), .ZN(n7190) );
  OAI211_X1 U8871 ( .C1(n9916), .C2(n7798), .A(n7191), .B(n7190), .ZN(n7192)
         );
  AOI21_X1 U8872 ( .B1(n9919), .B2(n9863), .A(n7192), .ZN(n7193) );
  OAI21_X1 U8873 ( .B1(n7194), .B2(n9855), .A(n7193), .ZN(P2_U3287) );
  XNOR2_X1 U8874 ( .A(n7195), .B(n7196), .ZN(n9666) );
  INV_X1 U8875 ( .A(n9666), .ZN(n7207) );
  OAI21_X1 U8876 ( .B1(n8111), .B2(n8212), .A(n7197), .ZN(n7198) );
  AOI22_X1 U8877 ( .A1(n7198), .A2(n9227), .B1(n9615), .B2(n7040), .ZN(n9664)
         );
  INV_X1 U8878 ( .A(n9664), .ZN(n7205) );
  OAI211_X1 U8879 ( .C1(n7200), .C2(n7199), .A(n9626), .B(n7282), .ZN(n9661)
         );
  NOR2_X1 U8880 ( .A1(n9661), .A2(n9239), .ZN(n7204) );
  NAND2_X1 U8881 ( .A1(n9622), .A2(n9660), .ZN(n7202) );
  AOI22_X1 U8882 ( .A1(n9620), .A2(P1_REG2_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n9646), .ZN(n7201) );
  OAI211_X1 U8883 ( .C1(n9235), .C2(n7142), .A(n7202), .B(n7201), .ZN(n7203)
         );
  AOI211_X1 U8884 ( .C1(n7205), .C2(n9219), .A(n7204), .B(n7203), .ZN(n7206)
         );
  OAI21_X1 U8885 ( .B1(n9222), .B2(n7207), .A(n7206), .ZN(P1_U3289) );
  MUX2_X1 U8886 ( .A(n6388), .B(n7208), .S(n8579), .Z(n7216) );
  NOR2_X1 U8887 ( .A1(n9866), .A2(n8539), .ZN(n8641) );
  INV_X1 U8888 ( .A(n7209), .ZN(n7214) );
  INV_X1 U8889 ( .A(n7210), .ZN(n7211) );
  OAI22_X1 U8890 ( .A1(n8693), .A2(n7212), .B1(n8556), .B2(n7211), .ZN(n7213)
         );
  AOI21_X1 U8891 ( .B1(n8641), .B2(n7214), .A(n7213), .ZN(n7215) );
  OAI211_X1 U8892 ( .C1(n7217), .C2(n8709), .A(n7216), .B(n7215), .ZN(P2_U3291) );
  INV_X1 U8893 ( .A(n7218), .ZN(n7221) );
  OAI222_X1 U8894 ( .A1(P2_U3152), .A2(n9870), .B1(n8844), .B2(n7221), .C1(
        n7219), .C2(n7714), .ZN(P2_U3334) );
  OAI222_X1 U8895 ( .A1(n7222), .A2(P1_U3084), .B1(n9391), .B2(n7221), .C1(
        n7220), .C2(n7688), .ZN(P1_U3329) );
  AOI22_X1 U8896 ( .A1(n9862), .A2(n7223), .B1(n9854), .B2(n5056), .ZN(n7224)
         );
  OAI21_X1 U8897 ( .B1(n8693), .B2(n7225), .A(n7224), .ZN(n7228) );
  MUX2_X1 U8898 ( .A(n7226), .B(P2_REG2_REG_3__SCAN_IN), .S(n9866), .Z(n7227)
         );
  AOI211_X1 U8899 ( .C1(n9863), .C2(n7229), .A(n7228), .B(n7227), .ZN(n7230)
         );
  INV_X1 U8900 ( .A(n7230), .ZN(P2_U3293) );
  NAND2_X1 U8901 ( .A1(n7364), .A2(n7353), .ZN(n7231) );
  XNOR2_X1 U8902 ( .A(n9926), .B(n4296), .ZN(n7320) );
  NAND2_X1 U8903 ( .A1(n8436), .A2(n6682), .ZN(n7318) );
  XNOR2_X1 U8904 ( .A(n7320), .B(n7318), .ZN(n7360) );
  NAND2_X1 U8905 ( .A1(n7231), .A2(n7360), .ZN(n7336) );
  OAI211_X1 U8906 ( .C1(n7231), .C2(n7360), .A(n7336), .B(n8352), .ZN(n7236)
         );
  NOR2_X1 U8907 ( .A1(n8404), .A2(n7232), .ZN(n7234) );
  OAI22_X1 U8908 ( .A1(n8403), .A2(n7412), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5179), .ZN(n7233) );
  AOI211_X1 U8909 ( .C1(n8375), .C2(n7431), .A(n7234), .B(n7233), .ZN(n7235)
         );
  OAI211_X1 U8910 ( .C1(n4559), .C2(n8360), .A(n7236), .B(n7235), .ZN(P2_U3238) );
  XOR2_X1 U8911 ( .A(n7238), .B(n7237), .Z(n7239) );
  XNOR2_X1 U8912 ( .A(n7240), .B(n7239), .ZN(n7249) );
  NOR2_X1 U8913 ( .A1(n7302), .A2(n9678), .ZN(n9715) );
  NAND2_X1 U8914 ( .A1(n9715), .A2(n7241), .ZN(n7247) );
  NAND2_X1 U8915 ( .A1(P1_U3084), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n9533) );
  INV_X1 U8916 ( .A(n9533), .ZN(n7242) );
  AOI21_X1 U8917 ( .B1(n8922), .B2(n8953), .A(n7242), .ZN(n7246) );
  INV_X1 U8918 ( .A(n7243), .ZN(n7300) );
  NAND2_X1 U8919 ( .A1(n8907), .A2(n7300), .ZN(n7245) );
  NAND2_X1 U8920 ( .A1(n8938), .A2(n8955), .ZN(n7244) );
  AND4_X1 U8921 ( .A1(n7247), .A2(n7246), .A3(n7245), .A4(n7244), .ZN(n7248)
         );
  OAI21_X1 U8922 ( .B1(n7249), .B2(n8944), .A(n7248), .ZN(P1_U3219) );
  INV_X1 U8923 ( .A(n7250), .ZN(n7251) );
  INV_X1 U8924 ( .A(n8215), .ZN(n7252) );
  NOR2_X1 U8925 ( .A1(n8011), .A2(n7252), .ZN(n7253) );
  NAND2_X1 U8926 ( .A1(n7253), .A2(n8112), .ZN(n7307) );
  OAI21_X1 U8927 ( .B1(n8112), .B2(n7253), .A(n7307), .ZN(n7254) );
  AOI22_X1 U8928 ( .A1(n7254), .A2(n9227), .B1(n9226), .B2(n9668), .ZN(n9692)
         );
  INV_X1 U8929 ( .A(n9235), .ZN(n7454) );
  AOI22_X1 U8930 ( .A1(n9620), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n7255), .B2(
        n9646), .ZN(n7256) );
  OAI21_X1 U8931 ( .B1(n9204), .B2(n7257), .A(n7256), .ZN(n7259) );
  OAI211_X1 U8932 ( .C1(n9625), .C2(n7257), .A(n7312), .B(n9626), .ZN(n9689)
         );
  NOR2_X1 U8933 ( .A1(n9689), .A2(n9239), .ZN(n7258) );
  AOI211_X1 U8934 ( .C1(n7454), .C2(n9687), .A(n7259), .B(n7258), .ZN(n7263)
         );
  NAND2_X1 U8935 ( .A1(n7261), .A2(n8112), .ZN(n9688) );
  NAND3_X1 U8936 ( .A1(n7260), .A2(n9688), .A3(n9231), .ZN(n7262) );
  OAI211_X1 U8937 ( .C1(n9692), .C2(n9620), .A(n7263), .B(n7262), .ZN(P1_U3286) );
  NAND2_X1 U8938 ( .A1(n9706), .A2(n7299), .ZN(n8149) );
  NAND2_X1 U8939 ( .A1(n8954), .A2(n7302), .ZN(n8029) );
  NAND2_X1 U8940 ( .A1(n7265), .A2(n8029), .ZN(n7695) );
  INV_X1 U8941 ( .A(n8953), .ZN(n7494) );
  NAND2_X1 U8942 ( .A1(n7494), .A2(n7468), .ZN(n8036) );
  INV_X1 U8943 ( .A(n8036), .ZN(n7266) );
  AND2_X1 U8944 ( .A1(n7393), .A2(n8953), .ZN(n8039) );
  OR2_X1 U8945 ( .A1(n7266), .A2(n8039), .ZN(n8121) );
  XNOR2_X1 U8946 ( .A(n7695), .B(n8121), .ZN(n7267) );
  AOI22_X1 U8947 ( .A1(n7267), .A2(n9227), .B1(n9226), .B2(n8954), .ZN(n7388)
         );
  NAND2_X1 U8948 ( .A1(n7294), .A2(n7269), .ZN(n7270) );
  NAND2_X1 U8949 ( .A1(n8954), .A2(n7299), .ZN(n7271) );
  NAND2_X1 U8950 ( .A1(n7292), .A2(n7271), .ZN(n7450) );
  XOR2_X1 U8951 ( .A(n7450), .B(n8121), .Z(n7390) );
  NAND2_X1 U8952 ( .A1(n7390), .A2(n9231), .ZN(n7278) );
  INV_X1 U8953 ( .A(n7466), .ZN(n7272) );
  AOI22_X1 U8954 ( .A1(n9620), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n7272), .B2(
        n9646), .ZN(n7273) );
  OAI21_X1 U8955 ( .B1(n9235), .B2(n7444), .A(n7273), .ZN(n7276) );
  OAI211_X1 U8956 ( .C1(n7274), .C2(n7393), .A(n9626), .B(n7481), .ZN(n7387)
         );
  NOR2_X1 U8957 ( .A1(n7387), .A2(n9239), .ZN(n7275) );
  AOI211_X1 U8958 ( .C1(n9622), .C2(n7468), .A(n7276), .B(n7275), .ZN(n7277)
         );
  OAI211_X1 U8959 ( .C1(n9620), .C2(n7388), .A(n7278), .B(n7277), .ZN(P1_U3282) );
  XOR2_X1 U8960 ( .A(n7279), .B(n8108), .Z(n9671) );
  XNOR2_X1 U8961 ( .A(n8108), .B(n8154), .ZN(n7281) );
  OAI22_X1 U8962 ( .A1(n7281), .A2(n9617), .B1(n7280), .B2(n9217), .ZN(n9673)
         );
  NAND2_X1 U8963 ( .A1(n9673), .A2(n9219), .ZN(n7289) );
  AOI21_X1 U8964 ( .B1(n7282), .B2(n9667), .A(n9236), .ZN(n7283) );
  NAND2_X1 U8965 ( .A1(n7283), .A2(n9624), .ZN(n9669) );
  NOR2_X1 U8966 ( .A1(n9669), .A2(n9239), .ZN(n7287) );
  AOI22_X1 U8967 ( .A1(n9620), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n9646), .B2(
        n5816), .ZN(n7284) );
  OAI21_X1 U8968 ( .B1(n9204), .B2(n7285), .A(n7284), .ZN(n7286) );
  AOI211_X1 U8969 ( .C1(n7454), .C2(n9668), .A(n7287), .B(n7286), .ZN(n7288)
         );
  OAI211_X1 U8970 ( .C1(n9222), .C2(n9671), .A(n7289), .B(n7288), .ZN(P1_U3288) );
  NAND2_X1 U8971 ( .A1(n7290), .A2(n8118), .ZN(n7291) );
  NAND2_X1 U8972 ( .A1(n7292), .A2(n7291), .ZN(n9713) );
  XNOR2_X1 U8973 ( .A(n7293), .B(n8118), .ZN(n7296) );
  OAI22_X1 U8974 ( .A1(n7494), .A2(n9705), .B1(n7294), .B2(n9217), .ZN(n7295)
         );
  AOI21_X1 U8975 ( .B1(n7296), .B2(n9227), .A(n7295), .ZN(n7297) );
  OAI21_X1 U8976 ( .B1(n9713), .B2(n9610), .A(n7297), .ZN(n9717) );
  NAND2_X1 U8977 ( .A1(n9717), .A2(n9219), .ZN(n7305) );
  AOI211_X1 U8978 ( .C1(n7299), .C2(n7298), .A(n9236), .B(n7274), .ZN(n9714)
         );
  AOI22_X1 U8979 ( .A1(n9620), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n7300), .B2(
        n9646), .ZN(n7301) );
  OAI21_X1 U8980 ( .B1(n9204), .B2(n7302), .A(n7301), .ZN(n7303) );
  AOI21_X1 U8981 ( .B1(n9714), .B2(n9629), .A(n7303), .ZN(n7304) );
  OAI211_X1 U8982 ( .C1(n9713), .C2(n7730), .A(n7305), .B(n7304), .ZN(P1_U3283) );
  INV_X1 U8983 ( .A(n8117), .ZN(n8013) );
  XNOR2_X1 U8984 ( .A(n7306), .B(n8013), .ZN(n9698) );
  NAND2_X1 U8985 ( .A1(n7307), .A2(n8155), .ZN(n7308) );
  XNOR2_X1 U8986 ( .A(n7308), .B(n8117), .ZN(n7309) );
  AOI222_X1 U8987 ( .A1(n9227), .A2(n7309), .B1(n8955), .B2(n9686), .C1(n9614), 
        .C2(n9226), .ZN(n9697) );
  MUX2_X1 U8988 ( .A(n7310), .B(n9697), .S(n9219), .Z(n7317) );
  AOI211_X1 U8989 ( .C1(n9694), .C2(n7312), .A(n9236), .B(n7311), .ZN(n9693)
         );
  OAI22_X1 U8990 ( .A1(n9204), .A2(n7314), .B1(n7313), .B2(n9206), .ZN(n7315)
         );
  AOI21_X1 U8991 ( .B1(n9693), .B2(n9629), .A(n7315), .ZN(n7316) );
  OAI211_X1 U8992 ( .C1(n9222), .C2(n9698), .A(n7317), .B(n7316), .ZN(P1_U3285) );
  INV_X1 U8993 ( .A(n9809), .ZN(n9938) );
  INV_X1 U8994 ( .A(n7318), .ZN(n7319) );
  NAND2_X1 U8995 ( .A1(n7320), .A2(n7319), .ZN(n7335) );
  NAND2_X1 U8996 ( .A1(n7336), .A2(n7335), .ZN(n7327) );
  XNOR2_X1 U8997 ( .A(n9809), .B(n7375), .ZN(n7322) );
  OR2_X1 U8998 ( .A1(n7412), .A2(n7321), .ZN(n7323) );
  NAND2_X1 U8999 ( .A1(n7322), .A2(n7323), .ZN(n7349) );
  INV_X1 U9000 ( .A(n7322), .ZN(n7325) );
  INV_X1 U9001 ( .A(n7323), .ZN(n7324) );
  NAND2_X1 U9002 ( .A1(n7325), .A2(n7324), .ZN(n7334) );
  NAND2_X1 U9003 ( .A1(n7349), .A2(n7334), .ZN(n7326) );
  XNOR2_X1 U9004 ( .A(n7327), .B(n7326), .ZN(n7328) );
  NAND2_X1 U9005 ( .A1(n7328), .A2(n8352), .ZN(n7333) );
  NAND2_X1 U9006 ( .A1(n8436), .A2(n8545), .ZN(n7330) );
  NAND2_X1 U9007 ( .A1(n8434), .A2(n8547), .ZN(n7329) );
  AND2_X1 U9008 ( .A1(n7330), .A2(n7329), .ZN(n9802) );
  OAI22_X1 U9009 ( .A1(n8417), .A2(n9802), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10078), .ZN(n7331) );
  AOI21_X1 U9010 ( .B1(n9804), .B2(n8375), .A(n7331), .ZN(n7332) );
  OAI211_X1 U9011 ( .C1(n9938), .C2(n8360), .A(n7333), .B(n7332), .ZN(P2_U3226) );
  AND2_X1 U9012 ( .A1(n7335), .A2(n7334), .ZN(n7351) );
  NAND2_X1 U9013 ( .A1(n7336), .A2(n7351), .ZN(n7337) );
  AND2_X1 U9014 ( .A1(n7337), .A2(n7349), .ZN(n7338) );
  XNOR2_X1 U9015 ( .A(n8796), .B(n4296), .ZN(n7356) );
  NAND2_X1 U9016 ( .A1(n8434), .A2(n6682), .ZN(n7354) );
  XNOR2_X1 U9017 ( .A(n7356), .B(n7354), .ZN(n7350) );
  XNOR2_X1 U9018 ( .A(n7338), .B(n7350), .ZN(n7343) );
  OAI22_X1 U9019 ( .A1(n8403), .A2(n7411), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5213), .ZN(n7341) );
  INV_X1 U9020 ( .A(n7419), .ZN(n7339) );
  OAI22_X1 U9021 ( .A1(n8404), .A2(n7412), .B1(n8411), .B2(n7339), .ZN(n7340)
         );
  AOI211_X1 U9022 ( .C1(n8796), .C2(n8420), .A(n7341), .B(n7340), .ZN(n7342)
         );
  OAI21_X1 U9023 ( .B1(n7343), .B2(n8422), .A(n7342), .ZN(P2_U3236) );
  XNOR2_X1 U9024 ( .A(n8791), .B(n7375), .ZN(n7344) );
  NAND2_X1 U9025 ( .A1(n8433), .A2(n6682), .ZN(n7345) );
  NAND2_X1 U9026 ( .A1(n7344), .A2(n7345), .ZN(n7373) );
  INV_X1 U9027 ( .A(n7344), .ZN(n7347) );
  INV_X1 U9028 ( .A(n7345), .ZN(n7346) );
  NAND2_X1 U9029 ( .A1(n7347), .A2(n7346), .ZN(n7348) );
  NAND2_X1 U9030 ( .A1(n7373), .A2(n7348), .ZN(n7367) );
  AND2_X1 U9031 ( .A1(n7353), .A2(n7358), .ZN(n7357) );
  INV_X1 U9032 ( .A(n7354), .ZN(n7355) );
  NAND2_X1 U9033 ( .A1(n7356), .A2(n7355), .ZN(n7362) );
  AND2_X1 U9034 ( .A1(n7357), .A2(n7362), .ZN(n7363) );
  AND2_X1 U9035 ( .A1(n7360), .A2(n7359), .ZN(n7361) );
  OR2_X2 U9036 ( .A1(n7365), .A2(n7367), .ZN(n7374) );
  INV_X1 U9037 ( .A(n7374), .ZN(n7366) );
  AOI21_X1 U9038 ( .B1(n7367), .B2(n7365), .A(n7366), .ZN(n7372) );
  OAI22_X1 U9039 ( .A1(n8403), .A2(n7607), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10091), .ZN(n7370) );
  INV_X1 U9040 ( .A(n7602), .ZN(n7368) );
  OAI22_X1 U9041 ( .A1(n8404), .A2(n7606), .B1(n8411), .B2(n7368), .ZN(n7369)
         );
  AOI211_X1 U9042 ( .C1(n8791), .C2(n8420), .A(n7370), .B(n7369), .ZN(n7371)
         );
  OAI21_X1 U9043 ( .B1(n7372), .B2(n8422), .A(n7371), .ZN(P2_U3217) );
  NAND2_X2 U9044 ( .A1(n7374), .A2(n7373), .ZN(n7552) );
  XNOR2_X1 U9045 ( .A(n8786), .B(n7375), .ZN(n7551) );
  NAND2_X1 U9046 ( .A1(n8432), .A2(n6682), .ZN(n7550) );
  XNOR2_X1 U9047 ( .A(n7551), .B(n7550), .ZN(n7376) );
  XNOR2_X1 U9048 ( .A(n7552), .B(n7376), .ZN(n7383) );
  INV_X1 U9049 ( .A(n8691), .ZN(n7380) );
  NOR2_X1 U9050 ( .A1(n7411), .A2(n9846), .ZN(n7378) );
  NOR2_X1 U9051 ( .A1(n8674), .A2(n9848), .ZN(n7377) );
  OR2_X1 U9052 ( .A1(n7378), .A2(n7377), .ZN(n8702) );
  AOI22_X1 U9053 ( .A1(n8364), .A2(n8702), .B1(P2_REG3_REG_15__SCAN_IN), .B2(
        P2_U3152), .ZN(n7379) );
  OAI21_X1 U9054 ( .B1(n7380), .B2(n8411), .A(n7379), .ZN(n7381) );
  AOI21_X1 U9055 ( .B1(n8786), .B2(n8420), .A(n7381), .ZN(n7382) );
  OAI21_X1 U9056 ( .B1(n7383), .B2(n8422), .A(n7382), .ZN(P2_U3243) );
  INV_X1 U9057 ( .A(n7384), .ZN(n7443) );
  AOI22_X1 U9058 ( .A1(n7385), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n9389), .ZN(n7386) );
  OAI21_X1 U9059 ( .B1(n7443), .B2(n9391), .A(n7386), .ZN(P1_U3327) );
  NAND2_X1 U9060 ( .A1(n4299), .A2(n8242), .ZN(n9712) );
  OAI211_X1 U9061 ( .C1(n7444), .C2(n9705), .A(n7388), .B(n7387), .ZN(n7389)
         );
  AOI21_X1 U9062 ( .B1(n7390), .B2(n9710), .A(n7389), .ZN(n7396) );
  OAI22_X1 U9063 ( .A1(n9342), .A2(n7393), .B1(n9733), .B2(n5912), .ZN(n7391)
         );
  INV_X1 U9064 ( .A(n7391), .ZN(n7392) );
  OAI21_X1 U9065 ( .B1(n7396), .B2(n9731), .A(n7392), .ZN(P1_U3532) );
  OAI22_X1 U9066 ( .A1(n9379), .A2(n7393), .B1(n9720), .B2(n5913), .ZN(n7394)
         );
  INV_X1 U9067 ( .A(n7394), .ZN(n7395) );
  OAI21_X1 U9068 ( .B1(n7396), .B2(n9718), .A(n7395), .ZN(P1_U3481) );
  INV_X1 U9069 ( .A(n7397), .ZN(n7401) );
  OAI222_X1 U9070 ( .A1(n7688), .A2(n10121), .B1(n7399), .B2(n7401), .C1(n7398), .C2(P1_U3084), .ZN(P1_U3328) );
  OAI222_X1 U9071 ( .A1(n7714), .A2(n7402), .B1(n8844), .B2(n7401), .C1(
        P2_U3152), .C2(n7400), .ZN(P2_U3333) );
  OR2_X1 U9072 ( .A1(n7179), .A2(n7403), .ZN(n7405) );
  AND2_X1 U9073 ( .A1(n7405), .A2(n7404), .ZN(n9805) );
  OR2_X1 U9074 ( .A1(n9805), .A2(n9800), .ZN(n9806) );
  AND2_X1 U9075 ( .A1(n9806), .A2(n7406), .ZN(n7408) );
  OAI21_X1 U9076 ( .B1(n7408), .B2(n7892), .A(n7407), .ZN(n7417) );
  OR2_X1 U9077 ( .A1(n7417), .A2(n8679), .ZN(n7416) );
  OAI21_X1 U9078 ( .B1(n7817), .B2(n7410), .A(n7409), .ZN(n7414) );
  OAI22_X1 U9079 ( .A1(n7412), .A2(n9846), .B1(n7411), .B2(n9848), .ZN(n7413)
         );
  AOI21_X1 U9080 ( .B1(n7414), .B2(n9818), .A(n7413), .ZN(n7415) );
  AND2_X1 U9081 ( .A1(n7416), .A2(n7415), .ZN(n8802) );
  INV_X1 U9082 ( .A(n7417), .ZN(n8800) );
  AND2_X1 U9083 ( .A1(n9811), .A2(n8796), .ZN(n7418) );
  OR2_X1 U9084 ( .A1(n7418), .A2(n7599), .ZN(n8798) );
  AOI22_X1 U9085 ( .A1(n9866), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n7419), .B2(
        n9854), .ZN(n7421) );
  NAND2_X1 U9086 ( .A1(n8796), .A2(n9856), .ZN(n7420) );
  OAI211_X1 U9087 ( .C1(n8798), .C2(n7798), .A(n7421), .B(n7420), .ZN(n7422)
         );
  AOI21_X1 U9088 ( .B1(n8800), .B2(n9863), .A(n7422), .ZN(n7423) );
  OAI21_X1 U9089 ( .B1(n8802), .B2(n9855), .A(n7423), .ZN(P2_U3283) );
  OR2_X1 U9090 ( .A1(n7179), .A2(n7424), .ZN(n7427) );
  AND2_X1 U9091 ( .A1(n7427), .A2(n7425), .ZN(n7429) );
  NAND2_X1 U9092 ( .A1(n7427), .A2(n7426), .ZN(n7428) );
  OAI21_X1 U9093 ( .B1(n7429), .B2(n7814), .A(n7428), .ZN(n9931) );
  INV_X1 U9094 ( .A(n9810), .ZN(n7430) );
  AOI21_X1 U9095 ( .B1(n9926), .B2(n9830), .A(n7430), .ZN(n9928) );
  AOI22_X1 U9096 ( .A1(n9866), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n7431), .B2(
        n9854), .ZN(n7432) );
  OAI21_X1 U9097 ( .B1(n8693), .B2(n4559), .A(n7432), .ZN(n7440) );
  OR2_X1 U9098 ( .A1(n7433), .A2(n9816), .ZN(n9819) );
  AND2_X1 U9099 ( .A1(n9819), .A2(n7885), .ZN(n7436) );
  NAND2_X1 U9100 ( .A1(n9819), .A2(n7434), .ZN(n7435) );
  OAI21_X1 U9101 ( .B1(n7437), .B2(n7436), .A(n7435), .ZN(n7438) );
  AOI222_X1 U9102 ( .A1(n9818), .A2(n7438), .B1(n4655), .B2(n8545), .C1(n8435), 
        .C2(n8547), .ZN(n9930) );
  NOR2_X1 U9103 ( .A1(n9930), .A2(n9855), .ZN(n7439) );
  AOI211_X1 U9104 ( .C1(n9928), .C2(n8707), .A(n7440), .B(n7439), .ZN(n7441)
         );
  OAI21_X1 U9105 ( .B1(n8709), .B2(n9931), .A(n7441), .ZN(P2_U3285) );
  OAI222_X1 U9106 ( .A1(P2_U3152), .A2(n9869), .B1(n8844), .B2(n7443), .C1(
        n7442), .C2(n7714), .ZN(P2_U3332) );
  NAND2_X1 U9107 ( .A1(n7500), .A2(n7444), .ZN(n8044) );
  NAND2_X1 U9108 ( .A1(n8041), .A2(n8044), .ZN(n8120) );
  OR2_X1 U9109 ( .A1(n8039), .A2(n8120), .ZN(n7693) );
  OR2_X1 U9110 ( .A1(n7695), .A2(n7693), .ZN(n7643) );
  OR2_X1 U9111 ( .A1(n8120), .A2(n8036), .ZN(n7445) );
  AND2_X1 U9112 ( .A1(n7643), .A2(n7445), .ZN(n7474) );
  NAND2_X1 U9113 ( .A1(n8044), .A2(n8036), .ZN(n8030) );
  NAND2_X1 U9114 ( .A1(n8030), .A2(n8041), .ZN(n7642) );
  NAND2_X1 U9115 ( .A1(n7474), .A2(n7642), .ZN(n7446) );
  OR2_X1 U9116 ( .A1(n7645), .A2(n8951), .ZN(n7651) );
  NAND2_X1 U9117 ( .A1(n7645), .A2(n8951), .ZN(n7649) );
  AND2_X1 U9118 ( .A1(n7651), .A2(n7649), .ZN(n8123) );
  INV_X1 U9119 ( .A(n8123), .ZN(n8043) );
  XNOR2_X1 U9120 ( .A(n7446), .B(n8043), .ZN(n7447) );
  AOI22_X1 U9121 ( .A1(n7447), .A2(n9227), .B1(n9615), .B2(n8952), .ZN(n7632)
         );
  OR2_X1 U9122 ( .A1(n8953), .A2(n7468), .ZN(n7449) );
  AND2_X1 U9123 ( .A1(n7468), .A2(n8953), .ZN(n7448) );
  XNOR2_X1 U9124 ( .A(n7650), .B(n8123), .ZN(n7634) );
  NAND2_X1 U9125 ( .A1(n7634), .A2(n9231), .ZN(n7459) );
  INV_X1 U9126 ( .A(n7645), .ZN(n7637) );
  INV_X1 U9127 ( .A(n7658), .ZN(n7451) );
  OAI211_X1 U9128 ( .C1(n7637), .C2(n7452), .A(n7451), .B(n9626), .ZN(n7631)
         );
  INV_X1 U9129 ( .A(n7631), .ZN(n7457) );
  OAI22_X1 U9130 ( .A1(n9219), .A2(n5947), .B1(n7591), .B2(n9206), .ZN(n7453)
         );
  AOI21_X1 U9131 ( .B1(n7454), .B2(n8950), .A(n7453), .ZN(n7455) );
  OAI21_X1 U9132 ( .B1(n7637), .B2(n9204), .A(n7455), .ZN(n7456) );
  AOI21_X1 U9133 ( .B1(n7457), .B2(n9629), .A(n7456), .ZN(n7458) );
  OAI211_X1 U9134 ( .C1(n9620), .C2(n7632), .A(n7459), .B(n7458), .ZN(P1_U3280) );
  INV_X1 U9135 ( .A(n7582), .ZN(n7461) );
  AOI21_X1 U9136 ( .B1(n7462), .B2(n7460), .A(n7461), .ZN(n7470) );
  NOR2_X1 U9137 ( .A1(n8905), .A2(n9706), .ZN(n7463) );
  AOI211_X1 U9138 ( .C1(n8922), .C2(n8952), .A(n7464), .B(n7463), .ZN(n7465)
         );
  OAI21_X1 U9139 ( .B1(n8940), .B2(n7466), .A(n7465), .ZN(n7467) );
  AOI21_X1 U9140 ( .B1(n8942), .B2(n7468), .A(n7467), .ZN(n7469) );
  OAI21_X1 U9141 ( .B1(n7470), .B2(n8944), .A(n7469), .ZN(P1_U3229) );
  OAI21_X1 U9142 ( .B1(n7472), .B2(n8120), .A(n7471), .ZN(n9452) );
  INV_X1 U9143 ( .A(n9452), .ZN(n7488) );
  INV_X1 U9144 ( .A(n8120), .ZN(n7476) );
  OR2_X1 U9145 ( .A1(n7695), .A2(n8039), .ZN(n7473) );
  NAND2_X1 U9146 ( .A1(n7473), .A2(n8036), .ZN(n7475) );
  OAI21_X1 U9147 ( .B1(n7476), .B2(n7475), .A(n7474), .ZN(n7478) );
  INV_X1 U9148 ( .A(n8951), .ZN(n7644) );
  OAI22_X1 U9149 ( .A1(n7494), .A2(n9217), .B1(n7644), .B2(n9705), .ZN(n7477)
         );
  AOI21_X1 U9150 ( .B1(n7478), .B2(n9227), .A(n7477), .ZN(n7479) );
  OAI21_X1 U9151 ( .B1(n7488), .B2(n9610), .A(n7479), .ZN(n9450) );
  NAND2_X1 U9152 ( .A1(n9450), .A2(n9219), .ZN(n7487) );
  OAI22_X1 U9153 ( .A1(n9219), .A2(n7480), .B1(n7498), .B2(n9206), .ZN(n7485)
         );
  INV_X1 U9154 ( .A(n7481), .ZN(n7483) );
  INV_X1 U9155 ( .A(n7500), .ZN(n9449) );
  OAI211_X1 U9156 ( .C1(n7483), .C2(n9449), .A(n9626), .B(n7482), .ZN(n9448)
         );
  NOR2_X1 U9157 ( .A1(n9448), .A2(n9239), .ZN(n7484) );
  AOI211_X1 U9158 ( .C1(n9622), .C2(n7500), .A(n7485), .B(n7484), .ZN(n7486)
         );
  OAI211_X1 U9159 ( .C1(n7488), .C2(n7730), .A(n7487), .B(n7486), .ZN(P1_U3281) );
  NAND2_X1 U9160 ( .A1(n7582), .A2(n7489), .ZN(n7492) );
  NAND2_X1 U9161 ( .A1(n7583), .A2(n7490), .ZN(n7491) );
  XNOR2_X1 U9162 ( .A(n7492), .B(n7491), .ZN(n7502) );
  INV_X1 U9163 ( .A(n7493), .ZN(n7496) );
  NOR2_X1 U9164 ( .A1(n8905), .A2(n7494), .ZN(n7495) );
  AOI211_X1 U9165 ( .C1(n8922), .C2(n8951), .A(n7496), .B(n7495), .ZN(n7497)
         );
  OAI21_X1 U9166 ( .B1(n8940), .B2(n7498), .A(n7497), .ZN(n7499) );
  AOI21_X1 U9167 ( .B1(n8942), .B2(n7500), .A(n7499), .ZN(n7501) );
  OAI21_X1 U9168 ( .B1(n7502), .B2(n8944), .A(n7501), .ZN(P1_U3215) );
  NOR2_X1 U9169 ( .A1(n7503), .A2(n7918), .ZN(n7504) );
  OR2_X1 U9170 ( .A1(n7505), .A2(n7504), .ZN(n8778) );
  OR2_X1 U9171 ( .A1(n7605), .A2(n7506), .ZN(n8696) );
  NAND2_X1 U9172 ( .A1(n8696), .A2(n7507), .ZN(n7508) );
  XNOR2_X1 U9173 ( .A(n7508), .B(n7918), .ZN(n7509) );
  NAND2_X1 U9174 ( .A1(n7509), .A2(n9818), .ZN(n7512) );
  NAND2_X1 U9175 ( .A1(n8432), .A2(n8545), .ZN(n7511) );
  NAND2_X1 U9176 ( .A1(n8430), .A2(n8547), .ZN(n7510) );
  AND2_X1 U9177 ( .A1(n7511), .A2(n7510), .ZN(n7559) );
  NAND2_X1 U9178 ( .A1(n7512), .A2(n7559), .ZN(n8780) );
  INV_X1 U9179 ( .A(n8834), .ZN(n7564) );
  NAND2_X1 U9180 ( .A1(n8689), .A2(n8834), .ZN(n7513) );
  NAND2_X1 U9181 ( .A1(n7513), .A2(n6686), .ZN(n7514) );
  NOR2_X1 U9182 ( .A1(n8665), .A2(n7514), .ZN(n8779) );
  NAND2_X1 U9183 ( .A1(n8779), .A2(n9862), .ZN(n7516) );
  AOI22_X1 U9184 ( .A1(n9866), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n7561), .B2(
        n9854), .ZN(n7515) );
  OAI211_X1 U9185 ( .C1(n7564), .C2(n8693), .A(n7516), .B(n7515), .ZN(n7517)
         );
  AOI21_X1 U9186 ( .B1(n8780), .B2(n8579), .A(n7517), .ZN(n7518) );
  OAI21_X1 U9187 ( .B1(n8778), .B2(n8709), .A(n7518), .ZN(P2_U3280) );
  INV_X1 U9188 ( .A(n7519), .ZN(n7521) );
  OAI222_X1 U9189 ( .A1(n7688), .A2(n7520), .B1(n9391), .B2(n7521), .C1(n9479), 
        .C2(P1_U3084), .ZN(P1_U3326) );
  OAI222_X1 U9190 ( .A1(n7714), .A2(n7522), .B1(n8844), .B2(n7521), .C1(n8002), 
        .C2(P2_U3152), .ZN(P2_U3331) );
  XNOR2_X1 U9191 ( .A(n7525), .B(n7524), .ZN(n7526) );
  XNOR2_X1 U9192 ( .A(n7523), .B(n7526), .ZN(n7532) );
  INV_X1 U9193 ( .A(n9225), .ZN(n8048) );
  OAI21_X1 U9194 ( .B1(n8936), .B2(n8048), .A(n7527), .ZN(n7528) );
  AOI21_X1 U9195 ( .B1(n8938), .B2(n8950), .A(n7528), .ZN(n7529) );
  OAI21_X1 U9196 ( .B1(n8940), .B2(n7724), .A(n7529), .ZN(n7530) );
  AOI21_X1 U9197 ( .B1(n8942), .B2(n7723), .A(n7530), .ZN(n7531) );
  OAI21_X1 U9198 ( .B1(n7532), .B2(n8944), .A(n7531), .ZN(P1_U3232) );
  NAND2_X1 U9199 ( .A1(n7582), .A2(n7533), .ZN(n7588) );
  NAND2_X1 U9200 ( .A1(n7588), .A2(n7534), .ZN(n7537) );
  AND2_X1 U9201 ( .A1(n7588), .A2(n7535), .ZN(n7536) );
  AOI21_X1 U9202 ( .B1(n7538), .B2(n7537), .A(n7536), .ZN(n7544) );
  INV_X1 U9203 ( .A(n9459), .ZN(n7698) );
  OAI21_X1 U9204 ( .B1(n8936), .B2(n7698), .A(n7539), .ZN(n7540) );
  AOI21_X1 U9205 ( .B1(n8938), .B2(n8951), .A(n7540), .ZN(n7541) );
  OAI21_X1 U9206 ( .B1(n8940), .B2(n7655), .A(n7541), .ZN(n7542) );
  AOI21_X1 U9207 ( .B1(n8942), .B2(n9460), .A(n7542), .ZN(n7543) );
  OAI21_X1 U9208 ( .B1(n7544), .B2(n8944), .A(n7543), .ZN(P1_U3222) );
  INV_X1 U9209 ( .A(n7545), .ZN(n7712) );
  AOI21_X1 U9210 ( .B1(n9389), .B2(P2_DATAO_REG_28__SCAN_IN), .A(n7546), .ZN(
        n7547) );
  OAI21_X1 U9211 ( .B1(n7712), .B2(n9391), .A(n7547), .ZN(P1_U3325) );
  NOR2_X1 U9212 ( .A1(n8674), .A2(n7321), .ZN(n7549) );
  XNOR2_X1 U9213 ( .A(n8834), .B(n4296), .ZN(n7548) );
  NOR2_X1 U9214 ( .A1(n7548), .A2(n7549), .ZN(n7623) );
  AOI21_X1 U9215 ( .B1(n7549), .B2(n7548), .A(n7623), .ZN(n7556) );
  INV_X1 U9216 ( .A(n7552), .ZN(n7555) );
  INV_X1 U9217 ( .A(n7551), .ZN(n7554) );
  OAI21_X1 U9218 ( .B1(n7556), .B2(n4377), .A(n7625), .ZN(n7557) );
  NAND2_X1 U9219 ( .A1(n7557), .A2(n8352), .ZN(n7563) );
  OAI22_X1 U9220 ( .A1(n8417), .A2(n7559), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7558), .ZN(n7560) );
  AOI21_X1 U9221 ( .B1(n7561), .B2(n8375), .A(n7560), .ZN(n7562) );
  OAI211_X1 U9222 ( .C1(n7564), .C2(n8360), .A(n7563), .B(n7562), .ZN(P2_U3228) );
  XNOR2_X1 U9223 ( .A(n7572), .B(P2_REG2_REG_17__SCAN_IN), .ZN(n9784) );
  OAI21_X1 U9224 ( .B1(n7566), .B2(n7571), .A(n7565), .ZN(n9785) );
  NAND2_X1 U9225 ( .A1(n9784), .A2(n9785), .ZN(n9782) );
  OAI21_X1 U9226 ( .B1(n7572), .B2(n7567), .A(n9782), .ZN(n8445) );
  XNOR2_X1 U9227 ( .A(n8445), .B(n8451), .ZN(n7568) );
  NAND2_X1 U9228 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n7568), .ZN(n8448) );
  OAI21_X1 U9229 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n7568), .A(n8448), .ZN(
        n7580) );
  INV_X1 U9230 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10186) );
  NAND2_X1 U9231 ( .A1(P2_U3152), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n7681) );
  OAI21_X1 U9232 ( .B1(n8464), .B2(n10186), .A(n7681), .ZN(n7577) );
  INV_X1 U9233 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8775) );
  INV_X1 U9234 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n7570) );
  AOI21_X1 U9235 ( .B1(n7571), .B2(n7570), .A(n7569), .ZN(n9789) );
  XNOR2_X1 U9236 ( .A(n7572), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n9788) );
  NAND2_X1 U9237 ( .A1(n9789), .A2(n9788), .ZN(n9787) );
  OAI21_X1 U9238 ( .B1(n7572), .B2(n8775), .A(n9787), .ZN(n7574) );
  INV_X1 U9239 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8452) );
  AOI22_X1 U9240 ( .A1(P2_REG1_REG_18__SCAN_IN), .A2(n8451), .B1(n8446), .B2(
        n8452), .ZN(n7573) );
  NOR2_X1 U9241 ( .A1(n7574), .A2(n7573), .ZN(n8450) );
  AOI21_X1 U9242 ( .B1(n7574), .B2(n7573), .A(n8450), .ZN(n7575) );
  NOR2_X1 U9243 ( .A1(n7575), .A2(n9735), .ZN(n7576) );
  AOI211_X1 U9244 ( .C1(n9791), .C2(n8446), .A(n7577), .B(n7576), .ZN(n7578)
         );
  OAI21_X1 U9245 ( .B1(n7580), .B2(n7579), .A(n7578), .ZN(P2_U3263) );
  NAND2_X1 U9246 ( .A1(n7582), .A2(n7581), .ZN(n7584) );
  AND2_X1 U9247 ( .A1(n7584), .A2(n7583), .ZN(n7586) );
  AOI21_X1 U9248 ( .B1(n7586), .B2(n7585), .A(n8944), .ZN(n7590) );
  AND2_X1 U9249 ( .A1(n7588), .A2(n7587), .ZN(n7589) );
  NAND2_X1 U9250 ( .A1(n7590), .A2(n7589), .ZN(n7595) );
  NOR2_X1 U9251 ( .A1(n8940), .A2(n7591), .ZN(n7593) );
  INV_X1 U9252 ( .A(n8950), .ZN(n7641) );
  NAND2_X1 U9253 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3084), .ZN(n9547) );
  OAI21_X1 U9254 ( .B1(n8936), .B2(n7641), .A(n9547), .ZN(n7592) );
  AOI211_X1 U9255 ( .C1(n8938), .C2(n8952), .A(n7593), .B(n7592), .ZN(n7594)
         );
  OAI211_X1 U9256 ( .C1(n7637), .C2(n8910), .A(n7595), .B(n7594), .ZN(P1_U3234) );
  OAI21_X1 U9257 ( .B1(n7597), .B2(n7902), .A(n7596), .ZN(n7598) );
  INV_X1 U9258 ( .A(n7598), .ZN(n8795) );
  INV_X1 U9259 ( .A(n7599), .ZN(n7601) );
  INV_X1 U9260 ( .A(n8690), .ZN(n7600) );
  AOI21_X1 U9261 ( .B1(n8791), .B2(n7601), .A(n7600), .ZN(n8792) );
  AOI22_X1 U9262 ( .A1(n9866), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n7602), .B2(
        n9854), .ZN(n7603) );
  OAI21_X1 U9263 ( .B1(n7604), .B2(n8693), .A(n7603), .ZN(n7611) );
  AOI21_X1 U9264 ( .B1(n7605), .B2(n7902), .A(n9843), .ZN(n7609) );
  OR2_X1 U9265 ( .A1(n7605), .A2(n7902), .ZN(n8701) );
  OAI22_X1 U9266 ( .A1(n7607), .A2(n9848), .B1(n7606), .B2(n9846), .ZN(n7608)
         );
  AOI21_X1 U9267 ( .B1(n7609), .B2(n8701), .A(n7608), .ZN(n8794) );
  NOR2_X1 U9268 ( .A1(n8794), .A2(n9855), .ZN(n7610) );
  AOI211_X1 U9269 ( .C1(n8792), .C2(n8707), .A(n7611), .B(n7610), .ZN(n7612)
         );
  OAI21_X1 U9270 ( .B1(n8795), .B2(n8709), .A(n7612), .ZN(P2_U3282) );
  XNOR2_X1 U9271 ( .A(n7615), .B(n7614), .ZN(n7616) );
  XNOR2_X1 U9272 ( .A(n7613), .B(n7616), .ZN(n7622) );
  NOR2_X1 U9273 ( .A1(n8905), .A2(n7698), .ZN(n7617) );
  AOI211_X1 U9274 ( .C1(n8922), .C2(n8949), .A(n7618), .B(n7617), .ZN(n7619)
         );
  OAI21_X1 U9275 ( .B1(n8940), .B2(n7705), .A(n7619), .ZN(n7620) );
  AOI21_X1 U9276 ( .B1(n8942), .B2(n8257), .A(n7620), .ZN(n7621) );
  OAI21_X1 U9277 ( .B1(n7622), .B2(n8944), .A(n7621), .ZN(P1_U3213) );
  INV_X1 U9278 ( .A(n7623), .ZN(n7624) );
  XNOR2_X1 U9279 ( .A(n8668), .B(n4296), .ZN(n7676) );
  NOR2_X1 U9280 ( .A1(n8654), .A2(n7321), .ZN(n7677) );
  XNOR2_X1 U9281 ( .A(n7676), .B(n7677), .ZN(n7678) );
  XNOR2_X1 U9282 ( .A(n7679), .B(n7678), .ZN(n7630) );
  OAI22_X1 U9283 ( .A1(n8403), .A2(n8675), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5278), .ZN(n7628) );
  INV_X1 U9284 ( .A(n8683), .ZN(n7626) );
  OAI22_X1 U9285 ( .A1(n8404), .A2(n8674), .B1(n8411), .B2(n7626), .ZN(n7627)
         );
  AOI211_X1 U9286 ( .C1(n8668), .C2(n8420), .A(n7628), .B(n7627), .ZN(n7629)
         );
  OAI21_X1 U9287 ( .B1(n7630), .B2(n8422), .A(n7629), .ZN(P2_U3230) );
  OAI211_X1 U9288 ( .C1(n7641), .C2(n9705), .A(n7632), .B(n7631), .ZN(n7633)
         );
  AOI21_X1 U9289 ( .B1(n7634), .B2(n9710), .A(n7633), .ZN(n7640) );
  AOI22_X1 U9290 ( .A1(n7645), .A2(n5756), .B1(n9731), .B2(
        P1_REG1_REG_11__SCAN_IN), .ZN(n7635) );
  OAI21_X1 U9291 ( .B1(n7640), .B2(n9731), .A(n7635), .ZN(P1_U3534) );
  INV_X1 U9292 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n7636) );
  OAI22_X1 U9293 ( .A1(n7637), .A2(n9379), .B1(n9720), .B2(n7636), .ZN(n7638)
         );
  INV_X1 U9294 ( .A(n7638), .ZN(n7639) );
  OAI21_X1 U9295 ( .B1(n7640), .B2(n9718), .A(n7639), .ZN(P1_U3487) );
  NAND2_X1 U9296 ( .A1(n9460), .A2(n7641), .ZN(n8165) );
  NAND2_X1 U9297 ( .A1(n7645), .A2(n7644), .ZN(n8007) );
  NAND2_X1 U9298 ( .A1(n7643), .A2(n8164), .ZN(n7646) );
  OR2_X1 U9299 ( .A1(n7645), .A2(n7644), .ZN(n7692) );
  NAND2_X1 U9300 ( .A1(n7646), .A2(n7692), .ZN(n7647) );
  XOR2_X1 U9301 ( .A(n8125), .B(n7647), .Z(n7648) );
  AOI22_X1 U9302 ( .A1(n7648), .A2(n9227), .B1(n9615), .B2(n8951), .ZN(n9463)
         );
  INV_X1 U9303 ( .A(n7690), .ZN(n7653) );
  AOI21_X1 U9304 ( .B1(n8125), .B2(n7654), .A(n7653), .ZN(n9465) );
  NAND2_X1 U9305 ( .A1(n9465), .A2(n9231), .ZN(n7663) );
  INV_X1 U9306 ( .A(n7655), .ZN(n7656) );
  AOI22_X1 U9307 ( .A1(n9620), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n7656), .B2(
        n9646), .ZN(n7657) );
  OAI21_X1 U9308 ( .B1(n9235), .B2(n7698), .A(n7657), .ZN(n7661) );
  OAI211_X1 U9309 ( .C1(n7659), .C2(n7658), .A(n4315), .B(n9626), .ZN(n9461)
         );
  NOR2_X1 U9310 ( .A1(n9461), .A2(n9239), .ZN(n7660) );
  AOI211_X1 U9311 ( .C1(n9622), .C2(n9460), .A(n7661), .B(n7660), .ZN(n7662)
         );
  OAI211_X1 U9312 ( .C1(n9620), .C2(n9463), .A(n7663), .B(n7662), .ZN(P1_U3279) );
  XOR2_X1 U9313 ( .A(n7665), .B(n7664), .Z(n7666) );
  XNOR2_X1 U9314 ( .A(n7667), .B(n7666), .ZN(n7672) );
  NAND2_X1 U9315 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9549) );
  OAI21_X1 U9316 ( .B1(n8905), .B2(n8048), .A(n9549), .ZN(n7668) );
  AOI21_X1 U9317 ( .B1(n8922), .B2(n8948), .A(n7668), .ZN(n7669) );
  OAI21_X1 U9318 ( .B1(n8940), .B2(n9232), .A(n7669), .ZN(n7670) );
  AOI21_X1 U9319 ( .B1(n9328), .B2(n8942), .A(n7670), .ZN(n7671) );
  OAI21_X1 U9320 ( .B1(n7672), .B2(n8944), .A(n7671), .ZN(P1_U3239) );
  INV_X1 U9321 ( .A(n7673), .ZN(n7687) );
  OAI222_X1 U9322 ( .A1(n8844), .A2(n7687), .B1(P2_U3152), .B2(n7675), .C1(
        n7674), .C2(n7714), .ZN(P2_U3329) );
  XNOR2_X1 U9323 ( .A(n8769), .B(n4296), .ZN(n7732) );
  NAND2_X1 U9324 ( .A1(n8429), .A2(n6682), .ZN(n7731) );
  XNOR2_X1 U9325 ( .A(n7732), .B(n7731), .ZN(n7734) );
  XNOR2_X1 U9326 ( .A(n7735), .B(n7734), .ZN(n7685) );
  AOI22_X1 U9327 ( .A1(n7680), .A2(n8430), .B1(n8375), .B2(n8659), .ZN(n7682)
         );
  OAI211_X1 U9328 ( .C1(n8655), .C2(n8403), .A(n7682), .B(n7681), .ZN(n7683)
         );
  AOI21_X1 U9329 ( .B1(n8769), .B2(n8420), .A(n7683), .ZN(n7684) );
  OAI21_X1 U9330 ( .B1(n7685), .B2(n8422), .A(n7684), .ZN(P2_U3240) );
  OAI222_X1 U9331 ( .A1(n7688), .A2(n10089), .B1(n9391), .B2(n7687), .C1(n7686), .C2(P1_U3084), .ZN(P1_U3324) );
  XNOR2_X1 U9332 ( .A(n8257), .B(n8048), .ZN(n8129) );
  NAND2_X1 U9333 ( .A1(n9460), .A2(n8950), .ZN(n7689) );
  OR2_X1 U9334 ( .A1(n7723), .A2(n9459), .ZN(n7691) );
  XOR2_X1 U9335 ( .A(n8129), .B(n8258), .Z(n9458) );
  INV_X1 U9336 ( .A(n9458), .ZN(n7711) );
  AND2_X1 U9337 ( .A1(n8034), .A2(n7692), .ZN(n8047) );
  INV_X1 U9338 ( .A(n8047), .ZN(n7696) );
  OR2_X1 U9339 ( .A1(n7693), .A2(n7696), .ZN(n7694) );
  OR2_X1 U9340 ( .A1(n7696), .A2(n8164), .ZN(n7716) );
  AND2_X1 U9341 ( .A1(n8165), .A2(n7716), .ZN(n7697) );
  NAND2_X1 U9342 ( .A1(n7717), .A2(n7697), .ZN(n7699) );
  OR2_X1 U9343 ( .A1(n7723), .A2(n7698), .ZN(n8049) );
  NAND2_X1 U9344 ( .A1(n7723), .A2(n7698), .ZN(n8008) );
  INV_X1 U9345 ( .A(n8129), .ZN(n7700) );
  NAND2_X1 U9346 ( .A1(n7701), .A2(n8129), .ZN(n7702) );
  NAND3_X1 U9347 ( .A1(n8296), .A2(n9227), .A3(n7702), .ZN(n7704) );
  AOI22_X1 U9348 ( .A1(n9226), .A2(n9459), .B1(n8949), .B2(n9686), .ZN(n7703)
         );
  NAND2_X1 U9349 ( .A1(n7704), .A2(n7703), .ZN(n9457) );
  OAI211_X1 U9350 ( .C1(n4381), .C2(n4584), .A(n9626), .B(n4852), .ZN(n9455)
         );
  OAI22_X1 U9351 ( .A1(n9219), .A2(n7706), .B1(n7705), .B2(n9206), .ZN(n7707)
         );
  AOI21_X1 U9352 ( .B1(n8257), .B2(n9622), .A(n7707), .ZN(n7708) );
  OAI21_X1 U9353 ( .B1(n9455), .B2(n9239), .A(n7708), .ZN(n7709) );
  AOI21_X1 U9354 ( .B1(n9457), .B2(n9219), .A(n7709), .ZN(n7710) );
  OAI21_X1 U9355 ( .B1(n7711), .B2(n9222), .A(n7710), .ZN(P1_U3277) );
  OAI222_X1 U9356 ( .A1(n7714), .A2(n7713), .B1(P2_U3152), .B2(n5459), .C1(
        n8844), .C2(n7712), .ZN(P2_U3330) );
  XOR2_X1 U9357 ( .A(n7715), .B(n8127), .Z(n9336) );
  AOI22_X1 U9358 ( .A1(n9615), .A2(n8950), .B1(n9225), .B2(n9686), .ZN(n7722)
         );
  INV_X1 U9359 ( .A(n8165), .ZN(n8046) );
  NOR3_X1 U9360 ( .A1(n4360), .A2(n8046), .A3(n8127), .ZN(n7720) );
  INV_X1 U9361 ( .A(n7718), .ZN(n7719) );
  OAI21_X1 U9362 ( .B1(n7720), .B2(n7719), .A(n9227), .ZN(n7721) );
  OAI211_X1 U9363 ( .C1(n9336), .C2(n9610), .A(n7722), .B(n7721), .ZN(n9337)
         );
  NAND2_X1 U9364 ( .A1(n9337), .A2(n9219), .ZN(n7729) );
  AOI211_X1 U9365 ( .C1(n7723), .C2(n4315), .A(n9236), .B(n4381), .ZN(n9338)
         );
  NOR2_X1 U9366 ( .A1(n9380), .A2(n9204), .ZN(n7727) );
  OAI22_X1 U9367 ( .A1(n9219), .A2(n7725), .B1(n7724), .B2(n9206), .ZN(n7726)
         );
  AOI211_X1 U9368 ( .C1(n9338), .C2(n9629), .A(n7727), .B(n7726), .ZN(n7728)
         );
  OAI211_X1 U9369 ( .C1(n7730), .C2(n9336), .A(n7729), .B(n7728), .ZN(P1_U3278) );
  INV_X1 U9370 ( .A(n7731), .ZN(n7733) );
  AND2_X1 U9371 ( .A1(n8428), .A2(n6682), .ZN(n7737) );
  XNOR2_X1 U9372 ( .A(n8639), .B(n4296), .ZN(n7736) );
  NOR2_X1 U9373 ( .A1(n7736), .A2(n7737), .ZN(n7738) );
  AOI21_X1 U9374 ( .B1(n7737), .B2(n7736), .A(n7738), .ZN(n8350) );
  NAND2_X1 U9375 ( .A1(n8351), .A2(n8350), .ZN(n8349) );
  INV_X1 U9376 ( .A(n7738), .ZN(n7739) );
  XNOR2_X1 U9377 ( .A(n8757), .B(n4296), .ZN(n7740) );
  NOR2_X1 U9378 ( .A1(n8638), .A2(n7321), .ZN(n7741) );
  XNOR2_X1 U9379 ( .A(n7740), .B(n7741), .ZN(n8391) );
  XNOR2_X1 U9380 ( .A(n8602), .B(n4296), .ZN(n7742) );
  NOR2_X1 U9381 ( .A1(n8617), .A2(n7321), .ZN(n7744) );
  XNOR2_X1 U9382 ( .A(n7742), .B(n7744), .ZN(n8361) );
  INV_X1 U9383 ( .A(n7742), .ZN(n7743) );
  NOR2_X1 U9384 ( .A1(n8363), .A2(n6686), .ZN(n8401) );
  NOR2_X1 U9385 ( .A1(n8400), .A2(n8401), .ZN(n8399) );
  NOR2_X1 U9386 ( .A1(n8399), .A2(n7746), .ZN(n7752) );
  XNOR2_X1 U9387 ( .A(n8819), .B(n4296), .ZN(n7753) );
  XNOR2_X1 U9388 ( .A(n8735), .B(n4296), .ZN(n8383) );
  AND2_X1 U9389 ( .A1(n8546), .A2(n6682), .ZN(n8380) );
  INV_X1 U9390 ( .A(n8383), .ZN(n7749) );
  NOR2_X1 U9391 ( .A1(n8372), .A2(n6686), .ZN(n8382) );
  INV_X1 U9392 ( .A(n8382), .ZN(n7748) );
  INV_X1 U9393 ( .A(n7752), .ZN(n7754) );
  OAI21_X1 U9394 ( .B1(n8382), .B2(n8383), .A(n8379), .ZN(n7755) );
  NAND2_X1 U9395 ( .A1(n7756), .A2(n7755), .ZN(n8371) );
  NOR2_X1 U9396 ( .A1(n8413), .A2(n7321), .ZN(n7758) );
  XNOR2_X1 U9397 ( .A(n8731), .B(n4296), .ZN(n7757) );
  XOR2_X1 U9398 ( .A(n7758), .B(n7757), .Z(n8370) );
  XNOR2_X1 U9399 ( .A(n8814), .B(n4296), .ZN(n7760) );
  NAND2_X1 U9400 ( .A1(n8504), .A2(n6682), .ZN(n7759) );
  XNOR2_X1 U9401 ( .A(n7760), .B(n7759), .ZN(n8409) );
  XNOR2_X1 U9402 ( .A(n8500), .B(n4296), .ZN(n7761) );
  NOR2_X1 U9403 ( .A1(n8412), .A2(n6686), .ZN(n7762) );
  XNOR2_X1 U9404 ( .A(n7761), .B(n7762), .ZN(n8333) );
  INV_X1 U9405 ( .A(n7761), .ZN(n7763) );
  NOR2_X1 U9406 ( .A1(n8336), .A2(n6686), .ZN(n7765) );
  XNOR2_X1 U9407 ( .A(n7765), .B(n4296), .ZN(n7766) );
  XNOR2_X1 U9408 ( .A(n7772), .B(n7766), .ZN(n7767) );
  NOR2_X1 U9409 ( .A1(n8484), .A2(n8411), .ZN(n7771) );
  OAI22_X1 U9410 ( .A1(n7769), .A2(n8417), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7768), .ZN(n7770) );
  AOI211_X1 U9411 ( .C1(n7772), .C2(n8420), .A(n7771), .B(n7770), .ZN(n7773)
         );
  OAI21_X1 U9412 ( .B1(n7774), .B2(n8422), .A(n7773), .ZN(P2_U3222) );
  XOR2_X1 U9413 ( .A(n7810), .B(n7775), .Z(n9900) );
  AOI211_X1 U9414 ( .C1(n9897), .C2(n4380), .A(n6682), .B(n7776), .ZN(n9896)
         );
  OAI22_X1 U9415 ( .A1(n8693), .A2(n7859), .B1(n8556), .B2(n7777), .ZN(n7778)
         );
  AOI21_X1 U9416 ( .B1(n9896), .B2(n9862), .A(n7778), .ZN(n7787) );
  INV_X1 U9417 ( .A(n7810), .ZN(n7779) );
  NAND3_X1 U9418 ( .A1(n7780), .A2(n7779), .A3(n7834), .ZN(n7781) );
  NAND2_X1 U9419 ( .A1(n7782), .A2(n7781), .ZN(n7785) );
  NAND2_X1 U9420 ( .A1(n8441), .A2(n8545), .ZN(n7783) );
  OAI21_X1 U9421 ( .B1(n9847), .B2(n9848), .A(n7783), .ZN(n7784) );
  AOI21_X1 U9422 ( .B1(n7785), .B2(n9818), .A(n7784), .ZN(n9899) );
  MUX2_X1 U9423 ( .A(n6456), .B(n9899), .S(n8579), .Z(n7786) );
  OAI211_X1 U9424 ( .C1(n9900), .C2(n8709), .A(n7787), .B(n7786), .ZN(P2_U3290) );
  NAND2_X1 U9425 ( .A1(n8840), .A2(n7792), .ZN(n7790) );
  NAND2_X1 U9426 ( .A1(n7788), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n7789) );
  NAND2_X1 U9427 ( .A1(n8810), .A2(n8466), .ZN(n8465) );
  NAND2_X1 U9428 ( .A1(n7791), .A2(n7792), .ZN(n7794) );
  NAND2_X1 U9429 ( .A1(n5092), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n7793) );
  XNOR2_X1 U9430 ( .A(n8465), .B(n7799), .ZN(n8710) );
  OR2_X1 U9431 ( .A1(n7988), .A2(n7795), .ZN(n8715) );
  NOR2_X1 U9432 ( .A1(n9866), .A2(n8715), .ZN(n8468) );
  INV_X1 U9433 ( .A(n7799), .ZN(n8806) );
  NOR2_X1 U9434 ( .A1(n8806), .A2(n8693), .ZN(n7796) );
  AOI211_X1 U9435 ( .C1(n9866), .C2(P2_REG2_REG_31__SCAN_IN), .A(n8468), .B(
        n7796), .ZN(n7797) );
  OAI21_X1 U9436 ( .B1(n8710), .B2(n7798), .A(n7797), .ZN(P2_U3265) );
  NAND2_X1 U9437 ( .A1(n7799), .A2(n7988), .ZN(n7993) );
  INV_X1 U9438 ( .A(n7800), .ZN(n8424) );
  NAND2_X1 U9439 ( .A1(n8810), .A2(n8424), .ZN(n7990) );
  NAND2_X1 U9440 ( .A1(n7993), .A2(n7990), .ZN(n7979) );
  INV_X1 U9441 ( .A(n7979), .ZN(n7827) );
  INV_X1 U9442 ( .A(n8810), .ZN(n7801) );
  NAND2_X1 U9443 ( .A1(n7801), .A2(n7800), .ZN(n7974) );
  NAND2_X1 U9444 ( .A1(n7982), .A2(n7974), .ZN(n7994) );
  INV_X1 U9445 ( .A(n7994), .ZN(n7977) );
  INV_X1 U9446 ( .A(n8530), .ZN(n8527) );
  INV_X1 U9447 ( .A(n7802), .ZN(n8632) );
  INV_X1 U9448 ( .A(n7803), .ZN(n7804) );
  NAND4_X1 U9449 ( .A1(n7848), .A2(n7805), .A3(n7804), .A4(n7829), .ZN(n7809)
         );
  NOR4_X1 U9450 ( .A1(n7809), .A2(n7808), .A3(n7807), .A4(n7806), .ZN(n7813)
         );
  INV_X1 U9451 ( .A(n7869), .ZN(n7812) );
  NAND4_X1 U9452 ( .A1(n7813), .A2(n7812), .A3(n7811), .A4(n7810), .ZN(n7815)
         );
  NOR4_X1 U9453 ( .A1(n7815), .A2(n7814), .A3(n9816), .A4(n9841), .ZN(n7816)
         );
  NAND3_X1 U9454 ( .A1(n7817), .A2(n9800), .A3(n7816), .ZN(n7818) );
  NOR4_X1 U9455 ( .A1(n7918), .A2(n7909), .A3(n7902), .A4(n7818), .ZN(n7819)
         );
  NAND4_X1 U9456 ( .A1(n8632), .A2(n8671), .A3(n8651), .A4(n7819), .ZN(n7820)
         );
  NOR4_X1 U9457 ( .A1(n8566), .A2(n8590), .A3(n8620), .A4(n7820), .ZN(n7821)
         );
  INV_X1 U9458 ( .A(n8597), .ZN(n8604) );
  NAND4_X1 U9459 ( .A1(n8527), .A2(n7822), .A3(n7821), .A4(n8604), .ZN(n7823)
         );
  NOR4_X1 U9460 ( .A1(n7824), .A2(n8501), .A3(n8515), .A4(n7823), .ZN(n7825)
         );
  NAND4_X1 U9461 ( .A1(n7827), .A2(n7826), .A3(n7977), .A4(n7825), .ZN(n7828)
         );
  XNOR2_X1 U9462 ( .A(n7828), .B(n8682), .ZN(n7830) );
  OAI22_X1 U9463 ( .A1(n7830), .A2(n7989), .B1(n7829), .B2(n6674), .ZN(n8000)
         );
  NOR2_X1 U9464 ( .A1(n7831), .A2(n8682), .ZN(n7832) );
  NAND2_X2 U9465 ( .A1(n7833), .A2(n7832), .ZN(n7978) );
  INV_X1 U9466 ( .A(n7929), .ZN(n7932) );
  NAND2_X1 U9467 ( .A1(n7834), .A2(n7839), .ZN(n7837) );
  NAND2_X1 U9468 ( .A1(n7835), .A2(n7860), .ZN(n7836) );
  AOI21_X1 U9469 ( .B1(n7839), .B2(n7838), .A(n7862), .ZN(n7841) );
  NOR3_X1 U9470 ( .A1(n7841), .A2(n7840), .A3(n7868), .ZN(n7851) );
  INV_X1 U9471 ( .A(n7978), .ZN(n7981) );
  INV_X1 U9472 ( .A(n7842), .ZN(n7843) );
  NOR2_X1 U9473 ( .A1(n7844), .A2(n7843), .ZN(n7852) );
  AOI21_X1 U9474 ( .B1(n7852), .B2(n7989), .A(n7845), .ZN(n7847) );
  INV_X1 U9475 ( .A(n7856), .ZN(n7846) );
  OAI211_X1 U9476 ( .C1(n7847), .C2(n7846), .A(n7854), .B(n7978), .ZN(n7849)
         );
  NAND2_X1 U9477 ( .A1(n7849), .A2(n7848), .ZN(n7850) );
  OAI22_X1 U9478 ( .A1(n7851), .A2(n7981), .B1(n7850), .B2(n7862), .ZN(n7865)
         );
  INV_X1 U9479 ( .A(n7852), .ZN(n7855) );
  NAND3_X1 U9480 ( .A1(n7855), .A2(n7854), .A3(n7853), .ZN(n7857) );
  NAND3_X1 U9481 ( .A1(n7857), .A2(n7981), .A3(n7856), .ZN(n7864) );
  AND2_X1 U9482 ( .A1(n7835), .A2(n7858), .ZN(n7861) );
  NAND2_X1 U9483 ( .A1(n8440), .A2(n7859), .ZN(n7866) );
  OAI211_X1 U9484 ( .C1(n7862), .C2(n7861), .A(n7860), .B(n7866), .ZN(n7863)
         );
  AOI22_X1 U9485 ( .A1(n7865), .A2(n7864), .B1(n7981), .B2(n7863), .ZN(n7871)
         );
  INV_X1 U9486 ( .A(n7866), .ZN(n7867) );
  MUX2_X1 U9487 ( .A(n7868), .B(n7867), .S(n7978), .Z(n7870) );
  MUX2_X1 U9488 ( .A(n7873), .B(n7872), .S(n7978), .Z(n7874) );
  INV_X1 U9489 ( .A(n7875), .ZN(n7878) );
  OAI21_X1 U9490 ( .B1(n7876), .B2(n9857), .A(n7880), .ZN(n7877) );
  MUX2_X1 U9491 ( .A(n7878), .B(n7877), .S(n7978), .Z(n7879) );
  INV_X1 U9492 ( .A(n7880), .ZN(n7883) );
  NAND2_X1 U9493 ( .A1(n7884), .A2(n7881), .ZN(n7882) );
  MUX2_X1 U9494 ( .A(n7883), .B(n7882), .S(n7978), .Z(n7889) );
  AND2_X1 U9495 ( .A1(n7890), .A2(n7884), .ZN(n7887) );
  AND2_X1 U9496 ( .A1(n7894), .A2(n7885), .ZN(n7886) );
  MUX2_X1 U9497 ( .A(n7887), .B(n7886), .S(n7978), .Z(n7888) );
  NAND3_X1 U9498 ( .A1(n7896), .A2(n7890), .A3(n7897), .ZN(n7891) );
  NAND2_X1 U9499 ( .A1(n7891), .A2(n7895), .ZN(n7893) );
  NAND3_X1 U9500 ( .A1(n7896), .A2(n7895), .A3(n7894), .ZN(n7898) );
  NAND2_X1 U9501 ( .A1(n7898), .A2(n7897), .ZN(n7899) );
  INV_X1 U9502 ( .A(n7902), .ZN(n7906) );
  MUX2_X1 U9503 ( .A(n7904), .B(n7903), .S(n7978), .Z(n7905) );
  INV_X1 U9504 ( .A(n7909), .ZN(n8699) );
  MUX2_X1 U9505 ( .A(n7910), .B(n8697), .S(n7978), .Z(n7911) );
  AND2_X1 U9506 ( .A1(n8786), .A2(n7978), .ZN(n7913) );
  NOR2_X1 U9507 ( .A1(n8786), .A2(n7978), .ZN(n7912) );
  MUX2_X1 U9508 ( .A(n7913), .B(n7912), .S(n8432), .Z(n7914) );
  MUX2_X1 U9509 ( .A(n8669), .B(n7915), .S(n7978), .Z(n7916) );
  AND2_X1 U9510 ( .A1(n7924), .A2(n7919), .ZN(n7921) );
  MUX2_X1 U9511 ( .A(n7921), .B(n7920), .S(n7978), .Z(n7922) );
  INV_X1 U9512 ( .A(n7924), .ZN(n7925) );
  OAI211_X1 U9513 ( .C1(n7934), .C2(n7925), .A(n8633), .B(n7935), .ZN(n7927)
         );
  NOR2_X1 U9514 ( .A1(n8751), .A2(n8617), .ZN(n7939) );
  INV_X1 U9515 ( .A(n7928), .ZN(n8587) );
  NAND2_X1 U9516 ( .A1(n7929), .A2(n8587), .ZN(n7930) );
  OAI21_X1 U9517 ( .B1(n7934), .B2(n7933), .A(n8613), .ZN(n7936) );
  NAND3_X1 U9518 ( .A1(n7936), .A2(n8615), .A3(n7935), .ZN(n7938) );
  NAND3_X1 U9519 ( .A1(n7938), .A2(n7937), .A3(n8587), .ZN(n7942) );
  NOR3_X1 U9520 ( .A1(n7940), .A2(n7939), .A3(n7978), .ZN(n7941) );
  INV_X1 U9521 ( .A(n7943), .ZN(n7950) );
  NAND2_X1 U9522 ( .A1(n8529), .A2(n7944), .ZN(n7947) );
  NAND2_X1 U9523 ( .A1(n7951), .A2(n7945), .ZN(n7946) );
  MUX2_X1 U9524 ( .A(n7947), .B(n7946), .S(n7978), .Z(n7948) );
  MUX2_X1 U9525 ( .A(n7951), .B(n8529), .S(n7978), .Z(n7952) );
  OAI211_X1 U9526 ( .C1(n8510), .C2(n7978), .A(n7953), .B(n7958), .ZN(n7957)
         );
  NAND2_X1 U9527 ( .A1(n7956), .A2(n7954), .ZN(n7955) );
  AOI22_X1 U9528 ( .A1(n7957), .A2(n7956), .B1(n7978), .B2(n7955), .ZN(n7960)
         );
  INV_X1 U9529 ( .A(n7958), .ZN(n7959) );
  INV_X1 U9530 ( .A(n7961), .ZN(n7964) );
  NAND2_X1 U9531 ( .A1(n7967), .A2(n7962), .ZN(n7963) );
  MUX2_X1 U9532 ( .A(n7964), .B(n7963), .S(n7978), .Z(n7965) );
  NAND2_X1 U9533 ( .A1(n8482), .A2(n7978), .ZN(n7968) );
  AOI22_X1 U9534 ( .A1(n7968), .A2(n7967), .B1(n8336), .B2(n7978), .ZN(n7969)
         );
  NAND2_X1 U9535 ( .A1(n7973), .A2(n7972), .ZN(n7975) );
  NAND3_X1 U9536 ( .A1(n7975), .A2(n7990), .A3(n7974), .ZN(n7976) );
  OAI21_X1 U9537 ( .B1(n7977), .B2(n7978), .A(n7976), .ZN(n7980) );
  AOI22_X1 U9538 ( .A1(n7980), .A2(n7993), .B1(n7979), .B2(n7978), .ZN(n7985)
         );
  NOR2_X1 U9539 ( .A1(n7982), .A2(n7981), .ZN(n7984) );
  INV_X1 U9540 ( .A(n7991), .ZN(n7992) );
  NOR4_X1 U9541 ( .A1(n9868), .A2(n9846), .A3(n8002), .A4(n8001), .ZN(n8004)
         );
  OAI21_X1 U9542 ( .B1(n8005), .B2(n5453), .A(P2_B_REG_SCAN_IN), .ZN(n8003) );
  OAI22_X1 U9543 ( .A1(n8006), .A2(n8005), .B1(n8004), .B2(n8003), .ZN(
        P2_U3244) );
  NAND2_X1 U9544 ( .A1(n8165), .A2(n8007), .ZN(n8033) );
  NAND2_X1 U9545 ( .A1(n8257), .A2(n8048), .ZN(n8050) );
  NAND2_X1 U9546 ( .A1(n8050), .A2(n8008), .ZN(n8170) );
  INV_X1 U9547 ( .A(n8009), .ZN(n8010) );
  NAND2_X1 U9548 ( .A1(n4299), .A2(n9127), .ZN(n8093) );
  NAND2_X1 U9549 ( .A1(n8215), .A2(n8012), .ZN(n8157) );
  OAI21_X1 U9550 ( .B1(n8019), .B2(n8157), .A(n8155), .ZN(n8015) );
  INV_X1 U9551 ( .A(n8093), .ZN(n8014) );
  AOI21_X1 U9552 ( .B1(n8015), .B2(n8014), .A(n8013), .ZN(n8023) );
  INV_X1 U9553 ( .A(n8023), .ZN(n8018) );
  AND2_X1 U9554 ( .A1(n8024), .A2(n8016), .ZN(n8159) );
  INV_X1 U9555 ( .A(n8148), .ZN(n8017) );
  AOI21_X1 U9556 ( .B1(n8018), .B2(n8159), .A(n8017), .ZN(n8028) );
  INV_X1 U9557 ( .A(n8156), .ZN(n8022) );
  INV_X1 U9558 ( .A(n8019), .ZN(n8020) );
  NAND2_X1 U9559 ( .A1(n8020), .A2(n8219), .ZN(n8021) );
  OAI211_X1 U9560 ( .C1(n8023), .C2(n8022), .A(n8021), .B(n8153), .ZN(n8026)
         );
  INV_X1 U9561 ( .A(n8024), .ZN(n8025) );
  AOI21_X1 U9562 ( .B1(n8026), .B2(n8148), .A(n8025), .ZN(n8027) );
  NAND2_X1 U9563 ( .A1(n8035), .A2(n8149), .ZN(n8031) );
  INV_X1 U9564 ( .A(n8029), .ZN(n8037) );
  NOR2_X1 U9565 ( .A1(n8039), .A2(n8037), .ZN(n8163) );
  AOI21_X1 U9566 ( .B1(n8031), .B2(n8163), .A(n8030), .ZN(n8032) );
  INV_X1 U9567 ( .A(n8041), .ZN(n8167) );
  INV_X1 U9568 ( .A(n8035), .ZN(n8038) );
  OAI211_X1 U9569 ( .C1(n8038), .C2(n8037), .A(n8036), .B(n8149), .ZN(n8042)
         );
  INV_X1 U9570 ( .A(n8039), .ZN(n8040) );
  NAND3_X1 U9571 ( .A1(n8042), .A2(n8041), .A3(n8040), .ZN(n8045) );
  OR2_X1 U9572 ( .A1(n8257), .A2(n8048), .ZN(n8295) );
  NAND2_X1 U9573 ( .A1(n8295), .A2(n8049), .ZN(n8051) );
  NAND2_X1 U9574 ( .A1(n8051), .A2(n8050), .ZN(n8169) );
  NAND2_X1 U9575 ( .A1(n8170), .A2(n8295), .ZN(n8052) );
  MUX2_X1 U9576 ( .A(n8169), .B(n8052), .S(n8093), .Z(n8053) );
  INV_X1 U9577 ( .A(n8949), .ZN(n9216) );
  OR2_X1 U9578 ( .A1(n9328), .A2(n9216), .ZN(n8297) );
  NAND2_X1 U9579 ( .A1(n9328), .A2(n9216), .ZN(n9211) );
  AND2_X1 U9580 ( .A1(n8297), .A2(n9211), .ZN(n9223) );
  NAND2_X1 U9581 ( .A1(n9325), .A2(n9331), .ZN(n8147) );
  NAND2_X1 U9582 ( .A1(n8299), .A2(n8147), .ZN(n9213) );
  INV_X1 U9583 ( .A(n9213), .ZN(n8131) );
  MUX2_X1 U9584 ( .A(n9211), .B(n8297), .S(n8093), .Z(n8054) );
  INV_X1 U9585 ( .A(n9169), .ZN(n9218) );
  OR2_X1 U9586 ( .A1(n9320), .A2(n9218), .ZN(n9165) );
  NAND2_X1 U9587 ( .A1(n9320), .A2(n9218), .ZN(n9167) );
  AND2_X1 U9588 ( .A1(n9165), .A2(n9167), .ZN(n9196) );
  MUX2_X1 U9589 ( .A(n8299), .B(n8147), .S(n8093), .Z(n8055) );
  NAND3_X1 U9590 ( .A1(n8056), .A2(n9196), .A3(n8055), .ZN(n8058) );
  INV_X1 U9591 ( .A(n8947), .ZN(n9199) );
  NAND2_X1 U9592 ( .A1(n9313), .A2(n9199), .ZN(n8302) );
  AND2_X1 U9593 ( .A1(n8302), .A2(n9167), .ZN(n8301) );
  OR2_X1 U9594 ( .A1(n9313), .A2(n9199), .ZN(n8107) );
  NAND2_X1 U9595 ( .A1(n8107), .A2(n9165), .ZN(n8303) );
  INV_X1 U9596 ( .A(n8303), .ZN(n8182) );
  MUX2_X1 U9597 ( .A(n8301), .B(n8182), .S(n8093), .Z(n8057) );
  NAND2_X1 U9598 ( .A1(n8058), .A2(n8057), .ZN(n8063) );
  INV_X1 U9599 ( .A(n9312), .ZN(n9178) );
  OR2_X1 U9600 ( .A1(n9157), .A2(n9178), .ZN(n8106) );
  INV_X1 U9601 ( .A(n9123), .ZN(n9153) );
  NAND2_X1 U9602 ( .A1(n9141), .A2(n9153), .ZN(n8105) );
  NAND2_X1 U9603 ( .A1(n9157), .A2(n9178), .ZN(n9133) );
  AND2_X1 U9604 ( .A1(n8105), .A2(n9133), .ZN(n8305) );
  OR2_X1 U9605 ( .A1(n9141), .A2(n9153), .ZN(n8306) );
  INV_X1 U9606 ( .A(n9104), .ZN(n9136) );
  NAND2_X1 U9607 ( .A1(n9296), .A2(n9136), .ZN(n8308) );
  INV_X1 U9608 ( .A(n9295), .ZN(n9120) );
  OR2_X1 U9609 ( .A1(n9286), .A2(n9120), .ZN(n8102) );
  OR2_X1 U9610 ( .A1(n9296), .A2(n9136), .ZN(n8104) );
  AND2_X1 U9611 ( .A1(n8102), .A2(n8104), .ZN(n8062) );
  NAND2_X1 U9612 ( .A1(n9286), .A2(n9120), .ZN(n8309) );
  INV_X1 U9613 ( .A(n9092), .ZN(n8877) );
  OR2_X1 U9614 ( .A1(n9278), .A2(n8877), .ZN(n9070) );
  NAND2_X1 U9615 ( .A1(n9070), .A2(n8312), .ZN(n8189) );
  INV_X1 U9616 ( .A(n9076), .ZN(n8060) );
  NAND2_X1 U9617 ( .A1(n9065), .A2(n8060), .ZN(n8314) );
  NAND2_X1 U9618 ( .A1(n9278), .A2(n8877), .ZN(n8313) );
  NAND2_X1 U9619 ( .A1(n9096), .A2(n9289), .ZN(n8103) );
  NAND2_X1 U9620 ( .A1(n8313), .A2(n8103), .ZN(n8067) );
  NAND2_X1 U9621 ( .A1(n8067), .A2(n9070), .ZN(n8059) );
  NAND2_X1 U9622 ( .A1(n8314), .A2(n8059), .ZN(n8190) );
  OAI21_X1 U9623 ( .B1(n8061), .B2(n8190), .A(n9043), .ZN(n8072) );
  AND2_X1 U9624 ( .A1(n9133), .A2(n8302), .ZN(n8178) );
  INV_X1 U9625 ( .A(n8062), .ZN(n8186) );
  NAND2_X1 U9626 ( .A1(n8306), .A2(n8106), .ZN(n8179) );
  AOI211_X1 U9627 ( .C1(n8063), .C2(n8178), .A(n8186), .B(n8179), .ZN(n8068)
         );
  INV_X1 U9628 ( .A(n8105), .ZN(n8064) );
  NAND2_X1 U9629 ( .A1(n8104), .A2(n8064), .ZN(n8065) );
  AND2_X1 U9630 ( .A1(n8065), .A2(n8308), .ZN(n8066) );
  NAND2_X1 U9631 ( .A1(n8309), .A2(n8066), .ZN(n8146) );
  AND2_X1 U9632 ( .A1(n8146), .A2(n8102), .ZN(n8183) );
  NOR3_X1 U9633 ( .A1(n8068), .A2(n8183), .A3(n8067), .ZN(n8070) );
  OAI21_X1 U9634 ( .B1(n4449), .B2(n4532), .A(n9043), .ZN(n8069) );
  OAI21_X1 U9635 ( .B1(n8070), .B2(n8069), .A(n8314), .ZN(n8071) );
  MUX2_X1 U9636 ( .A(n8072), .B(n8071), .S(n8093), .Z(n8077) );
  NOR2_X1 U9637 ( .A1(n9265), .A2(n9028), .ZN(n8278) );
  NAND2_X1 U9638 ( .A1(n9265), .A2(n9028), .ZN(n8284) );
  INV_X1 U9639 ( .A(n8284), .ZN(n8073) );
  INV_X1 U9640 ( .A(n9046), .ZN(n8076) );
  NAND2_X1 U9641 ( .A1(n9021), .A2(n8078), .ZN(n8100) );
  INV_X1 U9642 ( .A(n9028), .ZN(n9271) );
  NAND2_X1 U9643 ( .A1(n9265), .A2(n9271), .ZN(n8316) );
  AND2_X1 U9644 ( .A1(n8100), .A2(n8316), .ZN(n8074) );
  OR2_X1 U9645 ( .A1(n9265), .A2(n9271), .ZN(n8144) );
  MUX2_X1 U9646 ( .A(n8074), .B(n8144), .S(n8093), .Z(n8075) );
  INV_X1 U9647 ( .A(n9029), .ZN(n8288) );
  NAND2_X1 U9648 ( .A1(n9015), .A2(n8288), .ZN(n8320) );
  NAND2_X1 U9649 ( .A1(n8320), .A2(n8100), .ZN(n8143) );
  INV_X1 U9650 ( .A(n9010), .ZN(n8080) );
  NAND2_X1 U9651 ( .A1(n9248), .A2(n8080), .ZN(n8237) );
  INV_X1 U9652 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n8087) );
  INV_X1 U9653 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n8081) );
  OR2_X1 U9654 ( .A1(n8082), .A2(n8081), .ZN(n8086) );
  INV_X1 U9655 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n8083) );
  OR2_X1 U9656 ( .A1(n8084), .A2(n8083), .ZN(n8085) );
  OAI211_X1 U9657 ( .C1(n8088), .C2(n8087), .A(n8086), .B(n8085), .ZN(n8946)
         );
  NAND2_X1 U9658 ( .A1(n8946), .A2(n8097), .ZN(n8089) );
  NAND2_X1 U9659 ( .A1(n8999), .A2(n8089), .ZN(n8195) );
  MUX2_X1 U9660 ( .A(n8237), .B(n8194), .S(n8093), .Z(n8090) );
  NAND2_X1 U9661 ( .A1(n8195), .A2(n8090), .ZN(n8091) );
  NOR2_X1 U9662 ( .A1(n8092), .A2(n8195), .ZN(n8094) );
  MUX2_X1 U9663 ( .A(n8140), .B(n8094), .S(n8093), .Z(n8095) );
  INV_X1 U9664 ( .A(n8946), .ZN(n8099) );
  AND2_X1 U9665 ( .A1(n8999), .A2(n8099), .ZN(n8202) );
  OR2_X1 U9666 ( .A1(n9278), .A2(n9092), .ZN(n9056) );
  INV_X1 U9667 ( .A(n9056), .ZN(n8101) );
  AND2_X1 U9668 ( .A1(n9278), .A2(n9092), .ZN(n8275) );
  OR2_X1 U9669 ( .A1(n8101), .A2(n8275), .ZN(n9073) );
  NAND2_X1 U9670 ( .A1(n8312), .A2(n8103), .ZN(n8311) );
  NAND2_X1 U9671 ( .A1(n8106), .A2(n9133), .ZN(n9154) );
  INV_X1 U9672 ( .A(n9223), .ZN(n9230) );
  NOR2_X1 U9673 ( .A1(n8108), .A2(n9612), .ZN(n8113) );
  AND2_X1 U9674 ( .A1(n6638), .A2(n8109), .ZN(n8203) );
  NOR2_X1 U9675 ( .A1(n8110), .A2(n8203), .ZN(n9636) );
  NAND4_X1 U9676 ( .A1(n8113), .A2(n8112), .A3(n8111), .A4(n9636), .ZN(n8115)
         );
  NOR2_X1 U9677 ( .A1(n8115), .A2(n8114), .ZN(n8119) );
  NAND4_X1 U9678 ( .A1(n8119), .A2(n8118), .A3(n7162), .A4(n8117), .ZN(n8122)
         );
  OR3_X1 U9679 ( .A1(n8122), .A2(n8121), .A3(n8120), .ZN(n8124) );
  NOR2_X1 U9680 ( .A1(n8124), .A2(n8123), .ZN(n8126) );
  NAND3_X1 U9681 ( .A1(n8127), .A2(n8126), .A3(n8125), .ZN(n8128) );
  NOR3_X1 U9682 ( .A1(n9230), .A2(n8129), .A3(n8128), .ZN(n8130) );
  NAND4_X1 U9683 ( .A1(n9174), .A2(n8131), .A3(n9196), .A4(n8130), .ZN(n8132)
         );
  NOR2_X1 U9684 ( .A1(n9154), .A2(n8132), .ZN(n8133) );
  NAND3_X1 U9685 ( .A1(n9117), .A2(n9137), .A3(n8133), .ZN(n8134) );
  NOR2_X1 U9686 ( .A1(n8311), .A2(n8134), .ZN(n8135) );
  NAND3_X1 U9687 ( .A1(n9073), .A2(n9106), .A3(n8135), .ZN(n8136) );
  NOR2_X1 U9688 ( .A1(n8136), .A2(n9058), .ZN(n8137) );
  NAND4_X1 U9689 ( .A1(n9007), .A2(n9027), .A3(n8137), .A4(n9046), .ZN(n8138)
         );
  NOR4_X1 U9690 ( .A1(n8239), .A2(n8202), .A3(n8322), .A4(n8138), .ZN(n8139)
         );
  AOI21_X1 U9691 ( .B1(n8241), .B2(n8139), .A(n8206), .ZN(n8200) );
  INV_X1 U9692 ( .A(n8140), .ZN(n8199) );
  INV_X1 U9693 ( .A(n8316), .ZN(n8141) );
  AND2_X1 U9694 ( .A1(n8318), .A2(n8141), .ZN(n8142) );
  NOR2_X1 U9695 ( .A1(n8143), .A2(n8142), .ZN(n8231) );
  INV_X1 U9696 ( .A(n9133), .ZN(n8145) );
  OR2_X1 U9697 ( .A1(n8146), .A2(n8145), .ZN(n8226) );
  AND2_X1 U9698 ( .A1(n8147), .A2(n9211), .ZN(n8298) );
  NAND4_X1 U9699 ( .A1(n8165), .A2(n8164), .A3(n8149), .A4(n8148), .ZN(n8150)
         );
  NOR2_X1 U9700 ( .A1(n8170), .A2(n8150), .ZN(n8151) );
  AND2_X1 U9701 ( .A1(n8298), .A2(n8151), .ZN(n8152) );
  NAND2_X1 U9702 ( .A1(n8301), .A2(n8152), .ZN(n8223) );
  AND2_X1 U9703 ( .A1(n8153), .A2(n8159), .ZN(n8217) );
  NAND4_X1 U9704 ( .A1(n8154), .A2(n8217), .A3(n8215), .A4(n8209), .ZN(n8162)
         );
  NAND2_X1 U9705 ( .A1(n8219), .A2(n8213), .ZN(n8160) );
  NAND3_X1 U9706 ( .A1(n8157), .A2(n8156), .A3(n8155), .ZN(n8158) );
  NAND3_X1 U9707 ( .A1(n8160), .A2(n8159), .A3(n8158), .ZN(n8161) );
  NAND2_X1 U9708 ( .A1(n8162), .A2(n8161), .ZN(n8175) );
  INV_X1 U9709 ( .A(n8163), .ZN(n8166) );
  OAI211_X1 U9710 ( .C1(n8167), .C2(n8166), .A(n8165), .B(n8164), .ZN(n8168)
         );
  AND2_X1 U9711 ( .A1(n4358), .A2(n8168), .ZN(n8171) );
  OAI211_X1 U9712 ( .C1(n8171), .C2(n8170), .A(n8297), .B(n8169), .ZN(n8172)
         );
  NAND2_X1 U9713 ( .A1(n8298), .A2(n8172), .ZN(n8173) );
  NAND2_X1 U9714 ( .A1(n8173), .A2(n8299), .ZN(n8174) );
  NAND2_X1 U9715 ( .A1(n8301), .A2(n8174), .ZN(n8221) );
  OAI21_X1 U9716 ( .B1(n8223), .B2(n8175), .A(n8221), .ZN(n8176) );
  INV_X1 U9717 ( .A(n8176), .ZN(n8177) );
  NOR2_X1 U9718 ( .A1(n8226), .A2(n8177), .ZN(n8191) );
  INV_X1 U9719 ( .A(n8178), .ZN(n8181) );
  INV_X1 U9720 ( .A(n8179), .ZN(n8180) );
  OAI21_X1 U9721 ( .B1(n8182), .B2(n8181), .A(n8180), .ZN(n8185) );
  INV_X1 U9722 ( .A(n8183), .ZN(n8184) );
  OAI21_X1 U9723 ( .B1(n8186), .B2(n8185), .A(n8184), .ZN(n8187) );
  INV_X1 U9724 ( .A(n8187), .ZN(n8188) );
  OR2_X1 U9725 ( .A1(n8189), .A2(n8188), .ZN(n8228) );
  INV_X1 U9726 ( .A(n8190), .ZN(n8227) );
  OAI21_X1 U9727 ( .B1(n8191), .B2(n8228), .A(n8227), .ZN(n8192) );
  NAND3_X1 U9728 ( .A1(n8318), .A2(n8315), .A3(n8192), .ZN(n8193) );
  AND2_X1 U9729 ( .A1(n8231), .A2(n8193), .ZN(n8196) );
  NAND2_X1 U9730 ( .A1(n8194), .A2(n8319), .ZN(n8232) );
  OAI211_X1 U9731 ( .C1(n8196), .C2(n8232), .A(n8195), .B(n8237), .ZN(n8198)
         );
  INV_X1 U9732 ( .A(n8202), .ZN(n8238) );
  INV_X1 U9733 ( .A(n8203), .ZN(n8207) );
  NAND2_X1 U9734 ( .A1(n7040), .A2(n8204), .ZN(n8205) );
  NAND3_X1 U9735 ( .A1(n8207), .A2(n8206), .A3(n8205), .ZN(n8208) );
  NAND2_X1 U9736 ( .A1(n7158), .A2(n8208), .ZN(n8211) );
  OAI211_X1 U9737 ( .C1(n8212), .C2(n8211), .A(n8210), .B(n8209), .ZN(n8214)
         );
  NAND2_X1 U9738 ( .A1(n8214), .A2(n8213), .ZN(n8216) );
  NAND2_X1 U9739 ( .A1(n8216), .A2(n8215), .ZN(n8220) );
  INV_X1 U9740 ( .A(n8217), .ZN(n8218) );
  AOI21_X1 U9741 ( .B1(n8220), .B2(n8219), .A(n8218), .ZN(n8222) );
  OAI21_X1 U9742 ( .B1(n8223), .B2(n8222), .A(n8221), .ZN(n8224) );
  INV_X1 U9743 ( .A(n8224), .ZN(n8225) );
  NOR2_X1 U9744 ( .A1(n8226), .A2(n8225), .ZN(n8229) );
  OAI21_X1 U9745 ( .B1(n8229), .B2(n8228), .A(n8227), .ZN(n8230) );
  AND3_X1 U9746 ( .A1(n9027), .A2(n8315), .A3(n8230), .ZN(n8235) );
  INV_X1 U9747 ( .A(n8231), .ZN(n8234) );
  INV_X1 U9748 ( .A(n8232), .ZN(n8233) );
  OAI21_X1 U9749 ( .B1(n8235), .B2(n8234), .A(n8233), .ZN(n8236) );
  NAND3_X1 U9750 ( .A1(n8238), .A2(n8237), .A3(n8236), .ZN(n8240) );
  AOI21_X1 U9751 ( .B1(n8241), .B2(n8240), .A(n8239), .ZN(n8245) );
  INV_X1 U9752 ( .A(n8242), .ZN(n9644) );
  NAND2_X1 U9753 ( .A1(n8245), .A2(n8243), .ZN(n8244) );
  OAI211_X1 U9754 ( .C1(n8245), .C2(n9644), .A(n8244), .B(n8247), .ZN(n8251)
         );
  INV_X1 U9755 ( .A(n9654), .ZN(n8246) );
  NOR4_X1 U9756 ( .A1(n8246), .A2(n9634), .A3(n9479), .A4(n5718), .ZN(n8250)
         );
  INV_X1 U9757 ( .A(n8247), .ZN(n8248) );
  OAI21_X1 U9758 ( .B1(n5780), .B2(n8248), .A(P1_B_REG_SCAN_IN), .ZN(n8249) );
  INV_X1 U9759 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n8252) );
  NAND3_X1 U9760 ( .A1(n8252), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .ZN(n8256) );
  NAND2_X1 U9761 ( .A1(n7791), .A2(n8253), .ZN(n8255) );
  NAND2_X1 U9762 ( .A1(n8841), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n8254) );
  OAI211_X1 U9763 ( .C1(n5003), .C2(n8256), .A(n8255), .B(n8254), .ZN(P2_U3327) );
  NOR2_X1 U9764 ( .A1(n9328), .A2(n8949), .ZN(n8260) );
  NAND2_X1 U9765 ( .A1(n9328), .A2(n8949), .ZN(n8259) );
  OAI21_X1 U9766 ( .B1(n9229), .B2(n8260), .A(n8259), .ZN(n9202) );
  NAND2_X1 U9767 ( .A1(n9202), .A2(n9213), .ZN(n9187) );
  NAND2_X1 U9768 ( .A1(n9325), .A2(n8948), .ZN(n9186) );
  AND2_X1 U9769 ( .A1(n4378), .A2(n9186), .ZN(n8261) );
  NAND2_X1 U9770 ( .A1(n9187), .A2(n8261), .ZN(n8263) );
  OR2_X1 U9771 ( .A1(n9320), .A2(n9169), .ZN(n8262) );
  NAND2_X1 U9772 ( .A1(n8263), .A2(n8262), .ZN(n9173) );
  INV_X1 U9773 ( .A(n9173), .ZN(n8265) );
  NAND2_X1 U9774 ( .A1(n9313), .A2(n8947), .ZN(n8266) );
  OR2_X1 U9775 ( .A1(n9157), .A2(n9312), .ZN(n8267) );
  AND2_X1 U9776 ( .A1(n9141), .A2(n9123), .ZN(n8269) );
  INV_X1 U9777 ( .A(n9118), .ZN(n8271) );
  NAND2_X1 U9778 ( .A1(n9296), .A2(n9104), .ZN(n8272) );
  OR2_X1 U9779 ( .A1(n9286), .A2(n9295), .ZN(n8273) );
  NAND2_X1 U9780 ( .A1(n9358), .A2(n9289), .ZN(n8274) );
  INV_X1 U9781 ( .A(n8275), .ZN(n8276) );
  NAND2_X1 U9782 ( .A1(n9096), .A2(n9075), .ZN(n9068) );
  AND2_X1 U9783 ( .A1(n8276), .A2(n9068), .ZN(n9055) );
  AND2_X1 U9784 ( .A1(n9055), .A2(n9058), .ZN(n8277) );
  NAND2_X1 U9785 ( .A1(n9054), .A2(n8277), .ZN(n9036) );
  INV_X1 U9786 ( .A(n8278), .ZN(n8282) );
  INV_X1 U9787 ( .A(n9058), .ZN(n8279) );
  OR2_X1 U9788 ( .A1(n9065), .A2(n9076), .ZN(n8280) );
  NAND2_X1 U9789 ( .A1(n9036), .A2(n8283), .ZN(n8285) );
  INV_X1 U9790 ( .A(n9007), .ZN(n8287) );
  OAI21_X1 U9791 ( .B1(n9254), .B2(n8288), .A(n9004), .ZN(n8289) );
  AOI211_X1 U9792 ( .C1(n9248), .C2(n9013), .A(n9236), .B(n8996), .ZN(n9247)
         );
  NAND2_X1 U9793 ( .A1(n9248), .A2(n9622), .ZN(n8293) );
  INV_X1 U9794 ( .A(n8290), .ZN(n8291) );
  NAND3_X1 U9795 ( .A1(n8291), .A2(P1_REG3_REG_28__SCAN_IN), .A3(n9646), .ZN(
        n8292) );
  OAI211_X1 U9796 ( .C1(n9219), .C2(n8294), .A(n8293), .B(n8292), .ZN(n8331)
         );
  NAND2_X1 U9797 ( .A1(n9224), .A2(n8297), .ZN(n9212) );
  NAND2_X1 U9798 ( .A1(n9212), .A2(n8298), .ZN(n8300) );
  NAND2_X1 U9799 ( .A1(n8300), .A2(n8299), .ZN(n9197) );
  NAND2_X1 U9800 ( .A1(n8303), .A2(n8302), .ZN(n8304) );
  NAND2_X1 U9801 ( .A1(n8307), .A2(n8306), .ZN(n9122) );
  INV_X1 U9802 ( .A(n8309), .ZN(n8310) );
  AOI21_X1 U9803 ( .B1(n9103), .B2(n9106), .A(n8310), .ZN(n9091) );
  NAND2_X1 U9804 ( .A1(n9091), .A2(n9090), .ZN(n9089) );
  NAND2_X1 U9805 ( .A1(n9044), .A2(n8315), .ZN(n8317) );
  INV_X1 U9806 ( .A(n8319), .ZN(n8321) );
  XNOR2_X1 U9807 ( .A(n8324), .B(n8323), .ZN(n8329) );
  NAND2_X1 U9808 ( .A1(n9029), .A2(n9615), .ZN(n8327) );
  NOR2_X1 U9809 ( .A1(n9250), .A2(n9620), .ZN(n8330) );
  AOI211_X1 U9810 ( .C1(n9247), .C2(n9629), .A(n8331), .B(n8330), .ZN(n8332)
         );
  XNOR2_X1 U9811 ( .A(n8334), .B(n8333), .ZN(n8342) );
  OAI22_X1 U9812 ( .A1(n8336), .A2(n8403), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8335), .ZN(n8340) );
  INV_X1 U9813 ( .A(n8498), .ZN(n8337) );
  OAI22_X1 U9814 ( .A1(n8338), .A2(n8404), .B1(n8337), .B2(n8411), .ZN(n8339)
         );
  AOI211_X1 U9815 ( .C1(n8719), .C2(n8420), .A(n8340), .B(n8339), .ZN(n8341)
         );
  OAI21_X1 U9816 ( .B1(n8342), .B2(n8422), .A(n8341), .ZN(P2_U3216) );
  XNOR2_X1 U9817 ( .A(n8381), .B(n8380), .ZN(n8348) );
  INV_X1 U9818 ( .A(n8575), .ZN(n8344) );
  OAI22_X1 U9819 ( .A1(n8372), .A2(n9848), .B1(n8363), .B2(n9846), .ZN(n8569)
         );
  AOI22_X1 U9820 ( .A1(n8569), .A2(n8364), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3152), .ZN(n8343) );
  OAI21_X1 U9821 ( .B1(n8344), .B2(n8411), .A(n8343), .ZN(n8345) );
  AOI21_X1 U9822 ( .B1(n8346), .B2(n8420), .A(n8345), .ZN(n8347) );
  OAI21_X1 U9823 ( .B1(n8348), .B2(n8422), .A(n8347), .ZN(P2_U3218) );
  OAI21_X1 U9824 ( .B1(n8351), .B2(n8350), .A(n8349), .ZN(n8353) );
  NAND2_X1 U9825 ( .A1(n8353), .A2(n8352), .ZN(n8359) );
  INV_X1 U9826 ( .A(n8638), .ZN(n8427) );
  NOR2_X1 U9827 ( .A1(n8354), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8461) );
  INV_X1 U9828 ( .A(n8642), .ZN(n8355) );
  OAI22_X1 U9829 ( .A1(n8404), .A2(n8675), .B1(n8411), .B2(n8355), .ZN(n8356)
         );
  AOI211_X1 U9830 ( .C1(n8357), .C2(n8427), .A(n8461), .B(n8356), .ZN(n8358)
         );
  OAI211_X1 U9831 ( .C1(n4547), .C2(n8360), .A(n8359), .B(n8358), .ZN(P2_U3221) );
  XNOR2_X1 U9832 ( .A(n8362), .B(n8361), .ZN(n8369) );
  INV_X1 U9833 ( .A(n8607), .ZN(n8366) );
  OAI22_X1 U9834 ( .A1(n8363), .A2(n9848), .B1(n8638), .B2(n9846), .ZN(n8605)
         );
  AOI22_X1 U9835 ( .A1(n8364), .A2(n8605), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3152), .ZN(n8365) );
  OAI21_X1 U9836 ( .B1(n8366), .B2(n8411), .A(n8365), .ZN(n8367) );
  AOI21_X1 U9837 ( .B1(n8751), .B2(n8420), .A(n8367), .ZN(n8368) );
  OAI21_X1 U9838 ( .B1(n8369), .B2(n8422), .A(n8368), .ZN(P2_U3225) );
  XNOR2_X1 U9839 ( .A(n8371), .B(n8370), .ZN(n8378) );
  NOR2_X1 U9840 ( .A1(n8372), .A2(n9846), .ZN(n8373) );
  AOI21_X1 U9841 ( .B1(n8504), .B2(n8547), .A(n8373), .ZN(n8534) );
  OAI22_X1 U9842 ( .A1(n8534), .A2(n8417), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10142), .ZN(n8374) );
  AOI21_X1 U9843 ( .B1(n8537), .B2(n8375), .A(n8374), .ZN(n8377) );
  NAND2_X1 U9844 ( .A1(n8731), .A2(n8420), .ZN(n8376) );
  OAI211_X1 U9845 ( .C1(n8378), .C2(n8422), .A(n8377), .B(n8376), .ZN(P2_U3227) );
  AOI21_X1 U9846 ( .B1(n8381), .B2(n8380), .A(n8379), .ZN(n8385) );
  XNOR2_X1 U9847 ( .A(n8383), .B(n8382), .ZN(n8384) );
  XNOR2_X1 U9848 ( .A(n8385), .B(n8384), .ZN(n8390) );
  OAI22_X1 U9849 ( .A1(n8413), .A2(n8403), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8386), .ZN(n8388) );
  OAI22_X1 U9850 ( .A1(n8404), .A2(n8591), .B1(n8411), .B2(n8557), .ZN(n8387)
         );
  AOI211_X1 U9851 ( .C1(n8735), .C2(n8420), .A(n8388), .B(n8387), .ZN(n8389)
         );
  OAI21_X1 U9852 ( .B1(n8390), .B2(n8422), .A(n8389), .ZN(P2_U3231) );
  XNOR2_X1 U9853 ( .A(n8392), .B(n8391), .ZN(n8398) );
  OAI22_X1 U9854 ( .A1(n8403), .A2(n8617), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8393), .ZN(n8396) );
  OAI22_X1 U9855 ( .A1(n8404), .A2(n8655), .B1(n8411), .B2(n8394), .ZN(n8395)
         );
  AOI211_X1 U9856 ( .C1(n8757), .C2(n8420), .A(n8396), .B(n8395), .ZN(n8397)
         );
  OAI21_X1 U9857 ( .B1(n8398), .B2(n8422), .A(n8397), .ZN(P2_U3235) );
  AOI21_X1 U9858 ( .B1(n8401), .B2(n8400), .A(n8399), .ZN(n8408) );
  OAI22_X1 U9859 ( .A1(n8403), .A2(n8591), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8402), .ZN(n8406) );
  OAI22_X1 U9860 ( .A1(n8404), .A2(n8617), .B1(n8411), .B2(n8583), .ZN(n8405)
         );
  AOI211_X1 U9861 ( .C1(n8745), .C2(n8420), .A(n8406), .B(n8405), .ZN(n8407)
         );
  OAI21_X1 U9862 ( .B1(n8408), .B2(n8422), .A(n8407), .ZN(P2_U3237) );
  XNOR2_X1 U9863 ( .A(n8410), .B(n8409), .ZN(n8423) );
  NOR2_X1 U9864 ( .A1(n8521), .A2(n8411), .ZN(n8419) );
  OR2_X1 U9865 ( .A1(n8412), .A2(n9848), .ZN(n8415) );
  OR2_X1 U9866 ( .A1(n8413), .A2(n9846), .ZN(n8414) );
  AND2_X1 U9867 ( .A1(n8415), .A2(n8414), .ZN(n8513) );
  OAI22_X1 U9868 ( .A1(n8513), .A2(n8417), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8416), .ZN(n8418) );
  AOI211_X1 U9869 ( .C1(n8519), .C2(n8420), .A(n8419), .B(n8418), .ZN(n8421)
         );
  OAI21_X1 U9870 ( .B1(n8423), .B2(n8422), .A(n8421), .ZN(P2_U3242) );
  MUX2_X1 U9871 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8424), .S(P2_U3966), .Z(
        P2_U3582) );
  MUX2_X1 U9872 ( .A(n8503), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8444), .Z(
        P2_U3580) );
  MUX2_X1 U9873 ( .A(n8504), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8444), .Z(
        P2_U3578) );
  MUX2_X1 U9874 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8548), .S(P2_U3966), .Z(
        P2_U3577) );
  MUX2_X1 U9875 ( .A(n8425), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8444), .Z(
        P2_U3576) );
  MUX2_X1 U9876 ( .A(n8546), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8444), .Z(
        P2_U3575) );
  MUX2_X1 U9877 ( .A(n8426), .B(P2_DATAO_REG_21__SCAN_IN), .S(n8444), .Z(
        P2_U3573) );
  MUX2_X1 U9878 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8427), .S(P2_U3966), .Z(
        P2_U3572) );
  MUX2_X1 U9879 ( .A(n8428), .B(P2_DATAO_REG_19__SCAN_IN), .S(n8444), .Z(
        P2_U3571) );
  MUX2_X1 U9880 ( .A(n8429), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8444), .Z(
        P2_U3570) );
  MUX2_X1 U9881 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8430), .S(P2_U3966), .Z(
        P2_U3569) );
  MUX2_X1 U9882 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8431), .S(P2_U3966), .Z(
        P2_U3568) );
  MUX2_X1 U9883 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8432), .S(P2_U3966), .Z(
        P2_U3567) );
  MUX2_X1 U9884 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8433), .S(P2_U3966), .Z(
        P2_U3566) );
  MUX2_X1 U9885 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n8434), .S(P2_U3966), .Z(
        P2_U3565) );
  MUX2_X1 U9886 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n8435), .S(P2_U3966), .Z(
        P2_U3564) );
  MUX2_X1 U9887 ( .A(n8436), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8444), .Z(
        P2_U3563) );
  MUX2_X1 U9888 ( .A(n4655), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8444), .Z(
        P2_U3562) );
  MUX2_X1 U9889 ( .A(n8437), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8444), .Z(
        P2_U3561) );
  MUX2_X1 U9890 ( .A(n8438), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8444), .Z(
        P2_U3560) );
  MUX2_X1 U9891 ( .A(n8439), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8444), .Z(
        P2_U3559) );
  MUX2_X1 U9892 ( .A(n8440), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8444), .Z(
        P2_U3558) );
  MUX2_X1 U9893 ( .A(n8441), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8444), .Z(
        P2_U3557) );
  MUX2_X1 U9894 ( .A(n8442), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8444), .Z(
        P2_U3556) );
  MUX2_X1 U9895 ( .A(n8443), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8444), .Z(
        P2_U3555) );
  MUX2_X1 U9896 ( .A(n6687), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8444), .Z(
        P2_U3554) );
  MUX2_X1 U9897 ( .A(n6673), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8444), .Z(
        P2_U3553) );
  MUX2_X1 U9898 ( .A(n6701), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8444), .Z(
        P2_U3552) );
  NAND2_X1 U9899 ( .A1(n8446), .A2(n8445), .ZN(n8447) );
  NAND2_X1 U9900 ( .A1(n8448), .A2(n8447), .ZN(n8449) );
  XOR2_X1 U9901 ( .A(n8449), .B(P2_REG2_REG_19__SCAN_IN), .Z(n8458) );
  AOI21_X1 U9902 ( .B1(n8452), .B2(n8451), .A(n8450), .ZN(n8453) );
  XOR2_X1 U9903 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8453), .Z(n8457) );
  INV_X1 U9904 ( .A(n8457), .ZN(n8454) );
  NAND2_X1 U9905 ( .A1(n8454), .A2(n9786), .ZN(n8455) );
  OAI211_X1 U9906 ( .C1(n8458), .C2(n9736), .A(n8455), .B(n9734), .ZN(n8456)
         );
  INV_X1 U9907 ( .A(n8456), .ZN(n8460) );
  AOI22_X1 U9908 ( .A1(n8458), .A2(n9783), .B1(n8457), .B2(n9786), .ZN(n8459)
         );
  MUX2_X1 U9909 ( .A(n8460), .B(n8459), .S(n8682), .Z(n8463) );
  INV_X1 U9910 ( .A(n8461), .ZN(n8462) );
  OAI211_X1 U9911 ( .C1(n4750), .C2(n8464), .A(n8463), .B(n8462), .ZN(P2_U3264) );
  OAI211_X1 U9912 ( .C1(n8810), .C2(n8466), .A(n7321), .B(n8465), .ZN(n8716)
         );
  NOR2_X1 U9913 ( .A1(n8810), .A2(n8693), .ZN(n8467) );
  AOI211_X1 U9914 ( .C1(n9866), .C2(P2_REG2_REG_30__SCAN_IN), .A(n8468), .B(
        n8467), .ZN(n8469) );
  OAI21_X1 U9915 ( .B1(n9832), .B2(n8716), .A(n8469), .ZN(P2_U3266) );
  NAND2_X1 U9916 ( .A1(n8470), .A2(n9834), .ZN(n8478) );
  INV_X1 U9917 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n8471) );
  OAI22_X1 U9918 ( .A1(n8472), .A2(n8556), .B1(n8471), .B2(n8579), .ZN(n8475)
         );
  NOR2_X1 U9919 ( .A1(n8473), .A2(n9832), .ZN(n8474) );
  AOI211_X1 U9920 ( .C1(n9856), .C2(n8476), .A(n8475), .B(n8474), .ZN(n8477)
         );
  OAI211_X1 U9921 ( .C1(n8479), .C2(n9855), .A(n8478), .B(n8477), .ZN(P2_U3267) );
  INV_X1 U9922 ( .A(n8480), .ZN(n8490) );
  NAND2_X1 U9923 ( .A1(n8481), .A2(n9834), .ZN(n8489) );
  NOR2_X1 U9924 ( .A1(n8482), .A2(n8693), .ZN(n8486) );
  OAI22_X1 U9925 ( .A1(n8484), .A2(n8556), .B1(n8483), .B2(n8579), .ZN(n8485)
         );
  AOI211_X1 U9926 ( .C1(n8487), .C2(n9862), .A(n8486), .B(n8485), .ZN(n8488)
         );
  OAI211_X1 U9927 ( .C1(n8490), .C2(n9855), .A(n8489), .B(n8488), .ZN(P2_U3268) );
  NAND2_X1 U9928 ( .A1(n8516), .A2(n8515), .ZN(n8492) );
  NAND2_X1 U9929 ( .A1(n8492), .A2(n8491), .ZN(n8494) );
  XNOR2_X1 U9930 ( .A(n8494), .B(n8493), .ZN(n8723) );
  INV_X1 U9931 ( .A(n8517), .ZN(n8497) );
  INV_X1 U9932 ( .A(n8495), .ZN(n8496) );
  AOI21_X1 U9933 ( .B1(n8719), .B2(n8497), .A(n8496), .ZN(n8720) );
  AOI22_X1 U9934 ( .A1(n8498), .A2(n9854), .B1(P2_REG2_REG_27__SCAN_IN), .B2(
        n9855), .ZN(n8499) );
  OAI21_X1 U9935 ( .B1(n8500), .B2(n8693), .A(n8499), .ZN(n8507) );
  XNOR2_X1 U9936 ( .A(n8502), .B(n8501), .ZN(n8505) );
  AOI222_X1 U9937 ( .A1(n9818), .A2(n8505), .B1(n8504), .B2(n8545), .C1(n8503), 
        .C2(n8547), .ZN(n8722) );
  NOR2_X1 U9938 ( .A1(n8722), .A2(n9866), .ZN(n8506) );
  AOI211_X1 U9939 ( .C1(n8720), .C2(n8707), .A(n8507), .B(n8506), .ZN(n8508)
         );
  OAI21_X1 U9940 ( .B1(n8723), .B2(n8709), .A(n8508), .ZN(P2_U3269) );
  INV_X1 U9941 ( .A(n8509), .ZN(n8533) );
  NAND2_X1 U9942 ( .A1(n8533), .A2(n8510), .ZN(n8512) );
  AOI21_X1 U9943 ( .B1(n8515), .B2(n8512), .A(n8511), .ZN(n8514) );
  OAI21_X1 U9944 ( .B1(n8514), .B2(n9843), .A(n8513), .ZN(n8724) );
  INV_X1 U9945 ( .A(n8724), .ZN(n8526) );
  XNOR2_X1 U9946 ( .A(n8516), .B(n8515), .ZN(n8726) );
  NAND2_X1 U9947 ( .A1(n8726), .A2(n9834), .ZN(n8525) );
  INV_X1 U9948 ( .A(n8536), .ZN(n8518) );
  AOI211_X1 U9949 ( .C1(n8519), .C2(n8518), .A(n6682), .B(n8517), .ZN(n8725)
         );
  NOR2_X1 U9950 ( .A1(n8814), .A2(n8693), .ZN(n8523) );
  INV_X1 U9951 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8520) );
  OAI22_X1 U9952 ( .A1(n8521), .A2(n8556), .B1(n8520), .B2(n8579), .ZN(n8522)
         );
  AOI211_X1 U9953 ( .C1(n8725), .C2(n8641), .A(n8523), .B(n8522), .ZN(n8524)
         );
  OAI211_X1 U9954 ( .C1(n9866), .C2(n8526), .A(n8525), .B(n8524), .ZN(P2_U3270) );
  XNOR2_X1 U9955 ( .A(n8528), .B(n8527), .ZN(n8733) );
  AOI22_X1 U9956 ( .A1(n8731), .A2(n9856), .B1(n9866), .B2(
        P2_REG2_REG_25__SCAN_IN), .ZN(n8543) );
  NAND3_X1 U9957 ( .A1(n8531), .A2(n8530), .A3(n8529), .ZN(n8532) );
  NAND3_X1 U9958 ( .A1(n8533), .A2(n9818), .A3(n8532), .ZN(n8535) );
  NAND2_X1 U9959 ( .A1(n8535), .A2(n8534), .ZN(n8729) );
  AOI211_X1 U9960 ( .C1(n8731), .C2(n8553), .A(n6682), .B(n8536), .ZN(n8730)
         );
  INV_X1 U9961 ( .A(n8730), .ZN(n8540) );
  INV_X1 U9962 ( .A(n8537), .ZN(n8538) );
  OAI22_X1 U9963 ( .A1(n8540), .A2(n8539), .B1(n8556), .B2(n8538), .ZN(n8541)
         );
  OAI21_X1 U9964 ( .B1(n8729), .B2(n8541), .A(n8579), .ZN(n8542) );
  OAI211_X1 U9965 ( .C1(n8733), .C2(n8709), .A(n8543), .B(n8542), .ZN(P2_U3271) );
  XNOR2_X1 U9966 ( .A(n8544), .B(n8551), .ZN(n8549) );
  AOI222_X1 U9967 ( .A1(n9818), .A2(n8549), .B1(n8548), .B2(n8547), .C1(n8546), 
        .C2(n8545), .ZN(n8738) );
  OAI21_X1 U9968 ( .B1(n8552), .B2(n8551), .A(n8550), .ZN(n8734) );
  NAND2_X1 U9969 ( .A1(n8734), .A2(n9834), .ZN(n8562) );
  INV_X1 U9970 ( .A(n8553), .ZN(n8554) );
  AOI21_X1 U9971 ( .B1(n8735), .B2(n8572), .A(n8554), .ZN(n8736) );
  INV_X1 U9972 ( .A(n8735), .ZN(n8555) );
  NOR2_X1 U9973 ( .A1(n8555), .A2(n8693), .ZN(n8560) );
  OAI22_X1 U9974 ( .A1(n8579), .A2(n8558), .B1(n8557), .B2(n8556), .ZN(n8559)
         );
  AOI211_X1 U9975 ( .C1(n8736), .C2(n8707), .A(n8560), .B(n8559), .ZN(n8561)
         );
  OAI211_X1 U9976 ( .C1(n9866), .C2(n8738), .A(n8562), .B(n8561), .ZN(P2_U3272) );
  XOR2_X1 U9977 ( .A(n8566), .B(n8563), .Z(n8742) );
  INV_X1 U9978 ( .A(n8742), .ZN(n8581) );
  NAND2_X1 U9979 ( .A1(n8564), .A2(n8565), .ZN(n8567) );
  XNOR2_X1 U9980 ( .A(n8567), .B(n8566), .ZN(n8568) );
  NAND2_X1 U9981 ( .A1(n8568), .A2(n9818), .ZN(n8571) );
  INV_X1 U9982 ( .A(n8569), .ZN(n8570) );
  NAND2_X1 U9983 ( .A1(n8571), .A2(n8570), .ZN(n8740) );
  INV_X1 U9984 ( .A(n8572), .ZN(n8574) );
  AOI21_X1 U9985 ( .B1(n8599), .B2(n8586), .A(n8819), .ZN(n8573) );
  NOR3_X1 U9986 ( .A1(n8574), .A2(n8573), .A3(n6682), .ZN(n8741) );
  NAND2_X1 U9987 ( .A1(n8741), .A2(n9862), .ZN(n8577) );
  AOI22_X1 U9988 ( .A1(n9866), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n8575), .B2(
        n9854), .ZN(n8576) );
  OAI211_X1 U9989 ( .C1(n8819), .C2(n8693), .A(n8577), .B(n8576), .ZN(n8578)
         );
  AOI21_X1 U9990 ( .B1(n8740), .B2(n8579), .A(n8578), .ZN(n8580) );
  OAI21_X1 U9991 ( .B1(n8581), .B2(n8709), .A(n8580), .ZN(P2_U3273) );
  XOR2_X1 U9992 ( .A(n8590), .B(n8582), .Z(n8749) );
  XNOR2_X1 U9993 ( .A(n8599), .B(n8745), .ZN(n8746) );
  INV_X1 U9994 ( .A(n8583), .ZN(n8584) );
  AOI22_X1 U9995 ( .A1(n9866), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8584), .B2(
        n9854), .ZN(n8585) );
  OAI21_X1 U9996 ( .B1(n8586), .B2(n8693), .A(n8585), .ZN(n8595) );
  NAND2_X1 U9997 ( .A1(n8603), .A2(n8587), .ZN(n8589) );
  INV_X1 U9998 ( .A(n8564), .ZN(n8588) );
  AOI211_X1 U9999 ( .C1(n8590), .C2(n8589), .A(n9843), .B(n8588), .ZN(n8593)
         );
  OAI22_X1 U10000 ( .A1(n8591), .A2(n9848), .B1(n8617), .B2(n9846), .ZN(n8592)
         );
  NOR2_X1 U10001 ( .A1(n8593), .A2(n8592), .ZN(n8748) );
  NOR2_X1 U10002 ( .A1(n8748), .A2(n9855), .ZN(n8594) );
  AOI211_X1 U10003 ( .C1(n8746), .C2(n8707), .A(n8595), .B(n8594), .ZN(n8596)
         );
  OAI21_X1 U10004 ( .B1(n8749), .B2(n8709), .A(n8596), .ZN(P2_U3274) );
  XNOR2_X1 U10005 ( .A(n8598), .B(n8597), .ZN(n8754) );
  OAI21_X1 U10006 ( .B1(n8622), .B2(n8602), .A(n7321), .ZN(n8600) );
  NOR2_X1 U10007 ( .A1(n8600), .A2(n8599), .ZN(n8750) );
  INV_X1 U10008 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n8601) );
  OAI22_X1 U10009 ( .A1(n8602), .A2(n8693), .B1(n8579), .B2(n8601), .ZN(n8610)
         );
  OAI21_X1 U10010 ( .B1(n4365), .B2(n8604), .A(n8603), .ZN(n8606) );
  AOI21_X1 U10011 ( .B1(n8606), .B2(n9818), .A(n8605), .ZN(n8753) );
  NAND2_X1 U10012 ( .A1(n8607), .A2(n9854), .ZN(n8608) );
  AOI21_X1 U10013 ( .B1(n8753), .B2(n8608), .A(n9855), .ZN(n8609) );
  AOI211_X1 U10014 ( .C1(n8750), .C2(n9862), .A(n8610), .B(n8609), .ZN(n8611)
         );
  OAI21_X1 U10015 ( .B1(n8754), .B2(n8709), .A(n8611), .ZN(P2_U3275) );
  INV_X1 U10016 ( .A(n8612), .ZN(n8616) );
  AOI21_X1 U10017 ( .B1(n8631), .B2(n8613), .A(n4396), .ZN(n8614) );
  AOI211_X1 U10018 ( .C1(n8616), .C2(n8615), .A(n9843), .B(n8614), .ZN(n8619)
         );
  OAI22_X1 U10019 ( .A1(n8617), .A2(n9848), .B1(n8655), .B2(n9846), .ZN(n8618)
         );
  NOR2_X1 U10020 ( .A1(n8619), .A2(n8618), .ZN(n8760) );
  OR2_X1 U10021 ( .A1(n8621), .A2(n8620), .ZN(n8756) );
  NAND3_X1 U10022 ( .A1(n8756), .A2(n8755), .A3(n9834), .ZN(n8629) );
  AOI21_X1 U10023 ( .B1(n8757), .B2(n8623), .A(n8622), .ZN(n8758) );
  AOI22_X1 U10024 ( .A1(n9866), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8624), .B2(
        n9854), .ZN(n8625) );
  OAI21_X1 U10025 ( .B1(n8626), .B2(n8693), .A(n8625), .ZN(n8627) );
  AOI21_X1 U10026 ( .B1(n8758), .B2(n8707), .A(n8627), .ZN(n8628) );
  OAI211_X1 U10027 ( .C1(n9866), .C2(n8760), .A(n8629), .B(n8628), .ZN(
        P2_U3276) );
  XNOR2_X1 U10028 ( .A(n8630), .B(n8632), .ZN(n8764) );
  INV_X1 U10029 ( .A(n8764), .ZN(n8647) );
  INV_X1 U10030 ( .A(n8631), .ZN(n8636) );
  AOI21_X1 U10031 ( .B1(n8634), .B2(n8633), .A(n8632), .ZN(n8635) );
  NOR2_X1 U10032 ( .A1(n8636), .A2(n8635), .ZN(n8637) );
  OAI222_X1 U10033 ( .A1(n9848), .A2(n8638), .B1(n9846), .B2(n8675), .C1(n9843), .C2(n8637), .ZN(n8762) );
  XNOR2_X1 U10034 ( .A(n8656), .B(n8639), .ZN(n8640) );
  NOR2_X1 U10035 ( .A1(n8640), .A2(n6682), .ZN(n8763) );
  NAND2_X1 U10036 ( .A1(n8763), .A2(n8641), .ZN(n8644) );
  AOI22_X1 U10037 ( .A1(n9866), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n8642), .B2(
        n9854), .ZN(n8643) );
  OAI211_X1 U10038 ( .C1(n4547), .C2(n8693), .A(n8644), .B(n8643), .ZN(n8645)
         );
  AOI21_X1 U10039 ( .B1(n8762), .B2(n8579), .A(n8645), .ZN(n8646) );
  OAI21_X1 U10040 ( .B1(n8647), .B2(n8709), .A(n8646), .ZN(P2_U3277) );
  XNOR2_X1 U10041 ( .A(n8648), .B(n8651), .ZN(n8771) );
  AND2_X1 U10042 ( .A1(n8650), .A2(n8649), .ZN(n8652) );
  XNOR2_X1 U10043 ( .A(n8652), .B(n8651), .ZN(n8653) );
  OAI222_X1 U10044 ( .A1(n9848), .A2(n8655), .B1(n9846), .B2(n8654), .C1(n9843), .C2(n8653), .ZN(n8767) );
  INV_X1 U10045 ( .A(n8666), .ZN(n8658) );
  INV_X1 U10046 ( .A(n8656), .ZN(n8657) );
  AOI211_X1 U10047 ( .C1(n8769), .C2(n8658), .A(n6682), .B(n8657), .ZN(n8768)
         );
  NAND2_X1 U10048 ( .A1(n8768), .A2(n9862), .ZN(n8661) );
  AOI22_X1 U10049 ( .A1(n9866), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8659), .B2(
        n9854), .ZN(n8660) );
  OAI211_X1 U10050 ( .C1(n8662), .C2(n8693), .A(n8661), .B(n8660), .ZN(n8663)
         );
  AOI21_X1 U10051 ( .B1(n8767), .B2(n8579), .A(n8663), .ZN(n8664) );
  OAI21_X1 U10052 ( .B1(n8771), .B2(n8709), .A(n8664), .ZN(P2_U3278) );
  INV_X1 U10053 ( .A(n8665), .ZN(n8667) );
  AOI211_X1 U10054 ( .C1(n8668), .C2(n8667), .A(n6682), .B(n8666), .ZN(n8773)
         );
  NAND2_X1 U10055 ( .A1(n8670), .A2(n8669), .ZN(n8672) );
  XNOR2_X1 U10056 ( .A(n8672), .B(n8671), .ZN(n8673) );
  OAI222_X1 U10057 ( .A1(n9848), .A2(n8675), .B1(n9846), .B2(n8674), .C1(n9843), .C2(n8673), .ZN(n8772) );
  OAI21_X1 U10058 ( .B1(n8678), .B2(n8677), .A(n8676), .ZN(n8774) );
  INV_X1 U10059 ( .A(n8774), .ZN(n8680) );
  NOR2_X1 U10060 ( .A1(n8680), .A2(n8679), .ZN(n8681) );
  AOI211_X1 U10061 ( .C1(n8773), .C2(n8682), .A(n8772), .B(n8681), .ZN(n8687)
         );
  AOI22_X1 U10062 ( .A1(n9866), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n8683), .B2(
        n9854), .ZN(n8684) );
  OAI21_X1 U10063 ( .B1(n8830), .B2(n8693), .A(n8684), .ZN(n8685) );
  AOI21_X1 U10064 ( .B1(n8774), .B2(n9863), .A(n8685), .ZN(n8686) );
  OAI21_X1 U10065 ( .B1(n8687), .B2(n9855), .A(n8686), .ZN(P2_U3279) );
  XNOR2_X1 U10066 ( .A(n8688), .B(n8699), .ZN(n8790) );
  AOI21_X1 U10067 ( .B1(n8786), .B2(n8690), .A(n5436), .ZN(n8787) );
  AOI22_X1 U10068 ( .A1(n9866), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n8691), .B2(
        n9854), .ZN(n8692) );
  OAI21_X1 U10069 ( .B1(n8694), .B2(n8693), .A(n8692), .ZN(n8706) );
  AND2_X1 U10070 ( .A1(n8696), .A2(n8695), .ZN(n8704) );
  INV_X1 U10071 ( .A(n8697), .ZN(n8698) );
  NOR2_X1 U10072 ( .A1(n8699), .A2(n8698), .ZN(n8700) );
  AOI21_X1 U10073 ( .B1(n8701), .B2(n8700), .A(n9843), .ZN(n8703) );
  AOI21_X1 U10074 ( .B1(n8704), .B2(n8703), .A(n8702), .ZN(n8789) );
  NOR2_X1 U10075 ( .A1(n8789), .A2(n9866), .ZN(n8705) );
  AOI211_X1 U10076 ( .C1(n8787), .C2(n8707), .A(n8706), .B(n8705), .ZN(n8708)
         );
  OAI21_X1 U10077 ( .B1(n8709), .B2(n8790), .A(n8708), .ZN(P2_U3281) );
  INV_X1 U10078 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n8713) );
  MUX2_X1 U10079 ( .A(n8713), .B(n8804), .S(n9959), .Z(n8714) );
  OAI21_X1 U10080 ( .B1(n8806), .B2(n8777), .A(n8714), .ZN(P2_U3551) );
  INV_X1 U10081 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n8717) );
  MUX2_X1 U10082 ( .A(n8717), .B(n8807), .S(n9959), .Z(n8718) );
  OAI21_X1 U10083 ( .B1(n8810), .B2(n8777), .A(n8718), .ZN(P2_U3550) );
  AOI22_X1 U10084 ( .A1(n8720), .A2(n7321), .B1(n9927), .B2(n8719), .ZN(n8721)
         );
  OAI211_X1 U10085 ( .C1(n8723), .C2(n9932), .A(n8722), .B(n8721), .ZN(n8811)
         );
  MUX2_X1 U10086 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n8811), .S(n9959), .Z(
        P2_U3547) );
  INV_X1 U10087 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8727) );
  AOI211_X1 U10088 ( .C1(n8726), .C2(n9941), .A(n8725), .B(n8724), .ZN(n8812)
         );
  MUX2_X1 U10089 ( .A(n8727), .B(n8812), .S(n9959), .Z(n8728) );
  OAI21_X1 U10090 ( .B1(n8814), .B2(n8777), .A(n8728), .ZN(P2_U3546) );
  AOI211_X1 U10091 ( .C1(n9927), .C2(n8731), .A(n8730), .B(n8729), .ZN(n8732)
         );
  OAI21_X1 U10092 ( .B1(n8733), .B2(n9932), .A(n8732), .ZN(n8815) );
  MUX2_X1 U10093 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n8815), .S(n9959), .Z(
        P2_U3545) );
  INV_X1 U10094 ( .A(n8734), .ZN(n8739) );
  AOI22_X1 U10095 ( .A1(n8736), .A2(n7321), .B1(n9927), .B2(n8735), .ZN(n8737)
         );
  OAI211_X1 U10096 ( .C1(n8739), .C2(n9932), .A(n8738), .B(n8737), .ZN(n8816)
         );
  MUX2_X1 U10097 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8816), .S(n9959), .Z(
        P2_U3544) );
  INV_X1 U10098 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n8743) );
  AOI211_X1 U10099 ( .C1(n8742), .C2(n9941), .A(n8741), .B(n8740), .ZN(n8817)
         );
  MUX2_X1 U10100 ( .A(n8743), .B(n8817), .S(n9959), .Z(n8744) );
  OAI21_X1 U10101 ( .B1(n8819), .B2(n8777), .A(n8744), .ZN(P2_U3543) );
  AOI22_X1 U10102 ( .A1(n8746), .A2(n7321), .B1(n9927), .B2(n8745), .ZN(n8747)
         );
  OAI211_X1 U10103 ( .C1(n8749), .C2(n9932), .A(n8748), .B(n8747), .ZN(n8820)
         );
  MUX2_X1 U10104 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n8820), .S(n9959), .Z(
        P2_U3542) );
  AOI21_X1 U10105 ( .B1(n9927), .B2(n8751), .A(n8750), .ZN(n8752) );
  OAI211_X1 U10106 ( .C1(n8754), .C2(n9932), .A(n8753), .B(n8752), .ZN(n8821)
         );
  MUX2_X1 U10107 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n8821), .S(n9959), .Z(
        P2_U3541) );
  NAND3_X1 U10108 ( .A1(n8756), .A2(n8755), .A3(n9941), .ZN(n8761) );
  AOI22_X1 U10109 ( .A1(n8758), .A2(n7321), .B1(n9927), .B2(n8757), .ZN(n8759)
         );
  NAND3_X1 U10110 ( .A1(n8761), .A2(n8760), .A3(n8759), .ZN(n8822) );
  MUX2_X1 U10111 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n8822), .S(n9959), .Z(
        P2_U3540) );
  INV_X1 U10112 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8765) );
  AOI211_X1 U10113 ( .C1(n8764), .C2(n9941), .A(n8763), .B(n8762), .ZN(n8823)
         );
  MUX2_X1 U10114 ( .A(n8765), .B(n8823), .S(n9959), .Z(n8766) );
  OAI21_X1 U10115 ( .B1(n4547), .B2(n8777), .A(n8766), .ZN(P2_U3539) );
  AOI211_X1 U10116 ( .C1(n9927), .C2(n8769), .A(n8768), .B(n8767), .ZN(n8770)
         );
  OAI21_X1 U10117 ( .B1(n9932), .B2(n8771), .A(n8770), .ZN(n8826) );
  MUX2_X1 U10118 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n8826), .S(n9959), .Z(
        P2_U3538) );
  AOI211_X1 U10119 ( .C1(n8774), .C2(n9941), .A(n8773), .B(n8772), .ZN(n8827)
         );
  MUX2_X1 U10120 ( .A(n8775), .B(n8827), .S(n9959), .Z(n8776) );
  OAI21_X1 U10121 ( .B1(n8830), .B2(n8777), .A(n8776), .ZN(P2_U3537) );
  INV_X1 U10122 ( .A(n8777), .ZN(n8784) );
  OR2_X1 U10123 ( .A1(n8778), .A2(n9932), .ZN(n8782) );
  NOR2_X1 U10124 ( .A1(n8780), .A2(n8779), .ZN(n8781) );
  NAND2_X1 U10125 ( .A1(n8782), .A2(n8781), .ZN(n8832) );
  MUX2_X1 U10126 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n8832), .S(n9959), .Z(n8783) );
  AOI21_X1 U10127 ( .B1(n8784), .B2(n8834), .A(n8783), .ZN(n8785) );
  INV_X1 U10128 ( .A(n8785), .ZN(P2_U3536) );
  AOI22_X1 U10129 ( .A1(n8787), .A2(n7321), .B1(n9927), .B2(n8786), .ZN(n8788)
         );
  OAI211_X1 U10130 ( .C1(n8790), .C2(n9932), .A(n8789), .B(n8788), .ZN(n8837)
         );
  MUX2_X1 U10131 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n8837), .S(n9959), .Z(
        P2_U3535) );
  AOI22_X1 U10132 ( .A1(n8792), .A2(n7321), .B1(n9927), .B2(n8791), .ZN(n8793)
         );
  OAI211_X1 U10133 ( .C1(n8795), .C2(n9932), .A(n8794), .B(n8793), .ZN(n8838)
         );
  MUX2_X1 U10134 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n8838), .S(n9959), .Z(
        P2_U3534) );
  INV_X1 U10135 ( .A(n8796), .ZN(n8797) );
  OAI22_X1 U10136 ( .A1(n8798), .A2(n6682), .B1(n8797), .B2(n9937), .ZN(n8799)
         );
  AOI21_X1 U10137 ( .B1(n8800), .B2(n9920), .A(n8799), .ZN(n8801) );
  NAND2_X1 U10138 ( .A1(n8802), .A2(n8801), .ZN(n8839) );
  MUX2_X1 U10139 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n8839), .S(n9959), .Z(
        P2_U3533) );
  INV_X1 U10140 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n8803) );
  MUX2_X1 U10141 ( .A(n8804), .B(n8803), .S(n9942), .Z(n8805) );
  OAI21_X1 U10142 ( .B1(n8806), .B2(n8831), .A(n8805), .ZN(P2_U3519) );
  INV_X1 U10143 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n8808) );
  MUX2_X1 U10144 ( .A(n8808), .B(n8807), .S(n9944), .Z(n8809) );
  OAI21_X1 U10145 ( .B1(n8810), .B2(n8831), .A(n8809), .ZN(P2_U3518) );
  MUX2_X1 U10146 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n8811), .S(n9944), .Z(
        P2_U3515) );
  MUX2_X1 U10147 ( .A(n10077), .B(n8812), .S(n9944), .Z(n8813) );
  OAI21_X1 U10148 ( .B1(n8814), .B2(n8831), .A(n8813), .ZN(P2_U3514) );
  MUX2_X1 U10149 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n8815), .S(n9944), .Z(
        P2_U3513) );
  MUX2_X1 U10150 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n8816), .S(n9944), .Z(
        P2_U3512) );
  MUX2_X1 U10151 ( .A(n10075), .B(n8817), .S(n9944), .Z(n8818) );
  OAI21_X1 U10152 ( .B1(n8819), .B2(n8831), .A(n8818), .ZN(P2_U3511) );
  MUX2_X1 U10153 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n8820), .S(n9944), .Z(
        P2_U3510) );
  MUX2_X1 U10154 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n8821), .S(n9944), .Z(
        P2_U3509) );
  MUX2_X1 U10155 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n8822), .S(n9944), .Z(
        P2_U3508) );
  INV_X1 U10156 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n8824) );
  MUX2_X1 U10157 ( .A(n8824), .B(n8823), .S(n9944), .Z(n8825) );
  OAI21_X1 U10158 ( .B1(n4547), .B2(n8831), .A(n8825), .ZN(P2_U3507) );
  MUX2_X1 U10159 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n8826), .S(n9944), .Z(
        P2_U3505) );
  INV_X1 U10160 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n8828) );
  MUX2_X1 U10161 ( .A(n8828), .B(n8827), .S(n9944), .Z(n8829) );
  OAI21_X1 U10162 ( .B1(n8830), .B2(n8831), .A(n8829), .ZN(P2_U3502) );
  INV_X1 U10163 ( .A(n8831), .ZN(n8835) );
  MUX2_X1 U10164 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n8832), .S(n9944), .Z(n8833) );
  AOI21_X1 U10165 ( .B1(n8835), .B2(n8834), .A(n8833), .ZN(n8836) );
  INV_X1 U10166 ( .A(n8836), .ZN(P2_U3499) );
  MUX2_X1 U10167 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n8837), .S(n9944), .Z(
        P2_U3496) );
  MUX2_X1 U10168 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n8838), .S(n9944), .Z(
        P2_U3493) );
  MUX2_X1 U10169 ( .A(P2_REG0_REG_13__SCAN_IN), .B(n8839), .S(n9944), .Z(
        P2_U3490) );
  INV_X1 U10170 ( .A(n8840), .ZN(n9392) );
  AOI22_X1 U10171 ( .A1(n8842), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n8841), .ZN(n8843) );
  OAI21_X1 U10172 ( .B1(n9392), .B2(n8844), .A(n8843), .ZN(P2_U3328) );
  MUX2_X1 U10173 ( .A(n8845), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  NOR2_X1 U10174 ( .A1(n4332), .A2(n8846), .ZN(n8848) );
  XNOR2_X1 U10175 ( .A(n8848), .B(n8847), .ZN(n8853) );
  AOI22_X1 U10176 ( .A1(n8938), .A2(n9295), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3084), .ZN(n8850) );
  NAND2_X1 U10177 ( .A1(n8907), .A2(n9097), .ZN(n8849) );
  OAI211_X1 U10178 ( .C1(n8877), .C2(n8936), .A(n8850), .B(n8849), .ZN(n8851)
         );
  AOI21_X1 U10179 ( .B1(n9096), .B2(n8942), .A(n8851), .ZN(n8852) );
  OAI21_X1 U10180 ( .B1(n8853), .B2(n8944), .A(n8852), .ZN(P1_U3214) );
  INV_X1 U10181 ( .A(n8916), .ZN(n8854) );
  AOI21_X1 U10182 ( .B1(n8856), .B2(n8855), .A(n8854), .ZN(n8861) );
  NAND2_X1 U10183 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n8989) );
  OAI21_X1 U10184 ( .B1(n8936), .B2(n9153), .A(n8989), .ZN(n8857) );
  AOI21_X1 U10185 ( .B1(n8938), .B2(n8947), .A(n8857), .ZN(n8858) );
  OAI21_X1 U10186 ( .B1(n8940), .B2(n9158), .A(n8858), .ZN(n8859) );
  AOI21_X1 U10187 ( .B1(n9157), .B2(n8942), .A(n8859), .ZN(n8860) );
  OAI21_X1 U10188 ( .B1(n8861), .B2(n8944), .A(n8860), .ZN(P1_U3217) );
  OAI21_X1 U10189 ( .B1(n8864), .B2(n8863), .A(n8862), .ZN(n8865) );
  NAND2_X1 U10190 ( .A1(n8865), .A2(n8901), .ZN(n8870) );
  NOR2_X1 U10191 ( .A1(n8940), .A2(n9126), .ZN(n8868) );
  OAI22_X1 U10192 ( .A1(n8905), .A2(n9153), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8866), .ZN(n8867) );
  AOI211_X1 U10193 ( .C1(n8922), .C2(n9295), .A(n8868), .B(n8867), .ZN(n8869)
         );
  OAI211_X1 U10194 ( .C1(n9125), .C2(n8910), .A(n8870), .B(n8869), .ZN(
        P1_U3221) );
  OAI21_X1 U10195 ( .B1(n8873), .B2(n8872), .A(n8871), .ZN(n8874) );
  NAND2_X1 U10196 ( .A1(n8874), .A2(n8901), .ZN(n8880) );
  INV_X1 U10197 ( .A(n8875), .ZN(n9060) );
  AOI22_X1 U10198 ( .A1(n9028), .A2(n8922), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3084), .ZN(n8876) );
  OAI21_X1 U10199 ( .B1(n8877), .B2(n8905), .A(n8876), .ZN(n8878) );
  AOI21_X1 U10200 ( .B1(n9060), .B2(n8907), .A(n8878), .ZN(n8879) );
  OAI211_X1 U10201 ( .C1(n9354), .C2(n8910), .A(n8880), .B(n8879), .ZN(
        P1_U3223) );
  INV_X1 U10202 ( .A(n8881), .ZN(n8882) );
  AOI21_X1 U10203 ( .B1(n8884), .B2(n8883), .A(n8882), .ZN(n8889) );
  AND2_X1 U10204 ( .A1(P1_U3084), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9565) );
  NOR2_X1 U10205 ( .A1(n8905), .A2(n9216), .ZN(n8885) );
  AOI211_X1 U10206 ( .C1(n8922), .C2(n9169), .A(n9565), .B(n8885), .ZN(n8886)
         );
  OAI21_X1 U10207 ( .B1(n8940), .B2(n9207), .A(n8886), .ZN(n8887) );
  AOI21_X1 U10208 ( .B1(n9325), .B2(n8942), .A(n8887), .ZN(n8888) );
  OAI21_X1 U10209 ( .B1(n8889), .B2(n8944), .A(n8888), .ZN(P1_U3224) );
  OAI21_X1 U10210 ( .B1(n8892), .B2(n8890), .A(n8891), .ZN(n8893) );
  NAND2_X1 U10211 ( .A1(n8893), .A2(n8901), .ZN(n8897) );
  NOR2_X1 U10212 ( .A1(n8940), .A2(n9192), .ZN(n8895) );
  NAND2_X1 U10213 ( .A1(P1_U3084), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9581) );
  OAI21_X1 U10214 ( .B1(n8936), .B2(n9199), .A(n9581), .ZN(n8894) );
  AOI211_X1 U10215 ( .C1(n8938), .C2(n8948), .A(n8895), .B(n8894), .ZN(n8896)
         );
  OAI211_X1 U10216 ( .C1(n9191), .C2(n8910), .A(n8897), .B(n8896), .ZN(
        P1_U3226) );
  OAI21_X1 U10217 ( .B1(n8900), .B2(n8899), .A(n8898), .ZN(n8902) );
  NAND2_X1 U10218 ( .A1(n8902), .A2(n8901), .ZN(n8909) );
  INV_X1 U10219 ( .A(n8903), .ZN(n9082) );
  AOI22_X1 U10220 ( .A1(n9076), .A2(n8922), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3084), .ZN(n8904) );
  OAI21_X1 U10221 ( .B1(n9289), .B2(n8905), .A(n8904), .ZN(n8906) );
  AOI21_X1 U10222 ( .B1(n9082), .B2(n8907), .A(n8906), .ZN(n8908) );
  OAI211_X1 U10223 ( .C1(n9085), .C2(n8910), .A(n8909), .B(n8908), .ZN(
        P1_U3227) );
  AOI22_X1 U10224 ( .A1(n8922), .A2(n9104), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3084), .ZN(n8912) );
  NAND2_X1 U10225 ( .A1(n8938), .A2(n9312), .ZN(n8911) );
  OAI211_X1 U10226 ( .C1(n8940), .C2(n9142), .A(n8912), .B(n8911), .ZN(n8920)
         );
  INV_X1 U10227 ( .A(n8913), .ZN(n8914) );
  NAND3_X1 U10228 ( .A1(n8916), .A2(n8915), .A3(n8914), .ZN(n8917) );
  AOI21_X1 U10229 ( .B1(n8918), .B2(n8917), .A(n8944), .ZN(n8919) );
  AOI211_X1 U10230 ( .C1(n8942), .C2(n9141), .A(n8920), .B(n8919), .ZN(n8921)
         );
  INV_X1 U10231 ( .A(n8921), .ZN(P1_U3231) );
  AOI22_X1 U10232 ( .A1(n8938), .A2(n9104), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3084), .ZN(n8924) );
  NAND2_X1 U10233 ( .A1(n8922), .A2(n9075), .ZN(n8923) );
  OAI211_X1 U10234 ( .C1(n8940), .C2(n9108), .A(n8924), .B(n8923), .ZN(n8930)
         );
  AOI21_X1 U10235 ( .B1(n8928), .B2(n8925), .A(n8926), .ZN(n8927) );
  AOI211_X1 U10236 ( .C1(n4326), .C2(n8928), .A(n8944), .B(n8927), .ZN(n8929)
         );
  AOI211_X1 U10237 ( .C1(n8942), .C2(n9286), .A(n8930), .B(n8929), .ZN(n8931)
         );
  INV_X1 U10238 ( .A(n8931), .ZN(P1_U3233) );
  NAND2_X1 U10239 ( .A1(n8933), .A2(n8932), .ZN(n8934) );
  XOR2_X1 U10240 ( .A(n8935), .B(n8934), .Z(n8945) );
  NAND2_X1 U10241 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9597) );
  OAI21_X1 U10242 ( .B1(n8936), .B2(n9178), .A(n9597), .ZN(n8937) );
  AOI21_X1 U10243 ( .B1(n8938), .B2(n9169), .A(n8937), .ZN(n8939) );
  OAI21_X1 U10244 ( .B1(n8940), .B2(n9175), .A(n8939), .ZN(n8941) );
  AOI21_X1 U10245 ( .B1(n9313), .B2(n8942), .A(n8941), .ZN(n8943) );
  OAI21_X1 U10246 ( .B1(n8945), .B2(n8944), .A(n8943), .ZN(P1_U3236) );
  MUX2_X1 U10247 ( .A(n8946), .B(P1_DATAO_REG_30__SCAN_IN), .S(n8956), .Z(
        P1_U3585) );
  MUX2_X1 U10248 ( .A(n9010), .B(P1_DATAO_REG_29__SCAN_IN), .S(n8956), .Z(
        P1_U3584) );
  MUX2_X1 U10249 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9029), .S(P1_U4006), .Z(
        P1_U3583) );
  MUX2_X1 U10250 ( .A(n9047), .B(P1_DATAO_REG_27__SCAN_IN), .S(n8956), .Z(
        P1_U3582) );
  MUX2_X1 U10251 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9028), .S(P1_U4006), .Z(
        P1_U3581) );
  MUX2_X1 U10252 ( .A(n9076), .B(P1_DATAO_REG_25__SCAN_IN), .S(n8956), .Z(
        P1_U3580) );
  MUX2_X1 U10253 ( .A(n9092), .B(P1_DATAO_REG_24__SCAN_IN), .S(n8956), .Z(
        P1_U3579) );
  MUX2_X1 U10254 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9075), .S(P1_U4006), .Z(
        P1_U3578) );
  MUX2_X1 U10255 ( .A(n9295), .B(P1_DATAO_REG_22__SCAN_IN), .S(n8956), .Z(
        P1_U3577) );
  MUX2_X1 U10256 ( .A(n9104), .B(P1_DATAO_REG_21__SCAN_IN), .S(n8956), .Z(
        P1_U3576) );
  MUX2_X1 U10257 ( .A(n9123), .B(P1_DATAO_REG_20__SCAN_IN), .S(n8956), .Z(
        P1_U3575) );
  MUX2_X1 U10258 ( .A(n9312), .B(P1_DATAO_REG_19__SCAN_IN), .S(n8956), .Z(
        P1_U3574) );
  MUX2_X1 U10259 ( .A(n8947), .B(P1_DATAO_REG_18__SCAN_IN), .S(n8956), .Z(
        P1_U3573) );
  MUX2_X1 U10260 ( .A(n9169), .B(P1_DATAO_REG_17__SCAN_IN), .S(n8956), .Z(
        P1_U3572) );
  MUX2_X1 U10261 ( .A(n8948), .B(P1_DATAO_REG_16__SCAN_IN), .S(n8956), .Z(
        P1_U3571) );
  MUX2_X1 U10262 ( .A(n8949), .B(P1_DATAO_REG_15__SCAN_IN), .S(n8956), .Z(
        P1_U3570) );
  MUX2_X1 U10263 ( .A(n9225), .B(P1_DATAO_REG_14__SCAN_IN), .S(n8956), .Z(
        P1_U3569) );
  MUX2_X1 U10264 ( .A(n9459), .B(P1_DATAO_REG_13__SCAN_IN), .S(n8956), .Z(
        P1_U3568) );
  MUX2_X1 U10265 ( .A(n8950), .B(P1_DATAO_REG_12__SCAN_IN), .S(n8956), .Z(
        P1_U3567) );
  MUX2_X1 U10266 ( .A(n8951), .B(P1_DATAO_REG_11__SCAN_IN), .S(n8956), .Z(
        P1_U3566) );
  MUX2_X1 U10267 ( .A(n8952), .B(P1_DATAO_REG_10__SCAN_IN), .S(n8956), .Z(
        P1_U3565) );
  MUX2_X1 U10268 ( .A(n8953), .B(P1_DATAO_REG_9__SCAN_IN), .S(n8956), .Z(
        P1_U3564) );
  MUX2_X1 U10269 ( .A(n8954), .B(P1_DATAO_REG_8__SCAN_IN), .S(n8956), .Z(
        P1_U3563) );
  MUX2_X1 U10270 ( .A(n8955), .B(P1_DATAO_REG_7__SCAN_IN), .S(n8956), .Z(
        P1_U3562) );
  MUX2_X1 U10271 ( .A(n9687), .B(P1_DATAO_REG_6__SCAN_IN), .S(n8956), .Z(
        P1_U3561) );
  MUX2_X1 U10272 ( .A(n9614), .B(P1_DATAO_REG_5__SCAN_IN), .S(n8956), .Z(
        P1_U3560) );
  MUX2_X1 U10273 ( .A(n9668), .B(P1_DATAO_REG_4__SCAN_IN), .S(n8956), .Z(
        P1_U3559) );
  MUX2_X1 U10274 ( .A(n6792), .B(P1_DATAO_REG_3__SCAN_IN), .S(n8956), .Z(
        P1_U3558) );
  MUX2_X1 U10275 ( .A(n8957), .B(P1_DATAO_REG_2__SCAN_IN), .S(n8956), .Z(
        P1_U3557) );
  MUX2_X1 U10276 ( .A(n7040), .B(P1_DATAO_REG_1__SCAN_IN), .S(n8956), .Z(
        P1_U3556) );
  MUX2_X1 U10277 ( .A(n6638), .B(P1_DATAO_REG_0__SCAN_IN), .S(n8956), .Z(
        P1_U3555) );
  XNOR2_X1 U10278 ( .A(n8979), .B(P1_REG1_REG_18__SCAN_IN), .ZN(n9604) );
  INV_X1 U10279 ( .A(n8975), .ZN(n9583) );
  XNOR2_X1 U10280 ( .A(n9583), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n9588) );
  INV_X1 U10281 ( .A(n9566), .ZN(n8962) );
  INV_X1 U10282 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n8961) );
  XOR2_X1 U10283 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9566), .Z(n9569) );
  AOI21_X1 U10284 ( .B1(n8966), .B2(n6001), .A(n8958), .ZN(n8959) );
  NAND2_X1 U10285 ( .A1(n9555), .A2(n8959), .ZN(n8960) );
  XNOR2_X1 U10286 ( .A(n8959), .B(n8970), .ZN(n9557) );
  NAND2_X1 U10287 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n9557), .ZN(n9556) );
  NAND2_X1 U10288 ( .A1(n8960), .A2(n9556), .ZN(n9570) );
  NAND2_X1 U10289 ( .A1(n9569), .A2(n9570), .ZN(n9568) );
  OAI21_X1 U10290 ( .B1(n8962), .B2(n8961), .A(n9568), .ZN(n9587) );
  NAND2_X1 U10291 ( .A1(n9588), .A2(n9587), .ZN(n9586) );
  OAI21_X1 U10292 ( .B1(n9583), .B2(n8963), .A(n9586), .ZN(n9603) );
  NOR2_X1 U10293 ( .A1(n9604), .A2(n9603), .ZN(n9602) );
  AOI21_X1 U10294 ( .B1(n9600), .B2(n8964), .A(n9602), .ZN(n8965) );
  XOR2_X1 U10295 ( .A(n8965), .B(P1_REG1_REG_19__SCAN_IN), .Z(n8982) );
  NAND2_X1 U10296 ( .A1(n8967), .A2(n8966), .ZN(n8969) );
  NOR2_X1 U10297 ( .A1(n8970), .A2(n8971), .ZN(n8972) );
  INV_X1 U10298 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9551) );
  NAND2_X1 U10299 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n9566), .ZN(n8973) );
  OAI21_X1 U10300 ( .B1(n9566), .B2(P1_REG2_REG_16__SCAN_IN), .A(n8973), .ZN(
        n9562) );
  NOR2_X1 U10301 ( .A1(n9563), .A2(n9562), .ZN(n9561) );
  AOI21_X1 U10302 ( .B1(n9566), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9561), .ZN(
        n9574) );
  NAND2_X1 U10303 ( .A1(P1_REG2_REG_17__SCAN_IN), .A2(n8975), .ZN(n8974) );
  OAI21_X1 U10304 ( .B1(n8975), .B2(P1_REG2_REG_17__SCAN_IN), .A(n8974), .ZN(
        n9575) );
  NOR2_X1 U10305 ( .A1(n9574), .A2(n9575), .ZN(n9576) );
  OR2_X1 U10306 ( .A1(n8979), .A2(n8976), .ZN(n8978) );
  NAND2_X1 U10307 ( .A1(n8979), .A2(n8976), .ZN(n8977) );
  AND2_X1 U10308 ( .A1(n8978), .A2(n8977), .ZN(n9594) );
  NAND2_X1 U10309 ( .A1(n8984), .A2(n8980), .ZN(n8981) );
  OAI211_X1 U10310 ( .C1(n8982), .C2(n9605), .A(n8981), .B(n9599), .ZN(n8987)
         );
  INV_X1 U10311 ( .A(n8982), .ZN(n8983) );
  OAI22_X1 U10312 ( .A1(n8984), .A2(n9580), .B1(n8983), .B2(n9605), .ZN(n8986)
         );
  MUX2_X1 U10313 ( .A(n8987), .B(n8986), .S(n8985), .Z(n8988) );
  INV_X1 U10314 ( .A(n8988), .ZN(n8990) );
  OAI211_X1 U10315 ( .C1(n9394), .C2(n9609), .A(n8990), .B(n8989), .ZN(
        P1_U3260) );
  NAND2_X1 U10316 ( .A1(n8991), .A2(n9629), .ZN(n8994) );
  INV_X1 U10317 ( .A(n9244), .ZN(n8992) );
  NOR2_X1 U10318 ( .A1(n8992), .A2(n9620), .ZN(n9001) );
  AOI21_X1 U10319 ( .B1(n9620), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9001), .ZN(
        n8993) );
  OAI211_X1 U10320 ( .C1(n8995), .C2(n9204), .A(n8994), .B(n8993), .ZN(
        P1_U3261) );
  INV_X1 U10321 ( .A(n8996), .ZN(n9000) );
  INV_X1 U10322 ( .A(n8997), .ZN(n8998) );
  NAND2_X1 U10323 ( .A1(n9245), .A2(n9629), .ZN(n9003) );
  AOI21_X1 U10324 ( .B1(n9620), .B2(P1_REG2_REG_30__SCAN_IN), .A(n9001), .ZN(
        n9002) );
  OAI211_X1 U10325 ( .C1(n9345), .C2(n9204), .A(n9003), .B(n9002), .ZN(
        P1_U3262) );
  NAND2_X1 U10326 ( .A1(n9005), .A2(n9007), .ZN(n9006) );
  NAND2_X1 U10327 ( .A1(n9004), .A2(n9006), .ZN(n9252) );
  XNOR2_X1 U10328 ( .A(n9008), .B(n8287), .ZN(n9009) );
  NAND2_X1 U10329 ( .A1(n9009), .A2(n9227), .ZN(n9012) );
  AOI22_X1 U10330 ( .A1(n9047), .A2(n9226), .B1(n9686), .B2(n9010), .ZN(n9011)
         );
  NAND2_X1 U10331 ( .A1(n9012), .A2(n9011), .ZN(n9256) );
  OAI211_X1 U10332 ( .C1(n4321), .C2(n9254), .A(n9626), .B(n9013), .ZN(n9253)
         );
  AOI22_X1 U10333 ( .A1(n9014), .A2(n9646), .B1(P1_REG2_REG_28__SCAN_IN), .B2(
        n9620), .ZN(n9017) );
  NAND2_X1 U10334 ( .A1(n9015), .A2(n9622), .ZN(n9016) );
  OAI211_X1 U10335 ( .C1(n9253), .C2(n9239), .A(n9017), .B(n9016), .ZN(n9018)
         );
  AOI21_X1 U10336 ( .B1(n9256), .B2(n9219), .A(n9018), .ZN(n9019) );
  OAI21_X1 U10337 ( .B1(n9252), .B2(n9222), .A(n9019), .ZN(P1_U3263) );
  XNOR2_X1 U10338 ( .A(n9020), .B(n9027), .ZN(n9261) );
  INV_X1 U10339 ( .A(n9261), .ZN(n9034) );
  AOI211_X1 U10340 ( .C1(n9021), .C2(n9038), .A(n9236), .B(n4321), .ZN(n9260)
         );
  NOR2_X1 U10341 ( .A1(n4577), .A2(n9204), .ZN(n9025) );
  OAI22_X1 U10342 ( .A1(n9023), .A2(n9206), .B1(n9219), .B2(n9022), .ZN(n9024)
         );
  AOI211_X1 U10343 ( .C1(n9260), .C2(n9629), .A(n9025), .B(n9024), .ZN(n9033)
         );
  OAI211_X1 U10344 ( .C1(n4854), .C2(n9027), .A(n9026), .B(n9227), .ZN(n9031)
         );
  AOI22_X1 U10345 ( .A1(n9029), .A2(n9686), .B1(n9615), .B2(n9028), .ZN(n9030)
         );
  NAND2_X1 U10346 ( .A1(n9031), .A2(n9030), .ZN(n9259) );
  NAND2_X1 U10347 ( .A1(n9259), .A2(n9219), .ZN(n9032) );
  OAI211_X1 U10348 ( .C1(n9034), .C2(n9222), .A(n9033), .B(n9032), .ZN(
        P1_U3264) );
  NAND2_X1 U10349 ( .A1(n9036), .A2(n9035), .ZN(n9037) );
  XNOR2_X1 U10350 ( .A(n9037), .B(n9046), .ZN(n9268) );
  INV_X1 U10351 ( .A(n9038), .ZN(n9039) );
  AOI211_X1 U10352 ( .C1(n9265), .C2(n9062), .A(n9236), .B(n9039), .ZN(n9264)
         );
  AOI22_X1 U10353 ( .A1(n9040), .A2(n9646), .B1(P1_REG2_REG_26__SCAN_IN), .B2(
        n9620), .ZN(n9041) );
  OAI21_X1 U10354 ( .B1(n9042), .B2(n9204), .A(n9041), .ZN(n9050) );
  NAND2_X1 U10355 ( .A1(n9044), .A2(n9043), .ZN(n9045) );
  XOR2_X1 U10356 ( .A(n9046), .B(n9045), .Z(n9048) );
  AOI222_X1 U10357 ( .A1(n9227), .A2(n9048), .B1(n9047), .B2(n9686), .C1(n9076), .C2(n9615), .ZN(n9267) );
  NOR2_X1 U10358 ( .A1(n9267), .A2(n9620), .ZN(n9049) );
  AOI211_X1 U10359 ( .C1(n9264), .C2(n9629), .A(n9050), .B(n9049), .ZN(n9051)
         );
  OAI21_X1 U10360 ( .B1(n9222), .B2(n9268), .A(n9051), .ZN(P1_U3265) );
  XNOR2_X1 U10361 ( .A(n9052), .B(n9058), .ZN(n9053) );
  AOI22_X1 U10362 ( .A1(n9053), .A2(n9227), .B1(n9615), .B2(n9092), .ZN(n9270)
         );
  NAND2_X1 U10363 ( .A1(n9054), .A2(n9055), .ZN(n9057) );
  NAND2_X1 U10364 ( .A1(n9057), .A2(n9056), .ZN(n9059) );
  XNOR2_X1 U10365 ( .A(n9059), .B(n9058), .ZN(n9273) );
  NAND2_X1 U10366 ( .A1(n9273), .A2(n9231), .ZN(n9067) );
  AOI22_X1 U10367 ( .A1(n9060), .A2(n9646), .B1(n9620), .B2(
        P1_REG2_REG_25__SCAN_IN), .ZN(n9061) );
  OAI21_X1 U10368 ( .B1(n9271), .B2(n9235), .A(n9061), .ZN(n9064) );
  OAI211_X1 U10369 ( .C1(n9080), .C2(n9354), .A(n9062), .B(n9626), .ZN(n9269)
         );
  NOR2_X1 U10370 ( .A1(n9269), .A2(n9239), .ZN(n9063) );
  AOI211_X1 U10371 ( .C1(n9622), .C2(n9065), .A(n9064), .B(n9063), .ZN(n9066)
         );
  OAI211_X1 U10372 ( .C1(n9620), .C2(n9270), .A(n9067), .B(n9066), .ZN(
        P1_U3266) );
  NAND2_X1 U10373 ( .A1(n9054), .A2(n9068), .ZN(n9069) );
  XOR2_X1 U10374 ( .A(n9073), .B(n9069), .Z(n9280) );
  INV_X1 U10375 ( .A(n9070), .ZN(n9071) );
  NOR2_X1 U10376 ( .A1(n9072), .A2(n9071), .ZN(n9079) );
  OAI21_X1 U10377 ( .B1(n9074), .B2(n9073), .A(n9227), .ZN(n9078) );
  AOI22_X1 U10378 ( .A1(n9076), .A2(n9686), .B1(n9615), .B2(n9075), .ZN(n9077)
         );
  OAI21_X1 U10379 ( .B1(n9079), .B2(n9078), .A(n9077), .ZN(n9276) );
  INV_X1 U10380 ( .A(n9095), .ZN(n9081) );
  AOI211_X1 U10381 ( .C1(n9278), .C2(n9081), .A(n9236), .B(n9080), .ZN(n9277)
         );
  NAND2_X1 U10382 ( .A1(n9277), .A2(n9629), .ZN(n9084) );
  AOI22_X1 U10383 ( .A1(n9620), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n9082), .B2(
        n9646), .ZN(n9083) );
  OAI211_X1 U10384 ( .C1(n9085), .C2(n9204), .A(n9084), .B(n9083), .ZN(n9086)
         );
  AOI21_X1 U10385 ( .B1(n9276), .B2(n9219), .A(n9086), .ZN(n9087) );
  OAI21_X1 U10386 ( .B1(n9280), .B2(n9222), .A(n9087), .ZN(P1_U3267) );
  XNOR2_X1 U10387 ( .A(n9088), .B(n9090), .ZN(n9283) );
  INV_X1 U10388 ( .A(n9283), .ZN(n9102) );
  OAI211_X1 U10389 ( .C1(n9091), .C2(n9090), .A(n9089), .B(n9227), .ZN(n9094)
         );
  AOI22_X1 U10390 ( .A1(n9092), .A2(n9686), .B1(n9615), .B2(n9295), .ZN(n9093)
         );
  NAND2_X1 U10391 ( .A1(n9094), .A2(n9093), .ZN(n9281) );
  AOI211_X1 U10392 ( .C1(n9096), .C2(n4317), .A(n9236), .B(n9095), .ZN(n9282)
         );
  NAND2_X1 U10393 ( .A1(n9282), .A2(n9629), .ZN(n9099) );
  AOI22_X1 U10394 ( .A1(n9620), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n9097), .B2(
        n9646), .ZN(n9098) );
  OAI211_X1 U10395 ( .C1(n9358), .C2(n9204), .A(n9099), .B(n9098), .ZN(n9100)
         );
  AOI21_X1 U10396 ( .B1(n9219), .B2(n9281), .A(n9100), .ZN(n9101) );
  OAI21_X1 U10397 ( .B1(n9102), .B2(n9222), .A(n9101), .ZN(P1_U3268) );
  XNOR2_X1 U10398 ( .A(n9103), .B(n9106), .ZN(n9105) );
  AOI22_X1 U10399 ( .A1(n9105), .A2(n9227), .B1(n9615), .B2(n9104), .ZN(n9288)
         );
  XNOR2_X1 U10400 ( .A(n9107), .B(n9106), .ZN(n9291) );
  NAND2_X1 U10401 ( .A1(n9291), .A2(n9231), .ZN(n9115) );
  INV_X1 U10402 ( .A(n9108), .ZN(n9109) );
  AOI22_X1 U10403 ( .A1(n9620), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n9109), .B2(
        n9646), .ZN(n9110) );
  OAI21_X1 U10404 ( .B1(n9235), .B2(n9289), .A(n9110), .ZN(n9113) );
  AOI21_X1 U10405 ( .B1(n4361), .B2(n9286), .A(n9236), .ZN(n9111) );
  NAND2_X1 U10406 ( .A1(n9111), .A2(n4317), .ZN(n9287) );
  NOR2_X1 U10407 ( .A1(n9287), .A2(n9239), .ZN(n9112) );
  AOI211_X1 U10408 ( .C1(n9622), .C2(n9286), .A(n9113), .B(n9112), .ZN(n9114)
         );
  OAI211_X1 U10409 ( .C1(n9620), .C2(n9288), .A(n9115), .B(n9114), .ZN(
        P1_U3269) );
  NAND2_X1 U10410 ( .A1(n9118), .A2(n9117), .ZN(n9294) );
  NAND3_X1 U10411 ( .A1(n9116), .A2(n9294), .A3(n9231), .ZN(n9132) );
  OAI22_X1 U10412 ( .A1(n9235), .A2(n9120), .B1(n9119), .B2(n9219), .ZN(n9121)
         );
  AOI21_X1 U10413 ( .B1(n9296), .B2(n9622), .A(n9121), .ZN(n9131) );
  XNOR2_X1 U10414 ( .A(n9122), .B(n8270), .ZN(n9124) );
  AOI22_X1 U10415 ( .A1(n9124), .A2(n9227), .B1(n9226), .B2(n9123), .ZN(n9299)
         );
  INV_X1 U10416 ( .A(n9299), .ZN(n9129) );
  OAI211_X1 U10417 ( .C1(n9139), .C2(n9125), .A(n9626), .B(n4361), .ZN(n9297)
         );
  OAI22_X1 U10418 ( .A1(n9297), .A2(n9127), .B1(n9206), .B2(n9126), .ZN(n9128)
         );
  OAI21_X1 U10419 ( .B1(n9129), .B2(n9128), .A(n9219), .ZN(n9130) );
  NAND3_X1 U10420 ( .A1(n9132), .A2(n9131), .A3(n9130), .ZN(P1_U3270) );
  NAND2_X1 U10421 ( .A1(n9149), .A2(n9133), .ZN(n9134) );
  XOR2_X1 U10422 ( .A(n9134), .B(n9137), .Z(n9135) );
  OAI222_X1 U10423 ( .A1(n9705), .A2(n9136), .B1(n9217), .B2(n9178), .C1(n9135), .C2(n9617), .ZN(n9301) );
  INV_X1 U10424 ( .A(n9301), .ZN(n9148) );
  XNOR2_X1 U10425 ( .A(n9138), .B(n9137), .ZN(n9303) );
  NAND2_X1 U10426 ( .A1(n9303), .A2(n9231), .ZN(n9147) );
  INV_X1 U10427 ( .A(n9156), .ZN(n9140) );
  AOI211_X1 U10428 ( .C1(n9141), .C2(n9140), .A(n9236), .B(n9139), .ZN(n9302)
         );
  NOR2_X1 U10429 ( .A1(n9367), .A2(n9204), .ZN(n9145) );
  OAI22_X1 U10430 ( .A1(n9219), .A2(n9143), .B1(n9142), .B2(n9206), .ZN(n9144)
         );
  AOI211_X1 U10431 ( .C1(n9302), .C2(n9629), .A(n9145), .B(n9144), .ZN(n9146)
         );
  OAI211_X1 U10432 ( .C1(n9620), .C2(n9148), .A(n9147), .B(n9146), .ZN(
        P1_U3271) );
  INV_X1 U10433 ( .A(n9149), .ZN(n9150) );
  AOI21_X1 U10434 ( .B1(n9151), .B2(n9154), .A(n9150), .ZN(n9152) );
  OAI222_X1 U10435 ( .A1(n9705), .A2(n9153), .B1(n9217), .B2(n9199), .C1(n9617), .C2(n9152), .ZN(n9306) );
  INV_X1 U10436 ( .A(n9306), .ZN(n9164) );
  XOR2_X1 U10437 ( .A(n9155), .B(n9154), .Z(n9308) );
  NAND2_X1 U10438 ( .A1(n9308), .A2(n9231), .ZN(n9163) );
  AOI211_X1 U10439 ( .C1(n9157), .C2(n9180), .A(n9236), .B(n9156), .ZN(n9307)
         );
  INV_X1 U10440 ( .A(n9157), .ZN(n9371) );
  NOR2_X1 U10441 ( .A1(n9371), .A2(n9204), .ZN(n9161) );
  OAI22_X1 U10442 ( .A1(n9219), .A2(n9159), .B1(n9158), .B2(n9206), .ZN(n9160)
         );
  AOI211_X1 U10443 ( .C1(n9307), .C2(n9629), .A(n9161), .B(n9160), .ZN(n9162)
         );
  OAI211_X1 U10444 ( .C1(n9620), .C2(n9164), .A(n9163), .B(n9162), .ZN(
        P1_U3272) );
  INV_X1 U10445 ( .A(n9165), .ZN(n9166) );
  AOI21_X1 U10446 ( .B1(n9197), .B2(n9167), .A(n9166), .ZN(n9168) );
  XNOR2_X1 U10447 ( .A(n9168), .B(n9174), .ZN(n9170) );
  AOI22_X1 U10448 ( .A1(n9170), .A2(n9227), .B1(n9615), .B2(n9169), .ZN(n9316)
         );
  INV_X1 U10449 ( .A(n9171), .ZN(n9172) );
  AOI21_X1 U10450 ( .B1(n9174), .B2(n9173), .A(n9172), .ZN(n9311) );
  NAND2_X1 U10451 ( .A1(n9311), .A2(n9231), .ZN(n9185) );
  INV_X1 U10452 ( .A(n9175), .ZN(n9176) );
  AOI22_X1 U10453 ( .A1(n9620), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9176), .B2(
        n9646), .ZN(n9177) );
  OAI21_X1 U10454 ( .B1(n9235), .B2(n9178), .A(n9177), .ZN(n9183) );
  INV_X1 U10455 ( .A(n9179), .ZN(n9189) );
  INV_X1 U10456 ( .A(n9313), .ZN(n9181) );
  OAI211_X1 U10457 ( .C1(n9189), .C2(n9181), .A(n9626), .B(n9180), .ZN(n9314)
         );
  NOR2_X1 U10458 ( .A1(n9314), .A2(n9239), .ZN(n9182) );
  AOI211_X1 U10459 ( .C1(n9622), .C2(n9313), .A(n9183), .B(n9182), .ZN(n9184)
         );
  OAI211_X1 U10460 ( .C1(n9620), .C2(n9316), .A(n9185), .B(n9184), .ZN(
        P1_U3273) );
  NAND2_X1 U10461 ( .A1(n9187), .A2(n9186), .ZN(n9188) );
  XOR2_X1 U10462 ( .A(n9196), .B(n9188), .Z(n9322) );
  INV_X1 U10463 ( .A(n9203), .ZN(n9190) );
  AOI211_X1 U10464 ( .C1(n9320), .C2(n9190), .A(n9236), .B(n9189), .ZN(n9319)
         );
  NOR2_X1 U10465 ( .A1(n9191), .A2(n9204), .ZN(n9195) );
  OAI22_X1 U10466 ( .A1(n9219), .A2(n9193), .B1(n9192), .B2(n9206), .ZN(n9194)
         );
  AOI211_X1 U10467 ( .C1(n9319), .C2(n9629), .A(n9195), .B(n9194), .ZN(n9201)
         );
  XNOR2_X1 U10468 ( .A(n9197), .B(n9196), .ZN(n9198) );
  OAI222_X1 U10469 ( .A1(n9705), .A2(n9199), .B1(n9217), .B2(n9331), .C1(n9617), .C2(n9198), .ZN(n9318) );
  NAND2_X1 U10470 ( .A1(n9318), .A2(n9219), .ZN(n9200) );
  OAI211_X1 U10471 ( .C1(n9322), .C2(n9222), .A(n9201), .B(n9200), .ZN(
        P1_U3274) );
  XNOR2_X1 U10472 ( .A(n9202), .B(n9213), .ZN(n9327) );
  AOI211_X1 U10473 ( .C1(n9325), .C2(n9237), .A(n9236), .B(n9203), .ZN(n9324)
         );
  INV_X1 U10474 ( .A(n9325), .ZN(n9205) );
  NOR2_X1 U10475 ( .A1(n9205), .A2(n9204), .ZN(n9210) );
  OAI22_X1 U10476 ( .A1(n9219), .A2(n9208), .B1(n9207), .B2(n9206), .ZN(n9209)
         );
  AOI211_X1 U10477 ( .C1(n9324), .C2(n9629), .A(n9210), .B(n9209), .ZN(n9221)
         );
  NAND2_X1 U10478 ( .A1(n9212), .A2(n9211), .ZN(n9214) );
  XNOR2_X1 U10479 ( .A(n9214), .B(n9213), .ZN(n9215) );
  OAI222_X1 U10480 ( .A1(n9705), .A2(n9218), .B1(n9217), .B2(n9216), .C1(n9215), .C2(n9617), .ZN(n9323) );
  NAND2_X1 U10481 ( .A1(n9323), .A2(n9219), .ZN(n9220) );
  OAI211_X1 U10482 ( .C1(n9327), .C2(n9222), .A(n9221), .B(n9220), .ZN(
        P1_U3275) );
  XNOR2_X1 U10483 ( .A(n9224), .B(n9223), .ZN(n9228) );
  AOI22_X1 U10484 ( .A1(n9228), .A2(n9227), .B1(n9226), .B2(n9225), .ZN(n9330)
         );
  XNOR2_X1 U10485 ( .A(n9229), .B(n9230), .ZN(n9333) );
  NAND2_X1 U10486 ( .A1(n9333), .A2(n9231), .ZN(n9243) );
  INV_X1 U10487 ( .A(n9232), .ZN(n9233) );
  AOI22_X1 U10488 ( .A1(n9620), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n9233), .B2(
        n9646), .ZN(n9234) );
  OAI21_X1 U10489 ( .B1(n9235), .B2(n9331), .A(n9234), .ZN(n9241) );
  AOI21_X1 U10490 ( .B1(n4852), .B2(n9328), .A(n9236), .ZN(n9238) );
  NAND2_X1 U10491 ( .A1(n9238), .A2(n9237), .ZN(n9329) );
  NOR2_X1 U10492 ( .A1(n9329), .A2(n9239), .ZN(n9240) );
  AOI211_X1 U10493 ( .C1(n9622), .C2(n9328), .A(n9241), .B(n9240), .ZN(n9242)
         );
  OAI211_X1 U10494 ( .C1(n9620), .C2(n9330), .A(n9243), .B(n9242), .ZN(
        P1_U3276) );
  NOR2_X1 U10495 ( .A1(n9245), .A2(n9244), .ZN(n9343) );
  MUX2_X1 U10496 ( .A(n8081), .B(n9343), .S(n9733), .Z(n9246) );
  OAI21_X1 U10497 ( .B1(n9345), .B2(n9342), .A(n9246), .ZN(P1_U3553) );
  AOI21_X1 U10498 ( .B1(n9695), .B2(n9248), .A(n9247), .ZN(n9249) );
  OAI21_X1 U10499 ( .B1(n9251), .B2(n9699), .A(n4855), .ZN(n9346) );
  MUX2_X1 U10500 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9346), .S(n9733), .Z(
        P1_U3552) );
  OAI21_X1 U10501 ( .B1(n9254), .B2(n9678), .A(n9253), .ZN(n9255) );
  NOR2_X1 U10502 ( .A1(n9256), .A2(n9255), .ZN(n9257) );
  NAND2_X1 U10503 ( .A1(n9258), .A2(n9257), .ZN(n9347) );
  MUX2_X1 U10504 ( .A(n9347), .B(P1_REG1_REG_28__SCAN_IN), .S(n9731), .Z(
        P1_U3551) );
  INV_X1 U10505 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n9262) );
  AOI211_X1 U10506 ( .C1(n9261), .C2(n9710), .A(n9260), .B(n9259), .ZN(n9348)
         );
  MUX2_X1 U10507 ( .A(n9262), .B(n9348), .S(n9733), .Z(n9263) );
  OAI21_X1 U10508 ( .B1(n4577), .B2(n9342), .A(n9263), .ZN(P1_U3550) );
  AOI21_X1 U10509 ( .B1(n9695), .B2(n9265), .A(n9264), .ZN(n9266) );
  OAI211_X1 U10510 ( .C1(n9268), .C2(n9699), .A(n9267), .B(n9266), .ZN(n9351)
         );
  MUX2_X1 U10511 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9351), .S(n9733), .Z(
        P1_U3549) );
  INV_X1 U10512 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n9274) );
  OAI211_X1 U10513 ( .C1(n9271), .C2(n9705), .A(n9270), .B(n9269), .ZN(n9272)
         );
  AOI21_X1 U10514 ( .B1(n9273), .B2(n9710), .A(n9272), .ZN(n9352) );
  MUX2_X1 U10515 ( .A(n9274), .B(n9352), .S(n9733), .Z(n9275) );
  OAI21_X1 U10516 ( .B1(n9354), .B2(n9342), .A(n9275), .ZN(P1_U3548) );
  AOI211_X1 U10517 ( .C1(n9695), .C2(n9278), .A(n9277), .B(n9276), .ZN(n9279)
         );
  OAI21_X1 U10518 ( .B1(n9280), .B2(n9699), .A(n9279), .ZN(n9355) );
  MUX2_X1 U10519 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9355), .S(n9733), .Z(
        P1_U3547) );
  INV_X1 U10520 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n9284) );
  AOI211_X1 U10521 ( .C1(n9283), .C2(n9710), .A(n9282), .B(n9281), .ZN(n9356)
         );
  MUX2_X1 U10522 ( .A(n9284), .B(n9356), .S(n9733), .Z(n9285) );
  OAI21_X1 U10523 ( .B1(n9358), .B2(n9342), .A(n9285), .ZN(P1_U3546) );
  INV_X1 U10524 ( .A(n9286), .ZN(n9362) );
  INV_X1 U10525 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n9292) );
  OAI211_X1 U10526 ( .C1(n9289), .C2(n9705), .A(n9288), .B(n9287), .ZN(n9290)
         );
  AOI21_X1 U10527 ( .B1(n9291), .B2(n9710), .A(n9290), .ZN(n9359) );
  MUX2_X1 U10528 ( .A(n9292), .B(n9359), .S(n9733), .Z(n9293) );
  OAI21_X1 U10529 ( .B1(n9362), .B2(n9342), .A(n9293), .ZN(P1_U3545) );
  NAND3_X1 U10530 ( .A1(n9116), .A2(n9294), .A3(n9710), .ZN(n9300) );
  AOI22_X1 U10531 ( .A1(n9296), .A2(n9695), .B1(n9686), .B2(n9295), .ZN(n9298)
         );
  NAND4_X1 U10532 ( .A1(n9300), .A2(n9299), .A3(n9298), .A4(n9297), .ZN(n9363)
         );
  MUX2_X1 U10533 ( .A(n9363), .B(P1_REG1_REG_21__SCAN_IN), .S(n9731), .Z(
        P1_U3544) );
  AOI211_X1 U10534 ( .C1(n9303), .C2(n9710), .A(n9302), .B(n9301), .ZN(n9364)
         );
  MUX2_X1 U10535 ( .A(n9304), .B(n9364), .S(n9733), .Z(n9305) );
  OAI21_X1 U10536 ( .B1(n9367), .B2(n9342), .A(n9305), .ZN(P1_U3543) );
  AOI211_X1 U10537 ( .C1(n9308), .C2(n9710), .A(n9307), .B(n9306), .ZN(n9368)
         );
  MUX2_X1 U10538 ( .A(n9309), .B(n9368), .S(n9733), .Z(n9310) );
  OAI21_X1 U10539 ( .B1(n9371), .B2(n9342), .A(n9310), .ZN(P1_U3542) );
  NAND2_X1 U10540 ( .A1(n9311), .A2(n9710), .ZN(n9317) );
  AOI22_X1 U10541 ( .A1(n9313), .A2(n9695), .B1(n9686), .B2(n9312), .ZN(n9315)
         );
  NAND4_X1 U10542 ( .A1(n9317), .A2(n9316), .A3(n9315), .A4(n9314), .ZN(n9372)
         );
  MUX2_X1 U10543 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9372), .S(n9733), .Z(
        P1_U3541) );
  AOI211_X1 U10544 ( .C1(n9695), .C2(n9320), .A(n9319), .B(n9318), .ZN(n9321)
         );
  OAI21_X1 U10545 ( .B1(n9322), .B2(n9699), .A(n9321), .ZN(n9373) );
  MUX2_X1 U10546 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9373), .S(n9733), .Z(
        P1_U3540) );
  AOI211_X1 U10547 ( .C1(n9695), .C2(n9325), .A(n9324), .B(n9323), .ZN(n9326)
         );
  OAI21_X1 U10548 ( .B1(n9699), .B2(n9327), .A(n9326), .ZN(n9374) );
  MUX2_X1 U10549 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9374), .S(n9733), .Z(
        P1_U3539) );
  OAI211_X1 U10550 ( .C1(n9331), .C2(n9705), .A(n9330), .B(n9329), .ZN(n9332)
         );
  AOI21_X1 U10551 ( .B1(n9333), .B2(n9710), .A(n9332), .ZN(n9375) );
  MUX2_X1 U10552 ( .A(n9334), .B(n9375), .S(n9733), .Z(n9335) );
  OAI21_X1 U10553 ( .B1(n4583), .B2(n9342), .A(n9335), .ZN(P1_U3538) );
  INV_X1 U10554 ( .A(n9336), .ZN(n9339) );
  INV_X1 U10555 ( .A(n9712), .ZN(n9684) );
  AOI211_X1 U10556 ( .C1(n9339), .C2(n9684), .A(n9338), .B(n9337), .ZN(n9377)
         );
  MUX2_X1 U10557 ( .A(n9340), .B(n9377), .S(n9733), .Z(n9341) );
  OAI21_X1 U10558 ( .B1(n9380), .B2(n9342), .A(n9341), .ZN(P1_U3536) );
  MUX2_X1 U10559 ( .A(n8083), .B(n9343), .S(n9720), .Z(n9344) );
  OAI21_X1 U10560 ( .B1(n9345), .B2(n9379), .A(n9344), .ZN(P1_U3521) );
  MUX2_X1 U10561 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9346), .S(n9720), .Z(
        P1_U3520) );
  MUX2_X1 U10562 ( .A(n9347), .B(P1_REG0_REG_28__SCAN_IN), .S(n9718), .Z(
        P1_U3519) );
  INV_X1 U10563 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n9349) );
  MUX2_X1 U10564 ( .A(n9349), .B(n9348), .S(n9720), .Z(n9350) );
  OAI21_X1 U10565 ( .B1(n4577), .B2(n9379), .A(n9350), .ZN(P1_U3518) );
  MUX2_X1 U10566 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9351), .S(n9720), .Z(
        P1_U3517) );
  MUX2_X1 U10567 ( .A(n10158), .B(n9352), .S(n9720), .Z(n9353) );
  OAI21_X1 U10568 ( .B1(n9354), .B2(n9379), .A(n9353), .ZN(P1_U3516) );
  MUX2_X1 U10569 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9355), .S(n9720), .Z(
        P1_U3515) );
  MUX2_X1 U10570 ( .A(n10066), .B(n9356), .S(n9720), .Z(n9357) );
  OAI21_X1 U10571 ( .B1(n9358), .B2(n9379), .A(n9357), .ZN(P1_U3514) );
  INV_X1 U10572 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n9360) );
  MUX2_X1 U10573 ( .A(n9360), .B(n9359), .S(n9720), .Z(n9361) );
  OAI21_X1 U10574 ( .B1(n9362), .B2(n9379), .A(n9361), .ZN(P1_U3513) );
  MUX2_X1 U10575 ( .A(n9363), .B(P1_REG0_REG_21__SCAN_IN), .S(n9718), .Z(
        P1_U3512) );
  INV_X1 U10576 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n9365) );
  MUX2_X1 U10577 ( .A(n9365), .B(n9364), .S(n9720), .Z(n9366) );
  OAI21_X1 U10578 ( .B1(n9367), .B2(n9379), .A(n9366), .ZN(P1_U3511) );
  INV_X1 U10579 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n9369) );
  MUX2_X1 U10580 ( .A(n9369), .B(n9368), .S(n9720), .Z(n9370) );
  OAI21_X1 U10581 ( .B1(n9371), .B2(n9379), .A(n9370), .ZN(P1_U3510) );
  MUX2_X1 U10582 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9372), .S(n9720), .Z(
        P1_U3508) );
  MUX2_X1 U10583 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9373), .S(n9720), .Z(
        P1_U3505) );
  MUX2_X1 U10584 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9374), .S(n9720), .Z(
        P1_U3502) );
  MUX2_X1 U10585 ( .A(n10062), .B(n9375), .S(n9720), .Z(n9376) );
  OAI21_X1 U10586 ( .B1(n4583), .B2(n9379), .A(n9376), .ZN(P1_U3499) );
  MUX2_X1 U10587 ( .A(n5990), .B(n9377), .S(n9720), .Z(n9378) );
  OAI21_X1 U10588 ( .B1(n9380), .B2(n9379), .A(n9378), .ZN(P1_U3493) );
  AND2_X1 U10589 ( .A1(n9654), .A2(n9381), .ZN(n9650) );
  MUX2_X1 U10590 ( .A(P1_D_REG_0__SCAN_IN), .B(n9382), .S(n9650), .Z(P1_U3440)
         );
  INV_X1 U10591 ( .A(n7791), .ZN(n9388) );
  INV_X1 U10592 ( .A(n9383), .ZN(n9384) );
  NOR4_X1 U10593 ( .A1(n9384), .A2(P1_IR_REG_30__SCAN_IN), .A3(n9385), .A4(
        P1_U3084), .ZN(n9386) );
  AOI21_X1 U10594 ( .B1(n9389), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9386), .ZN(
        n9387) );
  OAI21_X1 U10595 ( .B1(n9388), .B2(n9391), .A(n9387), .ZN(P1_U3322) );
  AOI22_X1 U10596 ( .A1(n5771), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n9389), .ZN(n9390) );
  OAI21_X1 U10597 ( .B1(n9392), .B2(n9391), .A(n9390), .ZN(P1_U3323) );
  MUX2_X1 U10598 ( .A(n9393), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  MUX2_X1 U10599 ( .A(n9394), .B(P1_ADDR_REG_19__SCAN_IN), .S(
        P2_ADDR_REG_19__SCAN_IN), .Z(n9424) );
  NOR2_X1 U10600 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n9395) );
  AOI21_X1 U10601 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n9395), .ZN(n9967) );
  NOR2_X1 U10602 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n9396) );
  AOI21_X1 U10603 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n9396), .ZN(n9970) );
  NOR2_X1 U10604 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n9397) );
  AOI21_X1 U10605 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n9397), .ZN(n9973) );
  NOR2_X1 U10606 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n9398) );
  AOI21_X1 U10607 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n9398), .ZN(n9976) );
  NOR2_X1 U10608 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n9399) );
  AOI21_X1 U10609 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n9399), .ZN(n9979) );
  NOR2_X1 U10610 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n9405) );
  XNOR2_X1 U10611 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10198) );
  NAND2_X1 U10612 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n9403) );
  XOR2_X1 U10613 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10196) );
  NAND2_X1 U10614 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n9401) );
  INV_X1 U10615 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n9497) );
  XNOR2_X1 U10616 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(n9497), .ZN(n10194) );
  AOI21_X1 U10617 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9960) );
  NAND3_X1 U10618 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n9962) );
  OAI21_X1 U10619 ( .B1(n9960), .B2(n9964), .A(n9962), .ZN(n10193) );
  NAND2_X1 U10620 ( .A1(n10194), .A2(n10193), .ZN(n9400) );
  NAND2_X1 U10621 ( .A1(n9401), .A2(n9400), .ZN(n10195) );
  NAND2_X1 U10622 ( .A1(n10196), .A2(n10195), .ZN(n9402) );
  NAND2_X1 U10623 ( .A1(n9403), .A2(n9402), .ZN(n10197) );
  NOR2_X1 U10624 ( .A1(n10198), .A2(n10197), .ZN(n9404) );
  NOR2_X1 U10625 ( .A1(n9405), .A2(n9404), .ZN(n9406) );
  NOR2_X1 U10626 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n9406), .ZN(n10181) );
  AND2_X1 U10627 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n9406), .ZN(n10180) );
  NOR2_X1 U10628 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10180), .ZN(n9407) );
  NOR2_X1 U10629 ( .A1(n10181), .A2(n9407), .ZN(n9408) );
  NAND2_X1 U10630 ( .A1(n9408), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n9410) );
  INV_X1 U10631 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n10093) );
  XNOR2_X1 U10632 ( .A(n9408), .B(n10093), .ZN(n10179) );
  NAND2_X1 U10633 ( .A1(n10179), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n9409) );
  NAND2_X1 U10634 ( .A1(n9410), .A2(n9409), .ZN(n9411) );
  NAND2_X1 U10635 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n9411), .ZN(n9413) );
  XOR2_X1 U10636 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n9411), .Z(n10183) );
  NAND2_X1 U10637 ( .A1(n10183), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n9412) );
  NAND2_X1 U10638 ( .A1(n9413), .A2(n9412), .ZN(n9414) );
  NAND2_X1 U10639 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n9414), .ZN(n9416) );
  XOR2_X1 U10640 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n9414), .Z(n10189) );
  NAND2_X1 U10641 ( .A1(n10189), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n9415) );
  NAND2_X1 U10642 ( .A1(n9416), .A2(n9415), .ZN(n9417) );
  AND2_X1 U10643 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n9417), .ZN(n9418) );
  XNOR2_X1 U10644 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n9417), .ZN(n10191) );
  NOR2_X1 U10645 ( .A1(n10192), .A2(n10191), .ZN(n10190) );
  NOR2_X1 U10646 ( .A1(n9418), .A2(n10190), .ZN(n9988) );
  NAND2_X1 U10647 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n9419) );
  OAI21_X1 U10648 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n9419), .ZN(n9987) );
  NOR2_X1 U10649 ( .A1(n9988), .A2(n9987), .ZN(n9986) );
  AOI21_X1 U10650 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n9986), .ZN(n9985) );
  NAND2_X1 U10651 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n9420) );
  OAI21_X1 U10652 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n9420), .ZN(n9984) );
  NOR2_X1 U10653 ( .A1(n9985), .A2(n9984), .ZN(n9983) );
  AOI21_X1 U10654 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n9983), .ZN(n9982) );
  NOR2_X1 U10655 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n9421) );
  AOI21_X1 U10656 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n9421), .ZN(n9981) );
  NAND2_X1 U10657 ( .A1(n9982), .A2(n9981), .ZN(n9980) );
  OAI21_X1 U10658 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n9980), .ZN(n9978) );
  NAND2_X1 U10659 ( .A1(n9979), .A2(n9978), .ZN(n9977) );
  OAI21_X1 U10660 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n9977), .ZN(n9975) );
  NAND2_X1 U10661 ( .A1(n9976), .A2(n9975), .ZN(n9974) );
  OAI21_X1 U10662 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n9974), .ZN(n9972) );
  NAND2_X1 U10663 ( .A1(n9973), .A2(n9972), .ZN(n9971) );
  OAI21_X1 U10664 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n9971), .ZN(n9969) );
  NAND2_X1 U10665 ( .A1(n9970), .A2(n9969), .ZN(n9968) );
  OAI21_X1 U10666 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n9968), .ZN(n9966) );
  NAND2_X1 U10667 ( .A1(n9967), .A2(n9966), .ZN(n9965) );
  OAI21_X1 U10668 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n9965), .ZN(n10185) );
  NOR2_X1 U10669 ( .A1(n10186), .A2(n10185), .ZN(n9422) );
  NAND2_X1 U10670 ( .A1(n10186), .A2(n10185), .ZN(n10184) );
  OAI21_X1 U10671 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n9422), .A(n10184), .ZN(
        n9423) );
  XOR2_X1 U10672 ( .A(n9424), .B(n9423), .Z(ADD_1071_U4) );
  AOI22_X1 U10673 ( .A1(n9567), .A2(n9425), .B1(n9535), .B2(
        P1_ADDR_REG_3__SCAN_IN), .ZN(n9436) );
  AOI21_X1 U10674 ( .B1(n9428), .B2(n9427), .A(n9426), .ZN(n9429) );
  NAND2_X1 U10675 ( .A1(n9595), .A2(n9429), .ZN(n9434) );
  OAI211_X1 U10676 ( .C1(n9432), .C2(n9431), .A(n9585), .B(n9430), .ZN(n9433)
         );
  NAND4_X1 U10677 ( .A1(n9436), .A2(n9435), .A3(n9434), .A4(n9433), .ZN(
        P1_U3244) );
  AOI22_X1 U10678 ( .A1(n9781), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n9447) );
  NAND2_X1 U10679 ( .A1(n9791), .A2(n9437), .ZN(n9446) );
  OAI211_X1 U10680 ( .C1(n9440), .C2(n9439), .A(n9786), .B(n9438), .ZN(n9445)
         );
  OAI211_X1 U10681 ( .C1(n9443), .C2(n9442), .A(n9783), .B(n9441), .ZN(n9444)
         );
  NAND4_X1 U10682 ( .A1(n9447), .A2(n9446), .A3(n9445), .A4(n9444), .ZN(
        P2_U3247) );
  OAI21_X1 U10683 ( .B1(n9449), .B2(n9678), .A(n9448), .ZN(n9451) );
  AOI211_X1 U10684 ( .C1(n9684), .C2(n9452), .A(n9451), .B(n9450), .ZN(n9454)
         );
  AOI22_X1 U10685 ( .A1(n9720), .A2(n9454), .B1(n5960), .B2(n9718), .ZN(
        P1_U3484) );
  AOI22_X1 U10686 ( .A1(n9733), .A2(n9454), .B1(n9453), .B2(n9731), .ZN(
        P1_U3533) );
  OAI21_X1 U10687 ( .B1(n4584), .B2(n9678), .A(n9455), .ZN(n9456) );
  AOI211_X1 U10688 ( .C1(n9458), .C2(n9710), .A(n9457), .B(n9456), .ZN(n9467)
         );
  AOI22_X1 U10689 ( .A1(n9733), .A2(n9467), .B1(n6001), .B2(n9731), .ZN(
        P1_U3537) );
  AOI22_X1 U10690 ( .A1(n9460), .A2(n9695), .B1(n9686), .B2(n9459), .ZN(n9462)
         );
  NAND3_X1 U10691 ( .A1(n9463), .A2(n9462), .A3(n9461), .ZN(n9464) );
  AOI21_X1 U10692 ( .B1(n9465), .B2(n9710), .A(n9464), .ZN(n9468) );
  AOI22_X1 U10693 ( .A1(n9733), .A2(n9468), .B1(n5928), .B2(n9731), .ZN(
        P1_U3535) );
  INV_X1 U10694 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n9466) );
  AOI22_X1 U10695 ( .A1(n9720), .A2(n9467), .B1(n9466), .B2(n9718), .ZN(
        P1_U3496) );
  AOI22_X1 U10696 ( .A1(n9720), .A2(n9468), .B1(n5933), .B2(n9718), .ZN(
        P1_U3490) );
  XNOR2_X1 U10697 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U10698 ( .A(P2_RD_REG_SCAN_IN), .B(P1_RD_REG_SCAN_IN), .ZN(U126) );
  INV_X1 U10699 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n9476) );
  NOR2_X1 U10700 ( .A1(n9479), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n9469) );
  NOR2_X1 U10701 ( .A1(n9469), .A2(n5718), .ZN(n9470) );
  XNOR2_X1 U10702 ( .A(n9470), .B(n5573), .ZN(n9483) );
  NAND2_X1 U10703 ( .A1(n4568), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n9472) );
  AOI21_X1 U10704 ( .B1(n9479), .B2(n9472), .A(n9471), .ZN(n9473) );
  AOI22_X1 U10705 ( .A1(n9535), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(n9483), .B2(
        n9473), .ZN(n9475) );
  OR3_X1 U10706 ( .A1(n9605), .A2(P1_REG1_REG_0__SCAN_IN), .A3(n5573), .ZN(
        n9474) );
  OAI211_X1 U10707 ( .C1(P1_STATE_REG_SCAN_IN), .C2(n9476), .A(n9475), .B(
        n9474), .ZN(P1_U3241) );
  OAI21_X1 U10708 ( .B1(n9478), .B2(n9477), .A(n4624), .ZN(n9494) );
  NAND2_X1 U10709 ( .A1(n4568), .A2(n9479), .ZN(n9481) );
  OR2_X1 U10710 ( .A1(n9480), .A2(n9481), .ZN(n9486) );
  INV_X1 U10711 ( .A(n9481), .ZN(n9482) );
  OAI21_X1 U10712 ( .B1(n9483), .B2(n9482), .A(P1_U4006), .ZN(n9484) );
  INV_X1 U10713 ( .A(n9484), .ZN(n9485) );
  NAND2_X1 U10714 ( .A1(n9486), .A2(n9485), .ZN(n9508) );
  XNOR2_X1 U10715 ( .A(n9488), .B(n9487), .ZN(n9490) );
  INV_X1 U10716 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n9489) );
  OAI22_X1 U10717 ( .A1(n9605), .A2(n9490), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9489), .ZN(n9491) );
  AOI21_X1 U10718 ( .B1(n9567), .B2(n9492), .A(n9491), .ZN(n9493) );
  OAI211_X1 U10719 ( .C1(n9580), .C2(n9494), .A(n9508), .B(n9493), .ZN(n9495)
         );
  INV_X1 U10720 ( .A(n9495), .ZN(n9496) );
  OAI21_X1 U10721 ( .B1(n9609), .B2(n9497), .A(n9496), .ZN(P1_U3243) );
  OAI21_X1 U10722 ( .B1(n4334), .B2(n9499), .A(n9498), .ZN(n9500) );
  AOI22_X1 U10723 ( .A1(n9501), .A2(n9567), .B1(n9595), .B2(n9500), .ZN(n9510)
         );
  AOI21_X1 U10724 ( .B1(n9504), .B2(n9503), .A(n9502), .ZN(n9505) );
  NOR2_X1 U10725 ( .A1(n9605), .A2(n9505), .ZN(n9506) );
  AOI211_X1 U10726 ( .C1(P1_ADDR_REG_4__SCAN_IN), .C2(n9535), .A(n9507), .B(
        n9506), .ZN(n9509) );
  NAND3_X1 U10727 ( .A1(n9510), .A2(n9509), .A3(n9508), .ZN(P1_U3245) );
  AOI22_X1 U10728 ( .A1(n9567), .A2(n9511), .B1(n9535), .B2(
        P1_ADDR_REG_5__SCAN_IN), .ZN(n9522) );
  OAI21_X1 U10729 ( .B1(n9514), .B2(n9513), .A(n9512), .ZN(n9515) );
  NAND2_X1 U10730 ( .A1(n9595), .A2(n9515), .ZN(n9520) );
  OAI211_X1 U10731 ( .C1(n9518), .C2(n9517), .A(n9585), .B(n9516), .ZN(n9519)
         );
  NAND4_X1 U10732 ( .A1(n9522), .A2(n9521), .A3(n9520), .A4(n9519), .ZN(
        P1_U3246) );
  AOI22_X1 U10733 ( .A1(n9567), .A2(n9523), .B1(n9535), .B2(
        P1_ADDR_REG_8__SCAN_IN), .ZN(n9534) );
  OAI21_X1 U10734 ( .B1(n9526), .B2(n9525), .A(n9524), .ZN(n9527) );
  NAND2_X1 U10735 ( .A1(n9527), .A2(n9595), .ZN(n9532) );
  OAI211_X1 U10736 ( .C1(n9530), .C2(n9529), .A(n9585), .B(n9528), .ZN(n9531)
         );
  NAND4_X1 U10737 ( .A1(n9534), .A2(n9533), .A3(n9532), .A4(n9531), .ZN(
        P1_U3249) );
  AOI22_X1 U10738 ( .A1(n9567), .A2(n9536), .B1(n9535), .B2(
        P1_ADDR_REG_11__SCAN_IN), .ZN(n9548) );
  AOI21_X1 U10739 ( .B1(n9539), .B2(n9538), .A(n9537), .ZN(n9540) );
  OR2_X1 U10740 ( .A1(n9540), .A2(n9605), .ZN(n9546) );
  OAI21_X1 U10741 ( .B1(n9543), .B2(n9542), .A(n9541), .ZN(n9544) );
  NAND2_X1 U10742 ( .A1(n9544), .A2(n9595), .ZN(n9545) );
  NAND4_X1 U10743 ( .A1(n9548), .A2(n9547), .A3(n9546), .A4(n9545), .ZN(
        P1_U3252) );
  INV_X1 U10744 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n9560) );
  INV_X1 U10745 ( .A(n9549), .ZN(n9554) );
  AOI211_X1 U10746 ( .C1(n9552), .C2(n9551), .A(n9550), .B(n9580), .ZN(n9553)
         );
  AOI211_X1 U10747 ( .C1(n9567), .C2(n9555), .A(n9554), .B(n9553), .ZN(n9559)
         );
  OAI211_X1 U10748 ( .C1(n9557), .C2(P1_REG1_REG_15__SCAN_IN), .A(n9585), .B(
        n9556), .ZN(n9558) );
  OAI211_X1 U10749 ( .C1(n9560), .C2(n9609), .A(n9559), .B(n9558), .ZN(
        P1_U3256) );
  INV_X1 U10750 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n9573) );
  AOI211_X1 U10751 ( .C1(n9563), .C2(n9562), .A(n9561), .B(n9580), .ZN(n9564)
         );
  AOI211_X1 U10752 ( .C1(n9567), .C2(n9566), .A(n9565), .B(n9564), .ZN(n9572)
         );
  OAI211_X1 U10753 ( .C1(n9570), .C2(n9569), .A(n9585), .B(n9568), .ZN(n9571)
         );
  OAI211_X1 U10754 ( .C1(n9573), .C2(n9609), .A(n9572), .B(n9571), .ZN(
        P1_U3257) );
  INV_X1 U10755 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9591) );
  NAND2_X1 U10756 ( .A1(n9575), .A2(n9574), .ZN(n9578) );
  INV_X1 U10757 ( .A(n9576), .ZN(n9577) );
  NAND2_X1 U10758 ( .A1(n9578), .A2(n9577), .ZN(n9579) );
  OAI211_X1 U10759 ( .C1(n9599), .C2(n9583), .A(n9582), .B(n9581), .ZN(n9584)
         );
  INV_X1 U10760 ( .A(n9584), .ZN(n9590) );
  OAI211_X1 U10761 ( .C1(n9588), .C2(n9587), .A(n9586), .B(n9585), .ZN(n9589)
         );
  OAI211_X1 U10762 ( .C1(n9591), .C2(n9609), .A(n9590), .B(n9589), .ZN(
        P1_U3258) );
  INV_X1 U10763 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10187) );
  AOI21_X1 U10764 ( .B1(n9594), .B2(n9593), .A(n9592), .ZN(n9596) );
  NAND2_X1 U10765 ( .A1(n9596), .A2(n9595), .ZN(n9598) );
  OAI211_X1 U10766 ( .C1(n9600), .C2(n9599), .A(n9598), .B(n9597), .ZN(n9601)
         );
  INV_X1 U10767 ( .A(n9601), .ZN(n9608) );
  AOI21_X1 U10768 ( .B1(n9604), .B2(n9603), .A(n9602), .ZN(n9606) );
  OR2_X1 U10769 ( .A1(n9606), .A2(n9605), .ZN(n9607) );
  OAI211_X1 U10770 ( .C1(n10187), .C2(n9609), .A(n9608), .B(n9607), .ZN(
        P1_U3259) );
  INV_X1 U10771 ( .A(n9610), .ZN(n9675) );
  XNOR2_X1 U10772 ( .A(n9611), .B(n9612), .ZN(n9683) );
  XNOR2_X1 U10773 ( .A(n9613), .B(n9612), .ZN(n9618) );
  AOI22_X1 U10774 ( .A1(n9615), .A2(n6792), .B1(n9614), .B2(n9686), .ZN(n9616)
         );
  OAI21_X1 U10775 ( .B1(n9618), .B2(n9617), .A(n9616), .ZN(n9619) );
  AOI21_X1 U10776 ( .B1(n9675), .B2(n9683), .A(n9619), .ZN(n9680) );
  AOI222_X1 U10777 ( .A1(n9623), .A2(n9622), .B1(n9621), .B2(n9646), .C1(
        P1_REG2_REG_4__SCAN_IN), .C2(n9620), .ZN(n9632) );
  INV_X1 U10778 ( .A(n9625), .ZN(n9627) );
  OAI211_X1 U10779 ( .C1(n9679), .C2(n4588), .A(n9627), .B(n9626), .ZN(n9677)
         );
  INV_X1 U10780 ( .A(n9677), .ZN(n9628) );
  AOI22_X1 U10781 ( .A1(n9683), .A2(n9630), .B1(n9629), .B2(n9628), .ZN(n9631)
         );
  OAI211_X1 U10782 ( .C1(n9620), .C2(n9680), .A(n9632), .B(n9631), .ZN(
        P1_U3287) );
  NAND2_X1 U10783 ( .A1(n9634), .A2(n9633), .ZN(n9635) );
  OR2_X1 U10784 ( .A1(n9636), .A2(n9635), .ZN(n9638) );
  NAND2_X1 U10785 ( .A1(n7040), .A2(n9686), .ZN(n9637) );
  AND2_X1 U10786 ( .A1(n9638), .A2(n9637), .ZN(n9642) );
  INV_X1 U10787 ( .A(n9642), .ZN(n9645) );
  NAND2_X1 U10788 ( .A1(n9640), .A2(n9639), .ZN(n9641) );
  AND2_X1 U10789 ( .A1(n9642), .A2(n9641), .ZN(n9722) );
  INV_X1 U10790 ( .A(n9722), .ZN(n9643) );
  OAI21_X1 U10791 ( .B1(n9645), .B2(n9644), .A(n9643), .ZN(n9648) );
  AOI22_X1 U10792 ( .A1(P1_REG3_REG_0__SCAN_IN), .A2(n9646), .B1(
        P1_REG2_REG_0__SCAN_IN), .B2(n9620), .ZN(n9647) );
  OAI21_X1 U10793 ( .B1(n9620), .B2(n9648), .A(n9647), .ZN(P1_U3291) );
  AND2_X1 U10794 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9651), .ZN(P1_U3292) );
  AND2_X1 U10795 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9651), .ZN(P1_U3293) );
  AND2_X1 U10796 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9651), .ZN(P1_U3294) );
  AND2_X1 U10797 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9651), .ZN(P1_U3295) );
  AND2_X1 U10798 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9651), .ZN(P1_U3296) );
  AND2_X1 U10799 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9651), .ZN(P1_U3297) );
  AND2_X1 U10800 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9651), .ZN(P1_U3298) );
  AND2_X1 U10801 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9651), .ZN(P1_U3299) );
  AND2_X1 U10802 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9651), .ZN(P1_U3300) );
  AND2_X1 U10803 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9651), .ZN(P1_U3301) );
  AND2_X1 U10804 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9651), .ZN(P1_U3302) );
  AND2_X1 U10805 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9651), .ZN(P1_U3303) );
  AND2_X1 U10806 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9651), .ZN(P1_U3304) );
  AND2_X1 U10807 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9651), .ZN(P1_U3305) );
  AND2_X1 U10808 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9651), .ZN(P1_U3306) );
  AND2_X1 U10809 ( .A1(n9651), .A2(P1_D_REG_16__SCAN_IN), .ZN(P1_U3307) );
  AND2_X1 U10810 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9651), .ZN(P1_U3308) );
  INV_X1 U10811 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n10146) );
  NOR2_X1 U10812 ( .A1(n9650), .A2(n10146), .ZN(P1_U3309) );
  INV_X1 U10813 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n10064) );
  NOR2_X1 U10814 ( .A1(n9650), .A2(n10064), .ZN(P1_U3310) );
  AND2_X1 U10815 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9651), .ZN(P1_U3311) );
  INV_X1 U10816 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n10149) );
  NOR2_X1 U10817 ( .A1(n9650), .A2(n10149), .ZN(P1_U3312) );
  AND2_X1 U10818 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9651), .ZN(P1_U3313) );
  AND2_X1 U10819 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9651), .ZN(P1_U3314) );
  AND2_X1 U10820 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9651), .ZN(P1_U3315) );
  INV_X1 U10821 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n10141) );
  NOR2_X1 U10822 ( .A1(n9650), .A2(n10141), .ZN(P1_U3316) );
  AND2_X1 U10823 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9651), .ZN(P1_U3317) );
  AND2_X1 U10824 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9651), .ZN(P1_U3318) );
  AND2_X1 U10825 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n9651), .ZN(P1_U3319) );
  AND2_X1 U10826 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9651), .ZN(P1_U3320) );
  AND2_X1 U10827 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9651), .ZN(P1_U3321) );
  INV_X1 U10828 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n9653) );
  OAI21_X1 U10829 ( .B1(n9654), .B2(n9653), .A(n9652), .ZN(P1_U3441) );
  AOI22_X1 U10830 ( .A1(n9720), .A2(n9722), .B1(n5769), .B2(n9718), .ZN(
        P1_U3454) );
  OAI211_X1 U10831 ( .C1(n9657), .C2(n9712), .A(n9656), .B(n9655), .ZN(n9658)
         );
  NOR2_X1 U10832 ( .A1(n9659), .A2(n9658), .ZN(n9723) );
  AOI22_X1 U10833 ( .A1(n9720), .A2(n9723), .B1(n5786), .B2(n9718), .ZN(
        P1_U3457) );
  AOI22_X1 U10834 ( .A1(n6792), .A2(n9686), .B1(n9695), .B2(n9660), .ZN(n9663)
         );
  NAND2_X1 U10835 ( .A1(n9666), .A2(n9684), .ZN(n9662) );
  NAND4_X1 U10836 ( .A1(n9664), .A2(n9663), .A3(n9662), .A4(n9661), .ZN(n9665)
         );
  AOI21_X1 U10837 ( .B1(n9675), .B2(n9666), .A(n9665), .ZN(n9725) );
  AOI22_X1 U10838 ( .A1(n9720), .A2(n9725), .B1(n5802), .B2(n9718), .ZN(
        P1_U3460) );
  INV_X1 U10839 ( .A(n9671), .ZN(n9674) );
  AOI22_X1 U10840 ( .A1(n9668), .A2(n9686), .B1(n9695), .B2(n9667), .ZN(n9670)
         );
  OAI211_X1 U10841 ( .C1(n9671), .C2(n9712), .A(n9670), .B(n9669), .ZN(n9672)
         );
  AOI211_X1 U10842 ( .C1(n9675), .C2(n9674), .A(n9673), .B(n9672), .ZN(n9726)
         );
  INV_X1 U10843 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n9676) );
  AOI22_X1 U10844 ( .A1(n9720), .A2(n9726), .B1(n9676), .B2(n9718), .ZN(
        P1_U3463) );
  OAI21_X1 U10845 ( .B1(n9679), .B2(n9678), .A(n9677), .ZN(n9682) );
  INV_X1 U10846 ( .A(n9680), .ZN(n9681) );
  AOI211_X1 U10847 ( .C1(n9684), .C2(n9683), .A(n9682), .B(n9681), .ZN(n9727)
         );
  AOI22_X1 U10848 ( .A1(n9720), .A2(n9727), .B1(n5828), .B2(n9718), .ZN(
        P1_U3466) );
  AOI22_X1 U10849 ( .A1(n9687), .A2(n9686), .B1(n9695), .B2(n9685), .ZN(n9691)
         );
  NAND3_X1 U10850 ( .A1(n7260), .A2(n9688), .A3(n9710), .ZN(n9690) );
  AOI22_X1 U10851 ( .A1(n9720), .A2(n9728), .B1(n5844), .B2(n9718), .ZN(
        P1_U3469) );
  AOI21_X1 U10852 ( .B1(n9695), .B2(n9694), .A(n9693), .ZN(n9696) );
  OAI211_X1 U10853 ( .C1(n9699), .C2(n9698), .A(n9697), .B(n9696), .ZN(n9700)
         );
  INV_X1 U10854 ( .A(n9700), .ZN(n9729) );
  INV_X1 U10855 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9701) );
  AOI22_X1 U10856 ( .A1(n9720), .A2(n9729), .B1(n9701), .B2(n9718), .ZN(
        P1_U3472) );
  INV_X1 U10857 ( .A(n9702), .ZN(n9703) );
  OAI211_X1 U10858 ( .C1(n9706), .C2(n9705), .A(n9704), .B(n9703), .ZN(n9708)
         );
  AOI211_X1 U10859 ( .C1(n9710), .C2(n9709), .A(n9708), .B(n9707), .ZN(n9730)
         );
  INV_X1 U10860 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9711) );
  AOI22_X1 U10861 ( .A1(n9720), .A2(n9730), .B1(n9711), .B2(n9718), .ZN(
        P1_U3475) );
  NOR2_X1 U10862 ( .A1(n9713), .A2(n9712), .ZN(n9716) );
  NOR4_X1 U10863 ( .A1(n9717), .A2(n9716), .A3(n9715), .A4(n9714), .ZN(n9732)
         );
  INV_X1 U10864 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n9719) );
  AOI22_X1 U10865 ( .A1(n9720), .A2(n9732), .B1(n9719), .B2(n9718), .ZN(
        P1_U3478) );
  AOI22_X1 U10866 ( .A1(n9733), .A2(n9722), .B1(n9721), .B2(n9731), .ZN(
        P1_U3523) );
  AOI22_X1 U10867 ( .A1(n9733), .A2(n9723), .B1(n6305), .B2(n9731), .ZN(
        P1_U3524) );
  AOI22_X1 U10868 ( .A1(n9733), .A2(n9725), .B1(n9724), .B2(n9731), .ZN(
        P1_U3525) );
  AOI22_X1 U10869 ( .A1(n9733), .A2(n9726), .B1(n6304), .B2(n9731), .ZN(
        P1_U3526) );
  AOI22_X1 U10870 ( .A1(n9733), .A2(n9727), .B1(n5824), .B2(n9731), .ZN(
        P1_U3527) );
  AOI22_X1 U10871 ( .A1(n9733), .A2(n9728), .B1(n6303), .B2(n9731), .ZN(
        P1_U3528) );
  AOI22_X1 U10872 ( .A1(n9733), .A2(n9729), .B1(n5863), .B2(n9731), .ZN(
        P1_U3529) );
  AOI22_X1 U10873 ( .A1(n9733), .A2(n9730), .B1(n5877), .B2(n9731), .ZN(
        P1_U3530) );
  AOI22_X1 U10874 ( .A1(n9733), .A2(n9732), .B1(n6302), .B2(n9731), .ZN(
        P1_U3531) );
  AOI22_X1 U10875 ( .A1(n9783), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n9786), .ZN(n9741) );
  AOI22_X1 U10876 ( .A1(n9781), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n9740) );
  OAI21_X1 U10877 ( .B1(n9735), .B2(P2_REG1_REG_0__SCAN_IN), .A(n9734), .ZN(
        n9738) );
  NOR2_X1 U10878 ( .A1(n9736), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n9737) );
  OAI21_X1 U10879 ( .B1(n9738), .B2(n9737), .A(P2_IR_REG_0__SCAN_IN), .ZN(
        n9739) );
  OAI211_X1 U10880 ( .C1(P2_IR_REG_0__SCAN_IN), .C2(n9741), .A(n9740), .B(
        n9739), .ZN(P2_U3245) );
  INV_X1 U10881 ( .A(n9742), .ZN(n9743) );
  AOI21_X1 U10882 ( .B1(n9781), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n9743), .ZN(
        n9754) );
  NAND2_X1 U10883 ( .A1(n9791), .A2(n9744), .ZN(n9753) );
  OAI211_X1 U10884 ( .C1(n9747), .C2(n9746), .A(n9786), .B(n9745), .ZN(n9752)
         );
  OAI211_X1 U10885 ( .C1(n9750), .C2(n9749), .A(n9783), .B(n9748), .ZN(n9751)
         );
  NAND4_X1 U10886 ( .A1(n9754), .A2(n9753), .A3(n9752), .A4(n9751), .ZN(
        P2_U3248) );
  INV_X1 U10887 ( .A(n9755), .ZN(n9756) );
  AOI21_X1 U10888 ( .B1(n9781), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n9756), .ZN(
        n9767) );
  NAND2_X1 U10889 ( .A1(n9791), .A2(n9757), .ZN(n9766) );
  OAI211_X1 U10890 ( .C1(n9760), .C2(n9759), .A(n9786), .B(n9758), .ZN(n9765)
         );
  OAI211_X1 U10891 ( .C1(n9763), .C2(n9762), .A(n9783), .B(n9761), .ZN(n9764)
         );
  NAND4_X1 U10892 ( .A1(n9767), .A2(n9766), .A3(n9765), .A4(n9764), .ZN(
        P2_U3252) );
  INV_X1 U10893 ( .A(n9768), .ZN(n9769) );
  AOI21_X1 U10894 ( .B1(n9781), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n9769), .ZN(
        n9780) );
  NAND2_X1 U10895 ( .A1(n9791), .A2(n9770), .ZN(n9779) );
  OAI211_X1 U10896 ( .C1(n9773), .C2(n9772), .A(n9786), .B(n9771), .ZN(n9778)
         );
  OAI211_X1 U10897 ( .C1(n9776), .C2(n9775), .A(n9783), .B(n9774), .ZN(n9777)
         );
  NAND4_X1 U10898 ( .A1(n9780), .A2(n9779), .A3(n9778), .A4(n9777), .ZN(
        P2_U3255) );
  AOI22_X1 U10899 ( .A1(n9781), .A2(P2_ADDR_REG_17__SCAN_IN), .B1(
        P2_REG3_REG_17__SCAN_IN), .B2(P2_U3152), .ZN(n9795) );
  OAI211_X1 U10900 ( .C1(n9785), .C2(n9784), .A(n9783), .B(n9782), .ZN(n9794)
         );
  OAI211_X1 U10901 ( .C1(n9789), .C2(n9788), .A(n9787), .B(n9786), .ZN(n9793)
         );
  NAND2_X1 U10902 ( .A1(n9791), .A2(n9790), .ZN(n9792) );
  NAND4_X1 U10903 ( .A1(n9795), .A2(n9794), .A3(n9793), .A4(n9792), .ZN(
        P2_U3262) );
  OR2_X1 U10904 ( .A1(n7433), .A2(n9796), .ZN(n9798) );
  NAND2_X1 U10905 ( .A1(n9798), .A2(n9797), .ZN(n9801) );
  OAI211_X1 U10906 ( .C1(n9801), .C2(n9800), .A(n9799), .B(n9818), .ZN(n9803)
         );
  AND2_X1 U10907 ( .A1(n9803), .A2(n9802), .ZN(n9936) );
  AOI222_X1 U10908 ( .A1(n9809), .A2(n9856), .B1(P2_REG2_REG_12__SCAN_IN), 
        .B2(n9855), .C1(n9854), .C2(n9804), .ZN(n9815) );
  INV_X1 U10909 ( .A(n9805), .ZN(n9808) );
  OAI21_X1 U10910 ( .B1(n9808), .B2(n9807), .A(n9806), .ZN(n9940) );
  AOI21_X1 U10911 ( .B1(n9810), .B2(n9809), .A(n6682), .ZN(n9812) );
  NAND2_X1 U10912 ( .A1(n9812), .A2(n9811), .ZN(n9935) );
  INV_X1 U10913 ( .A(n9935), .ZN(n9813) );
  AOI22_X1 U10914 ( .A1(n9940), .A2(n9834), .B1(n9862), .B2(n9813), .ZN(n9814)
         );
  OAI211_X1 U10915 ( .C1(n9866), .C2(n9936), .A(n9815), .B(n9814), .ZN(
        P2_U3284) );
  NAND2_X1 U10916 ( .A1(n7433), .A2(n9816), .ZN(n9817) );
  NAND3_X1 U10917 ( .A1(n9819), .A2(n9818), .A3(n9817), .ZN(n9821) );
  AND2_X1 U10918 ( .A1(n9821), .A2(n9820), .ZN(n9922) );
  AOI222_X1 U10919 ( .A1(n9823), .A2(n9856), .B1(P2_REG2_REG_10__SCAN_IN), 
        .B2(n9855), .C1(n9854), .C2(n9822), .ZN(n9836) );
  NAND2_X1 U10920 ( .A1(n9825), .A2(n9824), .ZN(n9827) );
  OR2_X1 U10921 ( .A1(n9827), .A2(n9826), .ZN(n9829) );
  NAND2_X1 U10922 ( .A1(n9827), .A2(n9826), .ZN(n9828) );
  AND2_X1 U10923 ( .A1(n9829), .A2(n9828), .ZN(n9925) );
  OAI211_X1 U10924 ( .C1(n9831), .C2(n9923), .A(n7321), .B(n9830), .ZN(n9921)
         );
  NOR2_X1 U10925 ( .A1(n9921), .A2(n9832), .ZN(n9833) );
  AOI21_X1 U10926 ( .B1(n9925), .B2(n9834), .A(n9833), .ZN(n9835) );
  OAI211_X1 U10927 ( .C1(n9866), .C2(n9922), .A(n9836), .B(n9835), .ZN(
        P2_U3286) );
  INV_X1 U10928 ( .A(n9837), .ZN(n9838) );
  AOI21_X1 U10929 ( .B1(n9840), .B2(n9839), .A(n9838), .ZN(n9913) );
  NAND2_X1 U10930 ( .A1(n9842), .A2(n9841), .ZN(n9844) );
  AOI21_X1 U10931 ( .B1(n9845), .B2(n9844), .A(n9843), .ZN(n9851) );
  OAI22_X1 U10932 ( .A1(n9849), .A2(n9848), .B1(n9847), .B2(n9846), .ZN(n9850)
         );
  AOI211_X1 U10933 ( .C1(n9913), .C2(n9852), .A(n9851), .B(n9850), .ZN(n9910)
         );
  AOI222_X1 U10934 ( .A1(n9857), .A2(n9856), .B1(P2_REG2_REG_8__SCAN_IN), .B2(
        n9855), .C1(n9854), .C2(n9853), .ZN(n9865) );
  INV_X1 U10935 ( .A(n9859), .ZN(n9860) );
  OAI211_X1 U10936 ( .C1(n4563), .C2(n4560), .A(n9860), .B(n7321), .ZN(n9909)
         );
  INV_X1 U10937 ( .A(n9909), .ZN(n9861) );
  AOI22_X1 U10938 ( .A1(n9913), .A2(n9863), .B1(n9862), .B2(n9861), .ZN(n9864)
         );
  OAI211_X1 U10939 ( .C1(n9866), .C2(n9910), .A(n9865), .B(n9864), .ZN(
        P2_U3288) );
  NOR2_X1 U10940 ( .A1(n9868), .A2(n9867), .ZN(n9874) );
  AND2_X1 U10941 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n9989), .ZN(P2_U3297) );
  AND2_X1 U10942 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n9989), .ZN(P2_U3298) );
  AND2_X1 U10943 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n9989), .ZN(P2_U3299) );
  AND2_X1 U10944 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n9989), .ZN(P2_U3300) );
  AND2_X1 U10945 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n9989), .ZN(P2_U3301) );
  AND2_X1 U10946 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n9989), .ZN(P2_U3303) );
  AND2_X1 U10947 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n9989), .ZN(P2_U3304) );
  AND2_X1 U10948 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n9989), .ZN(P2_U3305) );
  INV_X1 U10949 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n10144) );
  NOR2_X1 U10950 ( .A1(n9874), .A2(n10144), .ZN(P2_U3306) );
  AND2_X1 U10951 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n9989), .ZN(P2_U3307) );
  AND2_X1 U10952 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n9989), .ZN(P2_U3308) );
  AND2_X1 U10953 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n9989), .ZN(P2_U3309) );
  AND2_X1 U10954 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n9989), .ZN(P2_U3310) );
  AND2_X1 U10955 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n9989), .ZN(P2_U3311) );
  AND2_X1 U10956 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n9989), .ZN(P2_U3312) );
  AND2_X1 U10957 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n9989), .ZN(P2_U3313) );
  AND2_X1 U10958 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n9989), .ZN(P2_U3314) );
  AND2_X1 U10959 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n9989), .ZN(P2_U3315) );
  AND2_X1 U10960 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n9989), .ZN(P2_U3316) );
  AND2_X1 U10961 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n9989), .ZN(P2_U3317) );
  AND2_X1 U10962 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n9989), .ZN(P2_U3318) );
  AND2_X1 U10963 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n9989), .ZN(P2_U3319) );
  AND2_X1 U10964 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n9989), .ZN(P2_U3320) );
  AND2_X1 U10965 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n9989), .ZN(P2_U3321) );
  AND2_X1 U10966 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n9989), .ZN(P2_U3322) );
  AND2_X1 U10967 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n9989), .ZN(P2_U3323) );
  AND2_X1 U10968 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n9989), .ZN(P2_U3324) );
  AND2_X1 U10969 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n9989), .ZN(P2_U3325) );
  AND2_X1 U10970 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n9989), .ZN(P2_U3326) );
  NAND2_X1 U10971 ( .A1(n9870), .A2(n9869), .ZN(n9872) );
  NAND2_X1 U10972 ( .A1(n9871), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9875) );
  OAI22_X1 U10973 ( .A1(n9872), .A2(n9875), .B1(P2_D_REG_0__SCAN_IN), .B2(
        n9874), .ZN(n9873) );
  INV_X1 U10974 ( .A(n9873), .ZN(P2_U3437) );
  OAI22_X1 U10975 ( .A1(n9876), .A2(n9875), .B1(P2_D_REG_1__SCAN_IN), .B2(
        n9874), .ZN(n9877) );
  INV_X1 U10976 ( .A(n9877), .ZN(P2_U3438) );
  INV_X1 U10977 ( .A(n9878), .ZN(n9883) );
  OAI22_X1 U10978 ( .A1(n9881), .A2(n9932), .B1(n9880), .B2(n9879), .ZN(n9882)
         );
  NOR2_X1 U10979 ( .A1(n9883), .A2(n9882), .ZN(n9945) );
  INV_X1 U10980 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n9884) );
  AOI22_X1 U10981 ( .A1(n9944), .A2(n9945), .B1(n9884), .B2(n9942), .ZN(
        P2_U3451) );
  OAI211_X1 U10982 ( .C1(n9887), .C2(n9937), .A(n9886), .B(n9885), .ZN(n9888)
         );
  AOI21_X1 U10983 ( .B1(n9889), .B2(n9941), .A(n9888), .ZN(n9946) );
  INV_X1 U10984 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10164) );
  AOI22_X1 U10985 ( .A1(n9944), .A2(n9946), .B1(n10164), .B2(n9942), .ZN(
        P2_U3457) );
  OAI21_X1 U10986 ( .B1(n9891), .B2(n9937), .A(n9890), .ZN(n9893) );
  AOI211_X1 U10987 ( .C1(n9941), .C2(n9894), .A(n9893), .B(n9892), .ZN(n9947)
         );
  INV_X1 U10988 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n9895) );
  AOI22_X1 U10989 ( .A1(n9944), .A2(n9947), .B1(n9895), .B2(n9942), .ZN(
        P2_U3463) );
  AOI21_X1 U10990 ( .B1(n9927), .B2(n9897), .A(n9896), .ZN(n9898) );
  OAI211_X1 U10991 ( .C1(n9900), .C2(n9932), .A(n9899), .B(n9898), .ZN(n9901)
         );
  INV_X1 U10992 ( .A(n9901), .ZN(n9948) );
  INV_X1 U10993 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n9902) );
  AOI22_X1 U10994 ( .A1(n9944), .A2(n9948), .B1(n9902), .B2(n9942), .ZN(
        P2_U3469) );
  OAI21_X1 U10995 ( .B1(n9904), .B2(n9937), .A(n9903), .ZN(n9906) );
  AOI211_X1 U10996 ( .C1(n9907), .C2(n9941), .A(n9906), .B(n9905), .ZN(n9949)
         );
  INV_X1 U10997 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n9908) );
  AOI22_X1 U10998 ( .A1(n9944), .A2(n9949), .B1(n9908), .B2(n9942), .ZN(
        P2_U3472) );
  OAI21_X1 U10999 ( .B1(n4563), .B2(n9937), .A(n9909), .ZN(n9912) );
  INV_X1 U11000 ( .A(n9910), .ZN(n9911) );
  AOI211_X1 U11001 ( .C1(n9920), .C2(n9913), .A(n9912), .B(n9911), .ZN(n9951)
         );
  INV_X1 U11002 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n9914) );
  AOI22_X1 U11003 ( .A1(n9944), .A2(n9951), .B1(n9914), .B2(n9942), .ZN(
        P2_U3475) );
  OAI22_X1 U11004 ( .A1(n9916), .A2(n6682), .B1(n9915), .B2(n9937), .ZN(n9918)
         );
  AOI211_X1 U11005 ( .C1(n9920), .C2(n9919), .A(n9918), .B(n9917), .ZN(n9953)
         );
  INV_X1 U11006 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10147) );
  AOI22_X1 U11007 ( .A1(n9944), .A2(n9953), .B1(n10147), .B2(n9942), .ZN(
        P2_U3478) );
  OAI211_X1 U11008 ( .C1(n9923), .C2(n9937), .A(n9922), .B(n9921), .ZN(n9924)
         );
  AOI21_X1 U11009 ( .B1(n9925), .B2(n9941), .A(n9924), .ZN(n9954) );
  AOI22_X1 U11010 ( .A1(n9944), .A2(n9954), .B1(n5168), .B2(n9942), .ZN(
        P2_U3481) );
  AOI22_X1 U11011 ( .A1(n9928), .A2(n7321), .B1(n9927), .B2(n9926), .ZN(n9929)
         );
  OAI211_X1 U11012 ( .C1(n9932), .C2(n9931), .A(n9930), .B(n9929), .ZN(n9933)
         );
  INV_X1 U11013 ( .A(n9933), .ZN(n9955) );
  INV_X1 U11014 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n9934) );
  AOI22_X1 U11015 ( .A1(n9944), .A2(n9955), .B1(n9934), .B2(n9942), .ZN(
        P2_U3484) );
  OAI211_X1 U11016 ( .C1(n9938), .C2(n9937), .A(n9936), .B(n9935), .ZN(n9939)
         );
  AOI21_X1 U11017 ( .B1(n9941), .B2(n9940), .A(n9939), .ZN(n9958) );
  INV_X1 U11018 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n9943) );
  AOI22_X1 U11019 ( .A1(n9944), .A2(n9958), .B1(n9943), .B2(n9942), .ZN(
        P2_U3487) );
  AOI22_X1 U11020 ( .A1(n9959), .A2(n9945), .B1(n6401), .B2(n9956), .ZN(
        P2_U3520) );
  AOI22_X1 U11021 ( .A1(n9959), .A2(n9946), .B1(n6403), .B2(n9956), .ZN(
        P2_U3522) );
  AOI22_X1 U11022 ( .A1(n9959), .A2(n9947), .B1(n6406), .B2(n9956), .ZN(
        P2_U3524) );
  AOI22_X1 U11023 ( .A1(n9959), .A2(n9948), .B1(n6410), .B2(n9956), .ZN(
        P2_U3526) );
  AOI22_X1 U11024 ( .A1(n9959), .A2(n9949), .B1(n6464), .B2(n9956), .ZN(
        P2_U3527) );
  AOI22_X1 U11025 ( .A1(n9959), .A2(n9951), .B1(n9950), .B2(n9956), .ZN(
        P2_U3528) );
  AOI22_X1 U11026 ( .A1(n9959), .A2(n9953), .B1(n9952), .B2(n9956), .ZN(
        P2_U3529) );
  AOI22_X1 U11027 ( .A1(n9959), .A2(n9954), .B1(n6463), .B2(n9956), .ZN(
        P2_U3530) );
  AOI22_X1 U11028 ( .A1(n9959), .A2(n9955), .B1(n6471), .B2(n9956), .ZN(
        P2_U3531) );
  AOI22_X1 U11029 ( .A1(n9959), .A2(n9958), .B1(n9957), .B2(n9956), .ZN(
        P2_U3532) );
  INV_X1 U11030 ( .A(n9960), .ZN(n9961) );
  NAND2_X1 U11031 ( .A1(n9962), .A2(n9961), .ZN(n9963) );
  XOR2_X1 U11032 ( .A(n9964), .B(n9963), .Z(ADD_1071_U5) );
  XOR2_X1 U11033 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  OAI21_X1 U11034 ( .B1(n9967), .B2(n9966), .A(n9965), .ZN(ADD_1071_U56) );
  OAI21_X1 U11035 ( .B1(n9970), .B2(n9969), .A(n9968), .ZN(ADD_1071_U57) );
  OAI21_X1 U11036 ( .B1(n9973), .B2(n9972), .A(n9971), .ZN(ADD_1071_U58) );
  OAI21_X1 U11037 ( .B1(n9976), .B2(n9975), .A(n9974), .ZN(ADD_1071_U59) );
  OAI21_X1 U11038 ( .B1(n9979), .B2(n9978), .A(n9977), .ZN(ADD_1071_U60) );
  OAI21_X1 U11039 ( .B1(n9982), .B2(n9981), .A(n9980), .ZN(ADD_1071_U61) );
  AOI21_X1 U11040 ( .B1(n9985), .B2(n9984), .A(n9983), .ZN(ADD_1071_U62) );
  AOI21_X1 U11041 ( .B1(n9988), .B2(n9987), .A(n9986), .ZN(ADD_1071_U63) );
  NAND2_X1 U11042 ( .A1(n9989), .A2(P2_D_REG_26__SCAN_IN), .ZN(n10178) );
  INV_X1 U11043 ( .A(SI_21_), .ZN(n10067) );
  OAI22_X1 U11044 ( .A1(n10067), .A2(keyinput23), .B1(n5844), .B2(keyinput24), 
        .ZN(n9990) );
  AOI221_X1 U11045 ( .B1(n10067), .B2(keyinput23), .C1(keyinput24), .C2(n5844), 
        .A(n9990), .ZN(n10001) );
  XNOR2_X1 U11046 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(keyinput62), .ZN(n9994) );
  XNOR2_X1 U11047 ( .A(P2_IR_REG_0__SCAN_IN), .B(keyinput29), .ZN(n9993) );
  XNOR2_X1 U11048 ( .A(P1_IR_REG_30__SCAN_IN), .B(keyinput8), .ZN(n9992) );
  XNOR2_X1 U11049 ( .A(P2_IR_REG_29__SCAN_IN), .B(keyinput55), .ZN(n9991) );
  NAND4_X1 U11050 ( .A1(n9994), .A2(n9993), .A3(n9992), .A4(n9991), .ZN(n9999)
         );
  XNOR2_X1 U11051 ( .A(n9995), .B(keyinput17), .ZN(n9998) );
  INV_X1 U11052 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n9996) );
  XNOR2_X1 U11053 ( .A(keyinput15), .B(n9996), .ZN(n9997) );
  NOR3_X1 U11054 ( .A1(n9999), .A2(n9998), .A3(n9997), .ZN(n10000) );
  NAND2_X1 U11055 ( .A1(n10001), .A2(n10000), .ZN(n10176) );
  INV_X1 U11056 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n10003) );
  OAI22_X1 U11057 ( .A1(n10004), .A2(keyinput1), .B1(n10003), .B2(keyinput7), 
        .ZN(n10002) );
  AOI221_X1 U11058 ( .B1(n10004), .B2(keyinput1), .C1(keyinput7), .C2(n10003), 
        .A(n10002), .ZN(n10012) );
  OAI22_X1 U11059 ( .A1(n10006), .A2(keyinput10), .B1(n10075), .B2(keyinput52), 
        .ZN(n10005) );
  AOI221_X1 U11060 ( .B1(n10006), .B2(keyinput10), .C1(keyinput52), .C2(n10075), .A(n10005), .ZN(n10011) );
  OAI22_X1 U11061 ( .A1(n10062), .A2(keyinput43), .B1(n10089), .B2(keyinput44), 
        .ZN(n10007) );
  AOI221_X1 U11062 ( .B1(n10062), .B2(keyinput43), .C1(keyinput44), .C2(n10089), .A(n10007), .ZN(n10010) );
  OAI22_X1 U11063 ( .A1(n10064), .A2(keyinput42), .B1(n10077), .B2(keyinput56), 
        .ZN(n10008) );
  AOI221_X1 U11064 ( .B1(n10064), .B2(keyinput42), .C1(keyinput56), .C2(n10077), .A(n10008), .ZN(n10009) );
  NAND4_X1 U11065 ( .A1(n10012), .A2(n10011), .A3(n10010), .A4(n10009), .ZN(
        n10175) );
  AOI22_X1 U11066 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(keyinput9), .B1(
        P1_REG0_REG_23__SCAN_IN), .B2(keyinput19), .ZN(n10013) );
  OAI221_X1 U11067 ( .B1(P2_REG3_REG_14__SCAN_IN), .B2(keyinput9), .C1(
        P1_REG0_REG_23__SCAN_IN), .C2(keyinput19), .A(n10013), .ZN(n10020) );
  AOI22_X1 U11068 ( .A1(P1_ADDR_REG_14__SCAN_IN), .A2(keyinput11), .B1(
        P2_IR_REG_15__SCAN_IN), .B2(keyinput0), .ZN(n10014) );
  OAI221_X1 U11069 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(keyinput11), .C1(
        P2_IR_REG_15__SCAN_IN), .C2(keyinput0), .A(n10014), .ZN(n10019) );
  AOI22_X1 U11070 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(keyinput13), .B1(
        P1_REG3_REG_11__SCAN_IN), .B2(keyinput22), .ZN(n10015) );
  OAI221_X1 U11071 ( .B1(P2_IR_REG_31__SCAN_IN), .B2(keyinput13), .C1(
        P1_REG3_REG_11__SCAN_IN), .C2(keyinput22), .A(n10015), .ZN(n10018) );
  AOI22_X1 U11072 ( .A1(P1_REG0_REG_10__SCAN_IN), .A2(keyinput51), .B1(
        P1_REG0_REG_26__SCAN_IN), .B2(keyinput49), .ZN(n10016) );
  OAI221_X1 U11073 ( .B1(P1_REG0_REG_10__SCAN_IN), .B2(keyinput51), .C1(
        P1_REG0_REG_26__SCAN_IN), .C2(keyinput49), .A(n10016), .ZN(n10017) );
  NOR4_X1 U11074 ( .A1(n10020), .A2(n10019), .A3(n10018), .A4(n10017), .ZN(
        n10048) );
  AOI22_X1 U11075 ( .A1(P1_REG0_REG_31__SCAN_IN), .A2(keyinput16), .B1(
        P1_REG0_REG_13__SCAN_IN), .B2(keyinput27), .ZN(n10021) );
  OAI221_X1 U11076 ( .B1(P1_REG0_REG_31__SCAN_IN), .B2(keyinput16), .C1(
        P1_REG0_REG_13__SCAN_IN), .C2(keyinput27), .A(n10021), .ZN(n10028) );
  AOI22_X1 U11077 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(keyinput61), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(keyinput26), .ZN(n10022) );
  OAI221_X1 U11078 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(keyinput61), .C1(
        P2_DATAO_REG_25__SCAN_IN), .C2(keyinput26), .A(n10022), .ZN(n10027) );
  AOI22_X1 U11079 ( .A1(P2_REG0_REG_10__SCAN_IN), .A2(keyinput60), .B1(
        P2_IR_REG_16__SCAN_IN), .B2(keyinput57), .ZN(n10023) );
  OAI221_X1 U11080 ( .B1(P2_REG0_REG_10__SCAN_IN), .B2(keyinput60), .C1(
        P2_IR_REG_16__SCAN_IN), .C2(keyinput57), .A(n10023), .ZN(n10026) );
  AOI22_X1 U11081 ( .A1(P1_REG2_REG_3__SCAN_IN), .A2(keyinput4), .B1(
        P1_REG0_REG_16__SCAN_IN), .B2(keyinput37), .ZN(n10024) );
  OAI221_X1 U11082 ( .B1(P1_REG2_REG_3__SCAN_IN), .B2(keyinput4), .C1(
        P1_REG0_REG_16__SCAN_IN), .C2(keyinput37), .A(n10024), .ZN(n10025) );
  NOR4_X1 U11083 ( .A1(n10028), .A2(n10027), .A3(n10026), .A4(n10025), .ZN(
        n10047) );
  AOI22_X1 U11084 ( .A1(P2_REG1_REG_11__SCAN_IN), .A2(keyinput36), .B1(
        P2_REG3_REG_12__SCAN_IN), .B2(keyinput63), .ZN(n10029) );
  OAI221_X1 U11085 ( .B1(P2_REG1_REG_11__SCAN_IN), .B2(keyinput36), .C1(
        P2_REG3_REG_12__SCAN_IN), .C2(keyinput63), .A(n10029), .ZN(n10036) );
  AOI22_X1 U11086 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(keyinput14), .B1(
        P1_REG3_REG_17__SCAN_IN), .B2(keyinput41), .ZN(n10030) );
  OAI221_X1 U11087 ( .B1(P2_REG3_REG_11__SCAN_IN), .B2(keyinput14), .C1(
        P1_REG3_REG_17__SCAN_IN), .C2(keyinput41), .A(n10030), .ZN(n10035) );
  AOI22_X1 U11088 ( .A1(P1_REG1_REG_28__SCAN_IN), .A2(keyinput20), .B1(
        P1_IR_REG_16__SCAN_IN), .B2(keyinput53), .ZN(n10031) );
  OAI221_X1 U11089 ( .B1(P1_REG1_REG_28__SCAN_IN), .B2(keyinput20), .C1(
        P1_IR_REG_16__SCAN_IN), .C2(keyinput53), .A(n10031), .ZN(n10034) );
  AOI22_X1 U11090 ( .A1(P1_REG0_REG_28__SCAN_IN), .A2(keyinput47), .B1(
        P2_ADDR_REG_19__SCAN_IN), .B2(keyinput58), .ZN(n10032) );
  OAI221_X1 U11091 ( .B1(P1_REG0_REG_28__SCAN_IN), .B2(keyinput47), .C1(
        P2_ADDR_REG_19__SCAN_IN), .C2(keyinput58), .A(n10032), .ZN(n10033) );
  NOR4_X1 U11092 ( .A1(n10036), .A2(n10035), .A3(n10034), .A4(n10033), .ZN(
        n10046) );
  AOI22_X1 U11093 ( .A1(P2_REG2_REG_26__SCAN_IN), .A2(keyinput32), .B1(
        P2_REG1_REG_31__SCAN_IN), .B2(keyinput33), .ZN(n10037) );
  OAI221_X1 U11094 ( .B1(P2_REG2_REG_26__SCAN_IN), .B2(keyinput32), .C1(
        P2_REG1_REG_31__SCAN_IN), .C2(keyinput33), .A(n10037), .ZN(n10044) );
  AOI22_X1 U11095 ( .A1(P2_REG0_REG_6__SCAN_IN), .A2(keyinput6), .B1(
        P1_REG2_REG_18__SCAN_IN), .B2(keyinput12), .ZN(n10038) );
  OAI221_X1 U11096 ( .B1(P2_REG0_REG_6__SCAN_IN), .B2(keyinput6), .C1(
        P1_REG2_REG_18__SCAN_IN), .C2(keyinput12), .A(n10038), .ZN(n10043) );
  AOI22_X1 U11097 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(keyinput34), .B1(
        P2_REG2_REG_10__SCAN_IN), .B2(keyinput39), .ZN(n10039) );
  OAI221_X1 U11098 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(keyinput34), .C1(
        P2_REG2_REG_10__SCAN_IN), .C2(keyinput39), .A(n10039), .ZN(n10042) );
  AOI22_X1 U11099 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(keyinput54), .B1(
        P1_DATAO_REG_21__SCAN_IN), .B2(keyinput25), .ZN(n10040) );
  OAI221_X1 U11100 ( .B1(P2_REG3_REG_19__SCAN_IN), .B2(keyinput54), .C1(
        P1_DATAO_REG_21__SCAN_IN), .C2(keyinput25), .A(n10040), .ZN(n10041) );
  NOR4_X1 U11101 ( .A1(n10044), .A2(n10043), .A3(n10042), .A4(n10041), .ZN(
        n10045) );
  NAND4_X1 U11102 ( .A1(n10048), .A2(n10047), .A3(n10046), .A4(n10045), .ZN(
        n10174) );
  AOI22_X1 U11103 ( .A1(n5990), .A2(keyinput91), .B1(n10156), .B2(keyinput112), 
        .ZN(n10049) );
  OAI221_X1 U11104 ( .B1(n5990), .B2(keyinput91), .C1(n10156), .C2(keyinput112), .A(n10049), .ZN(n10050) );
  INV_X1 U11105 ( .A(n10050), .ZN(n10060) );
  XNOR2_X1 U11106 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(keyinput122), .ZN(n10053)
         );
  XNOR2_X1 U11107 ( .A(P1_IR_REG_30__SCAN_IN), .B(keyinput72), .ZN(n10052) );
  XNOR2_X1 U11108 ( .A(P2_IR_REG_20__SCAN_IN), .B(keyinput81), .ZN(n10051) );
  AND3_X1 U11109 ( .A1(n10053), .A2(n10052), .A3(n10051), .ZN(n10059) );
  AOI22_X1 U11110 ( .A1(n10161), .A2(keyinput95), .B1(n5573), .B2(keyinput123), 
        .ZN(n10054) );
  OAI221_X1 U11111 ( .B1(n10161), .B2(keyinput95), .C1(n5573), .C2(keyinput123), .A(n10054), .ZN(n10055) );
  INV_X1 U11112 ( .A(n10055), .ZN(n10058) );
  INV_X1 U11113 ( .A(keyinput92), .ZN(n10056) );
  XNOR2_X1 U11114 ( .A(n10144), .B(n10056), .ZN(n10057) );
  AND4_X1 U11115 ( .A1(n10060), .A2(n10059), .A3(n10058), .A4(n10057), .ZN(
        n10101) );
  AOI22_X1 U11116 ( .A1(n10062), .A2(keyinput107), .B1(n6302), .B2(keyinput99), 
        .ZN(n10061) );
  OAI221_X1 U11117 ( .B1(n10062), .B2(keyinput107), .C1(n6302), .C2(keyinput99), .A(n10061), .ZN(n10073) );
  AOI22_X1 U11118 ( .A1(n10064), .A2(keyinput106), .B1(n10146), .B2(keyinput69), .ZN(n10063) );
  OAI221_X1 U11119 ( .B1(n10064), .B2(keyinput106), .C1(n10146), .C2(
        keyinput69), .A(n10063), .ZN(n10072) );
  AOI22_X1 U11120 ( .A1(n10067), .A2(keyinput87), .B1(keyinput83), .B2(n10066), 
        .ZN(n10065) );
  OAI221_X1 U11121 ( .B1(n10067), .B2(keyinput87), .C1(n10066), .C2(keyinput83), .A(n10065), .ZN(n10071) );
  XOR2_X1 U11122 ( .A(n5815), .B(keyinput68), .Z(n10069) );
  XNOR2_X1 U11123 ( .A(P2_IR_REG_29__SCAN_IN), .B(keyinput119), .ZN(n10068) );
  NAND2_X1 U11124 ( .A1(n10069), .A2(n10068), .ZN(n10070) );
  NOR4_X1 U11125 ( .A1(n10073), .A2(n10072), .A3(n10071), .A4(n10070), .ZN(
        n10100) );
  AOI22_X1 U11126 ( .A1(n10164), .A2(keyinput94), .B1(n10075), .B2(keyinput116), .ZN(n10074) );
  OAI221_X1 U11127 ( .B1(n10164), .B2(keyinput94), .C1(n10075), .C2(
        keyinput116), .A(n10074), .ZN(n10086) );
  AOI22_X1 U11128 ( .A1(n10078), .A2(keyinput127), .B1(keyinput120), .B2(
        n10077), .ZN(n10076) );
  OAI221_X1 U11129 ( .B1(n10078), .B2(keyinput127), .C1(n10077), .C2(
        keyinput120), .A(n10076), .ZN(n10085) );
  AOI22_X1 U11130 ( .A1(n6417), .A2(keyinput98), .B1(n10080), .B2(keyinput64), 
        .ZN(n10079) );
  OAI221_X1 U11131 ( .B1(n6417), .B2(keyinput98), .C1(n10080), .C2(keyinput64), 
        .A(n10079), .ZN(n10084) );
  AOI22_X1 U11132 ( .A1(n10082), .A2(keyinput89), .B1(keyinput96), .B2(n8520), 
        .ZN(n10081) );
  OAI221_X1 U11133 ( .B1(n10082), .B2(keyinput89), .C1(n8520), .C2(keyinput96), 
        .A(n10081), .ZN(n10083) );
  NOR4_X1 U11134 ( .A1(n10086), .A2(n10085), .A3(n10084), .A4(n10083), .ZN(
        n10099) );
  INV_X1 U11135 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n10150) );
  AOI22_X1 U11136 ( .A1(n8354), .A2(keyinput118), .B1(n10150), .B2(keyinput82), 
        .ZN(n10087) );
  OAI221_X1 U11137 ( .B1(n8354), .B2(keyinput118), .C1(n10150), .C2(keyinput82), .A(n10087), .ZN(n10097) );
  AOI22_X1 U11138 ( .A1(n10089), .A2(keyinput108), .B1(keyinput80), .B2(n5712), 
        .ZN(n10088) );
  OAI221_X1 U11139 ( .B1(n10089), .B2(keyinput108), .C1(n5712), .C2(keyinput80), .A(n10088), .ZN(n10096) );
  AOI22_X1 U11140 ( .A1(n10158), .A2(keyinput67), .B1(keyinput73), .B2(n10091), 
        .ZN(n10090) );
  OAI221_X1 U11141 ( .B1(n10158), .B2(keyinput67), .C1(n10091), .C2(keyinput73), .A(n10090), .ZN(n10095) );
  AOI22_X1 U11142 ( .A1(n5960), .A2(keyinput115), .B1(keyinput125), .B2(n10093), .ZN(n10092) );
  OAI221_X1 U11143 ( .B1(n5960), .B2(keyinput115), .C1(n10093), .C2(
        keyinput125), .A(n10092), .ZN(n10094) );
  NOR4_X1 U11144 ( .A1(n10097), .A2(n10096), .A3(n10095), .A4(n10094), .ZN(
        n10098) );
  NAND4_X1 U11145 ( .A1(n10101), .A2(n10100), .A3(n10099), .A4(n10098), .ZN(
        n10172) );
  AOI22_X1 U11146 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(keyinput79), .B1(
        P1_D_REG_16__SCAN_IN), .B2(keyinput102), .ZN(n10102) );
  OAI221_X1 U11147 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(keyinput79), .C1(
        P1_D_REG_16__SCAN_IN), .C2(keyinput102), .A(n10102), .ZN(n10109) );
  AOI22_X1 U11148 ( .A1(P2_REG0_REG_9__SCAN_IN), .A2(keyinput104), .B1(
        P1_REG3_REG_17__SCAN_IN), .B2(keyinput105), .ZN(n10103) );
  OAI221_X1 U11149 ( .B1(P2_REG0_REG_9__SCAN_IN), .B2(keyinput104), .C1(
        P1_REG3_REG_17__SCAN_IN), .C2(keyinput105), .A(n10103), .ZN(n10108) );
  AOI22_X1 U11150 ( .A1(P2_REG1_REG_20__SCAN_IN), .A2(keyinput71), .B1(
        P2_IR_REG_0__SCAN_IN), .B2(keyinput93), .ZN(n10104) );
  OAI221_X1 U11151 ( .B1(P2_REG1_REG_20__SCAN_IN), .B2(keyinput71), .C1(
        P2_IR_REG_0__SCAN_IN), .C2(keyinput93), .A(n10104), .ZN(n10107) );
  AOI22_X1 U11152 ( .A1(P1_REG0_REG_16__SCAN_IN), .A2(keyinput101), .B1(
        P1_REG0_REG_28__SCAN_IN), .B2(keyinput111), .ZN(n10105) );
  OAI221_X1 U11153 ( .B1(P1_REG0_REG_16__SCAN_IN), .B2(keyinput101), .C1(
        P1_REG0_REG_28__SCAN_IN), .C2(keyinput111), .A(n10105), .ZN(n10106) );
  NOR4_X1 U11154 ( .A1(n10109), .A2(n10108), .A3(n10107), .A4(n10106), .ZN(
        n10139) );
  AOI22_X1 U11155 ( .A1(P2_REG0_REG_10__SCAN_IN), .A2(keyinput124), .B1(
        P2_REG1_REG_11__SCAN_IN), .B2(keyinput100), .ZN(n10110) );
  OAI221_X1 U11156 ( .B1(P2_REG0_REG_10__SCAN_IN), .B2(keyinput124), .C1(
        P2_REG1_REG_11__SCAN_IN), .C2(keyinput100), .A(n10110), .ZN(n10117) );
  AOI22_X1 U11157 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(keyinput77), .B1(
        P1_REG0_REG_5__SCAN_IN), .B2(keyinput88), .ZN(n10111) );
  OAI221_X1 U11158 ( .B1(P2_IR_REG_31__SCAN_IN), .B2(keyinput77), .C1(
        P1_REG0_REG_5__SCAN_IN), .C2(keyinput88), .A(n10111), .ZN(n10116) );
  AOI22_X1 U11159 ( .A1(P2_REG2_REG_10__SCAN_IN), .A2(keyinput103), .B1(
        P2_REG3_REG_25__SCAN_IN), .B2(keyinput66), .ZN(n10112) );
  OAI221_X1 U11160 ( .B1(P2_REG2_REG_10__SCAN_IN), .B2(keyinput103), .C1(
        P2_REG3_REG_25__SCAN_IN), .C2(keyinput66), .A(n10112), .ZN(n10115) );
  AOI22_X1 U11161 ( .A1(P2_REG0_REG_6__SCAN_IN), .A2(keyinput70), .B1(
        P1_REG3_REG_11__SCAN_IN), .B2(keyinput86), .ZN(n10113) );
  OAI221_X1 U11162 ( .B1(P2_REG0_REG_6__SCAN_IN), .B2(keyinput70), .C1(
        P1_REG3_REG_11__SCAN_IN), .C2(keyinput86), .A(n10113), .ZN(n10114) );
  NOR4_X1 U11163 ( .A1(n10117), .A2(n10116), .A3(n10115), .A4(n10114), .ZN(
        n10138) );
  AOI22_X1 U11164 ( .A1(P1_REG1_REG_26__SCAN_IN), .A2(keyinput110), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(keyinput126), .ZN(n10118) );
  OAI221_X1 U11165 ( .B1(P1_REG1_REG_26__SCAN_IN), .B2(keyinput110), .C1(
        P2_DATAO_REG_9__SCAN_IN), .C2(keyinput126), .A(n10118), .ZN(n10127) );
  AOI22_X1 U11166 ( .A1(P2_REG1_REG_29__SCAN_IN), .A2(keyinput74), .B1(
        P2_IR_REG_16__SCAN_IN), .B2(keyinput121), .ZN(n10119) );
  OAI221_X1 U11167 ( .B1(P2_REG1_REG_29__SCAN_IN), .B2(keyinput74), .C1(
        P2_IR_REG_16__SCAN_IN), .C2(keyinput121), .A(n10119), .ZN(n10126) );
  AOI22_X1 U11168 ( .A1(n10121), .A2(keyinput90), .B1(n10149), .B2(keyinput109), .ZN(n10120) );
  OAI221_X1 U11169 ( .B1(n10121), .B2(keyinput90), .C1(n10149), .C2(
        keyinput109), .A(n10120), .ZN(n10125) );
  INV_X1 U11170 ( .A(SI_14_), .ZN(n10160) );
  AOI22_X1 U11171 ( .A1(n10123), .A2(keyinput113), .B1(n10160), .B2(
        keyinput114), .ZN(n10122) );
  OAI221_X1 U11172 ( .B1(n10123), .B2(keyinput113), .C1(n10160), .C2(
        keyinput114), .A(n10122), .ZN(n10124) );
  NOR4_X1 U11173 ( .A1(n10127), .A2(n10126), .A3(n10125), .A4(n10124), .ZN(
        n10137) );
  AOI22_X1 U11174 ( .A1(P1_ADDR_REG_14__SCAN_IN), .A2(keyinput75), .B1(
        P1_REG2_REG_18__SCAN_IN), .B2(keyinput76), .ZN(n10128) );
  OAI221_X1 U11175 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(keyinput75), .C1(
        P1_REG2_REG_18__SCAN_IN), .C2(keyinput76), .A(n10128), .ZN(n10135) );
  AOI22_X1 U11176 ( .A1(P2_REG1_REG_31__SCAN_IN), .A2(keyinput97), .B1(
        P1_DATAO_REG_10__SCAN_IN), .B2(keyinput65), .ZN(n10129) );
  OAI221_X1 U11177 ( .B1(P2_REG1_REG_31__SCAN_IN), .B2(keyinput97), .C1(
        P1_DATAO_REG_10__SCAN_IN), .C2(keyinput65), .A(n10129), .ZN(n10134) );
  AOI22_X1 U11178 ( .A1(P1_REG1_REG_28__SCAN_IN), .A2(keyinput84), .B1(
        P1_IR_REG_16__SCAN_IN), .B2(keyinput117), .ZN(n10130) );
  OAI221_X1 U11179 ( .B1(P1_REG1_REG_28__SCAN_IN), .B2(keyinput84), .C1(
        P1_IR_REG_16__SCAN_IN), .C2(keyinput117), .A(n10130), .ZN(n10133) );
  AOI22_X1 U11180 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(keyinput78), .B1(
        P1_D_REG_7__SCAN_IN), .B2(keyinput85), .ZN(n10131) );
  OAI221_X1 U11181 ( .B1(P2_REG3_REG_11__SCAN_IN), .B2(keyinput78), .C1(
        P1_D_REG_7__SCAN_IN), .C2(keyinput85), .A(n10131), .ZN(n10132) );
  NOR4_X1 U11182 ( .A1(n10135), .A2(n10134), .A3(n10133), .A4(n10132), .ZN(
        n10136) );
  NAND4_X1 U11183 ( .A1(n10139), .A2(n10138), .A3(n10137), .A4(n10136), .ZN(
        n10171) );
  AOI22_X1 U11184 ( .A1(n10142), .A2(keyinput2), .B1(n10141), .B2(keyinput21), 
        .ZN(n10140) );
  OAI221_X1 U11185 ( .B1(n10142), .B2(keyinput2), .C1(n10141), .C2(keyinput21), 
        .A(n10140), .ZN(n10154) );
  AOI22_X1 U11186 ( .A1(n6302), .A2(keyinput35), .B1(keyinput28), .B2(n10144), 
        .ZN(n10143) );
  OAI221_X1 U11187 ( .B1(n6302), .B2(keyinput35), .C1(n10144), .C2(keyinput28), 
        .A(n10143), .ZN(n10153) );
  AOI22_X1 U11188 ( .A1(n10147), .A2(keyinput40), .B1(n10146), .B2(keyinput5), 
        .ZN(n10145) );
  OAI221_X1 U11189 ( .B1(n10147), .B2(keyinput40), .C1(n10146), .C2(keyinput5), 
        .A(n10145), .ZN(n10152) );
  AOI22_X1 U11190 ( .A1(n10150), .A2(keyinput18), .B1(n10149), .B2(keyinput45), 
        .ZN(n10148) );
  OAI221_X1 U11191 ( .B1(n10150), .B2(keyinput18), .C1(n10149), .C2(keyinput45), .A(n10148), .ZN(n10151) );
  NOR4_X1 U11192 ( .A1(n10154), .A2(n10153), .A3(n10152), .A4(n10151), .ZN(
        n10170) );
  AOI22_X1 U11193 ( .A1(n10156), .A2(keyinput48), .B1(keyinput59), .B2(n5573), 
        .ZN(n10155) );
  OAI221_X1 U11194 ( .B1(n10156), .B2(keyinput48), .C1(n5573), .C2(keyinput59), 
        .A(n10155), .ZN(n10168) );
  AOI22_X1 U11195 ( .A1(P1_D_REG_16__SCAN_IN), .A2(keyinput38), .B1(n10158), 
        .B2(keyinput3), .ZN(n10157) );
  OAI221_X1 U11196 ( .B1(P1_D_REG_16__SCAN_IN), .B2(keyinput38), .C1(n10158), 
        .C2(keyinput3), .A(n10157), .ZN(n10167) );
  AOI22_X1 U11197 ( .A1(n10161), .A2(keyinput31), .B1(n10160), .B2(keyinput50), 
        .ZN(n10159) );
  OAI221_X1 U11198 ( .B1(n10161), .B2(keyinput31), .C1(n10160), .C2(keyinput50), .A(n10159), .ZN(n10166) );
  AOI22_X1 U11199 ( .A1(n10164), .A2(keyinput30), .B1(n10163), .B2(keyinput46), 
        .ZN(n10162) );
  OAI221_X1 U11200 ( .B1(n10164), .B2(keyinput30), .C1(n10163), .C2(keyinput46), .A(n10162), .ZN(n10165) );
  NOR4_X1 U11201 ( .A1(n10168), .A2(n10167), .A3(n10166), .A4(n10165), .ZN(
        n10169) );
  OAI211_X1 U11202 ( .C1(n10172), .C2(n10171), .A(n10170), .B(n10169), .ZN(
        n10173) );
  NOR4_X1 U11203 ( .A1(n10176), .A2(n10175), .A3(n10174), .A4(n10173), .ZN(
        n10177) );
  XNOR2_X1 U11204 ( .A(n10178), .B(n10177), .ZN(P2_U3302) );
  XOR2_X1 U11205 ( .A(n10179), .B(P2_ADDR_REG_6__SCAN_IN), .Z(ADD_1071_U50) );
  NOR2_X1 U11206 ( .A1(n10181), .A2(n10180), .ZN(n10182) );
  XOR2_X1 U11207 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n10182), .Z(ADD_1071_U51) );
  XOR2_X1 U11208 ( .A(n10183), .B(P2_ADDR_REG_7__SCAN_IN), .Z(ADD_1071_U49) );
  OAI21_X1 U11209 ( .B1(n10186), .B2(n10185), .A(n10184), .ZN(n10188) );
  XOR2_X1 U11210 ( .A(n10188), .B(n10187), .Z(ADD_1071_U55) );
  XOR2_X1 U11211 ( .A(n10189), .B(P2_ADDR_REG_8__SCAN_IN), .Z(ADD_1071_U48) );
  AOI21_X1 U11212 ( .B1(n10192), .B2(n10191), .A(n10190), .ZN(ADD_1071_U47) );
  XOR2_X1 U11213 ( .A(n10194), .B(n10193), .Z(ADD_1071_U54) );
  XOR2_X1 U11214 ( .A(n10196), .B(n10195), .Z(ADD_1071_U53) );
  XNOR2_X1 U11215 ( .A(n10198), .B(n10197), .ZN(ADD_1071_U52) );
  CLKBUF_X1 U4796 ( .A(n5806), .Z(n6139) );
  CLKBUF_X1 U4800 ( .A(n6690), .Z(n7375) );
  NAND2_X1 U4804 ( .A1(n5459), .A2(n8002), .ZN(n5050) );
  CLKBUF_X1 U4946 ( .A(n5799), .Z(n8082) );
  CLKBUF_X2 U5756 ( .A(n7153), .Z(n4298) );
  CLKBUF_X1 U6119 ( .A(n5826), .Z(n8088) );
  INV_X2 U6222 ( .A(n9219), .ZN(n9620) );
endmodule

