

module b14_C_SARLock_k_64_3 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, U3352, U3351, U3350, U3349, U3348, U3347, 
        U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, U3338, U3337, 
        U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, U3328, U3327, 
        U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, U3320, U3319, 
        U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, U3310, U3309, 
        U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, U3300, U3299, 
        U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, U3467, U3469, 
        U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, U3487, U3489, 
        U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, U3506, U3507, 
        U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, U3516, U3517, 
        U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, U3526, U3527, 
        U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, U3536, U3537, 
        U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, U3546, U3547, 
        U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, U3284, U3283, 
        U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, U3274, U3273, 
        U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, U3264, U3263, 
        U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, U3255, U3254, 
        U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, U3245, U3244, 
        U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, U3554, U3555, 
        U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, U3564, U3565, 
        U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, U3574, U3575, 
        U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, U3237, U3236, 
        U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, U3227, U3226, 
        U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, U3217, U3216, 
        U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, U4043 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038,
         n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048,
         n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058,
         n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068,
         n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078,
         n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088,
         n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098,
         n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108,
         n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118,
         n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128,
         n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138,
         n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148,
         n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158,
         n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168,
         n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178,
         n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188,
         n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198,
         n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208,
         n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218,
         n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228,
         n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238,
         n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248,
         n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258,
         n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268,
         n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278,
         n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288,
         n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298,
         n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308,
         n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318,
         n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328,
         n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338,
         n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348,
         n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358,
         n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368,
         n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378,
         n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388,
         n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398,
         n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408,
         n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418,
         n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428,
         n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438,
         n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448,
         n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458,
         n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468,
         n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478,
         n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488,
         n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498,
         n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508,
         n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518,
         n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528,
         n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538,
         n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548,
         n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558,
         n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568,
         n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578,
         n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588,
         n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598,
         n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608,
         n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618,
         n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628,
         n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638,
         n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648,
         n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658,
         n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668,
         n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678,
         n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688,
         n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698,
         n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708,
         n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718,
         n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728,
         n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738,
         n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748,
         n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758,
         n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768,
         n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778,
         n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788,
         n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798,
         n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808,
         n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818,
         n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828,
         n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838,
         n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848,
         n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858,
         n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868,
         n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878,
         n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888,
         n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898,
         n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908,
         n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918,
         n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928,
         n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938,
         n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948,
         n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958,
         n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968,
         n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978,
         n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988,
         n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998,
         n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008,
         n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018,
         n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028,
         n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038,
         n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048,
         n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058,
         n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068,
         n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078,
         n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088,
         n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098,
         n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108,
         n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118,
         n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128,
         n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138,
         n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148,
         n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158,
         n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168,
         n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178,
         n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188,
         n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198,
         n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208,
         n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218,
         n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
         n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
         n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248,
         n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258,
         n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268,
         n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278,
         n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288,
         n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298,
         n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308,
         n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318,
         n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328,
         n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338,
         n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348,
         n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358,
         n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368,
         n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378,
         n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388,
         n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398,
         n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408,
         n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418,
         n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428,
         n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438,
         n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448,
         n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458,
         n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468,
         n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478,
         n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488,
         n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498,
         n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508,
         n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518,
         n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528,
         n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538,
         n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548,
         n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558,
         n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568,
         n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578,
         n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588,
         n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598,
         n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608,
         n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618,
         n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628,
         n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638,
         n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648,
         n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658,
         n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668,
         n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678,
         n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688,
         n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698,
         n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708,
         n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718,
         n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728,
         n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738,
         n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748,
         n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758,
         n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768,
         n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778,
         n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788,
         n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798,
         n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808,
         n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818,
         n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828,
         n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838,
         n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848,
         n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858,
         n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868,
         n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878,
         n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888,
         n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898,
         n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908,
         n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918,
         n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928,
         n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938,
         n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948,
         n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958,
         n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968,
         n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978,
         n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988,
         n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998,
         n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008,
         n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018,
         n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028,
         n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038,
         n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048,
         n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058,
         n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068,
         n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078,
         n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088,
         n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098,
         n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108,
         n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118,
         n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128,
         n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138,
         n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148,
         n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158,
         n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168,
         n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178,
         n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188,
         n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198,
         n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208,
         n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218,
         n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228,
         n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238,
         n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248,
         n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258,
         n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268,
         n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278,
         n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288,
         n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298,
         n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308,
         n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318,
         n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328,
         n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338,
         n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348,
         n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
         n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368,
         n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378,
         n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
         n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
         n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
         n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
         n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
         n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
         n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
         n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
         n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
         n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
         n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
         n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
         n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
         n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
         n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
         n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
         n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
         n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
         n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
         n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
         n4579;

  CLKBUF_X2 U2272 ( .A(n2369), .Z(n2029) );
  CLKBUF_X2 U2273 ( .A(n2332), .Z(n2398) );
  INV_X1 U2274 ( .A(n2339), .ZN(n3190) );
  OR2_X1 U2275 ( .A1(n2339), .A2(n4540), .ZN(n2330) );
  INV_X1 U2276 ( .A(n2687), .ZN(n3193) );
  INV_X1 U2277 ( .A(n2378), .ZN(n2242) );
  XNOR2_X1 U2278 ( .A(n2299), .B(IR_REG_22__SCAN_IN), .ZN(n4258) );
  XNOR2_X2 U2279 ( .A(n2871), .B(n4266), .ZN(n2895) );
  AOI21_X2 U2280 ( .B1(n4502), .B2(REG1_REG_5__SCAN_IN), .A(n4282), .ZN(n2873)
         );
  NOR2_X2 U2281 ( .A1(n4284), .A2(n4283), .ZN(n4282) );
  OR2_X2 U2282 ( .A1(n4459), .A2(n4260), .ZN(n2841) );
  AND2_X4 U2283 ( .A1(n4255), .A2(n2852), .ZN(n2345) );
  NAND4_X1 U2284 ( .A1(n2350), .A2(n2349), .A3(n2348), .A4(n2347), .ZN(n3623)
         );
  AND2_X1 U2285 ( .A1(n2814), .A2(n2813), .ZN(n3827) );
  AND2_X1 U2286 ( .A1(n3304), .A2(n3443), .ZN(n2546) );
  AOI21_X1 U2287 ( .B1(n3844), .B2(n3540), .A(n3541), .ZN(n3825) );
  AND2_X1 U2288 ( .A1(n2207), .A2(n2206), .ZN(n4360) );
  NAND2_X1 U2289 ( .A1(n2804), .A2(n3465), .ZN(n3960) );
  OR2_X1 U2290 ( .A1(n3127), .A2(n3463), .ZN(n3156) );
  NAND2_X1 U2291 ( .A1(n4326), .A2(n2056), .ZN(n3072) );
  NAND2_X1 U2292 ( .A1(n2801), .A2(n3495), .ZN(n3142) );
  OR2_X1 U2293 ( .A1(n3045), .A2(n3044), .ZN(n2801) );
  NAND2_X1 U2294 ( .A1(n2114), .A2(n2113), .ZN(n2112) );
  NAND2_X1 U2295 ( .A1(n2049), .A2(n2034), .ZN(n2103) );
  OR2_X1 U2296 ( .A1(n2929), .A2(n2344), .ZN(n2114) );
  OAI211_X1 U2297 ( .C1(n2936), .C2(n2165), .A(n2757), .B(n2163), .ZN(n2979)
         );
  AOI21_X1 U2298 ( .B1(n2074), .B2(n2077), .A(n2072), .ZN(n2071) );
  AOI21_X1 U2299 ( .B1(n3457), .B2(n2076), .A(n2075), .ZN(n2074) );
  INV_X2 U2300 ( .A(n3388), .ZN(n3449) );
  AND2_X1 U2301 ( .A1(n2338), .A2(n2337), .ZN(n2342) );
  OR2_X1 U2302 ( .A1(n4447), .A2(n3534), .ZN(n4436) );
  INV_X1 U2303 ( .A(n2937), .ZN(n3622) );
  AND4_X1 U2304 ( .A1(n2362), .A2(n2361), .A3(n2360), .A4(n2359), .ZN(n2937)
         );
  INV_X1 U2305 ( .A(n2841), .ZN(n4540) );
  AND2_X1 U2306 ( .A1(n2908), .A2(REG1_REG_4__SCAN_IN), .ZN(n2918) );
  XNOR2_X1 U2307 ( .A(n2182), .B(n2921), .ZN(n2908) );
  NAND4_X1 U2308 ( .A1(n2321), .A2(n2320), .A3(n2319), .A4(n2318), .ZN(n2748)
         );
  NAND2_X2 U2309 ( .A1(n2951), .A2(n2714), .ZN(n2687) );
  NAND2_X1 U2310 ( .A1(n2301), .A2(n2300), .ZN(n4459) );
  OR2_X1 U2311 ( .A1(n2894), .A2(n2872), .ZN(n2182) );
  NAND2_X1 U2312 ( .A1(n2730), .A2(n4259), .ZN(n2951) );
  OR3_X2 U2313 ( .A1(n2690), .A2(n2704), .A3(n2096), .ZN(n2849) );
  INV_X1 U2314 ( .A(n2730), .ZN(n4260) );
  CLKBUF_X3 U2315 ( .A(n2346), .Z(n3518) );
  BUF_X2 U2316 ( .A(n2331), .Z(n3514) );
  XNOR2_X1 U2317 ( .A(n2295), .B(n2294), .ZN(n2730) );
  NAND2_X1 U2318 ( .A1(n2313), .A2(IR_REG_31__SCAN_IN), .ZN(n2295) );
  AND2_X1 U2319 ( .A1(n2298), .A2(n2040), .ZN(n4259) );
  XNOR2_X1 U2320 ( .A(n2277), .B(IR_REG_30__SCAN_IN), .ZN(n4255) );
  NAND2_X1 U2321 ( .A1(n2278), .A2(IR_REG_31__SCAN_IN), .ZN(n2277) );
  OAI21_X1 U2322 ( .B1(n2296), .B2(n2258), .A(IR_REG_31__SCAN_IN), .ZN(n2708)
         );
  OR2_X1 U2323 ( .A1(n2285), .A2(n2718), .ZN(n2291) );
  NAND2_X1 U2324 ( .A1(n3626), .A2(n3627), .ZN(n3641) );
  NOR2_X1 U2325 ( .A1(n2243), .A2(n2272), .ZN(n2241) );
  OAI211_X2 U2326 ( .C1(n2179), .C2(n4505), .A(n2180), .B(n2170), .ZN(n4268)
         );
  NAND2_X1 U2327 ( .A1(n2718), .A2(IR_REG_1__SCAN_IN), .ZN(n2180) );
  NAND2_X1 U2328 ( .A1(n4505), .A2(IR_REG_1__SCAN_IN), .ZN(n2170) );
  NAND2_X1 U2329 ( .A1(n2260), .A2(n2259), .ZN(n2258) );
  INV_X1 U2330 ( .A(IR_REG_0__SCAN_IN), .ZN(n2220) );
  NOR2_X1 U2331 ( .A1(IR_REG_8__SCAN_IN), .A2(IR_REG_7__SCAN_IN), .ZN(n2271)
         );
  NOR2_X1 U2332 ( .A1(IR_REG_16__SCAN_IN), .A2(IR_REG_15__SCAN_IN), .ZN(n2119)
         );
  NOR2_X1 U2333 ( .A1(IR_REG_14__SCAN_IN), .A2(IR_REG_13__SCAN_IN), .ZN(n2118)
         );
  NOR2_X1 U2334 ( .A1(IR_REG_12__SCAN_IN), .A2(IR_REG_11__SCAN_IN), .ZN(n2117)
         );
  NOR2_X1 U2335 ( .A1(IR_REG_10__SCAN_IN), .A2(IR_REG_9__SCAN_IN), .ZN(n2116)
         );
  NOR3_X1 U2336 ( .A1(IR_REG_20__SCAN_IN), .A2(IR_REG_19__SCAN_IN), .A3(
        IR_REG_18__SCAN_IN), .ZN(n2274) );
  INV_X1 U2337 ( .A(IR_REG_3__SCAN_IN), .ZN(n2363) );
  NOR2_X2 U2338 ( .A1(n4373), .A2(n3664), .ZN(n4382) );
  INV_X4 U2339 ( .A(n2330), .ZN(n3195) );
  AOI21_X1 U2340 ( .B1(n2224), .B2(n2226), .A(n2223), .ZN(n2222) );
  INV_X1 U2341 ( .A(n3219), .ZN(n2511) );
  AOI21_X1 U2342 ( .B1(n3265), .B2(n3264), .A(n2253), .ZN(n2252) );
  INV_X1 U2343 ( .A(n2414), .ZN(n2253) );
  NAND2_X1 U2344 ( .A1(n2305), .A2(n2849), .ZN(n2369) );
  NOR2_X1 U2345 ( .A1(n3766), .A2(n3588), .ZN(n3747) );
  NAND2_X1 U2346 ( .A1(n3226), .A2(n2634), .ZN(n3229) );
  NAND2_X1 U2347 ( .A1(n2115), .A2(n2649), .ZN(n3333) );
  NAND2_X1 U2348 ( .A1(n3229), .A2(n2647), .ZN(n2115) );
  AOI21_X1 U2349 ( .B1(n3254), .B2(n2107), .A(n2058), .ZN(n2106) );
  NAND2_X1 U2350 ( .A1(n3254), .A2(n2109), .ZN(n2108) );
  INV_X1 U2351 ( .A(n3409), .ZN(n2107) );
  MUX2_X1 U2352 ( .A(n4267), .B(DATAI_2_), .S(n2352), .Z(n2964) );
  NAND2_X1 U2353 ( .A1(n4324), .A2(n4325), .ZN(n4323) );
  OR2_X1 U2354 ( .A1(n3206), .A2(n2840), .ZN(n2130) );
  INV_X1 U2355 ( .A(n2790), .ZN(n2125) );
  INV_X1 U2356 ( .A(n2127), .ZN(n2126) );
  NAND2_X1 U2357 ( .A1(n2788), .A2(n2263), .ZN(n3728) );
  AND2_X1 U2358 ( .A1(n3904), .A2(n3891), .ZN(n2776) );
  OAI22_X1 U2359 ( .A1(n3132), .A2(n2768), .B1(n4404), .B2(n3128), .ZN(n3162)
         );
  AOI21_X1 U2360 ( .B1(n2141), .B2(n2144), .A(n2047), .ZN(n2140) );
  NOR2_X1 U2361 ( .A1(n2031), .A2(n2765), .ZN(n2141) );
  NAND2_X1 U2362 ( .A1(n2144), .A2(n2143), .ZN(n2142) );
  INV_X1 U2363 ( .A(n2765), .ZN(n2143) );
  AND2_X1 U2364 ( .A1(n2276), .A2(n2303), .ZN(n2256) );
  AND2_X1 U2365 ( .A1(n2273), .A2(n2275), .ZN(n2196) );
  NAND2_X1 U2366 ( .A1(n2748), .A2(n4453), .ZN(n3468) );
  OR2_X1 U2367 ( .A1(n2499), .A2(n2227), .ZN(n2226) );
  INV_X1 U2368 ( .A(n3397), .ZN(n2227) );
  NOR2_X1 U2369 ( .A1(n2235), .A2(n2231), .ZN(n2230) );
  INV_X1 U2370 ( .A(n2634), .ZN(n2231) );
  NOR2_X1 U2371 ( .A1(n3335), .A2(n2649), .ZN(n2235) );
  INV_X1 U2372 ( .A(n2645), .ZN(n2234) );
  OAI22_X1 U2373 ( .A1(n2937), .A2(n2029), .B1(n2339), .B2(n3000), .ZN(n2370)
         );
  INV_X1 U2374 ( .A(n3245), .ZN(n2113) );
  NAND2_X1 U2375 ( .A1(n2250), .A2(n2251), .ZN(n2248) );
  NAND2_X1 U2376 ( .A1(n3061), .A2(n2252), .ZN(n2249) );
  INV_X1 U2377 ( .A(n3265), .ZN(n2250) );
  NAND2_X1 U2378 ( .A1(n4505), .A2(n2183), .ZN(n2168) );
  NAND2_X1 U2379 ( .A1(n2179), .A2(IR_REG_0__SCAN_IN), .ZN(n2169) );
  OAI22_X1 U2380 ( .A1(n4348), .A2(n4344), .B1(REG2_REG_13__SCAN_IN), .B2(
        n4491), .ZN(n3074) );
  OR2_X1 U2381 ( .A1(n3513), .A2(n3572), .ZN(n3548) );
  AOI21_X1 U2382 ( .B1(n3827), .B2(n3582), .A(n2817), .ZN(n3766) );
  NOR2_X1 U2383 ( .A1(n3578), .A2(n2094), .ZN(n2093) );
  INV_X1 U2384 ( .A(n3579), .ZN(n2094) );
  AND2_X1 U2385 ( .A1(n2153), .A2(n2772), .ZN(n2147) );
  INV_X1 U2386 ( .A(n3475), .ZN(n2085) );
  AND2_X1 U2387 ( .A1(n2038), .A2(n3835), .ZN(n2195) );
  NOR2_X1 U2388 ( .A1(n3377), .A2(n3286), .ZN(n2193) );
  NAND2_X1 U2389 ( .A1(n3468), .A2(n2793), .ZN(n4447) );
  NOR2_X1 U2390 ( .A1(IR_REG_26__SCAN_IN), .A2(IR_REG_27__SCAN_IN), .ZN(n2276)
         );
  INV_X1 U2391 ( .A(n2258), .ZN(n2257) );
  INV_X1 U2392 ( .A(IR_REG_25__SCAN_IN), .ZN(n2275) );
  INV_X1 U2393 ( .A(IR_REG_23__SCAN_IN), .ZN(n2707) );
  INV_X1 U2394 ( .A(n2243), .ZN(n2240) );
  OAI22_X1 U2395 ( .A1(n2771), .A2(n2657), .B1(n2029), .B2(n2838), .ZN(n3216)
         );
  AND2_X1 U2396 ( .A1(n2607), .A2(n2606), .ZN(n3274) );
  INV_X1 U2397 ( .A(n2112), .ZN(n3346) );
  NAND2_X1 U2398 ( .A1(n2099), .A2(n2097), .ZN(n3115) );
  AND2_X1 U2399 ( .A1(n2103), .A2(n2098), .ZN(n2097) );
  INV_X1 U2400 ( .A(n3118), .ZN(n2098) );
  INV_X1 U2401 ( .A(n3358), .ZN(n2237) );
  INV_X1 U2402 ( .A(n3385), .ZN(n2621) );
  NAND2_X1 U2403 ( .A1(n3195), .A2(n2751), .ZN(n2337) );
  NAND2_X1 U2404 ( .A1(n4439), .A2(n3190), .ZN(n2322) );
  OAI22_X2 U2405 ( .A1(n3323), .A2(n2560), .B1(n3324), .B2(n2559), .ZN(n3411)
         );
  OR2_X1 U2406 ( .A1(n2650), .A2(n3298), .ZN(n2662) );
  INV_X1 U2407 ( .A(n2692), .ZN(n2096) );
  NAND2_X1 U2408 ( .A1(n2177), .A2(n4562), .ZN(n2176) );
  INV_X1 U2409 ( .A(n2180), .ZN(n2177) );
  NAND2_X1 U2410 ( .A1(n2168), .A2(n2169), .ZN(n2178) );
  XNOR2_X1 U2411 ( .A(n2881), .B(n2210), .ZN(n2897) );
  NAND2_X1 U2412 ( .A1(n2897), .A2(REG2_REG_3__SCAN_IN), .ZN(n2896) );
  NAND2_X1 U2413 ( .A1(n4287), .A2(n2046), .ZN(n2883) );
  NAND2_X1 U2414 ( .A1(n4264), .A2(REG2_REG_7__SCAN_IN), .ZN(n2204) );
  NAND2_X1 U2415 ( .A1(n4323), .A2(n2064), .ZN(n3092) );
  NAND2_X1 U2416 ( .A1(n3074), .A2(n3095), .ZN(n2208) );
  NAND2_X1 U2417 ( .A1(n4363), .A2(n2181), .ZN(n3663) );
  NAND2_X1 U2418 ( .A1(n3671), .A2(REG1_REG_15__SCAN_IN), .ZN(n2181) );
  AOI21_X1 U2419 ( .B1(n3671), .B2(REG2_REG_15__SCAN_IN), .A(n4358), .ZN(n3673) );
  OAI21_X1 U2420 ( .B1(n2293), .B2(IR_REG_18__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2314) );
  INV_X1 U2421 ( .A(IR_REG_19__SCAN_IN), .ZN(n4099) );
  NAND2_X1 U2422 ( .A1(n2314), .A2(n4099), .ZN(n2313) );
  AND2_X1 U2423 ( .A1(n4378), .A2(n2215), .ZN(n2213) );
  NOR2_X1 U2424 ( .A1(n2662), .A2(n3436), .ZN(n2679) );
  NOR2_X1 U2425 ( .A1(n3719), .A2(n2839), .ZN(n2790) );
  INV_X1 U2426 ( .A(n3548), .ZN(n3713) );
  NOR2_X1 U2427 ( .A1(n3797), .A2(n2037), .ZN(n3730) );
  OAI22_X1 U2428 ( .A1(n3825), .A2(n2156), .B1(n2158), .B2(n2783), .ZN(n3773)
         );
  AND2_X1 U2429 ( .A1(n2162), .A2(n2159), .ZN(n2158) );
  NAND2_X1 U2430 ( .A1(n2161), .A2(n2030), .ZN(n2156) );
  NAND2_X1 U2431 ( .A1(n2030), .A2(n2160), .ZN(n2159) );
  OR2_X1 U2432 ( .A1(n3923), .A2(n3911), .ZN(n2774) );
  AND2_X1 U2433 ( .A1(n2769), .A2(n2035), .ZN(n2153) );
  NAND2_X1 U2434 ( .A1(n2061), .A2(n2035), .ZN(n2151) );
  NAND2_X1 U2435 ( .A1(n2770), .A2(n2769), .ZN(n2155) );
  AOI21_X1 U2436 ( .B1(n2140), .B2(n2142), .A(n2138), .ZN(n2137) );
  AOI21_X1 U2437 ( .B1(n2031), .B2(n2764), .A(n2048), .ZN(n2144) );
  OAI21_X1 U2438 ( .B1(n3029), .B2(n2081), .A(n2078), .ZN(n3045) );
  AOI21_X1 U2439 ( .B1(n2080), .B2(n2082), .A(n2079), .ZN(n2078) );
  OAI21_X1 U2440 ( .B1(n2980), .B2(n2978), .A(n3485), .ZN(n3009) );
  OAI22_X1 U2441 ( .A1(n2979), .A2(n2758), .B1(n3317), .B2(n3621), .ZN(n3008)
         );
  NOR2_X1 U2442 ( .A1(n4524), .A2(n4259), .ZN(n2833) );
  NAND2_X1 U2443 ( .A1(n2083), .A2(n2939), .ZN(n2941) );
  NAND2_X1 U2444 ( .A1(n2938), .A2(n3469), .ZN(n2083) );
  OR2_X1 U2445 ( .A1(n4459), .A2(n2730), .ZN(n4403) );
  NAND2_X1 U2446 ( .A1(n3983), .A2(n2188), .ZN(n3992) );
  INV_X1 U2447 ( .A(n3269), .ZN(n3103) );
  INV_X1 U2448 ( .A(n4550), .ZN(n4535) );
  NAND2_X1 U2449 ( .A1(n2693), .A2(n2692), .ZN(n2854) );
  NAND2_X1 U2450 ( .A1(n2849), .A2(n4481), .ZN(n2862) );
  NAND2_X1 U2451 ( .A1(n2278), .A2(n2068), .ZN(n2280) );
  AOI21_X1 U2452 ( .B1(n2720), .B2(n2055), .A(n2069), .ZN(n2068) );
  NOR2_X1 U2453 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_29__SCAN_IN), .ZN(n2069)
         );
  AND2_X1 U2454 ( .A1(n2285), .A2(n2276), .ZN(n2717) );
  INV_X1 U2455 ( .A(IR_REG_24__SCAN_IN), .ZN(n2289) );
  NAND2_X1 U2456 ( .A1(n2269), .A2(n2261), .ZN(n2378) );
  INV_X1 U2457 ( .A(IR_REG_4__SCAN_IN), .ZN(n2268) );
  INV_X1 U2458 ( .A(n3618), .ZN(n3120) );
  OR2_X1 U2459 ( .A1(n2736), .A2(n2723), .ZN(n3387) );
  OR2_X1 U2460 ( .A1(n2736), .A2(n2733), .ZN(n3388) );
  NAND2_X1 U2461 ( .A1(n2200), .A2(n2198), .ZN(n3645) );
  NAND2_X1 U2462 ( .A1(n3641), .A2(n3642), .ZN(n2200) );
  XNOR2_X1 U2463 ( .A(n3092), .B(n2197), .ZN(n4341) );
  XNOR2_X1 U2464 ( .A(n3663), .B(n3672), .ZN(n4372) );
  NOR2_X1 U2465 ( .A1(n4372), .A2(REG1_REG_16__SCAN_IN), .ZN(n4373) );
  OAI21_X1 U2466 ( .B1(n2314), .B2(n4099), .A(n2313), .ZN(n3681) );
  AOI21_X1 U2467 ( .B1(n3728), .B2(n2042), .A(n2121), .ZN(n2187) );
  NAND2_X1 U2468 ( .A1(n2122), .A2(n2036), .ZN(n2121) );
  XNOR2_X1 U2469 ( .A(n3701), .B(n3700), .ZN(n3183) );
  NAND2_X1 U2470 ( .A1(n2120), .A2(n2123), .ZN(n3701) );
  NAND2_X1 U2471 ( .A1(n3728), .A2(n2127), .ZN(n2120) );
  NAND2_X1 U2472 ( .A1(n2089), .A2(n2087), .ZN(n4141) );
  AND2_X1 U2473 ( .A1(n3743), .A2(n2088), .ZN(n2087) );
  NAND2_X1 U2474 ( .A1(n2090), .A2(n4461), .ZN(n2089) );
  OR2_X1 U2475 ( .A1(n3768), .A2(n4443), .ZN(n2088) );
  INV_X1 U2476 ( .A(n3264), .ZN(n2251) );
  INV_X1 U2477 ( .A(IR_REG_22__SCAN_IN), .ZN(n2260) );
  INV_X1 U2478 ( .A(IR_REG_21__SCAN_IN), .ZN(n2259) );
  INV_X1 U2479 ( .A(n2225), .ZN(n2224) );
  OAI21_X1 U2480 ( .B1(n2226), .B2(n3398), .A(n2498), .ZN(n2225) );
  INV_X1 U2481 ( .A(n2541), .ZN(n2543) );
  CLKBUF_X1 U2482 ( .A(n2330), .Z(n2657) );
  NAND2_X1 U2483 ( .A1(n3675), .A2(REG2_REG_18__SCAN_IN), .ZN(n2215) );
  INV_X1 U2484 ( .A(n2779), .ZN(n2160) );
  INV_X1 U2485 ( .A(n3585), .ZN(n2092) );
  INV_X1 U2486 ( .A(n3459), .ZN(n2075) );
  INV_X1 U2487 ( .A(n3458), .ZN(n2076) );
  INV_X1 U2488 ( .A(n4401), .ZN(n2138) );
  INV_X1 U2489 ( .A(n2755), .ZN(n2164) );
  NAND2_X1 U2490 ( .A1(n3825), .A2(n2779), .ZN(n2157) );
  INV_X1 U2491 ( .A(n3969), .ZN(n2838) );
  INV_X1 U2492 ( .A(IR_REG_17__SCAN_IN), .ZN(n2273) );
  NAND2_X1 U2493 ( .A1(n2244), .A2(n2271), .ZN(n2243) );
  INV_X1 U2494 ( .A(n2245), .ZN(n2244) );
  INV_X1 U2495 ( .A(IR_REG_15__SCAN_IN), .ZN(n2523) );
  NAND2_X1 U2496 ( .A1(n2270), .A2(n2246), .ZN(n2245) );
  INV_X1 U2497 ( .A(IR_REG_6__SCAN_IN), .ZN(n2270) );
  INV_X1 U2498 ( .A(IR_REG_5__SCAN_IN), .ZN(n2246) );
  INV_X1 U2499 ( .A(IR_REG_2__SCAN_IN), .ZN(n2267) );
  NOR2_X1 U2500 ( .A1(n2614), .A2(n2613), .ZN(n2623) );
  NAND2_X1 U2501 ( .A1(n2412), .A2(n2413), .ZN(n2414) );
  OAI21_X1 U2502 ( .B1(n2352), .B2(n2132), .A(n2131), .ZN(n4439) );
  INV_X1 U2503 ( .A(n4268), .ZN(n2132) );
  NAND2_X1 U2504 ( .A1(n3396), .A2(n3398), .ZN(n2228) );
  AOI21_X1 U2505 ( .B1(n3335), .B2(n2234), .A(n2233), .ZN(n2232) );
  NOR2_X1 U2506 ( .A1(n2647), .A2(n2648), .ZN(n2233) );
  AND3_X1 U2507 ( .A1(REG3_REG_4__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .A3(
        REG3_REG_5__SCAN_IN), .ZN(n2384) );
  INV_X1 U2508 ( .A(n2547), .ZN(n2548) );
  NOR2_X1 U2509 ( .A1(n3344), .A2(n3345), .ZN(n2111) );
  NAND2_X1 U2510 ( .A1(n3419), .A2(n3420), .ZN(n2105) );
  NOR2_X1 U2511 ( .A1(n2102), .A2(n2101), .ZN(n2100) );
  INV_X1 U2512 ( .A(n3420), .ZN(n2101) );
  INV_X1 U2513 ( .A(n2049), .ZN(n2102) );
  AND2_X1 U2514 ( .A1(n2573), .A2(REG3_REG_19__SCAN_IN), .ZN(n2587) );
  NAND2_X1 U2515 ( .A1(n2587), .A2(REG3_REG_20__SCAN_IN), .ZN(n2614) );
  NAND2_X1 U2516 ( .A1(n3357), .A2(n3358), .ZN(n3355) );
  AND2_X1 U2517 ( .A1(n4258), .A2(n4259), .ZN(n2864) );
  AND2_X1 U2518 ( .A1(REG3_REG_17__SCAN_IN), .A2(n2548), .ZN(n2561) );
  OR2_X1 U2519 ( .A1(n2877), .A2(IR_REG_27__SCAN_IN), .ZN(n2134) );
  NAND2_X1 U2520 ( .A1(n2877), .A2(IR_REG_28__SCAN_IN), .ZN(n2133) );
  AND2_X1 U2521 ( .A1(n2514), .A2(REG3_REG_15__SCAN_IN), .ZN(n2532) );
  INV_X1 U2522 ( .A(n2054), .ZN(n2527) );
  AND4_X1 U2523 ( .A1(n2506), .A2(n2505), .A3(n2504), .A4(n2503), .ZN(n2771)
         );
  AND4_X1 U2524 ( .A1(n2454), .A2(n2453), .A3(n2452), .A4(n2451), .ZN(n3144)
         );
  NAND2_X1 U2525 ( .A1(n2332), .A2(REG0_REG_1__SCAN_IN), .ZN(n2321) );
  NAND2_X1 U2526 ( .A1(n2881), .A2(n4266), .ZN(n2209) );
  AND2_X1 U2527 ( .A1(n2167), .A2(n3082), .ZN(n3085) );
  NAND2_X1 U2528 ( .A1(n3084), .A2(n3083), .ZN(n2167) );
  XNOR2_X1 U2529 ( .A(n2203), .B(n2202), .ZN(n3654) );
  NAND2_X1 U2530 ( .A1(n3654), .A2(REG2_REG_8__SCAN_IN), .ZN(n3653) );
  NAND2_X1 U2531 ( .A1(n4314), .A2(n3090), .ZN(n4324) );
  XNOR2_X1 U2532 ( .A(n3072), .B(n2197), .ZN(n4336) );
  NAND2_X1 U2533 ( .A1(n4336), .A2(REG2_REG_12__SCAN_IN), .ZN(n4335) );
  NAND2_X1 U2534 ( .A1(n4352), .A2(n3094), .ZN(n3660) );
  NAND2_X1 U2535 ( .A1(n4386), .A2(n3915), .ZN(n2216) );
  INV_X1 U2536 ( .A(n2215), .ZN(n2211) );
  INV_X1 U2537 ( .A(n2216), .ZN(n2214) );
  NAND2_X1 U2538 ( .A1(n2124), .A2(n3700), .ZN(n2122) );
  INV_X1 U2539 ( .A(n3716), .ZN(n2129) );
  NOR2_X1 U2540 ( .A1(n2791), .A2(n2128), .ZN(n2127) );
  INV_X1 U2541 ( .A(n2789), .ZN(n2128) );
  AND2_X1 U2542 ( .A1(n2822), .A2(n2725), .ZN(n3210) );
  XNOR2_X1 U2543 ( .A(n3739), .B(n2091), .ZN(n2090) );
  INV_X1 U2544 ( .A(n3740), .ZN(n2091) );
  AND4_X1 U2545 ( .A1(n2619), .A2(n2618), .A3(n2617), .A4(n2616), .ZN(n3795)
         );
  OR2_X1 U2546 ( .A1(n3765), .A2(n3554), .ZN(n3789) );
  AND2_X1 U2547 ( .A1(n2195), .A2(n3820), .ZN(n2194) );
  NAND2_X1 U2548 ( .A1(n2095), .A2(n2093), .ZN(n3846) );
  AND4_X1 U2549 ( .A1(n2566), .A2(n2565), .A3(n2564), .A4(n2563), .ZN(n3904)
         );
  NAND2_X1 U2550 ( .A1(n2095), .A2(n3579), .ZN(n3902) );
  NAND2_X1 U2551 ( .A1(n2146), .A2(n2148), .ZN(n3920) );
  INV_X1 U2552 ( .A(n2149), .ZN(n2148) );
  OAI21_X1 U2553 ( .B1(n2151), .B2(n2150), .A(n2773), .ZN(n2149) );
  AND4_X1 U2554 ( .A1(n2553), .A2(n2552), .A3(n2551), .A4(n2550), .ZN(n3923)
         );
  AND4_X1 U2555 ( .A1(n2537), .A2(n2536), .A3(n2535), .A4(n2534), .ZN(n3942)
         );
  INV_X1 U2556 ( .A(n2193), .ZN(n2191) );
  INV_X1 U2557 ( .A(REG3_REG_13__SCAN_IN), .ZN(n2478) );
  OR2_X1 U2558 ( .A1(n2479), .A2(n2478), .ZN(n2501) );
  INV_X1 U2559 ( .A(REG3_REG_11__SCAN_IN), .ZN(n2448) );
  NAND2_X1 U2560 ( .A1(n2073), .A2(n3457), .ZN(n4402) );
  NAND2_X1 U2561 ( .A1(n3142), .A2(n3458), .ZN(n2073) );
  INV_X1 U2562 ( .A(REG3_REG_10__SCAN_IN), .ZN(n4059) );
  OR2_X1 U2563 ( .A1(n2434), .A2(n4059), .ZN(n2449) );
  INV_X1 U2564 ( .A(n4464), .ZN(n4441) );
  OR2_X1 U2565 ( .A1(n2424), .A2(n3119), .ZN(n2434) );
  INV_X1 U2566 ( .A(n3055), .ZN(n3030) );
  AND4_X1 U2567 ( .A1(n2404), .A2(n2403), .A3(n2402), .A4(n2401), .ZN(n3011)
         );
  NOR2_X1 U2568 ( .A1(n2085), .A2(n2795), .ZN(n2084) );
  OR2_X1 U2569 ( .A1(n2992), .A2(n3349), .ZN(n2993) );
  NAND2_X1 U2570 ( .A1(n2941), .A2(n3475), .ZN(n2997) );
  INV_X1 U2571 ( .A(n4461), .ZN(n4409) );
  AND2_X1 U2572 ( .A1(n3469), .A2(n3471), .ZN(n2960) );
  NOR2_X1 U2573 ( .A1(n3983), .A2(n3984), .ZN(n3982) );
  NOR3_X1 U2574 ( .A1(n3797), .A2(n3338), .A3(n3757), .ZN(n3758) );
  OR2_X1 U2575 ( .A1(n3796), .A2(n3791), .ZN(n3797) );
  AND2_X1 U2576 ( .A1(n3892), .A2(n2195), .ZN(n3833) );
  NAND2_X1 U2577 ( .A1(n3892), .A2(n2038), .ZN(n3853) );
  AND2_X1 U2578 ( .A1(n3909), .A2(n3891), .ZN(n3892) );
  NAND2_X1 U2579 ( .A1(n3892), .A2(n3876), .ZN(n3875) );
  NOR2_X1 U2580 ( .A1(n3927), .A2(n3328), .ZN(n3909) );
  OR2_X1 U2581 ( .A1(n3949), .A2(n3309), .ZN(n3927) );
  NOR2_X1 U2582 ( .A1(n4416), .A2(n2192), .ZN(n3968) );
  NAND2_X1 U2583 ( .A1(n2838), .A2(n2193), .ZN(n2192) );
  OR2_X1 U2584 ( .A1(n3099), .A2(n3050), .ZN(n3138) );
  NOR2_X1 U2585 ( .A1(n3138), .A2(n3240), .ZN(n4418) );
  OR2_X1 U2586 ( .A1(n3035), .A2(n3269), .ZN(n3099) );
  NOR2_X1 U2587 ( .A1(n2993), .A2(n3317), .ZN(n3015) );
  AND2_X1 U2588 ( .A1(n3015), .A2(n3010), .ZN(n3034) );
  NOR2_X1 U2589 ( .A1(n4452), .A2(n2964), .ZN(n4516) );
  NAND2_X1 U2590 ( .A1(n2189), .A2(IR_REG_31__SCAN_IN), .ZN(n2877) );
  NAND2_X1 U2591 ( .A1(n2285), .A2(n2190), .ZN(n2189) );
  INV_X1 U2592 ( .A(IR_REG_26__SCAN_IN), .ZN(n2190) );
  NAND2_X1 U2593 ( .A1(n2718), .A2(n2275), .ZN(n2287) );
  INV_X1 U2594 ( .A(n2285), .ZN(n2302) );
  OR3_X1 U2595 ( .A1(n2286), .A2(n2718), .A3(n2275), .ZN(n2288) );
  OAI21_X1 U2596 ( .B1(n2708), .B2(n2707), .A(n2706), .ZN(n2863) );
  INV_X1 U2597 ( .A(IR_REG_20__SCAN_IN), .ZN(n2294) );
  OR2_X1 U2598 ( .A1(n2488), .A2(n2487), .ZN(n2507) );
  NOR2_X1 U2599 ( .A1(IR_REG_11__SCAN_IN), .A2(IR_REG_10__SCAN_IN), .ZN(n2486)
         );
  OR2_X1 U2600 ( .A1(n2488), .A2(IR_REG_10__SCAN_IN), .ZN(n2455) );
  NAND2_X1 U2601 ( .A1(n2104), .A2(n3420), .ZN(n3060) );
  OR2_X1 U2602 ( .A1(n3418), .A2(n3419), .ZN(n2104) );
  CLKBUF_X1 U2603 ( .A(n3237), .Z(n3238) );
  INV_X1 U2604 ( .A(n2114), .ZN(n3246) );
  OAI21_X1 U2605 ( .B1(n3411), .B2(n3408), .A(n3409), .ZN(n3255) );
  INV_X1 U2606 ( .A(n4439), .ZN(n4453) );
  NAND2_X1 U2607 ( .A1(n3229), .A2(n2645), .ZN(n3334) );
  NAND2_X1 U2608 ( .A1(n2099), .A2(n2103), .ZN(n3117) );
  INV_X1 U2609 ( .A(n2837), .ZN(n4460) );
  AND4_X1 U2610 ( .A1(n2605), .A2(n2604), .A3(n2603), .A4(n2602), .ZN(n3849)
         );
  INV_X1 U2611 ( .A(n2781), .ZN(n3820) );
  INV_X1 U2612 ( .A(n2239), .ZN(n2238) );
  AOI21_X1 U2613 ( .B1(n2239), .B2(n2237), .A(n2059), .ZN(n2236) );
  AND2_X1 U2614 ( .A1(n3359), .A2(n2609), .ZN(n2239) );
  INV_X1 U2615 ( .A(n2964), .ZN(n2970) );
  INV_X1 U2616 ( .A(n3389), .ZN(n3448) );
  INV_X1 U2617 ( .A(n3387), .ZN(n3446) );
  NOR2_X1 U2618 ( .A1(n2029), .A2(n2716), .ZN(n3604) );
  INV_X1 U2619 ( .A(n3795), .ZN(n3830) );
  INV_X1 U2620 ( .A(n3923), .ZN(n3614) );
  INV_X1 U2621 ( .A(n3942), .ZN(n3906) );
  INV_X1 U2622 ( .A(n2771), .ZN(n3944) );
  INV_X1 U2623 ( .A(n3144), .ZN(n3616) );
  INV_X1 U2624 ( .A(n3011), .ZN(n3619) );
  NAND2_X1 U2625 ( .A1(n2398), .A2(REG0_REG_3__SCAN_IN), .ZN(n2350) );
  NAND4_X1 U2626 ( .A1(n2284), .A2(n2283), .A3(n2282), .A4(n2281), .ZN(n3625)
         );
  NAND2_X1 U2627 ( .A1(n2332), .A2(REG0_REG_0__SCAN_IN), .ZN(n2284) );
  OR2_X1 U2628 ( .A1(n2849), .A2(n2859), .ZN(n3624) );
  NAND2_X1 U2629 ( .A1(n2876), .A2(n2875), .ZN(n4280) );
  OAI21_X1 U2630 ( .B1(n4268), .B2(n2880), .A(n2201), .ZN(n3626) );
  NAND2_X1 U2631 ( .A1(n4268), .A2(n2880), .ZN(n2201) );
  NAND2_X1 U2632 ( .A1(n2178), .A2(n2174), .ZN(n2173) );
  NOR2_X1 U2633 ( .A1(n2918), .A2(n2043), .ZN(n4284) );
  XNOR2_X1 U2634 ( .A(n2883), .B(n4501), .ZN(n4300) );
  NAND2_X1 U2635 ( .A1(n4300), .A2(REG2_REG_6__SCAN_IN), .ZN(n4299) );
  XNOR2_X1 U2636 ( .A(n3085), .B(n2202), .ZN(n3651) );
  NAND2_X1 U2637 ( .A1(n3651), .A2(REG1_REG_8__SCAN_IN), .ZN(n3650) );
  INV_X1 U2638 ( .A(n4494), .ZN(n4331) );
  NAND2_X1 U2639 ( .A1(n4340), .A2(n3093), .ZN(n4353) );
  NAND2_X1 U2640 ( .A1(n4353), .A2(n4354), .ZN(n4352) );
  XNOR2_X1 U2641 ( .A(n3660), .B(n3095), .ZN(n3096) );
  AND2_X1 U2642 ( .A1(n2205), .A2(n2208), .ZN(n3668) );
  NOR2_X1 U2643 ( .A1(n3669), .A2(n3076), .ZN(n2205) );
  NAND2_X1 U2644 ( .A1(n2208), .A2(REG2_REG_14__SCAN_IN), .ZN(n2207) );
  NAND2_X1 U2645 ( .A1(n4377), .A2(n2216), .ZN(n4388) );
  NAND2_X1 U2646 ( .A1(n2212), .A2(n2067), .ZN(n3678) );
  AND2_X1 U2647 ( .A1(n2680), .A2(n2724), .ZN(n3723) );
  OAI21_X1 U2648 ( .B1(n3728), .B2(n2790), .A(n2789), .ZN(n3711) );
  NAND2_X1 U2649 ( .A1(n2152), .A2(n2151), .ZN(n3938) );
  NAND2_X1 U2650 ( .A1(n3162), .A2(n2153), .ZN(n2152) );
  NAND2_X1 U2651 ( .A1(n2154), .A2(n2769), .ZN(n3958) );
  OR2_X1 U2652 ( .A1(n3162), .A2(n2770), .ZN(n2154) );
  OR2_X1 U2653 ( .A1(n3101), .A2(n2142), .ZN(n2136) );
  NAND2_X1 U2654 ( .A1(n2139), .A2(n2144), .ZN(n3141) );
  NAND2_X1 U2655 ( .A1(n3101), .A2(n2031), .ZN(n2139) );
  NAND2_X1 U2656 ( .A1(n2145), .A2(n2763), .ZN(n3049) );
  OR2_X1 U2657 ( .A1(n3101), .A2(n2764), .ZN(n2145) );
  NAND2_X1 U2658 ( .A1(n2977), .A2(n2976), .ZN(n3808) );
  OR2_X1 U2659 ( .A1(n2862), .A2(n2731), .ZN(n4413) );
  INV_X1 U2660 ( .A(REG2_REG_2__SCAN_IN), .ZN(n4105) );
  AND2_X1 U2661 ( .A1(n3894), .A2(n4540), .ZN(n4455) );
  INV_X1 U2662 ( .A(n4413), .ZN(n4466) );
  INV_X2 U2663 ( .A(n4576), .ZN(n4579) );
  OR2_X1 U2664 ( .A1(n2844), .A2(n2946), .ZN(n4576) );
  INV_X1 U2665 ( .A(n2185), .ZN(n2184) );
  NOR2_X1 U2666 ( .A1(n4141), .A2(n2086), .ZN(n4143) );
  AND2_X1 U2667 ( .A1(n4142), .A2(n4540), .ZN(n2086) );
  INV_X2 U2668 ( .A(n4558), .ZN(n4560) );
  NAND2_X1 U2669 ( .A1(n2855), .A2(n2854), .ZN(n4480) );
  AND2_X1 U2670 ( .A1(n2256), .A2(n2255), .ZN(n2254) );
  INV_X1 U2671 ( .A(IR_REG_29__SCAN_IN), .ZN(n2255) );
  INV_X1 U2672 ( .A(n2280), .ZN(n2852) );
  NOR2_X1 U2673 ( .A1(n2722), .A2(n2721), .ZN(n4256) );
  NAND2_X1 U2674 ( .A1(n2706), .A2(IR_REG_31__SCAN_IN), .ZN(n2290) );
  AND2_X1 U2675 ( .A1(n2863), .A2(STATE_REG_SCAN_IN), .ZN(n4481) );
  INV_X1 U2676 ( .A(n3681), .ZN(n4261) );
  AND2_X1 U2677 ( .A1(n2408), .A2(n2421), .ZN(n4264) );
  NAND2_X1 U2678 ( .A1(IR_REG_31__SCAN_IN), .A2(n2219), .ZN(n2199) );
  NAND2_X1 U2679 ( .A1(n2183), .A2(n2220), .ZN(n2219) );
  OR2_X1 U2680 ( .A1(n3175), .A2(n4193), .ZN(n2847) );
  OR2_X1 U2681 ( .A1(n3849), .A2(n3835), .ZN(n2030) );
  INV_X2 U2682 ( .A(IR_REG_31__SCAN_IN), .ZN(n2718) );
  AND2_X1 U2683 ( .A1(n2763), .A2(n2044), .ZN(n2031) );
  AND2_X1 U2684 ( .A1(n4377), .A2(n2066), .ZN(n2032) );
  AND3_X1 U2685 ( .A1(n2257), .A2(n2274), .A3(n2053), .ZN(n2033) );
  NAND2_X1 U2686 ( .A1(n2105), .A2(n2252), .ZN(n2034) );
  INV_X1 U2687 ( .A(n3457), .ZN(n2077) );
  NAND2_X1 U2688 ( .A1(n2771), .A2(n2838), .ZN(n2035) );
  OR2_X1 U2689 ( .A1(n2129), .A2(n3207), .ZN(n2036) );
  OR3_X1 U2690 ( .A1(n3338), .A2(n3757), .A3(n3741), .ZN(n2037) );
  AND2_X1 U2691 ( .A1(n3876), .A2(n3854), .ZN(n2038) );
  INV_X1 U2692 ( .A(n3671), .ZN(n4490) );
  AND2_X1 U2693 ( .A1(n2538), .A2(n2525), .ZN(n3671) );
  INV_X1 U2694 ( .A(IR_REG_1__SCAN_IN), .ZN(n2183) );
  AND2_X1 U2695 ( .A1(n2896), .A2(n2209), .ZN(n2039) );
  OR2_X1 U2696 ( .A1(n2296), .A2(IR_REG_21__SCAN_IN), .ZN(n2040) );
  NAND2_X2 U2697 ( .A1(n2849), .A2(n2951), .ZN(n2339) );
  AND2_X1 U2698 ( .A1(n2372), .A2(n2371), .ZN(n2041) );
  AND3_X1 U2699 ( .A1(n2242), .A2(n2241), .A3(n2273), .ZN(n2292) );
  NOR2_X1 U2700 ( .A1(n4255), .A2(n2280), .ZN(n2331) );
  NAND2_X1 U2701 ( .A1(n2229), .A2(n2232), .ZN(n3292) );
  AND2_X1 U2702 ( .A1(n4255), .A2(n2280), .ZN(n2346) );
  AND2_X1 U2703 ( .A1(n2292), .A2(n2033), .ZN(n2286) );
  OAI21_X1 U2704 ( .B1(n3411), .B2(n2108), .A(n2106), .ZN(n3357) );
  NOR2_X1 U2705 ( .A1(n2378), .A2(IR_REG_5__SCAN_IN), .ZN(n2389) );
  AND2_X1 U2706 ( .A1(n3700), .A2(n2127), .ZN(n2042) );
  AND2_X1 U2707 ( .A1(n2182), .A2(n4265), .ZN(n2043) );
  OR2_X1 U2708 ( .A1(n3617), .A2(n3050), .ZN(n2044) );
  NOR2_X1 U2709 ( .A1(n3235), .A2(n3236), .ZN(n2045) );
  OAI21_X1 U2710 ( .B1(n3357), .B2(n2238), .A(n2236), .ZN(n3383) );
  OR2_X1 U2711 ( .A1(n4292), .A2(n2988), .ZN(n2046) );
  AND4_X1 U2712 ( .A1(n2336), .A2(n2335), .A3(n2334), .A4(n2333), .ZN(n2753)
         );
  AND2_X1 U2713 ( .A1(n2802), .A2(n3143), .ZN(n2047) );
  INV_X1 U2714 ( .A(n2081), .ZN(n2080) );
  OAI21_X1 U2715 ( .B1(n2082), .B2(n2799), .A(n3494), .ZN(n2081) );
  NAND2_X1 U2716 ( .A1(n3067), .A2(n2204), .ZN(n2203) );
  NOR2_X1 U2717 ( .A1(n3104), .A2(n3121), .ZN(n2048) );
  AND2_X1 U2718 ( .A1(n2249), .A2(n2248), .ZN(n2049) );
  INV_X1 U2719 ( .A(n2124), .ZN(n2123) );
  OAI21_X1 U2720 ( .B1(n2126), .B2(n2125), .A(n2130), .ZN(n2124) );
  AND2_X1 U2721 ( .A1(n2157), .A2(n2030), .ZN(n2050) );
  AND2_X1 U2722 ( .A1(n3355), .A2(n3359), .ZN(n2051) );
  AND2_X1 U2723 ( .A1(n2093), .A2(n2092), .ZN(n2052) );
  AND2_X1 U2724 ( .A1(n2707), .A2(n2289), .ZN(n2053) );
  INV_X1 U2725 ( .A(n2175), .ZN(n2174) );
  NAND2_X1 U2726 ( .A1(n2180), .A2(REG1_REG_1__SCAN_IN), .ZN(n2175) );
  AND2_X1 U2727 ( .A1(n2279), .A2(n2280), .ZN(n2332) );
  INV_X1 U2728 ( .A(n4263), .ZN(n2202) );
  NAND2_X1 U2729 ( .A1(n2228), .A2(n3397), .ZN(n3282) );
  INV_X1 U2730 ( .A(n3217), .ZN(n2223) );
  NOR2_X1 U2731 ( .A1(n2378), .A2(n2245), .ZN(n2391) );
  NAND2_X1 U2732 ( .A1(n2242), .A2(n2240), .ZN(n2430) );
  OAI21_X1 U2733 ( .B1(n2546), .B2(n2545), .A(n2544), .ZN(n3323) );
  NAND2_X1 U2734 ( .A1(n2136), .A2(n2140), .ZN(n4400) );
  NAND2_X1 U2735 ( .A1(n3059), .A2(n2414), .ZN(n3263) );
  NAND2_X1 U2736 ( .A1(n3237), .A2(n2447), .ZN(n3396) );
  XNOR2_X1 U2737 ( .A(n2687), .B(n2526), .ZN(n2054) );
  NOR2_X1 U2738 ( .A1(n3074), .A2(n3095), .ZN(n3669) );
  INV_X1 U2739 ( .A(n2783), .ZN(n2161) );
  AND2_X1 U2740 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_29__SCAN_IN), .ZN(n2055)
         );
  OR2_X1 U2741 ( .A1(n4331), .A2(n4412), .ZN(n2056) );
  INV_X1 U2742 ( .A(IR_REG_28__SCAN_IN), .ZN(n2303) );
  OR2_X1 U2743 ( .A1(n3797), .A2(n3338), .ZN(n2057) );
  AND2_X1 U2744 ( .A1(n2586), .A2(n2585), .ZN(n2058) );
  AND2_X1 U2745 ( .A1(n2611), .A2(n2610), .ZN(n2059) );
  NAND2_X1 U2746 ( .A1(n3199), .A2(n3434), .ZN(n2060) );
  NAND2_X1 U2747 ( .A1(n2155), .A2(n3957), .ZN(n2061) );
  INV_X1 U2748 ( .A(n2247), .ZN(n3059) );
  NOR2_X1 U2749 ( .A1(n3060), .A2(n3061), .ZN(n2247) );
  INV_X1 U2750 ( .A(n2772), .ZN(n2150) );
  OR2_X1 U2751 ( .A1(n3963), .A2(n3447), .ZN(n2772) );
  INV_X1 U2752 ( .A(n3091), .ZN(n2197) );
  XNOR2_X1 U2753 ( .A(n2291), .B(IR_REG_26__SCAN_IN), .ZN(n2692) );
  INV_X1 U2754 ( .A(n3408), .ZN(n2109) );
  OR2_X1 U2755 ( .A1(n4416), .A2(n2191), .ZN(n2062) );
  XNOR2_X1 U2756 ( .A(n2290), .B(n2289), .ZN(n2690) );
  INV_X1 U2757 ( .A(n3490), .ZN(n2079) );
  INV_X1 U2758 ( .A(n3461), .ZN(n2072) );
  OR2_X1 U2759 ( .A1(n4416), .A2(n3286), .ZN(n2063) );
  OR2_X1 U2760 ( .A1(n4331), .A2(n4577), .ZN(n2064) );
  NAND2_X1 U2761 ( .A1(n2242), .A2(n2241), .ZN(n2065) );
  INV_X1 U2762 ( .A(n2110), .ZN(n3343) );
  NAND2_X1 U2763 ( .A1(n2112), .A2(n2111), .ZN(n2110) );
  NAND2_X1 U2764 ( .A1(n2708), .A2(n2707), .ZN(n2706) );
  INV_X2 U2765 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  AND2_X2 U2766 ( .A1(n2950), .A2(n4413), .ZN(n4471) );
  NOR2_X1 U2767 ( .A1(n4389), .A2(n2214), .ZN(n2066) );
  INV_X1 U2768 ( .A(n3394), .ZN(n3434) );
  OR2_X1 U2769 ( .A1(n2066), .A2(n2211), .ZN(n2067) );
  INV_X1 U2770 ( .A(n4266), .ZN(n2210) );
  NAND2_X1 U2771 ( .A1(n3142), .A2(n2074), .ZN(n2070) );
  NAND2_X1 U2772 ( .A1(n2070), .A2(n2071), .ZN(n3127) );
  OAI21_X1 U2773 ( .B1(n3029), .B2(n2800), .A(n3489), .ZN(n3102) );
  INV_X1 U2774 ( .A(n3489), .ZN(n2082) );
  NAND2_X1 U2775 ( .A1(n2941), .A2(n2084), .ZN(n2796) );
  NAND2_X1 U2776 ( .A1(n3922), .A2(n3921), .ZN(n2095) );
  NAND2_X1 U2777 ( .A1(n2095), .A2(n2052), .ZN(n2814) );
  NAND2_X1 U2778 ( .A1(n3418), .A2(n2100), .ZN(n2099) );
  NOR2_X2 U2779 ( .A1(n2930), .A2(n2928), .ZN(n2929) );
  OAI21_X2 U2780 ( .B1(n3396), .B2(n2226), .A(n2224), .ZN(n3219) );
  NAND4_X1 U2781 ( .A1(n2119), .A2(n2118), .A3(n2117), .A4(n2116), .ZN(n2272)
         );
  NAND2_X1 U2782 ( .A1(n2352), .A2(DATAI_1_), .ZN(n2131) );
  NAND3_X4 U2783 ( .A1(n2134), .A2(n2133), .A3(n2304), .ZN(n2352) );
  NAND2_X1 U2784 ( .A1(n2135), .A2(n2137), .ZN(n2767) );
  NAND2_X1 U2785 ( .A1(n3101), .A2(n2140), .ZN(n2135) );
  NAND2_X1 U2786 ( .A1(n3162), .A2(n2147), .ZN(n2146) );
  AOI21_X2 U2787 ( .B1(n3773), .B2(n2785), .A(n2784), .ZN(n3746) );
  NOR2_X1 U2788 ( .A1(n2782), .A2(n3814), .ZN(n2162) );
  NAND2_X1 U2789 ( .A1(n3532), .A2(n2166), .ZN(n2165) );
  NAND2_X1 U2790 ( .A1(n2756), .A2(n2755), .ZN(n2166) );
  NAND3_X1 U2791 ( .A1(n3532), .A2(n2166), .A3(n2164), .ZN(n2163) );
  OAI21_X1 U2792 ( .B1(n2936), .B2(n2756), .A(n2755), .ZN(n2995) );
  AOI22_X1 U2793 ( .A1(n3861), .A2(n2778), .B1(n3258), .B2(n3887), .ZN(n3844)
         );
  AOI21_X1 U2794 ( .B1(n3883), .B2(n3885), .A(n2776), .ZN(n3861) );
  OAI21_X1 U2795 ( .B1(n3008), .B2(n2760), .A(n2759), .ZN(n3040) );
  AOI22_X1 U2796 ( .A1(n3920), .A2(n3558), .B1(n3309), .B2(n3906), .ZN(n3901)
         );
  NAND2_X1 U2797 ( .A1(n2959), .A2(n2754), .ZN(n2936) );
  NAND2_X1 U2798 ( .A1(n2752), .A2(n3530), .ZN(n2959) );
  NAND2_X1 U2799 ( .A1(n4445), .A2(n2750), .ZN(n2961) );
  NAND2_X1 U2800 ( .A1(n4327), .A2(n4328), .ZN(n4326) );
  NAND2_X1 U2801 ( .A1(n4288), .A2(n4289), .ZN(n4287) );
  NOR2_X2 U2802 ( .A1(n4294), .A2(n2874), .ZN(n3084) );
  NAND4_X1 U2803 ( .A1(n2168), .A2(n2176), .A3(n2169), .A4(REG1_REG_1__SCAN_IN), .ZN(n2171) );
  NAND3_X1 U2804 ( .A1(n2172), .A2(n2171), .A3(n3629), .ZN(n3628) );
  NAND3_X1 U2805 ( .A1(n2175), .A2(n2176), .A3(n2178), .ZN(n2172) );
  OAI211_X1 U2806 ( .C1(n2178), .C2(REG1_REG_1__SCAN_IN), .A(n2173), .B(n2176), 
        .ZN(n3630) );
  NAND2_X1 U2807 ( .A1(n2183), .A2(IR_REG_31__SCAN_IN), .ZN(n2179) );
  NAND3_X1 U2808 ( .A1(n2183), .A2(n2220), .A3(n2267), .ZN(n2351) );
  NAND2_X1 U2809 ( .A1(n2186), .A2(n2184), .ZN(n4211) );
  OAI21_X1 U2810 ( .B1(n3992), .B2(n2841), .A(n3993), .ZN(n2185) );
  NAND2_X1 U2811 ( .A1(n3991), .A2(n4550), .ZN(n2186) );
  XNOR2_X1 U2812 ( .A(n2187), .B(n3702), .ZN(n3991) );
  OR2_X1 U2813 ( .A1(n3706), .A2(n3705), .ZN(n2188) );
  NOR3_X4 U2814 ( .A1(n3797), .A2(n3722), .A3(n2037), .ZN(n3720) );
  NAND2_X1 U2815 ( .A1(n3892), .A2(n2194), .ZN(n3796) );
  AND4_X2 U2816 ( .A1(n2033), .A2(n2242), .A3(n2241), .A4(n2196), .ZN(n2285)
         );
  MUX2_X1 U2817 ( .A(REG2_REG_2__SCAN_IN), .B(n4105), .S(n4267), .Z(n2198) );
  XNOR2_X2 U2818 ( .A(n2199), .B(IR_REG_2__SCAN_IN), .ZN(n4267) );
  INV_X1 U2819 ( .A(n3669), .ZN(n2206) );
  NAND2_X1 U2820 ( .A1(n2206), .A2(n2208), .ZN(n3075) );
  NAND2_X1 U2821 ( .A1(n4376), .A2(n2213), .ZN(n2212) );
  NAND2_X1 U2822 ( .A1(n4376), .A2(n4378), .ZN(n4377) );
  OAI211_X1 U2823 ( .C1(n2218), .C2(n2060), .A(n2217), .B(n3215), .ZN(U3217)
         );
  NAND2_X1 U2824 ( .A1(n2218), .A2(n2265), .ZN(n2217) );
  NAND2_X1 U2825 ( .A1(n3189), .A2(n3188), .ZN(n2218) );
  NAND2_X1 U2826 ( .A1(n2221), .A2(n2222), .ZN(n2510) );
  NAND2_X1 U2827 ( .A1(n3396), .A2(n2224), .ZN(n2221) );
  NAND2_X1 U2828 ( .A1(n3226), .A2(n2230), .ZN(n2229) );
  NAND2_X1 U2829 ( .A1(n2285), .A2(n2256), .ZN(n2720) );
  NAND2_X1 U2830 ( .A1(n2285), .A2(n2254), .ZN(n2278) );
  NAND2_X1 U2831 ( .A1(n2292), .A2(n2274), .ZN(n2296) );
  AND2_X1 U2832 ( .A1(n3625), .A2(n2837), .ZN(n4446) );
  XNOR2_X1 U2833 ( .A(n3431), .B(n2266), .ZN(n3435) );
  AND2_X1 U2834 ( .A1(n2352), .A2(DATAI_30_), .ZN(n3984) );
  AND2_X1 U2835 ( .A1(n2352), .A2(DATAI_23_), .ZN(n3791) );
  AND2_X1 U2836 ( .A1(n2352), .A2(DATAI_21_), .ZN(n3829) );
  NAND2_X1 U2837 ( .A1(n2352), .A2(DATAI_28_), .ZN(n3207) );
  NAND2_X1 U2838 ( .A1(n2352), .A2(DATAI_26_), .ZN(n2839) );
  NAND2_X1 U2839 ( .A1(n2352), .A2(DATAI_24_), .ZN(n3774) );
  MUX2_X2 U2840 ( .A(REG1_REG_26__SCAN_IN), .B(n4213), .S(n4579), .Z(n4145) );
  INV_X1 U2841 ( .A(n2748), .ZN(n2749) );
  XNOR2_X1 U2842 ( .A(n2326), .B(n2327), .ZN(n2922) );
  OAI21_X1 U2843 ( .B1(n2342), .B2(n2341), .A(n2343), .ZN(n2930) );
  AND2_X2 U2844 ( .A1(n2741), .A2(STATE_REG_SCAN_IN), .ZN(n3450) );
  NAND2_X1 U2845 ( .A1(n2622), .A2(n2621), .ZN(n3226) );
  INV_X1 U2846 ( .A(IR_REG_30__SCAN_IN), .ZN(n3184) );
  INV_X1 U2847 ( .A(n3115), .ZN(n3116) );
  AND2_X1 U2848 ( .A1(n2268), .A2(n2363), .ZN(n2261) );
  OR2_X1 U2849 ( .A1(n2749), .A2(n2330), .ZN(n2262) );
  OR2_X1 U2850 ( .A1(n3768), .A2(n2787), .ZN(n2263) );
  INV_X1 U2851 ( .A(n3447), .ZN(n3947) );
  OR2_X1 U2852 ( .A1(n3614), .A2(n3328), .ZN(n2264) );
  AND3_X1 U2853 ( .A1(n3214), .A2(n3213), .A3(n3434), .ZN(n2265) );
  AND2_X1 U2854 ( .A1(n2352), .A2(DATAI_25_), .ZN(n3757) );
  AND2_X1 U2855 ( .A1(n3433), .A2(n3432), .ZN(n2266) );
  INV_X1 U2856 ( .A(n3768), .ZN(n3610) );
  OAI22_X1 U2857 ( .A1(n2923), .A2(n2922), .B1(n2329), .B2(n2328), .ZN(n2928)
         );
  INV_X1 U2858 ( .A(n2583), .ZN(n2586) );
  AND2_X1 U2859 ( .A1(n2647), .A2(n2648), .ZN(n2645) );
  INV_X1 U2860 ( .A(n3757), .ZN(n2787) );
  NAND2_X1 U2861 ( .A1(n2543), .A2(n2542), .ZN(n2544) );
  NAND2_X1 U2862 ( .A1(n2303), .A2(IR_REG_27__SCAN_IN), .ZN(n2304) );
  INV_X1 U2863 ( .A(REG3_REG_14__SCAN_IN), .ZN(n2500) );
  INV_X1 U2864 ( .A(REG3_REG_7__SCAN_IN), .ZN(n4039) );
  AND2_X1 U2865 ( .A1(n3756), .A2(n3774), .ZN(n2784) );
  AND2_X1 U2866 ( .A1(n2352), .A2(DATAI_22_), .ZN(n2781) );
  NAND2_X1 U2867 ( .A1(n3963), .A2(n3447), .ZN(n2773) );
  NOR2_X1 U2868 ( .A1(n2449), .A2(n2448), .ZN(n2463) );
  INV_X1 U2869 ( .A(n3402), .ZN(n4417) );
  AND2_X1 U2870 ( .A1(n4256), .A2(n2864), .ZN(n4407) );
  NOR2_X1 U2871 ( .A1(n2501), .A2(n2500), .ZN(n2514) );
  OR2_X1 U2872 ( .A1(n2638), .A2(n2637), .ZN(n2650) );
  AND2_X1 U2873 ( .A1(n2561), .A2(REG3_REG_18__SCAN_IN), .ZN(n2573) );
  INV_X1 U2874 ( .A(n3424), .ZN(n3389) );
  INV_X1 U2875 ( .A(REG3_REG_9__SCAN_IN), .ZN(n3119) );
  INV_X1 U2876 ( .A(n4403), .ZN(n4440) );
  INV_X1 U2877 ( .A(n3753), .ZN(n3719) );
  OR2_X1 U2878 ( .A1(n3753), .A2(n3741), .ZN(n2789) );
  AND2_X1 U2879 ( .A1(n3787), .A2(n2780), .ZN(n3814) );
  INV_X1 U2880 ( .A(n3558), .ZN(n3921) );
  INV_X1 U2881 ( .A(n4407), .ZN(n4443) );
  INV_X1 U2882 ( .A(n3567), .ZN(n3978) );
  INV_X1 U2883 ( .A(n3886), .ZN(n3891) );
  NAND2_X1 U2884 ( .A1(n2827), .A2(n2864), .ZN(n4464) );
  OR2_X1 U2885 ( .A1(n2430), .A2(IR_REG_9__SCAN_IN), .ZN(n2488) );
  AND2_X1 U2886 ( .A1(n2743), .A2(n2742), .ZN(n2744) );
  AND2_X1 U2887 ( .A1(n2317), .A2(n2316), .ZN(n2923) );
  AND2_X1 U2888 ( .A1(n2662), .A2(n2651), .ZN(n3760) );
  INV_X1 U2889 ( .A(n3774), .ZN(n3338) );
  INV_X1 U2890 ( .A(n3854), .ZN(n3362) );
  OR2_X1 U2891 ( .A1(n2946), .A2(n2705), .ZN(n2736) );
  INV_X1 U2892 ( .A(n2839), .ZN(n3741) );
  AND4_X1 U2893 ( .A1(n2655), .A2(n2654), .A3(n2653), .A4(n2652), .ZN(n3768)
         );
  AND4_X1 U2894 ( .A1(n2628), .A2(n2627), .A3(n2626), .A4(n2625), .ZN(n3816)
         );
  AND2_X1 U2895 ( .A1(n2352), .A2(n2865), .ZN(n2875) );
  INV_X1 U2896 ( .A(n4293), .ZN(n4394) );
  OR2_X1 U2897 ( .A1(n3686), .A2(n3687), .ZN(n3700) );
  INV_X1 U2898 ( .A(n4455), .ZN(n3952) );
  INV_X1 U2899 ( .A(n4448), .ZN(n4462) );
  INV_X1 U2900 ( .A(n4471), .ZN(n3935) );
  NAND2_X1 U2901 ( .A1(n2821), .A2(n2820), .ZN(n4461) );
  OAI22_X1 U2902 ( .A1(n2854), .A2(D_REG_0__SCAN_IN), .B1(n2856), .B2(n2692), 
        .ZN(n2946) );
  INV_X1 U2903 ( .A(n3240), .ZN(n3143) );
  NAND2_X1 U2904 ( .A1(n4448), .A2(n4524), .ZN(n4550) );
  INV_X1 U2905 ( .A(n4481), .ZN(n2859) );
  AND2_X1 U2906 ( .A1(n2432), .A2(n2488), .ZN(n3081) );
  AND2_X1 U2907 ( .A1(n2876), .A2(n2866), .ZN(n4392) );
  OR2_X1 U2908 ( .A1(n2736), .A2(n2712), .ZN(n3394) );
  NAND2_X1 U2909 ( .A1(n3435), .A2(n3434), .ZN(n3441) );
  NAND4_X1 U2910 ( .A1(n2667), .A2(n2666), .A3(n2665), .A4(n2664), .ZN(n3753)
         );
  INV_X1 U2911 ( .A(n3904), .ZN(n3872) );
  OR2_X1 U2912 ( .A1(n4280), .A2(n4256), .ZN(n4399) );
  INV_X1 U2913 ( .A(n3808), .ZN(n3955) );
  OR2_X1 U2914 ( .A1(n4576), .A2(n2841), .ZN(n4193) );
  OR2_X1 U2915 ( .A1(n3175), .A2(n4251), .ZN(n2842) );
  OR2_X1 U2916 ( .A1(n4558), .A2(n2841), .ZN(n4251) );
  OR2_X1 U2917 ( .A1(n2844), .A2(n2835), .ZN(n4558) );
  INV_X1 U2918 ( .A(n4480), .ZN(n4479) );
  INV_X1 U2919 ( .A(n3624), .ZN(U4043) );
  INV_X1 U2920 ( .A(n2351), .ZN(n2269) );
  INV_X1 U2921 ( .A(n4255), .ZN(n2279) );
  NAND2_X1 U2922 ( .A1(n2331), .A2(REG1_REG_0__SCAN_IN), .ZN(n2283) );
  NAND2_X1 U2923 ( .A1(n2345), .A2(REG3_REG_0__SCAN_IN), .ZN(n2282) );
  NAND2_X1 U2924 ( .A1(n2346), .A2(REG2_REG_0__SCAN_IN), .ZN(n2281) );
  NAND3_X1 U2925 ( .A1(n2302), .A2(n2288), .A3(n2287), .ZN(n2704) );
  INV_X1 U2926 ( .A(n2292), .ZN(n2293) );
  NAND2_X1 U2927 ( .A1(n2296), .A2(IR_REG_31__SCAN_IN), .ZN(n2297) );
  MUX2_X1 U2928 ( .A(IR_REG_31__SCAN_IN), .B(n2297), .S(IR_REG_21__SCAN_IN), 
        .Z(n2298) );
  NAND2_X1 U2929 ( .A1(n2040), .A2(IR_REG_31__SCAN_IN), .ZN(n2299) );
  INV_X1 U2930 ( .A(n4258), .ZN(n2301) );
  INV_X1 U2931 ( .A(n4259), .ZN(n2300) );
  NAND2_X1 U2932 ( .A1(n3625), .A2(n3195), .ZN(n2308) );
  MUX2_X1 U2933 ( .A(IR_REG_0__SCAN_IN), .B(DATAI_0_), .S(n2352), .Z(n2837) );
  INV_X1 U2934 ( .A(n2951), .ZN(n2305) );
  INV_X2 U2935 ( .A(n2369), .ZN(n2671) );
  INV_X1 U2936 ( .A(IR_REG_0__SCAN_IN), .ZN(n4505) );
  NOR2_X1 U2937 ( .A1(n2849), .A2(n4505), .ZN(n2306) );
  AOI21_X1 U2938 ( .B1(n2837), .B2(n2671), .A(n2306), .ZN(n2307) );
  NAND2_X1 U2939 ( .A1(n2308), .A2(n2307), .ZN(n2902) );
  NAND2_X1 U2940 ( .A1(n3625), .A2(n2671), .ZN(n2312) );
  INV_X1 U2941 ( .A(REG1_REG_0__SCAN_IN), .ZN(n2309) );
  NAND2_X1 U2942 ( .A1(n2837), .A2(n3190), .ZN(n2315) );
  OAI21_X1 U2943 ( .B1(n2849), .B2(n2309), .A(n2315), .ZN(n2310) );
  INV_X1 U2944 ( .A(n2310), .ZN(n2311) );
  NAND2_X1 U2945 ( .A1(n2312), .A2(n2311), .ZN(n2903) );
  NAND2_X1 U2946 ( .A1(n2902), .A2(n2903), .ZN(n2317) );
  NAND2_X1 U2947 ( .A1(n4258), .A2(n3681), .ZN(n2714) );
  NAND2_X1 U2948 ( .A1(n2315), .A2(n3193), .ZN(n2316) );
  NAND2_X1 U2949 ( .A1(n2345), .A2(REG3_REG_1__SCAN_IN), .ZN(n2320) );
  NAND2_X1 U2950 ( .A1(n2346), .A2(REG2_REG_1__SCAN_IN), .ZN(n2319) );
  NAND2_X1 U2951 ( .A1(n2331), .A2(REG1_REG_1__SCAN_IN), .ZN(n2318) );
  NAND2_X1 U2952 ( .A1(n2748), .A2(n2671), .ZN(n2323) );
  NAND2_X1 U2953 ( .A1(n2323), .A2(n2322), .ZN(n2324) );
  XNOR2_X1 U2954 ( .A(n2324), .B(n2687), .ZN(n2326) );
  NAND2_X1 U2955 ( .A1(n4439), .A2(n2671), .ZN(n2325) );
  NAND2_X1 U2956 ( .A1(n2262), .A2(n2325), .ZN(n2327) );
  INV_X1 U2957 ( .A(n2326), .ZN(n2329) );
  INV_X1 U2958 ( .A(n2327), .ZN(n2328) );
  NAND2_X1 U2959 ( .A1(n2964), .A2(n2671), .ZN(n2338) );
  NAND2_X1 U2960 ( .A1(n2331), .A2(REG1_REG_2__SCAN_IN), .ZN(n2336) );
  NAND2_X1 U2961 ( .A1(n2332), .A2(REG0_REG_2__SCAN_IN), .ZN(n2335) );
  NAND2_X1 U2962 ( .A1(n2345), .A2(REG3_REG_2__SCAN_IN), .ZN(n2334) );
  NAND2_X1 U2963 ( .A1(n2346), .A2(REG2_REG_2__SCAN_IN), .ZN(n2333) );
  OAI22_X1 U2964 ( .A1(n2753), .A2(n2029), .B1(n2339), .B2(n2970), .ZN(n2340)
         );
  XNOR2_X1 U2965 ( .A(n2340), .B(n3193), .ZN(n2341) );
  NAND2_X1 U2966 ( .A1(n2341), .A2(n2342), .ZN(n2343) );
  INV_X1 U2967 ( .A(n2343), .ZN(n2344) );
  NAND2_X1 U2968 ( .A1(n2331), .A2(REG1_REG_3__SCAN_IN), .ZN(n2349) );
  INV_X1 U2969 ( .A(REG3_REG_3__SCAN_IN), .ZN(n3249) );
  NAND2_X1 U2970 ( .A1(n2345), .A2(n3249), .ZN(n2348) );
  NAND2_X1 U2971 ( .A1(n2346), .A2(REG2_REG_3__SCAN_IN), .ZN(n2347) );
  NAND2_X1 U2972 ( .A1(n3623), .A2(n2671), .ZN(n2354) );
  NAND2_X1 U2973 ( .A1(n2351), .A2(IR_REG_31__SCAN_IN), .ZN(n2364) );
  XNOR2_X1 U2974 ( .A(n2364), .B(IR_REG_3__SCAN_IN), .ZN(n4266) );
  MUX2_X1 U2975 ( .A(n4266), .B(DATAI_3_), .S(n2352), .Z(n3474) );
  NAND2_X1 U2976 ( .A1(n3474), .A2(n3190), .ZN(n2353) );
  NAND2_X1 U2977 ( .A1(n2354), .A2(n2353), .ZN(n2355) );
  XNOR2_X1 U2978 ( .A(n2355), .B(n2687), .ZN(n2357) );
  INV_X1 U2979 ( .A(n3623), .ZN(n3473) );
  INV_X1 U2980 ( .A(n3474), .ZN(n2953) );
  OAI22_X1 U2981 ( .A1(n3473), .A2(n2657), .B1(n2029), .B2(n2953), .ZN(n2356)
         );
  XNOR2_X1 U2982 ( .A(n2357), .B(n2356), .ZN(n3245) );
  NOR2_X1 U2983 ( .A1(n2357), .A2(n2356), .ZN(n3345) );
  NAND2_X1 U2984 ( .A1(n2398), .A2(REG0_REG_4__SCAN_IN), .ZN(n2362) );
  NAND2_X1 U2985 ( .A1(n3514), .A2(REG1_REG_4__SCAN_IN), .ZN(n2361) );
  INV_X1 U2986 ( .A(REG3_REG_4__SCAN_IN), .ZN(n2358) );
  XNOR2_X1 U2987 ( .A(n2358), .B(REG3_REG_3__SCAN_IN), .ZN(n3350) );
  NAND2_X1 U2988 ( .A1(n2345), .A2(n3350), .ZN(n2360) );
  NAND2_X1 U2989 ( .A1(n3518), .A2(REG2_REG_4__SCAN_IN), .ZN(n2359) );
  OR2_X1 U2990 ( .A1(n2937), .A2(n2657), .ZN(n2368) );
  NAND2_X1 U2991 ( .A1(n2364), .A2(n2363), .ZN(n2365) );
  NAND2_X1 U2992 ( .A1(n2365), .A2(IR_REG_31__SCAN_IN), .ZN(n2366) );
  XNOR2_X1 U2993 ( .A(n2366), .B(IR_REG_4__SCAN_IN), .ZN(n4265) );
  MUX2_X1 U2994 ( .A(n4265), .B(DATAI_4_), .S(n2352), .Z(n3349) );
  NAND2_X1 U2995 ( .A1(n3349), .A2(n2671), .ZN(n2367) );
  NAND2_X1 U2996 ( .A1(n2368), .A2(n2367), .ZN(n2371) );
  INV_X1 U2997 ( .A(n3349), .ZN(n3000) );
  XNOR2_X1 U2998 ( .A(n2370), .B(n2687), .ZN(n2372) );
  XNOR2_X1 U2999 ( .A(n2371), .B(n2372), .ZN(n3344) );
  NOR2_X2 U3000 ( .A1(n3343), .A2(n2041), .ZN(n3314) );
  NAND2_X1 U3001 ( .A1(n3514), .A2(REG1_REG_5__SCAN_IN), .ZN(n2377) );
  NAND2_X1 U3002 ( .A1(n2398), .A2(REG0_REG_5__SCAN_IN), .ZN(n2376) );
  AOI21_X1 U3003 ( .B1(REG3_REG_3__SCAN_IN), .B2(REG3_REG_4__SCAN_IN), .A(
        REG3_REG_5__SCAN_IN), .ZN(n2373) );
  NOR2_X1 U3004 ( .A1(n2373), .A2(n2384), .ZN(n3318) );
  NAND2_X1 U3005 ( .A1(n2345), .A2(n3318), .ZN(n2375) );
  NAND2_X1 U3006 ( .A1(n3518), .A2(REG2_REG_5__SCAN_IN), .ZN(n2374) );
  NAND4_X1 U3007 ( .A1(n2377), .A2(n2376), .A3(n2375), .A4(n2374), .ZN(n3621)
         );
  INV_X1 U3008 ( .A(n3621), .ZN(n2797) );
  NAND2_X1 U3009 ( .A1(n2378), .A2(IR_REG_31__SCAN_IN), .ZN(n2379) );
  XNOR2_X1 U3010 ( .A(n2379), .B(IR_REG_5__SCAN_IN), .ZN(n4502) );
  MUX2_X1 U3011 ( .A(n4502), .B(DATAI_5_), .S(n2352), .Z(n3317) );
  INV_X1 U3012 ( .A(n3317), .ZN(n2981) );
  OAI22_X1 U3013 ( .A1(n2797), .A2(n2029), .B1(n2339), .B2(n2981), .ZN(n2380)
         );
  XNOR2_X1 U3014 ( .A(n2380), .B(n2687), .ZN(n2381) );
  AOI22_X1 U3015 ( .A1(n3621), .A2(n3195), .B1(n2671), .B2(n3317), .ZN(n2383)
         );
  XOR2_X1 U3016 ( .A(n2381), .B(n2383), .Z(n3315) );
  INV_X1 U3017 ( .A(n2381), .ZN(n2382) );
  OAI22_X1 U3018 ( .A1(n3314), .A2(n3315), .B1(n2383), .B2(n2382), .ZN(n3418)
         );
  NAND2_X1 U3019 ( .A1(n2398), .A2(REG0_REG_6__SCAN_IN), .ZN(n2388) );
  NAND2_X1 U3020 ( .A1(n3514), .A2(REG1_REG_6__SCAN_IN), .ZN(n2387) );
  NAND2_X1 U3021 ( .A1(n2384), .A2(REG3_REG_6__SCAN_IN), .ZN(n2399) );
  OAI21_X1 U3022 ( .B1(n2384), .B2(REG3_REG_6__SCAN_IN), .A(n2399), .ZN(n3017)
         );
  INV_X1 U3023 ( .A(n3017), .ZN(n3426) );
  NAND2_X1 U3024 ( .A1(n2345), .A2(n3426), .ZN(n2386) );
  NAND2_X1 U3025 ( .A1(n3518), .A2(REG2_REG_6__SCAN_IN), .ZN(n2385) );
  NAND4_X1 U3026 ( .A1(n2388), .A2(n2387), .A3(n2386), .A4(n2385), .ZN(n3620)
         );
  NAND2_X1 U3027 ( .A1(n3620), .A2(n2671), .ZN(n2394) );
  NOR2_X1 U3028 ( .A1(n2389), .A2(n2718), .ZN(n2390) );
  MUX2_X1 U3029 ( .A(n2718), .B(n2390), .S(IR_REG_6__SCAN_IN), .Z(n2392) );
  OR2_X1 U3030 ( .A1(n2392), .A2(n2391), .ZN(n4501) );
  INV_X1 U3031 ( .A(n4501), .ZN(n2884) );
  MUX2_X1 U3032 ( .A(n2884), .B(DATAI_6_), .S(n2352), .Z(n3425) );
  NAND2_X1 U3033 ( .A1(n3425), .A2(n3190), .ZN(n2393) );
  NAND2_X1 U3034 ( .A1(n2394), .A2(n2393), .ZN(n2395) );
  XNOR2_X1 U3035 ( .A(n2395), .B(n3193), .ZN(n2397) );
  AOI22_X1 U3036 ( .A1(n3620), .A2(n3195), .B1(n2671), .B2(n3425), .ZN(n2396)
         );
  NOR2_X1 U3037 ( .A1(n2397), .A2(n2396), .ZN(n3419) );
  NAND2_X1 U3038 ( .A1(n2397), .A2(n2396), .ZN(n3420) );
  NAND2_X1 U3039 ( .A1(n2398), .A2(REG0_REG_7__SCAN_IN), .ZN(n2404) );
  NAND2_X1 U3040 ( .A1(n3514), .A2(REG1_REG_7__SCAN_IN), .ZN(n2403) );
  NOR2_X1 U3041 ( .A1(n2399), .A2(n4039), .ZN(n2415) );
  AND2_X1 U3042 ( .A1(n2399), .A2(n4039), .ZN(n2400) );
  NOR2_X1 U3043 ( .A1(n2415), .A2(n2400), .ZN(n3064) );
  NAND2_X1 U3044 ( .A1(n2345), .A2(n3064), .ZN(n2402) );
  NAND2_X1 U3045 ( .A1(n3518), .A2(REG2_REG_7__SCAN_IN), .ZN(n2401) );
  OR2_X1 U3046 ( .A1(n3011), .A2(n2657), .ZN(n2410) );
  NOR2_X1 U3047 ( .A1(n2391), .A2(n2718), .ZN(n2405) );
  NAND2_X1 U3048 ( .A1(n2405), .A2(IR_REG_7__SCAN_IN), .ZN(n2408) );
  INV_X1 U3049 ( .A(n2405), .ZN(n2407) );
  INV_X1 U3050 ( .A(IR_REG_7__SCAN_IN), .ZN(n2406) );
  NAND2_X1 U3051 ( .A1(n2407), .A2(n2406), .ZN(n2421) );
  MUX2_X1 U3052 ( .A(n4264), .B(DATAI_7_), .S(n2352), .Z(n3055) );
  NAND2_X1 U3053 ( .A1(n3055), .A2(n2671), .ZN(n2409) );
  NAND2_X1 U3054 ( .A1(n2410), .A2(n2409), .ZN(n2413) );
  OAI22_X1 U3055 ( .A1(n3011), .A2(n2029), .B1(n2339), .B2(n3030), .ZN(n2411)
         );
  XNOR2_X1 U3056 ( .A(n2411), .B(n2687), .ZN(n2412) );
  XNOR2_X1 U3057 ( .A(n2413), .B(n2412), .ZN(n3061) );
  NAND2_X1 U3058 ( .A1(n3514), .A2(REG1_REG_8__SCAN_IN), .ZN(n2420) );
  NAND2_X1 U3059 ( .A1(n2398), .A2(REG0_REG_8__SCAN_IN), .ZN(n2419) );
  NAND2_X1 U3060 ( .A1(n2415), .A2(REG3_REG_8__SCAN_IN), .ZN(n2424) );
  OR2_X1 U3061 ( .A1(n2415), .A2(REG3_REG_8__SCAN_IN), .ZN(n2416) );
  AND2_X1 U3062 ( .A1(n2424), .A2(n2416), .ZN(n4429) );
  NAND2_X1 U3063 ( .A1(n2345), .A2(n4429), .ZN(n2418) );
  NAND2_X1 U3064 ( .A1(n3518), .A2(REG2_REG_8__SCAN_IN), .ZN(n2417) );
  NAND4_X1 U3065 ( .A1(n2420), .A2(n2419), .A3(n2418), .A4(n2417), .ZN(n3618)
         );
  NAND2_X1 U3066 ( .A1(n2421), .A2(IR_REG_31__SCAN_IN), .ZN(n2422) );
  XNOR2_X1 U3067 ( .A(n2422), .B(IR_REG_8__SCAN_IN), .ZN(n4263) );
  MUX2_X1 U3068 ( .A(n4263), .B(DATAI_8_), .S(n2352), .Z(n3269) );
  OAI22_X1 U3069 ( .A1(n3120), .A2(n2657), .B1(n2029), .B2(n3103), .ZN(n3264)
         );
  OAI22_X1 U3070 ( .A1(n3120), .A2(n2029), .B1(n2339), .B2(n3103), .ZN(n2423)
         );
  XNOR2_X1 U3071 ( .A(n2423), .B(n2687), .ZN(n3265) );
  NAND2_X1 U3072 ( .A1(n2398), .A2(REG0_REG_9__SCAN_IN), .ZN(n2429) );
  NAND2_X1 U3073 ( .A1(n3514), .A2(REG1_REG_9__SCAN_IN), .ZN(n2428) );
  NAND2_X1 U3074 ( .A1(n2424), .A2(n3119), .ZN(n2425) );
  AND2_X1 U3075 ( .A1(n2434), .A2(n2425), .ZN(n3123) );
  NAND2_X1 U3076 ( .A1(n2345), .A2(n3123), .ZN(n2427) );
  NAND2_X1 U3077 ( .A1(n3518), .A2(REG2_REG_9__SCAN_IN), .ZN(n2426) );
  NAND4_X1 U3078 ( .A1(n2429), .A2(n2428), .A3(n2427), .A4(n2426), .ZN(n3617)
         );
  INV_X1 U3079 ( .A(n3617), .ZN(n3104) );
  NAND2_X1 U3080 ( .A1(n2430), .A2(IR_REG_31__SCAN_IN), .ZN(n2431) );
  MUX2_X1 U3081 ( .A(IR_REG_31__SCAN_IN), .B(n2431), .S(IR_REG_9__SCAN_IN), 
        .Z(n2432) );
  MUX2_X1 U3082 ( .A(n3081), .B(DATAI_9_), .S(n2352), .Z(n3050) );
  INV_X1 U3083 ( .A(n3050), .ZN(n3121) );
  OAI22_X1 U3084 ( .A1(n3104), .A2(n2029), .B1(n2339), .B2(n3121), .ZN(n2433)
         );
  XNOR2_X1 U3085 ( .A(n2433), .B(n2687), .ZN(n2443) );
  OAI22_X1 U3086 ( .A1(n3104), .A2(n2657), .B1(n2029), .B2(n3121), .ZN(n2442)
         );
  XNOR2_X1 U3087 ( .A(n2443), .B(n2442), .ZN(n3118) );
  NAND2_X1 U3088 ( .A1(n3514), .A2(REG1_REG_10__SCAN_IN), .ZN(n2439) );
  NAND2_X1 U3089 ( .A1(n2398), .A2(REG0_REG_10__SCAN_IN), .ZN(n2438) );
  NAND2_X1 U3090 ( .A1(n2434), .A2(n4059), .ZN(n2435) );
  AND2_X1 U3091 ( .A1(n2449), .A2(n2435), .ZN(n4422) );
  NAND2_X1 U3092 ( .A1(n2345), .A2(n4422), .ZN(n2437) );
  NAND2_X1 U3093 ( .A1(n3518), .A2(REG2_REG_10__SCAN_IN), .ZN(n2436) );
  NAND4_X1 U3094 ( .A1(n2439), .A2(n2438), .A3(n2437), .A4(n2436), .ZN(n4406)
         );
  NAND2_X1 U3095 ( .A1(n2488), .A2(IR_REG_31__SCAN_IN), .ZN(n2440) );
  XNOR2_X1 U3096 ( .A(n2440), .B(IR_REG_10__SCAN_IN), .ZN(n3088) );
  MUX2_X1 U3097 ( .A(n3088), .B(DATAI_10_), .S(n2352), .Z(n3240) );
  AOI22_X1 U3098 ( .A1(n4406), .A2(n3195), .B1(n2671), .B2(n3240), .ZN(n2445)
         );
  INV_X1 U3099 ( .A(n4406), .ZN(n2802) );
  OAI22_X1 U3100 ( .A1(n2802), .A2(n2029), .B1(n2339), .B2(n3143), .ZN(n2441)
         );
  XNOR2_X1 U3101 ( .A(n2441), .B(n2687), .ZN(n2444) );
  XOR2_X1 U3102 ( .A(n2445), .B(n2444), .Z(n3235) );
  NOR2_X1 U3103 ( .A1(n2443), .A2(n2442), .ZN(n3236) );
  NAND2_X1 U3104 ( .A1(n3115), .A2(n2045), .ZN(n3237) );
  INV_X1 U3105 ( .A(n2444), .ZN(n2446) );
  OR2_X1 U3106 ( .A1(n2446), .A2(n2445), .ZN(n2447) );
  NAND2_X1 U3107 ( .A1(n3514), .A2(REG1_REG_11__SCAN_IN), .ZN(n2454) );
  NAND2_X1 U3108 ( .A1(n2398), .A2(REG0_REG_11__SCAN_IN), .ZN(n2453) );
  AND2_X1 U3109 ( .A1(n2449), .A2(n2448), .ZN(n2450) );
  OR2_X1 U3110 ( .A1(n2450), .A2(n2463), .ZN(n4414) );
  INV_X1 U3111 ( .A(n4414), .ZN(n3403) );
  NAND2_X1 U3112 ( .A1(n2345), .A2(n3403), .ZN(n2452) );
  NAND2_X1 U3113 ( .A1(n3518), .A2(REG2_REG_11__SCAN_IN), .ZN(n2451) );
  OR2_X1 U3114 ( .A1(n3144), .A2(n2657), .ZN(n2457) );
  NAND2_X1 U3115 ( .A1(n2455), .A2(IR_REG_31__SCAN_IN), .ZN(n2470) );
  XNOR2_X1 U3116 ( .A(n2470), .B(IR_REG_11__SCAN_IN), .ZN(n4494) );
  MUX2_X1 U3117 ( .A(n4494), .B(DATAI_11_), .S(n2352), .Z(n3402) );
  NAND2_X1 U3118 ( .A1(n3402), .A2(n2671), .ZN(n2456) );
  AND2_X1 U3119 ( .A1(n2457), .A2(n2456), .ZN(n2460) );
  OAI22_X1 U3120 ( .A1(n3144), .A2(n2029), .B1(n2339), .B2(n4417), .ZN(n2458)
         );
  XNOR2_X1 U3121 ( .A(n2458), .B(n3193), .ZN(n2459) );
  NAND2_X1 U3122 ( .A1(n2460), .A2(n2459), .ZN(n3398) );
  INV_X1 U3123 ( .A(n2459), .ZN(n2462) );
  INV_X1 U3124 ( .A(n2460), .ZN(n2461) );
  NAND2_X1 U3125 ( .A1(n2462), .A2(n2461), .ZN(n3397) );
  NAND2_X1 U3126 ( .A1(n2398), .A2(REG0_REG_12__SCAN_IN), .ZN(n2468) );
  NAND2_X1 U3127 ( .A1(n3514), .A2(REG1_REG_12__SCAN_IN), .ZN(n2467) );
  OR2_X1 U3128 ( .A1(n2463), .A2(REG3_REG_12__SCAN_IN), .ZN(n2464) );
  NAND2_X1 U3129 ( .A1(n2463), .A2(REG3_REG_12__SCAN_IN), .ZN(n2479) );
  AND2_X1 U3130 ( .A1(n2464), .A2(n2479), .ZN(n3287) );
  NAND2_X1 U3131 ( .A1(n2345), .A2(n3287), .ZN(n2466) );
  NAND2_X1 U3132 ( .A1(n3518), .A2(REG2_REG_12__SCAN_IN), .ZN(n2465) );
  NAND4_X1 U3133 ( .A1(n2468), .A2(n2467), .A3(n2466), .A4(n2465), .ZN(n3401)
         );
  NAND2_X1 U3134 ( .A1(n3401), .A2(n3195), .ZN(n2474) );
  INV_X1 U3135 ( .A(IR_REG_11__SCAN_IN), .ZN(n2469) );
  NAND2_X1 U3136 ( .A1(n2470), .A2(n2469), .ZN(n2471) );
  NAND2_X1 U3137 ( .A1(n2471), .A2(IR_REG_31__SCAN_IN), .ZN(n2472) );
  XNOR2_X1 U3138 ( .A(n2472), .B(IR_REG_12__SCAN_IN), .ZN(n3091) );
  MUX2_X1 U3139 ( .A(n3091), .B(DATAI_12_), .S(n2352), .Z(n3286) );
  NAND2_X1 U3140 ( .A1(n3286), .A2(n2671), .ZN(n2473) );
  NAND2_X1 U3141 ( .A1(n2474), .A2(n2473), .ZN(n3369) );
  INV_X1 U3142 ( .A(n3369), .ZN(n2494) );
  NAND2_X1 U3143 ( .A1(n3401), .A2(n2671), .ZN(n2476) );
  NAND2_X1 U3144 ( .A1(n3286), .A2(n3190), .ZN(n2475) );
  NAND2_X1 U3145 ( .A1(n2476), .A2(n2475), .ZN(n2477) );
  XNOR2_X1 U3146 ( .A(n2477), .B(n2687), .ZN(n3370) );
  INV_X1 U3147 ( .A(n3370), .ZN(n3372) );
  NAND2_X1 U31480 ( .A1(n3514), .A2(REG1_REG_13__SCAN_IN), .ZN(n2484) );
  NAND2_X1 U31490 ( .A1(n2398), .A2(REG0_REG_13__SCAN_IN), .ZN(n2483) );
  NAND2_X1 U3150 ( .A1(n2479), .A2(n2478), .ZN(n2480) );
  AND2_X1 U3151 ( .A1(n2501), .A2(n2480), .ZN(n3378) );
  NAND2_X1 U3152 ( .A1(n2345), .A2(n3378), .ZN(n2482) );
  NAND2_X1 U3153 ( .A1(n3518), .A2(REG2_REG_13__SCAN_IN), .ZN(n2481) );
  NAND4_X1 U3154 ( .A1(n2484), .A2(n2483), .A3(n2482), .A4(n2481), .ZN(n3615)
         );
  NAND2_X1 U3155 ( .A1(n3615), .A2(n2671), .ZN(n2491) );
  INV_X1 U3156 ( .A(IR_REG_12__SCAN_IN), .ZN(n2485) );
  NAND2_X1 U3157 ( .A1(n2486), .A2(n2485), .ZN(n2487) );
  NAND2_X1 U3158 ( .A1(n2507), .A2(IR_REG_31__SCAN_IN), .ZN(n2489) );
  XNOR2_X1 U3159 ( .A(n2489), .B(IR_REG_13__SCAN_IN), .ZN(n4491) );
  MUX2_X1 U3160 ( .A(n4491), .B(DATAI_13_), .S(n2352), .Z(n3377) );
  NAND2_X1 U3161 ( .A1(n3377), .A2(n3190), .ZN(n2490) );
  NAND2_X1 U3162 ( .A1(n2491), .A2(n2490), .ZN(n2492) );
  XNOR2_X1 U3163 ( .A(n2492), .B(n3193), .ZN(n2496) );
  AOI22_X1 U3164 ( .A1(n3615), .A2(n3195), .B1(n2671), .B2(n3377), .ZN(n2495)
         );
  NOR2_X1 U3165 ( .A1(n2496), .A2(n2495), .ZN(n3368) );
  INV_X1 U3166 ( .A(n3368), .ZN(n2493) );
  OAI21_X1 U3167 ( .B1(n2494), .B2(n3372), .A(n2493), .ZN(n2499) );
  NOR3_X1 U3168 ( .A1(n3368), .A2(n3369), .A3(n3370), .ZN(n2497) );
  AND2_X1 U3169 ( .A1(n2496), .A2(n2495), .ZN(n3367) );
  NOR2_X1 U3170 ( .A1(n2497), .A2(n3367), .ZN(n2498) );
  NAND2_X1 U3171 ( .A1(n3514), .A2(REG1_REG_14__SCAN_IN), .ZN(n2506) );
  NAND2_X1 U3172 ( .A1(n2398), .A2(REG0_REG_14__SCAN_IN), .ZN(n2505) );
  AND2_X1 U3173 ( .A1(n2501), .A2(n2500), .ZN(n2502) );
  NOR2_X1 U3174 ( .A1(n2514), .A2(n2502), .ZN(n3970) );
  NAND2_X1 U3175 ( .A1(n2345), .A2(n3970), .ZN(n2504) );
  NAND2_X1 U3176 ( .A1(n3518), .A2(REG2_REG_14__SCAN_IN), .ZN(n2503) );
  NOR2_X1 U3177 ( .A1(n2507), .A2(IR_REG_13__SCAN_IN), .ZN(n2521) );
  OR2_X1 U3178 ( .A1(n2521), .A2(n2718), .ZN(n2508) );
  XNOR2_X1 U3179 ( .A(n2508), .B(IR_REG_14__SCAN_IN), .ZN(n4262) );
  MUX2_X1 U3180 ( .A(n4262), .B(DATAI_14_), .S(n2352), .Z(n3969) );
  OAI22_X1 U3181 ( .A1(n2771), .A2(n2029), .B1(n2339), .B2(n2838), .ZN(n2509)
         );
  XOR2_X1 U3182 ( .A(n2687), .B(n2509), .Z(n3217) );
  NAND2_X1 U3183 ( .A1(n2510), .A2(n3216), .ZN(n2513) );
  NAND2_X1 U3184 ( .A1(n2511), .A2(n2223), .ZN(n2512) );
  NAND2_X1 U3185 ( .A1(n2513), .A2(n2512), .ZN(n2531) );
  INV_X1 U3186 ( .A(n2531), .ZN(n2528) );
  NAND2_X1 U3187 ( .A1(n2398), .A2(REG0_REG_15__SCAN_IN), .ZN(n2519) );
  NAND2_X1 U3188 ( .A1(n3514), .A2(REG1_REG_15__SCAN_IN), .ZN(n2518) );
  NOR2_X1 U3189 ( .A1(n2514), .A2(REG3_REG_15__SCAN_IN), .ZN(n2515) );
  NOR2_X1 U3190 ( .A1(n2532), .A2(n2515), .ZN(n3950) );
  NAND2_X1 U3191 ( .A1(n2345), .A2(n3950), .ZN(n2517) );
  NAND2_X1 U3192 ( .A1(n3518), .A2(REG2_REG_15__SCAN_IN), .ZN(n2516) );
  NAND4_X1 U3193 ( .A1(n2519), .A2(n2518), .A3(n2517), .A4(n2516), .ZN(n3963)
         );
  INV_X1 U3194 ( .A(n3963), .ZN(n2805) );
  INV_X1 U3195 ( .A(IR_REG_14__SCAN_IN), .ZN(n2520) );
  NAND2_X1 U3196 ( .A1(n2521), .A2(n2520), .ZN(n2522) );
  NAND2_X1 U3197 ( .A1(n2522), .A2(IR_REG_31__SCAN_IN), .ZN(n2524) );
  NAND2_X1 U3198 ( .A1(n2524), .A2(n2523), .ZN(n2538) );
  OR2_X1 U3199 ( .A1(n2524), .A2(n2523), .ZN(n2525) );
  MUX2_X1 U3200 ( .A(n3671), .B(DATAI_15_), .S(n2352), .Z(n3447) );
  OAI22_X1 U3201 ( .A1(n2805), .A2(n2029), .B1(n2339), .B2(n3947), .ZN(n2526)
         );
  NAND2_X1 U3202 ( .A1(n2528), .A2(n2527), .ZN(n3304) );
  NAND2_X1 U3203 ( .A1(n3963), .A2(n3195), .ZN(n2530) );
  NAND2_X1 U3204 ( .A1(n3447), .A2(n2671), .ZN(n2529) );
  NAND2_X1 U3205 ( .A1(n2530), .A2(n2529), .ZN(n3443) );
  NAND2_X1 U3206 ( .A1(n2531), .A2(n2054), .ZN(n3442) );
  NAND2_X1 U3207 ( .A1(n2332), .A2(REG0_REG_16__SCAN_IN), .ZN(n2537) );
  NAND2_X1 U3208 ( .A1(n3514), .A2(REG1_REG_16__SCAN_IN), .ZN(n2536) );
  OR2_X1 U3209 ( .A1(n2532), .A2(REG3_REG_16__SCAN_IN), .ZN(n2533) );
  NAND2_X1 U32100 ( .A1(n2532), .A2(REG3_REG_16__SCAN_IN), .ZN(n2547) );
  AND2_X1 U32110 ( .A1(n2533), .A2(n2547), .ZN(n3930) );
  NAND2_X1 U32120 ( .A1(n2345), .A2(n3930), .ZN(n2535) );
  NAND2_X1 U32130 ( .A1(n3518), .A2(REG2_REG_16__SCAN_IN), .ZN(n2534) );
  NAND2_X1 U32140 ( .A1(n2538), .A2(IR_REG_31__SCAN_IN), .ZN(n2539) );
  XNOR2_X1 U32150 ( .A(n2539), .B(IR_REG_16__SCAN_IN), .ZN(n3672) );
  MUX2_X1 U32160 ( .A(n3672), .B(DATAI_16_), .S(n2352), .Z(n3309) );
  INV_X1 U32170 ( .A(n3309), .ZN(n3928) );
  OAI22_X1 U32180 ( .A1(n3942), .A2(n2029), .B1(n2339), .B2(n3928), .ZN(n2540)
         );
  XNOR2_X1 U32190 ( .A(n2540), .B(n2687), .ZN(n2541) );
  AOI22_X1 U32200 ( .A1(n3906), .A2(n3195), .B1(n2671), .B2(n3309), .ZN(n2542)
         );
  XNOR2_X1 U32210 ( .A(n2541), .B(n2542), .ZN(n3306) );
  NAND2_X1 U32220 ( .A1(n3442), .A2(n3306), .ZN(n2545) );
  NAND2_X1 U32230 ( .A1(n3514), .A2(REG1_REG_17__SCAN_IN), .ZN(n2553) );
  NAND2_X1 U32240 ( .A1(n2398), .A2(REG0_REG_17__SCAN_IN), .ZN(n2552) );
  NOR2_X1 U32250 ( .A1(REG3_REG_17__SCAN_IN), .A2(n2548), .ZN(n2549) );
  NOR2_X1 U32260 ( .A1(n2561), .A2(n2549), .ZN(n3913) );
  NAND2_X1 U32270 ( .A1(n2345), .A2(n3913), .ZN(n2551) );
  NAND2_X1 U32280 ( .A1(n3518), .A2(REG2_REG_17__SCAN_IN), .ZN(n2550) );
  NAND2_X1 U32290 ( .A1(n2065), .A2(IR_REG_31__SCAN_IN), .ZN(n2554) );
  XNOR2_X1 U32300 ( .A(n2554), .B(IR_REG_17__SCAN_IN), .ZN(n4485) );
  MUX2_X1 U32310 ( .A(n4485), .B(DATAI_17_), .S(n2352), .Z(n3328) );
  INV_X1 U32320 ( .A(n3328), .ZN(n3911) );
  OAI22_X1 U32330 ( .A1(n3923), .A2(n2029), .B1(n2339), .B2(n3911), .ZN(n2555)
         );
  XNOR2_X1 U32340 ( .A(n2555), .B(n2687), .ZN(n3325) );
  OR2_X1 U32350 ( .A1(n3923), .A2(n2657), .ZN(n2557) );
  NAND2_X1 U32360 ( .A1(n3328), .A2(n2671), .ZN(n2556) );
  NAND2_X1 U32370 ( .A1(n2557), .A2(n2556), .ZN(n2558) );
  NOR2_X1 U32380 ( .A1(n3325), .A2(n2558), .ZN(n2560) );
  INV_X1 U32390 ( .A(n3325), .ZN(n2559) );
  INV_X1 U32400 ( .A(n2558), .ZN(n3324) );
  NAND2_X1 U32410 ( .A1(n3514), .A2(REG1_REG_18__SCAN_IN), .ZN(n2566) );
  NAND2_X1 U32420 ( .A1(n2398), .A2(REG0_REG_18__SCAN_IN), .ZN(n2565) );
  NOR2_X1 U32430 ( .A1(n2561), .A2(REG3_REG_18__SCAN_IN), .ZN(n2562) );
  NOR2_X1 U32440 ( .A1(n2573), .A2(n2562), .ZN(n3895) );
  NAND2_X1 U32450 ( .A1(n2345), .A2(n3895), .ZN(n2564) );
  NAND2_X1 U32460 ( .A1(n3518), .A2(REG2_REG_18__SCAN_IN), .ZN(n2563) );
  OR2_X1 U32470 ( .A1(n2292), .A2(n2718), .ZN(n2567) );
  XNOR2_X1 U32480 ( .A(n2567), .B(IR_REG_18__SCAN_IN), .ZN(n3675) );
  MUX2_X1 U32490 ( .A(n3675), .B(DATAI_18_), .S(n2352), .Z(n3886) );
  OAI22_X1 U32500 ( .A1(n3904), .A2(n2029), .B1(n2339), .B2(n3891), .ZN(n2568)
         );
  XNOR2_X1 U32510 ( .A(n2568), .B(n3193), .ZN(n2572) );
  OR2_X1 U32520 ( .A1(n3904), .A2(n2657), .ZN(n2570) );
  NAND2_X1 U32530 ( .A1(n3886), .A2(n2671), .ZN(n2569) );
  AND2_X1 U32540 ( .A1(n2570), .A2(n2569), .ZN(n2571) );
  NOR2_X1 U32550 ( .A1(n2572), .A2(n2571), .ZN(n3408) );
  NAND2_X1 U32560 ( .A1(n2572), .A2(n2571), .ZN(n3409) );
  NAND2_X1 U32570 ( .A1(n2332), .A2(REG0_REG_19__SCAN_IN), .ZN(n2578) );
  NAND2_X1 U32580 ( .A1(n3514), .A2(REG1_REG_19__SCAN_IN), .ZN(n2577) );
  NOR2_X1 U32590 ( .A1(n2573), .A2(REG3_REG_19__SCAN_IN), .ZN(n2574) );
  NOR2_X1 U32600 ( .A1(n2587), .A2(n2574), .ZN(n3877) );
  NAND2_X1 U32610 ( .A1(n2345), .A2(n3877), .ZN(n2576) );
  NAND2_X1 U32620 ( .A1(n3518), .A2(REG2_REG_19__SCAN_IN), .ZN(n2575) );
  NAND4_X1 U32630 ( .A1(n2578), .A2(n2577), .A3(n2576), .A4(n2575), .ZN(n3887)
         );
  INV_X1 U32640 ( .A(n3887), .ZN(n2777) );
  INV_X1 U32650 ( .A(DATAI_19_), .ZN(n2579) );
  MUX2_X1 U32660 ( .A(n3681), .B(n2579), .S(n2352), .Z(n3876) );
  OAI22_X1 U32670 ( .A1(n2777), .A2(n2657), .B1(n2029), .B2(n3876), .ZN(n2584)
         );
  NAND2_X1 U32680 ( .A1(n3887), .A2(n2671), .ZN(n2581) );
  INV_X1 U32690 ( .A(n3876), .ZN(n3258) );
  NAND2_X1 U32700 ( .A1(n3258), .A2(n3190), .ZN(n2580) );
  NAND2_X1 U32710 ( .A1(n2581), .A2(n2580), .ZN(n2582) );
  XNOR2_X1 U32720 ( .A(n2582), .B(n2687), .ZN(n2583) );
  XOR2_X1 U32730 ( .A(n2584), .B(n2583), .Z(n3254) );
  INV_X1 U32740 ( .A(n2584), .ZN(n2585) );
  NAND2_X1 U32750 ( .A1(n2398), .A2(REG0_REG_20__SCAN_IN), .ZN(n2592) );
  NAND2_X1 U32760 ( .A1(n3514), .A2(REG1_REG_20__SCAN_IN), .ZN(n2591) );
  OAI21_X1 U32770 ( .B1(n2587), .B2(REG3_REG_20__SCAN_IN), .A(n2614), .ZN(
        n2588) );
  INV_X1 U32780 ( .A(n2588), .ZN(n3856) );
  NAND2_X1 U32790 ( .A1(n2345), .A2(n3856), .ZN(n2590) );
  NAND2_X1 U32800 ( .A1(n3518), .A2(REG2_REG_20__SCAN_IN), .ZN(n2589) );
  NAND4_X1 U32810 ( .A1(n2592), .A2(n2591), .A3(n2590), .A4(n2589), .ZN(n3613)
         );
  NAND2_X1 U32820 ( .A1(n3613), .A2(n2671), .ZN(n2594) );
  NAND2_X1 U32830 ( .A1(n2352), .A2(DATAI_20_), .ZN(n3854) );
  NAND2_X1 U32840 ( .A1(n3190), .A2(n3362), .ZN(n2593) );
  NAND2_X1 U32850 ( .A1(n2594), .A2(n2593), .ZN(n2595) );
  XNOR2_X1 U32860 ( .A(n2595), .B(n2687), .ZN(n2598) );
  NAND2_X1 U32870 ( .A1(n3613), .A2(n3195), .ZN(n2597) );
  NAND2_X1 U32880 ( .A1(n2671), .A2(n3362), .ZN(n2596) );
  NAND2_X1 U32890 ( .A1(n2597), .A2(n2596), .ZN(n2599) );
  NAND2_X1 U32900 ( .A1(n2598), .A2(n2599), .ZN(n3358) );
  INV_X1 U32910 ( .A(n2598), .ZN(n2601) );
  INV_X1 U32920 ( .A(n2599), .ZN(n2600) );
  NAND2_X1 U32930 ( .A1(n2601), .A2(n2600), .ZN(n3359) );
  NAND2_X1 U32940 ( .A1(n2332), .A2(REG0_REG_21__SCAN_IN), .ZN(n2605) );
  NAND2_X1 U32950 ( .A1(n3514), .A2(REG1_REG_21__SCAN_IN), .ZN(n2604) );
  XNOR2_X1 U32960 ( .A(n2614), .B(REG3_REG_21__SCAN_IN), .ZN(n3837) );
  NAND2_X1 U32970 ( .A1(n2345), .A2(n3837), .ZN(n2603) );
  NAND2_X1 U32980 ( .A1(n3518), .A2(REG2_REG_21__SCAN_IN), .ZN(n2602) );
  OR2_X1 U32990 ( .A1(n3849), .A2(n2657), .ZN(n2607) );
  NAND2_X1 U33000 ( .A1(n2671), .A2(n3829), .ZN(n2606) );
  INV_X1 U33010 ( .A(n3829), .ZN(n3835) );
  OAI22_X1 U33020 ( .A1(n3849), .A2(n2029), .B1(n2339), .B2(n3835), .ZN(n2608)
         );
  XNOR2_X1 U33030 ( .A(n2608), .B(n3193), .ZN(n3275) );
  NAND2_X1 U33040 ( .A1(n3274), .A2(n3275), .ZN(n2609) );
  INV_X1 U33050 ( .A(n3275), .ZN(n2611) );
  INV_X1 U33060 ( .A(n3274), .ZN(n2610) );
  INV_X1 U33070 ( .A(n3383), .ZN(n2622) );
  NAND2_X1 U33080 ( .A1(n2398), .A2(REG0_REG_22__SCAN_IN), .ZN(n2619) );
  NAND2_X1 U33090 ( .A1(n3514), .A2(REG1_REG_22__SCAN_IN), .ZN(n2618) );
  INV_X1 U33100 ( .A(n2614), .ZN(n2612) );
  AOI21_X1 U33110 ( .B1(n2612), .B2(REG3_REG_21__SCAN_IN), .A(
        REG3_REG_22__SCAN_IN), .ZN(n2615) );
  NAND2_X1 U33120 ( .A1(REG3_REG_21__SCAN_IN), .A2(REG3_REG_22__SCAN_IN), .ZN(
        n2613) );
  OR2_X1 U33130 ( .A1(n2615), .A2(n2623), .ZN(n3809) );
  INV_X1 U33140 ( .A(n3809), .ZN(n3392) );
  NAND2_X1 U33150 ( .A1(n2345), .A2(n3392), .ZN(n2617) );
  NAND2_X1 U33160 ( .A1(n3518), .A2(REG2_REG_22__SCAN_IN), .ZN(n2616) );
  OAI22_X1 U33170 ( .A1(n3795), .A2(n2029), .B1(n2339), .B2(n3820), .ZN(n2620)
         );
  XNOR2_X1 U33180 ( .A(n2620), .B(n2687), .ZN(n2633) );
  OAI22_X1 U33190 ( .A1(n3795), .A2(n2657), .B1(n2029), .B2(n3820), .ZN(n2632)
         );
  XNOR2_X1 U33200 ( .A(n2633), .B(n2632), .ZN(n3385) );
  NAND2_X1 U33210 ( .A1(n3514), .A2(REG1_REG_23__SCAN_IN), .ZN(n2628) );
  NAND2_X1 U33220 ( .A1(n2332), .A2(REG0_REG_23__SCAN_IN), .ZN(n2627) );
  NAND2_X1 U33230 ( .A1(n2623), .A2(REG3_REG_23__SCAN_IN), .ZN(n2638) );
  OR2_X1 U33240 ( .A1(n2623), .A2(REG3_REG_23__SCAN_IN), .ZN(n2624) );
  AND2_X1 U33250 ( .A1(n2638), .A2(n2624), .ZN(n3799) );
  NAND2_X1 U33260 ( .A1(n2345), .A2(n3799), .ZN(n2626) );
  NAND2_X1 U33270 ( .A1(n3518), .A2(REG2_REG_23__SCAN_IN), .ZN(n2625) );
  INV_X1 U33280 ( .A(n3791), .ZN(n3798) );
  OAI22_X1 U33290 ( .A1(n3816), .A2(n2029), .B1(n2339), .B2(n3798), .ZN(n2629)
         );
  XNOR2_X1 U33300 ( .A(n2629), .B(n2687), .ZN(n2636) );
  OR2_X1 U33310 ( .A1(n3816), .A2(n2657), .ZN(n2631) );
  NAND2_X1 U33320 ( .A1(n2671), .A2(n3791), .ZN(n2630) );
  NAND2_X1 U33330 ( .A1(n2631), .A2(n2630), .ZN(n2635) );
  XNOR2_X1 U33340 ( .A(n2636), .B(n2635), .ZN(n3227) );
  NOR2_X1 U33350 ( .A1(n2633), .A2(n2632), .ZN(n3228) );
  NOR2_X1 U33360 ( .A1(n3227), .A2(n3228), .ZN(n2634) );
  NAND2_X1 U33370 ( .A1(n2636), .A2(n2635), .ZN(n2647) );
  NAND2_X1 U33380 ( .A1(n3514), .A2(REG1_REG_24__SCAN_IN), .ZN(n2643) );
  NAND2_X1 U33390 ( .A1(n2398), .A2(REG0_REG_24__SCAN_IN), .ZN(n2642) );
  INV_X1 U33400 ( .A(REG3_REG_24__SCAN_IN), .ZN(n2637) );
  NAND2_X1 U33410 ( .A1(n2638), .A2(n2637), .ZN(n2639) );
  AND2_X1 U33420 ( .A1(n2650), .A2(n2639), .ZN(n3776) );
  NAND2_X1 U33430 ( .A1(n2345), .A2(n3776), .ZN(n2641) );
  NAND2_X1 U33440 ( .A1(n3518), .A2(REG2_REG_24__SCAN_IN), .ZN(n2640) );
  NAND4_X1 U33450 ( .A1(n2643), .A2(n2642), .A3(n2641), .A4(n2640), .ZN(n3792)
         );
  NOR2_X1 U33460 ( .A1(n2029), .A2(n3774), .ZN(n2644) );
  AOI21_X1 U33470 ( .B1(n3792), .B2(n3195), .A(n2644), .ZN(n2648) );
  INV_X1 U33480 ( .A(n3792), .ZN(n3756) );
  OAI22_X1 U33490 ( .A1(n3756), .A2(n2029), .B1(n2339), .B2(n3774), .ZN(n2646)
         );
  XNOR2_X1 U33500 ( .A(n2646), .B(n2687), .ZN(n3335) );
  INV_X1 U33510 ( .A(n2648), .ZN(n2649) );
  NAND2_X1 U33520 ( .A1(n2398), .A2(REG0_REG_25__SCAN_IN), .ZN(n2655) );
  NAND2_X1 U3353 ( .A1(n3514), .A2(REG1_REG_25__SCAN_IN), .ZN(n2654) );
  INV_X1 U33540 ( .A(REG3_REG_25__SCAN_IN), .ZN(n3298) );
  NAND2_X1 U3355 ( .A1(n2650), .A2(n3298), .ZN(n2651) );
  NAND2_X1 U3356 ( .A1(n2345), .A2(n3760), .ZN(n2653) );
  NAND2_X1 U3357 ( .A1(n3518), .A2(REG2_REG_25__SCAN_IN), .ZN(n2652) );
  OAI22_X1 U3358 ( .A1(n3768), .A2(n2029), .B1(n2339), .B2(n2787), .ZN(n2656)
         );
  XNOR2_X1 U3359 ( .A(n2656), .B(n3193), .ZN(n2661) );
  OR2_X1 U3360 ( .A1(n3768), .A2(n2657), .ZN(n2659) );
  NAND2_X1 U3361 ( .A1(n2671), .A2(n3757), .ZN(n2658) );
  AND2_X1 U3362 ( .A1(n2659), .A2(n2658), .ZN(n2660) );
  NAND2_X1 U3363 ( .A1(n2661), .A2(n2660), .ZN(n3294) );
  NOR2_X1 U3364 ( .A1(n2661), .A2(n2660), .ZN(n3293) );
  AOI21_X1 U3365 ( .B1(n3292), .B2(n3294), .A(n3293), .ZN(n3431) );
  NAND2_X1 U3366 ( .A1(n3514), .A2(REG1_REG_26__SCAN_IN), .ZN(n2667) );
  NAND2_X1 U3367 ( .A1(n2398), .A2(REG0_REG_26__SCAN_IN), .ZN(n2666) );
  INV_X1 U3368 ( .A(REG3_REG_26__SCAN_IN), .ZN(n3436) );
  AND2_X1 U3369 ( .A1(n2662), .A2(n3436), .ZN(n2663) );
  NOR2_X1 U3370 ( .A1(n2679), .A2(n2663), .ZN(n3732) );
  NAND2_X1 U3371 ( .A1(n2345), .A2(n3732), .ZN(n2665) );
  NAND2_X1 U3372 ( .A1(n3518), .A2(REG2_REG_26__SCAN_IN), .ZN(n2664) );
  NAND2_X1 U3373 ( .A1(n3753), .A2(n2671), .ZN(n2669) );
  NAND2_X1 U3374 ( .A1(n3190), .A2(n3741), .ZN(n2668) );
  NAND2_X1 U3375 ( .A1(n2669), .A2(n2668), .ZN(n2670) );
  XNOR2_X1 U3376 ( .A(n2670), .B(n2687), .ZN(n2674) );
  NAND2_X1 U3377 ( .A1(n3753), .A2(n3195), .ZN(n2673) );
  NAND2_X1 U3378 ( .A1(n2671), .A2(n3741), .ZN(n2672) );
  NAND2_X1 U3379 ( .A1(n2673), .A2(n2672), .ZN(n2675) );
  NAND2_X1 U3380 ( .A1(n2674), .A2(n2675), .ZN(n3432) );
  NAND2_X1 U3381 ( .A1(n3431), .A2(n3432), .ZN(n2678) );
  INV_X1 U3382 ( .A(n2674), .ZN(n2677) );
  INV_X1 U3383 ( .A(n2675), .ZN(n2676) );
  NAND2_X1 U3384 ( .A1(n2677), .A2(n2676), .ZN(n3433) );
  NAND2_X1 U3385 ( .A1(n2678), .A2(n3433), .ZN(n3187) );
  NAND2_X1 U3386 ( .A1(n2398), .A2(REG0_REG_27__SCAN_IN), .ZN(n2684) );
  NAND2_X1 U3387 ( .A1(n3514), .A2(REG1_REG_27__SCAN_IN), .ZN(n2683) );
  OR2_X1 U3388 ( .A1(n2679), .A2(REG3_REG_27__SCAN_IN), .ZN(n2680) );
  NAND2_X1 U3389 ( .A1(n2679), .A2(REG3_REG_27__SCAN_IN), .ZN(n2724) );
  NAND2_X1 U3390 ( .A1(n2345), .A2(n3723), .ZN(n2682) );
  NAND2_X1 U3391 ( .A1(n3518), .A2(REG2_REG_27__SCAN_IN), .ZN(n2681) );
  NAND4_X1 U3392 ( .A1(n2684), .A2(n2683), .A3(n2682), .A4(n2681), .ZN(n3742)
         );
  NAND2_X1 U3393 ( .A1(n3742), .A2(n2671), .ZN(n2686) );
  NAND2_X1 U3394 ( .A1(n2352), .A2(DATAI_27_), .ZN(n2840) );
  INV_X1 U3395 ( .A(n2840), .ZN(n3722) );
  NAND2_X1 U3396 ( .A1(n3190), .A2(n3722), .ZN(n2685) );
  NAND2_X1 U3397 ( .A1(n2686), .A2(n2685), .ZN(n2688) );
  XNOR2_X1 U3398 ( .A(n2688), .B(n2687), .ZN(n3202) );
  NOR2_X1 U3399 ( .A1(n2029), .A2(n2840), .ZN(n2689) );
  AOI21_X1 U3400 ( .B1(n3742), .B2(n3195), .A(n2689), .ZN(n3200) );
  XNOR2_X1 U3401 ( .A(n3202), .B(n3200), .ZN(n3188) );
  XNOR2_X1 U3402 ( .A(n3187), .B(n3188), .ZN(n2713) );
  NAND2_X1 U3403 ( .A1(n2704), .A2(n2690), .ZN(n2691) );
  MUX2_X1 U3404 ( .A(n2690), .B(n2691), .S(B_REG_SCAN_IN), .Z(n2693) );
  INV_X1 U3405 ( .A(n2690), .ZN(n2856) );
  NOR4_X1 U3406 ( .A1(D_REG_31__SCAN_IN), .A2(D_REG_20__SCAN_IN), .A3(
        D_REG_3__SCAN_IN), .A4(D_REG_2__SCAN_IN), .ZN(n2702) );
  NOR4_X1 U3407 ( .A1(D_REG_4__SCAN_IN), .A2(D_REG_5__SCAN_IN), .A3(
        D_REG_6__SCAN_IN), .A4(D_REG_7__SCAN_IN), .ZN(n2701) );
  INV_X1 U3408 ( .A(D_REG_24__SCAN_IN), .ZN(n4474) );
  INV_X1 U3409 ( .A(D_REG_17__SCAN_IN), .ZN(n4476) );
  INV_X1 U3410 ( .A(D_REG_30__SCAN_IN), .ZN(n4473) );
  INV_X1 U3411 ( .A(D_REG_12__SCAN_IN), .ZN(n4477) );
  NAND4_X1 U3412 ( .A1(n4474), .A2(n4476), .A3(n4473), .A4(n4477), .ZN(n2699)
         );
  NOR4_X1 U3413 ( .A1(D_REG_13__SCAN_IN), .A2(D_REG_14__SCAN_IN), .A3(
        D_REG_15__SCAN_IN), .A4(D_REG_16__SCAN_IN), .ZN(n2697) );
  NOR4_X1 U3414 ( .A1(D_REG_10__SCAN_IN), .A2(D_REG_8__SCAN_IN), .A3(
        D_REG_9__SCAN_IN), .A4(D_REG_11__SCAN_IN), .ZN(n2696) );
  NOR4_X1 U3415 ( .A1(D_REG_23__SCAN_IN), .A2(D_REG_25__SCAN_IN), .A3(
        D_REG_26__SCAN_IN), .A4(D_REG_29__SCAN_IN), .ZN(n2695) );
  NOR4_X1 U3416 ( .A1(D_REG_18__SCAN_IN), .A2(D_REG_19__SCAN_IN), .A3(
        D_REG_21__SCAN_IN), .A4(D_REG_22__SCAN_IN), .ZN(n2694) );
  NAND4_X1 U3417 ( .A1(n2697), .A2(n2696), .A3(n2695), .A4(n2694), .ZN(n2698)
         );
  NOR4_X1 U3418 ( .A1(D_REG_27__SCAN_IN), .A2(D_REG_28__SCAN_IN), .A3(n2699), 
        .A4(n2698), .ZN(n2700) );
  AND3_X1 U3419 ( .A1(n2702), .A2(n2701), .A3(n2700), .ZN(n2703) );
  NOR2_X1 U3420 ( .A1(n2854), .A2(n2703), .ZN(n2831) );
  INV_X1 U3421 ( .A(n2704), .ZN(n4257) );
  OAI22_X1 U3422 ( .A1(n2854), .A2(D_REG_1__SCAN_IN), .B1(n4257), .B2(n2692), 
        .ZN(n2945) );
  OR2_X1 U3423 ( .A1(n2831), .A2(n2945), .ZN(n2705) );
  INV_X1 U3424 ( .A(n4459), .ZN(n2734) );
  NAND2_X1 U3425 ( .A1(n2730), .A2(n3681), .ZN(n2737) );
  NAND2_X1 U3426 ( .A1(n2734), .A2(n2737), .ZN(n2710) );
  INV_X1 U3427 ( .A(n2864), .ZN(n2709) );
  NAND2_X1 U3428 ( .A1(n2710), .A2(n2709), .ZN(n2711) );
  OR2_X1 U3429 ( .A1(n2862), .A2(n2711), .ZN(n2712) );
  NAND2_X1 U3430 ( .A1(n2713), .A2(n3434), .ZN(n2747) );
  INV_X1 U3431 ( .A(n2714), .ZN(n2715) );
  NAND2_X1 U3432 ( .A1(n4481), .A2(n2715), .ZN(n2716) );
  NOR2_X1 U3433 ( .A1(n2717), .A2(n2718), .ZN(n2719) );
  MUX2_X1 U3434 ( .A(n2718), .B(n2719), .S(IR_REG_28__SCAN_IN), .Z(n2722) );
  INV_X1 U3435 ( .A(n2720), .ZN(n2721) );
  INV_X1 U3436 ( .A(n4256), .ZN(n2827) );
  NAND2_X1 U3437 ( .A1(n3604), .A2(n2827), .ZN(n2723) );
  NAND2_X1 U3438 ( .A1(n2332), .A2(REG0_REG_28__SCAN_IN), .ZN(n2729) );
  NAND2_X1 U3439 ( .A1(n3514), .A2(REG1_REG_28__SCAN_IN), .ZN(n2728) );
  INV_X1 U3440 ( .A(REG3_REG_28__SCAN_IN), .ZN(n3204) );
  OR2_X1 U3441 ( .A1(n2724), .A2(n3204), .ZN(n2822) );
  NAND2_X1 U3442 ( .A1(n2724), .A2(n3204), .ZN(n2725) );
  NAND2_X1 U3443 ( .A1(n2345), .A2(n3210), .ZN(n2727) );
  NAND2_X1 U3444 ( .A1(n3518), .A2(REG2_REG_28__SCAN_IN), .ZN(n2726) );
  NAND4_X1 U3445 ( .A1(n2729), .A2(n2728), .A3(n2727), .A4(n2726), .ZN(n3716)
         );
  AOI22_X1 U3446 ( .A1(n3446), .A2(n3716), .B1(REG3_REG_27__SCAN_IN), .B2(
        U3149), .ZN(n2745) );
  OR2_X1 U3447 ( .A1(n2862), .A2(n4403), .ZN(n2732) );
  NAND2_X1 U3448 ( .A1(n2730), .A2(n4261), .ZN(n4465) );
  OR2_X1 U3449 ( .A1(n4465), .A2(n4258), .ZN(n4524) );
  INV_X1 U3450 ( .A(n2833), .ZN(n2731) );
  OAI21_X2 U3451 ( .B1(n2736), .B2(n2732), .A(n4413), .ZN(n3424) );
  NAND2_X1 U3452 ( .A1(n3604), .A2(n4256), .ZN(n2733) );
  AOI22_X1 U3453 ( .A1(n3722), .A2(n3424), .B1(n3449), .B2(n3753), .ZN(n2743)
         );
  NAND3_X1 U3454 ( .A1(n4403), .A2(n2734), .A3(n4261), .ZN(n2735) );
  NAND2_X1 U3455 ( .A1(n2736), .A2(n2735), .ZN(n2905) );
  AND2_X1 U3456 ( .A1(n2864), .A2(n2737), .ZN(n2832) );
  INV_X1 U3457 ( .A(n2863), .ZN(n2738) );
  NOR2_X1 U34580 ( .A1(n2832), .A2(n2738), .ZN(n2739) );
  AND2_X1 U34590 ( .A1(n2849), .A2(n2739), .ZN(n2740) );
  NAND2_X1 U3460 ( .A1(n2905), .A2(n2740), .ZN(n2741) );
  NAND2_X1 U3461 ( .A1(n3450), .A2(n3723), .ZN(n2742) );
  AND2_X1 U3462 ( .A1(n2745), .A2(n2744), .ZN(n2746) );
  NAND2_X1 U3463 ( .A1(n2747), .A2(n2746), .ZN(U3211) );
  NAND2_X1 U3464 ( .A1(n2749), .A2(n4439), .ZN(n2793) );
  NAND2_X1 U3465 ( .A1(n4447), .A2(n4446), .ZN(n4445) );
  NAND2_X1 U3466 ( .A1(n2748), .A2(n4439), .ZN(n2750) );
  INV_X1 U34670 ( .A(n2961), .ZN(n2752) );
  NAND2_X1 U3468 ( .A1(n2753), .A2(n2964), .ZN(n3469) );
  INV_X1 U34690 ( .A(n2753), .ZN(n2751) );
  NAND2_X1 U3470 ( .A1(n2751), .A2(n2970), .ZN(n3471) );
  INV_X1 U34710 ( .A(n2960), .ZN(n3530) );
  NAND2_X1 U3472 ( .A1(n2753), .A2(n2970), .ZN(n2754) );
  NOR2_X1 U34730 ( .A1(n3623), .A2(n3474), .ZN(n2756) );
  NAND2_X1 U3474 ( .A1(n3623), .A2(n3474), .ZN(n2755) );
  NAND2_X1 U34750 ( .A1(n2937), .A2(n3349), .ZN(n3476) );
  NAND2_X1 U3476 ( .A1(n3622), .A2(n3000), .ZN(n3479) );
  NAND2_X1 U34770 ( .A1(n3476), .A2(n3479), .ZN(n3532) );
  NAND2_X1 U3478 ( .A1(n3622), .A2(n3349), .ZN(n2757) );
  AND2_X1 U34790 ( .A1(n3621), .A2(n3317), .ZN(n2758) );
  NOR2_X1 U3480 ( .A1(n3620), .A2(n3425), .ZN(n2760) );
  NAND2_X1 U34810 ( .A1(n3620), .A2(n3425), .ZN(n2759) );
  NAND2_X1 U3482 ( .A1(n3011), .A2(n3055), .ZN(n2799) );
  NAND2_X1 U34830 ( .A1(n3619), .A2(n3030), .ZN(n3489) );
  NAND2_X1 U3484 ( .A1(n2799), .A2(n3489), .ZN(n3531) );
  NAND2_X1 U34850 ( .A1(n3040), .A2(n3531), .ZN(n2762) );
  NAND2_X1 U3486 ( .A1(n3619), .A2(n3055), .ZN(n2761) );
  NAND2_X1 U34870 ( .A1(n2762), .A2(n2761), .ZN(n3101) );
  AND2_X1 U3488 ( .A1(n3618), .A2(n3269), .ZN(n2764) );
  NAND2_X1 U34890 ( .A1(n3120), .A2(n3103), .ZN(n2763) );
  AND2_X1 U3490 ( .A1(n4406), .A2(n3240), .ZN(n2765) );
  NAND2_X1 U34910 ( .A1(n3144), .A2(n3402), .ZN(n3461) );
  NAND2_X1 U3492 ( .A1(n3616), .A2(n4417), .ZN(n3459) );
  NAND2_X1 U34930 ( .A1(n3461), .A2(n3459), .ZN(n4401) );
  NAND2_X1 U3494 ( .A1(n3144), .A2(n4417), .ZN(n2766) );
  NAND2_X1 U34950 ( .A1(n2767), .A2(n2766), .ZN(n3132) );
  NOR2_X1 U3496 ( .A1(n3401), .A2(n3286), .ZN(n2768) );
  INV_X1 U34970 ( .A(n3401), .ZN(n4404) );
  INV_X1 U3498 ( .A(n3286), .ZN(n3128) );
  AND2_X1 U34990 ( .A1(n3615), .A2(n3377), .ZN(n2770) );
  INV_X1 U3500 ( .A(n3615), .ZN(n3966) );
  INV_X1 U35010 ( .A(n3377), .ZN(n2803) );
  NAND2_X1 U3502 ( .A1(n3966), .A2(n2803), .ZN(n2769) );
  NAND2_X1 U35030 ( .A1(n2771), .A2(n3969), .ZN(n3939) );
  NAND2_X1 U3504 ( .A1(n3944), .A2(n2838), .ZN(n3455) );
  NAND2_X1 U35050 ( .A1(n3939), .A2(n3455), .ZN(n3957) );
  OR2_X1 U35060 ( .A1(n3942), .A2(n3309), .ZN(n3579) );
  NAND2_X1 U35070 ( .A1(n3942), .A2(n3309), .ZN(n3575) );
  NAND2_X1 U35080 ( .A1(n3579), .A2(n3575), .ZN(n3558) );
  NAND2_X1 U35090 ( .A1(n3901), .A2(n2774), .ZN(n2775) );
  NAND2_X1 U35100 ( .A1(n2775), .A2(n2264), .ZN(n3883) );
  NAND2_X1 U35110 ( .A1(n3904), .A2(n3886), .ZN(n3865) );
  NAND2_X1 U35120 ( .A1(n3872), .A2(n3891), .ZN(n3866) );
  NAND2_X1 U35130 ( .A1(n3865), .A2(n3866), .ZN(n3885) );
  NAND2_X1 U35140 ( .A1(n2777), .A2(n3876), .ZN(n2778) );
  NAND2_X1 U35150 ( .A1(n3613), .A2(n3362), .ZN(n3540) );
  NOR2_X1 U35160 ( .A1(n3613), .A2(n3362), .ZN(n3541) );
  NAND2_X1 U35170 ( .A1(n3849), .A2(n3835), .ZN(n2779) );
  INV_X1 U35180 ( .A(n3816), .ZN(n3611) );
  NOR2_X1 U35190 ( .A1(n3611), .A2(n3791), .ZN(n2782) );
  NAND2_X1 U35200 ( .A1(n3795), .A2(n2781), .ZN(n3787) );
  AND2_X1 U35210 ( .A1(n3830), .A2(n3820), .ZN(n2815) );
  INV_X1 U35220 ( .A(n2815), .ZN(n2780) );
  NAND2_X1 U35230 ( .A1(n3830), .A2(n2781), .ZN(n3783) );
  OAI22_X1 U35240 ( .A1(n2782), .A2(n3783), .B1(n3816), .B2(n3798), .ZN(n2783)
         );
  NAND2_X1 U35250 ( .A1(n3792), .A2(n3338), .ZN(n2785) );
  NAND2_X1 U35260 ( .A1(n3768), .A2(n2787), .ZN(n2786) );
  NAND2_X1 U35270 ( .A1(n3746), .A2(n2786), .ZN(n2788) );
  NOR2_X1 U35280 ( .A1(n3742), .A2(n3722), .ZN(n2791) );
  INV_X1 U35290 ( .A(n3742), .ZN(n3206) );
  AND2_X1 U35300 ( .A1(n3716), .A2(n3207), .ZN(n3686) );
  NOR2_X1 U35310 ( .A1(n3716), .A2(n3207), .ZN(n3687) );
  XNOR2_X1 U35320 ( .A(n2951), .B(n4258), .ZN(n2792) );
  NAND2_X1 U35330 ( .A1(n2792), .A2(n3681), .ZN(n4448) );
  INV_X1 U35340 ( .A(n3625), .ZN(n4444) );
  NAND2_X1 U35350 ( .A1(n4444), .A2(n2837), .ZN(n3534) );
  NAND2_X1 U35360 ( .A1(n4436), .A2(n2793), .ZN(n2794) );
  NAND2_X1 U35370 ( .A1(n2794), .A2(n2960), .ZN(n2938) );
  XNOR2_X1 U35380 ( .A(n3623), .B(n3474), .ZN(n2939) );
  NAND2_X1 U35390 ( .A1(n3473), .A2(n3474), .ZN(n3475) );
  INV_X1 U35400 ( .A(n3476), .ZN(n2795) );
  NAND2_X1 U35410 ( .A1(n2796), .A2(n3479), .ZN(n2980) );
  AND2_X1 U35420 ( .A1(n3621), .A2(n2981), .ZN(n2978) );
  NAND2_X1 U35430 ( .A1(n2797), .A2(n3317), .ZN(n3485) );
  INV_X1 U35440 ( .A(n3425), .ZN(n3010) );
  NAND2_X1 U35450 ( .A1(n3620), .A2(n3010), .ZN(n3484) );
  NAND2_X1 U35460 ( .A1(n3009), .A2(n3484), .ZN(n2798) );
  INV_X1 U35470 ( .A(n3620), .ZN(n2982) );
  NAND2_X1 U35480 ( .A1(n2982), .A2(n3425), .ZN(n3481) );
  NAND2_X1 U35490 ( .A1(n2798), .A2(n3481), .ZN(n3029) );
  INV_X1 U35500 ( .A(n2799), .ZN(n2800) );
  NAND2_X1 U35510 ( .A1(n3120), .A2(n3269), .ZN(n3494) );
  NAND2_X1 U35520 ( .A1(n3618), .A2(n3103), .ZN(n3490) );
  AND2_X1 U35530 ( .A1(n3617), .A2(n3121), .ZN(n3044) );
  NAND2_X1 U35540 ( .A1(n3104), .A2(n3050), .ZN(n3495) );
  NAND2_X1 U35550 ( .A1(n4406), .A2(n3143), .ZN(n3458) );
  NAND2_X1 U35560 ( .A1(n2802), .A2(n3240), .ZN(n3457) );
  NOR2_X1 U35570 ( .A1(n3401), .A2(n3128), .ZN(n3463) );
  NAND2_X1 U35580 ( .A1(n3615), .A2(n2803), .ZN(n3157) );
  NAND2_X1 U35590 ( .A1(n3401), .A2(n3128), .ZN(n3155) );
  AND2_X1 U35600 ( .A1(n3157), .A2(n3155), .ZN(n3462) );
  NAND2_X1 U35610 ( .A1(n3156), .A2(n3462), .ZN(n2804) );
  NAND2_X1 U35620 ( .A1(n3966), .A2(n3377), .ZN(n3465) );
  INV_X1 U35630 ( .A(n3957), .ZN(n3961) );
  NAND2_X1 U35640 ( .A1(n3960), .A2(n3961), .ZN(n3959) );
  NAND2_X1 U35650 ( .A1(n2805), .A2(n3447), .ZN(n3464) );
  NAND2_X1 U35660 ( .A1(n3963), .A2(n3947), .ZN(n3456) );
  NAND2_X1 U35670 ( .A1(n3464), .A2(n3456), .ZN(n3940) );
  INV_X1 U35680 ( .A(n3939), .ZN(n3574) );
  NOR2_X1 U35690 ( .A1(n3940), .A2(n3574), .ZN(n2806) );
  NAND2_X1 U35700 ( .A1(n3959), .A2(n2806), .ZN(n2807) );
  NAND2_X1 U35710 ( .A1(n2807), .A2(n3456), .ZN(n3922) );
  NAND2_X1 U35720 ( .A1(n3887), .A2(n3876), .ZN(n2808) );
  AND2_X1 U35730 ( .A1(n3866), .A2(n2808), .ZN(n2810) );
  OR2_X1 U35740 ( .A1(n3923), .A2(n3328), .ZN(n3862) );
  NAND2_X1 U35750 ( .A1(n2810), .A2(n3862), .ZN(n3578) );
  AND2_X1 U35760 ( .A1(n3613), .A2(n3854), .ZN(n3585) );
  NAND2_X1 U35770 ( .A1(n3923), .A2(n3328), .ZN(n3863) );
  NAND2_X1 U35780 ( .A1(n3865), .A2(n3863), .ZN(n2811) );
  NOR2_X1 U35790 ( .A1(n3887), .A2(n3876), .ZN(n2809) );
  AOI21_X1 U35800 ( .B1(n2811), .B2(n2810), .A(n2809), .ZN(n3845) );
  INV_X1 U35810 ( .A(n3613), .ZN(n3870) );
  NAND2_X1 U3582 ( .A1(n3870), .A2(n3362), .ZN(n2812) );
  AND2_X1 U3583 ( .A1(n3845), .A2(n2812), .ZN(n3584) );
  NOR2_X1 U3584 ( .A1(n3584), .A2(n3585), .ZN(n3504) );
  INV_X1 U3585 ( .A(n3504), .ZN(n2813) );
  NAND2_X1 U3586 ( .A1(n3849), .A2(n3829), .ZN(n3785) );
  AND2_X1 U3587 ( .A1(n3787), .A2(n3785), .ZN(n3582) );
  NOR2_X1 U3588 ( .A1(n3849), .A2(n3829), .ZN(n3786) );
  NOR2_X1 U3589 ( .A1(n3816), .A2(n3791), .ZN(n3554) );
  NOR2_X1 U3590 ( .A1(n3554), .A2(n2815), .ZN(n3508) );
  INV_X1 U3591 ( .A(n3508), .ZN(n2816) );
  AOI21_X1 U3592 ( .B1(n3786), .B2(n3787), .A(n2816), .ZN(n3587) );
  INV_X1 U3593 ( .A(n3587), .ZN(n2817) );
  NAND2_X1 U3594 ( .A1(n3816), .A2(n3791), .ZN(n3553) );
  NAND2_X1 U3595 ( .A1(n3756), .A2(n3338), .ZN(n3556) );
  NAND2_X1 U3596 ( .A1(n3553), .A2(n3556), .ZN(n3588) );
  NAND2_X1 U3597 ( .A1(n3768), .A2(n3757), .ZN(n3737) );
  NAND2_X1 U3598 ( .A1(n3719), .A2(n3741), .ZN(n3535) );
  NAND2_X1 U3599 ( .A1(n3737), .A2(n3535), .ZN(n3571) );
  INV_X1 U3600 ( .A(n3571), .ZN(n2818) );
  OR2_X1 U3601 ( .A1(n3768), .A2(n3757), .ZN(n3555) );
  NAND2_X1 U3602 ( .A1(n3792), .A2(n3774), .ZN(n3748) );
  AND2_X1 U3603 ( .A1(n3555), .A2(n3748), .ZN(n3736) );
  NAND2_X1 U3604 ( .A1(n3753), .A2(n2839), .ZN(n3568) );
  OAI21_X1 U3605 ( .B1(n3736), .B2(n3571), .A(n3568), .ZN(n3511) );
  AOI21_X1 U3606 ( .B1(n3747), .B2(n2818), .A(n3511), .ZN(n3714) );
  AND2_X1 U3607 ( .A1(n3742), .A2(n2840), .ZN(n3513) );
  NOR2_X1 U3608 ( .A1(n3742), .A2(n2840), .ZN(n3572) );
  NAND2_X1 U3609 ( .A1(n3714), .A2(n3713), .ZN(n3712) );
  INV_X1 U3610 ( .A(n3572), .ZN(n2819) );
  NAND2_X1 U3611 ( .A1(n3712), .A2(n2819), .ZN(n3689) );
  XOR2_X1 U3612 ( .A(n3700), .B(n3689), .Z(n2830) );
  NAND2_X1 U3613 ( .A1(n4260), .A2(n4259), .ZN(n2821) );
  NAND2_X1 U3614 ( .A1(n4258), .A2(n4261), .ZN(n2820) );
  NAND2_X1 U3615 ( .A1(n3514), .A2(REG1_REG_29__SCAN_IN), .ZN(n2826) );
  NAND2_X1 U3616 ( .A1(n2332), .A2(REG0_REG_29__SCAN_IN), .ZN(n2825) );
  INV_X1 U3617 ( .A(n2822), .ZN(n3698) );
  NAND2_X1 U3618 ( .A1(n2345), .A2(n3698), .ZN(n2824) );
  NAND2_X1 U3619 ( .A1(n3518), .A2(REG2_REG_29__SCAN_IN), .ZN(n2823) );
  NAND4_X1 U3620 ( .A1(n2826), .A2(n2825), .A3(n2824), .A4(n2823), .ZN(n3609)
         );
  INV_X1 U3621 ( .A(n3207), .ZN(n3699) );
  AOI22_X1 U3622 ( .A1(n3609), .A2(n4441), .B1(n4440), .B2(n3699), .ZN(n2828)
         );
  OAI21_X1 U3623 ( .B1(n3206), .B2(n4443), .A(n2828), .ZN(n2829) );
  AOI21_X1 U3624 ( .B1(n2830), .B2(n4461), .A(n2829), .ZN(n3178) );
  OAI21_X1 U3625 ( .B1(n3183), .B2(n4535), .A(n3178), .ZN(n2845) );
  INV_X1 U3626 ( .A(n2831), .ZN(n2947) );
  OR2_X1 U3627 ( .A1(n2862), .A2(n2832), .ZN(n2904) );
  NOR2_X1 U3628 ( .A1(n2904), .A2(n2833), .ZN(n2834) );
  NAND3_X1 U3629 ( .A1(n2947), .A2(n2834), .A3(n2945), .ZN(n2844) );
  INV_X1 U3630 ( .A(n2946), .ZN(n2835) );
  MUX2_X1 U3631 ( .A(REG0_REG_28__SCAN_IN), .B(n2845), .S(n4560), .Z(n2836) );
  INV_X1 U3632 ( .A(n2836), .ZN(n2843) );
  NAND2_X1 U3633 ( .A1(n4460), .A2(n4453), .ZN(n4452) );
  NAND2_X1 U3634 ( .A1(n4516), .A2(n2953), .ZN(n2992) );
  NAND2_X1 U3635 ( .A1(n3034), .A2(n3030), .ZN(n3035) );
  NAND2_X1 U3636 ( .A1(n4418), .A2(n4417), .ZN(n4416) );
  NAND2_X1 U3637 ( .A1(n3968), .A2(n3947), .ZN(n3949) );
  NAND2_X1 U3638 ( .A1(n3720), .A2(n3207), .ZN(n3704) );
  OAI21_X1 U3639 ( .B1(n3720), .B2(n3207), .A(n3704), .ZN(n3175) );
  NAND2_X1 U3640 ( .A1(n2843), .A2(n2842), .ZN(U3514) );
  MUX2_X1 U3641 ( .A(REG1_REG_28__SCAN_IN), .B(n2845), .S(n4579), .Z(n2846) );
  INV_X1 U3642 ( .A(n2846), .ZN(n2848) );
  NAND2_X1 U3643 ( .A1(n2848), .A2(n2847), .ZN(U3546) );
  INV_X1 U3644 ( .A(DATAI_24_), .ZN(n2850) );
  MUX2_X1 U3645 ( .A(n2690), .B(n2850), .S(U3149), .Z(n2851) );
  INV_X1 U3646 ( .A(n2851), .ZN(U3328) );
  INV_X1 U3647 ( .A(DATAI_29_), .ZN(n4030) );
  NAND2_X1 U3648 ( .A1(n2852), .A2(STATE_REG_SCAN_IN), .ZN(n2853) );
  OAI21_X1 U3649 ( .B1(STATE_REG_SCAN_IN), .B2(n4030), .A(n2853), .ZN(U3323)
         );
  INV_X1 U3650 ( .A(n2862), .ZN(n2855) );
  INV_X1 U3651 ( .A(D_REG_0__SCAN_IN), .ZN(n2858) );
  NOR3_X1 U3652 ( .A1(n2692), .A2(n2856), .A3(n2859), .ZN(n2857) );
  AOI21_X1 U3653 ( .B1(n4480), .B2(n2858), .A(n2857), .ZN(U3458) );
  INV_X1 U3654 ( .A(D_REG_1__SCAN_IN), .ZN(n2861) );
  NOR3_X1 U3655 ( .A1(n4257), .A2(n2692), .A3(n2859), .ZN(n2860) );
  AOI21_X1 U3656 ( .B1(n4480), .B2(n2861), .A(n2860), .ZN(U3459) );
  OR2_X1 U3657 ( .A1(n2863), .A2(U3149), .ZN(n3607) );
  NAND2_X1 U3658 ( .A1(n2862), .A2(n3607), .ZN(n2876) );
  NAND2_X1 U3659 ( .A1(n2864), .A2(n2863), .ZN(n2865) );
  INV_X1 U3660 ( .A(n2875), .ZN(n2866) );
  NOR2_X1 U3661 ( .A1(n4392), .A2(U4043), .ZN(U3148) );
  INV_X1 U3662 ( .A(DATAO_REG_12__SCAN_IN), .ZN(n2868) );
  NAND2_X1 U3663 ( .A1(n3401), .A2(U4043), .ZN(n2867) );
  OAI21_X1 U3664 ( .B1(U4043), .B2(n2868), .A(n2867), .ZN(U3562) );
  INV_X1 U3665 ( .A(REG1_REG_3__SCAN_IN), .ZN(n4566) );
  INV_X1 U3666 ( .A(REG1_REG_2__SCAN_IN), .ZN(n4564) );
  MUX2_X1 U3667 ( .A(REG1_REG_2__SCAN_IN), .B(n4564), .S(n4267), .Z(n3640) );
  INV_X1 U3668 ( .A(REG1_REG_1__SCAN_IN), .ZN(n4562) );
  AND2_X1 U3669 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n3629)
         );
  NAND2_X1 U3670 ( .A1(n4268), .A2(REG1_REG_1__SCAN_IN), .ZN(n2869) );
  NAND2_X1 U3671 ( .A1(n3628), .A2(n2869), .ZN(n3639) );
  NAND2_X1 U3672 ( .A1(n3640), .A2(n3639), .ZN(n3638) );
  NAND2_X1 U3673 ( .A1(n4267), .A2(REG1_REG_2__SCAN_IN), .ZN(n2870) );
  NAND2_X1 U3674 ( .A1(n3638), .A2(n2870), .ZN(n2871) );
  NOR2_X1 U3675 ( .A1(n4566), .A2(n2895), .ZN(n2894) );
  AND2_X1 U3676 ( .A1(n2871), .A2(n4266), .ZN(n2872) );
  INV_X1 U3677 ( .A(n4502), .ZN(n4292) );
  INV_X1 U3678 ( .A(REG1_REG_5__SCAN_IN), .ZN(n4570) );
  AOI22_X1 U3679 ( .A1(REG1_REG_5__SCAN_IN), .A2(n4292), .B1(n4502), .B2(n4570), .ZN(n4283) );
  NOR2_X1 U3680 ( .A1(n2873), .A2(n4501), .ZN(n2874) );
  INV_X1 U3681 ( .A(REG1_REG_6__SCAN_IN), .ZN(n4296) );
  XNOR2_X1 U3682 ( .A(n4501), .B(n2873), .ZN(n4295) );
  NOR2_X1 U3683 ( .A1(n4296), .A2(n4295), .ZN(n4294) );
  INV_X1 U3684 ( .A(n4264), .ZN(n2891) );
  INV_X1 U3685 ( .A(REG1_REG_7__SCAN_IN), .ZN(n4572) );
  NAND2_X1 U3686 ( .A1(n2891), .A2(n4572), .ZN(n3082) );
  NAND2_X1 U3687 ( .A1(n4264), .A2(REG1_REG_7__SCAN_IN), .ZN(n3083) );
  NAND2_X1 U3688 ( .A1(n3082), .A2(n3083), .ZN(n2879) );
  XNOR2_X1 U3689 ( .A(n2877), .B(IR_REG_27__SCAN_IN), .ZN(n4277) );
  OR2_X1 U3690 ( .A1(n4280), .A2(n4277), .ZN(n4293) );
  OAI21_X1 U3691 ( .B1(n3084), .B2(n2879), .A(n4394), .ZN(n2878) );
  AOI21_X1 U3692 ( .B1(n3084), .B2(n2879), .A(n2878), .ZN(n2893) );
  INV_X1 U3693 ( .A(REG2_REG_5__SCAN_IN), .ZN(n2988) );
  AOI22_X1 U3694 ( .A1(REG2_REG_5__SCAN_IN), .A2(n4502), .B1(n4292), .B2(n2988), .ZN(n4289) );
  INV_X1 U3695 ( .A(n4267), .ZN(n3636) );
  INV_X1 U3696 ( .A(REG2_REG_1__SCAN_IN), .ZN(n2880) );
  INV_X1 U3697 ( .A(REG2_REG_0__SCAN_IN), .ZN(n4469) );
  NOR2_X1 U3698 ( .A1(n4505), .A2(n4469), .ZN(n3627) );
  NAND2_X1 U3699 ( .A1(n4268), .A2(REG2_REG_1__SCAN_IN), .ZN(n3642) );
  OAI21_X1 U3700 ( .B1(n4105), .B2(n3636), .A(n3645), .ZN(n2881) );
  INV_X1 U3701 ( .A(n4265), .ZN(n2921) );
  XNOR2_X1 U3702 ( .A(n2039), .B(n2921), .ZN(n2909) );
  INV_X1 U3703 ( .A(REG2_REG_4__SCAN_IN), .ZN(n2882) );
  OAI22_X1 U3704 ( .A1(n2909), .A2(n2882), .B1(n2039), .B2(n2921), .ZN(n4288)
         );
  NAND2_X1 U3705 ( .A1(n2884), .A2(n2883), .ZN(n2885) );
  NAND2_X1 U3706 ( .A1(n2885), .A2(n4299), .ZN(n2888) );
  MUX2_X1 U3707 ( .A(REG2_REG_7__SCAN_IN), .B(n3038), .S(n4264), .Z(n2887) );
  AND2_X1 U3708 ( .A1(n4256), .A2(n4277), .ZN(n3603) );
  INV_X1 U3709 ( .A(n3603), .ZN(n2886) );
  NOR2_X2 U3710 ( .A1(n2886), .A2(n4280), .ZN(n4346) );
  NAND2_X1 U3711 ( .A1(n2887), .A2(n2888), .ZN(n3067) );
  OAI211_X1 U3712 ( .C1(n2888), .C2(n2887), .A(n4346), .B(n3067), .ZN(n2890)
         );
  NOR2_X1 U3713 ( .A1(n4039), .A2(STATE_REG_SCAN_IN), .ZN(n3056) );
  AOI21_X1 U3714 ( .B1(n4392), .B2(ADDR_REG_7__SCAN_IN), .A(n3056), .ZN(n2889)
         );
  OAI211_X1 U3715 ( .C1(n4399), .C2(n2891), .A(n2890), .B(n2889), .ZN(n2892)
         );
  OR2_X1 U3716 ( .A1(n2893), .A2(n2892), .ZN(U3247) );
  AOI211_X1 U3717 ( .C1(n4566), .C2(n2895), .A(n2894), .B(n4293), .ZN(n2901)
         );
  OAI211_X1 U3718 ( .C1(REG2_REG_3__SCAN_IN), .C2(n2897), .A(n4346), .B(n2896), 
        .ZN(n2899) );
  NOR2_X1 U3719 ( .A1(STATE_REG_SCAN_IN), .A2(n3249), .ZN(n3248) );
  AOI21_X1 U3720 ( .B1(n4392), .B2(ADDR_REG_3__SCAN_IN), .A(n3248), .ZN(n2898)
         );
  OAI211_X1 U3721 ( .C1(n4399), .C2(n2210), .A(n2899), .B(n2898), .ZN(n2900)
         );
  OR2_X1 U3722 ( .A1(n2901), .A2(n2900), .ZN(U3243) );
  XNOR2_X1 U3723 ( .A(n2903), .B(n2902), .ZN(n2913) );
  INV_X1 U3724 ( .A(n2904), .ZN(n2948) );
  NAND2_X1 U3725 ( .A1(n2905), .A2(n2948), .ZN(n2933) );
  OAI22_X1 U3726 ( .A1(n3389), .A2(n4460), .B1(n3387), .B2(n2749), .ZN(n2906)
         );
  AOI21_X1 U3727 ( .B1(REG3_REG_0__SCAN_IN), .B2(n2933), .A(n2906), .ZN(n2907)
         );
  OAI21_X1 U3728 ( .B1(n3394), .B2(n2913), .A(n2907), .ZN(U3229) );
  AND2_X1 U3729 ( .A1(U3149), .A2(REG3_REG_4__SCAN_IN), .ZN(n3348) );
  OAI21_X1 U3730 ( .B1(REG1_REG_4__SCAN_IN), .B2(n2908), .A(n4394), .ZN(n2917)
         );
  XNOR2_X1 U3731 ( .A(REG2_REG_4__SCAN_IN), .B(n2909), .ZN(n2910) );
  NAND2_X1 U3732 ( .A1(n4346), .A2(n2910), .ZN(n2916) );
  NAND2_X1 U3733 ( .A1(n4277), .A2(n4469), .ZN(n2911) );
  AND2_X1 U3734 ( .A1(n4256), .A2(n2911), .ZN(n4276) );
  INV_X1 U3735 ( .A(n4277), .ZN(n2912) );
  NAND3_X1 U3736 ( .A1(n2913), .A2(n4256), .A3(n2912), .ZN(n2915) );
  AOI21_X1 U3737 ( .B1(n3603), .B2(n3627), .A(n3624), .ZN(n2914) );
  OAI211_X1 U3738 ( .C1(IR_REG_0__SCAN_IN), .C2(n4276), .A(n2915), .B(n2914), 
        .ZN(n3649) );
  OAI211_X1 U3739 ( .C1(n2918), .C2(n2917), .A(n2916), .B(n3649), .ZN(n2919)
         );
  AOI211_X1 U3740 ( .C1(n4392), .C2(ADDR_REG_4__SCAN_IN), .A(n3348), .B(n2919), 
        .ZN(n2920) );
  OAI21_X1 U3741 ( .B1(n2921), .B2(n4399), .A(n2920), .ZN(U3244) );
  XNOR2_X1 U3742 ( .A(n2922), .B(n2923), .ZN(n2927) );
  AOI22_X1 U3743 ( .A1(n2751), .A2(n3446), .B1(n3449), .B2(n3625), .ZN(n2924)
         );
  OAI21_X1 U3744 ( .B1(n3389), .B2(n4453), .A(n2924), .ZN(n2925) );
  AOI21_X1 U3745 ( .B1(REG3_REG_1__SCAN_IN), .B2(n2933), .A(n2925), .ZN(n2926)
         );
  OAI21_X1 U3746 ( .B1(n2927), .B2(n3394), .A(n2926), .ZN(U3219) );
  AOI21_X1 U3747 ( .B1(n2928), .B2(n2930), .A(n2929), .ZN(n2935) );
  AOI22_X1 U3748 ( .A1(n2748), .A2(n3449), .B1(n3446), .B2(n3623), .ZN(n2931)
         );
  OAI21_X1 U3749 ( .B1(n3389), .B2(n2970), .A(n2931), .ZN(n2932) );
  AOI21_X1 U3750 ( .B1(REG3_REG_2__SCAN_IN), .B2(n2933), .A(n2932), .ZN(n2934)
         );
  OAI21_X1 U3751 ( .B1(n2935), .B2(n3394), .A(n2934), .ZN(U3234) );
  XNOR2_X1 U3752 ( .A(n2936), .B(n2939), .ZN(n4525) );
  OAI22_X1 U3753 ( .A1(n2937), .A2(n4464), .B1(n4403), .B2(n2953), .ZN(n2943)
         );
  INV_X1 U3754 ( .A(n2939), .ZN(n3564) );
  NAND3_X1 U3755 ( .A1(n2938), .A2(n3469), .A3(n3564), .ZN(n2940) );
  AOI21_X1 U3756 ( .B1(n2941), .B2(n2940), .A(n4409), .ZN(n2942) );
  AOI211_X1 U3757 ( .C1(n4407), .C2(n2751), .A(n2943), .B(n2942), .ZN(n2944)
         );
  OAI21_X1 U3758 ( .B1(n4525), .B2(n4448), .A(n2944), .ZN(n4527) );
  INV_X1 U3759 ( .A(n4527), .ZN(n2958) );
  INV_X1 U3760 ( .A(n2945), .ZN(n2949) );
  NAND4_X1 U3761 ( .A1(n2949), .A2(n2948), .A3(n2947), .A4(n2946), .ZN(n2950)
         );
  INV_X1 U3762 ( .A(n4525), .ZN(n2956) );
  NOR2_X1 U3763 ( .A1(n2951), .A2(n3681), .ZN(n2952) );
  NAND2_X1 U3764 ( .A1(n3935), .A2(n2952), .ZN(n2977) );
  INV_X1 U3765 ( .A(n2977), .ZN(n4467) );
  AND2_X1 U3766 ( .A1(n3935), .A2(n3681), .ZN(n3894) );
  OAI21_X1 U3767 ( .B1(n4516), .B2(n2953), .A(n2992), .ZN(n4523) );
  AOI22_X1 U3768 ( .A1(n4471), .A2(REG2_REG_3__SCAN_IN), .B1(n4466), .B2(n3249), .ZN(n2954) );
  OAI21_X1 U3769 ( .B1(n3952), .B2(n4523), .A(n2954), .ZN(n2955) );
  AOI21_X1 U3770 ( .B1(n2956), .B2(n4467), .A(n2955), .ZN(n2957) );
  OAI21_X1 U3771 ( .B1(n2958), .B2(n4471), .A(n2957), .ZN(U3287) );
  NAND2_X1 U3772 ( .A1(n2961), .A2(n2960), .ZN(n2962) );
  NAND2_X1 U3773 ( .A1(n2959), .A2(n2962), .ZN(n4521) );
  INV_X1 U3774 ( .A(n4521), .ZN(n2975) );
  NAND3_X1 U3775 ( .A1(n3530), .A2(n2793), .A3(n4436), .ZN(n2963) );
  NAND2_X1 U3776 ( .A1(n2938), .A2(n2963), .ZN(n2967) );
  AOI22_X1 U3777 ( .A1(n3623), .A2(n4441), .B1(n2964), .B2(n4440), .ZN(n2965)
         );
  OAI21_X1 U3778 ( .B1(n2749), .B2(n4443), .A(n2965), .ZN(n2966) );
  AOI21_X1 U3779 ( .B1(n2967), .B2(n4461), .A(n2966), .ZN(n2969) );
  NAND2_X1 U3780 ( .A1(n4521), .A2(n4462), .ZN(n2968) );
  AND2_X1 U3781 ( .A1(n2969), .A2(n2968), .ZN(n4518) );
  MUX2_X1 U3782 ( .A(n4518), .B(n4105), .S(n4471), .Z(n2974) );
  INV_X1 U3783 ( .A(n4452), .ZN(n2971) );
  NOR2_X1 U3784 ( .A1(n2971), .A2(n2970), .ZN(n4517) );
  NOR3_X1 U3785 ( .A1(n3952), .A2(n4516), .A3(n4517), .ZN(n2972) );
  AOI21_X1 U3786 ( .B1(n4466), .B2(REG3_REG_2__SCAN_IN), .A(n2972), .ZN(n2973)
         );
  OAI211_X1 U3787 ( .C1(n2975), .C2(n2977), .A(n2974), .B(n2973), .ZN(U3288)
         );
  NAND2_X1 U3788 ( .A1(n3935), .A2(n4462), .ZN(n2976) );
  INV_X1 U3789 ( .A(n2978), .ZN(n3478) );
  NAND2_X1 U3790 ( .A1(n3478), .A2(n3485), .ZN(n3551) );
  XNOR2_X1 U3791 ( .A(n2979), .B(n3551), .ZN(n4536) );
  XOR2_X1 U3792 ( .A(n3551), .B(n2980), .Z(n2985) );
  OAI22_X1 U3793 ( .A1(n2982), .A2(n4464), .B1(n4403), .B2(n2981), .ZN(n2983)
         );
  AOI21_X1 U3794 ( .B1(n4407), .B2(n3622), .A(n2983), .ZN(n2984) );
  OAI21_X1 U3795 ( .B1(n2985), .B2(n4409), .A(n2984), .ZN(n4537) );
  NAND2_X1 U3796 ( .A1(n4537), .A2(n3972), .ZN(n2991) );
  AND2_X1 U3797 ( .A1(n2993), .A2(n3317), .ZN(n2986) );
  NOR2_X1 U3798 ( .A1(n3015), .A2(n2986), .ZN(n4539) );
  INV_X1 U3799 ( .A(n3318), .ZN(n2987) );
  OAI22_X1 U3800 ( .A1(n3935), .A2(n2988), .B1(n2987), .B2(n4413), .ZN(n2989)
         );
  AOI21_X1 U3801 ( .B1(n4539), .B2(n4455), .A(n2989), .ZN(n2990) );
  OAI211_X1 U3802 ( .C1(n3955), .C2(n4536), .A(n2991), .B(n2990), .ZN(U3285)
         );
  AOI21_X1 U3803 ( .B1(n2992), .B2(n3349), .A(n2841), .ZN(n2994) );
  NAND2_X1 U3804 ( .A1(n2994), .A2(n2993), .ZN(n4530) );
  NOR2_X1 U3805 ( .A1(n4530), .A2(n4261), .ZN(n3005) );
  INV_X1 U3806 ( .A(n3532), .ZN(n2996) );
  XNOR2_X1 U3807 ( .A(n2995), .B(n2996), .ZN(n4529) );
  NAND2_X1 U3808 ( .A1(n4529), .A2(n4462), .ZN(n3004) );
  XNOR2_X1 U3809 ( .A(n2997), .B(n2996), .ZN(n3002) );
  NAND2_X1 U3810 ( .A1(n3623), .A2(n4407), .ZN(n2999) );
  NAND2_X1 U3811 ( .A1(n3621), .A2(n4441), .ZN(n2998) );
  OAI211_X1 U3812 ( .C1(n4403), .C2(n3000), .A(n2999), .B(n2998), .ZN(n3001)
         );
  AOI21_X1 U3813 ( .B1(n3002), .B2(n4461), .A(n3001), .ZN(n3003) );
  NAND2_X1 U3814 ( .A1(n3004), .A2(n3003), .ZN(n4533) );
  AOI211_X1 U3815 ( .C1(n4466), .C2(n3350), .A(n3005), .B(n4533), .ZN(n3007)
         );
  AOI22_X1 U3816 ( .A1(n4529), .A2(n4467), .B1(REG2_REG_4__SCAN_IN), .B2(n4471), .ZN(n3006) );
  OAI21_X1 U3817 ( .B1(n3007), .B2(n4471), .A(n3006), .ZN(U3286) );
  NAND2_X1 U3818 ( .A1(n3481), .A2(n3484), .ZN(n3528) );
  XNOR2_X1 U3819 ( .A(n3008), .B(n3528), .ZN(n3024) );
  INV_X1 U3820 ( .A(n3024), .ZN(n3022) );
  XNOR2_X1 U3821 ( .A(n3009), .B(n3528), .ZN(n3014) );
  OAI22_X1 U3822 ( .A1(n3011), .A2(n4464), .B1(n4403), .B2(n3010), .ZN(n3012)
         );
  AOI21_X1 U3823 ( .B1(n4407), .B2(n3621), .A(n3012), .ZN(n3013) );
  OAI21_X1 U3824 ( .B1(n3014), .B2(n4409), .A(n3013), .ZN(n3023) );
  NAND2_X1 U3825 ( .A1(n3023), .A2(n3972), .ZN(n3021) );
  INV_X1 U3826 ( .A(n3015), .ZN(n3016) );
  AOI21_X1 U3827 ( .B1(n3425), .B2(n3016), .A(n3034), .ZN(n3026) );
  INV_X1 U3828 ( .A(n4471), .ZN(n3972) );
  INV_X1 U3829 ( .A(REG2_REG_6__SCAN_IN), .ZN(n3018) );
  OAI22_X1 U3830 ( .A1(n3972), .A2(n3018), .B1(n3017), .B2(n4413), .ZN(n3019)
         );
  AOI21_X1 U3831 ( .B1(n3026), .B2(n4455), .A(n3019), .ZN(n3020) );
  OAI211_X1 U3832 ( .C1(n3955), .C2(n3022), .A(n3021), .B(n3020), .ZN(U3284)
         );
  AOI21_X1 U3833 ( .B1(n4550), .B2(n3024), .A(n3023), .ZN(n3028) );
  INV_X1 U3834 ( .A(n4251), .ZN(n4207) );
  AOI22_X1 U3835 ( .A1(n3026), .A2(n4207), .B1(n4558), .B2(REG0_REG_6__SCAN_IN), .ZN(n3025) );
  OAI21_X1 U3836 ( .B1(n3028), .B2(n4558), .A(n3025), .ZN(U3479) );
  INV_X1 U3837 ( .A(n4193), .ZN(n3985) );
  AOI22_X1 U3838 ( .A1(n3026), .A2(n3985), .B1(n4576), .B2(REG1_REG_6__SCAN_IN), .ZN(n3027) );
  OAI21_X1 U3839 ( .B1(n3028), .B2(n4576), .A(n3027), .ZN(U3524) );
  XNOR2_X1 U3840 ( .A(n3029), .B(n3531), .ZN(n3033) );
  OAI22_X1 U3841 ( .A1(n3120), .A2(n4464), .B1(n4403), .B2(n3030), .ZN(n3031)
         );
  AOI21_X1 U3842 ( .B1(n4407), .B2(n3620), .A(n3031), .ZN(n3032) );
  OAI21_X1 U3843 ( .B1(n3033), .B2(n4409), .A(n3032), .ZN(n4542) );
  INV_X1 U3844 ( .A(n4542), .ZN(n3043) );
  INV_X1 U3845 ( .A(n3034), .ZN(n3036) );
  INV_X1 U3846 ( .A(n3035), .ZN(n3100) );
  AOI211_X1 U3847 ( .C1(n3055), .C2(n3036), .A(n2841), .B(n3100), .ZN(n4543)
         );
  INV_X1 U3848 ( .A(REG2_REG_7__SCAN_IN), .ZN(n3038) );
  INV_X1 U3849 ( .A(n3064), .ZN(n3037) );
  OAI22_X1 U3850 ( .A1(n3935), .A2(n3038), .B1(n3037), .B2(n4413), .ZN(n3039)
         );
  AOI21_X1 U3851 ( .B1(n4543), .B2(n3894), .A(n3039), .ZN(n3042) );
  XOR2_X1 U3852 ( .A(n3040), .B(n3531), .Z(n4544) );
  NAND2_X1 U3853 ( .A1(n4544), .A2(n3808), .ZN(n3041) );
  OAI211_X1 U3854 ( .C1(n3043), .C2(n4471), .A(n3042), .B(n3041), .ZN(U3283)
         );
  INV_X1 U3855 ( .A(n3044), .ZN(n3496) );
  NAND2_X1 U3856 ( .A1(n3496), .A2(n3495), .ZN(n3552) );
  XNOR2_X1 U3857 ( .A(n3045), .B(n3552), .ZN(n3048) );
  AOI22_X1 U3858 ( .A1(n4406), .A2(n4441), .B1(n4440), .B2(n3050), .ZN(n3046)
         );
  OAI21_X1 U3859 ( .B1(n3120), .B2(n4443), .A(n3046), .ZN(n3047) );
  AOI21_X1 U3860 ( .B1(n3048), .B2(n4461), .A(n3047), .ZN(n4546) );
  XNOR2_X1 U3861 ( .A(n3049), .B(n3552), .ZN(n4549) );
  NAND2_X1 U3862 ( .A1(n3099), .A2(n3050), .ZN(n3051) );
  NAND2_X1 U3863 ( .A1(n3138), .A2(n3051), .ZN(n4547) );
  AOI22_X1 U3864 ( .A1(n4471), .A2(REG2_REG_9__SCAN_IN), .B1(n3123), .B2(n4466), .ZN(n3052) );
  OAI21_X1 U3865 ( .B1(n4547), .B2(n3952), .A(n3052), .ZN(n3053) );
  AOI21_X1 U3866 ( .B1(n4549), .B2(n3808), .A(n3053), .ZN(n3054) );
  OAI21_X1 U3867 ( .B1(n4546), .B2(n4471), .A(n3054), .ZN(U3281) );
  AOI22_X1 U3868 ( .A1(n3055), .A2(n3424), .B1(n3449), .B2(n3620), .ZN(n3058)
         );
  INV_X1 U3869 ( .A(n3056), .ZN(n3057) );
  OAI211_X1 U3870 ( .C1(n3120), .C2(n3387), .A(n3058), .B(n3057), .ZN(n3063)
         );
  AOI211_X1 U3871 ( .C1(n3061), .C2(n3060), .A(n3394), .B(n2247), .ZN(n3062)
         );
  AOI211_X1 U3872 ( .C1(n3450), .C2(n3064), .A(n3063), .B(n3062), .ZN(n3065)
         );
  INV_X1 U3873 ( .A(n3065), .ZN(U3210) );
  INV_X1 U3874 ( .A(REG2_REG_14__SCAN_IN), .ZN(n3076) );
  INV_X1 U3875 ( .A(n4262), .ZN(n3095) );
  INV_X1 U3876 ( .A(REG2_REG_11__SCAN_IN), .ZN(n4412) );
  AOI22_X1 U3877 ( .A1(n4494), .A2(REG2_REG_11__SCAN_IN), .B1(n4412), .B2(
        n4331), .ZN(n4328) );
  NAND2_X1 U3878 ( .A1(REG2_REG_9__SCAN_IN), .A2(n3081), .ZN(n3069) );
  INV_X1 U3879 ( .A(n3081), .ZN(n4499) );
  INV_X1 U3880 ( .A(REG2_REG_9__SCAN_IN), .ZN(n3066) );
  AOI22_X1 U3881 ( .A1(REG2_REG_9__SCAN_IN), .A2(n3081), .B1(n4499), .B2(n3066), .ZN(n4308) );
  NAND2_X1 U3882 ( .A1(n2203), .A2(n4263), .ZN(n3068) );
  NAND2_X1 U3883 ( .A1(n3068), .A2(n3653), .ZN(n4307) );
  NAND2_X1 U3884 ( .A1(n4308), .A2(n4307), .ZN(n4306) );
  NAND2_X1 U3885 ( .A1(n3069), .A2(n4306), .ZN(n3070) );
  NAND2_X1 U3886 ( .A1(n3088), .A2(n3070), .ZN(n3071) );
  INV_X1 U3887 ( .A(n3088), .ZN(n4497) );
  XNOR2_X1 U3888 ( .A(n3070), .B(n4497), .ZN(n4317) );
  NAND2_X1 U3889 ( .A1(REG2_REG_10__SCAN_IN), .A2(n4317), .ZN(n4316) );
  NAND2_X1 U3890 ( .A1(n3071), .A2(n4316), .ZN(n4327) );
  NAND2_X1 U3891 ( .A1(n3091), .A2(n3072), .ZN(n3073) );
  NAND2_X1 U3892 ( .A1(n3073), .A2(n4335), .ZN(n4348) );
  INV_X1 U3893 ( .A(n4491), .ZN(n4357) );
  INV_X1 U3894 ( .A(REG2_REG_13__SCAN_IN), .ZN(n4345) );
  NOR2_X1 U3895 ( .A1(n4357), .A2(n4345), .ZN(n4344) );
  INV_X1 U3896 ( .A(n4346), .ZN(n4387) );
  AOI211_X1 U3897 ( .C1(n3076), .C2(n3075), .A(n3668), .B(n4387), .ZN(n3079)
         );
  AND2_X1 U3898 ( .A1(REG3_REG_14__SCAN_IN), .A2(U3149), .ZN(n3221) );
  AOI21_X1 U3899 ( .B1(n4392), .B2(ADDR_REG_14__SCAN_IN), .A(n3221), .ZN(n3077) );
  OAI21_X1 U3900 ( .B1(n4399), .B2(n3095), .A(n3077), .ZN(n3078) );
  NOR2_X1 U3901 ( .A1(n3079), .A2(n3078), .ZN(n3098) );
  INV_X1 U3902 ( .A(REG1_REG_13__SCAN_IN), .ZN(n3080) );
  AOI22_X1 U3903 ( .A1(n4491), .A2(REG1_REG_13__SCAN_IN), .B1(n3080), .B2(
        n4357), .ZN(n4354) );
  INV_X1 U3904 ( .A(REG1_REG_11__SCAN_IN), .ZN(n4577) );
  AOI22_X1 U3905 ( .A1(n4494), .A2(REG1_REG_11__SCAN_IN), .B1(n4577), .B2(
        n4331), .ZN(n4325) );
  NAND2_X1 U3906 ( .A1(REG1_REG_9__SCAN_IN), .A2(n3081), .ZN(n3087) );
  INV_X1 U3907 ( .A(REG1_REG_9__SCAN_IN), .ZN(n4574) );
  AOI22_X1 U3908 ( .A1(REG1_REG_9__SCAN_IN), .A2(n3081), .B1(n4499), .B2(n4574), .ZN(n4305) );
  NAND2_X1 U3909 ( .A1(n3085), .A2(n4263), .ZN(n3086) );
  NAND2_X1 U3910 ( .A1(n3086), .A2(n3650), .ZN(n4304) );
  NAND2_X1 U3911 ( .A1(n4305), .A2(n4304), .ZN(n4303) );
  NAND2_X1 U3912 ( .A1(n3087), .A2(n4303), .ZN(n3089) );
  NAND2_X1 U3913 ( .A1(n3088), .A2(n3089), .ZN(n3090) );
  XNOR2_X1 U3914 ( .A(n3089), .B(n4497), .ZN(n4315) );
  NAND2_X1 U3915 ( .A1(REG1_REG_10__SCAN_IN), .A2(n4315), .ZN(n4314) );
  NAND2_X1 U3916 ( .A1(n3091), .A2(n3092), .ZN(n3093) );
  NAND2_X1 U3917 ( .A1(REG1_REG_12__SCAN_IN), .A2(n4341), .ZN(n4340) );
  NAND2_X1 U3918 ( .A1(n4491), .A2(REG1_REG_13__SCAN_IN), .ZN(n3094) );
  NAND2_X1 U3919 ( .A1(REG1_REG_14__SCAN_IN), .A2(n3096), .ZN(n3661) );
  OAI211_X1 U3920 ( .C1(n3096), .C2(REG1_REG_14__SCAN_IN), .A(n4394), .B(n3661), .ZN(n3097) );
  NAND2_X1 U3921 ( .A1(n3098), .A2(n3097), .ZN(U3254) );
  OAI21_X1 U3922 ( .B1(n3100), .B2(n3103), .A(n3099), .ZN(n4430) );
  INV_X1 U3923 ( .A(REG0_REG_8__SCAN_IN), .ZN(n3110) );
  INV_X1 U3924 ( .A(n4524), .ZN(n4557) );
  NAND2_X1 U3925 ( .A1(n3494), .A2(n3490), .ZN(n3549) );
  XOR2_X1 U3926 ( .A(n3549), .B(n3101), .Z(n4432) );
  XOR2_X1 U3927 ( .A(n3549), .B(n3102), .Z(n3107) );
  OAI22_X1 U3928 ( .A1(n3104), .A2(n4464), .B1(n4403), .B2(n3103), .ZN(n3105)
         );
  AOI21_X1 U3929 ( .B1(n4407), .B2(n3619), .A(n3105), .ZN(n3106) );
  OAI21_X1 U3930 ( .B1(n3107), .B2(n4409), .A(n3106), .ZN(n3108) );
  AOI21_X1 U3931 ( .B1(n4462), .B2(n4432), .A(n3108), .ZN(n4435) );
  INV_X1 U3932 ( .A(n4435), .ZN(n3109) );
  AOI21_X1 U3933 ( .B1(n4557), .B2(n4432), .A(n3109), .ZN(n3112) );
  MUX2_X1 U3934 ( .A(n3110), .B(n3112), .S(n4560), .Z(n3111) );
  OAI21_X1 U3935 ( .B1(n4430), .B2(n4251), .A(n3111), .ZN(U3483) );
  INV_X1 U3936 ( .A(REG1_REG_8__SCAN_IN), .ZN(n3113) );
  MUX2_X1 U3937 ( .A(n3113), .B(n3112), .S(n4579), .Z(n3114) );
  OAI21_X1 U3938 ( .B1(n4430), .B2(n4193), .A(n3114), .ZN(U3526) );
  AOI21_X1 U3939 ( .B1(n3118), .B2(n3117), .A(n3116), .ZN(n3126) );
  NOR2_X1 U3940 ( .A1(STATE_REG_SCAN_IN), .A2(n3119), .ZN(n4312) );
  OAI22_X1 U3941 ( .A1(n3389), .A2(n3121), .B1(n3388), .B2(n3120), .ZN(n3122)
         );
  AOI211_X1 U3942 ( .C1(n3446), .C2(n4406), .A(n4312), .B(n3122), .ZN(n3125)
         );
  NAND2_X1 U3943 ( .A1(n3450), .A2(n3123), .ZN(n3124) );
  OAI211_X1 U3944 ( .C1(n3126), .C2(n3394), .A(n3125), .B(n3124), .ZN(U3228)
         );
  XNOR2_X1 U3945 ( .A(n3401), .B(n3128), .ZN(n3563) );
  XNOR2_X1 U3946 ( .A(n3127), .B(n3563), .ZN(n3131) );
  OAI22_X1 U3947 ( .A1(n3966), .A2(n4464), .B1(n4403), .B2(n3128), .ZN(n3129)
         );
  AOI21_X1 U3948 ( .B1(n4407), .B2(n3616), .A(n3129), .ZN(n3130) );
  OAI21_X1 U3949 ( .B1(n3131), .B2(n4409), .A(n3130), .ZN(n3167) );
  INV_X1 U3950 ( .A(n3167), .ZN(n3137) );
  XNOR2_X1 U3951 ( .A(n3132), .B(n3563), .ZN(n3168) );
  NAND2_X1 U3952 ( .A1(n4416), .A2(n3286), .ZN(n3133) );
  NAND2_X1 U3953 ( .A1(n2063), .A2(n3133), .ZN(n3174) );
  AOI22_X1 U3954 ( .A1(n4471), .A2(REG2_REG_12__SCAN_IN), .B1(n3287), .B2(
        n4466), .ZN(n3134) );
  OAI21_X1 U3955 ( .B1(n3174), .B2(n3952), .A(n3134), .ZN(n3135) );
  AOI21_X1 U3956 ( .B1(n3168), .B2(n3808), .A(n3135), .ZN(n3136) );
  OAI21_X1 U3957 ( .B1(n3137), .B2(n4471), .A(n3136), .ZN(U3278) );
  INV_X1 U3958 ( .A(n3138), .ZN(n3140) );
  INV_X1 U3959 ( .A(n4418), .ZN(n3139) );
  OAI21_X1 U3960 ( .B1(n3140), .B2(n3143), .A(n3139), .ZN(n4423) );
  INV_X1 U3961 ( .A(REG1_REG_10__SCAN_IN), .ZN(n3150) );
  NAND2_X1 U3962 ( .A1(n3457), .A2(n3458), .ZN(n3550) );
  XOR2_X1 U3963 ( .A(n3550), .B(n3141), .Z(n4425) );
  XNOR2_X1 U3964 ( .A(n3142), .B(n3550), .ZN(n3147) );
  OAI22_X1 U3965 ( .A1(n3144), .A2(n4464), .B1(n4403), .B2(n3143), .ZN(n3145)
         );
  AOI21_X1 U3966 ( .B1(n4407), .B2(n3617), .A(n3145), .ZN(n3146) );
  OAI21_X1 U3967 ( .B1(n3147), .B2(n4409), .A(n3146), .ZN(n3148) );
  AOI21_X1 U3968 ( .B1(n4425), .B2(n4462), .A(n3148), .ZN(n4428) );
  INV_X1 U3969 ( .A(n4428), .ZN(n3149) );
  AOI21_X1 U3970 ( .B1(n4557), .B2(n4425), .A(n3149), .ZN(n3152) );
  MUX2_X1 U3971 ( .A(n3150), .B(n3152), .S(n4579), .Z(n3151) );
  OAI21_X1 U3972 ( .B1(n4423), .B2(n4193), .A(n3151), .ZN(U3528) );
  INV_X1 U3973 ( .A(REG0_REG_10__SCAN_IN), .ZN(n3153) );
  MUX2_X1 U3974 ( .A(n3153), .B(n3152), .S(n4560), .Z(n3154) );
  OAI21_X1 U3975 ( .B1(n4423), .B2(n4251), .A(n3154), .ZN(U3487) );
  NAND2_X1 U3976 ( .A1(n3156), .A2(n3155), .ZN(n3158) );
  NAND2_X1 U3977 ( .A1(n3465), .A2(n3157), .ZN(n3557) );
  XNOR2_X1 U3978 ( .A(n3158), .B(n3557), .ZN(n3161) );
  AOI22_X1 U3979 ( .A1(n3944), .A2(n4441), .B1(n4440), .B2(n3377), .ZN(n3159)
         );
  OAI21_X1 U3980 ( .B1(n4404), .B2(n4443), .A(n3159), .ZN(n3160) );
  AOI21_X1 U3981 ( .B1(n3161), .B2(n4461), .A(n3160), .ZN(n4201) );
  XOR2_X1 U3982 ( .A(n3557), .B(n3162), .Z(n4200) );
  NAND2_X1 U3983 ( .A1(n2063), .A2(n3377), .ZN(n3163) );
  NAND2_X1 U3984 ( .A1(n2062), .A2(n3163), .ZN(n4203) );
  AOI22_X1 U3985 ( .A1(n4471), .A2(REG2_REG_13__SCAN_IN), .B1(n3378), .B2(
        n4466), .ZN(n3164) );
  OAI21_X1 U3986 ( .B1(n4203), .B2(n3952), .A(n3164), .ZN(n3165) );
  AOI21_X1 U3987 ( .B1(n4200), .B2(n3808), .A(n3165), .ZN(n3166) );
  OAI21_X1 U3988 ( .B1(n4471), .B2(n4201), .A(n3166), .ZN(U3277) );
  INV_X1 U3989 ( .A(REG1_REG_12__SCAN_IN), .ZN(n3169) );
  AOI21_X1 U3990 ( .B1(n4550), .B2(n3168), .A(n3167), .ZN(n3171) );
  MUX2_X1 U3991 ( .A(n3169), .B(n3171), .S(n4579), .Z(n3170) );
  OAI21_X1 U3992 ( .B1(n3174), .B2(n4193), .A(n3170), .ZN(U3530) );
  INV_X1 U3993 ( .A(REG0_REG_12__SCAN_IN), .ZN(n3172) );
  MUX2_X1 U3994 ( .A(n3172), .B(n3171), .S(n4560), .Z(n3173) );
  OAI21_X1 U3995 ( .B1(n3174), .B2(n4251), .A(n3173), .ZN(U3491) );
  INV_X1 U3996 ( .A(n3175), .ZN(n3181) );
  INV_X1 U3997 ( .A(REG2_REG_28__SCAN_IN), .ZN(n3177) );
  INV_X1 U3998 ( .A(n3210), .ZN(n3176) );
  OAI22_X1 U3999 ( .A1(n3972), .A2(n3177), .B1(n3176), .B2(n4413), .ZN(n3180)
         );
  NOR2_X1 U4000 ( .A1(n3178), .A2(n4471), .ZN(n3179) );
  AOI211_X1 U4001 ( .C1(n4455), .C2(n3181), .A(n3180), .B(n3179), .ZN(n3182)
         );
  OAI21_X1 U4002 ( .B1(n3183), .B2(n3955), .A(n3182), .ZN(U3262) );
  NAND3_X1 U4003 ( .A1(n3184), .A2(STATE_REG_SCAN_IN), .A3(IR_REG_31__SCAN_IN), 
        .ZN(n3186) );
  INV_X1 U4004 ( .A(DATAI_31_), .ZN(n3185) );
  OAI22_X1 U4005 ( .A1(n2278), .A2(n3186), .B1(STATE_REG_SCAN_IN), .B2(n3185), 
        .ZN(U3321) );
  INV_X1 U4006 ( .A(n3187), .ZN(n3189) );
  NAND2_X1 U4007 ( .A1(n3716), .A2(n2671), .ZN(n3192) );
  NAND2_X1 U4008 ( .A1(n3190), .A2(n3699), .ZN(n3191) );
  NAND2_X1 U4009 ( .A1(n3192), .A2(n3191), .ZN(n3194) );
  XNOR2_X1 U4010 ( .A(n3194), .B(n3193), .ZN(n3198) );
  NAND2_X1 U4011 ( .A1(n3716), .A2(n3195), .ZN(n3196) );
  OAI21_X1 U4012 ( .B1(n3207), .B2(n2029), .A(n3196), .ZN(n3197) );
  XNOR2_X1 U4013 ( .A(n3198), .B(n3197), .ZN(n3214) );
  INV_X1 U4014 ( .A(n3214), .ZN(n3199) );
  INV_X1 U4015 ( .A(n3200), .ZN(n3201) );
  NAND2_X1 U4016 ( .A1(n3202), .A2(n3201), .ZN(n3213) );
  INV_X1 U4017 ( .A(n3213), .ZN(n3203) );
  NAND3_X1 U4018 ( .A1(n3199), .A2(n3434), .A3(n3203), .ZN(n3212) );
  INV_X1 U4019 ( .A(n3609), .ZN(n3205) );
  OAI22_X1 U4020 ( .A1(n3387), .A2(n3205), .B1(STATE_REG_SCAN_IN), .B2(n3204), 
        .ZN(n3209) );
  OAI22_X1 U4021 ( .A1(n3389), .A2(n3207), .B1(n3388), .B2(n3206), .ZN(n3208)
         );
  AOI211_X1 U4022 ( .C1(n3450), .C2(n3210), .A(n3209), .B(n3208), .ZN(n3211)
         );
  AND2_X1 U4023 ( .A1(n3212), .A2(n3211), .ZN(n3215) );
  XNOR2_X1 U4024 ( .A(n3217), .B(n3216), .ZN(n3218) );
  XNOR2_X1 U4025 ( .A(n3219), .B(n3218), .ZN(n3220) );
  NAND2_X1 U4026 ( .A1(n3220), .A2(n3434), .ZN(n3225) );
  AOI21_X1 U4027 ( .B1(n3446), .B2(n3963), .A(n3221), .ZN(n3224) );
  AOI22_X1 U4028 ( .A1(n3969), .A2(n3424), .B1(n3449), .B2(n3615), .ZN(n3223)
         );
  NAND2_X1 U4029 ( .A1(n3450), .A2(n3970), .ZN(n3222) );
  NAND4_X1 U4030 ( .A1(n3225), .A2(n3224), .A3(n3223), .A4(n3222), .ZN(U3212)
         );
  INV_X1 U4031 ( .A(n3226), .ZN(n3384) );
  OAI21_X1 U4032 ( .B1(n3384), .B2(n3228), .A(n3227), .ZN(n3230) );
  NAND3_X1 U4033 ( .A1(n3230), .A2(n3434), .A3(n3229), .ZN(n3234) );
  AOI22_X1 U4034 ( .A1(n3446), .A2(n3792), .B1(REG3_REG_23__SCAN_IN), .B2(
        U3149), .ZN(n3233) );
  AOI22_X1 U4035 ( .A1(n3830), .A2(n3449), .B1(n3448), .B2(n3791), .ZN(n3232)
         );
  NAND2_X1 U4036 ( .A1(n3450), .A2(n3799), .ZN(n3231) );
  NAND4_X1 U4037 ( .A1(n3234), .A2(n3233), .A3(n3232), .A4(n3231), .ZN(U3213)
         );
  OAI21_X1 U4038 ( .B1(n3116), .B2(n3236), .A(n3235), .ZN(n3239) );
  NAND3_X1 U4039 ( .A1(n3239), .A2(n3434), .A3(n3238), .ZN(n3244) );
  NOR2_X1 U4040 ( .A1(STATE_REG_SCAN_IN), .A2(n4059), .ZN(n4321) );
  AOI21_X1 U4041 ( .B1(n3616), .B2(n3446), .A(n4321), .ZN(n3243) );
  AOI22_X1 U4042 ( .A1(n3240), .A2(n3424), .B1(n3449), .B2(n3617), .ZN(n3242)
         );
  NAND2_X1 U40430 ( .A1(n3450), .A2(n4422), .ZN(n3241) );
  NAND4_X1 U4044 ( .A1(n3244), .A2(n3243), .A3(n3242), .A4(n3241), .ZN(U3214)
         );
  AOI21_X1 U4045 ( .B1(n3246), .B2(n3245), .A(n3346), .ZN(n3247) );
  OR2_X1 U4046 ( .A1(n3247), .A2(n3394), .ZN(n3253) );
  AOI21_X1 U4047 ( .B1(n3622), .B2(n3446), .A(n3248), .ZN(n3252) );
  AOI22_X1 U4048 ( .A1(n2751), .A2(n3449), .B1(n3448), .B2(n3474), .ZN(n3251)
         );
  NAND2_X1 U4049 ( .A1(n3450), .A2(n3249), .ZN(n3250) );
  NAND4_X1 U4050 ( .A1(n3253), .A2(n3252), .A3(n3251), .A4(n3250), .ZN(U3215)
         );
  XNOR2_X1 U4051 ( .A(n3255), .B(n3254), .ZN(n3256) );
  NAND2_X1 U4052 ( .A1(n3256), .A2(n3434), .ZN(n3262) );
  NAND2_X1 U4053 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n3680) );
  INV_X1 U4054 ( .A(n3680), .ZN(n3257) );
  AOI21_X1 U4055 ( .B1(n3446), .B2(n3613), .A(n3257), .ZN(n3261) );
  AOI22_X1 U4056 ( .A1(n3872), .A2(n3449), .B1(n3448), .B2(n3258), .ZN(n3260)
         );
  NAND2_X1 U4057 ( .A1(n3450), .A2(n3877), .ZN(n3259) );
  NAND4_X1 U4058 ( .A1(n3262), .A2(n3261), .A3(n3260), .A4(n3259), .ZN(U3216)
         );
  XNOR2_X1 U4059 ( .A(n3265), .B(n3264), .ZN(n3266) );
  XNOR2_X1 U4060 ( .A(n3263), .B(n3266), .ZN(n3267) );
  NAND2_X1 U4061 ( .A1(n3267), .A2(n3434), .ZN(n3273) );
  NAND2_X1 U4062 ( .A1(REG3_REG_8__SCAN_IN), .A2(U3149), .ZN(n3656) );
  INV_X1 U4063 ( .A(n3656), .ZN(n3268) );
  AOI21_X1 U4064 ( .B1(n3446), .B2(n3617), .A(n3268), .ZN(n3272) );
  AOI22_X1 U4065 ( .A1(n3619), .A2(n3449), .B1(n3448), .B2(n3269), .ZN(n3271)
         );
  NAND2_X1 U4066 ( .A1(n3450), .A2(n4429), .ZN(n3270) );
  NAND4_X1 U4067 ( .A1(n3273), .A2(n3272), .A3(n3271), .A4(n3270), .ZN(U3218)
         );
  XNOR2_X1 U4068 ( .A(n3275), .B(n3274), .ZN(n3276) );
  XNOR2_X1 U4069 ( .A(n2051), .B(n3276), .ZN(n3277) );
  NAND2_X1 U4070 ( .A1(n3277), .A2(n3434), .ZN(n3281) );
  AOI22_X1 U4071 ( .A1(n3830), .A2(n3446), .B1(REG3_REG_21__SCAN_IN), .B2(
        U3149), .ZN(n3280) );
  AOI22_X1 U4072 ( .A1(n3829), .A2(n3424), .B1(n3449), .B2(n3613), .ZN(n3279)
         );
  NAND2_X1 U4073 ( .A1(n3450), .A2(n3837), .ZN(n3278) );
  NAND4_X1 U4074 ( .A1(n3281), .A2(n3280), .A3(n3279), .A4(n3278), .ZN(U3220)
         );
  XNOR2_X1 U4075 ( .A(n3370), .B(n3369), .ZN(n3283) );
  XNOR2_X1 U4076 ( .A(n3282), .B(n3283), .ZN(n3284) );
  NAND2_X1 U4077 ( .A1(n3284), .A2(n3434), .ZN(n3291) );
  NAND2_X1 U4078 ( .A1(REG3_REG_12__SCAN_IN), .A2(U3149), .ZN(n4338) );
  INV_X1 U4079 ( .A(n4338), .ZN(n3285) );
  AOI21_X1 U4080 ( .B1(n3446), .B2(n3615), .A(n3285), .ZN(n3290) );
  AOI22_X1 U4081 ( .A1(n3616), .A2(n3449), .B1(n3448), .B2(n3286), .ZN(n3289)
         );
  NAND2_X1 U4082 ( .A1(n3450), .A2(n3287), .ZN(n3288) );
  NAND4_X1 U4083 ( .A1(n3291), .A2(n3290), .A3(n3289), .A4(n3288), .ZN(U3221)
         );
  INV_X1 U4084 ( .A(n3293), .ZN(n3295) );
  NAND2_X1 U4085 ( .A1(n3295), .A2(n3294), .ZN(n3296) );
  XNOR2_X1 U4086 ( .A(n3292), .B(n3296), .ZN(n3297) );
  NAND2_X1 U4087 ( .A1(n3297), .A2(n3434), .ZN(n3303) );
  NOR2_X1 U4088 ( .A1(n3298), .A2(STATE_REG_SCAN_IN), .ZN(n3299) );
  AOI21_X1 U4089 ( .B1(n3446), .B2(n3753), .A(n3299), .ZN(n3302) );
  AOI22_X1 U4090 ( .A1(n3757), .A2(n3424), .B1(n3449), .B2(n3792), .ZN(n3301)
         );
  NAND2_X1 U4091 ( .A1(n3450), .A2(n3760), .ZN(n3300) );
  NAND4_X1 U4092 ( .A1(n3303), .A2(n3302), .A3(n3301), .A4(n3300), .ZN(U3222)
         );
  INV_X1 U4093 ( .A(n3442), .ZN(n3305) );
  OAI21_X1 U4094 ( .B1(n3305), .B2(n3443), .A(n3304), .ZN(n3307) );
  XNOR2_X1 U4095 ( .A(n3307), .B(n3306), .ZN(n3308) );
  NAND2_X1 U4096 ( .A1(n3308), .A2(n3434), .ZN(n3313) );
  AND2_X1 U4097 ( .A1(REG3_REG_16__SCAN_IN), .A2(U3149), .ZN(n4371) );
  AOI21_X1 U4098 ( .B1(n3614), .B2(n3446), .A(n4371), .ZN(n3312) );
  AOI22_X1 U4099 ( .A1(n3309), .A2(n3424), .B1(n3449), .B2(n3963), .ZN(n3311)
         );
  NAND2_X1 U4100 ( .A1(n3450), .A2(n3930), .ZN(n3310) );
  NAND4_X1 U4101 ( .A1(n3313), .A2(n3312), .A3(n3311), .A4(n3310), .ZN(U3223)
         );
  XOR2_X1 U4102 ( .A(n3315), .B(n3314), .Z(n3316) );
  NAND2_X1 U4103 ( .A1(n3316), .A2(n3434), .ZN(n3322) );
  AND2_X1 U4104 ( .A1(U3149), .A2(REG3_REG_5__SCAN_IN), .ZN(n4286) );
  AOI21_X1 U4105 ( .B1(n3446), .B2(n3620), .A(n4286), .ZN(n3321) );
  AOI22_X1 U4106 ( .A1(n3622), .A2(n3449), .B1(n3448), .B2(n3317), .ZN(n3320)
         );
  NAND2_X1 U4107 ( .A1(n3450), .A2(n3318), .ZN(n3319) );
  NAND4_X1 U4108 ( .A1(n3322), .A2(n3321), .A3(n3320), .A4(n3319), .ZN(U3224)
         );
  XNOR2_X1 U4109 ( .A(n3325), .B(n3324), .ZN(n3326) );
  XNOR2_X1 U4110 ( .A(n3323), .B(n3326), .ZN(n3327) );
  NAND2_X1 U4111 ( .A1(n3327), .A2(n3434), .ZN(n3332) );
  AND2_X1 U4112 ( .A1(U3149), .A2(REG3_REG_17__SCAN_IN), .ZN(n4380) );
  AOI21_X1 U4113 ( .B1(n3872), .B2(n3446), .A(n4380), .ZN(n3331) );
  AOI22_X1 U4114 ( .A1(n3906), .A2(n3449), .B1(n3448), .B2(n3328), .ZN(n3330)
         );
  NAND2_X1 U4115 ( .A1(n3450), .A2(n3913), .ZN(n3329) );
  NAND4_X1 U4116 ( .A1(n3332), .A2(n3331), .A3(n3330), .A4(n3329), .ZN(U3225)
         );
  NAND2_X1 U4117 ( .A1(n3333), .A2(n3334), .ZN(n3336) );
  XNOR2_X1 U4118 ( .A(n3336), .B(n3335), .ZN(n3337) );
  NAND2_X1 U4119 ( .A1(n3337), .A2(n3434), .ZN(n3342) );
  AOI22_X1 U4120 ( .A1(n3610), .A2(n3446), .B1(REG3_REG_24__SCAN_IN), .B2(
        U3149), .ZN(n3341) );
  AOI22_X1 U4121 ( .A1(n3611), .A2(n3449), .B1(n3448), .B2(n3338), .ZN(n3340)
         );
  NAND2_X1 U4122 ( .A1(n3450), .A2(n3776), .ZN(n3339) );
  NAND4_X1 U4123 ( .A1(n3342), .A2(n3341), .A3(n3340), .A4(n3339), .ZN(U3226)
         );
  OAI21_X1 U4124 ( .B1(n3346), .B2(n3345), .A(n3344), .ZN(n3347) );
  NAND3_X1 U4125 ( .A1(n2110), .A2(n3434), .A3(n3347), .ZN(n3354) );
  AOI21_X1 U4126 ( .B1(n3446), .B2(n3621), .A(n3348), .ZN(n3353) );
  AOI22_X1 U4127 ( .A1(n3349), .A2(n3424), .B1(n3449), .B2(n3623), .ZN(n3352)
         );
  NAND2_X1 U4128 ( .A1(n3450), .A2(n3350), .ZN(n3351) );
  NAND4_X1 U4129 ( .A1(n3354), .A2(n3353), .A3(n3352), .A4(n3351), .ZN(U3227)
         );
  INV_X1 U4130 ( .A(n3359), .ZN(n3356) );
  NOR2_X1 U4131 ( .A1(n3355), .A2(n3356), .ZN(n3361) );
  AOI21_X1 U4132 ( .B1(n3359), .B2(n3358), .A(n3357), .ZN(n3360) );
  OAI21_X1 U4133 ( .B1(n3361), .B2(n3360), .A(n3434), .ZN(n3366) );
  INV_X1 U4134 ( .A(n3849), .ZN(n3612) );
  AOI22_X1 U4135 ( .A1(n3612), .A2(n3446), .B1(REG3_REG_20__SCAN_IN), .B2(
        U3149), .ZN(n3365) );
  AOI22_X1 U4136 ( .A1(n3362), .A2(n3424), .B1(n3449), .B2(n3887), .ZN(n3364)
         );
  NAND2_X1 U4137 ( .A1(n3450), .A2(n3856), .ZN(n3363) );
  NAND4_X1 U4138 ( .A1(n3366), .A2(n3365), .A3(n3364), .A4(n3363), .ZN(U3230)
         );
  NOR2_X1 U4139 ( .A1(n3368), .A2(n3367), .ZN(n3375) );
  INV_X1 U4140 ( .A(n3282), .ZN(n3373) );
  OAI21_X1 U4141 ( .B1(n3282), .B2(n3370), .A(n3369), .ZN(n3371) );
  OAI21_X1 U4142 ( .B1(n3373), .B2(n3372), .A(n3371), .ZN(n3374) );
  XOR2_X1 U4143 ( .A(n3375), .B(n3374), .Z(n3376) );
  NAND2_X1 U4144 ( .A1(n3376), .A2(n3434), .ZN(n3382) );
  AND2_X1 U4145 ( .A1(U3149), .A2(REG3_REG_13__SCAN_IN), .ZN(n4351) );
  AOI21_X1 U4146 ( .B1(n3944), .B2(n3446), .A(n4351), .ZN(n3381) );
  AOI22_X1 U4147 ( .A1(n3377), .A2(n3424), .B1(n3449), .B2(n3401), .ZN(n3380)
         );
  NAND2_X1 U4148 ( .A1(n3450), .A2(n3378), .ZN(n3379) );
  NAND4_X1 U4149 ( .A1(n3382), .A2(n3381), .A3(n3380), .A4(n3379), .ZN(U3231)
         );
  AOI21_X1 U4150 ( .B1(n3385), .B2(n3383), .A(n3384), .ZN(n3395) );
  INV_X1 U4151 ( .A(REG3_REG_22__SCAN_IN), .ZN(n3386) );
  OAI22_X1 U4152 ( .A1(n3387), .A2(n3816), .B1(STATE_REG_SCAN_IN), .B2(n3386), 
        .ZN(n3391) );
  OAI22_X1 U4153 ( .A1(n3389), .A2(n3820), .B1(n3388), .B2(n3849), .ZN(n3390)
         );
  AOI211_X1 U4154 ( .C1(n3392), .C2(n3450), .A(n3391), .B(n3390), .ZN(n3393)
         );
  OAI21_X1 U4155 ( .B1(n3395), .B2(n3394), .A(n3393), .ZN(U3232) );
  NAND2_X1 U4156 ( .A1(n3398), .A2(n3397), .ZN(n3399) );
  XNOR2_X1 U4157 ( .A(n3396), .B(n3399), .ZN(n3400) );
  NAND2_X1 U4158 ( .A1(n3400), .A2(n3434), .ZN(n3407) );
  AND2_X1 U4159 ( .A1(U3149), .A2(REG3_REG_11__SCAN_IN), .ZN(n4333) );
  AOI21_X1 U4160 ( .B1(n3446), .B2(n3401), .A(n4333), .ZN(n3406) );
  AOI22_X1 U4161 ( .A1(n3402), .A2(n3424), .B1(n3449), .B2(n4406), .ZN(n3405)
         );
  NAND2_X1 U4162 ( .A1(n3450), .A2(n3403), .ZN(n3404) );
  NAND4_X1 U4163 ( .A1(n3407), .A2(n3406), .A3(n3405), .A4(n3404), .ZN(U3233)
         );
  NAND2_X1 U4164 ( .A1(n2109), .A2(n3409), .ZN(n3410) );
  XNOR2_X1 U4165 ( .A(n3411), .B(n3410), .ZN(n3412) );
  NAND2_X1 U4166 ( .A1(n3412), .A2(n3434), .ZN(n3417) );
  INV_X1 U4167 ( .A(REG3_REG_18__SCAN_IN), .ZN(n3413) );
  NOR2_X1 U4168 ( .A1(STATE_REG_SCAN_IN), .A2(n3413), .ZN(n4391) );
  AOI21_X1 U4169 ( .B1(n3446), .B2(n3887), .A(n4391), .ZN(n3416) );
  AOI22_X1 U4170 ( .A1(n3614), .A2(n3449), .B1(n3448), .B2(n3886), .ZN(n3415)
         );
  NAND2_X1 U4171 ( .A1(n3450), .A2(n3895), .ZN(n3414) );
  NAND4_X1 U4172 ( .A1(n3417), .A2(n3416), .A3(n3415), .A4(n3414), .ZN(U3235)
         );
  INV_X1 U4173 ( .A(n3419), .ZN(n3421) );
  NAND2_X1 U4174 ( .A1(n3421), .A2(n3420), .ZN(n3422) );
  XNOR2_X1 U4175 ( .A(n3418), .B(n3422), .ZN(n3423) );
  NAND2_X1 U4176 ( .A1(n3423), .A2(n3434), .ZN(n3430) );
  INV_X1 U4177 ( .A(REG3_REG_6__SCAN_IN), .ZN(n4054) );
  NOR2_X1 U4178 ( .A1(STATE_REG_SCAN_IN), .A2(n4054), .ZN(n4298) );
  AOI21_X1 U4179 ( .B1(n3619), .B2(n3446), .A(n4298), .ZN(n3429) );
  AOI22_X1 U4180 ( .A1(n3425), .A2(n3424), .B1(n3449), .B2(n3621), .ZN(n3428)
         );
  NAND2_X1 U4181 ( .A1(n3450), .A2(n3426), .ZN(n3427) );
  NAND4_X1 U4182 ( .A1(n3430), .A2(n3429), .A3(n3428), .A4(n3427), .ZN(U3236)
         );
  NOR2_X1 U4183 ( .A1(n3436), .A2(STATE_REG_SCAN_IN), .ZN(n3437) );
  AOI21_X1 U4184 ( .B1(n3446), .B2(n3742), .A(n3437), .ZN(n3440) );
  AOI22_X1 U4185 ( .A1(n3610), .A2(n3449), .B1(n3448), .B2(n3741), .ZN(n3439)
         );
  NAND2_X1 U4186 ( .A1(n3450), .A2(n3732), .ZN(n3438) );
  NAND4_X1 U4187 ( .A1(n3441), .A2(n3440), .A3(n3439), .A4(n3438), .ZN(U3237)
         );
  NAND2_X1 U4188 ( .A1(n3442), .A2(n3304), .ZN(n3444) );
  XNOR2_X1 U4189 ( .A(n3444), .B(n3443), .ZN(n3445) );
  NAND2_X1 U4190 ( .A1(n3445), .A2(n3434), .ZN(n3454) );
  AND2_X1 U4191 ( .A1(REG3_REG_15__SCAN_IN), .A2(U3149), .ZN(n4362) );
  AOI21_X1 U4192 ( .B1(n3906), .B2(n3446), .A(n4362), .ZN(n3453) );
  AOI22_X1 U4193 ( .A1(n3944), .A2(n3449), .B1(n3448), .B2(n3447), .ZN(n3452)
         );
  NAND2_X1 U4194 ( .A1(n3450), .A2(n3950), .ZN(n3451) );
  NAND4_X1 U4195 ( .A1(n3454), .A2(n3453), .A3(n3452), .A4(n3451), .ZN(U3238)
         );
  INV_X1 U4196 ( .A(n3464), .ZN(n3573) );
  AND2_X1 U4197 ( .A1(n3456), .A2(n3455), .ZN(n3492) );
  NOR2_X1 U4198 ( .A1(n3573), .A2(n3492), .ZN(n3576) );
  AND2_X1 U4199 ( .A1(n3459), .A2(n3458), .ZN(n3460) );
  AND2_X1 U4200 ( .A1(n3462), .A2(n3460), .ZN(n3497) );
  OAI21_X1 U4201 ( .B1(n2072), .B2(n3463), .A(n3462), .ZN(n3466) );
  NAND4_X1 U4202 ( .A1(n3466), .A2(n3939), .A3(n3465), .A4(n3464), .ZN(n3467)
         );
  AOI21_X1 U4203 ( .B1(n2077), .B2(n3497), .A(n3467), .ZN(n3501) );
  INV_X1 U4204 ( .A(n3534), .ZN(n4437) );
  NAND2_X1 U4205 ( .A1(n3625), .A2(n4460), .ZN(n3533) );
  OAI211_X1 U4206 ( .C1(n4437), .C2(n4259), .A(n3533), .B(n3468), .ZN(n3470)
         );
  NAND3_X1 U4207 ( .A1(n3470), .A2(n3469), .A3(n2793), .ZN(n3472) );
  OAI211_X1 U4208 ( .C1(n3474), .C2(n3473), .A(n3472), .B(n3471), .ZN(n3477)
         );
  NAND3_X1 U4209 ( .A1(n3477), .A2(n3476), .A3(n3475), .ZN(n3480) );
  NAND4_X1 U4210 ( .A1(n3480), .A2(n3479), .A3(n3478), .A4(n3484), .ZN(n3483)
         );
  INV_X1 U4211 ( .A(n3531), .ZN(n3482) );
  NAND3_X1 U4212 ( .A1(n3483), .A2(n3482), .A3(n3481), .ZN(n3488) );
  INV_X1 U4213 ( .A(n3484), .ZN(n3486) );
  NOR3_X1 U4214 ( .A1(n3576), .A2(n3486), .A3(n3485), .ZN(n3487) );
  AOI21_X1 U4215 ( .B1(n3488), .B2(n3492), .A(n3487), .ZN(n3491) );
  NOR3_X1 U4216 ( .A1(n3491), .A2(n2082), .A3(n2079), .ZN(n3499) );
  INV_X1 U4217 ( .A(n3492), .ZN(n3493) );
  AOI21_X1 U4218 ( .B1(n3495), .B2(n3494), .A(n3493), .ZN(n3498) );
  OAI211_X1 U4219 ( .C1(n3499), .C2(n3498), .A(n3497), .B(n3496), .ZN(n3500)
         );
  OAI21_X1 U4220 ( .B1(n3576), .B2(n3501), .A(n3500), .ZN(n3502) );
  NAND2_X1 U4221 ( .A1(n3579), .A2(n3502), .ZN(n3503) );
  AOI211_X1 U4222 ( .C1(n3575), .C2(n3503), .A(n3585), .B(n3578), .ZN(n3505)
         );
  NOR2_X1 U4223 ( .A1(n3505), .A2(n3504), .ZN(n3506) );
  OAI21_X1 U4224 ( .B1(n3786), .B2(n3506), .A(n3582), .ZN(n3507) );
  AOI211_X1 U4225 ( .C1(n3508), .C2(n3507), .A(n3588), .B(n3571), .ZN(n3512)
         );
  NAND2_X1 U4226 ( .A1(n2352), .A2(DATAI_29_), .ZN(n3705) );
  AND2_X1 U4227 ( .A1(n3609), .A2(n3705), .ZN(n3509) );
  NOR2_X1 U4228 ( .A1(n3686), .A2(n3509), .ZN(n3569) );
  INV_X1 U4229 ( .A(n3569), .ZN(n3510) );
  OR4_X1 U4230 ( .A1(n3513), .A2(n3512), .A3(n3511), .A4(n3510), .ZN(n3527) );
  OR2_X1 U4231 ( .A1(n3687), .A2(n3572), .ZN(n3523) );
  NAND2_X1 U4232 ( .A1(n3514), .A2(REG1_REG_30__SCAN_IN), .ZN(n3517) );
  NAND2_X1 U4233 ( .A1(n3518), .A2(REG2_REG_30__SCAN_IN), .ZN(n3516) );
  NAND2_X1 U4234 ( .A1(n2332), .A2(REG0_REG_30__SCAN_IN), .ZN(n3515) );
  NAND3_X1 U4235 ( .A1(n3517), .A2(n3516), .A3(n3515), .ZN(n3692) );
  INV_X1 U4236 ( .A(n3984), .ZN(n3987) );
  NAND2_X1 U4237 ( .A1(n3514), .A2(REG1_REG_31__SCAN_IN), .ZN(n3521) );
  NAND2_X1 U4238 ( .A1(n3518), .A2(REG2_REG_31__SCAN_IN), .ZN(n3520) );
  NAND2_X1 U4239 ( .A1(n2398), .A2(REG0_REG_31__SCAN_IN), .ZN(n3519) );
  NAND3_X1 U4240 ( .A1(n3521), .A2(n3520), .A3(n3519), .ZN(n3977) );
  NAND2_X1 U4241 ( .A1(n2352), .A2(DATAI_31_), .ZN(n3567) );
  NAND2_X1 U4242 ( .A1(n3977), .A2(n3567), .ZN(n3525) );
  OAI21_X1 U4243 ( .B1(n3692), .B2(n3987), .A(n3525), .ZN(n3547) );
  INV_X1 U4244 ( .A(n3547), .ZN(n3522) );
  OAI21_X1 U4245 ( .B1(n3609), .B2(n3705), .A(n3522), .ZN(n3570) );
  AOI21_X1 U4246 ( .B1(n3523), .B2(n3569), .A(n3570), .ZN(n3592) );
  NOR2_X1 U4247 ( .A1(n3977), .A2(n3567), .ZN(n3596) );
  INV_X1 U4248 ( .A(n3692), .ZN(n3524) );
  NOR2_X1 U4249 ( .A1(n3524), .A2(n3984), .ZN(n3597) );
  NOR2_X1 U4250 ( .A1(n3596), .A2(n3597), .ZN(n3545) );
  INV_X1 U4251 ( .A(n3545), .ZN(n3526) );
  AOI22_X1 U4252 ( .A1(n3527), .A2(n3592), .B1(n3526), .B2(n3525), .ZN(n3601)
         );
  INV_X1 U4253 ( .A(n3814), .ZN(n3529) );
  NOR4_X1 U4254 ( .A1(n3530), .A2(n3529), .A3(n3957), .A4(n3528), .ZN(n3539)
         );
  XNOR2_X1 U4255 ( .A(n3609), .B(n3705), .ZN(n3702) );
  INV_X1 U4256 ( .A(n3702), .ZN(n3538) );
  NOR4_X1 U4257 ( .A1(n3885), .A2(n4401), .A3(n3532), .A4(n3531), .ZN(n3537)
         );
  NAND2_X1 U4258 ( .A1(n3534), .A2(n3533), .ZN(n4508) );
  NAND2_X1 U4259 ( .A1(n3535), .A2(n3568), .ZN(n3740) );
  NOR4_X1 U4260 ( .A1(n4447), .A2(n3940), .A3(n4508), .A4(n3740), .ZN(n3536)
         );
  NAND4_X1 U4261 ( .A1(n3539), .A2(n3538), .A3(n3537), .A4(n3536), .ZN(n3566)
         );
  INV_X1 U4262 ( .A(n3540), .ZN(n3542) );
  NOR2_X1 U4263 ( .A1(n3542), .A2(n3541), .ZN(n3847) );
  INV_X1 U4264 ( .A(n3785), .ZN(n3543) );
  OR2_X1 U4265 ( .A1(n3786), .A2(n3543), .ZN(n3826) );
  XNOR2_X1 U4266 ( .A(n3887), .B(n3876), .ZN(n3869) );
  NAND2_X1 U4267 ( .A1(n3862), .A2(n3863), .ZN(n3903) );
  NOR4_X1 U4268 ( .A1(n3847), .A2(n3826), .A3(n3869), .A4(n3903), .ZN(n3544)
         );
  NAND2_X1 U4269 ( .A1(n3545), .A2(n3544), .ZN(n3546) );
  NOR3_X1 U4270 ( .A1(n3548), .A2(n3547), .A3(n3546), .ZN(n3562) );
  NOR4_X1 U4271 ( .A1(n3552), .A2(n3551), .A3(n3550), .A4(n3549), .ZN(n3561)
         );
  INV_X1 U4272 ( .A(n3553), .ZN(n3765) );
  NAND2_X1 U4273 ( .A1(n3555), .A2(n3737), .ZN(n3750) );
  NAND2_X1 U4274 ( .A1(n3556), .A2(n3748), .ZN(n3772) );
  NOR4_X1 U4275 ( .A1(n3789), .A2(n3750), .A3(n3557), .A4(n3772), .ZN(n3560)
         );
  NOR2_X1 U4276 ( .A1(n3700), .A2(n3558), .ZN(n3559) );
  NAND4_X1 U4277 ( .A1(n3562), .A2(n3561), .A3(n3560), .A4(n3559), .ZN(n3565)
         );
  NOR4_X1 U4278 ( .A1(n3566), .A2(n3565), .A3(n3564), .A4(n3563), .ZN(n3599)
         );
  INV_X1 U4279 ( .A(n3977), .ZN(n3594) );
  NAND3_X1 U4280 ( .A1(n3713), .A2(n3569), .A3(n3568), .ZN(n3591) );
  NOR4_X1 U4281 ( .A1(n3687), .A2(n3572), .A3(n3571), .A4(n3570), .ZN(n3590)
         );
  NOR3_X1 U4282 ( .A1(n3960), .A2(n3574), .A3(n3573), .ZN(n3577) );
  OAI21_X1 U4283 ( .B1(n3577), .B2(n3576), .A(n3575), .ZN(n3581) );
  INV_X1 U4284 ( .A(n3578), .ZN(n3580) );
  NAND3_X1 U4285 ( .A1(n3581), .A2(n3580), .A3(n3579), .ZN(n3583) );
  OAI221_X1 U4286 ( .B1(n3585), .B2(n3584), .C1(n3585), .C2(n3583), .A(n3582), 
        .ZN(n3586) );
  OAI221_X1 U4287 ( .B1(n3588), .B2(n3587), .C1(n3588), .C2(n3586), .A(n3736), 
        .ZN(n3589) );
  AOI22_X1 U4288 ( .A1(n3592), .A2(n3591), .B1(n3590), .B2(n3589), .ZN(n3593)
         );
  AOI21_X1 U4289 ( .B1(n3984), .B2(n3594), .A(n3593), .ZN(n3595) );
  AOI211_X1 U4290 ( .C1(n3978), .C2(n3597), .A(n3596), .B(n3595), .ZN(n3598)
         );
  MUX2_X1 U4291 ( .A(n3599), .B(n3598), .S(n4259), .Z(n3600) );
  MUX2_X1 U4292 ( .A(n3601), .B(n3600), .S(n4260), .Z(n3602) );
  XNOR2_X1 U4293 ( .A(n3602), .B(n4261), .ZN(n3608) );
  NAND2_X1 U4294 ( .A1(n3604), .A2(n3603), .ZN(n3605) );
  OAI211_X1 U4295 ( .C1(n4258), .C2(n3607), .A(n3605), .B(B_REG_SCAN_IN), .ZN(
        n3606) );
  OAI21_X1 U4296 ( .B1(n3608), .B2(n3607), .A(n3606), .ZN(U3239) );
  MUX2_X1 U4297 ( .A(n3977), .B(DATAO_REG_31__SCAN_IN), .S(n3624), .Z(U3581)
         );
  MUX2_X1 U4298 ( .A(n3692), .B(DATAO_REG_30__SCAN_IN), .S(n3624), .Z(U3580)
         );
  MUX2_X1 U4299 ( .A(n3609), .B(DATAO_REG_29__SCAN_IN), .S(n3624), .Z(U3579)
         );
  MUX2_X1 U4300 ( .A(n3716), .B(DATAO_REG_28__SCAN_IN), .S(n3624), .Z(U3578)
         );
  MUX2_X1 U4301 ( .A(n3742), .B(DATAO_REG_27__SCAN_IN), .S(n3624), .Z(U3577)
         );
  MUX2_X1 U4302 ( .A(n3753), .B(DATAO_REG_26__SCAN_IN), .S(n3624), .Z(U3576)
         );
  MUX2_X1 U4303 ( .A(DATAO_REG_25__SCAN_IN), .B(n3610), .S(U4043), .Z(U3575)
         );
  MUX2_X1 U4304 ( .A(n3792), .B(DATAO_REG_24__SCAN_IN), .S(n3624), .Z(U3574)
         );
  MUX2_X1 U4305 ( .A(DATAO_REG_23__SCAN_IN), .B(n3611), .S(U4043), .Z(U3573)
         );
  MUX2_X1 U4306 ( .A(DATAO_REG_22__SCAN_IN), .B(n3830), .S(U4043), .Z(U3572)
         );
  MUX2_X1 U4307 ( .A(DATAO_REG_21__SCAN_IN), .B(n3612), .S(U4043), .Z(U3571)
         );
  MUX2_X1 U4308 ( .A(n3613), .B(DATAO_REG_20__SCAN_IN), .S(n3624), .Z(U3570)
         );
  MUX2_X1 U4309 ( .A(n3887), .B(DATAO_REG_19__SCAN_IN), .S(n3624), .Z(U3569)
         );
  MUX2_X1 U4310 ( .A(DATAO_REG_18__SCAN_IN), .B(n3872), .S(U4043), .Z(U3568)
         );
  MUX2_X1 U4311 ( .A(DATAO_REG_17__SCAN_IN), .B(n3614), .S(U4043), .Z(U3567)
         );
  MUX2_X1 U4312 ( .A(DATAO_REG_16__SCAN_IN), .B(n3906), .S(U4043), .Z(U3566)
         );
  MUX2_X1 U4313 ( .A(n3963), .B(DATAO_REG_15__SCAN_IN), .S(n3624), .Z(U3565)
         );
  MUX2_X1 U4314 ( .A(DATAO_REG_14__SCAN_IN), .B(n3944), .S(U4043), .Z(U3564)
         );
  MUX2_X1 U4315 ( .A(n3615), .B(DATAO_REG_13__SCAN_IN), .S(n3624), .Z(U3563)
         );
  MUX2_X1 U4316 ( .A(DATAO_REG_11__SCAN_IN), .B(n3616), .S(U4043), .Z(U3561)
         );
  MUX2_X1 U4317 ( .A(n4406), .B(DATAO_REG_10__SCAN_IN), .S(n3624), .Z(U3560)
         );
  MUX2_X1 U4318 ( .A(n3617), .B(DATAO_REG_9__SCAN_IN), .S(n3624), .Z(U3559) );
  MUX2_X1 U4319 ( .A(n3618), .B(DATAO_REG_8__SCAN_IN), .S(n3624), .Z(U3558) );
  MUX2_X1 U4320 ( .A(DATAO_REG_7__SCAN_IN), .B(n3619), .S(U4043), .Z(U3557) );
  MUX2_X1 U4321 ( .A(n3620), .B(DATAO_REG_6__SCAN_IN), .S(n3624), .Z(U3556) );
  MUX2_X1 U4322 ( .A(n3621), .B(DATAO_REG_5__SCAN_IN), .S(n3624), .Z(U3555) );
  MUX2_X1 U4323 ( .A(DATAO_REG_4__SCAN_IN), .B(n3622), .S(U4043), .Z(U3554) );
  MUX2_X1 U4324 ( .A(n3623), .B(DATAO_REG_3__SCAN_IN), .S(n3624), .Z(U3553) );
  MUX2_X1 U4325 ( .A(DATAO_REG_2__SCAN_IN), .B(n2751), .S(U4043), .Z(U3552) );
  MUX2_X1 U4326 ( .A(DATAO_REG_1__SCAN_IN), .B(n2748), .S(U4043), .Z(U3551) );
  MUX2_X1 U4327 ( .A(n3625), .B(DATAO_REG_0__SCAN_IN), .S(n3624), .Z(U3550) );
  OAI211_X1 U4328 ( .C1(n3627), .C2(n3626), .A(n4346), .B(n3641), .ZN(n3634)
         );
  OAI211_X1 U4329 ( .C1(n3630), .C2(n3629), .A(n4394), .B(n3628), .ZN(n3633)
         );
  AOI22_X1 U4330 ( .A1(n4392), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n3632) );
  INV_X1 U4331 ( .A(n4399), .ZN(n3652) );
  NAND2_X1 U4332 ( .A1(n3652), .A2(n4268), .ZN(n3631) );
  NAND4_X1 U4333 ( .A1(n3634), .A2(n3633), .A3(n3632), .A4(n3631), .ZN(U3241)
         );
  AOI22_X1 U4334 ( .A1(n4392), .A2(ADDR_REG_2__SCAN_IN), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n3635) );
  OAI21_X1 U4335 ( .B1(n3636), .B2(n4399), .A(n3635), .ZN(n3637) );
  INV_X1 U4336 ( .A(n3637), .ZN(n3648) );
  OAI211_X1 U4337 ( .C1(n3640), .C2(n3639), .A(n4394), .B(n3638), .ZN(n3647)
         );
  MUX2_X1 U4338 ( .A(n4105), .B(REG2_REG_2__SCAN_IN), .S(n4267), .Z(n3643) );
  NAND3_X1 U4339 ( .A1(n3643), .A2(n3642), .A3(n3641), .ZN(n3644) );
  NAND3_X1 U4340 ( .A1(n4346), .A2(n3645), .A3(n3644), .ZN(n3646) );
  NAND4_X1 U4341 ( .A1(n3649), .A2(n3648), .A3(n3647), .A4(n3646), .ZN(U3242)
         );
  OAI211_X1 U4342 ( .C1(n3651), .C2(REG1_REG_8__SCAN_IN), .A(n4394), .B(n3650), 
        .ZN(n3659) );
  AOI22_X1 U4343 ( .A1(n3652), .A2(n4263), .B1(n4392), .B2(ADDR_REG_8__SCAN_IN), .ZN(n3658) );
  OAI211_X1 U4344 ( .C1(REG2_REG_8__SCAN_IN), .C2(n3654), .A(n4346), .B(n3653), 
        .ZN(n3655) );
  AND2_X1 U4345 ( .A1(n3656), .A2(n3655), .ZN(n3657) );
  NAND3_X1 U4346 ( .A1(n3659), .A2(n3658), .A3(n3657), .ZN(U3248) );
  INV_X1 U4347 ( .A(REG1_REG_18__SCAN_IN), .ZN(n4080) );
  INV_X1 U4348 ( .A(n3675), .ZN(n4484) );
  AOI22_X1 U4349 ( .A1(n3675), .A2(REG1_REG_18__SCAN_IN), .B1(n4080), .B2(
        n4484), .ZN(n4396) );
  INV_X1 U4350 ( .A(REG1_REG_17__SCAN_IN), .ZN(n4183) );
  INV_X1 U4351 ( .A(n4485), .ZN(n4386) );
  INV_X1 U4352 ( .A(REG1_REG_15__SCAN_IN), .ZN(n4191) );
  AOI22_X1 U4353 ( .A1(REG1_REG_15__SCAN_IN), .A2(n3671), .B1(n4490), .B2(
        n4191), .ZN(n4365) );
  NAND2_X1 U4354 ( .A1(n3660), .A2(n4262), .ZN(n3662) );
  NAND2_X1 U4355 ( .A1(n3662), .A2(n3661), .ZN(n4364) );
  NAND2_X1 U4356 ( .A1(n4365), .A2(n4364), .ZN(n4363) );
  NOR2_X1 U4357 ( .A1(n3672), .A2(n3663), .ZN(n3664) );
  AOI22_X1 U4358 ( .A1(REG1_REG_17__SCAN_IN), .A2(n4386), .B1(n4485), .B2(
        n4183), .ZN(n4381) );
  NOR2_X1 U4359 ( .A1(n4382), .A2(n4381), .ZN(n4383) );
  AOI21_X1 U4360 ( .B1(n4183), .B2(n4386), .A(n4383), .ZN(n4395) );
  NAND2_X1 U4361 ( .A1(n4396), .A2(n4395), .ZN(n4393) );
  OAI21_X1 U4362 ( .B1(n4080), .B2(n4484), .A(n4393), .ZN(n3666) );
  XNOR2_X1 U4363 ( .A(n3681), .B(REG1_REG_19__SCAN_IN), .ZN(n3665) );
  XNOR2_X1 U4364 ( .A(n3666), .B(n3665), .ZN(n3685) );
  INV_X1 U4365 ( .A(REG2_REG_18__SCAN_IN), .ZN(n3667) );
  AOI22_X1 U4366 ( .A1(n3675), .A2(n3667), .B1(REG2_REG_18__SCAN_IN), .B2(
        n4484), .ZN(n4389) );
  INV_X1 U4367 ( .A(REG2_REG_17__SCAN_IN), .ZN(n3915) );
  AOI22_X1 U4368 ( .A1(REG2_REG_17__SCAN_IN), .A2(n4485), .B1(n4386), .B2(
        n3915), .ZN(n4378) );
  NAND2_X1 U4369 ( .A1(REG2_REG_15__SCAN_IN), .A2(n3671), .ZN(n3670) );
  OAI21_X1 U4370 ( .B1(REG2_REG_15__SCAN_IN), .B2(n3671), .A(n3670), .ZN(n4359) );
  NOR2_X1 U4371 ( .A1(n4360), .A2(n4359), .ZN(n4358) );
  INV_X1 U4372 ( .A(n3672), .ZN(n4488) );
  NAND2_X1 U4373 ( .A1(n3673), .A2(n4488), .ZN(n3674) );
  XOR2_X1 U4374 ( .A(n4488), .B(n3673), .Z(n4369) );
  NAND2_X1 U4375 ( .A1(n4369), .A2(n3932), .ZN(n4368) );
  NAND2_X1 U4376 ( .A1(n3674), .A2(n4368), .ZN(n4376) );
  INV_X1 U4377 ( .A(REG2_REG_19__SCAN_IN), .ZN(n3676) );
  MUX2_X1 U4378 ( .A(n3676), .B(REG2_REG_19__SCAN_IN), .S(n3681), .Z(n3677) );
  XNOR2_X1 U4379 ( .A(n3678), .B(n3677), .ZN(n3683) );
  NAND2_X1 U4380 ( .A1(n4392), .A2(ADDR_REG_19__SCAN_IN), .ZN(n3679) );
  OAI211_X1 U4381 ( .C1(n4399), .C2(n3681), .A(n3680), .B(n3679), .ZN(n3682)
         );
  AOI21_X1 U4382 ( .B1(n3683), .B2(n4346), .A(n3682), .ZN(n3684) );
  OAI21_X1 U4383 ( .B1(n3685), .B2(n4293), .A(n3684), .ZN(U3259) );
  INV_X1 U4384 ( .A(n3686), .ZN(n3688) );
  AOI21_X1 U4385 ( .B1(n3689), .B2(n3688), .A(n3687), .ZN(n3690) );
  XNOR2_X1 U4386 ( .A(n3690), .B(n3702), .ZN(n3696) );
  NAND2_X1 U4387 ( .A1(n3716), .A2(n4407), .ZN(n3694) );
  AND2_X1 U4388 ( .A1(n4277), .A2(B_REG_SCAN_IN), .ZN(n3691) );
  NOR2_X1 U4389 ( .A1(n4464), .A2(n3691), .ZN(n3976) );
  NAND2_X1 U4390 ( .A1(n3692), .A2(n3976), .ZN(n3693) );
  OAI211_X1 U4391 ( .C1(n3705), .C2(n4403), .A(n3694), .B(n3693), .ZN(n3695)
         );
  AOI21_X1 U4392 ( .B1(n3696), .B2(n4461), .A(n3695), .ZN(n3993) );
  INV_X1 U4393 ( .A(n3993), .ZN(n3697) );
  AOI21_X1 U4394 ( .B1(n3698), .B2(n4466), .A(n3697), .ZN(n3710) );
  NAND2_X1 U4395 ( .A1(n3991), .A2(n3808), .ZN(n3709) );
  INV_X1 U4396 ( .A(n3704), .ZN(n3706) );
  INV_X1 U4397 ( .A(n3705), .ZN(n3703) );
  OR2_X2 U4398 ( .A1(n3704), .A2(n3703), .ZN(n3983) );
  INV_X1 U4399 ( .A(n3992), .ZN(n3707) );
  AOI22_X1 U4400 ( .A1(n3707), .A2(n4455), .B1(REG2_REG_29__SCAN_IN), .B2(
        n4471), .ZN(n3708) );
  OAI211_X1 U4401 ( .C1(n4471), .C2(n3710), .A(n3709), .B(n3708), .ZN(U3354)
         );
  XNOR2_X1 U4402 ( .A(n3711), .B(n3713), .ZN(n3997) );
  OAI21_X1 U4403 ( .B1(n3714), .B2(n3713), .A(n3712), .ZN(n3715) );
  NAND2_X1 U4404 ( .A1(n3715), .A2(n4461), .ZN(n3718) );
  AOI22_X1 U4405 ( .A1(n3716), .A2(n4441), .B1(n3722), .B2(n4440), .ZN(n3717)
         );
  OAI211_X1 U4406 ( .C1(n3719), .C2(n4443), .A(n3718), .B(n3717), .ZN(n3994)
         );
  INV_X1 U4407 ( .A(n3730), .ZN(n3721) );
  AOI21_X1 U4408 ( .B1(n3722), .B2(n3721), .A(n3720), .ZN(n3995) );
  INV_X1 U4409 ( .A(n3995), .ZN(n3725) );
  AOI22_X1 U4410 ( .A1(n4471), .A2(REG2_REG_27__SCAN_IN), .B1(n3723), .B2(
        n4466), .ZN(n3724) );
  OAI21_X1 U4411 ( .B1(n3725), .B2(n3952), .A(n3724), .ZN(n3726) );
  AOI21_X1 U4412 ( .B1(n3994), .B2(n3972), .A(n3726), .ZN(n3727) );
  OAI21_X1 U4413 ( .B1(n3997), .B2(n3955), .A(n3727), .ZN(U3263) );
  INV_X1 U4414 ( .A(n3728), .ZN(n3729) );
  XOR2_X1 U4415 ( .A(n3740), .B(n3729), .Z(n4144) );
  INV_X1 U4416 ( .A(n3758), .ZN(n3731) );
  AOI21_X1 U4417 ( .B1(n3741), .B2(n3731), .A(n3730), .ZN(n4142) );
  INV_X1 U4418 ( .A(REG2_REG_26__SCAN_IN), .ZN(n3734) );
  INV_X1 U4419 ( .A(n3732), .ZN(n3733) );
  OAI22_X1 U4420 ( .A1(n3972), .A2(n3734), .B1(n3733), .B2(n4413), .ZN(n3735)
         );
  AOI21_X1 U4421 ( .B1(n4142), .B2(n4455), .A(n3735), .ZN(n3745) );
  INV_X1 U4422 ( .A(n3736), .ZN(n3738) );
  OAI21_X1 U4423 ( .B1(n3747), .B2(n3738), .A(n3737), .ZN(n3739) );
  AOI22_X1 U4424 ( .A1(n3742), .A2(n4441), .B1(n4440), .B2(n3741), .ZN(n3743)
         );
  NAND2_X1 U4425 ( .A1(n4141), .A2(n3972), .ZN(n3744) );
  OAI211_X1 U4426 ( .C1(n4144), .C2(n3955), .A(n3745), .B(n3744), .ZN(U3264)
         );
  XOR2_X1 U4427 ( .A(n3750), .B(n3746), .Z(n4148) );
  INV_X1 U4428 ( .A(n4148), .ZN(n3764) );
  INV_X1 U4429 ( .A(n3747), .ZN(n3749) );
  NAND2_X1 U4430 ( .A1(n3749), .A2(n3748), .ZN(n3751) );
  XNOR2_X1 U4431 ( .A(n3751), .B(n3750), .ZN(n3752) );
  NAND2_X1 U4432 ( .A1(n3752), .A2(n4461), .ZN(n3755) );
  AOI22_X1 U4433 ( .A1(n3753), .A2(n4441), .B1(n4440), .B2(n3757), .ZN(n3754)
         );
  OAI211_X1 U4434 ( .C1(n3756), .C2(n4443), .A(n3755), .B(n3754), .ZN(n4147)
         );
  AND2_X1 U4435 ( .A1(n2057), .A2(n3757), .ZN(n3759) );
  OR2_X1 U4436 ( .A1(n3759), .A2(n3758), .ZN(n4217) );
  AOI22_X1 U4437 ( .A1(n4471), .A2(REG2_REG_25__SCAN_IN), .B1(n3760), .B2(
        n4466), .ZN(n3761) );
  OAI21_X1 U4438 ( .B1(n4217), .B2(n3952), .A(n3761), .ZN(n3762) );
  AOI21_X1 U4439 ( .B1(n4147), .B2(n3972), .A(n3762), .ZN(n3763) );
  OAI21_X1 U4440 ( .B1(n3764), .B2(n3955), .A(n3763), .ZN(U3265) );
  NOR2_X1 U4441 ( .A1(n3766), .A2(n3765), .ZN(n3767) );
  XNOR2_X1 U4442 ( .A(n3767), .B(n3772), .ZN(n3771) );
  NOR2_X1 U4443 ( .A1(n3816), .A2(n4443), .ZN(n3770) );
  OAI22_X1 U4444 ( .A1(n3768), .A2(n4464), .B1(n4403), .B2(n3774), .ZN(n3769)
         );
  AOI211_X1 U4445 ( .C1(n3771), .C2(n4461), .A(n3770), .B(n3769), .ZN(n4151)
         );
  XNOR2_X1 U4446 ( .A(n3773), .B(n3772), .ZN(n4153) );
  NAND2_X1 U4447 ( .A1(n4153), .A2(n3808), .ZN(n3782) );
  INV_X1 U4448 ( .A(n3797), .ZN(n3775) );
  OAI21_X1 U4449 ( .B1(n3775), .B2(n3774), .A(n2057), .ZN(n4221) );
  INV_X1 U4450 ( .A(n4221), .ZN(n3780) );
  INV_X1 U4451 ( .A(REG2_REG_24__SCAN_IN), .ZN(n3778) );
  INV_X1 U4452 ( .A(n3776), .ZN(n3777) );
  OAI22_X1 U4453 ( .A1(n3972), .A2(n3778), .B1(n3777), .B2(n4413), .ZN(n3779)
         );
  AOI21_X1 U4454 ( .B1(n3780), .B2(n4455), .A(n3779), .ZN(n3781) );
  OAI211_X1 U4455 ( .C1(n4471), .C2(n4151), .A(n3782), .B(n3781), .ZN(U3266)
         );
  OR2_X1 U4456 ( .A1(n2050), .A2(n3814), .ZN(n3806) );
  NAND2_X1 U4457 ( .A1(n3806), .A2(n3783), .ZN(n3784) );
  XOR2_X1 U4458 ( .A(n3789), .B(n3784), .Z(n4157) );
  INV_X1 U4459 ( .A(n4157), .ZN(n3805) );
  OAI21_X1 U4460 ( .B1(n3827), .B2(n3786), .A(n3785), .ZN(n3813) );
  NAND2_X1 U4461 ( .A1(n3813), .A2(n3814), .ZN(n3812) );
  NAND2_X1 U4462 ( .A1(n3812), .A2(n3787), .ZN(n3788) );
  XOR2_X1 U4463 ( .A(n3789), .B(n3788), .Z(n3790) );
  NAND2_X1 U4464 ( .A1(n3790), .A2(n4461), .ZN(n3794) );
  AOI22_X1 U4465 ( .A1(n3792), .A2(n4441), .B1(n3791), .B2(n4440), .ZN(n3793)
         );
  OAI211_X1 U4466 ( .C1(n3795), .C2(n4443), .A(n3794), .B(n3793), .ZN(n4156)
         );
  INV_X1 U4467 ( .A(n3796), .ZN(n4160) );
  OAI21_X1 U4468 ( .B1(n4160), .B2(n3798), .A(n3797), .ZN(n4225) );
  NOR2_X1 U4469 ( .A1(n4225), .A2(n3952), .ZN(n3803) );
  INV_X1 U4470 ( .A(REG2_REG_23__SCAN_IN), .ZN(n3801) );
  INV_X1 U4471 ( .A(n3799), .ZN(n3800) );
  OAI22_X1 U4472 ( .A1(n3972), .A2(n3801), .B1(n3800), .B2(n4413), .ZN(n3802)
         );
  AOI211_X1 U4473 ( .C1(n4156), .C2(n3935), .A(n3803), .B(n3802), .ZN(n3804)
         );
  OAI21_X1 U4474 ( .B1(n3805), .B2(n3955), .A(n3804), .ZN(U3267) );
  INV_X1 U4475 ( .A(n3806), .ZN(n3807) );
  AOI21_X1 U4476 ( .B1(n3814), .B2(n2050), .A(n3807), .ZN(n4164) );
  NAND2_X1 U4477 ( .A1(n4164), .A2(n3808), .ZN(n3824) );
  INV_X1 U4478 ( .A(REG2_REG_22__SCAN_IN), .ZN(n3810) );
  OAI22_X1 U4479 ( .A1(n3972), .A2(n3810), .B1(n3809), .B2(n4413), .ZN(n3811)
         );
  INV_X1 U4480 ( .A(n3811), .ZN(n3823) );
  OAI21_X1 U4481 ( .B1(n3814), .B2(n3813), .A(n3812), .ZN(n3815) );
  NAND2_X1 U4482 ( .A1(n3815), .A2(n4461), .ZN(n3819) );
  OAI22_X1 U4483 ( .A1(n3816), .A2(n4464), .B1(n3820), .B2(n4403), .ZN(n3817)
         );
  INV_X1 U4484 ( .A(n3817), .ZN(n3818) );
  OAI211_X1 U4485 ( .C1(n3849), .C2(n4443), .A(n3819), .B(n3818), .ZN(n4162)
         );
  NAND2_X1 U4486 ( .A1(n4162), .A2(n3972), .ZN(n3822) );
  NOR2_X1 U4487 ( .A1(n3833), .A2(n3820), .ZN(n4161) );
  OR3_X1 U4488 ( .A1(n4161), .A2(n4160), .A3(n3952), .ZN(n3821) );
  NAND4_X1 U4489 ( .A1(n3824), .A2(n3823), .A3(n3822), .A4(n3821), .ZN(U3268)
         );
  XOR2_X1 U4490 ( .A(n3826), .B(n3825), .Z(n4167) );
  INV_X1 U4491 ( .A(n4167), .ZN(n3843) );
  XNOR2_X1 U4492 ( .A(n3827), .B(n3826), .ZN(n3828) );
  NAND2_X1 U4493 ( .A1(n3828), .A2(n4461), .ZN(n3832) );
  AOI22_X1 U4494 ( .A1(n3830), .A2(n4441), .B1(n4440), .B2(n3829), .ZN(n3831)
         );
  OAI211_X1 U4495 ( .C1(n3870), .C2(n4443), .A(n3832), .B(n3831), .ZN(n4166)
         );
  INV_X1 U4496 ( .A(n3853), .ZN(n3836) );
  INV_X1 U4497 ( .A(n3833), .ZN(n3834) );
  OAI21_X1 U4498 ( .B1(n3836), .B2(n3835), .A(n3834), .ZN(n4230) );
  NOR2_X1 U4499 ( .A1(n4230), .A2(n3952), .ZN(n3841) );
  INV_X1 U4500 ( .A(REG2_REG_21__SCAN_IN), .ZN(n3839) );
  INV_X1 U4501 ( .A(n3837), .ZN(n3838) );
  OAI22_X1 U4502 ( .A1(n3972), .A2(n3839), .B1(n3838), .B2(n4413), .ZN(n3840)
         );
  AOI211_X1 U4503 ( .C1(n4166), .C2(n3935), .A(n3841), .B(n3840), .ZN(n3842)
         );
  OAI21_X1 U4504 ( .B1(n3843), .B2(n3955), .A(n3842), .ZN(U3269) );
  XNOR2_X1 U4505 ( .A(n3844), .B(n3847), .ZN(n4171) );
  INV_X1 U4506 ( .A(n4171), .ZN(n3860) );
  NAND2_X1 U4507 ( .A1(n3846), .A2(n3845), .ZN(n3848) );
  XNOR2_X1 U4508 ( .A(n3848), .B(n3847), .ZN(n3852) );
  OAI22_X1 U4509 ( .A1(n3849), .A2(n4464), .B1(n4403), .B2(n3854), .ZN(n3850)
         );
  AOI21_X1 U4510 ( .B1(n4407), .B2(n3887), .A(n3850), .ZN(n3851) );
  OAI21_X1 U4511 ( .B1(n3852), .B2(n4409), .A(n3851), .ZN(n4170) );
  INV_X1 U4512 ( .A(n3875), .ZN(n3855) );
  OAI21_X1 U4513 ( .B1(n3855), .B2(n3854), .A(n3853), .ZN(n4234) );
  AOI22_X1 U4514 ( .A1(n4471), .A2(REG2_REG_20__SCAN_IN), .B1(n3856), .B2(
        n4466), .ZN(n3857) );
  OAI21_X1 U4515 ( .B1(n4234), .B2(n3952), .A(n3857), .ZN(n3858) );
  AOI21_X1 U4516 ( .B1(n4170), .B2(n3972), .A(n3858), .ZN(n3859) );
  OAI21_X1 U4517 ( .B1(n3860), .B2(n3955), .A(n3859), .ZN(U3270) );
  XOR2_X1 U4518 ( .A(n3869), .B(n3861), .Z(n4175) );
  INV_X1 U4519 ( .A(n4175), .ZN(n3882) );
  INV_X1 U4520 ( .A(n3862), .ZN(n3864) );
  OAI21_X1 U4521 ( .B1(n3902), .B2(n3864), .A(n3863), .ZN(n3884) );
  INV_X1 U4522 ( .A(n3865), .ZN(n3867) );
  OAI21_X1 U4523 ( .B1(n3884), .B2(n3867), .A(n3866), .ZN(n3868) );
  XOR2_X1 U4524 ( .A(n3869), .B(n3868), .Z(n3874) );
  OAI22_X1 U4525 ( .A1(n3870), .A2(n4464), .B1(n4403), .B2(n3876), .ZN(n3871)
         );
  AOI21_X1 U4526 ( .B1(n4407), .B2(n3872), .A(n3871), .ZN(n3873) );
  OAI21_X1 U4527 ( .B1(n3874), .B2(n4409), .A(n3873), .ZN(n4174) );
  OAI21_X1 U4528 ( .B1(n3892), .B2(n3876), .A(n3875), .ZN(n4238) );
  NOR2_X1 U4529 ( .A1(n4238), .A2(n3952), .ZN(n3880) );
  INV_X1 U4530 ( .A(n3877), .ZN(n3878) );
  OAI22_X1 U4531 ( .A1(n3972), .A2(n3676), .B1(n3878), .B2(n4413), .ZN(n3879)
         );
  AOI211_X1 U4532 ( .C1(n4174), .C2(n3935), .A(n3880), .B(n3879), .ZN(n3881)
         );
  OAI21_X1 U4533 ( .B1(n3882), .B2(n3955), .A(n3881), .ZN(U3271) );
  XOR2_X1 U4534 ( .A(n3885), .B(n3883), .Z(n4180) );
  XOR2_X1 U4535 ( .A(n3885), .B(n3884), .Z(n3890) );
  AOI22_X1 U4536 ( .A1(n3887), .A2(n4441), .B1(n3886), .B2(n4440), .ZN(n3888)
         );
  OAI21_X1 U4537 ( .B1(n3923), .B2(n4443), .A(n3888), .ZN(n3889) );
  AOI21_X1 U4538 ( .B1(n3890), .B2(n4461), .A(n3889), .ZN(n4179) );
  INV_X1 U4539 ( .A(n4179), .ZN(n3899) );
  OAI21_X1 U4540 ( .B1(n3909), .B2(n3891), .A(n4540), .ZN(n3893) );
  OR2_X1 U4541 ( .A1(n3893), .A2(n3892), .ZN(n4178) );
  INV_X1 U4542 ( .A(n3894), .ZN(n3897) );
  AOI22_X1 U4543 ( .A1(n4471), .A2(REG2_REG_18__SCAN_IN), .B1(n3895), .B2(
        n4466), .ZN(n3896) );
  OAI21_X1 U4544 ( .B1(n4178), .B2(n3897), .A(n3896), .ZN(n3898) );
  AOI21_X1 U4545 ( .B1(n3899), .B2(n3972), .A(n3898), .ZN(n3900) );
  OAI21_X1 U4546 ( .B1(n4180), .B2(n3955), .A(n3900), .ZN(U3272) );
  XNOR2_X1 U4547 ( .A(n3901), .B(n3903), .ZN(n4182) );
  INV_X1 U4548 ( .A(n4182), .ZN(n3919) );
  XOR2_X1 U4549 ( .A(n3903), .B(n3902), .Z(n3908) );
  OAI22_X1 U4550 ( .A1(n3904), .A2(n4464), .B1(n4403), .B2(n3911), .ZN(n3905)
         );
  AOI21_X1 U4551 ( .B1(n4407), .B2(n3906), .A(n3905), .ZN(n3907) );
  OAI21_X1 U4552 ( .B1(n3908), .B2(n4409), .A(n3907), .ZN(n4181) );
  INV_X1 U4553 ( .A(n3927), .ZN(n3912) );
  INV_X1 U4554 ( .A(n3909), .ZN(n3910) );
  OAI21_X1 U4555 ( .B1(n3912), .B2(n3911), .A(n3910), .ZN(n4243) );
  NOR2_X1 U4556 ( .A1(n4243), .A2(n3952), .ZN(n3917) );
  INV_X1 U4557 ( .A(n3913), .ZN(n3914) );
  OAI22_X1 U4558 ( .A1(n3972), .A2(n3915), .B1(n3914), .B2(n4413), .ZN(n3916)
         );
  AOI211_X1 U4559 ( .C1(n4181), .C2(n3935), .A(n3917), .B(n3916), .ZN(n3918)
         );
  OAI21_X1 U4560 ( .B1(n3919), .B2(n3955), .A(n3918), .ZN(U3273) );
  XNOR2_X1 U4561 ( .A(n3920), .B(n3921), .ZN(n4186) );
  INV_X1 U4562 ( .A(n4186), .ZN(n3937) );
  XNOR2_X1 U4563 ( .A(n3922), .B(n3921), .ZN(n3926) );
  OAI22_X1 U4564 ( .A1(n3923), .A2(n4464), .B1(n4403), .B2(n3928), .ZN(n3924)
         );
  AOI21_X1 U4565 ( .B1(n4407), .B2(n3963), .A(n3924), .ZN(n3925) );
  OAI21_X1 U4566 ( .B1(n3926), .B2(n4409), .A(n3925), .ZN(n4185) );
  INV_X1 U4567 ( .A(n3949), .ZN(n3929) );
  OAI21_X1 U4568 ( .B1(n3929), .B2(n3928), .A(n3927), .ZN(n4247) );
  NOR2_X1 U4569 ( .A1(n4247), .A2(n3952), .ZN(n3934) );
  INV_X1 U4570 ( .A(REG2_REG_16__SCAN_IN), .ZN(n3932) );
  INV_X1 U4571 ( .A(n3930), .ZN(n3931) );
  OAI22_X1 U4572 ( .A1(n3935), .A2(n3932), .B1(n3931), .B2(n4413), .ZN(n3933)
         );
  AOI211_X1 U4573 ( .C1(n4185), .C2(n3935), .A(n3934), .B(n3933), .ZN(n3936)
         );
  OAI21_X1 U4574 ( .B1(n3937), .B2(n3955), .A(n3936), .ZN(U3274) );
  XOR2_X1 U4575 ( .A(n3938), .B(n3940), .Z(n4190) );
  INV_X1 U4576 ( .A(n4190), .ZN(n3956) );
  NAND2_X1 U4577 ( .A1(n3959), .A2(n3939), .ZN(n3941) );
  XNOR2_X1 U4578 ( .A(n3941), .B(n3940), .ZN(n3946) );
  OAI22_X1 U4579 ( .A1(n3942), .A2(n4464), .B1(n4403), .B2(n3947), .ZN(n3943)
         );
  AOI21_X1 U4580 ( .B1(n4407), .B2(n3944), .A(n3943), .ZN(n3945) );
  OAI21_X1 U4581 ( .B1(n3946), .B2(n4409), .A(n3945), .ZN(n4189) );
  OR2_X1 U4582 ( .A1(n3968), .A2(n3947), .ZN(n3948) );
  NAND2_X1 U4583 ( .A1(n3949), .A2(n3948), .ZN(n4252) );
  AOI22_X1 U4584 ( .A1(n4471), .A2(REG2_REG_15__SCAN_IN), .B1(n3950), .B2(
        n4466), .ZN(n3951) );
  OAI21_X1 U4585 ( .B1(n4252), .B2(n3952), .A(n3951), .ZN(n3953) );
  AOI21_X1 U4586 ( .B1(n4189), .B2(n3972), .A(n3953), .ZN(n3954) );
  OAI21_X1 U4587 ( .B1(n3956), .B2(n3955), .A(n3954), .ZN(U3275) );
  XNOR2_X1 U4588 ( .A(n3958), .B(n3957), .ZN(n4194) );
  OAI21_X1 U4589 ( .B1(n3961), .B2(n3960), .A(n3959), .ZN(n3962) );
  NAND2_X1 U4590 ( .A1(n3962), .A2(n4461), .ZN(n3965) );
  AOI22_X1 U4591 ( .A1(n3963), .A2(n4441), .B1(n4440), .B2(n3969), .ZN(n3964)
         );
  OAI211_X1 U4592 ( .C1(n3966), .C2(n4443), .A(n3965), .B(n3964), .ZN(n3967)
         );
  AOI21_X1 U4593 ( .B1(n4194), .B2(n4462), .A(n3967), .ZN(n4198) );
  INV_X1 U4594 ( .A(n3968), .ZN(n4196) );
  NAND2_X1 U4595 ( .A1(n2062), .A2(n3969), .ZN(n4195) );
  AND3_X1 U4596 ( .A1(n4196), .A2(n4455), .A3(n4195), .ZN(n3974) );
  INV_X1 U4597 ( .A(n3970), .ZN(n3971) );
  OAI22_X1 U4598 ( .A1(n3972), .A2(n3076), .B1(n3971), .B2(n4413), .ZN(n3973)
         );
  AOI211_X1 U4599 ( .C1(n4194), .C2(n4467), .A(n3974), .B(n3973), .ZN(n3975)
         );
  OAI21_X1 U4600 ( .B1(n4198), .B2(n4471), .A(n3975), .ZN(U3276) );
  XNOR2_X1 U4601 ( .A(n3982), .B(n3978), .ZN(n4269) );
  INV_X1 U4602 ( .A(n4269), .ZN(n4206) );
  NAND2_X1 U4603 ( .A1(n3977), .A2(n3976), .ZN(n3986) );
  NAND2_X1 U4604 ( .A1(n3978), .A2(n4440), .ZN(n3979) );
  AND2_X1 U4605 ( .A1(n3986), .A2(n3979), .ZN(n4271) );
  INV_X1 U4606 ( .A(REG1_REG_31__SCAN_IN), .ZN(n3980) );
  MUX2_X1 U4607 ( .A(n4271), .B(n3980), .S(n4576), .Z(n3981) );
  OAI21_X1 U4608 ( .B1(n4206), .B2(n4193), .A(n3981), .ZN(U3549) );
  INV_X1 U4609 ( .A(REG1_REG_30__SCAN_IN), .ZN(n3990) );
  AOI21_X1 U4610 ( .B1(n3984), .B2(n3983), .A(n3982), .ZN(n4273) );
  NAND2_X1 U4611 ( .A1(n4273), .A2(n3985), .ZN(n3989) );
  OAI21_X1 U4612 ( .B1(n3987), .B2(n4403), .A(n3986), .ZN(n4272) );
  NAND2_X1 U4613 ( .A1(n4579), .A2(n4272), .ZN(n3988) );
  OAI211_X1 U4614 ( .C1(n4579), .C2(n3990), .A(n3989), .B(n3988), .ZN(U3548)
         );
  MUX2_X1 U4615 ( .A(REG1_REG_29__SCAN_IN), .B(n4211), .S(n4579), .Z(U3547) );
  AOI21_X1 U4616 ( .B1(n4540), .B2(n3995), .A(n3994), .ZN(n3996) );
  OAI21_X1 U4617 ( .B1(n3997), .B2(n4535), .A(n3996), .ZN(n4212) );
  MUX2_X1 U4618 ( .A(REG1_REG_27__SCAN_IN), .B(n4212), .S(n4579), .Z(U3545) );
  NOR2_X1 U4619 ( .A1(keyinput54), .A2(keyinput25), .ZN(n4008) );
  NAND3_X1 U4620 ( .A1(keyinput56), .A2(keyinput3), .A3(keyinput49), .ZN(n4000) );
  NAND4_X1 U4621 ( .A1(keyinput55), .A2(keyinput22), .A3(keyinput47), .A4(
        keyinput1), .ZN(n3999) );
  NAND4_X1 U4622 ( .A1(keyinput50), .A2(keyinput10), .A3(keyinput21), .A4(
        keyinput33), .ZN(n3998) );
  NOR4_X1 U4623 ( .A1(keyinput5), .A2(n4000), .A3(n3999), .A4(n3998), .ZN(
        n4007) );
  NAND4_X1 U4624 ( .A1(keyinput17), .A2(keyinput30), .A3(keyinput27), .A4(
        keyinput11), .ZN(n4005) );
  NAND3_X1 U4625 ( .A1(keyinput38), .A2(keyinput46), .A3(keyinput60), .ZN(
        n4004) );
  NOR3_X1 U4626 ( .A1(keyinput2), .A2(keyinput32), .A3(keyinput16), .ZN(n4002)
         );
  NOR3_X1 U4627 ( .A1(keyinput36), .A2(keyinput8), .A3(keyinput41), .ZN(n4001)
         );
  NAND4_X1 U4628 ( .A1(keyinput42), .A2(n4002), .A3(keyinput45), .A4(n4001), 
        .ZN(n4003) );
  NOR4_X1 U4629 ( .A1(keyinput44), .A2(n4005), .A3(n4004), .A4(n4003), .ZN(
        n4006) );
  NAND4_X1 U4630 ( .A1(keyinput26), .A2(n4008), .A3(n4007), .A4(n4006), .ZN(
        n4023) );
  NAND4_X1 U4631 ( .A1(keyinput58), .A2(keyinput39), .A3(keyinput23), .A4(
        keyinput24), .ZN(n4010) );
  NAND2_X1 U4632 ( .A1(keyinput31), .A2(keyinput48), .ZN(n4009) );
  NOR4_X1 U4633 ( .A1(keyinput7), .A2(keyinput15), .A3(n4010), .A4(n4009), 
        .ZN(n4021) );
  NAND3_X1 U4634 ( .A1(keyinput9), .A2(keyinput28), .A3(keyinput59), .ZN(n4012) );
  NAND3_X1 U4635 ( .A1(keyinput29), .A2(keyinput53), .A3(keyinput43), .ZN(
        n4011) );
  NOR4_X1 U4636 ( .A1(keyinput14), .A2(keyinput40), .A3(n4012), .A4(n4011), 
        .ZN(n4020) );
  NAND3_X1 U4637 ( .A1(keyinput0), .A2(keyinput20), .A3(keyinput51), .ZN(n4014) );
  NAND3_X1 U4638 ( .A1(keyinput34), .A2(keyinput12), .A3(keyinput4), .ZN(n4013) );
  NOR4_X1 U4639 ( .A1(keyinput37), .A2(keyinput19), .A3(n4014), .A4(n4013), 
        .ZN(n4019) );
  NAND2_X1 U4640 ( .A1(keyinput6), .A2(keyinput35), .ZN(n4017) );
  INV_X1 U4641 ( .A(keyinput57), .ZN(n4015) );
  NAND4_X1 U4642 ( .A1(keyinput18), .A2(keyinput61), .A3(keyinput63), .A4(
        n4015), .ZN(n4016) );
  NOR4_X1 U4643 ( .A1(keyinput62), .A2(keyinput52), .A3(n4017), .A4(n4016), 
        .ZN(n4018) );
  NAND4_X1 U4644 ( .A1(n4021), .A2(n4020), .A3(n4019), .A4(n4018), .ZN(n4022)
         );
  OAI21_X1 U4645 ( .B1(n4023), .B2(n4022), .A(keyinput13), .ZN(n4140) );
  INV_X1 U4646 ( .A(B_REG_SCAN_IN), .ZN(n4026) );
  INV_X1 U4647 ( .A(keyinput22), .ZN(n4025) );
  AOI22_X1 U4648 ( .A1(n4026), .A2(keyinput47), .B1(DATAO_REG_9__SCAN_IN), 
        .B2(n4025), .ZN(n4024) );
  OAI221_X1 U4649 ( .B1(n4026), .B2(keyinput47), .C1(n4025), .C2(
        DATAO_REG_9__SCAN_IN), .A(n4024), .ZN(n4037) );
  INV_X1 U4650 ( .A(REG2_REG_30__SCAN_IN), .ZN(n4275) );
  AOI22_X1 U4651 ( .A1(n4275), .A2(keyinput1), .B1(n3810), .B2(keyinput50), 
        .ZN(n4027) );
  OAI221_X1 U4652 ( .B1(n4275), .B2(keyinput1), .C1(n3810), .C2(keyinput50), 
        .A(n4027), .ZN(n4036) );
  INV_X1 U4653 ( .A(keyinput10), .ZN(n4029) );
  AOI22_X1 U4654 ( .A1(n4030), .A2(keyinput21), .B1(REG0_REG_31__SCAN_IN), 
        .B2(n4029), .ZN(n4028) );
  OAI221_X1 U4655 ( .B1(n4030), .B2(keyinput21), .C1(n4029), .C2(
        REG0_REG_31__SCAN_IN), .A(n4028), .ZN(n4035) );
  INV_X1 U4656 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4033) );
  INV_X1 U4657 ( .A(REG3_REG_12__SCAN_IN), .ZN(n4032) );
  AOI22_X1 U4658 ( .A1(n4033), .A2(keyinput33), .B1(n4032), .B2(keyinput9), 
        .ZN(n4031) );
  OAI221_X1 U4659 ( .B1(n4033), .B2(keyinput33), .C1(n4032), .C2(keyinput9), 
        .A(n4031), .ZN(n4034) );
  NOR4_X1 U4660 ( .A1(n4037), .A2(n4036), .A3(n4035), .A4(n4034), .ZN(n4078)
         );
  INV_X1 U4661 ( .A(DATAI_10_), .ZN(n4496) );
  AOI22_X1 U4662 ( .A1(n4039), .A2(keyinput11), .B1(keyinput38), .B2(n4496), 
        .ZN(n4038) );
  OAI221_X1 U4663 ( .B1(n4039), .B2(keyinput11), .C1(n4496), .C2(keyinput38), 
        .A(n4038), .ZN(n4042) );
  INV_X1 U4664 ( .A(D_REG_31__SCAN_IN), .ZN(n4472) );
  AOI22_X1 U4665 ( .A1(n4477), .A2(keyinput42), .B1(keyinput32), .B2(n4472), 
        .ZN(n4040) );
  OAI221_X1 U4666 ( .B1(n4477), .B2(keyinput42), .C1(n4472), .C2(keyinput32), 
        .A(n4040), .ZN(n4041) );
  NOR2_X1 U4667 ( .A1(n4042), .A2(n4041), .ZN(n4052) );
  INV_X1 U4668 ( .A(REG0_REG_9__SCAN_IN), .ZN(n4551) );
  INV_X1 U4669 ( .A(REG0_REG_6__SCAN_IN), .ZN(n4044) );
  AOI22_X1 U4670 ( .A1(n4551), .A2(keyinput62), .B1(keyinput52), .B2(n4044), 
        .ZN(n4043) );
  OAI221_X1 U4671 ( .B1(n4551), .B2(keyinput62), .C1(n4044), .C2(keyinput52), 
        .A(n4043), .ZN(n4050) );
  XNOR2_X1 U4672 ( .A(IR_REG_14__SCAN_IN), .B(keyinput44), .ZN(n4048) );
  XNOR2_X1 U4673 ( .A(IR_REG_23__SCAN_IN), .B(keyinput30), .ZN(n4047) );
  XNOR2_X1 U4674 ( .A(IR_REG_21__SCAN_IN), .B(keyinput46), .ZN(n4046) );
  XNOR2_X1 U4675 ( .A(IR_REG_24__SCAN_IN), .B(keyinput36), .ZN(n4045) );
  NAND4_X1 U4676 ( .A1(n4048), .A2(n4047), .A3(n4046), .A4(n4045), .ZN(n4049)
         );
  NOR2_X1 U4677 ( .A1(n4050), .A2(n4049), .ZN(n4051) );
  AND2_X1 U4678 ( .A1(n4052), .A2(n4051), .ZN(n4077) );
  AOI22_X1 U4679 ( .A1(n4054), .A2(keyinput35), .B1(keyinput61), .B2(n4469), 
        .ZN(n4053) );
  OAI221_X1 U4680 ( .B1(n4054), .B2(keyinput35), .C1(n4469), .C2(keyinput61), 
        .A(n4053), .ZN(n4057) );
  INV_X1 U4681 ( .A(D_REG_20__SCAN_IN), .ZN(n4475) );
  INV_X1 U4682 ( .A(D_REG_3__SCAN_IN), .ZN(n4478) );
  AOI22_X1 U4683 ( .A1(n4475), .A2(keyinput16), .B1(keyinput17), .B2(n4478), 
        .ZN(n4055) );
  OAI221_X1 U4684 ( .B1(n4475), .B2(keyinput16), .C1(n4478), .C2(keyinput17), 
        .A(n4055), .ZN(n4056) );
  NOR2_X1 U4685 ( .A1(n4057), .A2(n4056), .ZN(n4076) );
  INV_X1 U4686 ( .A(DATAI_0_), .ZN(n4504) );
  AOI22_X1 U4687 ( .A1(n4504), .A2(keyinput25), .B1(n4059), .B2(keyinput45), 
        .ZN(n4058) );
  OAI221_X1 U4688 ( .B1(n4504), .B2(keyinput25), .C1(n4059), .C2(keyinput45), 
        .A(n4058), .ZN(n4063) );
  XNOR2_X1 U4689 ( .A(REG0_REG_20__SCAN_IN), .B(keyinput0), .ZN(n4061) );
  XNOR2_X1 U4690 ( .A(keyinput18), .B(REG0_REG_1__SCAN_IN), .ZN(n4060) );
  NAND2_X1 U4691 ( .A1(n4061), .A2(n4060), .ZN(n4062) );
  NOR2_X1 U4692 ( .A1(n4063), .A2(n4062), .ZN(n4074) );
  INV_X1 U4693 ( .A(DATAI_8_), .ZN(n4066) );
  INV_X1 U4694 ( .A(DATAI_20_), .ZN(n4065) );
  AOI22_X1 U4695 ( .A1(n4066), .A2(keyinput8), .B1(n4065), .B2(keyinput41), 
        .ZN(n4064) );
  OAI221_X1 U4696 ( .B1(n4066), .B2(keyinput8), .C1(n4065), .C2(keyinput41), 
        .A(n4064), .ZN(n4072) );
  XNOR2_X1 U4697 ( .A(IR_REG_1__SCAN_IN), .B(keyinput63), .ZN(n4070) );
  XNOR2_X1 U4698 ( .A(IR_REG_4__SCAN_IN), .B(keyinput60), .ZN(n4069) );
  XNOR2_X1 U4699 ( .A(IR_REG_8__SCAN_IN), .B(keyinput27), .ZN(n4068) );
  XNOR2_X1 U4700 ( .A(IR_REG_7__SCAN_IN), .B(keyinput57), .ZN(n4067) );
  NAND4_X1 U4701 ( .A1(n4070), .A2(n4069), .A3(n4068), .A4(n4067), .ZN(n4071)
         );
  NOR2_X1 U4702 ( .A1(n4072), .A2(n4071), .ZN(n4073) );
  AND2_X1 U4703 ( .A1(n4074), .A2(n4073), .ZN(n4075) );
  NAND4_X1 U4704 ( .A1(n4078), .A2(n4077), .A3(n4076), .A4(n4075), .ZN(n4139)
         );
  AOI22_X1 U4705 ( .A1(keyinput26), .A2(n4080), .B1(keyinput13), .B2(n4183), 
        .ZN(n4079) );
  OAI21_X1 U4706 ( .B1(n4080), .B2(keyinput26), .A(n4079), .ZN(n4093) );
  INV_X1 U4707 ( .A(REG2_REG_25__SCAN_IN), .ZN(n4083) );
  INV_X1 U4708 ( .A(keyinput56), .ZN(n4082) );
  AOI22_X1 U4709 ( .A1(n4083), .A2(keyinput54), .B1(DATAI_30_), .B2(n4082), 
        .ZN(n4081) );
  OAI221_X1 U4710 ( .B1(n4083), .B2(keyinput54), .C1(n4082), .C2(DATAI_30_), 
        .A(n4081), .ZN(n4092) );
  INV_X1 U4711 ( .A(keyinput5), .ZN(n4086) );
  INV_X1 U4712 ( .A(keyinput3), .ZN(n4085) );
  AOI22_X1 U4713 ( .A1(n4086), .A2(DATAO_REG_8__SCAN_IN), .B1(
        DATAO_REG_12__SCAN_IN), .B2(n4085), .ZN(n4084) );
  OAI221_X1 U4714 ( .B1(n4086), .B2(DATAO_REG_8__SCAN_IN), .C1(n4085), .C2(
        DATAO_REG_12__SCAN_IN), .A(n4084), .ZN(n4091) );
  INV_X1 U4715 ( .A(keyinput49), .ZN(n4089) );
  INV_X1 U4716 ( .A(keyinput55), .ZN(n4088) );
  AOI22_X1 U4717 ( .A1(n4089), .A2(DATAO_REG_3__SCAN_IN), .B1(
        DATAO_REG_5__SCAN_IN), .B2(n4088), .ZN(n4087) );
  OAI221_X1 U4718 ( .B1(n4089), .B2(DATAO_REG_3__SCAN_IN), .C1(n4088), .C2(
        DATAO_REG_5__SCAN_IN), .A(n4087), .ZN(n4090) );
  NOR4_X1 U4719 ( .A1(n4093), .A2(n4092), .A3(n4091), .A4(n4090), .ZN(n4137)
         );
  INV_X1 U4720 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4149) );
  INV_X1 U4721 ( .A(DATAI_25_), .ZN(n4095) );
  AOI22_X1 U4722 ( .A1(n4149), .A2(keyinput51), .B1(keyinput34), .B2(n4095), 
        .ZN(n4094) );
  OAI221_X1 U4723 ( .B1(n4149), .B2(keyinput51), .C1(n4095), .C2(keyinput34), 
        .A(n4094), .ZN(n4103) );
  INV_X1 U4724 ( .A(DATAI_23_), .ZN(n4482) );
  INV_X1 U4725 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4154) );
  AOI22_X1 U4726 ( .A1(n4482), .A2(keyinput20), .B1(n4154), .B2(keyinput37), 
        .ZN(n4096) );
  OAI221_X1 U4727 ( .B1(n4482), .B2(keyinput20), .C1(n4154), .C2(keyinput37), 
        .A(n4096), .ZN(n4102) );
  AOI22_X1 U4728 ( .A1(n4476), .A2(keyinput4), .B1(keyinput2), .B2(n4473), 
        .ZN(n4097) );
  OAI221_X1 U4729 ( .B1(n4476), .B2(keyinput4), .C1(n4473), .C2(keyinput2), 
        .A(n4097), .ZN(n4101) );
  AOI22_X1 U4730 ( .A1(n4099), .A2(keyinput19), .B1(keyinput12), .B2(n4474), 
        .ZN(n4098) );
  OAI221_X1 U4731 ( .B1(n4099), .B2(keyinput19), .C1(n4474), .C2(keyinput12), 
        .A(n4098), .ZN(n4100) );
  NOR4_X1 U4732 ( .A1(n4103), .A2(n4102), .A3(n4101), .A4(n4100), .ZN(n4136)
         );
  AOI22_X1 U4733 ( .A1(n4345), .A2(keyinput31), .B1(n4105), .B2(keyinput48), 
        .ZN(n4104) );
  OAI221_X1 U4734 ( .B1(n4345), .B2(keyinput31), .C1(n4105), .C2(keyinput48), 
        .A(n4104), .ZN(n4117) );
  INV_X1 U4735 ( .A(keyinput7), .ZN(n4108) );
  INV_X1 U4736 ( .A(keyinput40), .ZN(n4107) );
  AOI22_X1 U4737 ( .A1(n4108), .A2(DATAI_31_), .B1(DATAO_REG_16__SCAN_IN), 
        .B2(n4107), .ZN(n4106) );
  OAI221_X1 U4738 ( .B1(n4108), .B2(DATAI_31_), .C1(n4107), .C2(
        DATAO_REG_16__SCAN_IN), .A(n4106), .ZN(n4116) );
  INV_X1 U4739 ( .A(REG0_REG_28__SCAN_IN), .ZN(n4111) );
  INV_X1 U4740 ( .A(keyinput29), .ZN(n4110) );
  AOI22_X1 U4741 ( .A1(n4111), .A2(keyinput53), .B1(DATAO_REG_22__SCAN_IN), 
        .B2(n4110), .ZN(n4109) );
  OAI221_X1 U4742 ( .B1(n4111), .B2(keyinput53), .C1(n4110), .C2(
        DATAO_REG_22__SCAN_IN), .A(n4109), .ZN(n4115) );
  INV_X1 U4743 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4210) );
  INV_X1 U4744 ( .A(keyinput6), .ZN(n4113) );
  AOI22_X1 U4745 ( .A1(n4210), .A2(keyinput43), .B1(REG1_REG_31__SCAN_IN), 
        .B2(n4113), .ZN(n4112) );
  OAI221_X1 U4746 ( .B1(n4210), .B2(keyinput43), .C1(n4113), .C2(
        REG1_REG_31__SCAN_IN), .A(n4112), .ZN(n4114) );
  NOR4_X1 U4747 ( .A1(n4117), .A2(n4116), .A3(n4115), .A4(n4114), .ZN(n4135)
         );
  INV_X1 U4748 ( .A(REG3_REG_2__SCAN_IN), .ZN(n4120) );
  INV_X1 U4749 ( .A(keyinput59), .ZN(n4119) );
  AOI22_X1 U4750 ( .A1(n4120), .A2(keyinput28), .B1(ADDR_REG_2__SCAN_IN), .B2(
        n4119), .ZN(n4118) );
  OAI221_X1 U4751 ( .B1(n4120), .B2(keyinput28), .C1(n4119), .C2(
        ADDR_REG_2__SCAN_IN), .A(n4118), .ZN(n4133) );
  INV_X1 U4752 ( .A(keyinput14), .ZN(n4123) );
  INV_X1 U4753 ( .A(keyinput58), .ZN(n4122) );
  AOI22_X1 U4754 ( .A1(n4123), .A2(ADDR_REG_5__SCAN_IN), .B1(
        ADDR_REG_6__SCAN_IN), .B2(n4122), .ZN(n4121) );
  OAI221_X1 U4755 ( .B1(n4123), .B2(ADDR_REG_5__SCAN_IN), .C1(n4122), .C2(
        ADDR_REG_6__SCAN_IN), .A(n4121), .ZN(n4132) );
  INV_X1 U4756 ( .A(keyinput39), .ZN(n4126) );
  INV_X1 U4757 ( .A(keyinput23), .ZN(n4125) );
  AOI22_X1 U4758 ( .A1(n4126), .A2(ADDR_REG_8__SCAN_IN), .B1(
        ADDR_REG_11__SCAN_IN), .B2(n4125), .ZN(n4124) );
  OAI221_X1 U4759 ( .B1(n4126), .B2(ADDR_REG_8__SCAN_IN), .C1(n4125), .C2(
        ADDR_REG_11__SCAN_IN), .A(n4124), .ZN(n4131) );
  INV_X1 U4760 ( .A(REG2_REG_12__SCAN_IN), .ZN(n4129) );
  INV_X1 U4761 ( .A(keyinput15), .ZN(n4128) );
  AOI22_X1 U4762 ( .A1(n4129), .A2(keyinput24), .B1(ADDR_REG_12__SCAN_IN), 
        .B2(n4128), .ZN(n4127) );
  OAI221_X1 U4763 ( .B1(n4129), .B2(keyinput24), .C1(n4128), .C2(
        ADDR_REG_12__SCAN_IN), .A(n4127), .ZN(n4130) );
  NOR4_X1 U4764 ( .A1(n4133), .A2(n4132), .A3(n4131), .A4(n4130), .ZN(n4134)
         );
  NAND4_X1 U4765 ( .A1(n4137), .A2(n4136), .A3(n4135), .A4(n4134), .ZN(n4138)
         );
  AOI211_X1 U4766 ( .C1(REG1_REG_17__SCAN_IN), .C2(n4140), .A(n4139), .B(n4138), .ZN(n4146) );
  OAI21_X1 U4767 ( .B1(n4144), .B2(n4535), .A(n4143), .ZN(n4213) );
  XOR2_X1 U4768 ( .A(n4146), .B(n4145), .Z(U3544) );
  AOI21_X1 U4769 ( .B1(n4148), .B2(n4550), .A(n4147), .ZN(n4214) );
  MUX2_X1 U4770 ( .A(n4149), .B(n4214), .S(n4579), .Z(n4150) );
  OAI21_X1 U4771 ( .B1(n4193), .B2(n4217), .A(n4150), .ZN(U3543) );
  INV_X1 U4772 ( .A(n4151), .ZN(n4152) );
  AOI21_X1 U4773 ( .B1(n4153), .B2(n4550), .A(n4152), .ZN(n4218) );
  MUX2_X1 U4774 ( .A(n4154), .B(n4218), .S(n4579), .Z(n4155) );
  OAI21_X1 U4775 ( .B1(n4193), .B2(n4221), .A(n4155), .ZN(U3542) );
  INV_X1 U4776 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4158) );
  AOI21_X1 U4777 ( .B1(n4157), .B2(n4550), .A(n4156), .ZN(n4222) );
  MUX2_X1 U4778 ( .A(n4158), .B(n4222), .S(n4579), .Z(n4159) );
  OAI21_X1 U4779 ( .B1(n4193), .B2(n4225), .A(n4159), .ZN(U3541) );
  NOR3_X1 U4780 ( .A1(n4161), .A2(n4160), .A3(n2841), .ZN(n4163) );
  AOI211_X1 U4781 ( .C1(n4164), .C2(n4550), .A(n4163), .B(n4162), .ZN(n4165)
         );
  INV_X1 U4782 ( .A(n4165), .ZN(n4226) );
  MUX2_X1 U4783 ( .A(REG1_REG_22__SCAN_IN), .B(n4226), .S(n4579), .Z(U3540) );
  INV_X1 U4784 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4168) );
  AOI21_X1 U4785 ( .B1(n4167), .B2(n4550), .A(n4166), .ZN(n4227) );
  MUX2_X1 U4786 ( .A(n4168), .B(n4227), .S(n4579), .Z(n4169) );
  OAI21_X1 U4787 ( .B1(n4193), .B2(n4230), .A(n4169), .ZN(U3539) );
  INV_X1 U4788 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4172) );
  AOI21_X1 U4789 ( .B1(n4171), .B2(n4550), .A(n4170), .ZN(n4231) );
  MUX2_X1 U4790 ( .A(n4172), .B(n4231), .S(n4579), .Z(n4173) );
  OAI21_X1 U4791 ( .B1(n4193), .B2(n4234), .A(n4173), .ZN(U3538) );
  INV_X1 U4792 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4176) );
  AOI21_X1 U4793 ( .B1(n4175), .B2(n4550), .A(n4174), .ZN(n4235) );
  MUX2_X1 U4794 ( .A(n4176), .B(n4235), .S(n4579), .Z(n4177) );
  OAI21_X1 U4795 ( .B1(n4193), .B2(n4238), .A(n4177), .ZN(U3537) );
  OAI211_X1 U4796 ( .C1(n4180), .C2(n4535), .A(n4179), .B(n4178), .ZN(n4239)
         );
  MUX2_X1 U4797 ( .A(REG1_REG_18__SCAN_IN), .B(n4239), .S(n4579), .Z(U3536) );
  AOI21_X1 U4798 ( .B1(n4182), .B2(n4550), .A(n4181), .ZN(n4240) );
  MUX2_X1 U4799 ( .A(n4183), .B(n4240), .S(n4579), .Z(n4184) );
  OAI21_X1 U4800 ( .B1(n4193), .B2(n4243), .A(n4184), .ZN(U3535) );
  INV_X1 U4801 ( .A(REG1_REG_16__SCAN_IN), .ZN(n4187) );
  AOI21_X1 U4802 ( .B1(n4186), .B2(n4550), .A(n4185), .ZN(n4244) );
  MUX2_X1 U4803 ( .A(n4187), .B(n4244), .S(n4579), .Z(n4188) );
  OAI21_X1 U4804 ( .B1(n4193), .B2(n4247), .A(n4188), .ZN(U3534) );
  AOI21_X1 U4805 ( .B1(n4190), .B2(n4550), .A(n4189), .ZN(n4248) );
  MUX2_X1 U4806 ( .A(n4191), .B(n4248), .S(n4579), .Z(n4192) );
  OAI21_X1 U4807 ( .B1(n4193), .B2(n4252), .A(n4192), .ZN(U3533) );
  INV_X1 U4808 ( .A(n4194), .ZN(n4199) );
  NAND3_X1 U4809 ( .A1(n4196), .A2(n4540), .A3(n4195), .ZN(n4197) );
  OAI211_X1 U4810 ( .C1(n4199), .C2(n4524), .A(n4198), .B(n4197), .ZN(n4253)
         );
  MUX2_X1 U4811 ( .A(REG1_REG_14__SCAN_IN), .B(n4253), .S(n4579), .Z(U3532) );
  NAND2_X1 U4812 ( .A1(n4200), .A2(n4550), .ZN(n4202) );
  OAI211_X1 U4813 ( .C1(n2841), .C2(n4203), .A(n4202), .B(n4201), .ZN(n4254)
         );
  MUX2_X1 U4814 ( .A(REG1_REG_13__SCAN_IN), .B(n4254), .S(n4579), .Z(U3531) );
  INV_X1 U4815 ( .A(REG0_REG_31__SCAN_IN), .ZN(n4204) );
  MUX2_X1 U4816 ( .A(n4271), .B(n4204), .S(n4558), .Z(n4205) );
  OAI21_X1 U4817 ( .B1(n4206), .B2(n4251), .A(n4205), .ZN(U3517) );
  NAND2_X1 U4818 ( .A1(n4273), .A2(n4207), .ZN(n4209) );
  NAND2_X1 U4819 ( .A1(n4560), .A2(n4272), .ZN(n4208) );
  OAI211_X1 U4820 ( .C1(n4560), .C2(n4210), .A(n4209), .B(n4208), .ZN(U3516)
         );
  MUX2_X1 U4821 ( .A(REG0_REG_29__SCAN_IN), .B(n4211), .S(n4560), .Z(U3515) );
  MUX2_X1 U4822 ( .A(REG0_REG_27__SCAN_IN), .B(n4212), .S(n4560), .Z(U3513) );
  MUX2_X1 U4823 ( .A(REG0_REG_26__SCAN_IN), .B(n4213), .S(n4560), .Z(U3512) );
  INV_X1 U4824 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4215) );
  MUX2_X1 U4825 ( .A(n4215), .B(n4214), .S(n4560), .Z(n4216) );
  OAI21_X1 U4826 ( .B1(n4217), .B2(n4251), .A(n4216), .ZN(U3511) );
  INV_X1 U4827 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4219) );
  MUX2_X1 U4828 ( .A(n4219), .B(n4218), .S(n4560), .Z(n4220) );
  OAI21_X1 U4829 ( .B1(n4221), .B2(n4251), .A(n4220), .ZN(U3510) );
  INV_X1 U4830 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4223) );
  MUX2_X1 U4831 ( .A(n4223), .B(n4222), .S(n4560), .Z(n4224) );
  OAI21_X1 U4832 ( .B1(n4225), .B2(n4251), .A(n4224), .ZN(U3509) );
  MUX2_X1 U4833 ( .A(REG0_REG_22__SCAN_IN), .B(n4226), .S(n4560), .Z(U3508) );
  INV_X1 U4834 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4228) );
  MUX2_X1 U4835 ( .A(n4228), .B(n4227), .S(n4560), .Z(n4229) );
  OAI21_X1 U4836 ( .B1(n4230), .B2(n4251), .A(n4229), .ZN(U3507) );
  INV_X1 U4837 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4232) );
  MUX2_X1 U4838 ( .A(n4232), .B(n4231), .S(n4560), .Z(n4233) );
  OAI21_X1 U4839 ( .B1(n4234), .B2(n4251), .A(n4233), .ZN(U3506) );
  INV_X1 U4840 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4236) );
  MUX2_X1 U4841 ( .A(n4236), .B(n4235), .S(n4560), .Z(n4237) );
  OAI21_X1 U4842 ( .B1(n4238), .B2(n4251), .A(n4237), .ZN(U3505) );
  MUX2_X1 U4843 ( .A(REG0_REG_18__SCAN_IN), .B(n4239), .S(n4560), .Z(U3503) );
  INV_X1 U4844 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4241) );
  MUX2_X1 U4845 ( .A(n4241), .B(n4240), .S(n4560), .Z(n4242) );
  OAI21_X1 U4846 ( .B1(n4243), .B2(n4251), .A(n4242), .ZN(U3501) );
  INV_X1 U4847 ( .A(REG0_REG_16__SCAN_IN), .ZN(n4245) );
  MUX2_X1 U4848 ( .A(n4245), .B(n4244), .S(n4560), .Z(n4246) );
  OAI21_X1 U4849 ( .B1(n4247), .B2(n4251), .A(n4246), .ZN(U3499) );
  INV_X1 U4850 ( .A(REG0_REG_15__SCAN_IN), .ZN(n4249) );
  MUX2_X1 U4851 ( .A(n4249), .B(n4248), .S(n4560), .Z(n4250) );
  OAI21_X1 U4852 ( .B1(n4252), .B2(n4251), .A(n4250), .ZN(U3497) );
  MUX2_X1 U4853 ( .A(REG0_REG_14__SCAN_IN), .B(n4253), .S(n4560), .Z(U3495) );
  MUX2_X1 U4854 ( .A(REG0_REG_13__SCAN_IN), .B(n4254), .S(n4560), .Z(U3493) );
  MUX2_X1 U4855 ( .A(DATAI_30_), .B(n4255), .S(STATE_REG_SCAN_IN), .Z(U3322)
         );
  MUX2_X1 U4856 ( .A(DATAI_28_), .B(n4256), .S(STATE_REG_SCAN_IN), .Z(U3324)
         );
  MUX2_X1 U4857 ( .A(n4277), .B(DATAI_27_), .S(U3149), .Z(U3325) );
  MUX2_X1 U4858 ( .A(n2692), .B(DATAI_26_), .S(U3149), .Z(U3326) );
  MUX2_X1 U4859 ( .A(DATAI_25_), .B(n4257), .S(STATE_REG_SCAN_IN), .Z(U3327)
         );
  MUX2_X1 U4860 ( .A(n4258), .B(DATAI_22_), .S(U3149), .Z(U3330) );
  MUX2_X1 U4861 ( .A(n4259), .B(DATAI_21_), .S(U3149), .Z(U3331) );
  MUX2_X1 U4862 ( .A(DATAI_20_), .B(n4260), .S(STATE_REG_SCAN_IN), .Z(U3332)
         );
  MUX2_X1 U4863 ( .A(DATAI_19_), .B(n4261), .S(STATE_REG_SCAN_IN), .Z(U3333)
         );
  MUX2_X1 U4864 ( .A(n4262), .B(DATAI_14_), .S(U3149), .Z(U3338) );
  MUX2_X1 U4865 ( .A(n4263), .B(DATAI_8_), .S(U3149), .Z(U3344) );
  MUX2_X1 U4866 ( .A(n4264), .B(DATAI_7_), .S(U3149), .Z(U3345) );
  MUX2_X1 U4867 ( .A(DATAI_4_), .B(n4265), .S(STATE_REG_SCAN_IN), .Z(U3348) );
  MUX2_X1 U4868 ( .A(DATAI_3_), .B(n4266), .S(STATE_REG_SCAN_IN), .Z(U3349) );
  MUX2_X1 U4869 ( .A(n4267), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  MUX2_X1 U4870 ( .A(n4268), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  AOI22_X1 U4871 ( .A1(n4269), .A2(n4455), .B1(n4471), .B2(
        REG2_REG_31__SCAN_IN), .ZN(n4270) );
  OAI21_X1 U4872 ( .B1(n4471), .B2(n4271), .A(n4270), .ZN(U3260) );
  AOI22_X1 U4873 ( .A1(n4273), .A2(n4455), .B1(n3972), .B2(n4272), .ZN(n4274)
         );
  OAI21_X1 U4874 ( .B1(n4275), .B2(n3972), .A(n4274), .ZN(U3261) );
  OAI21_X1 U4875 ( .B1(REG1_REG_0__SCAN_IN), .B2(n4277), .A(n4276), .ZN(n4278)
         );
  XNOR2_X1 U4876 ( .A(n4278), .B(n4505), .ZN(n4281) );
  AOI22_X1 U4877 ( .A1(ADDR_REG_0__SCAN_IN), .A2(n4392), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n4279) );
  OAI21_X1 U4878 ( .B1(n4281), .B2(n4280), .A(n4279), .ZN(U3240) );
  AOI211_X1 U4879 ( .C1(n4284), .C2(n4283), .A(n4282), .B(n4293), .ZN(n4285)
         );
  AOI211_X1 U4880 ( .C1(n4392), .C2(ADDR_REG_5__SCAN_IN), .A(n4286), .B(n4285), 
        .ZN(n4291) );
  OAI211_X1 U4881 ( .C1(n4289), .C2(n4288), .A(n4346), .B(n4287), .ZN(n4290)
         );
  OAI211_X1 U4882 ( .C1(n4399), .C2(n4292), .A(n4291), .B(n4290), .ZN(U3245)
         );
  AOI211_X1 U4883 ( .C1(n4296), .C2(n4295), .A(n4294), .B(n4293), .ZN(n4297)
         );
  AOI211_X1 U4884 ( .C1(n4392), .C2(ADDR_REG_6__SCAN_IN), .A(n4298), .B(n4297), 
        .ZN(n4302) );
  OAI211_X1 U4885 ( .C1(REG2_REG_6__SCAN_IN), .C2(n4300), .A(n4346), .B(n4299), 
        .ZN(n4301) );
  OAI211_X1 U4886 ( .C1(n4399), .C2(n4501), .A(n4302), .B(n4301), .ZN(U3246)
         );
  OAI211_X1 U4887 ( .C1(n4305), .C2(n4304), .A(n4394), .B(n4303), .ZN(n4310)
         );
  OAI211_X1 U4888 ( .C1(n4308), .C2(n4307), .A(n4346), .B(n4306), .ZN(n4309)
         );
  OAI211_X1 U4889 ( .C1(n4399), .C2(n4499), .A(n4310), .B(n4309), .ZN(n4311)
         );
  AOI211_X1 U4890 ( .C1(n4392), .C2(ADDR_REG_9__SCAN_IN), .A(n4312), .B(n4311), 
        .ZN(n4313) );
  INV_X1 U4891 ( .A(n4313), .ZN(U3249) );
  OAI211_X1 U4892 ( .C1(REG1_REG_10__SCAN_IN), .C2(n4315), .A(n4394), .B(n4314), .ZN(n4319) );
  OAI211_X1 U4893 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4317), .A(n4346), .B(n4316), .ZN(n4318) );
  OAI211_X1 U4894 ( .C1(n4399), .C2(n4497), .A(n4319), .B(n4318), .ZN(n4320)
         );
  AOI211_X1 U4895 ( .C1(n4392), .C2(ADDR_REG_10__SCAN_IN), .A(n4321), .B(n4320), .ZN(n4322) );
  INV_X1 U4896 ( .A(n4322), .ZN(U3250) );
  OAI211_X1 U4897 ( .C1(n4325), .C2(n4324), .A(n4394), .B(n4323), .ZN(n4330)
         );
  OAI211_X1 U4898 ( .C1(n4328), .C2(n4327), .A(n4346), .B(n4326), .ZN(n4329)
         );
  OAI211_X1 U4899 ( .C1(n4399), .C2(n4331), .A(n4330), .B(n4329), .ZN(n4332)
         );
  AOI211_X1 U4900 ( .C1(n4392), .C2(ADDR_REG_11__SCAN_IN), .A(n4333), .B(n4332), .ZN(n4334) );
  INV_X1 U4901 ( .A(n4334), .ZN(U3251) );
  OAI211_X1 U4902 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4336), .A(n4346), .B(n4335), .ZN(n4337) );
  NAND2_X1 U4903 ( .A1(n4338), .A2(n4337), .ZN(n4339) );
  AOI21_X1 U4904 ( .B1(n4392), .B2(ADDR_REG_12__SCAN_IN), .A(n4339), .ZN(n4343) );
  OAI211_X1 U4905 ( .C1(REG1_REG_12__SCAN_IN), .C2(n4341), .A(n4394), .B(n4340), .ZN(n4342) );
  OAI211_X1 U4906 ( .C1(n4399), .C2(n2197), .A(n4343), .B(n4342), .ZN(U3252)
         );
  AOI21_X1 U4907 ( .B1(n4357), .B2(n4345), .A(n4344), .ZN(n4349) );
  OAI21_X1 U4908 ( .B1(n4349), .B2(n4348), .A(n4346), .ZN(n4347) );
  AOI21_X1 U4909 ( .B1(n4349), .B2(n4348), .A(n4347), .ZN(n4350) );
  AOI211_X1 U4910 ( .C1(n4392), .C2(ADDR_REG_13__SCAN_IN), .A(n4351), .B(n4350), .ZN(n4356) );
  OAI211_X1 U4911 ( .C1(n4354), .C2(n4353), .A(n4394), .B(n4352), .ZN(n4355)
         );
  OAI211_X1 U4912 ( .C1(n4399), .C2(n4357), .A(n4356), .B(n4355), .ZN(U3253)
         );
  AOI211_X1 U4913 ( .C1(n4360), .C2(n4359), .A(n4358), .B(n4387), .ZN(n4361)
         );
  AOI211_X1 U4914 ( .C1(n4392), .C2(ADDR_REG_15__SCAN_IN), .A(n4362), .B(n4361), .ZN(n4367) );
  OAI211_X1 U4915 ( .C1(n4365), .C2(n4364), .A(n4394), .B(n4363), .ZN(n4366)
         );
  OAI211_X1 U4916 ( .C1(n4399), .C2(n4490), .A(n4367), .B(n4366), .ZN(U3255)
         );
  AOI221_X1 U4917 ( .B1(n4369), .B2(n4368), .C1(n3932), .C2(n4368), .A(n4387), 
        .ZN(n4370) );
  AOI211_X1 U4918 ( .C1(n4392), .C2(ADDR_REG_16__SCAN_IN), .A(n4371), .B(n4370), .ZN(n4375) );
  OAI221_X1 U4919 ( .B1(n4373), .B2(REG1_REG_16__SCAN_IN), .C1(n4373), .C2(
        n4372), .A(n4394), .ZN(n4374) );
  OAI211_X1 U4920 ( .C1(n4399), .C2(n4488), .A(n4375), .B(n4374), .ZN(U3256)
         );
  AOI221_X1 U4921 ( .B1(n4378), .B2(n4377), .C1(n4376), .C2(n4377), .A(n4387), 
        .ZN(n4379) );
  AOI211_X1 U4922 ( .C1(n4392), .C2(ADDR_REG_17__SCAN_IN), .A(n4380), .B(n4379), .ZN(n4385) );
  OAI221_X1 U4923 ( .B1(n4383), .B2(n4382), .C1(n4383), .C2(n4381), .A(n4394), 
        .ZN(n4384) );
  OAI211_X1 U4924 ( .C1(n4399), .C2(n4386), .A(n4385), .B(n4384), .ZN(U3257)
         );
  AOI211_X1 U4925 ( .C1(n4389), .C2(n4388), .A(n2032), .B(n4387), .ZN(n4390)
         );
  AOI211_X1 U4926 ( .C1(n4392), .C2(ADDR_REG_18__SCAN_IN), .A(n4391), .B(n4390), .ZN(n4398) );
  OAI211_X1 U4927 ( .C1(n4396), .C2(n4395), .A(n4394), .B(n4393), .ZN(n4397)
         );
  OAI211_X1 U4928 ( .C1(n4399), .C2(n4484), .A(n4398), .B(n4397), .ZN(U3258)
         );
  XNOR2_X1 U4929 ( .A(n4400), .B(n4401), .ZN(n4556) );
  XNOR2_X1 U4930 ( .A(n4402), .B(n4401), .ZN(n4410) );
  OAI22_X1 U4931 ( .A1(n4404), .A2(n4464), .B1(n4417), .B2(n4403), .ZN(n4405)
         );
  AOI21_X1 U4932 ( .B1(n4407), .B2(n4406), .A(n4405), .ZN(n4408) );
  OAI21_X1 U4933 ( .B1(n4410), .B2(n4409), .A(n4408), .ZN(n4411) );
  AOI21_X1 U4934 ( .B1(n4462), .B2(n4556), .A(n4411), .ZN(n4553) );
  OAI22_X1 U4935 ( .A1(n4414), .A2(n4413), .B1(n4412), .B2(n3972), .ZN(n4415)
         );
  INV_X1 U4936 ( .A(n4415), .ZN(n4421) );
  OAI21_X1 U4937 ( .B1(n4418), .B2(n4417), .A(n4416), .ZN(n4552) );
  INV_X1 U4938 ( .A(n4552), .ZN(n4419) );
  AOI22_X1 U4939 ( .A1(n4556), .A2(n4467), .B1(n4455), .B2(n4419), .ZN(n4420)
         );
  OAI211_X1 U4940 ( .C1(n4471), .C2(n4553), .A(n4421), .B(n4420), .ZN(U3279)
         );
  AOI22_X1 U4941 ( .A1(n4422), .A2(n4466), .B1(REG2_REG_10__SCAN_IN), .B2(
        n4471), .ZN(n4427) );
  INV_X1 U4942 ( .A(n4423), .ZN(n4424) );
  AOI22_X1 U4943 ( .A1(n4425), .A2(n4467), .B1(n4455), .B2(n4424), .ZN(n4426)
         );
  OAI211_X1 U4944 ( .C1(n4471), .C2(n4428), .A(n4427), .B(n4426), .ZN(U3280)
         );
  AOI22_X1 U4945 ( .A1(n4429), .A2(n4466), .B1(REG2_REG_8__SCAN_IN), .B2(n4471), .ZN(n4434) );
  INV_X1 U4946 ( .A(n4430), .ZN(n4431) );
  AOI22_X1 U4947 ( .A1(n4432), .A2(n4467), .B1(n4455), .B2(n4431), .ZN(n4433)
         );
  OAI211_X1 U4948 ( .C1(n4471), .C2(n4435), .A(n4434), .B(n4433), .ZN(U3282)
         );
  INV_X1 U4949 ( .A(n4447), .ZN(n4438) );
  OAI21_X1 U4950 ( .B1(n4438), .B2(n4437), .A(n4436), .ZN(n4451) );
  AOI22_X1 U4951 ( .A1(n2751), .A2(n4441), .B1(n4440), .B2(n4439), .ZN(n4442)
         );
  OAI21_X1 U4952 ( .B1(n4444), .B2(n4443), .A(n4442), .ZN(n4450) );
  OAI21_X1 U4953 ( .B1(n4447), .B2(n4446), .A(n4445), .ZN(n4512) );
  NOR2_X1 U4954 ( .A1(n4512), .A2(n4448), .ZN(n4449) );
  AOI211_X1 U4955 ( .C1(n4461), .C2(n4451), .A(n4450), .B(n4449), .ZN(n4510)
         );
  AOI22_X1 U4956 ( .A1(REG3_REG_1__SCAN_IN), .A2(n4466), .B1(
        REG2_REG_1__SCAN_IN), .B2(n4471), .ZN(n4458) );
  INV_X1 U4957 ( .A(n4512), .ZN(n4456) );
  OAI21_X1 U4958 ( .B1(n4453), .B2(n4460), .A(n4452), .ZN(n4511) );
  INV_X1 U4959 ( .A(n4511), .ZN(n4454) );
  AOI22_X1 U4960 ( .A1(n4456), .A2(n4467), .B1(n4455), .B2(n4454), .ZN(n4457)
         );
  OAI211_X1 U4961 ( .C1(n4471), .C2(n4510), .A(n4458), .B(n4457), .ZN(U3289)
         );
  NOR2_X1 U4962 ( .A1(n4460), .A2(n4459), .ZN(n4507) );
  OAI21_X1 U4963 ( .B1(n4462), .B2(n4461), .A(n4508), .ZN(n4463) );
  OAI21_X1 U4964 ( .B1(n2749), .B2(n4464), .A(n4463), .ZN(n4506) );
  AOI21_X1 U4965 ( .B1(n4507), .B2(n4465), .A(n4506), .ZN(n4470) );
  AOI22_X1 U4966 ( .A1(n4467), .A2(n4508), .B1(REG3_REG_0__SCAN_IN), .B2(n4466), .ZN(n4468) );
  OAI221_X1 U4967 ( .B1(n4471), .B2(n4470), .C1(n3972), .C2(n4469), .A(n4468), 
        .ZN(U3290) );
  NOR2_X1 U4968 ( .A1(n4479), .A2(n4472), .ZN(U3291) );
  NOR2_X1 U4969 ( .A1(n4479), .A2(n4473), .ZN(U3292) );
  AND2_X1 U4970 ( .A1(D_REG_29__SCAN_IN), .A2(n4480), .ZN(U3293) );
  AND2_X1 U4971 ( .A1(D_REG_28__SCAN_IN), .A2(n4480), .ZN(U3294) );
  AND2_X1 U4972 ( .A1(D_REG_27__SCAN_IN), .A2(n4480), .ZN(U3295) );
  AND2_X1 U4973 ( .A1(D_REG_26__SCAN_IN), .A2(n4480), .ZN(U3296) );
  AND2_X1 U4974 ( .A1(D_REG_25__SCAN_IN), .A2(n4480), .ZN(U3297) );
  NOR2_X1 U4975 ( .A1(n4479), .A2(n4474), .ZN(U3298) );
  AND2_X1 U4976 ( .A1(D_REG_23__SCAN_IN), .A2(n4480), .ZN(U3299) );
  AND2_X1 U4977 ( .A1(D_REG_22__SCAN_IN), .A2(n4480), .ZN(U3300) );
  AND2_X1 U4978 ( .A1(D_REG_21__SCAN_IN), .A2(n4480), .ZN(U3301) );
  NOR2_X1 U4979 ( .A1(n4479), .A2(n4475), .ZN(U3302) );
  AND2_X1 U4980 ( .A1(D_REG_19__SCAN_IN), .A2(n4480), .ZN(U3303) );
  AND2_X1 U4981 ( .A1(D_REG_18__SCAN_IN), .A2(n4480), .ZN(U3304) );
  NOR2_X1 U4982 ( .A1(n4479), .A2(n4476), .ZN(U3305) );
  AND2_X1 U4983 ( .A1(D_REG_16__SCAN_IN), .A2(n4480), .ZN(U3306) );
  AND2_X1 U4984 ( .A1(D_REG_15__SCAN_IN), .A2(n4480), .ZN(U3307) );
  AND2_X1 U4985 ( .A1(D_REG_14__SCAN_IN), .A2(n4480), .ZN(U3308) );
  AND2_X1 U4986 ( .A1(D_REG_13__SCAN_IN), .A2(n4480), .ZN(U3309) );
  NOR2_X1 U4987 ( .A1(n4479), .A2(n4477), .ZN(U3310) );
  AND2_X1 U4988 ( .A1(D_REG_11__SCAN_IN), .A2(n4480), .ZN(U3311) );
  AND2_X1 U4989 ( .A1(D_REG_10__SCAN_IN), .A2(n4480), .ZN(U3312) );
  AND2_X1 U4990 ( .A1(D_REG_9__SCAN_IN), .A2(n4480), .ZN(U3313) );
  AND2_X1 U4991 ( .A1(D_REG_8__SCAN_IN), .A2(n4480), .ZN(U3314) );
  AND2_X1 U4992 ( .A1(D_REG_7__SCAN_IN), .A2(n4480), .ZN(U3315) );
  AND2_X1 U4993 ( .A1(D_REG_6__SCAN_IN), .A2(n4480), .ZN(U3316) );
  AND2_X1 U4994 ( .A1(D_REG_5__SCAN_IN), .A2(n4480), .ZN(U3317) );
  AND2_X1 U4995 ( .A1(D_REG_4__SCAN_IN), .A2(n4480), .ZN(U3318) );
  NOR2_X1 U4996 ( .A1(n4479), .A2(n4478), .ZN(U3319) );
  AND2_X1 U4997 ( .A1(D_REG_2__SCAN_IN), .A2(n4480), .ZN(U3320) );
  AOI21_X1 U4998 ( .B1(U3149), .B2(n4482), .A(n4481), .ZN(U3329) );
  INV_X1 U4999 ( .A(DATAI_18_), .ZN(n4483) );
  AOI22_X1 U5000 ( .A1(STATE_REG_SCAN_IN), .A2(n4484), .B1(n4483), .B2(U3149), 
        .ZN(U3334) );
  OAI22_X1 U5001 ( .A1(U3149), .A2(n4485), .B1(DATAI_17_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4486) );
  INV_X1 U5002 ( .A(n4486), .ZN(U3335) );
  INV_X1 U5003 ( .A(DATAI_16_), .ZN(n4487) );
  AOI22_X1 U5004 ( .A1(STATE_REG_SCAN_IN), .A2(n4488), .B1(n4487), .B2(U3149), 
        .ZN(U3336) );
  INV_X1 U5005 ( .A(DATAI_15_), .ZN(n4489) );
  AOI22_X1 U5006 ( .A1(STATE_REG_SCAN_IN), .A2(n4490), .B1(n4489), .B2(U3149), 
        .ZN(U3337) );
  OAI22_X1 U5007 ( .A1(U3149), .A2(n4491), .B1(DATAI_13_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4492) );
  INV_X1 U5008 ( .A(n4492), .ZN(U3339) );
  INV_X1 U5009 ( .A(DATAI_12_), .ZN(n4493) );
  AOI22_X1 U5010 ( .A1(STATE_REG_SCAN_IN), .A2(n2197), .B1(n4493), .B2(U3149), 
        .ZN(U3340) );
  OAI22_X1 U5011 ( .A1(U3149), .A2(n4494), .B1(DATAI_11_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4495) );
  INV_X1 U5012 ( .A(n4495), .ZN(U3341) );
  AOI22_X1 U5013 ( .A1(STATE_REG_SCAN_IN), .A2(n4497), .B1(n4496), .B2(U3149), 
        .ZN(U3342) );
  INV_X1 U5014 ( .A(DATAI_9_), .ZN(n4498) );
  AOI22_X1 U5015 ( .A1(STATE_REG_SCAN_IN), .A2(n4499), .B1(n4498), .B2(U3149), 
        .ZN(U3343) );
  INV_X1 U5016 ( .A(DATAI_6_), .ZN(n4500) );
  AOI22_X1 U5017 ( .A1(STATE_REG_SCAN_IN), .A2(n4501), .B1(n4500), .B2(U3149), 
        .ZN(U3346) );
  OAI22_X1 U5018 ( .A1(U3149), .A2(n4502), .B1(DATAI_5_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4503) );
  INV_X1 U5019 ( .A(n4503), .ZN(U3347) );
  AOI22_X1 U5020 ( .A1(STATE_REG_SCAN_IN), .A2(n4505), .B1(n4504), .B2(U3149), 
        .ZN(U3352) );
  AOI211_X1 U5021 ( .C1(n4557), .C2(n4508), .A(n4507), .B(n4506), .ZN(n4561)
         );
  INV_X1 U5022 ( .A(REG0_REG_0__SCAN_IN), .ZN(n4509) );
  AOI22_X1 U5023 ( .A1(n4560), .A2(n4561), .B1(n4509), .B2(n4558), .ZN(U3467)
         );
  INV_X1 U5024 ( .A(n4510), .ZN(n4514) );
  OAI22_X1 U5025 ( .A1(n4512), .A2(n4524), .B1(n2841), .B2(n4511), .ZN(n4513)
         );
  NOR2_X1 U5026 ( .A1(n4514), .A2(n4513), .ZN(n4563) );
  INV_X1 U5027 ( .A(REG0_REG_1__SCAN_IN), .ZN(n4515) );
  AOI22_X1 U5028 ( .A1(n4560), .A2(n4563), .B1(n4515), .B2(n4558), .ZN(U3469)
         );
  NOR3_X1 U5029 ( .A1(n4517), .A2(n4516), .A3(n2841), .ZN(n4520) );
  INV_X1 U5030 ( .A(n4518), .ZN(n4519) );
  AOI211_X1 U5031 ( .C1(n4557), .C2(n4521), .A(n4520), .B(n4519), .ZN(n4565)
         );
  INV_X1 U5032 ( .A(REG0_REG_2__SCAN_IN), .ZN(n4522) );
  AOI22_X1 U5033 ( .A1(n4560), .A2(n4565), .B1(n4522), .B2(n4558), .ZN(U3471)
         );
  OAI22_X1 U5034 ( .A1(n4525), .A2(n4524), .B1(n2841), .B2(n4523), .ZN(n4526)
         );
  NOR2_X1 U5035 ( .A1(n4527), .A2(n4526), .ZN(n4567) );
  INV_X1 U5036 ( .A(REG0_REG_3__SCAN_IN), .ZN(n4528) );
  AOI22_X1 U5037 ( .A1(n4560), .A2(n4567), .B1(n4528), .B2(n4558), .ZN(U3473)
         );
  NAND2_X1 U5038 ( .A1(n4529), .A2(n4557), .ZN(n4531) );
  NAND2_X1 U5039 ( .A1(n4531), .A2(n4530), .ZN(n4532) );
  NOR2_X1 U5040 ( .A1(n4533), .A2(n4532), .ZN(n4569) );
  INV_X1 U5041 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4534) );
  AOI22_X1 U5042 ( .A1(n4560), .A2(n4569), .B1(n4534), .B2(n4558), .ZN(U3475)
         );
  NOR2_X1 U5043 ( .A1(n4536), .A2(n4535), .ZN(n4538) );
  AOI211_X1 U5044 ( .C1(n4540), .C2(n4539), .A(n4538), .B(n4537), .ZN(n4571)
         );
  INV_X1 U5045 ( .A(REG0_REG_5__SCAN_IN), .ZN(n4541) );
  AOI22_X1 U5046 ( .A1(n4560), .A2(n4571), .B1(n4541), .B2(n4558), .ZN(U3477)
         );
  AOI211_X1 U5047 ( .C1(n4544), .C2(n4550), .A(n4543), .B(n4542), .ZN(n4573)
         );
  INV_X1 U5048 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4545) );
  AOI22_X1 U5049 ( .A1(n4560), .A2(n4573), .B1(n4545), .B2(n4558), .ZN(U3481)
         );
  OAI21_X1 U5050 ( .B1(n2841), .B2(n4547), .A(n4546), .ZN(n4548) );
  AOI21_X1 U5051 ( .B1(n4550), .B2(n4549), .A(n4548), .ZN(n4575) );
  AOI22_X1 U5052 ( .A1(n4560), .A2(n4575), .B1(n4551), .B2(n4558), .ZN(U3485)
         );
  NOR2_X1 U5053 ( .A1(n4552), .A2(n2841), .ZN(n4555) );
  INV_X1 U5054 ( .A(n4553), .ZN(n4554) );
  AOI211_X1 U5055 ( .C1(n4557), .C2(n4556), .A(n4555), .B(n4554), .ZN(n4578)
         );
  INV_X1 U5056 ( .A(REG0_REG_11__SCAN_IN), .ZN(n4559) );
  AOI22_X1 U5057 ( .A1(n4560), .A2(n4578), .B1(n4559), .B2(n4558), .ZN(U3489)
         );
  AOI22_X1 U5058 ( .A1(n4579), .A2(n4561), .B1(n2309), .B2(n4576), .ZN(U3518)
         );
  AOI22_X1 U5059 ( .A1(n4579), .A2(n4563), .B1(n4562), .B2(n4576), .ZN(U3519)
         );
  AOI22_X1 U5060 ( .A1(n4579), .A2(n4565), .B1(n4564), .B2(n4576), .ZN(U3520)
         );
  AOI22_X1 U5061 ( .A1(n4579), .A2(n4567), .B1(n4566), .B2(n4576), .ZN(U3521)
         );
  INV_X1 U5062 ( .A(REG1_REG_4__SCAN_IN), .ZN(n4568) );
  AOI22_X1 U5063 ( .A1(n4579), .A2(n4569), .B1(n4568), .B2(n4576), .ZN(U3522)
         );
  AOI22_X1 U5064 ( .A1(n4579), .A2(n4571), .B1(n4570), .B2(n4576), .ZN(U3523)
         );
  AOI22_X1 U5065 ( .A1(n4579), .A2(n4573), .B1(n4572), .B2(n4576), .ZN(U3525)
         );
  AOI22_X1 U5066 ( .A1(n4579), .A2(n4575), .B1(n4574), .B2(n4576), .ZN(U3527)
         );
  AOI22_X1 U5067 ( .A1(n4579), .A2(n4578), .B1(n4577), .B2(n4576), .ZN(U3529)
         );
endmodule

