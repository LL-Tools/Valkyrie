

module b14_C_2inp_gates_syn ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, U3352, U3351, U3350, U3349, 
        U3348, U3347, U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, 
        U3338, U3337, U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, 
        U3328, U3327, U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, 
        U3320, U3319, U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, 
        U3310, U3309, U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, 
        U3300, U3299, U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, 
        U3467, U3469, U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, 
        U3487, U3489, U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, 
        U3506, U3507, U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, 
        U3516, U3517, U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, 
        U3526, U3527, U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, 
        U3536, U3537, U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, 
        U3546, U3547, U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, 
        U3284, U3283, U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, 
        U3274, U3273, U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, 
        U3264, U3263, U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, 
        U3255, U3254, U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, 
        U3245, U3244, U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, 
        U3554, U3555, U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, 
        U3564, U3565, U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, 
        U3574, U3575, U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, 
        U3237, U3236, U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, 
        U3227, U3226, U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, 
        U3217, U3216, U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, 
        U4043, keyinput127, keyinput126, keyinput125, keyinput124, keyinput123, 
        keyinput122, keyinput121, keyinput120, keyinput119, keyinput118, 
        keyinput117, keyinput116, keyinput115, keyinput114, keyinput113, 
        keyinput112, keyinput111, keyinput110, keyinput109, keyinput108, 
        keyinput107, keyinput106, keyinput105, keyinput104, keyinput103, 
        keyinput102, keyinput101, keyinput100, keyinput99, keyinput98, 
        keyinput97, keyinput96, keyinput95, keyinput94, keyinput93, keyinput92, 
        keyinput91, keyinput90, keyinput89, keyinput88, keyinput87, keyinput86, 
        keyinput85, keyinput84, keyinput83, keyinput82, keyinput81, keyinput80, 
        keyinput79, keyinput78, keyinput77, keyinput76, keyinput75, keyinput74, 
        keyinput73, keyinput72, keyinput71, keyinput70, keyinput69, keyinput68, 
        keyinput67, keyinput66, keyinput65, keyinput64, keyinput63, keyinput62, 
        keyinput61, keyinput60, keyinput59, keyinput58, keyinput57, keyinput56, 
        keyinput55, keyinput54, keyinput53, keyinput52, keyinput51, keyinput50, 
        keyinput49, keyinput48, keyinput47, keyinput46, keyinput45, keyinput44, 
        keyinput43, keyinput42, keyinput41, keyinput40, keyinput39, keyinput38, 
        keyinput37, keyinput36, keyinput35, keyinput34, keyinput33, keyinput32, 
        keyinput31, keyinput30, keyinput29, keyinput28, keyinput27, keyinput26, 
        keyinput25, keyinput24, keyinput23, keyinput22, keyinput21, keyinput20, 
        keyinput19, keyinput18, keyinput17, keyinput16, keyinput15, keyinput14, 
        keyinput13, keyinput12, keyinput11, keyinput10, keyinput9, keyinput8, 
        keyinput7, keyinput6, keyinput5, keyinput4, keyinput3, keyinput2, 
        keyinput1, keyinput0 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput127, keyinput126, keyinput125,
         keyinput124, keyinput123, keyinput122, keyinput121, keyinput120,
         keyinput119, keyinput118, keyinput117, keyinput116, keyinput115,
         keyinput114, keyinput113, keyinput112, keyinput111, keyinput110,
         keyinput109, keyinput108, keyinput107, keyinput106, keyinput105,
         keyinput104, keyinput103, keyinput102, keyinput101, keyinput100,
         keyinput99, keyinput98, keyinput97, keyinput96, keyinput95,
         keyinput94, keyinput93, keyinput92, keyinput91, keyinput90,
         keyinput89, keyinput88, keyinput87, keyinput86, keyinput85,
         keyinput84, keyinput83, keyinput82, keyinput81, keyinput80,
         keyinput79, keyinput78, keyinput77, keyinput76, keyinput75,
         keyinput74, keyinput73, keyinput72, keyinput71, keyinput70,
         keyinput69, keyinput68, keyinput67, keyinput66, keyinput65,
         keyinput64, keyinput63, keyinput62, keyinput61, keyinput60,
         keyinput59, keyinput58, keyinput57, keyinput56, keyinput55,
         keyinput54, keyinput53, keyinput52, keyinput51, keyinput50,
         keyinput49, keyinput48, keyinput47, keyinput46, keyinput45,
         keyinput44, keyinput43, keyinput42, keyinput41, keyinput40,
         keyinput39, keyinput38, keyinput37, keyinput36, keyinput35,
         keyinput34, keyinput33, keyinput32, keyinput31, keyinput30,
         keyinput29, keyinput28, keyinput27, keyinput26, keyinput25,
         keyinput24, keyinput23, keyinput22, keyinput21, keyinput20,
         keyinput19, keyinput18, keyinput17, keyinput16, keyinput15,
         keyinput14, keyinput13, keyinput12, keyinput11, keyinput10, keyinput9,
         keyinput8, keyinput7, keyinput6, keyinput5, keyinput4, keyinput3,
         keyinput2, keyinput1, keyinput0;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
         n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
         n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
         n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
         n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872;

  OAI21_X1 U2374 ( .B1(n4403), .B2(n2301), .A(n2300), .ZN(n4411) );
  INV_X2 U2375 ( .A(n3530), .ZN(n3487) );
  AND2_X1 U2376 ( .A1(n2298), .A2(n2150), .ZN(n4394) );
  NAND2_X1 U2377 ( .A1(n4130), .A2(n2594), .ZN(n4103) );
  CLKBUF_X3 U2378 ( .A(n2405), .Z(n3684) );
  NAND3_X1 U2379 ( .A1(n4353), .A2(n4355), .A3(n4354), .ZN(n2891) );
  NAND2_X1 U2380 ( .A1(n2896), .A2(n4534), .ZN(n3455) );
  INV_X1 U2381 ( .A(n3455), .ZN(n3533) );
  CLKBUF_X3 U2382 ( .A(n3533), .Z(n2135) );
  INV_X2 U2383 ( .A(n3276), .ZN(n2133) );
  NOR2_X2 U2384 ( .A1(n4431), .A2(n2304), .ZN(n3895) );
  AOI21_X2 U2385 ( .B1(n3512), .B2(n3437), .A(n3436), .ZN(n3556) );
  OAI21_X2 U2386 ( .B1(n3591), .B2(n3594), .A(n3592), .ZN(n3512) );
  OAI21_X2 U2387 ( .B1(n3218), .B2(n3243), .A(n2515), .ZN(n3245) );
  OAI21_X2 U2388 ( .B1(n3189), .B2(n2497), .A(n2496), .ZN(n3218) );
  XNOR2_X2 U2389 ( .A(n2822), .B(n2813), .ZN(n2821) );
  AOI21_X2 U2391 ( .B1(n3901), .B2(REG1_REG_11__SCAN_IN), .A(n4392), .ZN(n3890) );
  OR2_X1 U2392 ( .A1(n2761), .A2(n2751), .ZN(n2316) );
  AOI22_X1 U2393 ( .A1(n3931), .A2(n3930), .B1(n3929), .B2(n3938), .ZN(n3932)
         );
  XNOR2_X1 U2394 ( .A(n3931), .B(n3930), .ZN(n3387) );
  NAND2_X1 U2395 ( .A1(n2650), .A2(n2331), .ZN(n2330) );
  AND2_X1 U2396 ( .A1(n3723), .A2(n2418), .ZN(n2328) );
  NAND2_X1 U2397 ( .A1(n3762), .A2(n3765), .ZN(n3723) );
  CLKBUF_X2 U2398 ( .A(n2911), .Z(n3532) );
  NAND2_X2 U2399 ( .A1(n3756), .A2(n3759), .ZN(n3722) );
  INV_X2 U2400 ( .A(n3445), .ZN(n2896) );
  OR2_X1 U2401 ( .A1(n2794), .A2(n2421), .ZN(n2430) );
  INV_X1 U2402 ( .A(n3842), .ZN(n2385) );
  NAND2_X2 U2403 ( .A1(n2676), .A2(n2708), .ZN(n2892) );
  NAND2_X1 U2404 ( .A1(n4352), .A2(n2387), .ZN(n2405) );
  NAND2_X1 U2405 ( .A1(n4352), .A2(n2367), .ZN(n2423) );
  OAI21_X1 U2407 ( .B1(n2761), .B2(n4541), .A(n2205), .ZN(n2763) );
  AND2_X1 U2408 ( .A1(n2330), .A2(n2333), .ZN(n3953) );
  NAND2_X1 U2409 ( .A1(n2330), .A2(n2329), .ZN(n2663) );
  AOI21_X2 U2410 ( .B1(n3421), .B2(n3420), .A(n3419), .ZN(n3591) );
  OR2_X1 U2411 ( .A1(n3378), .A2(n4302), .ZN(n2757) );
  OR2_X1 U2412 ( .A1(n4384), .A2(n2499), .ZN(n2298) );
  NOR2_X1 U2413 ( .A1(n3888), .A2(n2160), .ZN(n3889) );
  NOR2_X1 U2414 ( .A1(n2655), .A2(n2162), .ZN(n2329) );
  NAND2_X1 U2415 ( .A1(n2751), .A2(n2664), .ZN(n2315) );
  NOR2_X1 U2416 ( .A1(n2279), .A2(n2275), .ZN(n2274) );
  OAI21_X1 U2417 ( .B1(n2855), .B2(n2834), .A(n2836), .ZN(n2880) );
  OAI21_X2 U2418 ( .B1(n2934), .B2(n4275), .A(n4169), .ZN(n2935) );
  AND2_X1 U2419 ( .A1(n2684), .A2(n3776), .ZN(n3768) );
  XNOR2_X1 U2420 ( .A(n2831), .B(n2848), .ZN(n2846) );
  NAND2_X1 U2421 ( .A1(n2867), .A2(n2830), .ZN(n2831) );
  NAND2_X1 U2422 ( .A1(n2756), .A2(n2755), .ZN(n4534) );
  INV_X2 U2423 ( .A(n3276), .ZN(n2911) );
  NAND2_X1 U2424 ( .A1(n2146), .A2(n2412), .ZN(n2890) );
  OR2_X2 U2425 ( .A1(n2892), .A2(n2902), .ZN(n3276) );
  NAND2_X2 U2426 ( .A1(n2892), .A2(n2936), .ZN(n3530) );
  BUF_X2 U2427 ( .A(n2410), .Z(n2411) );
  INV_X2 U2428 ( .A(n3856), .ZN(U4043) );
  INV_X4 U2429 ( .A(n3677), .ZN(n3679) );
  XNOR2_X1 U2430 ( .A(n2364), .B(IR_REG_30__SCAN_IN), .ZN(n2367) );
  AND2_X1 U2431 ( .A1(n2379), .A2(n2378), .ZN(n3677) );
  NAND2_X1 U2432 ( .A1(n2769), .A2(IR_REG_31__SCAN_IN), .ZN(n2364) );
  NAND2_X1 U2433 ( .A1(n2185), .A2(IR_REG_31__SCAN_IN), .ZN(n2374) );
  NAND2_X1 U2434 ( .A1(n2725), .A2(IR_REG_31__SCAN_IN), .ZN(n2731) );
  AND3_X1 U2435 ( .A1(n2323), .A2(n2296), .A3(n2346), .ZN(n2545) );
  AND2_X1 U2436 ( .A1(n2297), .A2(n2347), .ZN(n2296) );
  INV_X1 U2437 ( .A(n2136), .ZN(n2334) );
  NOR2_X1 U2438 ( .A1(n2350), .A2(IR_REG_10__SCAN_IN), .ZN(n2297) );
  AND2_X1 U2439 ( .A1(n2340), .A2(n2154), .ZN(n2323) );
  NAND2_X1 U2440 ( .A1(n4821), .A2(n2349), .ZN(n2350) );
  INV_X1 U2441 ( .A(IR_REG_12__SCAN_IN), .ZN(n2349) );
  INV_X1 U2442 ( .A(IR_REG_14__SCAN_IN), .ZN(n4608) );
  INV_X1 U2443 ( .A(IR_REG_19__SCAN_IN), .ZN(n2216) );
  INV_X1 U2444 ( .A(IR_REG_18__SCAN_IN), .ZN(n2602) );
  INV_X1 U2445 ( .A(IR_REG_21__SCAN_IN), .ZN(n2721) );
  INV_X1 U2446 ( .A(IR_REG_4__SCAN_IN), .ZN(n2433) );
  INV_X1 U2447 ( .A(IR_REG_5__SCAN_IN), .ZN(n2326) );
  INV_X1 U2448 ( .A(IR_REG_3__SCAN_IN), .ZN(n2414) );
  NOR2_X2 U2449 ( .A1(IR_REG_0__SCAN_IN), .A2(IR_REG_1__SCAN_IN), .ZN(n2399)
         );
  INV_X1 U2450 ( .A(IR_REG_11__SCAN_IN), .ZN(n4821) );
  AOI21_X2 U2451 ( .B1(n3912), .B2(REG1_REG_13__SCAN_IN), .A(n4411), .ZN(n3893) );
  XNOR2_X1 U2452 ( .A(n2180), .B(IR_REG_2__SCAN_IN), .ZN(n3872) );
  XNOR2_X2 U2453 ( .A(n2722), .B(n2721), .ZN(n2708) );
  AND3_X1 U2454 ( .A1(n2323), .A2(n2346), .A3(n2181), .ZN(n2183) );
  AND2_X1 U2455 ( .A1(n2347), .A2(n2182), .ZN(n2181) );
  AND2_X1 U2456 ( .A1(n2348), .A2(n2356), .ZN(n2182) );
  AND2_X1 U2457 ( .A1(n3402), .A2(n2287), .ZN(n2282) );
  INV_X1 U2458 ( .A(n3771), .ZN(n2204) );
  OR2_X1 U2459 ( .A1(n3841), .A2(n2952), .ZN(n3756) );
  OR2_X1 U2460 ( .A1(n2771), .A2(n2745), .ZN(n2924) );
  NAND2_X1 U2461 ( .A1(n2336), .A2(n4814), .ZN(n2335) );
  INV_X1 U2462 ( .A(n2350), .ZN(n2336) );
  INV_X1 U2463 ( .A(IR_REG_23__SCAN_IN), .ZN(n2730) );
  INV_X1 U2464 ( .A(IR_REG_9__SCAN_IN), .ZN(n2324) );
  NAND2_X1 U2465 ( .A1(n2399), .A2(n2400), .ZN(n2413) );
  INV_X1 U2466 ( .A(n3554), .ZN(n2255) );
  AND2_X1 U2467 ( .A1(n2708), .A2(n4356), .ZN(n2927) );
  NAND2_X1 U2468 ( .A1(n2802), .A2(n2236), .ZN(n3869) );
  NOR2_X1 U2469 ( .A1(n2332), .A2(n2342), .ZN(n2331) );
  INV_X1 U2470 ( .A(n2649), .ZN(n2332) );
  OR2_X1 U2471 ( .A1(n2311), .A2(n2635), .ZN(n2309) );
  AND2_X1 U2472 ( .A1(n2312), .A2(n2339), .ZN(n2311) );
  OR2_X1 U2473 ( .A1(n4055), .A2(n2313), .ZN(n2312) );
  NAND2_X1 U2474 ( .A1(n4143), .A2(n2581), .ZN(n2327) );
  OR2_X1 U2475 ( .A1(n3642), .A2(n3598), .ZN(n2581) );
  XNOR2_X1 U2476 ( .A(n3935), .B(n3930), .ZN(n2715) );
  AND2_X1 U2477 ( .A1(n4368), .A2(n2927), .ZN(n4289) );
  AND2_X1 U2478 ( .A1(n2710), .A2(n2358), .ZN(n2359) );
  NAND2_X1 U2479 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_28__SCAN_IN), .ZN(n2358) );
  INV_X1 U2480 ( .A(n2473), .ZN(n2321) );
  INV_X1 U2481 ( .A(n3816), .ZN(n2194) );
  NAND2_X1 U2482 ( .A1(n2149), .A2(n3527), .ZN(n2262) );
  INV_X1 U2483 ( .A(n3528), .ZN(n2263) );
  AOI21_X1 U2484 ( .B1(n2284), .B2(n3402), .A(n2170), .ZN(n2283) );
  INV_X1 U2485 ( .A(n2285), .ZN(n2284) );
  AND2_X1 U2486 ( .A1(n4440), .A2(REG1_REG_15__SCAN_IN), .ZN(n2304) );
  INV_X1 U2487 ( .A(n3987), .ZN(n2197) );
  OAI21_X1 U2488 ( .B1(n2309), .B2(n2155), .A(n2142), .ZN(n2307) );
  OR2_X1 U2489 ( .A1(n4105), .A2(n4024), .ZN(n4080) );
  AOI21_X1 U2490 ( .B1(n4164), .B2(n2191), .A(n2190), .ZN(n2189) );
  INV_X1 U2491 ( .A(n3689), .ZN(n2191) );
  AOI21_X1 U2492 ( .B1(n2203), .B2(n2202), .A(n2201), .ZN(n2200) );
  INV_X1 U2493 ( .A(n3776), .ZN(n2202) );
  INV_X1 U2494 ( .A(n3775), .ZN(n2201) );
  NAND2_X1 U2495 ( .A1(n2199), .A2(n2203), .ZN(n2198) );
  NAND2_X1 U2496 ( .A1(n2215), .A2(n3764), .ZN(n2211) );
  NAND2_X1 U2497 ( .A1(n3764), .A2(n2210), .ZN(n2209) );
  AND2_X1 U2498 ( .A1(n2682), .A2(n3765), .ZN(n2210) );
  AND2_X1 U2499 ( .A1(n3722), .A2(n2392), .ZN(n2322) );
  INV_X1 U2500 ( .A(n3111), .ZN(n2278) );
  NOR2_X1 U2501 ( .A1(n3110), .A2(n3111), .ZN(n2279) );
  INV_X1 U2502 ( .A(n3580), .ZN(n2275) );
  INV_X1 U2503 ( .A(n3048), .ZN(n2280) );
  AOI21_X1 U2504 ( .B1(n2268), .B2(n2267), .A(n2157), .ZN(n2266) );
  INV_X1 U2505 ( .A(n2164), .ZN(n2267) );
  AND2_X1 U2506 ( .A1(n3014), .A2(n3012), .ZN(n2291) );
  NAND2_X1 U2507 ( .A1(n3304), .A2(n3303), .ZN(n2294) );
  OR2_X1 U2508 ( .A1(n3304), .A2(n3303), .ZN(n2295) );
  NAND2_X1 U2509 ( .A1(n2252), .A2(n2253), .ZN(n2257) );
  AND2_X1 U2510 ( .A1(n2943), .A2(n2932), .ZN(n3366) );
  NAND2_X1 U2511 ( .A1(n2133), .A2(n3842), .ZN(n2909) );
  AOI22_X1 U2512 ( .A1(n3841), .A2(n3533), .B1(n3368), .B2(n2911), .ZN(n2922)
         );
  NAND2_X1 U2513 ( .A1(n2917), .A2(n2916), .ZN(n2918) );
  NAND2_X1 U2514 ( .A1(n2271), .A2(n2272), .ZN(n2270) );
  NAND2_X1 U2515 ( .A1(n2366), .A2(n2387), .ZN(n2420) );
  NAND2_X1 U2516 ( .A1(n3845), .A2(n2800), .ZN(n2236) );
  NAND2_X1 U2517 ( .A1(n2242), .A2(n2816), .ZN(n2817) );
  NAND2_X1 U2518 ( .A1(n2814), .A2(REG2_REG_3__SCAN_IN), .ZN(n2242) );
  XNOR2_X1 U2519 ( .A(n2817), .B(n3877), .ZN(n2818) );
  NAND2_X1 U2520 ( .A1(n2179), .A2(n2178), .ZN(n2244) );
  NAND2_X1 U2521 ( .A1(n2820), .A2(n4362), .ZN(n2178) );
  NAND2_X1 U2522 ( .A1(n2845), .A2(REG2_REG_6__SCAN_IN), .ZN(n2179) );
  XNOR2_X1 U2523 ( .A(n3889), .B(n2299), .ZN(n4384) );
  XNOR2_X1 U2524 ( .A(n3895), .B(n2303), .ZN(n4451) );
  NAND2_X1 U2525 ( .A1(n4451), .A2(n4450), .ZN(n4449) );
  NAND2_X1 U2526 ( .A1(n2171), .A2(n4459), .ZN(n2173) );
  INV_X1 U2527 ( .A(n4447), .ZN(n2171) );
  INV_X1 U2528 ( .A(n2175), .ZN(n2174) );
  OAI21_X1 U2529 ( .B1(n3917), .B2(n2176), .A(n2241), .ZN(n2175) );
  OR2_X1 U2530 ( .A1(n3918), .A2(REG2_REG_17__SCAN_IN), .ZN(n2241) );
  NAND3_X1 U2531 ( .A1(n2173), .A2(n2172), .A3(n2174), .ZN(n2240) );
  INV_X1 U2532 ( .A(n4480), .ZN(n2172) );
  NAND2_X1 U2533 ( .A1(n3947), .A2(n3946), .ZN(n4201) );
  NAND2_X1 U2534 ( .A1(n2197), .A2(n2196), .ZN(n3968) );
  AND2_X1 U2535 ( .A1(n2706), .A2(n2707), .ZN(n3960) );
  AND2_X1 U2536 ( .A1(n2642), .A2(REG3_REG_25__SCAN_IN), .ZN(n2657) );
  OR2_X1 U2537 ( .A1(n3973), .A2(n2234), .ZN(n2648) );
  NAND2_X1 U2538 ( .A1(n2314), .A2(n2627), .ZN(n2310) );
  OR2_X1 U2539 ( .A1(n4245), .A2(n4074), .ZN(n4069) );
  AND2_X1 U2540 ( .A1(n3631), .A2(n4238), .ZN(n2620) );
  NAND2_X1 U2541 ( .A1(n4049), .A2(n4055), .ZN(n4048) );
  NAND2_X1 U2542 ( .A1(n2327), .A2(n2161), .ZN(n4130) );
  OR2_X1 U2543 ( .A1(n4185), .A2(n4184), .ZN(n4188) );
  INV_X1 U2544 ( .A(n3117), .ZN(n3127) );
  INV_X1 U2545 ( .A(n4187), .ZN(n4167) );
  NAND2_X1 U2546 ( .A1(n3676), .A2(n2709), .ZN(n4162) );
  NAND2_X1 U2547 ( .A1(n3366), .A2(n2924), .ZN(n2966) );
  NOR3_X1 U2548 ( .A1(n4069), .A2(n2232), .A3(n2234), .ZN(n3995) );
  NOR2_X1 U2549 ( .A1(n4069), .A2(n2232), .ZN(n4010) );
  NAND2_X1 U2550 ( .A1(n4554), .A2(n4508), .ZN(n4527) );
  NAND2_X1 U2551 ( .A1(n2735), .A2(n4353), .ZN(n2771) );
  INV_X1 U2552 ( .A(IR_REG_27__SCAN_IN), .ZN(n2377) );
  NAND2_X1 U2553 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_27__SCAN_IN), .ZN(n2710) );
  NOR2_X1 U2554 ( .A1(n2335), .A2(n2355), .ZN(n2143) );
  INV_X1 U2555 ( .A(IR_REG_25__SCAN_IN), .ZN(n2728) );
  NAND2_X1 U2556 ( .A1(n2731), .A2(n2730), .ZN(n2733) );
  AND2_X1 U2557 ( .A1(n2347), .A2(n2348), .ZN(n2186) );
  INV_X2 U2558 ( .A(n2413), .ZN(n2346) );
  NAND2_X1 U2559 ( .A1(n3619), .A2(n2287), .ZN(n2286) );
  AND2_X1 U2560 ( .A1(n2254), .A2(n2251), .ZN(n2250) );
  NAND2_X1 U2561 ( .A1(n2258), .A2(n3611), .ZN(n2251) );
  NAND2_X1 U2562 ( .A1(n2938), .A2(n4368), .ZN(n3653) );
  INV_X1 U2563 ( .A(n2935), .ZN(n3668) );
  NAND4_X1 U2564 ( .A1(n2654), .A2(n2653), .A3(n2652), .A4(n2651), .ZN(n3961)
         );
  NAND4_X1 U2565 ( .A1(n2634), .A2(n2633), .A3(n2632), .A4(n2631), .ZN(n4057)
         );
  INV_X1 U2566 ( .A(n2240), .ZN(n4478) );
  NAND2_X1 U2567 ( .A1(n2174), .A2(n2173), .ZN(n4479) );
  INV_X1 U2568 ( .A(n4471), .ZN(n4476) );
  OR2_X1 U2569 ( .A1(n4381), .A2(n3853), .ZN(n4485) );
  NAND2_X1 U2570 ( .A1(n4201), .A2(n2231), .ZN(n4207) );
  OR2_X1 U2571 ( .A1(n3947), .A2(n3946), .ZN(n2231) );
  NAND2_X1 U2572 ( .A1(n3382), .A2(n2206), .ZN(n2761) );
  INV_X1 U2573 ( .A(n2207), .ZN(n2206) );
  OAI21_X1 U2574 ( .B1(n3387), .B2(n4522), .A(n2723), .ZN(n2207) );
  INV_X1 U2575 ( .A(n4354), .ZN(n2774) );
  INV_X1 U2576 ( .A(n3919), .ZN(n4490) );
  NOR2_X1 U2577 ( .A1(n4435), .A2(n2246), .ZN(n3916) );
  AND2_X1 U2578 ( .A1(n4440), .A2(REG2_REG_15__SCAN_IN), .ZN(n2246) );
  OR2_X1 U2579 ( .A1(n4144), .A2(n4023), .ZN(n4105) );
  OR2_X1 U2580 ( .A1(n2570), .A2(n4599), .ZN(n2584) );
  AND2_X1 U2581 ( .A1(n3327), .A2(n3324), .ZN(n3791) );
  OR3_X1 U2582 ( .A1(n2531), .A2(n2530), .A3(n2529), .ZN(n2539) );
  INV_X1 U2583 ( .A(REG3_REG_12__SCAN_IN), .ZN(n2530) );
  NAND2_X1 U2584 ( .A1(n2507), .A2(REG3_REG_11__SCAN_IN), .ZN(n2531) );
  INV_X1 U2585 ( .A(n2320), .ZN(n2319) );
  OAI21_X1 U2586 ( .B1(n2471), .B2(n2321), .A(n2484), .ZN(n2320) );
  NAND2_X1 U2587 ( .A1(n2319), .A2(n2321), .ZN(n2318) );
  INV_X1 U2588 ( .A(REG3_REG_14__SCAN_IN), .ZN(n4805) );
  INV_X1 U2589 ( .A(REG3_REG_8__SCAN_IN), .ZN(n4597) );
  INV_X1 U2590 ( .A(IR_REG_22__SCAN_IN), .ZN(n4814) );
  AOI21_X1 U2591 ( .B1(n2197), .B2(n2140), .A(n2192), .ZN(n3935) );
  NAND2_X1 U2592 ( .A1(n2193), .A2(n2707), .ZN(n2192) );
  NAND2_X1 U2593 ( .A1(n2137), .A2(n2194), .ZN(n2193) );
  OR2_X1 U2594 ( .A1(n3977), .A2(n3957), .ZN(n2752) );
  OR2_X1 U2595 ( .A1(n2233), .A2(n2235), .ZN(n2232) );
  OR2_X1 U2596 ( .A1(n4050), .A2(n4039), .ZN(n2233) );
  NOR2_X1 U2597 ( .A1(n2223), .A2(n4181), .ZN(n2222) );
  NAND2_X1 U2598 ( .A1(n2222), .A2(n4151), .ZN(n2221) );
  AND2_X1 U2599 ( .A1(n3211), .A2(n3299), .ZN(n2226) );
  NAND2_X1 U2600 ( .A1(n3020), .A2(n2681), .ZN(n2230) );
  INV_X1 U2601 ( .A(n3073), .ZN(n2229) );
  INV_X1 U2602 ( .A(IR_REG_17__SCAN_IN), .ZN(n2590) );
  INV_X1 U2603 ( .A(n3649), .ZN(n2269) );
  NAND2_X1 U2604 ( .A1(n2288), .A2(n2289), .ZN(n2287) );
  INV_X1 U2605 ( .A(n3621), .ZN(n2288) );
  NAND2_X1 U2606 ( .A1(n3621), .A2(n3620), .ZN(n2285) );
  AND2_X1 U2607 ( .A1(n3630), .A2(n2255), .ZN(n2254) );
  NAND2_X1 U2608 ( .A1(n3261), .A2(n3260), .ZN(n3266) );
  NOR2_X1 U2609 ( .A1(n2584), .A2(n3643), .ZN(n2595) );
  NAND2_X1 U2610 ( .A1(n3602), .A2(n2145), .ZN(n2260) );
  INV_X1 U2611 ( .A(REG3_REG_24__SCAN_IN), .ZN(n4600) );
  NAND2_X1 U2612 ( .A1(n3008), .A2(n3007), .ZN(n2292) );
  INV_X1 U2613 ( .A(n3516), .ZN(n3435) );
  INV_X1 U2614 ( .A(REG3_REG_18__SCAN_IN), .ZN(n3643) );
  OR2_X1 U2615 ( .A1(n2716), .A2(n4012), .ZN(n2638) );
  OR2_X1 U2616 ( .A1(n2405), .A2(n2406), .ZN(n2407) );
  NAND2_X1 U2617 ( .A1(n3869), .A2(n2803), .ZN(n2815) );
  NOR2_X1 U2618 ( .A1(n2864), .A2(n2245), .ZN(n2819) );
  AND2_X1 U2619 ( .A1(n2829), .A2(REG2_REG_5__SCAN_IN), .ZN(n2245) );
  XNOR2_X1 U2620 ( .A(n2880), .B(n2840), .ZN(n2837) );
  OR2_X1 U2621 ( .A1(n3902), .A2(n2237), .ZN(n3906) );
  NOR2_X1 U2622 ( .A1(n3903), .A2(n3904), .ZN(n2237) );
  NAND2_X1 U2623 ( .A1(n2302), .A2(REG1_REG_12__SCAN_IN), .ZN(n2301) );
  NAND2_X1 U2624 ( .A1(n3891), .A2(n2302), .ZN(n2300) );
  INV_X1 U2625 ( .A(n4412), .ZN(n2302) );
  NOR2_X1 U2626 ( .A1(n4403), .A2(n4692), .ZN(n4402) );
  NAND2_X1 U2627 ( .A1(n4397), .A2(n3908), .ZN(n3910) );
  OR2_X1 U2628 ( .A1(n4423), .A2(n3914), .ZN(n2248) );
  XNOR2_X1 U2629 ( .A(n3916), .B(n2303), .ZN(n4448) );
  NAND2_X1 U2630 ( .A1(n4449), .A2(n3896), .ZN(n4461) );
  NAND2_X1 U2631 ( .A1(n3973), .A2(n2234), .ZN(n2649) );
  INV_X1 U2632 ( .A(n2305), .ZN(n3985) );
  OR2_X1 U2633 ( .A1(n2155), .A2(n2310), .ZN(n2308) );
  INV_X1 U2634 ( .A(n2307), .ZN(n2306) );
  NAND2_X1 U2635 ( .A1(n2188), .A2(n2187), .ZN(n2704) );
  NOR2_X1 U2636 ( .A1(n2158), .A2(n2141), .ZN(n2187) );
  NAND2_X1 U2637 ( .A1(n3679), .A2(DATAI_23_), .ZN(n4033) );
  NOR2_X1 U2638 ( .A1(n4596), .A2(n2613), .ZN(n2628) );
  AND2_X1 U2639 ( .A1(n3804), .A2(n4028), .ZN(n4067) );
  AND2_X1 U2640 ( .A1(n2595), .A2(REG3_REG_19__SCAN_IN), .ZN(n2606) );
  INV_X1 U2641 ( .A(n4095), .ZN(n3441) );
  NOR2_X1 U2642 ( .A1(n4133), .A2(n3522), .ZN(n4094) );
  OAI21_X1 U2643 ( .B1(n4188), .B2(n4160), .A(n2189), .ZN(n4144) );
  AOI21_X1 U2644 ( .B1(n4177), .B2(n2556), .A(n2555), .ZN(n4161) );
  INV_X1 U2645 ( .A(n3396), .ZN(n3624) );
  NOR2_X1 U2646 ( .A1(n3241), .A2(n2341), .ZN(n2515) );
  NOR2_X1 U2647 ( .A1(n3249), .A2(n3299), .ZN(n2341) );
  NAND2_X1 U2648 ( .A1(n2198), .A2(n2139), .ZN(n2686) );
  NOR2_X1 U2649 ( .A1(n2487), .A2(n4771), .ZN(n2500) );
  NAND2_X1 U2650 ( .A1(n3185), .A2(n3211), .ZN(n3223) );
  NAND2_X1 U2651 ( .A1(n2198), .A2(n2200), .ZN(n3180) );
  NOR2_X1 U2652 ( .A1(n2213), .A2(n2214), .ZN(n2212) );
  NAND2_X1 U2653 ( .A1(n2211), .A2(n2209), .ZN(n2208) );
  INV_X1 U2654 ( .A(n3765), .ZN(n2214) );
  NOR2_X1 U2655 ( .A1(n3073), .A2(n2230), .ZN(n3086) );
  OR2_X1 U2656 ( .A1(n2972), .A2(n3368), .ZN(n3073) );
  NOR2_X1 U2657 ( .A1(n3073), .A2(n3074), .ZN(n3072) );
  NAND2_X1 U2658 ( .A1(n3679), .A2(n2382), .ZN(n2383) );
  NAND2_X1 U2659 ( .A1(IR_REG_1__SCAN_IN), .A2(n2144), .ZN(n4824) );
  NOR2_X1 U2660 ( .A1(n4201), .A2(n4204), .ZN(n4200) );
  NOR2_X1 U2661 ( .A1(n2752), .A2(n3929), .ZN(n3947) );
  NAND2_X1 U2662 ( .A1(n3679), .A2(DATAI_27_), .ZN(n4210) );
  NAND2_X1 U2663 ( .A1(n3679), .A2(DATAI_26_), .ZN(n3978) );
  NAND2_X1 U2664 ( .A1(n3995), .A2(n3978), .ZN(n3977) );
  NOR2_X1 U2665 ( .A1(n4069), .A2(n2233), .ZN(n4040) );
  NOR2_X1 U2666 ( .A1(n4178), .A2(n2220), .ZN(n4168) );
  INV_X1 U2667 ( .A(n2222), .ZN(n2220) );
  OR2_X1 U2668 ( .A1(n3345), .A2(n3500), .ZN(n4178) );
  NOR2_X1 U2669 ( .A1(n3255), .A2(n4287), .ZN(n3336) );
  NAND2_X1 U2670 ( .A1(n3185), .A2(n2225), .ZN(n3255) );
  AND2_X1 U2671 ( .A1(n2226), .A2(n3287), .ZN(n2225) );
  NAND2_X1 U2672 ( .A1(n3185), .A2(n2226), .ZN(n3253) );
  NOR2_X1 U2673 ( .A1(n3128), .A2(n3127), .ZN(n3167) );
  AND2_X1 U2674 ( .A1(n3167), .A2(n3192), .ZN(n3185) );
  INV_X1 U2675 ( .A(n3171), .ZN(n3192) );
  NAND2_X1 U2676 ( .A1(n2228), .A2(n2229), .ZN(n3128) );
  NOR3_X1 U2677 ( .A1(n3080), .A2(n2230), .A3(n3092), .ZN(n2228) );
  NAND2_X1 U2678 ( .A1(n2229), .A2(n2227), .ZN(n3085) );
  NOR2_X1 U2679 ( .A1(n3080), .A2(n2230), .ZN(n2227) );
  INV_X1 U2680 ( .A(n4275), .ZN(n4288) );
  NAND2_X1 U2681 ( .A1(n2402), .A2(n2401), .ZN(n2952) );
  NAND2_X1 U2682 ( .A1(n3677), .A2(n2134), .ZN(n2401) );
  INV_X1 U2683 ( .A(n4508), .ZN(n4540) );
  AND2_X1 U2684 ( .A1(n2973), .A2(n2392), .ZN(n2951) );
  INV_X1 U2685 ( .A(n4289), .ZN(n4276) );
  NOR2_X1 U2686 ( .A1(n2966), .A2(n2748), .ZN(n2760) );
  INV_X1 U2687 ( .A(n4527), .ZN(n4522) );
  INV_X1 U2688 ( .A(n4162), .ZN(n4553) );
  INV_X1 U2689 ( .A(n4355), .ZN(n2749) );
  AND2_X1 U2690 ( .A1(n2891), .A2(n4488), .ZN(n2932) );
  NAND2_X1 U2691 ( .A1(n2733), .A2(n2732), .ZN(n2942) );
  XNOR2_X1 U2692 ( .A(n2290), .B(IR_REG_20__SCAN_IN), .ZN(n2676) );
  XNOR2_X1 U2693 ( .A(n2580), .B(IR_REG_17__SCAN_IN), .ZN(n3918) );
  INV_X1 U2694 ( .A(IR_REG_16__SCAN_IN), .ZN(n2576) );
  AND2_X1 U2695 ( .A1(n2340), .A2(n2326), .ZN(n2325) );
  NAND2_X1 U2696 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_6__SCAN_IN), .ZN(n4817)
         );
  AOI21_X1 U2697 ( .B1(n2147), .B2(n3110), .A(n2277), .ZN(n2276) );
  NOR2_X1 U2698 ( .A1(n3048), .A2(n2278), .ZN(n2277) );
  INV_X1 U2699 ( .A(n3961), .ZN(n3988) );
  XNOR2_X1 U2700 ( .A(n3526), .B(n3525), .ZN(n3528) );
  INV_X1 U2701 ( .A(n4274), .ZN(n3500) );
  INV_X1 U2702 ( .A(n4033), .ZN(n4039) );
  NOR2_X1 U2703 ( .A1(n3613), .A2(n3557), .ZN(n3560) );
  NAND2_X1 U2704 ( .A1(n3679), .A2(DATAI_21_), .ZN(n4238) );
  INV_X1 U2705 ( .A(n3836), .ZN(n4111) );
  OR2_X1 U2706 ( .A1(n2657), .A2(n2643), .ZN(n3996) );
  NAND2_X1 U2707 ( .A1(n3581), .A2(n3580), .ZN(n3579) );
  INV_X1 U2708 ( .A(n4057), .ZN(n4008) );
  INV_X1 U2709 ( .A(n4563), .ZN(n3375) );
  INV_X1 U2710 ( .A(n2257), .ZN(n3613) );
  NAND2_X1 U2711 ( .A1(n2293), .A2(n2163), .ZN(n3392) );
  NAND2_X1 U2712 ( .A1(n2257), .A2(n2258), .ZN(n2256) );
  AND2_X1 U2713 ( .A1(n2930), .A2(n2929), .ZN(n3635) );
  INV_X1 U2714 ( .A(n4134), .ZN(n4124) );
  NAND2_X1 U2715 ( .A1(n3579), .A2(n3048), .ZN(n3112) );
  NAND2_X1 U2716 ( .A1(n2938), .A2(n3853), .ZN(n3655) );
  NAND2_X1 U2717 ( .A1(n2270), .A2(n2164), .ZN(n2265) );
  INV_X1 U2718 ( .A(n3654), .ZN(n3666) );
  INV_X1 U2719 ( .A(n3653), .ZN(n3671) );
  OR2_X1 U2720 ( .A1(n2420), .A2(n2393), .ZN(n2397) );
  OR2_X1 U2721 ( .A1(n2405), .A2(n4543), .ZN(n2372) );
  OR2_X1 U2722 ( .A1(n2420), .A2(n4666), .ZN(n2388) );
  OR2_X1 U2723 ( .A1(n2423), .A2(n2386), .ZN(n2390) );
  INV_X1 U2724 ( .A(n2236), .ZN(n3867) );
  XNOR2_X1 U2725 ( .A(n2815), .B(n2813), .ZN(n2814) );
  INV_X1 U2726 ( .A(n2818), .ZN(n3882) );
  XNOR2_X1 U2727 ( .A(n2819), .B(n4362), .ZN(n2845) );
  NAND2_X1 U2728 ( .A1(n2244), .A2(n2243), .ZN(n2860) );
  INV_X1 U2729 ( .A(n2856), .ZN(n2243) );
  INV_X1 U2730 ( .A(n2244), .ZN(n2857) );
  NAND2_X1 U2731 ( .A1(n2833), .A2(n2832), .ZN(n2855) );
  XNOR2_X1 U2732 ( .A(n3906), .B(n2299), .ZN(n4389) );
  NAND2_X1 U2733 ( .A1(n4389), .A2(REG2_REG_10__SCAN_IN), .ZN(n4388) );
  INV_X1 U2734 ( .A(n2298), .ZN(n4383) );
  NAND2_X1 U2735 ( .A1(n4398), .A2(n4399), .ZN(n4397) );
  XNOR2_X1 U2736 ( .A(n3910), .B(n4500), .ZN(n4408) );
  NAND2_X1 U2737 ( .A1(n4408), .A2(REG2_REG_12__SCAN_IN), .ZN(n4407) );
  XNOR2_X1 U2738 ( .A(n2177), .B(n4427), .ZN(n4424) );
  INV_X1 U2739 ( .A(n3913), .ZN(n2177) );
  NOR2_X1 U2740 ( .A1(n4424), .A2(n3347), .ZN(n4423) );
  XNOR2_X1 U2741 ( .A(n2566), .B(IR_REG_15__SCAN_IN), .ZN(n4440) );
  AND2_X1 U2742 ( .A1(n2248), .A2(n2247), .ZN(n4435) );
  INV_X1 U2743 ( .A(n4436), .ZN(n2247) );
  INV_X1 U2744 ( .A(n2248), .ZN(n4437) );
  NAND2_X1 U2745 ( .A1(n4447), .A2(n3917), .ZN(n4458) );
  NAND2_X1 U2746 ( .A1(n4458), .A2(n4459), .ZN(n4457) );
  AND2_X1 U2747 ( .A1(n2240), .A2(n2239), .ZN(n3922) );
  NAND2_X1 U2748 ( .A1(n3919), .A2(REG2_REG_18__SCAN_IN), .ZN(n2239) );
  NAND2_X1 U2749 ( .A1(n3968), .A2(n3816), .ZN(n2195) );
  OAI21_X1 U2750 ( .B1(n4049), .B2(n2310), .A(n2309), .ZN(n4002) );
  NAND2_X1 U2751 ( .A1(n4048), .A2(n2627), .ZN(n4021) );
  NAND2_X1 U2752 ( .A1(n2327), .A2(n2582), .ZN(n4129) );
  NAND2_X1 U2753 ( .A1(n4165), .A2(n4164), .ZN(n4163) );
  NAND2_X1 U2754 ( .A1(n4188), .A2(n3689), .ZN(n4165) );
  NAND2_X1 U2755 ( .A1(n3133), .A2(n2473), .ZN(n3176) );
  INV_X1 U2756 ( .A(n4193), .ZN(n4139) );
  NAND2_X1 U2757 ( .A1(n2419), .A2(n2418), .ZN(n2989) );
  INV_X1 U2758 ( .A(n4568), .ZN(n4169) );
  AND2_X1 U2759 ( .A1(n4372), .A2(n4288), .ZN(n4552) );
  INV_X1 U2760 ( .A(n2952), .ZN(n3368) );
  AND2_X1 U2761 ( .A1(n4171), .A2(n2982), .ZN(n4100) );
  OAI211_X1 U2762 ( .C1(n4534), .C2(n4207), .A(n4208), .B(n4209), .ZN(n4307)
         );
  OR2_X1 U2763 ( .A1(n3995), .A2(n3994), .ZN(n4316) );
  NAND2_X1 U2764 ( .A1(n2771), .A2(n2932), .ZN(n4486) );
  INV_X1 U2765 ( .A(n2185), .ZN(n2363) );
  INV_X1 U2766 ( .A(n2366), .ZN(n4352) );
  MUX2_X1 U2767 ( .A(n2712), .B(n2711), .S(IR_REG_28__SCAN_IN), .Z(n4368) );
  XNOR2_X1 U2768 ( .A(n2724), .B(IR_REG_26__SCAN_IN), .ZN(n4353) );
  NAND2_X1 U2769 ( .A1(n2138), .A2(IR_REG_31__SCAN_IN), .ZN(n2724) );
  INV_X1 U2770 ( .A(n2513), .ZN(n2184) );
  XNOR2_X1 U2771 ( .A(n2729), .B(n2728), .ZN(n4354) );
  XNOR2_X1 U2772 ( .A(n2726), .B(IR_REG_24__SCAN_IN), .ZN(n4355) );
  NAND2_X1 U2773 ( .A1(n2733), .A2(IR_REG_31__SCAN_IN), .ZN(n2726) );
  AND2_X1 U2774 ( .A1(n2942), .A2(STATE_REG_SCAN_IN), .ZN(n4488) );
  XNOR2_X1 U2775 ( .A(n2674), .B(IR_REG_22__SCAN_IN), .ZN(n4356) );
  INV_X1 U2776 ( .A(n2676), .ZN(n4357) );
  INV_X1 U2777 ( .A(n3901), .ZN(n4501) );
  AND2_X1 U2778 ( .A1(n2432), .A2(n2416), .ZN(n4364) );
  AOI21_X1 U2779 ( .B1(n4477), .B2(n4476), .A(n4475), .ZN(n4484) );
  OR2_X1 U2780 ( .A1(n4542), .A2(REG0_REG_28__SCAN_IN), .ZN(n2205) );
  OR2_X1 U2781 ( .A1(n2354), .A2(n2353), .ZN(n2136) );
  INV_X1 U2782 ( .A(n3764), .ZN(n2213) );
  AND2_X1 U2783 ( .A1(n3960), .A2(n3743), .ZN(n2137) );
  NAND3_X1 U2784 ( .A1(n2184), .A2(n2334), .A3(n2143), .ZN(n2138) );
  AND2_X1 U2785 ( .A1(n2200), .A2(n2168), .ZN(n2139) );
  AND2_X1 U2786 ( .A1(n2137), .A2(n2196), .ZN(n2140) );
  AND2_X1 U2787 ( .A1(n2256), .A2(n2255), .ZN(n3629) );
  NAND2_X1 U2788 ( .A1(n2384), .A2(n2383), .ZN(n2978) );
  NAND2_X1 U2789 ( .A1(n4026), .A2(n3808), .ZN(n2141) );
  NAND2_X1 U2790 ( .A1(n4034), .A2(n4224), .ZN(n2142) );
  INV_X1 U2791 ( .A(n4260), .ZN(n2223) );
  AND2_X1 U2792 ( .A1(n3553), .A2(n2259), .ZN(n2258) );
  NAND2_X1 U2793 ( .A1(n2292), .A2(n3012), .ZN(n3013) );
  AND3_X1 U2794 ( .A1(n4821), .A2(IR_REG_18__SCAN_IN), .A3(IR_REG_12__SCAN_IN), 
        .ZN(n2144) );
  NAND4_X1 U2795 ( .A1(n2391), .A2(n2390), .A3(n2389), .A4(n2388), .ZN(n2897)
         );
  XNOR2_X1 U2796 ( .A(n2360), .B(IR_REG_29__SCAN_IN), .ZN(n2366) );
  NAND2_X1 U2797 ( .A1(n2265), .A2(n3566), .ZN(n3648) );
  NAND2_X1 U2798 ( .A1(n2264), .A2(n2266), .ZN(n3529) );
  AND2_X1 U2799 ( .A1(n2346), .A2(n2325), .ZN(n2455) );
  NAND2_X2 U2800 ( .A1(n2892), .A2(n2891), .ZN(n3445) );
  INV_X1 U2801 ( .A(IR_REG_2__SCAN_IN), .ZN(n2400) );
  AND2_X1 U2802 ( .A1(n2262), .A2(n3605), .ZN(n2145) );
  NAND2_X1 U2803 ( .A1(n2346), .A2(n2340), .ZN(n2442) );
  AND3_X1 U2804 ( .A1(n2409), .A2(n2408), .A3(n2407), .ZN(n2146) );
  OR2_X1 U2805 ( .A1(n2280), .A2(n3111), .ZN(n2147) );
  OR3_X1 U2806 ( .A1(n2513), .A2(n2136), .A3(n2350), .ZN(n2148) );
  INV_X1 U2807 ( .A(IR_REG_10__SCAN_IN), .ZN(n2348) );
  NAND2_X1 U2808 ( .A1(n2266), .A2(n2263), .ZN(n2149) );
  NAND2_X1 U2809 ( .A1(n2604), .A2(IR_REG_31__SCAN_IN), .ZN(n2673) );
  OR2_X1 U2810 ( .A1(n3889), .A2(n2299), .ZN(n2150) );
  AND2_X1 U2811 ( .A1(n2195), .A2(n3743), .ZN(n2151) );
  AND2_X1 U2812 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2152)
         );
  AND2_X1 U2813 ( .A1(n2318), .A2(n2485), .ZN(n2153) );
  AND2_X1 U2814 ( .A1(n2326), .A2(n2324), .ZN(n2154) );
  INV_X1 U2815 ( .A(IR_REG_31__SCAN_IN), .ZN(n2357) );
  INV_X1 U2816 ( .A(n3905), .ZN(n2299) );
  NAND2_X1 U2817 ( .A1(n2545), .A2(n2351), .ZN(n2579) );
  AND2_X1 U2818 ( .A1(n3990), .A2(n2235), .ZN(n2155) );
  NAND2_X1 U2819 ( .A1(n2293), .A2(n2294), .ZN(n3388) );
  OR2_X1 U2820 ( .A1(n4069), .A2(n4050), .ZN(n2156) );
  AND2_X1 U2821 ( .A1(n3566), .A2(n2269), .ZN(n2268) );
  INV_X1 U2822 ( .A(IR_REG_20__SCAN_IN), .ZN(n2671) );
  AND2_X1 U2823 ( .A1(n3484), .A2(n3483), .ZN(n2157) );
  INV_X1 U2824 ( .A(n3620), .ZN(n2289) );
  INV_X1 U2825 ( .A(n3270), .ZN(n3299) );
  AND2_X1 U2826 ( .A1(n2189), .A2(n4160), .ZN(n2158) );
  NOR2_X1 U2827 ( .A1(n4402), .A2(n3891), .ZN(n2159) );
  AND2_X1 U2828 ( .A1(n4359), .A2(REG1_REG_9__SCAN_IN), .ZN(n2160) );
  AND2_X1 U2829 ( .A1(n3720), .A2(n2582), .ZN(n2161) );
  NOR2_X1 U2830 ( .A1(n3972), .A2(n3957), .ZN(n2162) );
  INV_X1 U2831 ( .A(n2627), .ZN(n2313) );
  NAND2_X1 U2832 ( .A1(n4036), .A2(n4050), .ZN(n2627) );
  AND2_X1 U2833 ( .A1(n3390), .A2(n2294), .ZN(n2163) );
  NAND2_X1 U2834 ( .A1(n3478), .A2(n3477), .ZN(n2164) );
  NAND3_X1 U2835 ( .A1(n2323), .A2(n2346), .A3(n2347), .ZN(n2165) );
  INV_X1 U2836 ( .A(n3728), .ZN(n2196) );
  AND2_X1 U2837 ( .A1(n2286), .A2(n2285), .ZN(n2166) );
  INV_X1 U2838 ( .A(n3287), .ZN(n3252) );
  INV_X1 U2839 ( .A(n2635), .ZN(n2314) );
  INV_X1 U2840 ( .A(n2655), .ZN(n2333) );
  NAND2_X1 U2841 ( .A1(n2268), .A2(n3527), .ZN(n2167) );
  INV_X1 U2842 ( .A(n3557), .ZN(n2259) );
  NAND2_X1 U2843 ( .A1(n2472), .A2(n2471), .ZN(n3133) );
  NAND2_X1 U2844 ( .A1(n3297), .A2(n3211), .ZN(n2168) );
  INV_X1 U2845 ( .A(n3611), .ZN(n2253) );
  INV_X1 U2846 ( .A(n3799), .ZN(n2190) );
  OAI21_X1 U2847 ( .B1(n3203), .B2(n3202), .A(n3204), .ZN(n3261) );
  NAND2_X1 U2848 ( .A1(n3147), .A2(n3146), .ZN(n3203) );
  NAND2_X1 U2849 ( .A1(n2273), .A2(n2276), .ZN(n3142) );
  NAND2_X1 U2850 ( .A1(n3679), .A2(DATAI_24_), .ZN(n4224) );
  INV_X1 U2851 ( .A(n4224), .ZN(n2235) );
  OR2_X1 U2852 ( .A1(n4178), .A2(n4181), .ZN(n2169) );
  AND2_X1 U2853 ( .A1(n3406), .A2(n3405), .ZN(n2170) );
  NOR3_X1 U2854 ( .A1(n4178), .A2(n2221), .A3(n4124), .ZN(n2224) );
  NAND2_X1 U2855 ( .A1(n2292), .A2(n2291), .ZN(n3041) );
  INV_X1 U2856 ( .A(n2219), .ZN(n4150) );
  NOR2_X1 U2857 ( .A1(n4178), .A2(n2221), .ZN(n2219) );
  INV_X1 U2858 ( .A(IR_REG_15__SCAN_IN), .ZN(n2577) );
  XNOR2_X1 U2859 ( .A(n2568), .B(n2576), .ZN(n4494) );
  INV_X1 U2860 ( .A(n4494), .ZN(n2303) );
  NAND4_X2 U2861 ( .A1(n2372), .A2(n2371), .A3(n2369), .A4(n2370), .ZN(n3842)
         );
  INV_X1 U2862 ( .A(n3993), .ZN(n2234) );
  NAND2_X1 U2863 ( .A1(n2950), .A2(n2403), .ZN(n3063) );
  INV_X1 U2864 ( .A(n4459), .ZN(n2176) );
  INV_X1 U2865 ( .A(IR_REG_0__SCAN_IN), .ZN(n2217) );
  INV_X1 U2866 ( .A(DATAI_0_), .ZN(n2218) );
  INV_X1 U2867 ( .A(n4555), .ZN(n4358) );
  NAND2_X1 U2868 ( .A1(n4555), .A2(n4356), .ZN(n2936) );
  NOR2_X1 U2869 ( .A1(n2399), .A2(n2357), .ZN(n2180) );
  AOI22_X1 U2870 ( .A1(n3533), .A2(n3842), .B1(n2911), .B2(n3549), .ZN(n2913)
         );
  NAND3_X1 U2871 ( .A1(n2186), .A2(n2323), .A3(n2346), .ZN(n2513) );
  NAND3_X1 U2872 ( .A1(n2183), .A2(n2334), .A3(n2143), .ZN(n2185) );
  NAND2_X1 U2873 ( .A1(n4188), .A2(n2189), .ZN(n2188) );
  INV_X1 U2874 ( .A(n3123), .ZN(n2199) );
  OAI21_X1 U2875 ( .B1(n3123), .B2(n2685), .A(n3776), .ZN(n3164) );
  AOI21_X1 U2876 ( .B1(n2685), .B2(n3776), .A(n2204), .ZN(n2203) );
  AOI21_X1 U2877 ( .B1(n2993), .B2(n2212), .A(n2208), .ZN(n3025) );
  INV_X1 U2878 ( .A(n3774), .ZN(n2215) );
  OAI21_X1 U2879 ( .B1(n2993), .B2(n2682), .A(n3765), .ZN(n3079) );
  NAND4_X1 U2880 ( .A1(n2721), .A2(n2671), .A3(n2577), .A4(n2216), .ZN(n2353)
         );
  AOI21_X1 U2881 ( .B1(n2673), .B2(n2216), .A(n2357), .ZN(n2290) );
  XNOR2_X1 U2882 ( .A(n2673), .B(n2216), .ZN(n4555) );
  MUX2_X1 U2883 ( .A(n2218), .B(n2217), .S(n3677), .Z(n4563) );
  INV_X1 U2884 ( .A(n2224), .ZN(n4133) );
  NOR3_X4 U2885 ( .A1(IR_REG_6__SCAN_IN), .A2(IR_REG_8__SCAN_IN), .A3(
        IR_REG_7__SCAN_IN), .ZN(n2347) );
  NAND2_X1 U2886 ( .A1(n4607), .A2(IR_REG_31__SCAN_IN), .ZN(n2238) );
  OAI21_X1 U2887 ( .B1(n2152), .B2(n4607), .A(n2238), .ZN(n2381) );
  INV_X1 U2888 ( .A(n3556), .ZN(n2252) );
  NAND2_X1 U2889 ( .A1(n2249), .A2(n2250), .ZN(n3504) );
  NAND2_X1 U2890 ( .A1(n3556), .A2(n2258), .ZN(n2249) );
  NAND2_X1 U2891 ( .A1(n3602), .A2(n3605), .ZN(n2271) );
  INV_X1 U2892 ( .A(n3604), .ZN(n2272) );
  NAND2_X1 U2893 ( .A1(n2261), .A2(n2260), .ZN(n3537) );
  OAI21_X1 U2894 ( .B1(n3604), .B2(n2167), .A(n2262), .ZN(n2261) );
  NAND3_X1 U2895 ( .A1(n2271), .A2(n2272), .A3(n2268), .ZN(n2264) );
  INV_X1 U2896 ( .A(n2270), .ZN(n3565) );
  NAND2_X1 U2897 ( .A1(n3581), .A2(n2274), .ZN(n2273) );
  NAND2_X1 U2898 ( .A1(n3619), .A2(n2282), .ZN(n2281) );
  NAND2_X1 U2899 ( .A1(n2281), .A2(n2283), .ZN(n3414) );
  NAND2_X1 U2900 ( .A1(n3305), .A2(n2295), .ZN(n2293) );
  OAI21_X1 U2901 ( .B1(n4049), .B2(n2308), .A(n2306), .ZN(n2305) );
  NAND2_X1 U2902 ( .A1(n2316), .A2(n2315), .ZN(n2758) );
  NAND2_X1 U2903 ( .A1(n2472), .A2(n2319), .ZN(n2317) );
  NAND2_X1 U2904 ( .A1(n2317), .A2(n2153), .ZN(n3189) );
  NAND2_X1 U2905 ( .A1(n2322), .A2(n2973), .ZN(n2950) );
  NAND2_X1 U2906 ( .A1(n2677), .A2(n2974), .ZN(n2973) );
  NAND3_X1 U2907 ( .A1(n2325), .A2(n2346), .A3(n2347), .ZN(n2493) );
  NAND2_X1 U2908 ( .A1(n2991), .A2(n2435), .ZN(n3084) );
  NAND2_X1 U2909 ( .A1(n2419), .A2(n2328), .ZN(n2991) );
  NAND2_X1 U2910 ( .A1(n2650), .A2(n2649), .ZN(n3966) );
  OR3_X1 U2911 ( .A1(n2513), .A2(n2335), .A3(n2136), .ZN(n2725) );
  NAND2_X1 U2912 ( .A1(n4094), .A2(n3441), .ZN(n4245) );
  AOI21_X1 U2913 ( .B1(n3375), .B2(n2911), .A(n2903), .ZN(n2904) );
  AND2_X1 U2914 ( .A1(n2897), .A2(n3375), .ZN(n2974) );
  OR2_X1 U2915 ( .A1(n2891), .A2(n2900), .ZN(n2337) );
  OR2_X1 U2916 ( .A1(n2891), .A2(n2764), .ZN(n3856) );
  OR2_X1 U2917 ( .A1(n3652), .A2(n4210), .ZN(n2338) );
  OR2_X1 U2918 ( .A1(n4057), .A2(n4039), .ZN(n2339) );
  AND2_X1 U2919 ( .A1(n2414), .A2(n2433), .ZN(n2340) );
  AND2_X1 U2920 ( .A1(n3961), .A2(n3658), .ZN(n2342) );
  OR3_X1 U2921 ( .A1(n3517), .A2(n3638), .A3(n3639), .ZN(n2343) );
  NAND2_X1 U2922 ( .A1(n3679), .A2(DATAI_22_), .ZN(n4060) );
  XNOR2_X1 U2923 ( .A(n2895), .B(n3530), .ZN(n3009) );
  NAND2_X1 U2924 ( .A1(n2971), .A2(n4169), .ZN(n4372) );
  INV_X1 U2925 ( .A(n4142), .ZN(n4171) );
  AND2_X1 U2926 ( .A1(n4290), .A2(n3396), .ZN(n2344) );
  OR2_X1 U2927 ( .A1(n4290), .A2(n3396), .ZN(n2345) );
  NAND2_X1 U2928 ( .A1(n3679), .A2(DATAI_25_), .ZN(n3993) );
  INV_X1 U2929 ( .A(n3973), .ZN(n4225) );
  INV_X1 U2930 ( .A(n4036), .ZN(n4239) );
  INV_X1 U2931 ( .A(n3720), .ZN(n4132) );
  INV_X1 U2932 ( .A(IR_REG_13__SCAN_IN), .ZN(n2351) );
  INV_X1 U2933 ( .A(IR_REG_28__SCAN_IN), .ZN(n2373) );
  INV_X1 U2934 ( .A(n3295), .ZN(n3271) );
  OR2_X1 U2935 ( .A1(n2374), .A2(n2373), .ZN(n2375) );
  INV_X1 U2936 ( .A(IR_REG_24__SCAN_IN), .ZN(n4815) );
  INV_X1 U2937 ( .A(n2891), .ZN(n2902) );
  INV_X1 U2938 ( .A(REG3_REG_13__SCAN_IN), .ZN(n2529) );
  NOR2_X1 U2939 ( .A1(n4008), .A2(n4033), .ZN(n2635) );
  AND2_X1 U2940 ( .A1(n3505), .A2(n3506), .ZN(n3465) );
  OR2_X1 U2941 ( .A1(n3526), .A2(n3525), .ZN(n3527) );
  INV_X1 U2942 ( .A(REG3_REG_21__SCAN_IN), .ZN(n4596) );
  INV_X1 U2943 ( .A(n3016), .ZN(n3014) );
  NAND2_X1 U2944 ( .A1(n2343), .A2(n3435), .ZN(n3436) );
  NOR2_X1 U2945 ( .A1(n2539), .A2(n4805), .ZN(n2560) );
  NOR2_X1 U2946 ( .A1(n2636), .A2(n4600), .ZN(n2642) );
  OR2_X1 U2947 ( .A1(n2476), .A2(n4597), .ZN(n2487) );
  AND2_X1 U2948 ( .A1(n2657), .A2(n2656), .ZN(n2665) );
  NAND2_X1 U2949 ( .A1(n2606), .A2(REG3_REG_20__SCAN_IN), .ZN(n2613) );
  AND2_X1 U2950 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .ZN(
        n2437) );
  AND2_X1 U2951 ( .A1(n2932), .A2(n2931), .ZN(n2933) );
  INV_X1 U2952 ( .A(n4238), .ZN(n4074) );
  INV_X1 U2953 ( .A(n3768), .ZN(n2471) );
  AND2_X1 U2954 ( .A1(n2466), .A2(n4817), .ZN(n2468) );
  AND2_X1 U2955 ( .A1(n2500), .A2(REG3_REG_10__SCAN_IN), .ZN(n2507) );
  INV_X1 U2956 ( .A(n3990), .ZN(n4034) );
  INV_X1 U2957 ( .A(n3080), .ZN(n3585) );
  NOR2_X1 U2958 ( .A1(n2941), .A2(n3831), .ZN(n2938) );
  INV_X1 U2959 ( .A(REG3_REG_6__SCAN_IN), .ZN(n4768) );
  OR2_X1 U2960 ( .A1(n2665), .A2(n2658), .ZN(n3955) );
  OR2_X1 U2961 ( .A1(n2716), .A2(n3979), .ZN(n2651) );
  INV_X1 U2962 ( .A(REG3_REG_9__SCAN_IN), .ZN(n4771) );
  NOR2_X1 U2963 ( .A1(n3894), .A2(n4421), .ZN(n4433) );
  INV_X1 U2964 ( .A(REG3_REG_17__SCAN_IN), .ZN(n4599) );
  OR2_X1 U2965 ( .A1(n3745), .A2(n3744), .ZN(n3937) );
  AND2_X1 U2966 ( .A1(n3988), .A2(n3978), .ZN(n2655) );
  INV_X1 U2967 ( .A(n4060), .ZN(n4050) );
  INV_X1 U2968 ( .A(n3208), .ZN(n3211) );
  INV_X1 U2969 ( .A(n3723), .ZN(n2992) );
  AND2_X1 U2970 ( .A1(n4540), .A2(n2933), .ZN(n4568) );
  OR2_X1 U2971 ( .A1(n2771), .A2(D_REG_0__SCAN_IN), .ZN(n2750) );
  INV_X1 U2972 ( .A(n4357), .ZN(n2756) );
  XNOR2_X1 U2973 ( .A(n3143), .B(n3144), .ZN(n3141) );
  INV_X1 U2974 ( .A(n4210), .ZN(n3957) );
  INV_X1 U2975 ( .A(n2754), .ZN(n3929) );
  NAND2_X1 U2976 ( .A1(n2945), .A2(STATE_REG_SCAN_IN), .ZN(n3654) );
  AND2_X1 U2977 ( .A1(n3679), .A2(DATAI_20_), .ZN(n4095) );
  NAND2_X1 U2978 ( .A1(n3293), .A2(n3275), .ZN(n3305) );
  INV_X1 U2979 ( .A(n3655), .ZN(n3667) );
  OR2_X1 U2980 ( .A1(n2716), .A2(n3955), .ZN(n2659) );
  OR2_X1 U2981 ( .A1(n2716), .A2(n3996), .ZN(n2645) );
  INV_X1 U2982 ( .A(n4468), .ZN(n4464) );
  AOI21_X1 U2983 ( .B1(n4470), .B2(n4469), .A(n4468), .ZN(n4477) );
  NOR2_X2 U2984 ( .A1(n4368), .A2(n2713), .ZN(n4187) );
  INV_X1 U2985 ( .A(n4152), .ZN(n4373) );
  AND2_X1 U2986 ( .A1(n2750), .A2(n2775), .ZN(n2968) );
  OR3_X1 U2987 ( .A1(n4357), .A2(n4356), .A3(n4555), .ZN(n4508) );
  INV_X1 U2988 ( .A(n3598), .ZN(n4151) );
  INV_X1 U2989 ( .A(n4534), .ZN(n4529) );
  INV_X1 U2990 ( .A(n2968), .ZN(n2759) );
  AND2_X1 U2991 ( .A1(n2778), .A2(n2798), .ZN(n4473) );
  INV_X1 U2992 ( .A(n3635), .ZN(n3674) );
  NAND4_X1 U2993 ( .A1(n2662), .A2(n2661), .A3(n2660), .A4(n2659), .ZN(n3972)
         );
  NAND4_X1 U2994 ( .A1(n2647), .A2(n2646), .A3(n2645), .A4(n2644), .ZN(n3973)
         );
  INV_X1 U2995 ( .A(n4482), .ZN(n4434) );
  OR2_X1 U2996 ( .A1(n4381), .A2(n4378), .ZN(n4468) );
  NAND2_X1 U2997 ( .A1(n4171), .A2(n3029), .ZN(n4193) );
  OR2_X1 U3000 ( .A1(n4137), .A2(n4534), .ZN(n4152) );
  NAND2_X1 U3001 ( .A1(n4551), .A2(n4529), .ZN(n4302) );
  AND2_X2 U3002 ( .A1(n2760), .A2(n2968), .ZN(n4551) );
  OR2_X1 U3003 ( .A1(n3378), .A2(n4350), .ZN(n2762) );
  NAND2_X1 U3004 ( .A1(n4542), .A2(n4529), .ZN(n4350) );
  AND2_X2 U3005 ( .A1(n2760), .A2(n2759), .ZN(n4542) );
  INV_X1 U3006 ( .A(n4542), .ZN(n4541) );
  INV_X1 U3007 ( .A(n4486), .ZN(n4487) );
  INV_X1 U3008 ( .A(n4427), .ZN(n4497) );
  AND2_X1 U3009 ( .A1(n2457), .A2(n2456), .ZN(n4362) );
  NOR2_X1 U3010 ( .A1(IR_REG_17__SCAN_IN), .A2(IR_REG_16__SCAN_IN), .ZN(n2352)
         );
  NAND4_X1 U3011 ( .A1(n2352), .A2(n2602), .A3(n2351), .A4(n4608), .ZN(n2354)
         );
  NAND3_X1 U3012 ( .A1(n4815), .A2(n2730), .A3(n2728), .ZN(n2355) );
  INV_X1 U3013 ( .A(IR_REG_26__SCAN_IN), .ZN(n2356) );
  NAND2_X1 U3014 ( .A1(n2374), .A2(n2359), .ZN(n2360) );
  NOR2_X1 U3015 ( .A1(IR_REG_29__SCAN_IN), .A2(IR_REG_28__SCAN_IN), .ZN(n2361)
         );
  AND2_X1 U3016 ( .A1(n2361), .A2(n2377), .ZN(n2362) );
  NAND2_X1 U3017 ( .A1(n2363), .A2(n2362), .ZN(n2769) );
  INV_X1 U3018 ( .A(n2367), .ZN(n2387) );
  INV_X1 U3019 ( .A(n2423), .ZN(n2365) );
  INV_X1 U3020 ( .A(REG3_REG_1__SCAN_IN), .ZN(n2983) );
  NAND2_X1 U3021 ( .A1(n2365), .A2(REG3_REG_1__SCAN_IN), .ZN(n2371) );
  AND2_X2 U3022 ( .A1(n2366), .A2(n2367), .ZN(n2410) );
  NAND2_X1 U3023 ( .A1(n2410), .A2(REG2_REG_1__SCAN_IN), .ZN(n2370) );
  INV_X1 U3024 ( .A(REG0_REG_1__SCAN_IN), .ZN(n4826) );
  NOR2_X1 U3025 ( .A1(n4826), .A2(n4352), .ZN(n2368) );
  NAND2_X1 U3026 ( .A1(n2368), .A2(n2387), .ZN(n2369) );
  NAND2_X1 U3027 ( .A1(n2374), .A2(n2377), .ZN(n2376) );
  NAND2_X1 U3028 ( .A1(n2376), .A2(n2375), .ZN(n2379) );
  NAND2_X1 U3029 ( .A1(n2377), .A2(IR_REG_28__SCAN_IN), .ZN(n2378) );
  INV_X1 U3030 ( .A(IR_REG_1__SCAN_IN), .ZN(n4607) );
  INV_X1 U3031 ( .A(n2399), .ZN(n2380) );
  NAND2_X1 U3032 ( .A1(n2381), .A2(n2380), .ZN(n2804) );
  NAND2_X1 U3033 ( .A1(n3677), .A2(n2804), .ZN(n2384) );
  INV_X1 U3034 ( .A(DATAI_1_), .ZN(n2382) );
  INV_X1 U3035 ( .A(n2978), .ZN(n3549) );
  NAND2_X1 U3036 ( .A1(n2385), .A2(n3549), .ZN(n2678) );
  NAND2_X1 U3037 ( .A1(n3842), .A2(n2978), .ZN(n3754) );
  NAND2_X1 U3038 ( .A1(n2678), .A2(n3754), .ZN(n2677) );
  INV_X1 U3039 ( .A(REG1_REG_0__SCAN_IN), .ZN(n2900) );
  OR2_X1 U3040 ( .A1(n2405), .A2(n2900), .ZN(n2391) );
  INV_X1 U3041 ( .A(REG3_REG_0__SCAN_IN), .ZN(n2386) );
  NAND2_X1 U3042 ( .A1(n2410), .A2(REG2_REG_0__SCAN_IN), .ZN(n2389) );
  NAND2_X1 U3043 ( .A1(n3842), .A2(n3549), .ZN(n2392) );
  INV_X1 U3044 ( .A(REG1_REG_2__SCAN_IN), .ZN(n2805) );
  OR2_X1 U3045 ( .A1(n2405), .A2(n2805), .ZN(n2398) );
  INV_X1 U3046 ( .A(REG0_REG_2__SCAN_IN), .ZN(n2393) );
  NAND2_X1 U3047 ( .A1(n2410), .A2(REG2_REG_2__SCAN_IN), .ZN(n2396) );
  INV_X1 U3048 ( .A(REG3_REG_2__SCAN_IN), .ZN(n2394) );
  OR2_X1 U3049 ( .A1(n2423), .A2(n2394), .ZN(n2395) );
  NAND4_X4 U3050 ( .A1(n2398), .A2(n2397), .A3(n2396), .A4(n2395), .ZN(n3841)
         );
  INV_X1 U3051 ( .A(DATAI_2_), .ZN(n4827) );
  OR2_X1 U3052 ( .A1(n3677), .A2(DATAI_2_), .ZN(n2402) );
  NAND2_X1 U3053 ( .A1(n3841), .A2(n2952), .ZN(n3759) );
  OR2_X1 U3054 ( .A1(n3841), .A2(n3368), .ZN(n2403) );
  OR2_X1 U3055 ( .A1(n2423), .A2(REG3_REG_3__SCAN_IN), .ZN(n2409) );
  INV_X1 U3056 ( .A(REG0_REG_3__SCAN_IN), .ZN(n2404) );
  OR2_X1 U3057 ( .A1(n2420), .A2(n2404), .ZN(n2408) );
  INV_X1 U3058 ( .A(REG1_REG_3__SCAN_IN), .ZN(n2406) );
  NAND2_X1 U3059 ( .A1(n2411), .A2(REG2_REG_3__SCAN_IN), .ZN(n2412) );
  NAND2_X1 U3060 ( .A1(n2413), .A2(IR_REG_31__SCAN_IN), .ZN(n2415) );
  NAND2_X1 U3061 ( .A1(n2415), .A2(n2414), .ZN(n2432) );
  OR2_X1 U3062 ( .A1(n2415), .A2(n2414), .ZN(n2416) );
  MUX2_X1 U3063 ( .A(n4364), .B(DATAI_3_), .S(n3679), .Z(n3074) );
  NAND2_X1 U3064 ( .A1(n2890), .A2(n3074), .ZN(n2417) );
  NAND2_X1 U3065 ( .A1(n3063), .A2(n2417), .ZN(n2419) );
  OR2_X1 U3066 ( .A1(n2890), .A2(n3074), .ZN(n2418) );
  NAND2_X1 U3067 ( .A1(n2411), .A2(REG2_REG_4__SCAN_IN), .ZN(n2431) );
  INV_X1 U3068 ( .A(n2420), .ZN(n3682) );
  INV_X2 U3069 ( .A(n3682), .ZN(n2794) );
  INV_X1 U3070 ( .A(REG0_REG_4__SCAN_IN), .ZN(n2421) );
  INV_X1 U3071 ( .A(REG1_REG_4__SCAN_IN), .ZN(n2422) );
  OR2_X1 U3072 ( .A1(n2405), .A2(n2422), .ZN(n2429) );
  CLKBUF_X3 U3073 ( .A(n2423), .Z(n2716) );
  INV_X1 U3074 ( .A(n2437), .ZN(n2427) );
  INV_X1 U3075 ( .A(REG3_REG_4__SCAN_IN), .ZN(n2425) );
  INV_X1 U3076 ( .A(REG3_REG_3__SCAN_IN), .ZN(n2424) );
  NAND2_X1 U3077 ( .A1(n2425), .A2(n2424), .ZN(n2426) );
  NAND2_X1 U3078 ( .A1(n2427), .A2(n2426), .ZN(n3017) );
  OR2_X1 U3079 ( .A1(n2716), .A2(n3017), .ZN(n2428) );
  NAND4_X4 U3080 ( .A1(n2431), .A2(n2430), .A3(n2429), .A4(n2428), .ZN(n3840)
         );
  NAND2_X1 U3081 ( .A1(n2432), .A2(IR_REG_31__SCAN_IN), .ZN(n2434) );
  XNOR2_X1 U3082 ( .A(n2434), .B(n2433), .ZN(n3877) );
  INV_X1 U3083 ( .A(DATAI_4_), .ZN(n4825) );
  MUX2_X1 U3084 ( .A(n3877), .B(n4825), .S(n3679), .Z(n3020) );
  OR2_X2 U3085 ( .A1(n3840), .A2(n3020), .ZN(n3762) );
  NAND2_X1 U3086 ( .A1(n3840), .A2(n3020), .ZN(n3765) );
  INV_X1 U3087 ( .A(n3020), .ZN(n3006) );
  NAND2_X1 U3088 ( .A1(n3840), .A2(n3006), .ZN(n2435) );
  NAND2_X1 U3089 ( .A1(n2411), .A2(REG2_REG_5__SCAN_IN), .ZN(n2441) );
  INV_X1 U3090 ( .A(REG0_REG_5__SCAN_IN), .ZN(n2436) );
  OR2_X1 U3091 ( .A1(n2794), .A2(n2436), .ZN(n2440) );
  INV_X1 U3092 ( .A(REG1_REG_5__SCAN_IN), .ZN(n2828) );
  OR2_X1 U3093 ( .A1(n3684), .A2(n2828), .ZN(n2439) );
  NAND2_X1 U3094 ( .A1(n2437), .A2(REG3_REG_5__SCAN_IN), .ZN(n2449) );
  OAI21_X1 U3095 ( .B1(n2437), .B2(REG3_REG_5__SCAN_IN), .A(n2449), .ZN(n3582)
         );
  OR2_X1 U3096 ( .A1(n2716), .A2(n3582), .ZN(n2438) );
  NAND4_X1 U3097 ( .A1(n2441), .A2(n2440), .A3(n2439), .A4(n2438), .ZN(n3059)
         );
  NAND2_X1 U3098 ( .A1(n2442), .A2(IR_REG_31__SCAN_IN), .ZN(n2443) );
  XNOR2_X1 U3099 ( .A(n2443), .B(IR_REG_5__SCAN_IN), .ZN(n2829) );
  MUX2_X1 U3100 ( .A(n2829), .B(DATAI_5_), .S(n3679), .Z(n3080) );
  OR2_X1 U3101 ( .A1(n3059), .A2(n3080), .ZN(n2444) );
  NAND2_X1 U3102 ( .A1(n3084), .A2(n2444), .ZN(n2446) );
  NAND2_X1 U3103 ( .A1(n3059), .A2(n3080), .ZN(n2445) );
  NAND2_X1 U3104 ( .A1(n2446), .A2(n2445), .ZN(n3027) );
  NAND2_X1 U3105 ( .A1(n2411), .A2(REG2_REG_6__SCAN_IN), .ZN(n2454) );
  INV_X1 U3106 ( .A(REG0_REG_6__SCAN_IN), .ZN(n2447) );
  OR2_X1 U3107 ( .A1(n2794), .A2(n2447), .ZN(n2453) );
  INV_X1 U3108 ( .A(REG1_REG_6__SCAN_IN), .ZN(n2448) );
  OR2_X1 U3109 ( .A1(n3684), .A2(n2448), .ZN(n2452) );
  AND2_X1 U3110 ( .A1(n2449), .A2(n4768), .ZN(n2450) );
  NOR2_X1 U3111 ( .A1(n2449), .A2(n4768), .ZN(n2460) );
  OR2_X1 U3112 ( .A1(n2450), .A2(n2460), .ZN(n3031) );
  OR2_X1 U3113 ( .A1(n2716), .A2(n3031), .ZN(n2451) );
  NAND4_X1 U3114 ( .A1(n2454), .A2(n2453), .A3(n2452), .A4(n2451), .ZN(n3584)
         );
  OR2_X1 U3115 ( .A1(n2455), .A2(n2357), .ZN(n2466) );
  INV_X1 U3116 ( .A(IR_REG_6__SCAN_IN), .ZN(n4606) );
  NAND2_X1 U3117 ( .A1(n2466), .A2(n4606), .ZN(n2457) );
  OR2_X1 U3118 ( .A1(n2455), .A2(n4817), .ZN(n2456) );
  MUX2_X1 U3119 ( .A(n4362), .B(DATAI_6_), .S(n3679), .Z(n3092) );
  AND2_X1 U3120 ( .A1(n3584), .A2(n3092), .ZN(n2458) );
  OAI22_X1 U3121 ( .A1(n3027), .A2(n2458), .B1(n3092), .B2(n3584), .ZN(n3134)
         );
  INV_X1 U3122 ( .A(n3134), .ZN(n2472) );
  NAND2_X1 U3123 ( .A1(n2411), .A2(REG2_REG_7__SCAN_IN), .ZN(n2465) );
  INV_X1 U3124 ( .A(REG0_REG_7__SCAN_IN), .ZN(n2459) );
  OR2_X1 U3125 ( .A1(n2794), .A2(n2459), .ZN(n2464) );
  INV_X1 U3126 ( .A(REG1_REG_7__SCAN_IN), .ZN(n2835) );
  OR2_X1 U3127 ( .A1(n3684), .A2(n2835), .ZN(n2463) );
  NAND2_X1 U3128 ( .A1(n2460), .A2(REG3_REG_7__SCAN_IN), .ZN(n2476) );
  OR2_X1 U3129 ( .A1(n2460), .A2(REG3_REG_7__SCAN_IN), .ZN(n2461) );
  NAND2_X1 U3130 ( .A1(n2476), .A2(n2461), .ZN(n3131) );
  OR2_X1 U3131 ( .A1(n2716), .A2(n3131), .ZN(n2462) );
  NAND4_X1 U3132 ( .A1(n2465), .A2(n2464), .A3(n2463), .A4(n2462), .ZN(n3839)
         );
  INV_X1 U3133 ( .A(IR_REG_7__SCAN_IN), .ZN(n2467) );
  NAND2_X1 U3134 ( .A1(n2468), .A2(n2467), .ZN(n2482) );
  INV_X1 U3135 ( .A(n2468), .ZN(n2469) );
  NAND2_X1 U3136 ( .A1(n2469), .A2(IR_REG_7__SCAN_IN), .ZN(n2470) );
  NAND2_X1 U3137 ( .A1(n2482), .A2(n2470), .ZN(n4360) );
  INV_X1 U3138 ( .A(DATAI_7_), .ZN(n4583) );
  MUX2_X1 U3139 ( .A(n4360), .B(n4583), .S(n3679), .Z(n3117) );
  OR2_X1 U3140 ( .A1(n3839), .A2(n3117), .ZN(n2684) );
  NAND2_X1 U3141 ( .A1(n3839), .A2(n3117), .ZN(n3776) );
  NAND2_X1 U3142 ( .A1(n3839), .A2(n3127), .ZN(n2473) );
  NAND2_X1 U3143 ( .A1(n2411), .A2(REG2_REG_8__SCAN_IN), .ZN(n2481) );
  INV_X1 U3144 ( .A(REG0_REG_8__SCAN_IN), .ZN(n2474) );
  OR2_X1 U3145 ( .A1(n2794), .A2(n2474), .ZN(n2480) );
  INV_X1 U3146 ( .A(REG1_REG_8__SCAN_IN), .ZN(n2475) );
  OR2_X1 U3147 ( .A1(n3684), .A2(n2475), .ZN(n2479) );
  NAND2_X1 U31480 ( .A1(n2476), .A2(n4597), .ZN(n2477) );
  NAND2_X1 U31490 ( .A1(n2487), .A2(n2477), .ZN(n3169) );
  OR2_X1 U3150 ( .A1(n2716), .A2(n3169), .ZN(n2478) );
  NAND4_X1 U3151 ( .A1(n2481), .A2(n2480), .A3(n2479), .A4(n2478), .ZN(n3838)
         );
  NAND2_X1 U3152 ( .A1(n2482), .A2(IR_REG_31__SCAN_IN), .ZN(n2483) );
  XNOR2_X1 U3153 ( .A(n2483), .B(IR_REG_8__SCAN_IN), .ZN(n2882) );
  MUX2_X1 U3154 ( .A(n2882), .B(DATAI_8_), .S(n3679), .Z(n3171) );
  OR2_X1 U3155 ( .A1(n3838), .A2(n3171), .ZN(n2484) );
  NAND2_X1 U3156 ( .A1(n3838), .A2(n3171), .ZN(n2485) );
  NAND2_X1 U3157 ( .A1(n2411), .A2(REG2_REG_9__SCAN_IN), .ZN(n2492) );
  INV_X1 U3158 ( .A(REG0_REG_9__SCAN_IN), .ZN(n2486) );
  OR2_X1 U3159 ( .A1(n2794), .A2(n2486), .ZN(n2491) );
  INV_X1 U3160 ( .A(REG1_REG_9__SCAN_IN), .ZN(n2884) );
  OR2_X1 U3161 ( .A1(n3684), .A2(n2884), .ZN(n2490) );
  AND2_X1 U3162 ( .A1(n2487), .A2(n4771), .ZN(n2488) );
  OR2_X1 U3163 ( .A1(n2488), .A2(n2500), .ZN(n3209) );
  OR2_X1 U3164 ( .A1(n2716), .A2(n3209), .ZN(n2489) );
  NAND4_X1 U3165 ( .A1(n2492), .A2(n2491), .A3(n2490), .A4(n2489), .ZN(n3297)
         );
  NAND2_X1 U3166 ( .A1(n2493), .A2(IR_REG_31__SCAN_IN), .ZN(n2494) );
  MUX2_X1 U3167 ( .A(IR_REG_31__SCAN_IN), .B(n2494), .S(IR_REG_9__SCAN_IN), 
        .Z(n2495) );
  AND2_X1 U3168 ( .A1(n2495), .A2(n2165), .ZN(n4359) );
  MUX2_X1 U3169 ( .A(n4359), .B(DATAI_9_), .S(n3679), .Z(n3208) );
  AND2_X1 U3170 ( .A1(n3297), .A2(n3208), .ZN(n2497) );
  OR2_X1 U3171 ( .A1(n3297), .A2(n3208), .ZN(n2496) );
  NAND2_X1 U3172 ( .A1(n2410), .A2(REG2_REG_10__SCAN_IN), .ZN(n2505) );
  INV_X1 U3173 ( .A(REG0_REG_10__SCAN_IN), .ZN(n2498) );
  OR2_X1 U3174 ( .A1(n2794), .A2(n2498), .ZN(n2504) );
  INV_X1 U3175 ( .A(REG1_REG_10__SCAN_IN), .ZN(n2499) );
  OR2_X1 U3176 ( .A1(n3684), .A2(n2499), .ZN(n2503) );
  NOR2_X1 U3177 ( .A1(n2500), .A2(REG3_REG_10__SCAN_IN), .ZN(n2501) );
  OR2_X1 U3178 ( .A1(n2507), .A2(n2501), .ZN(n3296) );
  OR2_X1 U3179 ( .A1(n2716), .A2(n3296), .ZN(n2502) );
  NAND4_X1 U3180 ( .A1(n2505), .A2(n2504), .A3(n2503), .A4(n2502), .ZN(n3285)
         );
  NAND2_X1 U3181 ( .A1(n2165), .A2(IR_REG_31__SCAN_IN), .ZN(n2506) );
  XNOR2_X1 U3182 ( .A(n2506), .B(IR_REG_10__SCAN_IN), .ZN(n3905) );
  MUX2_X1 U3183 ( .A(n3905), .B(DATAI_10_), .S(n3679), .Z(n3270) );
  NOR2_X1 U3184 ( .A1(n3285), .A2(n3270), .ZN(n3243) );
  NAND2_X1 U3185 ( .A1(n2411), .A2(REG2_REG_11__SCAN_IN), .ZN(n2512) );
  INV_X1 U3186 ( .A(REG0_REG_11__SCAN_IN), .ZN(n4847) );
  OR2_X1 U3187 ( .A1(n2794), .A2(n4847), .ZN(n2511) );
  INV_X1 U3188 ( .A(REG1_REG_11__SCAN_IN), .ZN(n4300) );
  OR2_X1 U3189 ( .A1(n3684), .A2(n4300), .ZN(n2510) );
  OR2_X1 U3190 ( .A1(n2507), .A2(REG3_REG_11__SCAN_IN), .ZN(n2508) );
  NAND2_X1 U3191 ( .A1(n2531), .A2(n2508), .ZN(n3256) );
  OR2_X1 U3192 ( .A1(n2716), .A2(n3256), .ZN(n2509) );
  NAND4_X1 U3193 ( .A1(n2512), .A2(n2511), .A3(n2510), .A4(n2509), .ZN(n3279)
         );
  NAND2_X1 U3194 ( .A1(n2513), .A2(IR_REG_31__SCAN_IN), .ZN(n2522) );
  XNOR2_X1 U3195 ( .A(n2522), .B(IR_REG_11__SCAN_IN), .ZN(n3901) );
  INV_X1 U3196 ( .A(DATAI_11_), .ZN(n2514) );
  MUX2_X1 U3197 ( .A(n4501), .B(n2514), .S(n3679), .Z(n3287) );
  OR2_X1 U3198 ( .A1(n3279), .A2(n3287), .ZN(n3787) );
  NAND2_X1 U3199 ( .A1(n3279), .A2(n3287), .ZN(n3786) );
  NAND2_X1 U3200 ( .A1(n3787), .A2(n3786), .ZN(n3718) );
  INV_X1 U3201 ( .A(n3718), .ZN(n3241) );
  INV_X1 U3202 ( .A(n3285), .ZN(n3249) );
  OR2_X1 U3203 ( .A1(n3279), .A2(n3252), .ZN(n2516) );
  NAND2_X1 U3204 ( .A1(n3245), .A2(n2516), .ZN(n3234) );
  NAND2_X1 U3205 ( .A1(n2410), .A2(REG2_REG_12__SCAN_IN), .ZN(n2521) );
  INV_X1 U3206 ( .A(REG0_REG_12__SCAN_IN), .ZN(n2517) );
  OR2_X1 U3207 ( .A1(n2794), .A2(n2517), .ZN(n2520) );
  INV_X1 U3208 ( .A(REG1_REG_12__SCAN_IN), .ZN(n4692) );
  OR2_X1 U3209 ( .A1(n3684), .A2(n4692), .ZN(n2519) );
  XNOR2_X1 U32100 ( .A(n2531), .B(n2530), .ZN(n3318) );
  OR2_X1 U32110 ( .A1(n2716), .A2(n3318), .ZN(n2518) );
  NAND4_X1 U32120 ( .A1(n2521), .A2(n2520), .A3(n2519), .A4(n2518), .ZN(n3837)
         );
  NAND2_X1 U32130 ( .A1(n2522), .A2(n4821), .ZN(n2523) );
  NAND2_X1 U32140 ( .A1(n2523), .A2(IR_REG_31__SCAN_IN), .ZN(n2524) );
  XNOR2_X1 U32150 ( .A(n2524), .B(IR_REG_12__SCAN_IN), .ZN(n3909) );
  MUX2_X1 U32160 ( .A(n3909), .B(DATAI_12_), .S(n3679), .Z(n4287) );
  NAND2_X1 U32170 ( .A1(n3837), .A2(n4287), .ZN(n2525) );
  NAND2_X1 U32180 ( .A1(n3234), .A2(n2525), .ZN(n2527) );
  OR2_X1 U32190 ( .A1(n3837), .A2(n4287), .ZN(n2526) );
  NAND2_X1 U32200 ( .A1(n2527), .A2(n2526), .ZN(n3323) );
  INV_X1 U32210 ( .A(n3323), .ZN(n2538) );
  NAND2_X1 U32220 ( .A1(n2410), .A2(REG2_REG_13__SCAN_IN), .ZN(n2536) );
  INV_X1 U32230 ( .A(REG0_REG_13__SCAN_IN), .ZN(n2528) );
  OR2_X1 U32240 ( .A1(n2794), .A2(n2528), .ZN(n2535) );
  INV_X1 U32250 ( .A(REG1_REG_13__SCAN_IN), .ZN(n3892) );
  OR2_X1 U32260 ( .A1(n3684), .A2(n3892), .ZN(n2534) );
  OAI21_X1 U32270 ( .B1(n2531), .B2(n2530), .A(n2529), .ZN(n2532) );
  NAND2_X1 U32280 ( .A1(n2532), .A2(n2539), .ZN(n3338) );
  OR2_X1 U32290 ( .A1(n2716), .A2(n3338), .ZN(n2533) );
  NAND4_X1 U32300 ( .A1(n2536), .A2(n2535), .A3(n2534), .A4(n2533), .ZN(n4290)
         );
  OR2_X1 U32310 ( .A1(n2545), .A2(n2357), .ZN(n2537) );
  XNOR2_X1 U32320 ( .A(n2537), .B(IR_REG_13__SCAN_IN), .ZN(n3912) );
  MUX2_X1 U32330 ( .A(n3912), .B(DATAI_13_), .S(n3679), .Z(n3396) );
  AOI21_X1 U32340 ( .B1(n2538), .B2(n2345), .A(n2344), .ZN(n3344) );
  NAND2_X1 U32350 ( .A1(n2410), .A2(REG2_REG_14__SCAN_IN), .ZN(n2544) );
  INV_X1 U32360 ( .A(REG0_REG_14__SCAN_IN), .ZN(n4680) );
  OR2_X1 U32370 ( .A1(n2794), .A2(n4680), .ZN(n2543) );
  INV_X1 U32380 ( .A(REG1_REG_14__SCAN_IN), .ZN(n4849) );
  OR2_X1 U32390 ( .A1(n3684), .A2(n4849), .ZN(n2542) );
  AND2_X1 U32400 ( .A1(n2539), .A2(n4805), .ZN(n2540) );
  OR2_X1 U32410 ( .A1(n2540), .A2(n2560), .ZN(n3497) );
  OR2_X1 U32420 ( .A1(n2716), .A2(n3497), .ZN(n2541) );
  NAND4_X1 U32430 ( .A1(n2544), .A2(n2543), .A3(n2542), .A4(n2541), .ZN(n4186)
         );
  NAND2_X1 U32440 ( .A1(n2579), .A2(IR_REG_31__SCAN_IN), .ZN(n2546) );
  XNOR2_X1 U32450 ( .A(n2546), .B(IR_REG_14__SCAN_IN), .ZN(n4427) );
  INV_X1 U32460 ( .A(DATAI_14_), .ZN(n2547) );
  MUX2_X1 U32470 ( .A(n4497), .B(n2547), .S(n3679), .Z(n4274) );
  OR2_X1 U32480 ( .A1(n4186), .A2(n4274), .ZN(n3687) );
  NAND2_X1 U32490 ( .A1(n4186), .A2(n4274), .ZN(n3688) );
  NAND2_X1 U32500 ( .A1(n3687), .A2(n3688), .ZN(n3719) );
  NAND2_X1 U32510 ( .A1(n3344), .A2(n3719), .ZN(n3343) );
  OR2_X1 U32520 ( .A1(n4186), .A2(n3500), .ZN(n2548) );
  NAND2_X1 U32530 ( .A1(n3343), .A2(n2548), .ZN(n4177) );
  NAND2_X1 U32540 ( .A1(n2410), .A2(REG2_REG_15__SCAN_IN), .ZN(n2553) );
  INV_X1 U32550 ( .A(REG0_REG_15__SCAN_IN), .ZN(n2549) );
  OR2_X1 U32560 ( .A1(n2794), .A2(n2549), .ZN(n2552) );
  INV_X1 U32570 ( .A(REG1_REG_15__SCAN_IN), .ZN(n4850) );
  OR2_X1 U32580 ( .A1(n3684), .A2(n4850), .ZN(n2551) );
  XNOR2_X1 U32590 ( .A(n2560), .B(REG3_REG_15__SCAN_IN), .ZN(n3665) );
  OR2_X1 U32600 ( .A1(n2716), .A2(n3665), .ZN(n2550) );
  NAND4_X1 U32610 ( .A1(n2553), .A2(n2552), .A3(n2551), .A4(n2550), .ZN(n3415)
         );
  OR2_X1 U32620 ( .A1(n2579), .A2(IR_REG_14__SCAN_IN), .ZN(n2554) );
  NAND2_X1 U32630 ( .A1(n2554), .A2(IR_REG_31__SCAN_IN), .ZN(n2566) );
  MUX2_X1 U32640 ( .A(n4440), .B(DATAI_15_), .S(n3679), .Z(n4181) );
  NAND2_X1 U32650 ( .A1(n3415), .A2(n4181), .ZN(n2556) );
  NOR2_X1 U32660 ( .A1(n3415), .A2(n4181), .ZN(n2555) );
  NAND2_X1 U32670 ( .A1(n2410), .A2(REG2_REG_16__SCAN_IN), .ZN(n2565) );
  INV_X1 U32680 ( .A(REG0_REG_16__SCAN_IN), .ZN(n4679) );
  OR2_X1 U32690 ( .A1(n2794), .A2(n4679), .ZN(n2564) );
  INV_X1 U32700 ( .A(REG1_REG_16__SCAN_IN), .ZN(n4450) );
  OR2_X1 U32710 ( .A1(n3684), .A2(n4450), .ZN(n2563) );
  NAND2_X1 U32720 ( .A1(n2560), .A2(REG3_REG_15__SCAN_IN), .ZN(n2558) );
  INV_X1 U32730 ( .A(REG3_REG_16__SCAN_IN), .ZN(n2557) );
  NAND2_X1 U32740 ( .A1(n2558), .A2(n2557), .ZN(n2561) );
  AND2_X1 U32750 ( .A1(REG3_REG_16__SCAN_IN), .A2(REG3_REG_15__SCAN_IN), .ZN(
        n2559) );
  NAND2_X1 U32760 ( .A1(n2560), .A2(n2559), .ZN(n2570) );
  NAND2_X1 U32770 ( .A1(n2561), .A2(n2570), .ZN(n4170) );
  OR2_X1 U32780 ( .A1(n2716), .A2(n4170), .ZN(n2562) );
  NAND4_X1 U32790 ( .A1(n2565), .A2(n2564), .A3(n2563), .A4(n2562), .ZN(n4179)
         );
  NAND2_X1 U32800 ( .A1(n2566), .A2(n2577), .ZN(n2567) );
  NAND2_X1 U32810 ( .A1(n2567), .A2(IR_REG_31__SCAN_IN), .ZN(n2568) );
  INV_X1 U32820 ( .A(DATAI_16_), .ZN(n4493) );
  MUX2_X1 U32830 ( .A(n4494), .B(n4493), .S(n3679), .Z(n4260) );
  OR2_X1 U32840 ( .A1(n4179), .A2(n4260), .ZN(n3797) );
  NAND2_X1 U32850 ( .A1(n4179), .A2(n4260), .ZN(n3799) );
  NAND2_X1 U32860 ( .A1(n3797), .A2(n3799), .ZN(n4160) );
  NAND2_X1 U32870 ( .A1(n4161), .A2(n4160), .ZN(n4159) );
  NAND2_X1 U32880 ( .A1(n4179), .A2(n2223), .ZN(n2569) );
  NAND2_X1 U32890 ( .A1(n4159), .A2(n2569), .ZN(n4143) );
  NAND2_X1 U32900 ( .A1(n2410), .A2(REG2_REG_17__SCAN_IN), .ZN(n2575) );
  INV_X1 U32910 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4334) );
  OR2_X1 U32920 ( .A1(n2794), .A2(n4334), .ZN(n2574) );
  INV_X1 U32930 ( .A(REG1_REG_17__SCAN_IN), .ZN(n4858) );
  OR2_X1 U32940 ( .A1(n3684), .A2(n4858), .ZN(n2573) );
  NAND2_X1 U32950 ( .A1(n2570), .A2(n4599), .ZN(n2571) );
  NAND2_X1 U32960 ( .A1(n2584), .A2(n2571), .ZN(n4153) );
  OR2_X1 U32970 ( .A1(n2716), .A2(n4153), .ZN(n2572) );
  NAND4_X1 U32980 ( .A1(n2575), .A2(n2574), .A3(n2573), .A4(n2572), .ZN(n3642)
         );
  NAND3_X1 U32990 ( .A1(n2577), .A2(n4608), .A3(n2576), .ZN(n2578) );
  NOR2_X2 U33000 ( .A1(n2579), .A2(n2578), .ZN(n2591) );
  OR2_X1 U33010 ( .A1(n2591), .A2(n2357), .ZN(n2580) );
  MUX2_X1 U33020 ( .A(n3918), .B(DATAI_17_), .S(n3679), .Z(n3598) );
  NAND2_X1 U33030 ( .A1(n3642), .A2(n3598), .ZN(n2582) );
  NAND2_X1 U33040 ( .A1(n2410), .A2(REG2_REG_18__SCAN_IN), .ZN(n2589) );
  INV_X1 U33050 ( .A(REG0_REG_18__SCAN_IN), .ZN(n2583) );
  OR2_X1 U33060 ( .A1(n2794), .A2(n2583), .ZN(n2588) );
  INV_X1 U33070 ( .A(REG1_REG_18__SCAN_IN), .ZN(n4695) );
  OR2_X1 U33080 ( .A1(n3684), .A2(n4695), .ZN(n2587) );
  AND2_X1 U33090 ( .A1(n2584), .A2(n3643), .ZN(n2585) );
  OR2_X1 U33100 ( .A1(n2585), .A2(n2595), .ZN(n3641) );
  OR2_X1 U33110 ( .A1(n2716), .A2(n3641), .ZN(n2586) );
  NAND4_X1 U33120 ( .A1(n2589), .A2(n2588), .A3(n2587), .A4(n2586), .ZN(n4113)
         );
  NAND2_X1 U33130 ( .A1(n2591), .A2(n2590), .ZN(n2601) );
  NAND2_X1 U33140 ( .A1(n2601), .A2(IR_REG_31__SCAN_IN), .ZN(n2592) );
  XNOR2_X1 U33150 ( .A(n2592), .B(IR_REG_18__SCAN_IN), .ZN(n3919) );
  INV_X1 U33160 ( .A(DATAI_18_), .ZN(n2593) );
  MUX2_X1 U33170 ( .A(n4490), .B(n2593), .S(n3679), .Z(n4134) );
  OR2_X1 U33180 ( .A1(n4113), .A2(n4134), .ZN(n4106) );
  NAND2_X1 U33190 ( .A1(n4113), .A2(n4134), .ZN(n4107) );
  NAND2_X1 U33200 ( .A1(n4106), .A2(n4107), .ZN(n3720) );
  OR2_X1 U33210 ( .A1(n4113), .A2(n4124), .ZN(n2594) );
  NAND2_X1 U33220 ( .A1(n2410), .A2(REG2_REG_19__SCAN_IN), .ZN(n2600) );
  INV_X1 U33230 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4329) );
  OR2_X1 U33240 ( .A1(n2794), .A2(n4329), .ZN(n2599) );
  INV_X1 U33250 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4252) );
  OR2_X1 U33260 ( .A1(n3684), .A2(n4252), .ZN(n2598) );
  NOR2_X1 U33270 ( .A1(n2595), .A2(REG3_REG_19__SCAN_IN), .ZN(n2596) );
  OR2_X1 U33280 ( .A1(n2606), .A2(n2596), .ZN(n4118) );
  OR2_X1 U33290 ( .A1(n2716), .A2(n4118), .ZN(n2597) );
  NAND4_X1 U33300 ( .A1(n2600), .A2(n2599), .A3(n2598), .A4(n2597), .ZN(n4125)
         );
  INV_X1 U33310 ( .A(n2601), .ZN(n2603) );
  NAND2_X1 U33320 ( .A1(n2603), .A2(n2602), .ZN(n2604) );
  MUX2_X1 U33330 ( .A(n4358), .B(DATAI_19_), .S(n3679), .Z(n3522) );
  NOR2_X1 U33340 ( .A1(n4125), .A2(n3522), .ZN(n4086) );
  NAND2_X1 U33350 ( .A1(n2410), .A2(REG2_REG_20__SCAN_IN), .ZN(n2611) );
  INV_X1 U33360 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4848) );
  OR2_X1 U33370 ( .A1(n2794), .A2(n4848), .ZN(n2610) );
  INV_X1 U33380 ( .A(REG1_REG_20__SCAN_IN), .ZN(n2605) );
  OR2_X1 U33390 ( .A1(n3684), .A2(n2605), .ZN(n2609) );
  OR2_X1 U33400 ( .A1(n2606), .A2(REG3_REG_20__SCAN_IN), .ZN(n2607) );
  NAND2_X1 U33410 ( .A1(n2613), .A2(n2607), .ZN(n4096) );
  OR2_X1 U33420 ( .A1(n2716), .A2(n4096), .ZN(n2608) );
  NAND4_X1 U33430 ( .A1(n2611), .A2(n2610), .A3(n2609), .A4(n2608), .ZN(n3836)
         );
  NAND2_X1 U33440 ( .A1(n3836), .A2(n4095), .ZN(n3738) );
  NAND2_X1 U33450 ( .A1(n4125), .A2(n3522), .ZN(n4085) );
  OAI211_X1 U33460 ( .C1(n4103), .C2(n4086), .A(n3738), .B(n4085), .ZN(n2612)
         );
  NAND2_X1 U33470 ( .A1(n4111), .A2(n3441), .ZN(n3739) );
  NAND2_X1 U33480 ( .A1(n2612), .A2(n3739), .ZN(n4065) );
  NAND2_X1 U33490 ( .A1(n2411), .A2(REG2_REG_21__SCAN_IN), .ZN(n2619) );
  INV_X1 U33500 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4682) );
  OR2_X1 U33510 ( .A1(n2794), .A2(n4682), .ZN(n2618) );
  INV_X1 U33520 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4704) );
  OR2_X1 U3353 ( .A1(n3684), .A2(n4704), .ZN(n2617) );
  NAND2_X1 U33540 ( .A1(n2613), .A2(n4596), .ZN(n2615) );
  INV_X1 U3355 ( .A(n2628), .ZN(n2614) );
  NAND2_X1 U3356 ( .A1(n2615), .A2(n2614), .ZN(n4071) );
  OR2_X1 U3357 ( .A1(n2716), .A2(n4071), .ZN(n2616) );
  NAND4_X1 U3358 ( .A1(n2619), .A2(n2618), .A3(n2617), .A4(n2616), .ZN(n4082)
         );
  NAND2_X1 U3359 ( .A1(n4082), .A2(n4074), .ZN(n2621) );
  INV_X1 U3360 ( .A(n4082), .ZN(n3631) );
  AOI21_X2 U3361 ( .B1(n4065), .B2(n2621), .A(n2620), .ZN(n4049) );
  NAND2_X1 U3362 ( .A1(n2411), .A2(REG2_REG_22__SCAN_IN), .ZN(n2626) );
  XNOR2_X1 U3363 ( .A(REG3_REG_22__SCAN_IN), .B(n2628), .ZN(n4051) );
  OR2_X1 U3364 ( .A1(n2716), .A2(n4051), .ZN(n2625) );
  INV_X1 U3365 ( .A(REG1_REG_22__SCAN_IN), .ZN(n2622) );
  OR2_X1 U3366 ( .A1(n3684), .A2(n2622), .ZN(n2624) );
  INV_X1 U3367 ( .A(REG0_REG_22__SCAN_IN), .ZN(n4845) );
  OR2_X1 U3368 ( .A1(n2794), .A2(n4845), .ZN(n2623) );
  NAND4_X1 U3369 ( .A1(n2626), .A2(n2625), .A3(n2624), .A4(n2623), .ZN(n4036)
         );
  OR2_X1 U3370 ( .A1(n4036), .A2(n4060), .ZN(n4030) );
  NAND2_X1 U3371 ( .A1(n4036), .A2(n4060), .ZN(n2701) );
  NAND2_X1 U3372 ( .A1(n4030), .A2(n2701), .ZN(n4055) );
  NAND2_X1 U3373 ( .A1(n2410), .A2(REG2_REG_23__SCAN_IN), .ZN(n2634) );
  INV_X1 U3374 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4322) );
  OR2_X1 U3375 ( .A1(n2794), .A2(n4322), .ZN(n2633) );
  INV_X1 U3376 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4703) );
  OR2_X1 U3377 ( .A1(n3684), .A2(n4703), .ZN(n2632) );
  NAND3_X1 U3378 ( .A1(REG3_REG_22__SCAN_IN), .A2(REG3_REG_23__SCAN_IN), .A3(
        n2628), .ZN(n2636) );
  INV_X1 U3379 ( .A(REG3_REG_23__SCAN_IN), .ZN(n4810) );
  NAND2_X1 U3380 ( .A1(REG3_REG_22__SCAN_IN), .A2(n2628), .ZN(n2629) );
  NAND2_X1 U3381 ( .A1(n4810), .A2(n2629), .ZN(n2630) );
  NAND2_X1 U3382 ( .A1(n2636), .A2(n2630), .ZN(n4042) );
  OR2_X1 U3383 ( .A1(n2716), .A2(n4042), .ZN(n2631) );
  NAND2_X1 U3384 ( .A1(n2411), .A2(REG2_REG_24__SCAN_IN), .ZN(n2641) );
  INV_X1 U3385 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4318) );
  OR2_X1 U3386 ( .A1(n2794), .A2(n4318), .ZN(n2640) );
  INV_X1 U3387 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4229) );
  OR2_X1 U3388 ( .A1(n3684), .A2(n4229), .ZN(n2639) );
  AND2_X1 U3389 ( .A1(n2636), .A2(n4600), .ZN(n2637) );
  OR2_X1 U3390 ( .A1(n2637), .A2(n2642), .ZN(n4012) );
  NAND4_X1 U3391 ( .A1(n2641), .A2(n2640), .A3(n2639), .A4(n2638), .ZN(n3990)
         );
  NAND2_X1 U3392 ( .A1(n2411), .A2(REG2_REG_25__SCAN_IN), .ZN(n2647) );
  INV_X1 U3393 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4222) );
  OR2_X1 U3394 ( .A1(n3684), .A2(n4222), .ZN(n2646) );
  NOR2_X1 U3395 ( .A1(n2642), .A2(REG3_REG_25__SCAN_IN), .ZN(n2643) );
  INV_X1 U3396 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4314) );
  OR2_X1 U3397 ( .A1(n2794), .A2(n4314), .ZN(n2644) );
  NAND2_X1 U3398 ( .A1(n3985), .A2(n2648), .ZN(n2650) );
  NAND2_X1 U3399 ( .A1(n2411), .A2(REG2_REG_26__SCAN_IN), .ZN(n2654) );
  INV_X1 U3400 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4310) );
  OR2_X1 U3401 ( .A1(n2794), .A2(n4310), .ZN(n2653) );
  INV_X1 U3402 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4859) );
  OR2_X1 U3403 ( .A1(n3684), .A2(n4859), .ZN(n2652) );
  XNOR2_X1 U3404 ( .A(n2657), .B(REG3_REG_26__SCAN_IN), .ZN(n3979) );
  INV_X1 U3405 ( .A(n3978), .ZN(n3658) );
  NAND2_X1 U3406 ( .A1(n2411), .A2(REG2_REG_27__SCAN_IN), .ZN(n2662) );
  INV_X1 U3407 ( .A(REG0_REG_27__SCAN_IN), .ZN(n4684) );
  OR2_X1 U3408 ( .A1(n2794), .A2(n4684), .ZN(n2661) );
  INV_X1 U3409 ( .A(REG1_REG_27__SCAN_IN), .ZN(n4706) );
  OR2_X1 U3410 ( .A1(n3684), .A2(n4706), .ZN(n2660) );
  AND2_X1 U3411 ( .A1(REG3_REG_27__SCAN_IN), .A2(REG3_REG_26__SCAN_IN), .ZN(
        n2656) );
  AOI21_X1 U3412 ( .B1(n2657), .B2(REG3_REG_26__SCAN_IN), .A(
        REG3_REG_27__SCAN_IN), .ZN(n2658) );
  INV_X1 U3413 ( .A(n3972), .ZN(n3652) );
  NAND2_X2 U3414 ( .A1(n2663), .A2(n2338), .ZN(n3931) );
  NAND2_X1 U3415 ( .A1(n2411), .A2(REG2_REG_28__SCAN_IN), .ZN(n2670) );
  INV_X1 U3416 ( .A(REG0_REG_28__SCAN_IN), .ZN(n4846) );
  OR2_X1 U3417 ( .A1(n2794), .A2(n4846), .ZN(n2669) );
  INV_X1 U3418 ( .A(REG1_REG_28__SCAN_IN), .ZN(n2664) );
  OR2_X1 U3419 ( .A1(n3684), .A2(n2664), .ZN(n2668) );
  NAND2_X1 U3420 ( .A1(n2665), .A2(REG3_REG_28__SCAN_IN), .ZN(n3945) );
  OR2_X1 U3421 ( .A1(n2665), .A2(REG3_REG_28__SCAN_IN), .ZN(n2666) );
  NAND2_X1 U3422 ( .A1(n3945), .A2(n2666), .ZN(n3540) );
  OR2_X1 U3423 ( .A1(n2716), .A2(n3540), .ZN(n2667) );
  NAND4_X1 U3424 ( .A1(n2670), .A2(n2669), .A3(n2668), .A4(n2667), .ZN(n3938)
         );
  NAND2_X1 U3425 ( .A1(n3679), .A2(DATAI_28_), .ZN(n2754) );
  OR2_X1 U3426 ( .A1(n3938), .A2(n2754), .ZN(n3933) );
  NAND2_X1 U3427 ( .A1(n3938), .A2(n2754), .ZN(n3680) );
  NAND2_X1 U3428 ( .A1(n3933), .A2(n3680), .ZN(n3930) );
  OAI21_X1 U3429 ( .B1(IR_REG_19__SCAN_IN), .B2(IR_REG_20__SCAN_IN), .A(
        IR_REG_31__SCAN_IN), .ZN(n2672) );
  NAND2_X1 U3430 ( .A1(n2673), .A2(n2672), .ZN(n2722) );
  NAND2_X1 U3431 ( .A1(n2148), .A2(IR_REG_31__SCAN_IN), .ZN(n2674) );
  XNOR2_X1 U3432 ( .A(n2892), .B(n4356), .ZN(n2675) );
  NAND2_X1 U3433 ( .A1(n2675), .A2(n4555), .ZN(n4554) );
  INV_X1 U3434 ( .A(n2677), .ZN(n3747) );
  OR2_X1 U3435 ( .A1(n2897), .A2(n4563), .ZN(n3357) );
  INV_X1 U3436 ( .A(n3357), .ZN(n3755) );
  NAND2_X1 U3437 ( .A1(n3747), .A2(n3755), .ZN(n2975) );
  NAND2_X1 U3438 ( .A1(n2975), .A2(n2678), .ZN(n2680) );
  INV_X1 U3439 ( .A(n3722), .ZN(n2679) );
  NAND2_X1 U3440 ( .A1(n2680), .A2(n2679), .ZN(n2954) );
  NAND2_X1 U3441 ( .A1(n2954), .A2(n3756), .ZN(n3065) );
  INV_X1 U3442 ( .A(n3074), .ZN(n2681) );
  OR2_X1 U3443 ( .A1(n2890), .A2(n2681), .ZN(n3761) );
  NAND2_X1 U3444 ( .A1(n2890), .A2(n2681), .ZN(n3758) );
  NAND2_X1 U3445 ( .A1(n3761), .A2(n3758), .ZN(n3721) );
  INV_X1 U3446 ( .A(n3721), .ZN(n3066) );
  NAND2_X1 U3447 ( .A1(n3065), .A2(n3066), .ZN(n3064) );
  NAND2_X1 U3448 ( .A1(n3064), .A2(n3761), .ZN(n2993) );
  INV_X1 U3449 ( .A(n3762), .ZN(n2682) );
  OR2_X1 U3450 ( .A1(n3059), .A2(n3585), .ZN(n3774) );
  NAND2_X1 U3451 ( .A1(n3059), .A2(n3585), .ZN(n3764) );
  INV_X1 U3452 ( .A(n3092), .ZN(n3056) );
  AND2_X1 U3453 ( .A1(n3584), .A2(n3056), .ZN(n3024) );
  OR2_X1 U3454 ( .A1(n3025), .A2(n3024), .ZN(n2683) );
  OR2_X1 U3455 ( .A1(n3584), .A2(n3056), .ZN(n3767) );
  NAND2_X1 U3456 ( .A1(n2683), .A2(n3767), .ZN(n3123) );
  INV_X1 U3457 ( .A(n2684), .ZN(n2685) );
  OR2_X1 U34580 ( .A1(n3838), .A2(n3192), .ZN(n3771) );
  NAND2_X1 U34590 ( .A1(n3838), .A2(n3192), .ZN(n3775) );
  OR2_X1 U3460 ( .A1(n3297), .A2(n3211), .ZN(n3772) );
  NAND2_X1 U3461 ( .A1(n2686), .A2(n3772), .ZN(n3217) );
  NAND2_X1 U3462 ( .A1(n3285), .A2(n3299), .ZN(n3785) );
  NAND2_X1 U3463 ( .A1(n3217), .A2(n3785), .ZN(n2687) );
  OR2_X1 U3464 ( .A1(n3285), .A2(n3299), .ZN(n3781) );
  NAND2_X1 U3465 ( .A1(n2687), .A2(n3781), .ZN(n3242) );
  NAND2_X1 U3466 ( .A1(n3242), .A2(n3786), .ZN(n2688) );
  NAND2_X1 U34670 ( .A1(n2688), .A2(n3787), .ZN(n3329) );
  INV_X1 U3468 ( .A(n4287), .ZN(n2689) );
  NAND2_X1 U34690 ( .A1(n3837), .A2(n2689), .ZN(n3327) );
  NAND2_X1 U3470 ( .A1(n4290), .A2(n3624), .ZN(n3324) );
  NAND2_X1 U34710 ( .A1(n3329), .A2(n3791), .ZN(n2690) );
  NOR2_X1 U3472 ( .A1(n3837), .A2(n2689), .ZN(n3328) );
  NOR2_X1 U34730 ( .A1(n4290), .A2(n3624), .ZN(n3326) );
  AOI21_X1 U3474 ( .B1(n3791), .B2(n3328), .A(n3326), .ZN(n3788) );
  NAND2_X1 U34750 ( .A1(n2690), .A2(n3788), .ZN(n3691) );
  INV_X1 U3476 ( .A(n3719), .ZN(n2691) );
  NAND2_X1 U34770 ( .A1(n3691), .A2(n2691), .ZN(n2692) );
  NAND2_X1 U3478 ( .A1(n2692), .A2(n3687), .ZN(n4185) );
  INV_X1 U34790 ( .A(n4181), .ZN(n4267) );
  OR2_X1 U3480 ( .A1(n3415), .A2(n4267), .ZN(n3690) );
  NAND2_X1 U34810 ( .A1(n3415), .A2(n4267), .ZN(n3689) );
  NAND2_X1 U3482 ( .A1(n3690), .A2(n3689), .ZN(n4184) );
  INV_X1 U34830 ( .A(n4160), .ZN(n4164) );
  INV_X1 U3484 ( .A(n3522), .ZN(n4117) );
  NAND2_X1 U34850 ( .A1(n4125), .A2(n4117), .ZN(n2693) );
  AND2_X1 U3486 ( .A1(n4107), .A2(n2693), .ZN(n2698) );
  OR2_X1 U34870 ( .A1(n3642), .A2(n4151), .ZN(n4104) );
  NAND2_X1 U3488 ( .A1(n4106), .A2(n4104), .ZN(n2695) );
  NOR2_X1 U34890 ( .A1(n4125), .A2(n4117), .ZN(n2694) );
  AOI21_X1 U3490 ( .B1(n2698), .B2(n2695), .A(n2694), .ZN(n4079) );
  NAND2_X1 U34910 ( .A1(n4111), .A2(n4095), .ZN(n2696) );
  NAND2_X1 U3492 ( .A1(n4079), .A2(n2696), .ZN(n2697) );
  NAND2_X1 U34930 ( .A1(n3836), .A2(n3441), .ZN(n4025) );
  NAND2_X1 U3494 ( .A1(n2697), .A2(n4025), .ZN(n4026) );
  OR2_X1 U34950 ( .A1(n4082), .A2(n4238), .ZN(n4028) );
  AND2_X1 U3496 ( .A1(n4030), .A2(n4028), .ZN(n3808) );
  INV_X1 U34970 ( .A(n2698), .ZN(n4024) );
  NAND2_X1 U3498 ( .A1(n3642), .A2(n4151), .ZN(n4022) );
  NAND2_X1 U34990 ( .A1(n4025), .A2(n4022), .ZN(n2699) );
  NOR2_X1 U3500 ( .A1(n4024), .A2(n2699), .ZN(n3801) );
  OR2_X1 U35010 ( .A1(n2141), .A2(n3801), .ZN(n2703) );
  AND2_X1 U3502 ( .A1(n4082), .A2(n4238), .ZN(n3709) );
  NAND2_X1 U35030 ( .A1(n4057), .A2(n4033), .ZN(n2700) );
  NAND2_X1 U3504 ( .A1(n2701), .A2(n2700), .ZN(n3806) );
  AOI21_X1 U35050 ( .B1(n3709), .B2(n4030), .A(n3806), .ZN(n2702) );
  AND2_X1 U35060 ( .A1(n2703), .A2(n2702), .ZN(n3693) );
  NAND2_X1 U35070 ( .A1(n2704), .A2(n3693), .ZN(n4005) );
  OR2_X1 U35080 ( .A1(n3990), .A2(n4224), .ZN(n3732) );
  OR2_X1 U35090 ( .A1(n4057), .A2(n4033), .ZN(n4004) );
  NAND2_X1 U35100 ( .A1(n3732), .A2(n4004), .ZN(n3810) );
  INV_X1 U35110 ( .A(n3810), .ZN(n3696) );
  NAND2_X1 U35120 ( .A1(n4005), .A2(n3696), .ZN(n2705) );
  NAND2_X1 U35130 ( .A1(n3990), .A2(n4224), .ZN(n3731) );
  NAND2_X1 U35140 ( .A1(n2705), .A2(n3731), .ZN(n3987) );
  AND2_X1 U35150 ( .A1(n3973), .A2(n3993), .ZN(n3728) );
  OR2_X1 U35160 ( .A1(n3973), .A2(n3993), .ZN(n3967) );
  OR2_X1 U35170 ( .A1(n3961), .A2(n3978), .ZN(n3742) );
  AND2_X1 U35180 ( .A1(n3967), .A2(n3742), .ZN(n3816) );
  AND2_X1 U35190 ( .A1(n3961), .A2(n3978), .ZN(n3741) );
  AND2_X1 U35200 ( .A1(n3972), .A2(n4210), .ZN(n3814) );
  INV_X1 U35210 ( .A(n3814), .ZN(n2706) );
  OR2_X1 U35220 ( .A1(n3972), .A2(n4210), .ZN(n2707) );
  INV_X1 U35230 ( .A(n2707), .ZN(n3701) );
  NAND2_X1 U35240 ( .A1(n4357), .A2(n2708), .ZN(n3676) );
  NAND2_X1 U35250 ( .A1(n4358), .A2(n4356), .ZN(n2709) );
  AND2_X1 U35260 ( .A1(n2374), .A2(n2710), .ZN(n2712) );
  INV_X1 U35270 ( .A(n2712), .ZN(n2711) );
  INV_X1 U35280 ( .A(n2927), .ZN(n2713) );
  AND2_X1 U35290 ( .A1(n3972), .A2(n4187), .ZN(n2714) );
  AOI21_X1 U35300 ( .B1(n2715), .B2(n4162), .A(n2714), .ZN(n3382) );
  NAND2_X1 U35310 ( .A1(n2411), .A2(REG2_REG_29__SCAN_IN), .ZN(n2720) );
  INV_X1 U35320 ( .A(REG0_REG_29__SCAN_IN), .ZN(n4852) );
  OR2_X1 U35330 ( .A1(n2794), .A2(n4852), .ZN(n2719) );
  INV_X1 U35340 ( .A(REG1_REG_29__SCAN_IN), .ZN(n4701) );
  OR2_X1 U35350 ( .A1(n3684), .A2(n4701), .ZN(n2718) );
  OR2_X1 U35360 ( .A1(n2716), .A2(n3945), .ZN(n2717) );
  NAND4_X1 U35370 ( .A1(n2720), .A2(n2719), .A3(n2718), .A4(n2717), .ZN(n3835)
         );
  XOR2_X1 U35380 ( .A(n2722), .B(n2721), .Z(n2931) );
  INV_X1 U35390 ( .A(n4356), .ZN(n3828) );
  NAND2_X1 U35400 ( .A1(n2931), .A2(n3828), .ZN(n3356) );
  OR2_X1 U35410 ( .A1(n3356), .A2(n2756), .ZN(n4275) );
  AOI22_X1 U35420 ( .A1(n3835), .A2(n4289), .B1(n3929), .B2(n4288), .ZN(n2723)
         );
  NAND2_X1 U35430 ( .A1(n2756), .A2(n4555), .ZN(n2928) );
  NAND2_X1 U35440 ( .A1(n2928), .A2(n2927), .ZN(n2943) );
  OAI21_X1 U35450 ( .B1(IR_REG_23__SCAN_IN), .B2(IR_REG_24__SCAN_IN), .A(
        IR_REG_31__SCAN_IN), .ZN(n2727) );
  NAND2_X1 U35460 ( .A1(n2731), .A2(n2727), .ZN(n2729) );
  OR2_X1 U35470 ( .A1(n2731), .A2(n2730), .ZN(n2732) );
  NAND2_X1 U35480 ( .A1(n2749), .A2(n2774), .ZN(n2734) );
  MUX2_X1 U35490 ( .A(n2749), .B(n2734), .S(B_REG_SCAN_IN), .Z(n2735) );
  INV_X1 U35500 ( .A(D_REG_2__SCAN_IN), .ZN(n4639) );
  INV_X1 U35510 ( .A(D_REG_3__SCAN_IN), .ZN(n4638) );
  INV_X1 U35520 ( .A(D_REG_25__SCAN_IN), .ZN(n4664) );
  INV_X1 U35530 ( .A(D_REG_7__SCAN_IN), .ZN(n4634) );
  NAND4_X1 U35540 ( .A1(n4639), .A2(n4638), .A3(n4664), .A4(n4634), .ZN(n2736)
         );
  NOR4_X1 U35550 ( .A1(D_REG_13__SCAN_IN), .A2(D_REG_17__SCAN_IN), .A3(
        D_REG_22__SCAN_IN), .A4(n2736), .ZN(n4788) );
  NOR4_X1 U35560 ( .A1(D_REG_23__SCAN_IN), .A2(D_REG_15__SCAN_IN), .A3(
        D_REG_20__SCAN_IN), .A4(D_REG_16__SCAN_IN), .ZN(n2737) );
  INV_X1 U35570 ( .A(D_REG_14__SCAN_IN), .ZN(n4648) );
  INV_X1 U35580 ( .A(D_REG_11__SCAN_IN), .ZN(n4633) );
  NAND3_X1 U35590 ( .A1(n2737), .A2(n4648), .A3(n4633), .ZN(n2743) );
  NOR4_X1 U35600 ( .A1(D_REG_5__SCAN_IN), .A2(D_REG_6__SCAN_IN), .A3(
        D_REG_12__SCAN_IN), .A4(D_REG_9__SCAN_IN), .ZN(n2741) );
  NOR4_X1 U35610 ( .A1(D_REG_4__SCAN_IN), .A2(D_REG_28__SCAN_IN), .A3(
        D_REG_30__SCAN_IN), .A4(D_REG_8__SCAN_IN), .ZN(n2740) );
  NOR4_X1 U35620 ( .A1(D_REG_27__SCAN_IN), .A2(D_REG_24__SCAN_IN), .A3(
        D_REG_26__SCAN_IN), .A4(D_REG_29__SCAN_IN), .ZN(n2739) );
  NOR4_X1 U35630 ( .A1(D_REG_10__SCAN_IN), .A2(D_REG_21__SCAN_IN), .A3(
        D_REG_18__SCAN_IN), .A4(D_REG_19__SCAN_IN), .ZN(n2738) );
  NAND4_X1 U35640 ( .A1(n2741), .A2(n2740), .A3(n2739), .A4(n2738), .ZN(n2742)
         );
  NOR3_X1 U35650 ( .A1(D_REG_31__SCAN_IN), .A2(n2743), .A3(n2742), .ZN(n2744)
         );
  AND2_X1 U35660 ( .A1(n4788), .A2(n2744), .ZN(n2745) );
  OR2_X1 U35670 ( .A1(n2771), .A2(D_REG_1__SCAN_IN), .ZN(n2747) );
  INV_X1 U35680 ( .A(n4353), .ZN(n2772) );
  NAND2_X1 U35690 ( .A1(n2772), .A2(n2774), .ZN(n2746) );
  NAND2_X1 U35700 ( .A1(n2747), .A2(n2746), .ZN(n2967) );
  OAI21_X1 U35710 ( .B1(n2708), .B2(n4508), .A(n2967), .ZN(n2748) );
  NAND2_X1 U35720 ( .A1(n2749), .A2(n2772), .ZN(n2775) );
  INV_X1 U35730 ( .A(n4551), .ZN(n2751) );
  NAND2_X1 U35740 ( .A1(n2978), .A2(n4563), .ZN(n2972) );
  NAND2_X1 U35750 ( .A1(n3336), .A2(n3624), .ZN(n3345) );
  INV_X1 U35760 ( .A(n2752), .ZN(n3954) );
  INV_X1 U35770 ( .A(n3947), .ZN(n2753) );
  OAI21_X1 U35780 ( .B1(n3954), .B2(n2754), .A(n2753), .ZN(n3378) );
  INV_X1 U35790 ( .A(n3356), .ZN(n2755) );
  NAND2_X1 U35800 ( .A1(n2758), .A2(n2757), .ZN(U3546) );
  NAND2_X1 U35810 ( .A1(n2763), .A2(n2762), .ZN(U3514) );
  INV_X1 U3582 ( .A(n4488), .ZN(n2764) );
  INV_X2 U3583 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  INV_X1 U3584 ( .A(n2829), .ZN(n2872) );
  INV_X1 U3585 ( .A(DATAI_5_), .ZN(n2765) );
  MUX2_X1 U3586 ( .A(n2872), .B(n2765), .S(U3149), .Z(n2766) );
  INV_X1 U3587 ( .A(n2766), .ZN(U3347) );
  INV_X1 U3588 ( .A(DATAI_8_), .ZN(n2767) );
  INV_X1 U3589 ( .A(n2882), .ZN(n2840) );
  MUX2_X1 U3590 ( .A(n2767), .B(n2840), .S(STATE_REG_SCAN_IN), .Z(n2768) );
  INV_X1 U3591 ( .A(n2768), .ZN(U3344) );
  INV_X1 U3592 ( .A(IR_REG_30__SCAN_IN), .ZN(n4640) );
  NAND3_X1 U3593 ( .A1(IR_REG_31__SCAN_IN), .A2(STATE_REG_SCAN_IN), .A3(n4640), 
        .ZN(n2770) );
  INV_X1 U3594 ( .A(DATAI_31_), .ZN(n4835) );
  OAI22_X1 U3595 ( .A1(n2769), .A2(n2770), .B1(STATE_REG_SCAN_IN), .B2(n4835), 
        .ZN(U3321) );
  INV_X1 U3596 ( .A(D_REG_1__SCAN_IN), .ZN(n4836) );
  AND2_X1 U3597 ( .A1(n2772), .A2(n4488), .ZN(n2773) );
  AOI22_X1 U3598 ( .A1(n4486), .A2(n4836), .B1(n2774), .B2(n2773), .ZN(U3459)
         );
  INV_X1 U3599 ( .A(D_REG_0__SCAN_IN), .ZN(n4636) );
  INV_X1 U3600 ( .A(n2775), .ZN(n2776) );
  AOI22_X1 U3601 ( .A1(n4486), .A2(n4636), .B1(n2776), .B2(n4488), .ZN(U3458)
         );
  NOR2_X1 U3602 ( .A1(n2942), .A2(U3149), .ZN(n3829) );
  NOR2_X1 U3603 ( .A1(n2932), .A2(n3829), .ZN(n2799) );
  INV_X1 U3604 ( .A(n2799), .ZN(n2778) );
  NAND2_X1 U3605 ( .A1(n2927), .A2(n2942), .ZN(n2777) );
  NAND2_X1 U3606 ( .A1(n2777), .A2(n3679), .ZN(n2798) );
  NOR2_X1 U3607 ( .A1(n4473), .A2(U4043), .ZN(U3148) );
  INV_X1 U3608 ( .A(DATAO_REG_11__SCAN_IN), .ZN(n4790) );
  NAND2_X1 U3609 ( .A1(n3279), .A2(U4043), .ZN(n2779) );
  OAI21_X1 U3610 ( .B1(U4043), .B2(n4790), .A(n2779), .ZN(U3561) );
  INV_X1 U3611 ( .A(DATAO_REG_6__SCAN_IN), .ZN(n4793) );
  NAND2_X1 U3612 ( .A1(n3584), .A2(U4043), .ZN(n2780) );
  OAI21_X1 U3613 ( .B1(U4043), .B2(n4793), .A(n2780), .ZN(U3556) );
  INV_X1 U3614 ( .A(DATAO_REG_14__SCAN_IN), .ZN(n4754) );
  NAND2_X1 U3615 ( .A1(n4186), .A2(U4043), .ZN(n2781) );
  OAI21_X1 U3616 ( .B1(U4043), .B2(n4754), .A(n2781), .ZN(U3564) );
  INV_X1 U3617 ( .A(DATAO_REG_16__SCAN_IN), .ZN(n4757) );
  NAND2_X1 U3618 ( .A1(n4179), .A2(U4043), .ZN(n2782) );
  OAI21_X1 U3619 ( .B1(U4043), .B2(n4757), .A(n2782), .ZN(U3566) );
  INV_X1 U3620 ( .A(DATAO_REG_5__SCAN_IN), .ZN(n4744) );
  NAND2_X1 U3621 ( .A1(n3059), .A2(U4043), .ZN(n2783) );
  OAI21_X1 U3622 ( .B1(U4043), .B2(n4744), .A(n2783), .ZN(U3555) );
  INV_X1 U3623 ( .A(DATAO_REG_17__SCAN_IN), .ZN(n4756) );
  NAND2_X1 U3624 ( .A1(n3642), .A2(U4043), .ZN(n2784) );
  OAI21_X1 U3625 ( .B1(U4043), .B2(n4756), .A(n2784), .ZN(U3567) );
  INV_X1 U3626 ( .A(DATAO_REG_10__SCAN_IN), .ZN(n4751) );
  NAND2_X1 U3627 ( .A1(n3285), .A2(U4043), .ZN(n2785) );
  OAI21_X1 U3628 ( .B1(U4043), .B2(n4751), .A(n2785), .ZN(U3560) );
  INV_X1 U3629 ( .A(DATAO_REG_15__SCAN_IN), .ZN(n4753) );
  NAND2_X1 U3630 ( .A1(n3415), .A2(U4043), .ZN(n2786) );
  OAI21_X1 U3631 ( .B1(U4043), .B2(n4753), .A(n2786), .ZN(U3565) );
  INV_X1 U3632 ( .A(DATAO_REG_9__SCAN_IN), .ZN(n4794) );
  NAND2_X1 U3633 ( .A1(n3297), .A2(U4043), .ZN(n2787) );
  OAI21_X1 U3634 ( .B1(U4043), .B2(n4794), .A(n2787), .ZN(U3559) );
  INV_X1 U3635 ( .A(DATAO_REG_18__SCAN_IN), .ZN(n4760) );
  NAND2_X1 U3636 ( .A1(n4113), .A2(U4043), .ZN(n2788) );
  OAI21_X1 U3637 ( .B1(U4043), .B2(n4760), .A(n2788), .ZN(U3568) );
  INV_X1 U3638 ( .A(DATAO_REG_21__SCAN_IN), .ZN(n4759) );
  NAND2_X1 U3639 ( .A1(n4082), .A2(U4043), .ZN(n2789) );
  OAI21_X1 U3640 ( .B1(U4043), .B2(n4759), .A(n2789), .ZN(U3571) );
  INV_X1 U3641 ( .A(DATAO_REG_30__SCAN_IN), .ZN(n4769) );
  INV_X1 U3642 ( .A(REG0_REG_30__SCAN_IN), .ZN(n2793) );
  NAND2_X1 U3643 ( .A1(n2411), .A2(REG2_REG_30__SCAN_IN), .ZN(n2792) );
  INV_X1 U3644 ( .A(REG1_REG_30__SCAN_IN), .ZN(n2790) );
  OR2_X1 U3645 ( .A1(n3684), .A2(n2790), .ZN(n2791) );
  OAI211_X1 U3646 ( .C1(n2794), .C2(n2793), .A(n2792), .B(n2791), .ZN(n3940)
         );
  NAND2_X1 U3647 ( .A1(n3940), .A2(U4043), .ZN(n2795) );
  OAI21_X1 U3648 ( .B1(U4043), .B2(n4769), .A(n2795), .ZN(U3580) );
  INV_X1 U3649 ( .A(DATAO_REG_23__SCAN_IN), .ZN(n4789) );
  NAND2_X1 U3650 ( .A1(n4057), .A2(U4043), .ZN(n2796) );
  OAI21_X1 U3651 ( .B1(U4043), .B2(n4789), .A(n2796), .ZN(U3573) );
  INV_X1 U3652 ( .A(DATAO_REG_0__SCAN_IN), .ZN(n4795) );
  NAND2_X1 U3653 ( .A1(n2897), .A2(U4043), .ZN(n2797) );
  OAI21_X1 U3654 ( .B1(U4043), .B2(n4795), .A(n2797), .ZN(U3550) );
  INV_X1 U3655 ( .A(n4364), .ZN(n2813) );
  OR2_X1 U3656 ( .A1(n2799), .A2(n2798), .ZN(n4381) );
  INV_X1 U3657 ( .A(n4368), .ZN(n3853) );
  XNOR2_X1 U3658 ( .A(n2374), .B(IR_REG_27__SCAN_IN), .ZN(n4378) );
  INV_X1 U3659 ( .A(n4378), .ZN(n3852) );
  OR2_X1 U3660 ( .A1(n4368), .A2(n3852), .ZN(n3855) );
  NOR2_X2 U3661 ( .A1(n4381), .A2(n3855), .ZN(n4482) );
  XNOR2_X1 U3662 ( .A(n2804), .B(REG2_REG_1__SCAN_IN), .ZN(n3846) );
  AND2_X1 U3663 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n3857)
         );
  NAND2_X1 U3664 ( .A1(n3846), .A2(n3857), .ZN(n3845) );
  INV_X1 U3665 ( .A(n2804), .ZN(n4366) );
  NAND2_X1 U3666 ( .A1(n4366), .A2(REG2_REG_1__SCAN_IN), .ZN(n2800) );
  INV_X1 U3667 ( .A(REG2_REG_2__SCAN_IN), .ZN(n2801) );
  MUX2_X1 U3668 ( .A(n2801), .B(REG2_REG_2__SCAN_IN), .S(n2134), .Z(n2802) );
  INV_X1 U3669 ( .A(n2134), .ZN(n4365) );
  NAND2_X1 U3670 ( .A1(n4365), .A2(REG2_REG_2__SCAN_IN), .ZN(n2803) );
  INV_X1 U3671 ( .A(REG2_REG_3__SCAN_IN), .ZN(n3075) );
  XNOR2_X1 U3672 ( .A(n2814), .B(n3075), .ZN(n2810) );
  MUX2_X1 U3673 ( .A(n4543), .B(REG1_REG_1__SCAN_IN), .S(n2804), .Z(n3843) );
  AND2_X1 U3674 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n3844)
         );
  NAND2_X1 U3675 ( .A1(n3843), .A2(n3844), .ZN(n3863) );
  NAND2_X1 U3676 ( .A1(n4366), .A2(REG1_REG_1__SCAN_IN), .ZN(n3862) );
  NAND2_X1 U3677 ( .A1(n3863), .A2(n3862), .ZN(n2807) );
  MUX2_X1 U3678 ( .A(n2805), .B(REG1_REG_2__SCAN_IN), .S(n3872), .Z(n2806) );
  NAND2_X1 U3679 ( .A1(n2807), .A2(n2806), .ZN(n3865) );
  NAND2_X1 U3680 ( .A1(n4365), .A2(REG1_REG_2__SCAN_IN), .ZN(n2808) );
  NAND2_X1 U3681 ( .A1(n3865), .A2(n2808), .ZN(n2822) );
  XOR2_X1 U3682 ( .A(REG1_REG_3__SCAN_IN), .B(n2821), .Z(n2809) );
  AOI22_X1 U3683 ( .A1(n4482), .A2(n2810), .B1(n4464), .B2(n2809), .ZN(n2812)
         );
  AOI22_X1 U3684 ( .A1(n4473), .A2(ADDR_REG_3__SCAN_IN), .B1(
        REG3_REG_3__SCAN_IN), .B2(U3149), .ZN(n2811) );
  OAI211_X1 U3685 ( .C1(n2813), .C2(n4485), .A(n2812), .B(n2811), .ZN(U3243)
         );
  INV_X1 U3686 ( .A(REG2_REG_7__SCAN_IN), .ZN(n3132) );
  NAND2_X1 U3687 ( .A1(n2815), .A2(n4364), .ZN(n2816) );
  INV_X1 U3688 ( .A(n3877), .ZN(n4363) );
  AOI22_X1 U3689 ( .A1(n2818), .A2(REG2_REG_4__SCAN_IN), .B1(n4363), .B2(n2817), .ZN(n2866) );
  INV_X1 U3690 ( .A(REG2_REG_5__SCAN_IN), .ZN(n3087) );
  MUX2_X1 U3691 ( .A(n3087), .B(REG2_REG_5__SCAN_IN), .S(n2829), .Z(n2865) );
  NOR2_X1 U3692 ( .A1(n2866), .A2(n2865), .ZN(n2864) );
  INV_X1 U3693 ( .A(n2819), .ZN(n2820) );
  MUX2_X1 U3694 ( .A(REG2_REG_7__SCAN_IN), .B(n3132), .S(n4360), .Z(n2856) );
  OAI21_X1 U3695 ( .B1(n3132), .B2(n4360), .A(n2860), .ZN(n2875) );
  XNOR2_X1 U3696 ( .A(n2875), .B(n2840), .ZN(n2876) );
  XOR2_X1 U3697 ( .A(REG2_REG_8__SCAN_IN), .B(n2876), .Z(n2843) );
  NAND2_X1 U3698 ( .A1(n2821), .A2(REG1_REG_3__SCAN_IN), .ZN(n2824) );
  NAND2_X1 U3699 ( .A1(n2822), .A2(n4364), .ZN(n2823) );
  NAND2_X1 U3700 ( .A1(n2824), .A2(n2823), .ZN(n2825) );
  XNOR2_X1 U3701 ( .A(n2825), .B(n3877), .ZN(n3878) );
  NAND2_X1 U3702 ( .A1(n3878), .A2(REG1_REG_4__SCAN_IN), .ZN(n2827) );
  NAND2_X1 U3703 ( .A1(n2825), .A2(n4363), .ZN(n2826) );
  NAND2_X1 U3704 ( .A1(n2827), .A2(n2826), .ZN(n2868) );
  MUX2_X1 U3705 ( .A(REG1_REG_5__SCAN_IN), .B(n2828), .S(n2829), .Z(n2869) );
  NAND2_X1 U3706 ( .A1(n2868), .A2(n2869), .ZN(n2867) );
  NAND2_X1 U3707 ( .A1(n2829), .A2(REG1_REG_5__SCAN_IN), .ZN(n2830) );
  INV_X1 U3708 ( .A(n4362), .ZN(n2848) );
  NAND2_X1 U3709 ( .A1(n2846), .A2(REG1_REG_6__SCAN_IN), .ZN(n2833) );
  NAND2_X1 U3710 ( .A1(n2831), .A2(n4362), .ZN(n2832) );
  NOR2_X1 U3711 ( .A1(n4360), .A2(n2835), .ZN(n2834) );
  NAND2_X1 U3712 ( .A1(n4360), .A2(n2835), .ZN(n2836) );
  NOR2_X1 U3713 ( .A1(n2837), .A2(n2475), .ZN(n2881) );
  AOI211_X1 U3714 ( .C1(n2475), .C2(n2837), .A(n4468), .B(n2881), .ZN(n2842)
         );
  NAND2_X1 U3715 ( .A1(REG3_REG_8__SCAN_IN), .A2(U3149), .ZN(n3159) );
  INV_X1 U3716 ( .A(n3159), .ZN(n2838) );
  AOI21_X1 U3717 ( .B1(n4473), .B2(ADDR_REG_8__SCAN_IN), .A(n2838), .ZN(n2839)
         );
  OAI21_X1 U3718 ( .B1(n2840), .B2(n4485), .A(n2839), .ZN(n2841) );
  AOI211_X1 U3719 ( .C1(n2843), .C2(n4482), .A(n2842), .B(n2841), .ZN(n2844)
         );
  INV_X1 U3720 ( .A(n2844), .ZN(U3248) );
  XNOR2_X1 U3721 ( .A(n2845), .B(REG2_REG_6__SCAN_IN), .ZN(n2852) );
  XOR2_X1 U3722 ( .A(n2846), .B(REG1_REG_6__SCAN_IN), .Z(n2850) );
  NOR2_X1 U3723 ( .A1(STATE_REG_SCAN_IN), .A2(n4768), .ZN(n3058) );
  AOI21_X1 U3724 ( .B1(n4473), .B2(ADDR_REG_6__SCAN_IN), .A(n3058), .ZN(n2847)
         );
  OAI21_X1 U3725 ( .B1(n2848), .B2(n4485), .A(n2847), .ZN(n2849) );
  AOI21_X1 U3726 ( .B1(n4464), .B2(n2850), .A(n2849), .ZN(n2851) );
  OAI21_X1 U3727 ( .B1(n2852), .B2(n4434), .A(n2851), .ZN(U3246) );
  INV_X1 U3728 ( .A(DATAO_REG_26__SCAN_IN), .ZN(n4766) );
  NAND2_X1 U3729 ( .A1(n3961), .A2(U4043), .ZN(n2853) );
  OAI21_X1 U3730 ( .B1(U4043), .B2(n4766), .A(n2853), .ZN(U3576) );
  XOR2_X1 U3731 ( .A(n2835), .B(n4360), .Z(n2854) );
  XNOR2_X1 U3732 ( .A(n2855), .B(n2854), .ZN(n2863) );
  AOI21_X1 U3733 ( .B1(n2857), .B2(n2856), .A(n4434), .ZN(n2861) );
  INV_X1 U3734 ( .A(REG3_REG_7__SCAN_IN), .ZN(n4581) );
  NOR2_X1 U3735 ( .A1(STATE_REG_SCAN_IN), .A2(n4581), .ZN(n3119) );
  AOI21_X1 U3736 ( .B1(n4473), .B2(ADDR_REG_7__SCAN_IN), .A(n3119), .ZN(n2858)
         );
  OAI21_X1 U3737 ( .B1(n4360), .B2(n4485), .A(n2858), .ZN(n2859) );
  AOI21_X1 U3738 ( .B1(n2861), .B2(n2860), .A(n2859), .ZN(n2862) );
  OAI21_X1 U3739 ( .B1(n4468), .B2(n2863), .A(n2862), .ZN(U3247) );
  AOI211_X1 U3740 ( .C1(n2866), .C2(n2865), .A(n2864), .B(n4434), .ZN(n2874)
         );
  OAI211_X1 U3741 ( .C1(n2869), .C2(n2868), .A(n4464), .B(n2867), .ZN(n2871)
         );
  AND2_X1 U3742 ( .A1(U3149), .A2(REG3_REG_5__SCAN_IN), .ZN(n3587) );
  AOI21_X1 U3743 ( .B1(n4473), .B2(ADDR_REG_5__SCAN_IN), .A(n3587), .ZN(n2870)
         );
  OAI211_X1 U3744 ( .C1(n4485), .C2(n2872), .A(n2871), .B(n2870), .ZN(n2873)
         );
  OR2_X1 U3745 ( .A1(n2874), .A2(n2873), .ZN(U3245) );
  INV_X1 U3746 ( .A(n4359), .ZN(n3903) );
  AOI22_X1 U3747 ( .A1(n2876), .A2(REG2_REG_8__SCAN_IN), .B1(n2882), .B2(n2875), .ZN(n2878) );
  INV_X1 U3748 ( .A(REG2_REG_9__SCAN_IN), .ZN(n3904) );
  MUX2_X1 U3749 ( .A(n3904), .B(REG2_REG_9__SCAN_IN), .S(n4359), .Z(n2877) );
  NOR2_X1 U3750 ( .A1(n2878), .A2(n2877), .ZN(n3902) );
  AOI211_X1 U3751 ( .C1(n2878), .C2(n2877), .A(n4434), .B(n3902), .ZN(n2879)
         );
  INV_X1 U3752 ( .A(n2879), .ZN(n2889) );
  NOR2_X1 U3753 ( .A1(STATE_REG_SCAN_IN), .A2(n4771), .ZN(n3213) );
  INV_X1 U3754 ( .A(n2880), .ZN(n2883) );
  AOI21_X1 U3755 ( .B1(n2883), .B2(n2882), .A(n2881), .ZN(n2886) );
  MUX2_X1 U3756 ( .A(n2884), .B(REG1_REG_9__SCAN_IN), .S(n4359), .Z(n2885) );
  NOR2_X1 U3757 ( .A1(n2886), .A2(n2885), .ZN(n3888) );
  AOI211_X1 U3758 ( .C1(n2886), .C2(n2885), .A(n3888), .B(n4468), .ZN(n2887)
         );
  AOI211_X1 U3759 ( .C1(n4473), .C2(ADDR_REG_9__SCAN_IN), .A(n3213), .B(n2887), 
        .ZN(n2888) );
  OAI211_X1 U3760 ( .C1(n4485), .C2(n3903), .A(n2889), .B(n2888), .ZN(U3249)
         );
  NAND2_X1 U3761 ( .A1(n2890), .A2(n2911), .ZN(n2894) );
  NAND2_X1 U3762 ( .A1(n3074), .A2(n2896), .ZN(n2893) );
  NAND2_X1 U3763 ( .A1(n2894), .A2(n2893), .ZN(n2895) );
  AOI22_X1 U3764 ( .A1(n2890), .A2(n2135), .B1(n2911), .B2(n3074), .ZN(n3010)
         );
  XNOR2_X1 U3765 ( .A(n3009), .B(n3010), .ZN(n3007) );
  NAND2_X1 U3766 ( .A1(n3375), .A2(n2896), .ZN(n2899) );
  NAND2_X1 U3767 ( .A1(n2897), .A2(n2133), .ZN(n2898) );
  NAND2_X1 U3768 ( .A1(n2899), .A2(n2898), .ZN(n2906) );
  INV_X1 U3769 ( .A(n2906), .ZN(n2901) );
  NAND2_X1 U3770 ( .A1(n2901), .A2(n2337), .ZN(n3374) );
  NAND2_X1 U3771 ( .A1(n2897), .A2(n3533), .ZN(n2905) );
  AND2_X1 U3772 ( .A1(n2902), .A2(IR_REG_0__SCAN_IN), .ZN(n2903) );
  NAND2_X1 U3773 ( .A1(n2905), .A2(n2904), .ZN(n3373) );
  NAND2_X1 U3774 ( .A1(n3374), .A2(n3373), .ZN(n3372) );
  OR2_X1 U3775 ( .A1(n2906), .A2(n3530), .ZN(n2907) );
  NAND2_X1 U3776 ( .A1(n3372), .A2(n2907), .ZN(n3547) );
  NAND2_X1 U3777 ( .A1(n3549), .A2(n2896), .ZN(n2908) );
  NAND2_X1 U3778 ( .A1(n2909), .A2(n2908), .ZN(n2910) );
  XNOR2_X1 U3779 ( .A(n2910), .B(n3530), .ZN(n2912) );
  XNOR2_X1 U3780 ( .A(n2912), .B(n2913), .ZN(n3545) );
  NAND2_X1 U3781 ( .A1(n3547), .A2(n3545), .ZN(n3546) );
  INV_X1 U3782 ( .A(n2912), .ZN(n2914) );
  OR2_X1 U3783 ( .A1(n2914), .A2(n2913), .ZN(n2915) );
  NAND2_X1 U3784 ( .A1(n3546), .A2(n2915), .ZN(n3362) );
  INV_X1 U3785 ( .A(n3362), .ZN(n2920) );
  OR2_X1 U3786 ( .A1(n2952), .A2(n3445), .ZN(n2917) );
  NAND2_X1 U3787 ( .A1(n3841), .A2(n2911), .ZN(n2916) );
  XNOR2_X1 U3788 ( .A(n2918), .B(n3487), .ZN(n2921) );
  XNOR2_X1 U3789 ( .A(n2921), .B(n2922), .ZN(n3365) );
  INV_X1 U3790 ( .A(n3365), .ZN(n2919) );
  NAND2_X1 U3791 ( .A1(n2920), .A2(n2919), .ZN(n3363) );
  NAND2_X1 U3792 ( .A1(n2921), .A2(n2922), .ZN(n2923) );
  NAND2_X1 U3793 ( .A1(n3363), .A2(n2923), .ZN(n3008) );
  XOR2_X1 U3794 ( .A(n3007), .B(n3008), .Z(n2949) );
  INV_X1 U3795 ( .A(n2967), .ZN(n2925) );
  NAND3_X1 U3796 ( .A1(n2925), .A2(n2968), .A3(n2924), .ZN(n2941) );
  INV_X1 U3797 ( .A(n2932), .ZN(n2926) );
  NOR2_X1 U3798 ( .A1(n2941), .A2(n2926), .ZN(n2930) );
  AOI21_X1 U3799 ( .B1(n2755), .B2(n2928), .A(n2927), .ZN(n2929) );
  INV_X1 U3800 ( .A(n2930), .ZN(n2934) );
  INV_X1 U3801 ( .A(n3841), .ZN(n3068) );
  INV_X1 U3802 ( .A(n2936), .ZN(n2937) );
  NAND3_X1 U3803 ( .A1(n3532), .A2(n2937), .A3(n4488), .ZN(n3831) );
  INV_X1 U3804 ( .A(n3840), .ZN(n2939) );
  OAI22_X1 U3805 ( .A1(n3068), .A2(n3655), .B1(n3653), .B2(n2939), .ZN(n2947)
         );
  NAND3_X1 U3806 ( .A1(n4275), .A2(n4358), .A3(n2755), .ZN(n2940) );
  NAND2_X1 U3807 ( .A1(n2941), .A2(n2940), .ZN(n3367) );
  AND3_X1 U3808 ( .A1(n2943), .A2(n2891), .A3(n2942), .ZN(n2944) );
  NAND2_X1 U3809 ( .A1(n3367), .A2(n2944), .ZN(n2945) );
  MUX2_X1 U3810 ( .A(n3666), .B(U3149), .S(REG3_REG_3__SCAN_IN), .Z(n2946) );
  AOI211_X1 U3811 ( .C1(n3074), .C2(n2935), .A(n2947), .B(n2946), .ZN(n2948)
         );
  OAI21_X1 U3812 ( .B1(n2949), .B2(n3674), .A(n2948), .ZN(U3215) );
  OAI21_X1 U3813 ( .B1(n2951), .B2(n3722), .A(n2950), .ZN(n3104) );
  INV_X1 U3814 ( .A(n2890), .ZN(n3107) );
  OAI22_X1 U3815 ( .A1(n3107), .A2(n4276), .B1(n2952), .B2(n4275), .ZN(n2958)
         );
  INV_X1 U3816 ( .A(n4554), .ZN(n3335) );
  NAND2_X1 U3817 ( .A1(n3104), .A2(n3335), .ZN(n2957) );
  NAND3_X1 U3818 ( .A1(n2975), .A2(n3722), .A3(n2678), .ZN(n2953) );
  NAND2_X1 U3819 ( .A1(n2954), .A2(n2953), .ZN(n2955) );
  NAND2_X1 U3820 ( .A1(n2955), .A2(n4162), .ZN(n2956) );
  OAI211_X1 U3821 ( .C1(n2385), .C2(n4167), .A(n2957), .B(n2956), .ZN(n3102)
         );
  AOI211_X1 U3822 ( .C1(n4540), .C2(n3104), .A(n2958), .B(n3102), .ZN(n2965)
         );
  NAND2_X1 U3823 ( .A1(n2972), .A2(n3368), .ZN(n2959) );
  AND2_X1 U3824 ( .A1(n3073), .A2(n2959), .ZN(n3103) );
  INV_X1 U3825 ( .A(n3103), .ZN(n2962) );
  OAI22_X1 U3826 ( .A1(n4302), .A2(n2962), .B1(n4551), .B2(n2805), .ZN(n2960)
         );
  INV_X1 U3827 ( .A(n2960), .ZN(n2961) );
  OAI21_X1 U3828 ( .B1(n2965), .B2(n2751), .A(n2961), .ZN(U3520) );
  OAI22_X1 U3829 ( .A1(n4350), .A2(n2962), .B1(n4542), .B2(n2393), .ZN(n2963)
         );
  INV_X1 U3830 ( .A(n2963), .ZN(n2964) );
  OAI21_X1 U3831 ( .B1(n2965), .B2(n4541), .A(n2964), .ZN(U3471) );
  INV_X1 U3832 ( .A(n2966), .ZN(n2970) );
  NOR2_X1 U3833 ( .A1(n2968), .A2(n2967), .ZN(n2969) );
  NAND2_X1 U3834 ( .A1(n2970), .A2(n2969), .ZN(n2971) );
  NAND2_X1 U3835 ( .A1(n4372), .A2(n4555), .ZN(n4137) );
  OAI21_X1 U3836 ( .B1(n4563), .B2(n2978), .A(n2972), .ZN(n4504) );
  OAI21_X1 U3837 ( .B1(n2677), .B2(n2974), .A(n2973), .ZN(n4505) );
  OAI21_X1 U3838 ( .B1(n3747), .B2(n3755), .A(n2975), .ZN(n2980) );
  NAND2_X1 U3839 ( .A1(n2897), .A2(n4187), .ZN(n2977) );
  NAND2_X1 U3840 ( .A1(n3841), .A2(n4289), .ZN(n2976) );
  OAI211_X1 U3841 ( .C1(n4275), .C2(n2978), .A(n2977), .B(n2976), .ZN(n2979)
         );
  AOI21_X1 U3842 ( .B1(n2980), .B2(n4162), .A(n2979), .ZN(n2981) );
  OAI21_X1 U3843 ( .B1(n4554), .B2(n4505), .A(n2981), .ZN(n4507) );
  NAND2_X1 U3844 ( .A1(n4507), .A2(n4372), .ZN(n2988) );
  INV_X1 U3845 ( .A(n4505), .ZN(n2986) );
  OR2_X1 U3846 ( .A1(n2892), .A2(n4555), .ZN(n3028) );
  INV_X1 U3847 ( .A(n3028), .ZN(n2982) );
  INV_X1 U3848 ( .A(REG2_REG_1__SCAN_IN), .ZN(n2984) );
  OAI22_X1 U3849 ( .A1(n4171), .A2(n2984), .B1(n2983), .B2(n4169), .ZN(n2985)
         );
  AOI21_X1 U3850 ( .B1(n2986), .B2(n4100), .A(n2985), .ZN(n2987) );
  OAI211_X1 U3851 ( .C1(n4152), .C2(n4504), .A(n2988), .B(n2987), .ZN(U3289)
         );
  NAND2_X1 U3852 ( .A1(n2989), .A2(n2992), .ZN(n2990) );
  NAND2_X1 U3853 ( .A1(n2991), .A2(n2990), .ZN(n4513) );
  INV_X1 U3854 ( .A(n4100), .ZN(n4565) );
  XNOR2_X1 U3855 ( .A(n2993), .B(n2992), .ZN(n2997) );
  AOI22_X1 U3856 ( .A1(n2890), .A2(n4187), .B1(n3006), .B2(n4288), .ZN(n2995)
         );
  NAND2_X1 U3857 ( .A1(n3059), .A2(n4289), .ZN(n2994) );
  OAI211_X1 U3858 ( .C1(n4513), .C2(n4554), .A(n2995), .B(n2994), .ZN(n2996)
         );
  AOI21_X1 U3859 ( .B1(n2997), .B2(n4162), .A(n2996), .ZN(n2998) );
  INV_X1 U3860 ( .A(n2998), .ZN(n4515) );
  INV_X1 U3861 ( .A(n3086), .ZN(n2999) );
  OAI211_X1 U3862 ( .C1(n3072), .C2(n3020), .A(n2999), .B(n4529), .ZN(n4514)
         );
  OAI22_X1 U3863 ( .A1(n4514), .A2(n4358), .B1(n4169), .B2(n3017), .ZN(n3000)
         );
  OAI21_X1 U3864 ( .B1(n4515), .B2(n3000), .A(n4372), .ZN(n3002) );
  NAND2_X1 U3865 ( .A1(n4142), .A2(REG2_REG_4__SCAN_IN), .ZN(n3001) );
  OAI211_X1 U3866 ( .C1(n4513), .C2(n4565), .A(n3002), .B(n3001), .ZN(U3286)
         );
  NAND2_X1 U3867 ( .A1(n3840), .A2(n2911), .ZN(n3004) );
  OR2_X1 U3868 ( .A1(n3020), .A2(n3445), .ZN(n3003) );
  NAND2_X1 U3869 ( .A1(n3004), .A2(n3003), .ZN(n3005) );
  XNOR2_X1 U3870 ( .A(n3005), .B(n3487), .ZN(n3039) );
  AOI22_X1 U3871 ( .A1(n3840), .A2(n2135), .B1(n3006), .B2(n2911), .ZN(n3038)
         );
  XNOR2_X1 U3872 ( .A(n3039), .B(n3038), .ZN(n3016) );
  INV_X1 U3873 ( .A(n3009), .ZN(n3011) );
  NAND2_X1 U3874 ( .A1(n3011), .A2(n3010), .ZN(n3012) );
  INV_X1 U3875 ( .A(n3041), .ZN(n3015) );
  AOI211_X1 U3876 ( .C1(n3016), .C2(n3013), .A(n3674), .B(n3015), .ZN(n3023)
         );
  INV_X1 U3877 ( .A(n3059), .ZN(n3018) );
  OAI22_X1 U3878 ( .A1(n3653), .A2(n3018), .B1(n3654), .B2(n3017), .ZN(n3022)
         );
  NAND2_X1 U3879 ( .A1(REG3_REG_4__SCAN_IN), .A2(U3149), .ZN(n3876) );
  NAND2_X1 U3880 ( .A1(n3667), .A2(n2890), .ZN(n3019) );
  OAI211_X1 U3881 ( .C1(n3668), .C2(n3020), .A(n3876), .B(n3019), .ZN(n3021)
         );
  OR3_X1 U3882 ( .A1(n3023), .A2(n3022), .A3(n3021), .ZN(U3227) );
  INV_X1 U3883 ( .A(n3024), .ZN(n3777) );
  NAND2_X1 U3884 ( .A1(n3777), .A2(n3767), .ZN(n3711) );
  XNOR2_X1 U3885 ( .A(n3025), .B(n3711), .ZN(n3026) );
  AOI22_X1 U3886 ( .A1(n3026), .A2(n4162), .B1(n4187), .B2(n3059), .ZN(n3094)
         );
  XNOR2_X1 U3887 ( .A(n3027), .B(n3711), .ZN(n3095) );
  INV_X1 U3888 ( .A(n3095), .ZN(n3036) );
  NAND2_X1 U3889 ( .A1(n4554), .A2(n3028), .ZN(n3029) );
  NAND2_X1 U3890 ( .A1(n3085), .A2(n3092), .ZN(n3030) );
  NAND2_X1 U3891 ( .A1(n3128), .A2(n3030), .ZN(n3098) );
  INV_X1 U3892 ( .A(n3839), .ZN(n3165) );
  NAND2_X1 U3893 ( .A1(n4372), .A2(n4289), .ZN(n4559) );
  INV_X1 U3894 ( .A(n3031), .ZN(n3055) );
  AOI22_X1 U3895 ( .A1(n4142), .A2(REG2_REG_6__SCAN_IN), .B1(n3055), .B2(n4568), .ZN(n3032) );
  OAI21_X1 U3896 ( .B1(n3165), .B2(n4559), .A(n3032), .ZN(n3033) );
  AOI21_X1 U3897 ( .B1(n3092), .B2(n4552), .A(n3033), .ZN(n3034) );
  OAI21_X1 U3898 ( .B1(n3098), .B2(n4152), .A(n3034), .ZN(n3035) );
  AOI21_X1 U3899 ( .B1(n3036), .B2(n4139), .A(n3035), .ZN(n3037) );
  OAI21_X1 U3900 ( .B1(n3094), .B2(n4142), .A(n3037), .ZN(U3284) );
  OR2_X1 U3901 ( .A1(n3039), .A2(n3038), .ZN(n3040) );
  NAND2_X1 U3902 ( .A1(n3041), .A2(n3040), .ZN(n3581) );
  NAND2_X1 U3903 ( .A1(n3059), .A2(n2133), .ZN(n3043) );
  NAND2_X1 U3904 ( .A1(n3080), .A2(n2896), .ZN(n3042) );
  NAND2_X1 U3905 ( .A1(n3043), .A2(n3042), .ZN(n3044) );
  XNOR2_X1 U3906 ( .A(n3044), .B(n3530), .ZN(n3045) );
  AOI22_X1 U3907 ( .A1(n3059), .A2(n2135), .B1(n2133), .B2(n3080), .ZN(n3046)
         );
  XNOR2_X1 U3908 ( .A(n3045), .B(n3046), .ZN(n3580) );
  INV_X1 U3909 ( .A(n3045), .ZN(n3047) );
  OR2_X1 U3910 ( .A1(n3047), .A2(n3046), .ZN(n3048) );
  NAND2_X1 U3911 ( .A1(n3584), .A2(n2135), .ZN(n3050) );
  NAND2_X1 U3912 ( .A1(n3092), .A2(n2911), .ZN(n3049) );
  NAND2_X1 U3913 ( .A1(n3050), .A2(n3049), .ZN(n3111) );
  NAND2_X1 U3914 ( .A1(n3584), .A2(n2911), .ZN(n3052) );
  NAND2_X1 U3915 ( .A1(n3092), .A2(n2896), .ZN(n3051) );
  NAND2_X1 U3916 ( .A1(n3052), .A2(n3051), .ZN(n3053) );
  XNOR2_X1 U3917 ( .A(n3053), .B(n3530), .ZN(n3110) );
  XOR2_X1 U3918 ( .A(n3111), .B(n3110), .Z(n3054) );
  XNOR2_X1 U3919 ( .A(n3112), .B(n3054), .ZN(n3062) );
  AOI22_X1 U3920 ( .A1(n3671), .A2(n3839), .B1(n3666), .B2(n3055), .ZN(n3061)
         );
  NOR2_X1 U3921 ( .A1(n3668), .A2(n3056), .ZN(n3057) );
  AOI211_X1 U3922 ( .C1(n3667), .C2(n3059), .A(n3058), .B(n3057), .ZN(n3060)
         );
  OAI211_X1 U3923 ( .C1(n3062), .C2(n3674), .A(n3061), .B(n3060), .ZN(U3236)
         );
  XNOR2_X1 U3924 ( .A(n3063), .B(n3066), .ZN(n4509) );
  OAI21_X1 U3925 ( .B1(n3066), .B2(n3065), .A(n3064), .ZN(n3070) );
  AOI22_X1 U3926 ( .A1(n3840), .A2(n4289), .B1(n4288), .B2(n3074), .ZN(n3067)
         );
  OAI21_X1 U3927 ( .B1(n3068), .B2(n4167), .A(n3067), .ZN(n3069) );
  AOI21_X1 U3928 ( .B1(n3070), .B2(n4162), .A(n3069), .ZN(n3071) );
  OAI21_X1 U3929 ( .B1(n4509), .B2(n4554), .A(n3071), .ZN(n4510) );
  NAND2_X1 U3930 ( .A1(n4510), .A2(n4372), .ZN(n3078) );
  AOI21_X1 U3931 ( .B1(n3074), .B2(n3073), .A(n3072), .ZN(n4512) );
  OAI22_X1 U3932 ( .A1(n4372), .A2(n3075), .B1(REG3_REG_3__SCAN_IN), .B2(n4169), .ZN(n3076) );
  AOI21_X1 U3933 ( .B1(n4512), .B2(n4373), .A(n3076), .ZN(n3077) );
  OAI211_X1 U3934 ( .C1(n4509), .C2(n4565), .A(n3078), .B(n3077), .ZN(U3287)
         );
  NAND2_X1 U3935 ( .A1(n3774), .A2(n3764), .ZN(n3717) );
  XOR2_X1 U3936 ( .A(n3717), .B(n3079), .Z(n3083) );
  AOI22_X1 U3937 ( .A1(n3584), .A2(n4289), .B1(n4288), .B2(n3080), .ZN(n3082)
         );
  NAND2_X1 U3938 ( .A1(n3840), .A2(n4187), .ZN(n3081) );
  OAI211_X1 U3939 ( .C1(n3083), .C2(n4553), .A(n3082), .B(n3081), .ZN(n4519)
         );
  INV_X1 U3940 ( .A(n4519), .ZN(n3091) );
  XOR2_X1 U3941 ( .A(n3084), .B(n3717), .Z(n4521) );
  OAI21_X1 U3942 ( .B1(n3086), .B2(n3585), .A(n3085), .ZN(n4518) );
  NOR2_X1 U3943 ( .A1(n4518), .A2(n4152), .ZN(n3089) );
  OAI22_X1 U3944 ( .A1(n4372), .A2(n3087), .B1(n3582), .B2(n4169), .ZN(n3088)
         );
  AOI211_X1 U3945 ( .C1(n4521), .C2(n4139), .A(n3089), .B(n3088), .ZN(n3090)
         );
  OAI21_X1 U3946 ( .B1(n3091), .B2(n4142), .A(n3090), .ZN(U3285) );
  AOI22_X1 U3947 ( .A1(n3839), .A2(n4289), .B1(n3092), .B2(n4288), .ZN(n3093)
         );
  OAI211_X1 U3948 ( .C1(n4522), .C2(n3095), .A(n3094), .B(n3093), .ZN(n3100)
         );
  OAI22_X1 U3949 ( .A1(n3098), .A2(n4302), .B1(n4551), .B2(n2448), .ZN(n3096)
         );
  AOI21_X1 U3950 ( .B1(n3100), .B2(n4551), .A(n3096), .ZN(n3097) );
  INV_X1 U3951 ( .A(n3097), .ZN(U3524) );
  OAI22_X1 U3952 ( .A1(n3098), .A2(n4350), .B1(n4542), .B2(n2447), .ZN(n3099)
         );
  AOI21_X1 U3953 ( .B1(n3100), .B2(n4542), .A(n3099), .ZN(n3101) );
  INV_X1 U3954 ( .A(n3101), .ZN(U3479) );
  MUX2_X1 U3955 ( .A(n3102), .B(REG2_REG_2__SCAN_IN), .S(n4142), .Z(n3109) );
  AOI22_X1 U3956 ( .A1(n3104), .A2(n4100), .B1(n4373), .B2(n3103), .ZN(n3106)
         );
  AOI22_X1 U3957 ( .A1(n4552), .A2(n3368), .B1(REG3_REG_2__SCAN_IN), .B2(n4568), .ZN(n3105) );
  OAI211_X1 U3958 ( .C1(n3107), .C2(n4559), .A(n3106), .B(n3105), .ZN(n3108)
         );
  OR2_X1 U3959 ( .A1(n3109), .A2(n3108), .ZN(U3288) );
  NAND2_X1 U3960 ( .A1(n3839), .A2(n2133), .ZN(n3114) );
  OR2_X1 U3961 ( .A1(n3117), .A2(n3445), .ZN(n3113) );
  NAND2_X1 U3962 ( .A1(n3114), .A2(n3113), .ZN(n3115) );
  XNOR2_X1 U3963 ( .A(n3115), .B(n3530), .ZN(n3143) );
  AOI22_X1 U3964 ( .A1(n3839), .A2(n2135), .B1(n3127), .B2(n2133), .ZN(n3144)
         );
  XNOR2_X1 U3965 ( .A(n3142), .B(n3141), .ZN(n3122) );
  INV_X1 U3966 ( .A(n3131), .ZN(n3116) );
  AOI22_X1 U3967 ( .A1(n3671), .A2(n3838), .B1(n3666), .B2(n3116), .ZN(n3121)
         );
  NOR2_X1 U3968 ( .A1(n3668), .A2(n3117), .ZN(n3118) );
  AOI211_X1 U3969 ( .C1(n3667), .C2(n3584), .A(n3119), .B(n3118), .ZN(n3120)
         );
  OAI211_X1 U3970 ( .C1(n3122), .C2(n3674), .A(n3121), .B(n3120), .ZN(U3210)
         );
  XOR2_X1 U3971 ( .A(n3768), .B(n3123), .Z(n3126) );
  AOI22_X1 U3972 ( .A1(n3838), .A2(n4289), .B1(n3127), .B2(n4288), .ZN(n3125)
         );
  NAND2_X1 U3973 ( .A1(n3584), .A2(n4187), .ZN(n3124) );
  OAI211_X1 U3974 ( .C1(n3126), .C2(n4553), .A(n3125), .B(n3124), .ZN(n4524)
         );
  INV_X1 U3975 ( .A(n4524), .ZN(n3140) );
  INV_X1 U3976 ( .A(n4137), .ZN(n3138) );
  NAND2_X1 U3977 ( .A1(n3128), .A2(n3127), .ZN(n3129) );
  NAND2_X1 U3978 ( .A1(n3129), .A2(n4529), .ZN(n3130) );
  NOR2_X1 U3979 ( .A1(n3167), .A2(n3130), .ZN(n4525) );
  OAI22_X1 U3980 ( .A1(n4171), .A2(n3132), .B1(n3131), .B2(n4169), .ZN(n3137)
         );
  INV_X1 U3981 ( .A(n3133), .ZN(n3135) );
  AND2_X1 U3982 ( .A1(n3134), .A2(n3768), .ZN(n4523) );
  NOR3_X1 U3983 ( .A1(n3135), .A2(n4523), .A3(n4193), .ZN(n3136) );
  AOI211_X1 U3984 ( .C1(n3138), .C2(n4525), .A(n3137), .B(n3136), .ZN(n3139)
         );
  OAI21_X1 U3985 ( .B1(n4142), .B2(n3140), .A(n3139), .ZN(U3283) );
  NAND2_X1 U3986 ( .A1(n3142), .A2(n3141), .ZN(n3147) );
  INV_X1 U3987 ( .A(n3143), .ZN(n3145) );
  OR2_X1 U3988 ( .A1(n3145), .A2(n3144), .ZN(n3146) );
  NAND2_X1 U3989 ( .A1(n3838), .A2(n2911), .ZN(n3149) );
  NAND2_X1 U3990 ( .A1(n3171), .A2(n2896), .ZN(n3148) );
  NAND2_X1 U3991 ( .A1(n3149), .A2(n3148), .ZN(n3150) );
  XNOR2_X1 U3992 ( .A(n3150), .B(n3530), .ZN(n3156) );
  INV_X1 U3993 ( .A(n3156), .ZN(n3154) );
  NAND2_X1 U3994 ( .A1(n3838), .A2(n2135), .ZN(n3152) );
  NAND2_X1 U3995 ( .A1(n3171), .A2(n2133), .ZN(n3151) );
  NAND2_X1 U3996 ( .A1(n3152), .A2(n3151), .ZN(n3155) );
  INV_X1 U3997 ( .A(n3155), .ZN(n3153) );
  NAND2_X1 U3998 ( .A1(n3154), .A2(n3153), .ZN(n3204) );
  INV_X1 U3999 ( .A(n3204), .ZN(n3157) );
  AND2_X1 U4000 ( .A1(n3156), .A2(n3155), .ZN(n3202) );
  NOR2_X1 U4001 ( .A1(n3157), .A2(n3202), .ZN(n3158) );
  XNOR2_X1 U4002 ( .A(n3203), .B(n3158), .ZN(n3163) );
  OAI21_X1 U4003 ( .B1(n3655), .B2(n3165), .A(n3159), .ZN(n3161) );
  INV_X1 U4004 ( .A(n3297), .ZN(n3193) );
  OAI22_X1 U4005 ( .A1(n3653), .A2(n3193), .B1(n3654), .B2(n3169), .ZN(n3160)
         );
  AOI211_X1 U4006 ( .C1(n3171), .C2(n2935), .A(n3161), .B(n3160), .ZN(n3162)
         );
  OAI21_X1 U4007 ( .B1(n3163), .B2(n3674), .A(n3162), .ZN(U3218) );
  NAND2_X1 U4008 ( .A1(n3771), .A2(n3775), .ZN(n3710) );
  XOR2_X1 U4009 ( .A(n3710), .B(n3164), .Z(n3166) );
  OAI22_X1 U4010 ( .A1(n3166), .A2(n4553), .B1(n3165), .B2(n4167), .ZN(n3194)
         );
  INV_X1 U4011 ( .A(n3194), .ZN(n3179) );
  INV_X1 U4012 ( .A(n3167), .ZN(n3168) );
  AOI21_X1 U4013 ( .B1(n3171), .B2(n3168), .A(n3185), .ZN(n3199) );
  INV_X1 U4014 ( .A(n3169), .ZN(n3170) );
  AOI22_X1 U4015 ( .A1(n4142), .A2(REG2_REG_8__SCAN_IN), .B1(n3170), .B2(n4568), .ZN(n3173) );
  NAND2_X1 U4016 ( .A1(n4552), .A2(n3171), .ZN(n3172) );
  OAI211_X1 U4017 ( .C1(n3193), .C2(n4559), .A(n3173), .B(n3172), .ZN(n3174)
         );
  AOI21_X1 U4018 ( .B1(n3199), .B2(n4373), .A(n3174), .ZN(n3178) );
  INV_X1 U4019 ( .A(n3710), .ZN(n3175) );
  XNOR2_X1 U4020 ( .A(n3176), .B(n3175), .ZN(n3196) );
  NAND2_X1 U4021 ( .A1(n3196), .A2(n4139), .ZN(n3177) );
  OAI211_X1 U4022 ( .C1(n3179), .C2(n4142), .A(n3178), .B(n3177), .ZN(U3282)
         );
  NAND2_X1 U4023 ( .A1(n2168), .A2(n3772), .ZN(n3716) );
  XNOR2_X1 U4024 ( .A(n3180), .B(n3716), .ZN(n3184) );
  NAND2_X1 U4025 ( .A1(n3838), .A2(n4187), .ZN(n3182) );
  NAND2_X1 U4026 ( .A1(n3285), .A2(n4289), .ZN(n3181) );
  OAI211_X1 U4027 ( .C1(n4275), .C2(n3211), .A(n3182), .B(n3181), .ZN(n3183)
         );
  AOI21_X1 U4028 ( .B1(n3184), .B2(n4162), .A(n3183), .ZN(n4533) );
  OR2_X1 U4029 ( .A1(n3185), .A2(n3211), .ZN(n3186) );
  AND2_X1 U4030 ( .A1(n3223), .A2(n3186), .ZN(n4530) );
  OAI22_X1 U4031 ( .A1(n4171), .A2(n3904), .B1(n3209), .B2(n4169), .ZN(n3187)
         );
  AOI21_X1 U4032 ( .B1(n4530), .B2(n4373), .A(n3187), .ZN(n3191) );
  INV_X1 U4033 ( .A(n3716), .ZN(n3188) );
  XNOR2_X1 U4034 ( .A(n3189), .B(n3188), .ZN(n4528) );
  NAND2_X1 U4035 ( .A1(n4528), .A2(n4139), .ZN(n3190) );
  OAI211_X1 U4036 ( .C1(n4533), .C2(n4142), .A(n3191), .B(n3190), .ZN(U3281)
         );
  OAI22_X1 U4037 ( .A1(n3193), .A2(n4276), .B1(n3192), .B2(n4275), .ZN(n3195)
         );
  AOI211_X1 U4038 ( .C1(n3196), .C2(n4527), .A(n3195), .B(n3194), .ZN(n3201)
         );
  INV_X1 U4039 ( .A(n4350), .ZN(n4345) );
  NOR2_X1 U4040 ( .A1(n4542), .A2(n2474), .ZN(n3197) );
  AOI21_X1 U4041 ( .B1(n3199), .B2(n4345), .A(n3197), .ZN(n3198) );
  OAI21_X1 U4042 ( .B1(n3201), .B2(n4541), .A(n3198), .ZN(U3483) );
  INV_X1 U40430 ( .A(n4302), .ZN(n4295) );
  AOI22_X1 U4044 ( .A1(n3199), .A2(n4295), .B1(n2751), .B2(REG1_REG_8__SCAN_IN), .ZN(n3200) );
  OAI21_X1 U4045 ( .B1(n3201), .B2(n2751), .A(n3200), .ZN(U3526) );
  NAND2_X1 U4046 ( .A1(n3297), .A2(n2133), .ZN(n3206) );
  NAND2_X1 U4047 ( .A1(n3208), .A2(n2896), .ZN(n3205) );
  NAND2_X1 U4048 ( .A1(n3206), .A2(n3205), .ZN(n3207) );
  XNOR2_X1 U4049 ( .A(n3207), .B(n3530), .ZN(n3262) );
  AOI22_X1 U4050 ( .A1(n3297), .A2(n2135), .B1(n2911), .B2(n3208), .ZN(n3263)
         );
  XNOR2_X1 U4051 ( .A(n3262), .B(n3263), .ZN(n3260) );
  XOR2_X1 U4052 ( .A(n3261), .B(n3260), .Z(n3216) );
  INV_X1 U4053 ( .A(n3209), .ZN(n3210) );
  AOI22_X1 U4054 ( .A1(n3671), .A2(n3285), .B1(n3666), .B2(n3210), .ZN(n3215)
         );
  NOR2_X1 U4055 ( .A1(n3668), .A2(n3211), .ZN(n3212) );
  AOI211_X1 U4056 ( .C1(n3667), .C2(n3838), .A(n3213), .B(n3212), .ZN(n3214)
         );
  OAI211_X1 U4057 ( .C1(n3216), .C2(n3674), .A(n3215), .B(n3214), .ZN(U3228)
         );
  NAND2_X1 U4058 ( .A1(n3781), .A2(n3785), .ZN(n3714) );
  XNOR2_X1 U4059 ( .A(n3217), .B(n3714), .ZN(n3222) );
  XNOR2_X1 U4060 ( .A(n3218), .B(n3714), .ZN(n4539) );
  NAND2_X1 U4061 ( .A1(n4539), .A2(n3335), .ZN(n3221) );
  INV_X1 U4062 ( .A(n3279), .ZN(n3317) );
  OAI22_X1 U4063 ( .A1(n3317), .A2(n4276), .B1(n4275), .B2(n3299), .ZN(n3219)
         );
  AOI21_X1 U4064 ( .B1(n4187), .B2(n3297), .A(n3219), .ZN(n3220) );
  OAI211_X1 U4065 ( .C1(n4553), .C2(n3222), .A(n3221), .B(n3220), .ZN(n4537)
         );
  INV_X1 U4066 ( .A(n4537), .ZN(n3229) );
  INV_X1 U4067 ( .A(n3223), .ZN(n3224) );
  NOR2_X1 U4068 ( .A1(n3224), .A2(n3299), .ZN(n4536) );
  INV_X1 U4069 ( .A(n3253), .ZN(n4535) );
  NOR3_X1 U4070 ( .A1(n4536), .A2(n4535), .A3(n4152), .ZN(n3227) );
  INV_X1 U4071 ( .A(REG2_REG_10__SCAN_IN), .ZN(n3225) );
  OAI22_X1 U4072 ( .A1(n4171), .A2(n3225), .B1(n3296), .B2(n4169), .ZN(n3226)
         );
  AOI211_X1 U4073 ( .C1(n4539), .C2(n4100), .A(n3227), .B(n3226), .ZN(n3228)
         );
  OAI21_X1 U4074 ( .B1(n3229), .B2(n4142), .A(n3228), .ZN(U3280) );
  INV_X1 U4075 ( .A(n3327), .ZN(n3230) );
  OR2_X1 U4076 ( .A1(n3328), .A2(n3230), .ZN(n3715) );
  INV_X1 U4077 ( .A(n3715), .ZN(n3231) );
  XNOR2_X1 U4078 ( .A(n3329), .B(n3231), .ZN(n3233) );
  AND2_X1 U4079 ( .A1(n3279), .A2(n4187), .ZN(n3232) );
  AOI21_X1 U4080 ( .B1(n3233), .B2(n4162), .A(n3232), .ZN(n4292) );
  XNOR2_X1 U4081 ( .A(n3234), .B(n3715), .ZN(n4286) );
  INV_X1 U4082 ( .A(n4290), .ZN(n3496) );
  AOI21_X1 U4083 ( .B1(n4287), .B2(n3255), .A(n3336), .ZN(n4346) );
  NAND2_X1 U4084 ( .A1(n4346), .A2(n4373), .ZN(n3238) );
  INV_X1 U4085 ( .A(REG2_REG_12__SCAN_IN), .ZN(n3235) );
  OAI22_X1 U4086 ( .A1(n4171), .A2(n3235), .B1(n3318), .B2(n4169), .ZN(n3236)
         );
  AOI21_X1 U4087 ( .B1(n4287), .B2(n4552), .A(n3236), .ZN(n3237) );
  OAI211_X1 U4088 ( .C1(n3496), .C2(n4559), .A(n3238), .B(n3237), .ZN(n3239)
         );
  AOI21_X1 U4089 ( .B1(n4286), .B2(n4139), .A(n3239), .ZN(n3240) );
  OAI21_X1 U4090 ( .B1(n4292), .B2(n4142), .A(n3240), .ZN(U3278) );
  XNOR2_X1 U4091 ( .A(n3242), .B(n3241), .ZN(n3251) );
  OAI22_X1 U4092 ( .A1(n3218), .A2(n3243), .B1(n3249), .B2(n3299), .ZN(n3244)
         );
  INV_X1 U4093 ( .A(n3244), .ZN(n3246) );
  OAI21_X1 U4094 ( .B1(n3246), .B2(n3718), .A(n3245), .ZN(n4299) );
  NAND2_X1 U4095 ( .A1(n4299), .A2(n3335), .ZN(n3248) );
  AOI22_X1 U4096 ( .A1(n3837), .A2(n4289), .B1(n3252), .B2(n4288), .ZN(n3247)
         );
  OAI211_X1 U4097 ( .C1(n3249), .C2(n4167), .A(n3248), .B(n3247), .ZN(n3250)
         );
  AOI21_X1 U4098 ( .B1(n3251), .B2(n4162), .A(n3250), .ZN(n4297) );
  NAND2_X1 U4099 ( .A1(n3253), .A2(n3252), .ZN(n3254) );
  NAND2_X1 U4100 ( .A1(n3255), .A2(n3254), .ZN(n4351) );
  INV_X1 U4101 ( .A(n3256), .ZN(n3284) );
  AOI22_X1 U4102 ( .A1(n4142), .A2(REG2_REG_11__SCAN_IN), .B1(n3284), .B2(
        n4568), .ZN(n3257) );
  OAI21_X1 U4103 ( .B1(n4351), .B2(n4152), .A(n3257), .ZN(n3258) );
  AOI21_X1 U4104 ( .B1(n4299), .B2(n4100), .A(n3258), .ZN(n3259) );
  OAI21_X1 U4105 ( .B1(n4297), .B2(n4142), .A(n3259), .ZN(U3279) );
  INV_X1 U4106 ( .A(n3262), .ZN(n3264) );
  NAND2_X1 U4107 ( .A1(n3264), .A2(n3263), .ZN(n3265) );
  NAND2_X1 U4108 ( .A1(n3266), .A2(n3265), .ZN(n3292) );
  INV_X1 U4109 ( .A(n3292), .ZN(n3272) );
  NAND2_X1 U4110 ( .A1(n3285), .A2(n3532), .ZN(n3268) );
  NAND2_X1 U4111 ( .A1(n3270), .A2(n2896), .ZN(n3267) );
  NAND2_X1 U4112 ( .A1(n3268), .A2(n3267), .ZN(n3269) );
  XNOR2_X1 U4113 ( .A(n3269), .B(n3487), .ZN(n3274) );
  AOI22_X1 U4114 ( .A1(n3285), .A2(n2135), .B1(n3532), .B2(n3270), .ZN(n3273)
         );
  XNOR2_X1 U4115 ( .A(n3274), .B(n3273), .ZN(n3295) );
  NAND2_X1 U4116 ( .A1(n3272), .A2(n3271), .ZN(n3293) );
  OR2_X1 U4117 ( .A1(n3274), .A2(n3273), .ZN(n3275) );
  NAND2_X1 U4118 ( .A1(n3279), .A2(n2135), .ZN(n3278) );
  OR2_X1 U4119 ( .A1(n3287), .A2(n3276), .ZN(n3277) );
  NAND2_X1 U4120 ( .A1(n3278), .A2(n3277), .ZN(n3304) );
  NAND2_X1 U4121 ( .A1(n3279), .A2(n3532), .ZN(n3281) );
  OR2_X1 U4122 ( .A1(n3287), .A2(n3445), .ZN(n3280) );
  NAND2_X1 U4123 ( .A1(n3281), .A2(n3280), .ZN(n3282) );
  XNOR2_X1 U4124 ( .A(n3282), .B(n3530), .ZN(n3303) );
  XOR2_X1 U4125 ( .A(n3304), .B(n3303), .Z(n3283) );
  XNOR2_X1 U4126 ( .A(n3305), .B(n3283), .ZN(n3291) );
  AOI22_X1 U4127 ( .A1(n3667), .A2(n3285), .B1(n3666), .B2(n3284), .ZN(n3290)
         );
  INV_X1 U4128 ( .A(REG3_REG_11__SCAN_IN), .ZN(n3286) );
  NOR2_X1 U4129 ( .A1(STATE_REG_SCAN_IN), .A2(n3286), .ZN(n4395) );
  NOR2_X1 U4130 ( .A1(n3668), .A2(n3287), .ZN(n3288) );
  AOI211_X1 U4131 ( .C1(n3671), .C2(n3837), .A(n4395), .B(n3288), .ZN(n3289)
         );
  OAI211_X1 U4132 ( .C1(n3291), .C2(n3674), .A(n3290), .B(n3289), .ZN(U3233)
         );
  INV_X1 U4133 ( .A(n3293), .ZN(n3294) );
  AOI211_X1 U4134 ( .C1(n3295), .C2(n3292), .A(n3674), .B(n3294), .ZN(n3302)
         );
  OAI22_X1 U4135 ( .A1(n3653), .A2(n3317), .B1(n3654), .B2(n3296), .ZN(n3301)
         );
  NAND2_X1 U4136 ( .A1(REG3_REG_10__SCAN_IN), .A2(U3149), .ZN(n4385) );
  NAND2_X1 U4137 ( .A1(n3667), .A2(n3297), .ZN(n3298) );
  OAI211_X1 U4138 ( .C1(n3668), .C2(n3299), .A(n4385), .B(n3298), .ZN(n3300)
         );
  OR3_X1 U4139 ( .A1(n3302), .A2(n3301), .A3(n3300), .ZN(U3214) );
  NAND2_X1 U4140 ( .A1(n3837), .A2(n3532), .ZN(n3307) );
  NAND2_X1 U4141 ( .A1(n4287), .A2(n2896), .ZN(n3306) );
  NAND2_X1 U4142 ( .A1(n3307), .A2(n3306), .ZN(n3308) );
  XNOR2_X1 U4143 ( .A(n3308), .B(n3530), .ZN(n3314) );
  INV_X1 U4144 ( .A(n3314), .ZN(n3312) );
  NAND2_X1 U4145 ( .A1(n3837), .A2(n2135), .ZN(n3310) );
  NAND2_X1 U4146 ( .A1(n4287), .A2(n3532), .ZN(n3309) );
  NAND2_X1 U4147 ( .A1(n3310), .A2(n3309), .ZN(n3313) );
  INV_X1 U4148 ( .A(n3313), .ZN(n3311) );
  NAND2_X1 U4149 ( .A1(n3312), .A2(n3311), .ZN(n3391) );
  INV_X1 U4150 ( .A(n3391), .ZN(n3315) );
  AND2_X1 U4151 ( .A1(n3314), .A2(n3313), .ZN(n3389) );
  NOR2_X1 U4152 ( .A1(n3315), .A2(n3389), .ZN(n3316) );
  XNOR2_X1 U4153 ( .A(n3388), .B(n3316), .ZN(n3322) );
  NAND2_X1 U4154 ( .A1(REG3_REG_12__SCAN_IN), .A2(U3149), .ZN(n4404) );
  OAI21_X1 U4155 ( .B1(n3655), .B2(n3317), .A(n4404), .ZN(n3320) );
  OAI22_X1 U4156 ( .A1(n3653), .A2(n3496), .B1(n3654), .B2(n3318), .ZN(n3319)
         );
  AOI211_X1 U4157 ( .C1(n4287), .C2(n2935), .A(n3320), .B(n3319), .ZN(n3321)
         );
  OAI21_X1 U4158 ( .B1(n3322), .B2(n3674), .A(n3321), .ZN(U3221) );
  INV_X1 U4159 ( .A(n3324), .ZN(n3325) );
  OR2_X1 U4160 ( .A1(n3326), .A2(n3325), .ZN(n3733) );
  XNOR2_X1 U4161 ( .A(n3323), .B(n3733), .ZN(n4282) );
  OAI21_X1 U4162 ( .B1(n3329), .B2(n3328), .A(n3327), .ZN(n3330) );
  XOR2_X1 U4163 ( .A(n3733), .B(n3330), .Z(n3333) );
  AOI22_X1 U4164 ( .A1(n4186), .A2(n4289), .B1(n4288), .B2(n3396), .ZN(n3332)
         );
  NAND2_X1 U4165 ( .A1(n3837), .A2(n4187), .ZN(n3331) );
  OAI211_X1 U4166 ( .C1(n3333), .C2(n4553), .A(n3332), .B(n3331), .ZN(n3334)
         );
  AOI21_X1 U4167 ( .B1(n3335), .B2(n4282), .A(n3334), .ZN(n4284) );
  OR2_X1 U4168 ( .A1(n3336), .A2(n3624), .ZN(n3337) );
  NAND2_X1 U4169 ( .A1(n3345), .A2(n3337), .ZN(n4285) );
  INV_X1 U4170 ( .A(n3338), .ZN(n3623) );
  AOI22_X1 U4171 ( .A1(n4142), .A2(REG2_REG_13__SCAN_IN), .B1(n3623), .B2(
        n4568), .ZN(n3339) );
  OAI21_X1 U4172 ( .B1(n4285), .B2(n4152), .A(n3339), .ZN(n3340) );
  AOI21_X1 U4173 ( .B1(n4282), .B2(n4100), .A(n3340), .ZN(n3341) );
  OAI21_X1 U4174 ( .B1(n4284), .B2(n4142), .A(n3341), .ZN(U3277) );
  XNOR2_X1 U4175 ( .A(n3691), .B(n3719), .ZN(n3342) );
  OAI22_X1 U4176 ( .A1(n3342), .A2(n4553), .B1(n3496), .B2(n4167), .ZN(n4278)
         );
  INV_X1 U4177 ( .A(n4278), .ZN(n3353) );
  OAI21_X1 U4178 ( .B1(n3344), .B2(n3719), .A(n3343), .ZN(n4280) );
  INV_X1 U4179 ( .A(n3345), .ZN(n3346) );
  OAI21_X1 U4180 ( .B1(n3346), .B2(n4274), .A(n4178), .ZN(n4341) );
  INV_X1 U4181 ( .A(REG2_REG_14__SCAN_IN), .ZN(n3347) );
  OAI22_X1 U4182 ( .A1(n4171), .A2(n3347), .B1(n3497), .B2(n4169), .ZN(n3349)
         );
  INV_X1 U4183 ( .A(n3415), .ZN(n4277) );
  NOR2_X1 U4184 ( .A1(n4559), .A2(n4277), .ZN(n3348) );
  AOI211_X1 U4185 ( .C1(n4552), .C2(n3500), .A(n3349), .B(n3348), .ZN(n3350)
         );
  OAI21_X1 U4186 ( .B1(n4341), .B2(n4152), .A(n3350), .ZN(n3351) );
  AOI21_X1 U4187 ( .B1(n4280), .B2(n4139), .A(n3351), .ZN(n3352) );
  OAI21_X1 U4188 ( .B1(n4142), .B2(n3353), .A(n3352), .ZN(U3276) );
  INV_X1 U4189 ( .A(DATAI_30_), .ZN(n3355) );
  NAND2_X1 U4190 ( .A1(n2367), .A2(STATE_REG_SCAN_IN), .ZN(n3354) );
  OAI21_X1 U4191 ( .B1(STATE_REG_SCAN_IN), .B2(n3355), .A(n3354), .ZN(U3322)
         );
  NOR2_X1 U4192 ( .A1(n4563), .A2(n3356), .ZN(n4556) );
  NAND2_X1 U4193 ( .A1(n2897), .A2(n4563), .ZN(n3753) );
  NAND2_X1 U4194 ( .A1(n3357), .A2(n3753), .ZN(n4558) );
  INV_X1 U4195 ( .A(n4558), .ZN(n4564) );
  AOI21_X1 U4196 ( .B1(n4553), .B2(n4522), .A(n4564), .ZN(n3358) );
  AOI211_X1 U4197 ( .C1(n4289), .C2(n3842), .A(n4556), .B(n3358), .ZN(n3361)
         );
  INV_X1 U4198 ( .A(REG0_REG_0__SCAN_IN), .ZN(n4666) );
  NAND2_X1 U4199 ( .A1(n4541), .A2(REG0_REG_0__SCAN_IN), .ZN(n3359) );
  OAI21_X1 U4200 ( .B1(n3361), .B2(n4541), .A(n3359), .ZN(U3467) );
  NAND2_X1 U4201 ( .A1(n2751), .A2(REG1_REG_0__SCAN_IN), .ZN(n3360) );
  OAI21_X1 U4202 ( .B1(n3361), .B2(n2751), .A(n3360), .ZN(U3518) );
  INV_X1 U4203 ( .A(n3363), .ZN(n3364) );
  AOI21_X1 U4204 ( .B1(n3365), .B2(n3362), .A(n3364), .ZN(n3371) );
  NAND2_X1 U4205 ( .A1(n3367), .A2(n3366), .ZN(n3548) );
  AOI22_X1 U4206 ( .A1(n3667), .A2(n3842), .B1(REG3_REG_2__SCAN_IN), .B2(n3548), .ZN(n3370) );
  AOI22_X1 U4207 ( .A1(n3671), .A2(n2890), .B1(n2935), .B2(n3368), .ZN(n3369)
         );
  OAI211_X1 U4208 ( .C1(n3371), .C2(n3674), .A(n3370), .B(n3369), .ZN(U3234)
         );
  OAI21_X1 U4209 ( .B1(n3374), .B2(n3373), .A(n3372), .ZN(n3854) );
  AOI22_X1 U4210 ( .A1(n3671), .A2(n3842), .B1(REG3_REG_0__SCAN_IN), .B2(n3548), .ZN(n3377) );
  NAND2_X1 U4211 ( .A1(n2935), .A2(n3375), .ZN(n3376) );
  OAI211_X1 U4212 ( .C1(n3674), .C2(n3854), .A(n3377), .B(n3376), .ZN(U3229)
         );
  INV_X1 U4213 ( .A(n3378), .ZN(n3385) );
  INV_X1 U4214 ( .A(n3835), .ZN(n3539) );
  INV_X1 U4215 ( .A(REG2_REG_28__SCAN_IN), .ZN(n3379) );
  OAI22_X1 U4216 ( .A1(n4171), .A2(n3379), .B1(n3540), .B2(n4169), .ZN(n3380)
         );
  AOI21_X1 U4217 ( .B1(n3929), .B2(n4552), .A(n3380), .ZN(n3381) );
  OAI21_X1 U4218 ( .B1(n3539), .B2(n4559), .A(n3381), .ZN(n3384) );
  NOR2_X1 U4219 ( .A1(n3382), .A2(n4142), .ZN(n3383) );
  AOI211_X1 U4220 ( .C1(n4373), .C2(n3385), .A(n3384), .B(n3383), .ZN(n3386)
         );
  OAI21_X1 U4221 ( .B1(n3387), .B2(n4193), .A(n3386), .ZN(U3262) );
  INV_X1 U4222 ( .A(n3389), .ZN(n3390) );
  NAND2_X1 U4223 ( .A1(n3392), .A2(n3391), .ZN(n3619) );
  NAND2_X1 U4224 ( .A1(n4290), .A2(n3532), .ZN(n3394) );
  NAND2_X1 U4225 ( .A1(n3396), .A2(n2896), .ZN(n3393) );
  NAND2_X1 U4226 ( .A1(n3394), .A2(n3393), .ZN(n3395) );
  XNOR2_X1 U4227 ( .A(n3395), .B(n3487), .ZN(n3621) );
  AOI22_X1 U4228 ( .A1(n4290), .A2(n2135), .B1(n3532), .B2(n3396), .ZN(n3620)
         );
  NAND2_X1 U4229 ( .A1(n4186), .A2(n3532), .ZN(n3398) );
  OR2_X1 U4230 ( .A1(n4274), .A2(n3445), .ZN(n3397) );
  NAND2_X1 U4231 ( .A1(n3398), .A2(n3397), .ZN(n3399) );
  XNOR2_X1 U4232 ( .A(n3399), .B(n3530), .ZN(n3403) );
  NAND2_X1 U4233 ( .A1(n4186), .A2(n2135), .ZN(n3401) );
  OR2_X1 U4234 ( .A1(n4274), .A2(n3276), .ZN(n3400) );
  NAND2_X1 U4235 ( .A1(n3401), .A2(n3400), .ZN(n3404) );
  AND2_X1 U4236 ( .A1(n3403), .A2(n3404), .ZN(n3494) );
  INV_X1 U4237 ( .A(n3494), .ZN(n3402) );
  INV_X1 U4238 ( .A(n3403), .ZN(n3406) );
  INV_X1 U4239 ( .A(n3404), .ZN(n3405) );
  NAND2_X1 U4240 ( .A1(n3415), .A2(n3532), .ZN(n3408) );
  NAND2_X1 U4241 ( .A1(n4181), .A2(n2896), .ZN(n3407) );
  NAND2_X1 U4242 ( .A1(n3408), .A2(n3407), .ZN(n3409) );
  XNOR2_X1 U4243 ( .A(n3409), .B(n3487), .ZN(n3413) );
  NOR2_X1 U4244 ( .A1(n3414), .A2(n3413), .ZN(n3572) );
  AOI22_X1 U4245 ( .A1(n4179), .A2(n3532), .B1(n2223), .B2(n2896), .ZN(n3410)
         );
  XNOR2_X1 U4246 ( .A(n3410), .B(n3530), .ZN(n3412) );
  AOI22_X1 U4247 ( .A1(n4179), .A2(n2135), .B1(n2223), .B2(n3532), .ZN(n3411)
         );
  NAND2_X1 U4248 ( .A1(n3412), .A2(n3411), .ZN(n3418) );
  OAI21_X1 U4249 ( .B1(n3412), .B2(n3411), .A(n3418), .ZN(n3573) );
  NOR2_X1 U4250 ( .A1(n3572), .A2(n3573), .ZN(n3421) );
  NAND2_X1 U4251 ( .A1(n3414), .A2(n3413), .ZN(n3661) );
  NAND2_X1 U4252 ( .A1(n3415), .A2(n2135), .ZN(n3417) );
  NAND2_X1 U4253 ( .A1(n4181), .A2(n3532), .ZN(n3416) );
  NAND2_X1 U4254 ( .A1(n3417), .A2(n3416), .ZN(n3663) );
  NAND2_X1 U4255 ( .A1(n3661), .A2(n3663), .ZN(n3420) );
  INV_X1 U4256 ( .A(n3418), .ZN(n3419) );
  AOI22_X1 U4257 ( .A1(n3642), .A2(n3532), .B1(n2896), .B2(n3598), .ZN(n3422)
         );
  XNOR2_X1 U4258 ( .A(n3422), .B(n3530), .ZN(n3424) );
  AOI22_X1 U4259 ( .A1(n3642), .A2(n2135), .B1(n3532), .B2(n3598), .ZN(n3423)
         );
  NOR2_X1 U4260 ( .A1(n3424), .A2(n3423), .ZN(n3594) );
  NAND2_X1 U4261 ( .A1(n3424), .A2(n3423), .ZN(n3592) );
  NAND2_X1 U4262 ( .A1(n4113), .A2(n2135), .ZN(n3426) );
  OR2_X1 U4263 ( .A1(n4134), .A2(n3276), .ZN(n3425) );
  NAND2_X1 U4264 ( .A1(n3426), .A2(n3425), .ZN(n3638) );
  NAND2_X1 U4265 ( .A1(n4113), .A2(n3532), .ZN(n3428) );
  OR2_X1 U4266 ( .A1(n4134), .A2(n3445), .ZN(n3427) );
  NAND2_X1 U4267 ( .A1(n3428), .A2(n3427), .ZN(n3429) );
  XNOR2_X1 U4268 ( .A(n3429), .B(n3530), .ZN(n3639) );
  NAND2_X1 U4269 ( .A1(n4125), .A2(n3532), .ZN(n3431) );
  NAND2_X1 U4270 ( .A1(n3522), .A2(n2896), .ZN(n3430) );
  NAND2_X1 U4271 ( .A1(n3431), .A2(n3430), .ZN(n3432) );
  XNOR2_X1 U4272 ( .A(n3432), .B(n3487), .ZN(n3434) );
  AOI22_X1 U4273 ( .A1(n4125), .A2(n2135), .B1(n3532), .B2(n3522), .ZN(n3433)
         );
  NOR2_X1 U4274 ( .A1(n3434), .A2(n3433), .ZN(n3517) );
  AOI21_X1 U4275 ( .B1(n3638), .B2(n3639), .A(n3517), .ZN(n3437) );
  AND2_X1 U4276 ( .A1(n3434), .A2(n3433), .ZN(n3516) );
  NAND2_X1 U4277 ( .A1(n3836), .A2(n3532), .ZN(n3439) );
  NAND2_X1 U4278 ( .A1(n2896), .A2(n4095), .ZN(n3438) );
  NAND2_X1 U4279 ( .A1(n3439), .A2(n3438), .ZN(n3440) );
  XNOR2_X1 U4280 ( .A(n3440), .B(n3487), .ZN(n3444) );
  NOR2_X1 U4281 ( .A1(n3441), .A2(n3276), .ZN(n3442) );
  AOI21_X1 U4282 ( .B1(n3836), .B2(n2135), .A(n3442), .ZN(n3443) );
  NOR2_X1 U4283 ( .A1(n3444), .A2(n3443), .ZN(n3611) );
  AND2_X1 U4284 ( .A1(n3444), .A2(n3443), .ZN(n3557) );
  NAND2_X1 U4285 ( .A1(n4082), .A2(n3532), .ZN(n3447) );
  OR2_X1 U4286 ( .A1(n3445), .A2(n4238), .ZN(n3446) );
  NAND2_X1 U4287 ( .A1(n3447), .A2(n3446), .ZN(n3448) );
  XNOR2_X1 U4288 ( .A(n3448), .B(n3530), .ZN(n3454) );
  INV_X1 U4289 ( .A(n3454), .ZN(n3452) );
  NAND2_X1 U4290 ( .A1(n4082), .A2(n2135), .ZN(n3450) );
  NAND2_X1 U4291 ( .A1(n3532), .A2(n4074), .ZN(n3449) );
  NAND2_X1 U4292 ( .A1(n3450), .A2(n3449), .ZN(n3453) );
  INV_X1 U4293 ( .A(n3453), .ZN(n3451) );
  NAND2_X1 U4294 ( .A1(n3452), .A2(n3451), .ZN(n3553) );
  AND2_X1 U4295 ( .A1(n3454), .A2(n3453), .ZN(n3554) );
  OAI22_X1 U4296 ( .A1(n4239), .A2(n3455), .B1(n3276), .B2(n4060), .ZN(n3462)
         );
  OAI22_X1 U4297 ( .A1(n4239), .A2(n3276), .B1(n3445), .B2(n4060), .ZN(n3456)
         );
  XNOR2_X1 U4298 ( .A(n3456), .B(n3530), .ZN(n3461) );
  XOR2_X1 U4299 ( .A(n3462), .B(n3461), .Z(n3630) );
  NAND2_X1 U4300 ( .A1(n4057), .A2(n3532), .ZN(n3458) );
  OR2_X1 U4301 ( .A1(n3445), .A2(n4033), .ZN(n3457) );
  NAND2_X1 U4302 ( .A1(n3458), .A2(n3457), .ZN(n3459) );
  XNOR2_X1 U4303 ( .A(n3459), .B(n3530), .ZN(n3467) );
  NOR2_X1 U4304 ( .A1(n3276), .A2(n4033), .ZN(n3460) );
  AOI21_X1 U4305 ( .B1(n4057), .B2(n2135), .A(n3460), .ZN(n3468) );
  XNOR2_X1 U4306 ( .A(n3467), .B(n3468), .ZN(n3505) );
  INV_X1 U4307 ( .A(n3461), .ZN(n3464) );
  INV_X1 U4308 ( .A(n3462), .ZN(n3463) );
  NAND2_X1 U4309 ( .A1(n3464), .A2(n3463), .ZN(n3506) );
  NAND2_X1 U4310 ( .A1(n3504), .A2(n3465), .ZN(n3503) );
  NOR2_X1 U4311 ( .A1(n3276), .A2(n4224), .ZN(n3466) );
  AOI21_X1 U4312 ( .B1(n3990), .B2(n2135), .A(n3466), .ZN(n3471) );
  INV_X1 U4313 ( .A(n3467), .ZN(n3469) );
  OR2_X1 U4314 ( .A1(n3469), .A2(n3468), .ZN(n3472) );
  NAND3_X1 U4315 ( .A1(n3503), .A2(n3471), .A3(n3472), .ZN(n3602) );
  OAI22_X1 U4316 ( .A1(n4034), .A2(n3276), .B1(n3445), .B2(n4224), .ZN(n3470)
         );
  XNOR2_X1 U4317 ( .A(n3470), .B(n3530), .ZN(n3605) );
  AOI21_X1 U4318 ( .B1(n3503), .B2(n3472), .A(n3471), .ZN(n3604) );
  NAND2_X1 U4319 ( .A1(n3973), .A2(n3532), .ZN(n3474) );
  OR2_X1 U4320 ( .A1(n3445), .A2(n3993), .ZN(n3473) );
  NAND2_X1 U4321 ( .A1(n3474), .A2(n3473), .ZN(n3475) );
  XNOR2_X1 U4322 ( .A(n3475), .B(n3487), .ZN(n3478) );
  NOR2_X1 U4323 ( .A1(n3276), .A2(n3993), .ZN(n3476) );
  AOI21_X1 U4324 ( .B1(n3973), .B2(n2135), .A(n3476), .ZN(n3477) );
  OR2_X1 U4325 ( .A1(n3478), .A2(n3477), .ZN(n3566) );
  NAND2_X1 U4326 ( .A1(n3961), .A2(n3532), .ZN(n3480) );
  OR2_X1 U4327 ( .A1(n3445), .A2(n3978), .ZN(n3479) );
  NAND2_X1 U4328 ( .A1(n3480), .A2(n3479), .ZN(n3481) );
  XNOR2_X1 U4329 ( .A(n3481), .B(n3487), .ZN(n3484) );
  NOR2_X1 U4330 ( .A1(n3276), .A2(n3978), .ZN(n3482) );
  AOI21_X1 U4331 ( .B1(n3961), .B2(n2135), .A(n3482), .ZN(n3483) );
  NOR2_X1 U4332 ( .A1(n3484), .A2(n3483), .ZN(n3649) );
  NAND2_X1 U4333 ( .A1(n3972), .A2(n3532), .ZN(n3486) );
  OR2_X1 U4334 ( .A1(n3445), .A2(n4210), .ZN(n3485) );
  NAND2_X1 U4335 ( .A1(n3486), .A2(n3485), .ZN(n3488) );
  XNOR2_X1 U4336 ( .A(n3488), .B(n3487), .ZN(n3526) );
  NOR2_X1 U4337 ( .A1(n3276), .A2(n4210), .ZN(n3489) );
  AOI21_X1 U4338 ( .B1(n3972), .B2(n2135), .A(n3489), .ZN(n3525) );
  XNOR2_X1 U4339 ( .A(n3529), .B(n3528), .ZN(n3493) );
  INV_X1 U4340 ( .A(n3938), .ZN(n4211) );
  INV_X1 U4341 ( .A(REG3_REG_27__SCAN_IN), .ZN(n4592) );
  OAI22_X1 U4342 ( .A1(n3653), .A2(n4211), .B1(STATE_REG_SCAN_IN), .B2(n4592), 
        .ZN(n3491) );
  OAI22_X1 U4343 ( .A1(n3655), .A2(n3988), .B1(n3654), .B2(n3955), .ZN(n3490)
         );
  AOI211_X1 U4344 ( .C1(n3957), .C2(n2935), .A(n3491), .B(n3490), .ZN(n3492)
         );
  OAI21_X1 U4345 ( .B1(n3493), .B2(n3674), .A(n3492), .ZN(U3211) );
  NOR2_X1 U4346 ( .A1(n2170), .A2(n3494), .ZN(n3495) );
  XNOR2_X1 U4347 ( .A(n2166), .B(n3495), .ZN(n3502) );
  NAND2_X1 U4348 ( .A1(REG3_REG_14__SCAN_IN), .A2(U3149), .ZN(n4428) );
  OAI21_X1 U4349 ( .B1(n3655), .B2(n3496), .A(n4428), .ZN(n3499) );
  OAI22_X1 U4350 ( .A1(n3653), .A2(n4277), .B1(n3654), .B2(n3497), .ZN(n3498)
         );
  AOI211_X1 U4351 ( .C1(n3500), .C2(n2935), .A(n3499), .B(n3498), .ZN(n3501)
         );
  OAI21_X1 U4352 ( .B1(n3502), .B2(n3674), .A(n3501), .ZN(U3212) );
  NAND2_X1 U4353 ( .A1(n3503), .A2(n3635), .ZN(n3511) );
  AOI21_X1 U4354 ( .B1(n3504), .B2(n3506), .A(n3505), .ZN(n3510) );
  OAI22_X1 U4355 ( .A1(n3653), .A2(n4034), .B1(STATE_REG_SCAN_IN), .B2(n4810), 
        .ZN(n3508) );
  OAI22_X1 U4356 ( .A1(n3655), .A2(n4239), .B1(n3654), .B2(n4042), .ZN(n3507)
         );
  AOI211_X1 U4357 ( .C1(n4039), .C2(n2935), .A(n3508), .B(n3507), .ZN(n3509)
         );
  OAI21_X1 U4358 ( .B1(n3511), .B2(n3510), .A(n3509), .ZN(U3213) );
  INV_X1 U4359 ( .A(n3638), .ZN(n3515) );
  INV_X1 U4360 ( .A(n3512), .ZN(n3513) );
  OAI21_X1 U4361 ( .B1(n3513), .B2(n3638), .A(n3639), .ZN(n3514) );
  OAI21_X1 U4362 ( .B1(n3515), .B2(n3512), .A(n3514), .ZN(n3519) );
  NOR2_X1 U4363 ( .A1(n3517), .A2(n3516), .ZN(n3518) );
  XNOR2_X1 U4364 ( .A(n3519), .B(n3518), .ZN(n3524) );
  NAND2_X1 U4365 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n3923) );
  OAI21_X1 U4366 ( .B1(n3653), .B2(n4111), .A(n3923), .ZN(n3521) );
  INV_X1 U4367 ( .A(n4113), .ZN(n4146) );
  OAI22_X1 U4368 ( .A1(n3655), .A2(n4146), .B1(n3654), .B2(n4118), .ZN(n3520)
         );
  AOI211_X1 U4369 ( .C1(n3522), .C2(n2935), .A(n3521), .B(n3520), .ZN(n3523)
         );
  OAI21_X1 U4370 ( .B1(n3524), .B2(n3674), .A(n3523), .ZN(U3216) );
  AOI22_X1 U4371 ( .A1(n3938), .A2(n3532), .B1(n2896), .B2(n3929), .ZN(n3531)
         );
  XNOR2_X1 U4372 ( .A(n3531), .B(n3530), .ZN(n3535) );
  AOI22_X1 U4373 ( .A1(n3938), .A2(n2135), .B1(n3532), .B2(n3929), .ZN(n3534)
         );
  XNOR2_X1 U4374 ( .A(n3535), .B(n3534), .ZN(n3536) );
  XNOR2_X1 U4375 ( .A(n3537), .B(n3536), .ZN(n3538) );
  NAND2_X1 U4376 ( .A1(n3538), .A2(n3635), .ZN(n3544) );
  INV_X1 U4377 ( .A(REG3_REG_28__SCAN_IN), .ZN(n4594) );
  OAI22_X1 U4378 ( .A1(n3653), .A2(n3539), .B1(STATE_REG_SCAN_IN), .B2(n4594), 
        .ZN(n3542) );
  OAI22_X1 U4379 ( .A1(n3655), .A2(n3652), .B1(n3654), .B2(n3540), .ZN(n3541)
         );
  AOI211_X1 U4380 ( .C1(n3929), .C2(n2935), .A(n3542), .B(n3541), .ZN(n3543)
         );
  NAND2_X1 U4381 ( .A1(n3544), .A2(n3543), .ZN(U3217) );
  OAI211_X1 U4382 ( .C1(n3545), .C2(n3547), .A(n3546), .B(n3635), .ZN(n3552)
         );
  AOI22_X1 U4383 ( .A1(n3667), .A2(n2897), .B1(n3548), .B2(REG3_REG_1__SCAN_IN), .ZN(n3551) );
  AOI22_X1 U4384 ( .A1(n3671), .A2(n3841), .B1(n2935), .B2(n3549), .ZN(n3550)
         );
  NAND3_X1 U4385 ( .A1(n3552), .A2(n3551), .A3(n3550), .ZN(U3219) );
  INV_X1 U4386 ( .A(n3553), .ZN(n3555) );
  NOR2_X1 U4387 ( .A1(n3555), .A2(n3554), .ZN(n3559) );
  AOI211_X1 U4388 ( .C1(n3556), .C2(n2259), .A(n3611), .B(n3559), .ZN(n3558)
         );
  AOI211_X1 U4389 ( .C1(n3560), .C2(n3559), .A(n3674), .B(n3558), .ZN(n3564)
         );
  OAI22_X1 U4390 ( .A1(n3655), .A2(n4111), .B1(n3654), .B2(n4071), .ZN(n3563)
         );
  AOI22_X1 U4391 ( .A1(n3671), .A2(n4036), .B1(REG3_REG_21__SCAN_IN), .B2(
        U3149), .ZN(n3561) );
  OAI21_X1 U4392 ( .B1(n3668), .B2(n4238), .A(n3561), .ZN(n3562) );
  OR3_X1 U4393 ( .A1(n3564), .A2(n3563), .A3(n3562), .ZN(U3220) );
  NAND2_X1 U4394 ( .A1(n2164), .A2(n3566), .ZN(n3567) );
  XNOR2_X1 U4395 ( .A(n3565), .B(n3567), .ZN(n3571) );
  INV_X1 U4396 ( .A(REG3_REG_25__SCAN_IN), .ZN(n4822) );
  OAI22_X1 U4397 ( .A1(n3653), .A2(n3988), .B1(STATE_REG_SCAN_IN), .B2(n4822), 
        .ZN(n3569) );
  OAI22_X1 U4398 ( .A1(n3655), .A2(n4034), .B1(n3654), .B2(n3996), .ZN(n3568)
         );
  AOI211_X1 U4399 ( .C1(n2234), .C2(n2935), .A(n3569), .B(n3568), .ZN(n3570)
         );
  OAI21_X1 U4400 ( .B1(n3571), .B2(n3674), .A(n3570), .ZN(U3222) );
  OAI21_X1 U4401 ( .B1(n3572), .B2(n3663), .A(n3661), .ZN(n3574) );
  XNOR2_X1 U4402 ( .A(n3574), .B(n3573), .ZN(n3578) );
  INV_X1 U4403 ( .A(n3642), .ZN(n4261) );
  NAND2_X1 U4404 ( .A1(U3149), .A2(REG3_REG_16__SCAN_IN), .ZN(n4445) );
  OAI21_X1 U4405 ( .B1(n3653), .B2(n4261), .A(n4445), .ZN(n3576) );
  OAI22_X1 U4406 ( .A1(n3655), .A2(n4277), .B1(n3654), .B2(n4170), .ZN(n3575)
         );
  AOI211_X1 U4407 ( .C1(n2223), .C2(n2935), .A(n3576), .B(n3575), .ZN(n3577)
         );
  OAI21_X1 U4408 ( .B1(n3578), .B2(n3674), .A(n3577), .ZN(U3223) );
  OAI211_X1 U4409 ( .C1(n3581), .C2(n3580), .A(n3579), .B(n3635), .ZN(n3590)
         );
  INV_X1 U4410 ( .A(n3582), .ZN(n3583) );
  AOI22_X1 U4411 ( .A1(n3671), .A2(n3584), .B1(n3666), .B2(n3583), .ZN(n3589)
         );
  NOR2_X1 U4412 ( .A1(n3668), .A2(n3585), .ZN(n3586) );
  AOI211_X1 U4413 ( .C1(n3667), .C2(n3840), .A(n3587), .B(n3586), .ZN(n3588)
         );
  NAND3_X1 U4414 ( .A1(n3590), .A2(n3589), .A3(n3588), .ZN(U3224) );
  INV_X1 U4415 ( .A(n3592), .ZN(n3593) );
  NOR2_X1 U4416 ( .A1(n3594), .A2(n3593), .ZN(n3595) );
  XNOR2_X1 U4417 ( .A(n3591), .B(n3595), .ZN(n3601) );
  INV_X1 U4418 ( .A(n4153), .ZN(n3596) );
  AOI22_X1 U4419 ( .A1(n3667), .A2(n4179), .B1(n3666), .B2(n3596), .ZN(n3600)
         );
  NOR2_X1 U4420 ( .A1(STATE_REG_SCAN_IN), .A2(n4599), .ZN(n4456) );
  NOR2_X1 U4421 ( .A1(n3653), .A2(n4146), .ZN(n3597) );
  AOI211_X1 U4422 ( .C1(n3598), .C2(n2935), .A(n4456), .B(n3597), .ZN(n3599)
         );
  OAI211_X1 U4423 ( .C1(n3601), .C2(n3674), .A(n3600), .B(n3599), .ZN(U3225)
         );
  INV_X1 U4424 ( .A(n3602), .ZN(n3603) );
  NOR2_X1 U4425 ( .A1(n3604), .A2(n3603), .ZN(n3606) );
  XNOR2_X1 U4426 ( .A(n3606), .B(n3605), .ZN(n3610) );
  OAI22_X1 U4427 ( .A1(n3653), .A2(n4225), .B1(STATE_REG_SCAN_IN), .B2(n4600), 
        .ZN(n3608) );
  OAI22_X1 U4428 ( .A1(n3655), .A2(n4008), .B1(n3654), .B2(n4012), .ZN(n3607)
         );
  AOI211_X1 U4429 ( .C1(n2235), .C2(n2935), .A(n3608), .B(n3607), .ZN(n3609)
         );
  OAI21_X1 U4430 ( .B1(n3610), .B2(n3674), .A(n3609), .ZN(U3226) );
  NAND2_X1 U4431 ( .A1(n2253), .A2(n2259), .ZN(n3612) );
  AOI22_X1 U4432 ( .A1(n3613), .A2(n2259), .B1(n3556), .B2(n3612), .ZN(n3618)
         );
  INV_X1 U4433 ( .A(REG3_REG_20__SCAN_IN), .ZN(n3614) );
  OAI22_X1 U4434 ( .A1(n3653), .A2(n3631), .B1(STATE_REG_SCAN_IN), .B2(n3614), 
        .ZN(n3616) );
  INV_X1 U4435 ( .A(n4125), .ZN(n4084) );
  OAI22_X1 U4436 ( .A1(n3655), .A2(n4084), .B1(n3654), .B2(n4096), .ZN(n3615)
         );
  AOI211_X1 U4437 ( .C1(n4095), .C2(n2935), .A(n3616), .B(n3615), .ZN(n3617)
         );
  OAI21_X1 U4438 ( .B1(n3618), .B2(n3674), .A(n3617), .ZN(U3230) );
  XNOR2_X1 U4439 ( .A(n3621), .B(n3620), .ZN(n3622) );
  XNOR2_X1 U4440 ( .A(n3619), .B(n3622), .ZN(n3628) );
  AOI22_X1 U4441 ( .A1(n3667), .A2(n3837), .B1(n3666), .B2(n3623), .ZN(n3627)
         );
  AND2_X1 U4442 ( .A1(U3149), .A2(REG3_REG_13__SCAN_IN), .ZN(n4413) );
  NOR2_X1 U4443 ( .A1(n3668), .A2(n3624), .ZN(n3625) );
  AOI211_X1 U4444 ( .C1(n3671), .C2(n4186), .A(n4413), .B(n3625), .ZN(n3626)
         );
  OAI211_X1 U4445 ( .C1(n3628), .C2(n3674), .A(n3627), .B(n3626), .ZN(U3231)
         );
  OAI21_X1 U4446 ( .B1(n3630), .B2(n3629), .A(n3504), .ZN(n3636) );
  OAI22_X1 U4447 ( .A1(n3655), .A2(n3631), .B1(n3654), .B2(n4051), .ZN(n3634)
         );
  AOI22_X1 U4448 ( .A1(n3671), .A2(n4057), .B1(REG3_REG_22__SCAN_IN), .B2(
        U3149), .ZN(n3632) );
  OAI21_X1 U4449 ( .B1(n3668), .B2(n4060), .A(n3632), .ZN(n3633) );
  AOI211_X1 U4450 ( .C1(n3636), .C2(n3635), .A(n3634), .B(n3633), .ZN(n3637)
         );
  INV_X1 U4451 ( .A(n3637), .ZN(U3232) );
  XNOR2_X1 U4452 ( .A(n3639), .B(n3638), .ZN(n3640) );
  XNOR2_X1 U4453 ( .A(n3512), .B(n3640), .ZN(n3647) );
  INV_X1 U4454 ( .A(n3641), .ZN(n4135) );
  AOI22_X1 U4455 ( .A1(n3667), .A2(n3642), .B1(n3666), .B2(n4135), .ZN(n3646)
         );
  NOR2_X1 U4456 ( .A1(n3643), .A2(STATE_REG_SCAN_IN), .ZN(n4472) );
  NOR2_X1 U4457 ( .A1(n3653), .A2(n4084), .ZN(n3644) );
  AOI211_X1 U4458 ( .C1(n4124), .C2(n2935), .A(n4472), .B(n3644), .ZN(n3645)
         );
  OAI211_X1 U4459 ( .C1(n3647), .C2(n3674), .A(n3646), .B(n3645), .ZN(U3235)
         );
  NOR2_X1 U4460 ( .A1(n3649), .A2(n2157), .ZN(n3650) );
  XNOR2_X1 U4461 ( .A(n3648), .B(n3650), .ZN(n3660) );
  INV_X1 U4462 ( .A(REG3_REG_26__SCAN_IN), .ZN(n3651) );
  OAI22_X1 U4463 ( .A1(n3653), .A2(n3652), .B1(STATE_REG_SCAN_IN), .B2(n3651), 
        .ZN(n3657) );
  OAI22_X1 U4464 ( .A1(n3655), .A2(n4225), .B1(n3654), .B2(n3979), .ZN(n3656)
         );
  AOI211_X1 U4465 ( .C1(n3658), .C2(n2935), .A(n3657), .B(n3656), .ZN(n3659)
         );
  OAI21_X1 U4466 ( .B1(n3660), .B2(n3674), .A(n3659), .ZN(U3237) );
  INV_X1 U4467 ( .A(n3661), .ZN(n3662) );
  NOR2_X1 U4468 ( .A1(n3572), .A2(n3662), .ZN(n3664) );
  XNOR2_X1 U4469 ( .A(n3664), .B(n3663), .ZN(n3675) );
  INV_X1 U4470 ( .A(n3665), .ZN(n4180) );
  AOI22_X1 U4471 ( .A1(n3667), .A2(n4186), .B1(n3666), .B2(n4180), .ZN(n3673)
         );
  NAND2_X1 U4472 ( .A1(U3149), .A2(REG3_REG_15__SCAN_IN), .ZN(n4442) );
  INV_X1 U4473 ( .A(n4442), .ZN(n3670) );
  NOR2_X1 U4474 ( .A1(n3668), .A2(n4267), .ZN(n3669) );
  AOI211_X1 U4475 ( .C1(n3671), .C2(n4179), .A(n3670), .B(n3669), .ZN(n3672)
         );
  OAI211_X1 U4476 ( .C1(n3675), .C2(n3674), .A(n3673), .B(n3672), .ZN(U3238)
         );
  INV_X1 U4477 ( .A(n3676), .ZN(n3826) );
  NOR2_X1 U4478 ( .A1(n3677), .A2(n4835), .ZN(n4194) );
  INV_X1 U4479 ( .A(n4194), .ZN(n4197) );
  INV_X1 U4480 ( .A(n3940), .ZN(n3678) );
  AND2_X1 U4481 ( .A1(n3679), .A2(DATAI_30_), .ZN(n4204) );
  NOR2_X1 U4482 ( .A1(n3678), .A2(n4204), .ZN(n3736) );
  INV_X1 U4483 ( .A(n3736), .ZN(n3708) );
  NAND2_X1 U4484 ( .A1(n3679), .A2(DATAI_29_), .ZN(n3946) );
  NAND2_X1 U4485 ( .A1(n3835), .A2(n3946), .ZN(n3681) );
  INV_X1 U4486 ( .A(n3681), .ZN(n3744) );
  INV_X1 U4487 ( .A(n3680), .ZN(n3934) );
  NOR3_X1 U4488 ( .A1(n3744), .A2(n3934), .A3(n3741), .ZN(n3812) );
  INV_X1 U4489 ( .A(n3933), .ZN(n3702) );
  NOR2_X1 U4490 ( .A1(n3702), .A2(n3701), .ZN(n3686) );
  NAND2_X1 U4491 ( .A1(n3681), .A2(n3680), .ZN(n3685) );
  NOR2_X1 U4492 ( .A1(n3835), .A2(n3946), .ZN(n3745) );
  INV_X1 U4493 ( .A(n4204), .ZN(n3703) );
  AOI22_X1 U4494 ( .A1(n3682), .A2(REG0_REG_31__SCAN_IN), .B1(n2411), .B2(
        REG2_REG_31__SCAN_IN), .ZN(n3683) );
  OAI21_X1 U4495 ( .B1(n3684), .B2(n4857), .A(n3683), .ZN(n4196) );
  NAND2_X1 U4496 ( .A1(n4196), .A2(n4197), .ZN(n3817) );
  OAI21_X1 U4497 ( .B1(n3703), .B2(n3940), .A(n3817), .ZN(n3712) );
  NOR2_X1 U4498 ( .A1(n3745), .A2(n3712), .ZN(n3698) );
  OAI21_X1 U4499 ( .B1(n3686), .B2(n3685), .A(n3698), .ZN(n3820) );
  AOI21_X1 U4500 ( .B1(n3960), .B2(n3812), .A(n3820), .ZN(n3705) );
  AND2_X1 U4501 ( .A1(n2196), .A2(n3731), .ZN(n3809) );
  INV_X1 U4502 ( .A(n3809), .ZN(n3697) );
  NAND2_X1 U4503 ( .A1(n3687), .A2(n3690), .ZN(n3790) );
  NAND2_X1 U4504 ( .A1(n3689), .A2(n3688), .ZN(n3779) );
  NAND2_X1 U4505 ( .A1(n3779), .A2(n3690), .ZN(n3782) );
  OAI21_X1 U4506 ( .B1(n3691), .B2(n3790), .A(n3782), .ZN(n3692) );
  AOI21_X1 U4507 ( .B1(n3797), .B2(n3692), .A(n2190), .ZN(n3694) );
  OAI21_X1 U4508 ( .B1(n3694), .B2(n2141), .A(n3693), .ZN(n3695) );
  OAI221_X1 U4509 ( .B1(n3697), .B2(n3696), .C1(n3697), .C2(n3695), .A(n3816), 
        .ZN(n3700) );
  INV_X1 U4510 ( .A(n3698), .ZN(n3699) );
  NOR4_X1 U4511 ( .A1(n3702), .A2(n3701), .A3(n3700), .A4(n3699), .ZN(n3704)
         );
  OAI22_X1 U4512 ( .A1(n3705), .A2(n3704), .B1(n3703), .B2(n4196), .ZN(n3707)
         );
  NOR2_X1 U4513 ( .A1(n4196), .A2(n4197), .ZN(n3737) );
  INV_X1 U4514 ( .A(n3737), .ZN(n3706) );
  OAI211_X1 U4515 ( .C1(n4197), .C2(n3708), .A(n3707), .B(n3706), .ZN(n3825)
         );
  INV_X1 U4516 ( .A(n3709), .ZN(n3804) );
  INV_X1 U4517 ( .A(n4067), .ZN(n3713) );
  NOR4_X1 U4518 ( .A1(n3713), .A2(n3712), .A3(n3711), .A4(n3710), .ZN(n3727)
         );
  NAND2_X1 U4519 ( .A1(n4104), .A2(n4022), .ZN(n4145) );
  NOR4_X1 U4520 ( .A1(n3716), .A2(n3715), .A3(n4145), .A4(n3714), .ZN(n3726)
         );
  NOR4_X1 U4521 ( .A1(n3720), .A2(n3719), .A3(n3718), .A4(n3717), .ZN(n3725)
         );
  NOR4_X1 U4522 ( .A1(n3723), .A2(n3722), .A3(n4184), .A4(n3721), .ZN(n3724)
         );
  NAND4_X1 U4523 ( .A1(n3727), .A2(n3726), .A3(n3725), .A4(n3724), .ZN(n3751)
         );
  INV_X1 U4524 ( .A(n3967), .ZN(n3729) );
  NOR2_X1 U4525 ( .A1(n3729), .A2(n3728), .ZN(n3986) );
  INV_X1 U4526 ( .A(n3986), .ZN(n3735) );
  INV_X1 U4527 ( .A(n4085), .ZN(n3730) );
  OR2_X1 U4528 ( .A1(n4086), .A2(n3730), .ZN(n4109) );
  INV_X1 U4529 ( .A(n4109), .ZN(n3734) );
  NAND2_X1 U4530 ( .A1(n3732), .A2(n3731), .ZN(n4006) );
  NOR4_X1 U4531 ( .A1(n3735), .A2(n3734), .A3(n3733), .A4(n4006), .ZN(n3740)
         );
  NOR2_X1 U4532 ( .A1(n3737), .A2(n3736), .ZN(n3819) );
  NAND2_X1 U4533 ( .A1(n3739), .A2(n3738), .ZN(n4089) );
  NAND4_X1 U4534 ( .A1(n3740), .A2(n3960), .A3(n3819), .A4(n4089), .ZN(n3750)
         );
  INV_X1 U4535 ( .A(n3741), .ZN(n3743) );
  NAND2_X1 U4536 ( .A1(n3743), .A2(n3742), .ZN(n3969) );
  NOR4_X1 U4537 ( .A1(n3969), .A2(n3937), .A3(n3930), .A4(n4558), .ZN(n3748)
         );
  NOR2_X1 U4538 ( .A1(n4160), .A2(n4055), .ZN(n3746) );
  NAND4_X1 U4539 ( .A1(n3748), .A2(n3768), .A3(n3747), .A4(n3746), .ZN(n3749)
         );
  XNOR2_X1 U4540 ( .A(n4057), .B(n4039), .ZN(n4020) );
  INV_X1 U4541 ( .A(n4020), .ZN(n4031) );
  NOR4_X1 U4542 ( .A1(n3751), .A2(n3750), .A3(n3749), .A4(n4031), .ZN(n3752)
         );
  NOR2_X1 U4543 ( .A1(n3752), .A2(n2708), .ZN(n3823) );
  OAI211_X1 U4544 ( .C1(n3755), .C2(n2708), .A(n3754), .B(n3753), .ZN(n3757)
         );
  NAND3_X1 U4545 ( .A1(n3757), .A2(n3756), .A3(n2678), .ZN(n3760) );
  NAND3_X1 U4546 ( .A1(n3760), .A2(n3759), .A3(n3758), .ZN(n3763) );
  NAND3_X1 U4547 ( .A1(n3763), .A2(n3762), .A3(n3761), .ZN(n3766) );
  NAND4_X1 U4548 ( .A1(n3766), .A2(n3765), .A3(n3777), .A4(n3764), .ZN(n3769)
         );
  NAND3_X1 U4549 ( .A1(n3769), .A2(n3768), .A3(n3767), .ZN(n3770) );
  NAND3_X1 U4550 ( .A1(n3770), .A2(n3776), .A3(n3775), .ZN(n3773) );
  AND3_X1 U4551 ( .A1(n3773), .A2(n3772), .A3(n3771), .ZN(n3780) );
  INV_X1 U4552 ( .A(n3782), .ZN(n3794) );
  NAND4_X1 U4553 ( .A1(n3777), .A2(n2215), .A3(n3776), .A4(n3775), .ZN(n3778)
         );
  OAI22_X1 U4554 ( .A1(n3780), .A2(n3779), .B1(n3794), .B2(n3778), .ZN(n3784)
         );
  INV_X1 U4555 ( .A(n3781), .ZN(n3783) );
  AOI22_X1 U4556 ( .A1(n3784), .A2(n2168), .B1(n3783), .B2(n3782), .ZN(n3796)
         );
  NAND3_X1 U4557 ( .A1(n3791), .A2(n3786), .A3(n3785), .ZN(n3795) );
  INV_X1 U4558 ( .A(n3787), .ZN(n3792) );
  INV_X1 U4559 ( .A(n3788), .ZN(n3789) );
  AOI211_X1 U4560 ( .C1(n3792), .C2(n3791), .A(n3790), .B(n3789), .ZN(n3793)
         );
  OAI22_X1 U4561 ( .A1(n3796), .A2(n3795), .B1(n3794), .B2(n3793), .ZN(n3800)
         );
  INV_X1 U4562 ( .A(n3797), .ZN(n3798) );
  AOI21_X1 U4563 ( .B1(n3800), .B2(n3799), .A(n3798), .ZN(n3803) );
  INV_X1 U4564 ( .A(n3801), .ZN(n3802) );
  OAI21_X1 U4565 ( .B1(n3803), .B2(n3802), .A(n4026), .ZN(n3805) );
  NAND2_X1 U4566 ( .A1(n3805), .A2(n3804), .ZN(n3807) );
  AOI21_X1 U4567 ( .B1(n3808), .B2(n3807), .A(n3806), .ZN(n3811) );
  OAI21_X1 U4568 ( .B1(n3811), .B2(n3810), .A(n3809), .ZN(n3815) );
  INV_X1 U4569 ( .A(n3812), .ZN(n3813) );
  AOI211_X1 U4570 ( .C1(n3816), .C2(n3815), .A(n3814), .B(n3813), .ZN(n3821)
         );
  INV_X1 U4571 ( .A(n3817), .ZN(n3818) );
  OAI22_X1 U4572 ( .A1(n3821), .A2(n3820), .B1(n3819), .B2(n3818), .ZN(n3822)
         );
  MUX2_X1 U4573 ( .A(n3823), .B(n3822), .S(n2756), .Z(n3824) );
  AOI21_X1 U4574 ( .B1(n3826), .B2(n3825), .A(n3824), .ZN(n3827) );
  XNOR2_X1 U4575 ( .A(n3827), .B(n4358), .ZN(n3834) );
  INV_X1 U4576 ( .A(n3829), .ZN(n3833) );
  NAND2_X1 U4577 ( .A1(n3829), .A2(n3828), .ZN(n3830) );
  OAI211_X1 U4578 ( .C1(n3831), .C2(n3855), .A(B_REG_SCAN_IN), .B(n3830), .ZN(
        n3832) );
  OAI21_X1 U4579 ( .B1(n3834), .B2(n3833), .A(n3832), .ZN(U3239) );
  MUX2_X1 U4580 ( .A(DATAO_REG_31__SCAN_IN), .B(n4196), .S(U4043), .Z(U3581)
         );
  MUX2_X1 U4581 ( .A(n3835), .B(DATAO_REG_29__SCAN_IN), .S(n3856), .Z(U3579)
         );
  MUX2_X1 U4582 ( .A(n3938), .B(DATAO_REG_28__SCAN_IN), .S(n3856), .Z(U3578)
         );
  MUX2_X1 U4583 ( .A(n3972), .B(DATAO_REG_27__SCAN_IN), .S(n3856), .Z(U3577)
         );
  MUX2_X1 U4584 ( .A(n3973), .B(DATAO_REG_25__SCAN_IN), .S(n3856), .Z(U3575)
         );
  MUX2_X1 U4585 ( .A(n3990), .B(DATAO_REG_24__SCAN_IN), .S(n3856), .Z(U3574)
         );
  MUX2_X1 U4586 ( .A(n4036), .B(DATAO_REG_22__SCAN_IN), .S(n3856), .Z(U3572)
         );
  MUX2_X1 U4587 ( .A(n3836), .B(DATAO_REG_20__SCAN_IN), .S(n3856), .Z(U3570)
         );
  MUX2_X1 U4588 ( .A(n4125), .B(DATAO_REG_19__SCAN_IN), .S(n3856), .Z(U3569)
         );
  MUX2_X1 U4589 ( .A(n4290), .B(DATAO_REG_13__SCAN_IN), .S(n3856), .Z(U3563)
         );
  MUX2_X1 U4590 ( .A(n3837), .B(DATAO_REG_12__SCAN_IN), .S(n3856), .Z(U3562)
         );
  MUX2_X1 U4591 ( .A(n3838), .B(DATAO_REG_8__SCAN_IN), .S(n3856), .Z(U3558) );
  MUX2_X1 U4592 ( .A(n3839), .B(DATAO_REG_7__SCAN_IN), .S(n3856), .Z(U3557) );
  MUX2_X1 U4593 ( .A(n3840), .B(DATAO_REG_4__SCAN_IN), .S(n3856), .Z(U3554) );
  MUX2_X1 U4594 ( .A(n2890), .B(DATAO_REG_3__SCAN_IN), .S(n3856), .Z(U3553) );
  MUX2_X1 U4595 ( .A(n3841), .B(DATAO_REG_2__SCAN_IN), .S(n3856), .Z(U3552) );
  MUX2_X1 U4596 ( .A(n3842), .B(DATAO_REG_1__SCAN_IN), .S(n3856), .Z(U3551) );
  OAI211_X1 U4597 ( .C1(n3844), .C2(n3843), .A(n4464), .B(n3863), .ZN(n3850)
         );
  OAI211_X1 U4598 ( .C1(n3846), .C2(n3857), .A(n4482), .B(n3845), .ZN(n3849)
         );
  AOI22_X1 U4599 ( .A1(n4473), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n3848) );
  INV_X1 U4600 ( .A(n4485), .ZN(n4441) );
  NAND2_X1 U4601 ( .A1(n4441), .A2(n4366), .ZN(n3847) );
  NAND4_X1 U4602 ( .A1(n3850), .A2(n3849), .A3(n3848), .A4(n3847), .ZN(U3241)
         );
  INV_X1 U4603 ( .A(REG2_REG_0__SCAN_IN), .ZN(n4804) );
  AND2_X1 U4604 ( .A1(n4378), .A2(n4804), .ZN(n3851) );
  NOR2_X1 U4605 ( .A1(n4368), .A2(n3851), .ZN(n4377) );
  NAND3_X1 U4606 ( .A1(n3854), .A2(n3853), .A3(n3852), .ZN(n3860) );
  INV_X1 U4607 ( .A(n3855), .ZN(n3858) );
  AOI21_X1 U4608 ( .B1(n3858), .B2(n3857), .A(n3856), .ZN(n3859) );
  OAI211_X1 U4609 ( .C1(IR_REG_0__SCAN_IN), .C2(n4377), .A(n3860), .B(n3859), 
        .ZN(n3887) );
  AOI22_X1 U4610 ( .A1(ADDR_REG_2__SCAN_IN), .A2(n4473), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n3875) );
  MUX2_X1 U4611 ( .A(REG1_REG_2__SCAN_IN), .B(n2805), .S(n2134), .Z(n3861) );
  NAND3_X1 U4612 ( .A1(n3863), .A2(n3862), .A3(n3861), .ZN(n3864) );
  NAND3_X1 U4613 ( .A1(n4464), .A2(n3865), .A3(n3864), .ZN(n3871) );
  MUX2_X1 U4614 ( .A(REG2_REG_2__SCAN_IN), .B(n2801), .S(n2134), .Z(n3866) );
  NAND2_X1 U4615 ( .A1(n3867), .A2(n3866), .ZN(n3868) );
  NAND3_X1 U4616 ( .A1(n4482), .A2(n3869), .A3(n3868), .ZN(n3870) );
  OAI211_X1 U4617 ( .C1(n4485), .C2(n2134), .A(n3871), .B(n3870), .ZN(n3873)
         );
  INV_X1 U4618 ( .A(n3873), .ZN(n3874) );
  NAND3_X1 U4619 ( .A1(n3887), .A2(n3875), .A3(n3874), .ZN(U3242) );
  NAND2_X1 U4620 ( .A1(n4473), .A2(ADDR_REG_4__SCAN_IN), .ZN(n3886) );
  OAI21_X1 U4621 ( .B1(n4485), .B2(n3877), .A(n3876), .ZN(n3881) );
  XNOR2_X1 U4622 ( .A(n3878), .B(REG1_REG_4__SCAN_IN), .ZN(n3879) );
  NOR2_X1 U4623 ( .A1(n4468), .A2(n3879), .ZN(n3880) );
  NOR2_X1 U4624 ( .A1(n3881), .A2(n3880), .ZN(n3885) );
  XNOR2_X1 U4625 ( .A(n3882), .B(REG2_REG_4__SCAN_IN), .ZN(n3883) );
  NAND2_X1 U4626 ( .A1(n4482), .A2(n3883), .ZN(n3884) );
  NAND4_X1 U4627 ( .A1(n3887), .A2(n3886), .A3(n3885), .A4(n3884), .ZN(U3244)
         );
  AOI22_X1 U4628 ( .A1(REG1_REG_18__SCAN_IN), .A2(n4490), .B1(n3919), .B2(
        n4695), .ZN(n4469) );
  INV_X1 U4629 ( .A(n3918), .ZN(n4492) );
  AOI22_X1 U4630 ( .A1(n3918), .A2(REG1_REG_17__SCAN_IN), .B1(n4858), .B2(
        n4492), .ZN(n4462) );
  AOI22_X1 U4631 ( .A1(REG1_REG_11__SCAN_IN), .A2(n4501), .B1(n3901), .B2(
        n4300), .ZN(n4393) );
  NOR2_X1 U4632 ( .A1(n4394), .A2(n4393), .ZN(n4392) );
  INV_X1 U4633 ( .A(n3909), .ZN(n4500) );
  NOR2_X1 U4634 ( .A1(n3890), .A2(n4500), .ZN(n3891) );
  INV_X1 U4635 ( .A(n3912), .ZN(n4499) );
  AOI22_X1 U4636 ( .A1(REG1_REG_13__SCAN_IN), .A2(n4499), .B1(n3912), .B2(
        n3892), .ZN(n4412) );
  NOR2_X1 U4637 ( .A1(n3893), .A2(n4497), .ZN(n3894) );
  XOR2_X1 U4638 ( .A(n4427), .B(n3893), .Z(n4422) );
  NOR2_X1 U4639 ( .A1(n4849), .A2(n4422), .ZN(n4421) );
  INV_X1 U4640 ( .A(n4440), .ZN(n4496) );
  AOI22_X1 U4641 ( .A1(REG1_REG_15__SCAN_IN), .A2(n4496), .B1(n4440), .B2(
        n4850), .ZN(n4432) );
  NOR2_X1 U4642 ( .A1(n4433), .A2(n4432), .ZN(n4431) );
  NAND2_X1 U4643 ( .A1(n3895), .A2(n4494), .ZN(n3896) );
  NAND2_X1 U4644 ( .A1(n4462), .A2(n4461), .ZN(n4460) );
  OAI21_X1 U4645 ( .B1(n3918), .B2(REG1_REG_17__SCAN_IN), .A(n4460), .ZN(n4470) );
  NOR2_X1 U4646 ( .A1(n4469), .A2(n4470), .ZN(n4471) );
  AOI21_X1 U4647 ( .B1(n3919), .B2(REG1_REG_18__SCAN_IN), .A(n4471), .ZN(n3898) );
  XNOR2_X1 U4648 ( .A(n4555), .B(n4252), .ZN(n3897) );
  XNOR2_X1 U4649 ( .A(n3898), .B(n3897), .ZN(n3928) );
  NAND2_X1 U4650 ( .A1(REG2_REG_18__SCAN_IN), .A2(n3919), .ZN(n3899) );
  OAI21_X1 U4651 ( .B1(REG2_REG_18__SCAN_IN), .B2(n3919), .A(n3899), .ZN(n4480) );
  NOR2_X1 U4652 ( .A1(n3918), .A2(REG2_REG_17__SCAN_IN), .ZN(n3900) );
  AOI21_X1 U4653 ( .B1(REG2_REG_17__SCAN_IN), .B2(n3918), .A(n3900), .ZN(n4459) );
  INV_X1 U4654 ( .A(REG2_REG_13__SCAN_IN), .ZN(n4862) );
  NOR2_X1 U4655 ( .A1(n4862), .A2(n4499), .ZN(n4415) );
  NAND2_X1 U4656 ( .A1(REG2_REG_11__SCAN_IN), .A2(n3901), .ZN(n3908) );
  INV_X1 U4657 ( .A(REG2_REG_11__SCAN_IN), .ZN(n4861) );
  AOI22_X1 U4658 ( .A1(REG2_REG_11__SCAN_IN), .A2(n3901), .B1(n4501), .B2(
        n4861), .ZN(n4399) );
  NAND2_X1 U4659 ( .A1(n3905), .A2(n3906), .ZN(n3907) );
  NAND2_X1 U4660 ( .A1(n3907), .A2(n4388), .ZN(n4398) );
  NAND2_X1 U4661 ( .A1(n3909), .A2(n3910), .ZN(n3911) );
  NAND2_X1 U4662 ( .A1(n3911), .A2(n4407), .ZN(n4417) );
  OAI22_X1 U4663 ( .A1(n4415), .A2(n4417), .B1(REG2_REG_13__SCAN_IN), .B2(
        n3912), .ZN(n3913) );
  NOR2_X1 U4664 ( .A1(n4497), .A2(n3913), .ZN(n3914) );
  INV_X1 U4665 ( .A(REG2_REG_15__SCAN_IN), .ZN(n3915) );
  AOI22_X1 U4666 ( .A1(REG2_REG_15__SCAN_IN), .A2(n4496), .B1(n4440), .B2(
        n3915), .ZN(n4436) );
  NAND2_X1 U4667 ( .A1(n3916), .A2(n4494), .ZN(n3917) );
  INV_X1 U4668 ( .A(REG2_REG_16__SCAN_IN), .ZN(n4717) );
  NAND2_X1 U4669 ( .A1(n4448), .A2(n4717), .ZN(n4447) );
  INV_X1 U4670 ( .A(REG2_REG_19__SCAN_IN), .ZN(n3920) );
  MUX2_X1 U4671 ( .A(n3920), .B(REG2_REG_19__SCAN_IN), .S(n4555), .Z(n3921) );
  XNOR2_X1 U4672 ( .A(n3922), .B(n3921), .ZN(n3926) );
  NAND2_X1 U4673 ( .A1(n4473), .A2(ADDR_REG_19__SCAN_IN), .ZN(n3924) );
  OAI211_X1 U4674 ( .C1(n4485), .C2(n4555), .A(n3924), .B(n3923), .ZN(n3925)
         );
  AOI21_X1 U4675 ( .B1(n3926), .B2(n4482), .A(n3925), .ZN(n3927) );
  OAI21_X1 U4676 ( .B1(n3928), .B2(n4468), .A(n3927), .ZN(U3259) );
  XNOR2_X1 U4677 ( .A(n3932), .B(n3937), .ZN(n4206) );
  INV_X1 U4678 ( .A(n4206), .ZN(n3952) );
  OAI21_X1 U4679 ( .B1(n3935), .B2(n3934), .A(n3933), .ZN(n3936) );
  XOR2_X1 U4680 ( .A(n3937), .B(n3936), .Z(n3944) );
  NAND2_X1 U4681 ( .A1(n3938), .A2(n4187), .ZN(n3942) );
  NAND2_X1 U4682 ( .A1(n4378), .A2(B_REG_SCAN_IN), .ZN(n3939) );
  AND2_X1 U4683 ( .A1(n4289), .A2(n3939), .ZN(n4195) );
  NAND2_X1 U4684 ( .A1(n3940), .A2(n4195), .ZN(n3941) );
  OAI211_X1 U4685 ( .C1(n3946), .C2(n4275), .A(n3942), .B(n3941), .ZN(n3943)
         );
  AOI21_X1 U4686 ( .B1(n3944), .B2(n4162), .A(n3943), .ZN(n4208) );
  OAI21_X1 U4687 ( .B1(n3945), .B2(n4169), .A(n4208), .ZN(n3950) );
  INV_X1 U4688 ( .A(REG2_REG_29__SCAN_IN), .ZN(n3948) );
  OAI22_X1 U4689 ( .A1(n4207), .A2(n4152), .B1(n3948), .B2(n4372), .ZN(n3949)
         );
  AOI21_X1 U4690 ( .B1(n3950), .B2(n4372), .A(n3949), .ZN(n3951) );
  OAI21_X1 U4691 ( .B1(n3952), .B2(n4193), .A(n3951), .ZN(U3354) );
  XOR2_X1 U4692 ( .A(n3960), .B(n3953), .Z(n4216) );
  AOI21_X1 U4693 ( .B1(n3957), .B2(n3977), .A(n3954), .ZN(n4213) );
  INV_X1 U4694 ( .A(n3955), .ZN(n3956) );
  AOI22_X1 U4695 ( .A1(n4142), .A2(REG2_REG_27__SCAN_IN), .B1(n3956), .B2(
        n4568), .ZN(n3959) );
  NAND2_X1 U4696 ( .A1(n4552), .A2(n3957), .ZN(n3958) );
  OAI211_X1 U4697 ( .C1(n4211), .C2(n4559), .A(n3959), .B(n3958), .ZN(n3964)
         );
  XNOR2_X1 U4698 ( .A(n2151), .B(n3960), .ZN(n3962) );
  AOI22_X1 U4699 ( .A1(n3962), .A2(n4162), .B1(n4187), .B2(n3961), .ZN(n4215)
         );
  NOR2_X1 U4700 ( .A1(n4215), .A2(n4142), .ZN(n3963) );
  AOI211_X1 U4701 ( .C1(n4373), .C2(n4213), .A(n3964), .B(n3963), .ZN(n3965)
         );
  OAI21_X1 U4702 ( .B1(n4216), .B2(n4193), .A(n3965), .ZN(U3263) );
  XOR2_X1 U4703 ( .A(n3969), .B(n3966), .Z(n4218) );
  INV_X1 U4704 ( .A(n4218), .ZN(n3984) );
  NAND2_X1 U4705 ( .A1(n3968), .A2(n3967), .ZN(n3970) );
  XNOR2_X1 U4706 ( .A(n3970), .B(n3969), .ZN(n3976) );
  NOR2_X1 U4707 ( .A1(n4275), .A2(n3978), .ZN(n3971) );
  AOI21_X1 U4708 ( .B1(n3972), .B2(n4289), .A(n3971), .ZN(n3975) );
  NAND2_X1 U4709 ( .A1(n3973), .A2(n4187), .ZN(n3974) );
  OAI211_X1 U4710 ( .C1(n3976), .C2(n4553), .A(n3975), .B(n3974), .ZN(n4217)
         );
  OAI21_X1 U4711 ( .B1(n3995), .B2(n3978), .A(n3977), .ZN(n4312) );
  NOR2_X1 U4712 ( .A1(n4312), .A2(n4152), .ZN(n3982) );
  INV_X1 U4713 ( .A(REG2_REG_26__SCAN_IN), .ZN(n3980) );
  OAI22_X1 U4714 ( .A1(n4171), .A2(n3980), .B1(n3979), .B2(n4169), .ZN(n3981)
         );
  AOI211_X1 U4715 ( .C1(n4217), .C2(n4372), .A(n3982), .B(n3981), .ZN(n3983)
         );
  OAI21_X1 U4716 ( .B1(n3984), .B2(n4193), .A(n3983), .ZN(U3264) );
  XNOR2_X1 U4717 ( .A(n3985), .B(n3986), .ZN(n4221) );
  INV_X1 U4718 ( .A(n4221), .ZN(n4001) );
  XNOR2_X1 U4719 ( .A(n3987), .B(n3986), .ZN(n3992) );
  OAI22_X1 U4720 ( .A1(n3988), .A2(n4276), .B1(n4275), .B2(n3993), .ZN(n3989)
         );
  AOI21_X1 U4721 ( .B1(n4187), .B2(n3990), .A(n3989), .ZN(n3991) );
  OAI21_X1 U4722 ( .B1(n3992), .B2(n4553), .A(n3991), .ZN(n4220) );
  NOR2_X1 U4723 ( .A1(n4010), .A2(n3993), .ZN(n3994) );
  INV_X1 U4724 ( .A(n3996), .ZN(n3997) );
  AOI22_X1 U4725 ( .A1(n4142), .A2(REG2_REG_25__SCAN_IN), .B1(n3997), .B2(
        n4568), .ZN(n3998) );
  OAI21_X1 U4726 ( .B1(n4316), .B2(n4152), .A(n3998), .ZN(n3999) );
  AOI21_X1 U4727 ( .B1(n4220), .B2(n4372), .A(n3999), .ZN(n4000) );
  OAI21_X1 U4728 ( .B1(n4001), .B2(n4193), .A(n4000), .ZN(U3265) );
  INV_X1 U4729 ( .A(n4002), .ZN(n4003) );
  XOR2_X1 U4730 ( .A(n4006), .B(n4003), .Z(n4228) );
  INV_X1 U4731 ( .A(n4228), .ZN(n4019) );
  NAND2_X1 U4732 ( .A1(n4005), .A2(n4004), .ZN(n4007) );
  XNOR2_X1 U4733 ( .A(n4007), .B(n4006), .ZN(n4009) );
  OAI22_X1 U4734 ( .A1(n4009), .A2(n4553), .B1(n4008), .B2(n4167), .ZN(n4227)
         );
  INV_X1 U4735 ( .A(n4010), .ZN(n4011) );
  OAI21_X1 U4736 ( .B1(n4040), .B2(n4224), .A(n4011), .ZN(n4320) );
  INV_X1 U4737 ( .A(REG2_REG_24__SCAN_IN), .ZN(n4013) );
  OAI22_X1 U4738 ( .A1(n4171), .A2(n4013), .B1(n4012), .B2(n4169), .ZN(n4015)
         );
  NOR2_X1 U4739 ( .A1(n4559), .A2(n4225), .ZN(n4014) );
  AOI211_X1 U4740 ( .C1(n4552), .C2(n2235), .A(n4015), .B(n4014), .ZN(n4016)
         );
  OAI21_X1 U4741 ( .B1(n4320), .B2(n4152), .A(n4016), .ZN(n4017) );
  AOI21_X1 U4742 ( .B1(n4227), .B2(n4372), .A(n4017), .ZN(n4018) );
  OAI21_X1 U4743 ( .B1(n4019), .B2(n4193), .A(n4018), .ZN(U3266) );
  XNOR2_X1 U4744 ( .A(n4021), .B(n4020), .ZN(n4232) );
  INV_X1 U4745 ( .A(n4232), .ZN(n4047) );
  INV_X1 U4746 ( .A(n4022), .ZN(n4023) );
  INV_X1 U4747 ( .A(n4025), .ZN(n4027) );
  OAI21_X1 U4748 ( .B1(n4080), .B2(n4027), .A(n4026), .ZN(n4066) );
  INV_X1 U4749 ( .A(n4028), .ZN(n4029) );
  AOI21_X1 U4750 ( .B1(n4066), .B2(n4067), .A(n4029), .ZN(n4056) );
  OAI21_X1 U4751 ( .B1(n4056), .B2(n4055), .A(n4030), .ZN(n4032) );
  XNOR2_X1 U4752 ( .A(n4032), .B(n4031), .ZN(n4038) );
  OAI22_X1 U4753 ( .A1(n4034), .A2(n4276), .B1(n4033), .B2(n4275), .ZN(n4035)
         );
  AOI21_X1 U4754 ( .B1(n4187), .B2(n4036), .A(n4035), .ZN(n4037) );
  OAI21_X1 U4755 ( .B1(n4038), .B2(n4553), .A(n4037), .ZN(n4231) );
  AND2_X1 U4756 ( .A1(n2156), .A2(n4039), .ZN(n4041) );
  OR2_X1 U4757 ( .A1(n4041), .A2(n4040), .ZN(n4324) );
  INV_X1 U4758 ( .A(n4042), .ZN(n4043) );
  AOI22_X1 U4759 ( .A1(n4142), .A2(REG2_REG_23__SCAN_IN), .B1(n4043), .B2(
        n4568), .ZN(n4044) );
  OAI21_X1 U4760 ( .B1(n4324), .B2(n4152), .A(n4044), .ZN(n4045) );
  AOI21_X1 U4761 ( .B1(n4231), .B2(n4372), .A(n4045), .ZN(n4046) );
  OAI21_X1 U4762 ( .B1(n4047), .B2(n4193), .A(n4046), .ZN(U3267) );
  OAI21_X1 U4763 ( .B1(n4049), .B2(n4055), .A(n4048), .ZN(n4237) );
  NAND2_X1 U4764 ( .A1(n4069), .A2(n4050), .ZN(n4234) );
  AND2_X1 U4765 ( .A1(n4234), .A2(n4373), .ZN(n4054) );
  INV_X1 U4766 ( .A(REG2_REG_22__SCAN_IN), .ZN(n4052) );
  OAI22_X1 U4767 ( .A1(n4372), .A2(n4052), .B1(n4051), .B2(n4169), .ZN(n4053)
         );
  AOI21_X1 U4768 ( .B1(n4054), .B2(n2156), .A(n4053), .ZN(n4064) );
  XNOR2_X1 U4769 ( .A(n4056), .B(n4055), .ZN(n4062) );
  NAND2_X1 U4770 ( .A1(n4082), .A2(n4187), .ZN(n4059) );
  NAND2_X1 U4771 ( .A1(n4057), .A2(n4289), .ZN(n4058) );
  OAI211_X1 U4772 ( .C1(n4275), .C2(n4060), .A(n4059), .B(n4058), .ZN(n4061)
         );
  AOI21_X1 U4773 ( .B1(n4062), .B2(n4162), .A(n4061), .ZN(n4236) );
  OR2_X1 U4774 ( .A1(n4236), .A2(n4142), .ZN(n4063) );
  OAI211_X1 U4775 ( .C1(n4237), .C2(n4193), .A(n4064), .B(n4063), .ZN(U3268)
         );
  XNOR2_X1 U4776 ( .A(n4065), .B(n4067), .ZN(n4244) );
  XOR2_X1 U4777 ( .A(n4067), .B(n4066), .Z(n4068) );
  OAI22_X1 U4778 ( .A1(n4068), .A2(n4553), .B1(n4111), .B2(n4167), .ZN(n4240)
         );
  INV_X1 U4779 ( .A(n4069), .ZN(n4070) );
  AOI21_X1 U4780 ( .B1(n4074), .B2(n4245), .A(n4070), .ZN(n4242) );
  NAND2_X1 U4781 ( .A1(n4242), .A2(n4373), .ZN(n4076) );
  INV_X1 U4782 ( .A(REG2_REG_21__SCAN_IN), .ZN(n4072) );
  OAI22_X1 U4783 ( .A1(n4171), .A2(n4072), .B1(n4071), .B2(n4169), .ZN(n4073)
         );
  AOI21_X1 U4784 ( .B1(n4074), .B2(n4552), .A(n4073), .ZN(n4075) );
  OAI211_X1 U4785 ( .C1(n4239), .C2(n4559), .A(n4076), .B(n4075), .ZN(n4077)
         );
  AOI21_X1 U4786 ( .B1(n4240), .B2(n4372), .A(n4077), .ZN(n4078) );
  OAI21_X1 U4787 ( .B1(n4244), .B2(n4193), .A(n4078), .ZN(U3269) );
  NAND2_X1 U4788 ( .A1(n4080), .A2(n4079), .ZN(n4081) );
  XNOR2_X1 U4789 ( .A(n4081), .B(n4089), .ZN(n4093) );
  AOI22_X1 U4790 ( .A1(n4082), .A2(n4289), .B1(n4288), .B2(n4095), .ZN(n4083)
         );
  OAI21_X1 U4791 ( .B1(n4084), .B2(n4167), .A(n4083), .ZN(n4092) );
  NAND2_X1 U4792 ( .A1(n4103), .A2(n4085), .ZN(n4088) );
  INV_X1 U4793 ( .A(n4086), .ZN(n4087) );
  NAND2_X1 U4794 ( .A1(n4088), .A2(n4087), .ZN(n4090) );
  XNOR2_X1 U4795 ( .A(n4090), .B(n4089), .ZN(n4249) );
  NOR2_X1 U4796 ( .A1(n4249), .A2(n4554), .ZN(n4091) );
  AOI211_X1 U4797 ( .C1(n4162), .C2(n4093), .A(n4092), .B(n4091), .ZN(n4248)
         );
  INV_X1 U4798 ( .A(n4249), .ZN(n4101) );
  INV_X1 U4799 ( .A(n4094), .ZN(n4116) );
  NAND2_X1 U4800 ( .A1(n4116), .A2(n4095), .ZN(n4246) );
  AND3_X1 U4801 ( .A1(n4246), .A2(n4373), .A3(n4245), .ZN(n4099) );
  INV_X1 U4802 ( .A(REG2_REG_20__SCAN_IN), .ZN(n4097) );
  OAI22_X1 U4803 ( .A1(n4171), .A2(n4097), .B1(n4096), .B2(n4169), .ZN(n4098)
         );
  AOI211_X1 U4804 ( .C1(n4101), .C2(n4100), .A(n4099), .B(n4098), .ZN(n4102)
         );
  OAI21_X1 U4805 ( .B1(n4248), .B2(n4142), .A(n4102), .ZN(U3270) );
  XOR2_X1 U4806 ( .A(n4109), .B(n4103), .Z(n4251) );
  INV_X1 U4807 ( .A(n4251), .ZN(n4122) );
  NAND2_X1 U4808 ( .A1(n4105), .A2(n4104), .ZN(n4123) );
  INV_X1 U4809 ( .A(n4106), .ZN(n4108) );
  OAI21_X1 U4810 ( .B1(n4123), .B2(n4108), .A(n4107), .ZN(n4110) );
  XNOR2_X1 U4811 ( .A(n4110), .B(n4109), .ZN(n4115) );
  OAI22_X1 U4812 ( .A1(n4111), .A2(n4276), .B1(n4275), .B2(n4117), .ZN(n4112)
         );
  AOI21_X1 U4813 ( .B1(n4187), .B2(n4113), .A(n4112), .ZN(n4114) );
  OAI21_X1 U4814 ( .B1(n4115), .B2(n4553), .A(n4114), .ZN(n4250) );
  OAI21_X1 U4815 ( .B1(n2224), .B2(n4117), .A(n4116), .ZN(n4331) );
  NOR2_X1 U4816 ( .A1(n4331), .A2(n4152), .ZN(n4120) );
  OAI22_X1 U4817 ( .A1(n4171), .A2(n3920), .B1(n4118), .B2(n4169), .ZN(n4119)
         );
  AOI211_X1 U4818 ( .C1(n4250), .C2(n4372), .A(n4120), .B(n4119), .ZN(n4121)
         );
  OAI21_X1 U4819 ( .B1(n4122), .B2(n4193), .A(n4121), .ZN(U3271) );
  XNOR2_X1 U4820 ( .A(n4123), .B(n4132), .ZN(n4128) );
  AOI22_X1 U4821 ( .A1(n4125), .A2(n4289), .B1(n4124), .B2(n4288), .ZN(n4126)
         );
  OAI21_X1 U4822 ( .B1(n4261), .B2(n4167), .A(n4126), .ZN(n4127) );
  AOI21_X1 U4823 ( .B1(n4128), .B2(n4162), .A(n4127), .ZN(n4255) );
  INV_X1 U4824 ( .A(n4130), .ZN(n4131) );
  AOI21_X1 U4825 ( .B1(n4132), .B2(n4129), .A(n4131), .ZN(n4256) );
  INV_X1 U4826 ( .A(n4256), .ZN(n4140) );
  OAI211_X1 U4827 ( .C1(n2219), .C2(n4134), .A(n4529), .B(n4133), .ZN(n4254)
         );
  AOI22_X1 U4828 ( .A1(n4142), .A2(REG2_REG_18__SCAN_IN), .B1(n4135), .B2(
        n4568), .ZN(n4136) );
  OAI21_X1 U4829 ( .B1(n4254), .B2(n4137), .A(n4136), .ZN(n4138) );
  AOI21_X1 U4830 ( .B1(n4140), .B2(n4139), .A(n4138), .ZN(n4141) );
  OAI21_X1 U4831 ( .B1(n4142), .B2(n4255), .A(n4141), .ZN(U3272) );
  XOR2_X1 U4832 ( .A(n4145), .B(n4143), .Z(n4258) );
  INV_X1 U4833 ( .A(n4258), .ZN(n4158) );
  XOR2_X1 U4834 ( .A(n4145), .B(n4144), .Z(n4149) );
  OAI22_X1 U4835 ( .A1(n4146), .A2(n4276), .B1(n4151), .B2(n4275), .ZN(n4147)
         );
  AOI21_X1 U4836 ( .B1(n4187), .B2(n4179), .A(n4147), .ZN(n4148) );
  OAI21_X1 U4837 ( .B1(n4149), .B2(n4553), .A(n4148), .ZN(n4257) );
  OAI21_X1 U4838 ( .B1(n4168), .B2(n4151), .A(n4150), .ZN(n4336) );
  NOR2_X1 U4839 ( .A1(n4336), .A2(n4152), .ZN(n4156) );
  INV_X1 U4840 ( .A(REG2_REG_17__SCAN_IN), .ZN(n4154) );
  OAI22_X1 U4841 ( .A1(n4171), .A2(n4154), .B1(n4153), .B2(n4169), .ZN(n4155)
         );
  AOI211_X1 U4842 ( .C1(n4257), .C2(n4372), .A(n4156), .B(n4155), .ZN(n4157)
         );
  OAI21_X1 U4843 ( .B1(n4158), .B2(n4193), .A(n4157), .ZN(U3273) );
  OAI21_X1 U4844 ( .B1(n4161), .B2(n4160), .A(n4159), .ZN(n4266) );
  OAI211_X1 U4845 ( .C1(n4165), .C2(n4164), .A(n4163), .B(n4162), .ZN(n4166)
         );
  OAI21_X1 U4846 ( .B1(n4277), .B2(n4167), .A(n4166), .ZN(n4262) );
  AOI21_X1 U4847 ( .B1(n2223), .B2(n2169), .A(n4168), .ZN(n4264) );
  NAND2_X1 U4848 ( .A1(n4264), .A2(n4373), .ZN(n4174) );
  OAI22_X1 U4849 ( .A1(n4171), .A2(n4717), .B1(n4170), .B2(n4169), .ZN(n4172)
         );
  AOI21_X1 U4850 ( .B1(n2223), .B2(n4552), .A(n4172), .ZN(n4173) );
  OAI211_X1 U4851 ( .C1(n4261), .C2(n4559), .A(n4174), .B(n4173), .ZN(n4175)
         );
  AOI21_X1 U4852 ( .B1(n4262), .B2(n4372), .A(n4175), .ZN(n4176) );
  OAI21_X1 U4853 ( .B1(n4266), .B2(n4193), .A(n4176), .ZN(U3274) );
  XOR2_X1 U4854 ( .A(n4184), .B(n4177), .Z(n4273) );
  XNOR2_X1 U4855 ( .A(n4178), .B(n4267), .ZN(n4270) );
  INV_X1 U4856 ( .A(n4179), .ZN(n4268) );
  AOI22_X1 U4857 ( .A1(n4142), .A2(REG2_REG_15__SCAN_IN), .B1(n4180), .B2(
        n4568), .ZN(n4183) );
  NAND2_X1 U4858 ( .A1(n4552), .A2(n4181), .ZN(n4182) );
  OAI211_X1 U4859 ( .C1(n4268), .C2(n4559), .A(n4183), .B(n4182), .ZN(n4191)
         );
  AOI21_X1 U4860 ( .B1(n4185), .B2(n4184), .A(n4553), .ZN(n4189) );
  AOI22_X1 U4861 ( .A1(n4189), .A2(n4188), .B1(n4187), .B2(n4186), .ZN(n4272)
         );
  NOR2_X1 U4862 ( .A1(n4272), .A2(n4142), .ZN(n4190) );
  AOI211_X1 U4863 ( .C1(n4373), .C2(n4270), .A(n4191), .B(n4190), .ZN(n4192)
         );
  OAI21_X1 U4864 ( .B1(n4273), .B2(n4193), .A(n4192), .ZN(U3275) );
  INV_X1 U4865 ( .A(REG1_REG_31__SCAN_IN), .ZN(n4857) );
  XNOR2_X1 U4866 ( .A(n4200), .B(n4194), .ZN(n4370) );
  NAND2_X1 U4867 ( .A1(n4370), .A2(n4295), .ZN(n4199) );
  NAND2_X1 U4868 ( .A1(n4196), .A2(n4195), .ZN(n4202) );
  OAI21_X1 U4869 ( .B1(n4197), .B2(n4275), .A(n4202), .ZN(n4369) );
  NAND2_X1 U4870 ( .A1(n4369), .A2(n4551), .ZN(n4198) );
  OAI211_X1 U4871 ( .C1(n4551), .C2(n4857), .A(n4199), .B(n4198), .ZN(U3549)
         );
  AOI21_X1 U4872 ( .B1(n4204), .B2(n4201), .A(n4200), .ZN(n4374) );
  INV_X1 U4873 ( .A(n4374), .ZN(n4306) );
  INV_X1 U4874 ( .A(n4202), .ZN(n4203) );
  AOI21_X1 U4875 ( .B1(n4204), .B2(n4288), .A(n4203), .ZN(n4376) );
  MUX2_X1 U4876 ( .A(n2790), .B(n4376), .S(n4551), .Z(n4205) );
  OAI21_X1 U4877 ( .B1(n4306), .B2(n4302), .A(n4205), .ZN(U3548) );
  NAND2_X1 U4878 ( .A1(n4206), .A2(n4527), .ZN(n4209) );
  MUX2_X1 U4879 ( .A(REG1_REG_29__SCAN_IN), .B(n4307), .S(n4551), .Z(U3547) );
  OAI22_X1 U4880 ( .A1(n4211), .A2(n4276), .B1(n4210), .B2(n4275), .ZN(n4212)
         );
  AOI21_X1 U4881 ( .B1(n4213), .B2(n4529), .A(n4212), .ZN(n4214) );
  OAI211_X1 U4882 ( .C1(n4216), .C2(n4522), .A(n4215), .B(n4214), .ZN(n4308)
         );
  MUX2_X1 U4883 ( .A(REG1_REG_27__SCAN_IN), .B(n4308), .S(n4551), .Z(U3545) );
  AOI21_X1 U4884 ( .B1(n4218), .B2(n4527), .A(n4217), .ZN(n4309) );
  MUX2_X1 U4885 ( .A(n4859), .B(n4309), .S(n4551), .Z(n4219) );
  OAI21_X1 U4886 ( .B1(n4302), .B2(n4312), .A(n4219), .ZN(U3544) );
  AOI21_X1 U4887 ( .B1(n4221), .B2(n4527), .A(n4220), .ZN(n4313) );
  MUX2_X1 U4888 ( .A(n4222), .B(n4313), .S(n4551), .Z(n4223) );
  OAI21_X1 U4889 ( .B1(n4302), .B2(n4316), .A(n4223), .ZN(U3543) );
  OAI22_X1 U4890 ( .A1(n4225), .A2(n4276), .B1(n4275), .B2(n4224), .ZN(n4226)
         );
  AOI211_X1 U4891 ( .C1(n4228), .C2(n4527), .A(n4227), .B(n4226), .ZN(n4317)
         );
  MUX2_X1 U4892 ( .A(n4229), .B(n4317), .S(n4551), .Z(n4230) );
  OAI21_X1 U4893 ( .B1(n4302), .B2(n4320), .A(n4230), .ZN(U3542) );
  AOI21_X1 U4894 ( .B1(n4232), .B2(n4527), .A(n4231), .ZN(n4321) );
  MUX2_X1 U4895 ( .A(n4703), .B(n4321), .S(n4551), .Z(n4233) );
  OAI21_X1 U4896 ( .B1(n4302), .B2(n4324), .A(n4233), .ZN(U3541) );
  NAND3_X1 U4897 ( .A1(n2156), .A2(n4529), .A3(n4234), .ZN(n4235) );
  OAI211_X1 U4898 ( .C1(n4237), .C2(n4522), .A(n4236), .B(n4235), .ZN(n4325)
         );
  MUX2_X1 U4899 ( .A(REG1_REG_22__SCAN_IN), .B(n4325), .S(n4551), .Z(U3540) );
  OAI22_X1 U4900 ( .A1(n4239), .A2(n4276), .B1(n4275), .B2(n4238), .ZN(n4241)
         );
  AOI211_X1 U4901 ( .C1(n4529), .C2(n4242), .A(n4241), .B(n4240), .ZN(n4243)
         );
  OAI21_X1 U4902 ( .B1(n4522), .B2(n4244), .A(n4243), .ZN(n4326) );
  MUX2_X1 U4903 ( .A(REG1_REG_21__SCAN_IN), .B(n4326), .S(n4551), .Z(U3539) );
  NAND3_X1 U4904 ( .A1(n4246), .A2(n4529), .A3(n4245), .ZN(n4247) );
  OAI211_X1 U4905 ( .C1(n4249), .C2(n4508), .A(n4248), .B(n4247), .ZN(n4327)
         );
  MUX2_X1 U4906 ( .A(REG1_REG_20__SCAN_IN), .B(n4327), .S(n4551), .Z(U3538) );
  AOI21_X1 U4907 ( .B1(n4251), .B2(n4527), .A(n4250), .ZN(n4328) );
  MUX2_X1 U4908 ( .A(n4252), .B(n4328), .S(n4551), .Z(n4253) );
  OAI21_X1 U4909 ( .B1(n4302), .B2(n4331), .A(n4253), .ZN(U3537) );
  OAI211_X1 U4910 ( .C1(n4256), .C2(n4522), .A(n4255), .B(n4254), .ZN(n4332)
         );
  MUX2_X1 U4911 ( .A(REG1_REG_18__SCAN_IN), .B(n4332), .S(n4551), .Z(U3536) );
  AOI21_X1 U4912 ( .B1(n4258), .B2(n4527), .A(n4257), .ZN(n4333) );
  MUX2_X1 U4913 ( .A(n4858), .B(n4333), .S(n4551), .Z(n4259) );
  OAI21_X1 U4914 ( .B1(n4302), .B2(n4336), .A(n4259), .ZN(U3535) );
  OAI22_X1 U4915 ( .A1(n4261), .A2(n4276), .B1(n4275), .B2(n4260), .ZN(n4263)
         );
  AOI211_X1 U4916 ( .C1(n4529), .C2(n4264), .A(n4263), .B(n4262), .ZN(n4265)
         );
  OAI21_X1 U4917 ( .B1(n4522), .B2(n4266), .A(n4265), .ZN(n4337) );
  MUX2_X1 U4918 ( .A(REG1_REG_16__SCAN_IN), .B(n4337), .S(n4551), .Z(U3534) );
  OAI22_X1 U4919 ( .A1(n4268), .A2(n4276), .B1(n4275), .B2(n4267), .ZN(n4269)
         );
  AOI21_X1 U4920 ( .B1(n4270), .B2(n4529), .A(n4269), .ZN(n4271) );
  OAI211_X1 U4921 ( .C1(n4273), .C2(n4522), .A(n4272), .B(n4271), .ZN(n4338)
         );
  MUX2_X1 U4922 ( .A(REG1_REG_15__SCAN_IN), .B(n4338), .S(n4551), .Z(U3533) );
  OAI22_X1 U4923 ( .A1(n4277), .A2(n4276), .B1(n4275), .B2(n4274), .ZN(n4279)
         );
  AOI211_X1 U4924 ( .C1(n4280), .C2(n4527), .A(n4279), .B(n4278), .ZN(n4339)
         );
  MUX2_X1 U4925 ( .A(n4849), .B(n4339), .S(n4551), .Z(n4281) );
  OAI21_X1 U4926 ( .B1(n4302), .B2(n4341), .A(n4281), .ZN(U3532) );
  NAND2_X1 U4927 ( .A1(n4282), .A2(n4540), .ZN(n4283) );
  OAI211_X1 U4928 ( .C1(n4534), .C2(n4285), .A(n4284), .B(n4283), .ZN(n4342)
         );
  MUX2_X1 U4929 ( .A(REG1_REG_13__SCAN_IN), .B(n4342), .S(n4551), .Z(U3531) );
  NAND2_X1 U4930 ( .A1(n4286), .A2(n4527), .ZN(n4293) );
  AOI22_X1 U4931 ( .A1(n4290), .A2(n4289), .B1(n4288), .B2(n4287), .ZN(n4291)
         );
  NAND3_X1 U4932 ( .A1(n4293), .A2(n4292), .A3(n4291), .ZN(n4343) );
  MUX2_X1 U4933 ( .A(REG1_REG_12__SCAN_IN), .B(n4343), .S(n4551), .Z(n4294) );
  AOI21_X1 U4934 ( .B1(n4295), .B2(n4346), .A(n4294), .ZN(n4296) );
  INV_X1 U4935 ( .A(n4296), .ZN(U3530) );
  INV_X1 U4936 ( .A(n4297), .ZN(n4298) );
  AOI21_X1 U4937 ( .B1(n4540), .B2(n4299), .A(n4298), .ZN(n4348) );
  MUX2_X1 U4938 ( .A(n4300), .B(n4348), .S(n4551), .Z(n4301) );
  OAI21_X1 U4939 ( .B1(n4302), .B2(n4351), .A(n4301), .ZN(U3529) );
  INV_X1 U4940 ( .A(REG0_REG_31__SCAN_IN), .ZN(n4851) );
  NAND2_X1 U4941 ( .A1(n4370), .A2(n4345), .ZN(n4304) );
  NAND2_X1 U4942 ( .A1(n4369), .A2(n4542), .ZN(n4303) );
  OAI211_X1 U4943 ( .C1(n4542), .C2(n4851), .A(n4304), .B(n4303), .ZN(U3517)
         );
  MUX2_X1 U4944 ( .A(n2793), .B(n4376), .S(n4542), .Z(n4305) );
  OAI21_X1 U4945 ( .B1(n4306), .B2(n4350), .A(n4305), .ZN(U3516) );
  MUX2_X1 U4946 ( .A(REG0_REG_29__SCAN_IN), .B(n4307), .S(n4542), .Z(U3515) );
  MUX2_X1 U4947 ( .A(REG0_REG_27__SCAN_IN), .B(n4308), .S(n4542), .Z(U3513) );
  MUX2_X1 U4948 ( .A(n4310), .B(n4309), .S(n4542), .Z(n4311) );
  OAI21_X1 U4949 ( .B1(n4312), .B2(n4350), .A(n4311), .ZN(U3512) );
  MUX2_X1 U4950 ( .A(n4314), .B(n4313), .S(n4542), .Z(n4315) );
  OAI21_X1 U4951 ( .B1(n4316), .B2(n4350), .A(n4315), .ZN(U3511) );
  MUX2_X1 U4952 ( .A(n4318), .B(n4317), .S(n4542), .Z(n4319) );
  OAI21_X1 U4953 ( .B1(n4320), .B2(n4350), .A(n4319), .ZN(U3510) );
  MUX2_X1 U4954 ( .A(n4322), .B(n4321), .S(n4542), .Z(n4323) );
  OAI21_X1 U4955 ( .B1(n4324), .B2(n4350), .A(n4323), .ZN(U3509) );
  MUX2_X1 U4956 ( .A(REG0_REG_22__SCAN_IN), .B(n4325), .S(n4542), .Z(U3508) );
  MUX2_X1 U4957 ( .A(REG0_REG_21__SCAN_IN), .B(n4326), .S(n4542), .Z(U3507) );
  MUX2_X1 U4958 ( .A(REG0_REG_20__SCAN_IN), .B(n4327), .S(n4542), .Z(U3506) );
  MUX2_X1 U4959 ( .A(n4329), .B(n4328), .S(n4542), .Z(n4330) );
  OAI21_X1 U4960 ( .B1(n4331), .B2(n4350), .A(n4330), .ZN(U3505) );
  MUX2_X1 U4961 ( .A(REG0_REG_18__SCAN_IN), .B(n4332), .S(n4542), .Z(U3503) );
  MUX2_X1 U4962 ( .A(n4334), .B(n4333), .S(n4542), .Z(n4335) );
  OAI21_X1 U4963 ( .B1(n4336), .B2(n4350), .A(n4335), .ZN(U3501) );
  MUX2_X1 U4964 ( .A(REG0_REG_16__SCAN_IN), .B(n4337), .S(n4542), .Z(U3499) );
  MUX2_X1 U4965 ( .A(REG0_REG_15__SCAN_IN), .B(n4338), .S(n4542), .Z(U3497) );
  MUX2_X1 U4966 ( .A(n4680), .B(n4339), .S(n4542), .Z(n4340) );
  OAI21_X1 U4967 ( .B1(n4341), .B2(n4350), .A(n4340), .ZN(U3495) );
  MUX2_X1 U4968 ( .A(REG0_REG_13__SCAN_IN), .B(n4342), .S(n4542), .Z(U3493) );
  MUX2_X1 U4969 ( .A(REG0_REG_12__SCAN_IN), .B(n4343), .S(n4542), .Z(n4344) );
  AOI21_X1 U4970 ( .B1(n4346), .B2(n4345), .A(n4344), .ZN(n4347) );
  INV_X1 U4971 ( .A(n4347), .ZN(U3491) );
  MUX2_X1 U4972 ( .A(n4847), .B(n4348), .S(n4542), .Z(n4349) );
  OAI21_X1 U4973 ( .B1(n4351), .B2(n4350), .A(n4349), .ZN(U3489) );
  MUX2_X1 U4974 ( .A(DATAI_29_), .B(n4352), .S(STATE_REG_SCAN_IN), .Z(U3323)
         );
  MUX2_X1 U4975 ( .A(n4378), .B(DATAI_27_), .S(U3149), .Z(U3325) );
  MUX2_X1 U4976 ( .A(n4353), .B(DATAI_26_), .S(U3149), .Z(U3326) );
  MUX2_X1 U4977 ( .A(n4354), .B(DATAI_25_), .S(U3149), .Z(U3327) );
  MUX2_X1 U4978 ( .A(DATAI_24_), .B(n4355), .S(STATE_REG_SCAN_IN), .Z(U3328)
         );
  MUX2_X1 U4979 ( .A(n4356), .B(DATAI_22_), .S(U3149), .Z(U3330) );
  MUX2_X1 U4980 ( .A(n2708), .B(DATAI_21_), .S(U3149), .Z(U3331) );
  MUX2_X1 U4981 ( .A(DATAI_20_), .B(n4357), .S(STATE_REG_SCAN_IN), .Z(U3332)
         );
  MUX2_X1 U4982 ( .A(DATAI_19_), .B(n4358), .S(STATE_REG_SCAN_IN), .Z(U3333)
         );
  MUX2_X1 U4983 ( .A(n4359), .B(DATAI_9_), .S(U3149), .Z(U3343) );
  INV_X1 U4984 ( .A(n4360), .ZN(n4361) );
  MUX2_X1 U4985 ( .A(DATAI_7_), .B(n4361), .S(STATE_REG_SCAN_IN), .Z(U3345) );
  MUX2_X1 U4986 ( .A(n4362), .B(DATAI_6_), .S(U3149), .Z(U3346) );
  MUX2_X1 U4987 ( .A(DATAI_4_), .B(n4363), .S(STATE_REG_SCAN_IN), .Z(U3348) );
  MUX2_X1 U4988 ( .A(n4364), .B(DATAI_3_), .S(U3149), .Z(U3349) );
  MUX2_X1 U4989 ( .A(n4365), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  MUX2_X1 U4990 ( .A(n4366), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  INV_X1 U4991 ( .A(DATAI_28_), .ZN(n4367) );
  AOI22_X1 U4992 ( .A1(STATE_REG_SCAN_IN), .A2(n4368), .B1(n4367), .B2(U3149), 
        .ZN(U3324) );
  INV_X1 U4993 ( .A(REG2_REG_31__SCAN_IN), .ZN(n4792) );
  AOI22_X1 U4994 ( .A1(n4370), .A2(n4373), .B1(n4372), .B2(n4369), .ZN(n4371)
         );
  OAI21_X1 U4995 ( .B1(n4372), .B2(n4792), .A(n4371), .ZN(U3260) );
  AOI22_X1 U4996 ( .A1(n4374), .A2(n4373), .B1(REG2_REG_30__SCAN_IN), .B2(
        n4142), .ZN(n4375) );
  OAI21_X1 U4997 ( .B1(n4142), .B2(n4376), .A(n4375), .ZN(U3261) );
  OAI21_X1 U4998 ( .B1(REG1_REG_0__SCAN_IN), .B2(n4378), .A(n4377), .ZN(n4379)
         );
  XOR2_X1 U4999 ( .A(n4379), .B(IR_REG_0__SCAN_IN), .Z(n4382) );
  AOI22_X1 U5000 ( .A1(ADDR_REG_0__SCAN_IN), .A2(n4473), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n4380) );
  OAI21_X1 U5001 ( .B1(n4382), .B2(n4381), .A(n4380), .ZN(U3240) );
  AOI211_X1 U5002 ( .C1(n2499), .C2(n4384), .A(n4383), .B(n4468), .ZN(n4387)
         );
  INV_X1 U5003 ( .A(n4385), .ZN(n4386) );
  AOI211_X1 U5004 ( .C1(n4473), .C2(ADDR_REG_10__SCAN_IN), .A(n4387), .B(n4386), .ZN(n4391) );
  OAI211_X1 U5005 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4389), .A(n4482), .B(n4388), .ZN(n4390) );
  OAI211_X1 U5006 ( .C1(n4485), .C2(n2299), .A(n4391), .B(n4390), .ZN(U3250)
         );
  AOI211_X1 U5007 ( .C1(n4394), .C2(n4393), .A(n4392), .B(n4468), .ZN(n4396)
         );
  AOI211_X1 U5008 ( .C1(n4473), .C2(ADDR_REG_11__SCAN_IN), .A(n4396), .B(n4395), .ZN(n4401) );
  OAI211_X1 U5009 ( .C1(n4399), .C2(n4398), .A(n4482), .B(n4397), .ZN(n4400)
         );
  OAI211_X1 U5010 ( .C1(n4485), .C2(n4501), .A(n4401), .B(n4400), .ZN(U3251)
         );
  AOI211_X1 U5011 ( .C1(n4692), .C2(n4403), .A(n4402), .B(n4468), .ZN(n4406)
         );
  INV_X1 U5012 ( .A(n4404), .ZN(n4405) );
  AOI211_X1 U5013 ( .C1(n4473), .C2(ADDR_REG_12__SCAN_IN), .A(n4406), .B(n4405), .ZN(n4410) );
  OAI211_X1 U5014 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4408), .A(n4482), .B(n4407), .ZN(n4409) );
  OAI211_X1 U5015 ( .C1(n4485), .C2(n4500), .A(n4410), .B(n4409), .ZN(U3252)
         );
  AOI211_X1 U5016 ( .C1(n2159), .C2(n4412), .A(n4411), .B(n4468), .ZN(n4414)
         );
  AOI211_X1 U5017 ( .C1(n4473), .C2(ADDR_REG_13__SCAN_IN), .A(n4414), .B(n4413), .ZN(n4420) );
  AOI21_X1 U5018 ( .B1(n4862), .B2(n4499), .A(n4415), .ZN(n4418) );
  AOI21_X1 U5019 ( .B1(n4418), .B2(n4417), .A(n4434), .ZN(n4416) );
  OAI21_X1 U5020 ( .B1(n4418), .B2(n4417), .A(n4416), .ZN(n4419) );
  OAI211_X1 U5021 ( .C1(n4485), .C2(n4499), .A(n4420), .B(n4419), .ZN(U3253)
         );
  NAND2_X1 U5022 ( .A1(ADDR_REG_14__SCAN_IN), .A2(n4473), .ZN(n4430) );
  AOI211_X1 U5023 ( .C1(n4849), .C2(n4422), .A(n4421), .B(n4468), .ZN(n4426)
         );
  AOI211_X1 U5024 ( .C1(n3347), .C2(n4424), .A(n4423), .B(n4434), .ZN(n4425)
         );
  AOI211_X1 U5025 ( .C1(n4441), .C2(n4427), .A(n4426), .B(n4425), .ZN(n4429)
         );
  NAND3_X1 U5026 ( .A1(n4430), .A2(n4429), .A3(n4428), .ZN(U3254) );
  INV_X1 U5027 ( .A(n4473), .ZN(n4444) );
  INV_X1 U5028 ( .A(ADDR_REG_15__SCAN_IN), .ZN(n4791) );
  AOI211_X1 U5029 ( .C1(n4433), .C2(n4432), .A(n4431), .B(n4468), .ZN(n4439)
         );
  AOI211_X1 U5030 ( .C1(n4437), .C2(n4436), .A(n4435), .B(n4434), .ZN(n4438)
         );
  AOI211_X1 U5031 ( .C1(n4441), .C2(n4440), .A(n4439), .B(n4438), .ZN(n4443)
         );
  OAI211_X1 U5032 ( .C1(n4444), .C2(n4791), .A(n4443), .B(n4442), .ZN(U3255)
         );
  INV_X1 U5033 ( .A(n4445), .ZN(n4446) );
  AOI21_X1 U5034 ( .B1(n4473), .B2(ADDR_REG_16__SCAN_IN), .A(n4446), .ZN(n4455) );
  OAI21_X1 U5035 ( .B1(n4448), .B2(n4717), .A(n4447), .ZN(n4453) );
  OAI21_X1 U5036 ( .B1(n4451), .B2(n4450), .A(n4449), .ZN(n4452) );
  AOI22_X1 U5037 ( .A1(n4482), .A2(n4453), .B1(n4464), .B2(n4452), .ZN(n4454)
         );
  OAI211_X1 U5038 ( .C1(n4494), .C2(n4485), .A(n4455), .B(n4454), .ZN(U3256)
         );
  AOI21_X1 U5039 ( .B1(n4473), .B2(ADDR_REG_17__SCAN_IN), .A(n4456), .ZN(n4467) );
  OAI21_X1 U5040 ( .B1(n4459), .B2(n4458), .A(n4457), .ZN(n4465) );
  OAI21_X1 U5041 ( .B1(n4462), .B2(n4461), .A(n4460), .ZN(n4463) );
  AOI22_X1 U5042 ( .A1(n4482), .A2(n4465), .B1(n4464), .B2(n4463), .ZN(n4466)
         );
  OAI211_X1 U5043 ( .C1(n4492), .C2(n4485), .A(n4467), .B(n4466), .ZN(U3257)
         );
  AOI21_X1 U5044 ( .B1(n4473), .B2(ADDR_REG_18__SCAN_IN), .A(n4472), .ZN(n4474) );
  INV_X1 U5045 ( .A(n4474), .ZN(n4475) );
  AOI21_X1 U5046 ( .B1(n4480), .B2(n4479), .A(n4478), .ZN(n4481) );
  NAND2_X1 U5047 ( .A1(n4482), .A2(n4481), .ZN(n4483) );
  OAI211_X1 U5048 ( .C1(n4485), .C2(n4490), .A(n4484), .B(n4483), .ZN(U3258)
         );
  AND2_X1 U5049 ( .A1(D_REG_31__SCAN_IN), .A2(n4486), .ZN(U3291) );
  INV_X1 U5050 ( .A(D_REG_30__SCAN_IN), .ZN(n4667) );
  NOR2_X1 U5051 ( .A1(n4487), .A2(n4667), .ZN(U3292) );
  AND2_X1 U5052 ( .A1(D_REG_29__SCAN_IN), .A2(n4486), .ZN(U3293) );
  INV_X1 U5053 ( .A(D_REG_28__SCAN_IN), .ZN(n4663) );
  NOR2_X1 U5054 ( .A1(n4487), .A2(n4663), .ZN(U3294) );
  AND2_X1 U5055 ( .A1(D_REG_27__SCAN_IN), .A2(n4486), .ZN(U3295) );
  AND2_X1 U5056 ( .A1(D_REG_26__SCAN_IN), .A2(n4486), .ZN(U3296) );
  NOR2_X1 U5057 ( .A1(n4487), .A2(n4664), .ZN(U3297) );
  AND2_X1 U5058 ( .A1(D_REG_24__SCAN_IN), .A2(n4486), .ZN(U3298) );
  INV_X1 U5059 ( .A(D_REG_23__SCAN_IN), .ZN(n4656) );
  NOR2_X1 U5060 ( .A1(n4487), .A2(n4656), .ZN(U3299) );
  INV_X1 U5061 ( .A(D_REG_22__SCAN_IN), .ZN(n4657) );
  NOR2_X1 U5062 ( .A1(n4487), .A2(n4657), .ZN(U3300) );
  AND2_X1 U5063 ( .A1(D_REG_21__SCAN_IN), .A2(n4486), .ZN(U3301) );
  INV_X1 U5064 ( .A(D_REG_20__SCAN_IN), .ZN(n4653) );
  NOR2_X1 U5065 ( .A1(n4487), .A2(n4653), .ZN(U3302) );
  AND2_X1 U5066 ( .A1(D_REG_19__SCAN_IN), .A2(n4486), .ZN(U3303) );
  AND2_X1 U5067 ( .A1(D_REG_18__SCAN_IN), .A2(n4486), .ZN(U3304) );
  INV_X1 U5068 ( .A(D_REG_17__SCAN_IN), .ZN(n4654) );
  NOR2_X1 U5069 ( .A1(n4487), .A2(n4654), .ZN(U3305) );
  INV_X1 U5070 ( .A(D_REG_16__SCAN_IN), .ZN(n4651) );
  NOR2_X1 U5071 ( .A1(n4487), .A2(n4651), .ZN(U3306) );
  INV_X1 U5072 ( .A(D_REG_15__SCAN_IN), .ZN(n4803) );
  NOR2_X1 U5073 ( .A1(n4487), .A2(n4803), .ZN(U3307) );
  NOR2_X1 U5074 ( .A1(n4487), .A2(n4648), .ZN(U3308) );
  INV_X1 U5075 ( .A(D_REG_13__SCAN_IN), .ZN(n4649) );
  NOR2_X1 U5076 ( .A1(n4487), .A2(n4649), .ZN(U3309) );
  AND2_X1 U5077 ( .A1(D_REG_12__SCAN_IN), .A2(n4486), .ZN(U3310) );
  NOR2_X1 U5078 ( .A1(n4487), .A2(n4633), .ZN(U3311) );
  AND2_X1 U5079 ( .A1(D_REG_10__SCAN_IN), .A2(n4486), .ZN(U3312) );
  AND2_X1 U5080 ( .A1(D_REG_9__SCAN_IN), .A2(n4486), .ZN(U3313) );
  AND2_X1 U5081 ( .A1(D_REG_8__SCAN_IN), .A2(n4486), .ZN(U3314) );
  NOR2_X1 U5082 ( .A1(n4487), .A2(n4634), .ZN(U3315) );
  AND2_X1 U5083 ( .A1(D_REG_6__SCAN_IN), .A2(n4486), .ZN(U3316) );
  AND2_X1 U5084 ( .A1(D_REG_5__SCAN_IN), .A2(n4486), .ZN(U3317) );
  AND2_X1 U5085 ( .A1(D_REG_4__SCAN_IN), .A2(n4486), .ZN(U3318) );
  NOR2_X1 U5086 ( .A1(n4487), .A2(n4638), .ZN(U3319) );
  NOR2_X1 U5087 ( .A1(n4487), .A2(n4639), .ZN(U3320) );
  INV_X1 U5088 ( .A(DATAI_23_), .ZN(n4489) );
  AOI21_X1 U5089 ( .B1(U3149), .B2(n4489), .A(n4488), .ZN(U3329) );
  AOI22_X1 U5090 ( .A1(STATE_REG_SCAN_IN), .A2(n4490), .B1(n2593), .B2(U3149), 
        .ZN(U3334) );
  INV_X1 U5091 ( .A(DATAI_17_), .ZN(n4491) );
  AOI22_X1 U5092 ( .A1(STATE_REG_SCAN_IN), .A2(n4492), .B1(n4491), .B2(U3149), 
        .ZN(U3335) );
  AOI22_X1 U5093 ( .A1(STATE_REG_SCAN_IN), .A2(n4494), .B1(n4493), .B2(U3149), 
        .ZN(U3336) );
  INV_X1 U5094 ( .A(DATAI_15_), .ZN(n4495) );
  AOI22_X1 U5095 ( .A1(STATE_REG_SCAN_IN), .A2(n4496), .B1(n4495), .B2(U3149), 
        .ZN(U3337) );
  AOI22_X1 U5096 ( .A1(STATE_REG_SCAN_IN), .A2(n4497), .B1(n2547), .B2(U3149), 
        .ZN(U3338) );
  INV_X1 U5097 ( .A(DATAI_13_), .ZN(n4498) );
  AOI22_X1 U5098 ( .A1(STATE_REG_SCAN_IN), .A2(n4499), .B1(n4498), .B2(U3149), 
        .ZN(U3339) );
  INV_X1 U5099 ( .A(DATAI_12_), .ZN(n4839) );
  AOI22_X1 U5100 ( .A1(STATE_REG_SCAN_IN), .A2(n4500), .B1(n4839), .B2(U3149), 
        .ZN(U3340) );
  AOI22_X1 U5101 ( .A1(STATE_REG_SCAN_IN), .A2(n4501), .B1(n2514), .B2(U3149), 
        .ZN(U3341) );
  INV_X1 U5102 ( .A(DATAI_10_), .ZN(n4502) );
  AOI22_X1 U5103 ( .A1(STATE_REG_SCAN_IN), .A2(n2299), .B1(n4502), .B2(U3149), 
        .ZN(U3342) );
  AOI22_X1 U5104 ( .A1(STATE_REG_SCAN_IN), .A2(n2217), .B1(n2218), .B2(U3149), 
        .ZN(U3352) );
  OAI22_X1 U5105 ( .A1(n4505), .A2(n4508), .B1(n4534), .B2(n4504), .ZN(n4506)
         );
  NOR2_X1 U5106 ( .A1(n4507), .A2(n4506), .ZN(n4544) );
  AOI22_X1 U5107 ( .A1(n4542), .A2(n4544), .B1(n4826), .B2(n4541), .ZN(U3469)
         );
  NOR2_X1 U5108 ( .A1(n4509), .A2(n4508), .ZN(n4511) );
  AOI211_X1 U5109 ( .C1(n4529), .C2(n4512), .A(n4511), .B(n4510), .ZN(n4545)
         );
  AOI22_X1 U5110 ( .A1(n4542), .A2(n4545), .B1(n2404), .B2(n4541), .ZN(U3473)
         );
  INV_X1 U5111 ( .A(n4513), .ZN(n4517) );
  INV_X1 U5112 ( .A(n4514), .ZN(n4516) );
  AOI211_X1 U5113 ( .C1(n4517), .C2(n4540), .A(n4516), .B(n4515), .ZN(n4546)
         );
  AOI22_X1 U5114 ( .A1(n4542), .A2(n4546), .B1(n2421), .B2(n4541), .ZN(U3475)
         );
  NOR2_X1 U5115 ( .A1(n4518), .A2(n4534), .ZN(n4520) );
  AOI211_X1 U5116 ( .C1(n4521), .C2(n4527), .A(n4520), .B(n4519), .ZN(n4547)
         );
  AOI22_X1 U5117 ( .A1(n4542), .A2(n4547), .B1(n2436), .B2(n4541), .ZN(U3477)
         );
  NOR2_X1 U5118 ( .A1(n4523), .A2(n4522), .ZN(n4526) );
  AOI211_X1 U5119 ( .C1(n4526), .C2(n3133), .A(n4525), .B(n4524), .ZN(n4548)
         );
  AOI22_X1 U5120 ( .A1(n4542), .A2(n4548), .B1(n2459), .B2(n4541), .ZN(U3481)
         );
  NAND2_X1 U5121 ( .A1(n4528), .A2(n4527), .ZN(n4532) );
  NAND2_X1 U5122 ( .A1(n4530), .A2(n4529), .ZN(n4531) );
  AND3_X1 U5123 ( .A1(n4533), .A2(n4532), .A3(n4531), .ZN(n4549) );
  AOI22_X1 U5124 ( .A1(n4542), .A2(n4549), .B1(n2486), .B2(n4541), .ZN(U3485)
         );
  NOR3_X1 U5125 ( .A1(n4536), .A2(n4535), .A3(n4534), .ZN(n4538) );
  AOI211_X1 U5126 ( .C1(n4540), .C2(n4539), .A(n4538), .B(n4537), .ZN(n4550)
         );
  AOI22_X1 U5127 ( .A1(n4542), .A2(n4550), .B1(n2498), .B2(n4541), .ZN(U3487)
         );
  INV_X1 U5128 ( .A(REG1_REG_1__SCAN_IN), .ZN(n4543) );
  AOI22_X1 U5129 ( .A1(n4551), .A2(n4544), .B1(n4543), .B2(n2751), .ZN(U3519)
         );
  AOI22_X1 U5130 ( .A1(n4551), .A2(n4545), .B1(n2406), .B2(n2751), .ZN(U3521)
         );
  AOI22_X1 U5131 ( .A1(n4551), .A2(n4546), .B1(n2422), .B2(n2751), .ZN(U3522)
         );
  AOI22_X1 U5132 ( .A1(n4551), .A2(n4547), .B1(n2828), .B2(n2751), .ZN(U3523)
         );
  AOI22_X1 U5133 ( .A1(n4551), .A2(n4548), .B1(n2835), .B2(n2751), .ZN(U3525)
         );
  AOI22_X1 U5134 ( .A1(n4551), .A2(n4549), .B1(n2884), .B2(n2751), .ZN(U3527)
         );
  AOI22_X1 U5135 ( .A1(n4551), .A2(n4550), .B1(n2499), .B2(n2751), .ZN(U3528)
         );
  INV_X1 U5136 ( .A(n4552), .ZN(n4562) );
  NAND2_X1 U5137 ( .A1(n4554), .A2(n4553), .ZN(n4557) );
  AOI22_X1 U5138 ( .A1(n4558), .A2(n4557), .B1(n4556), .B2(n4555), .ZN(n4560)
         );
  OAI222_X1 U5139 ( .A1(n4563), .A2(n4562), .B1(n4142), .B2(n4560), .C1(n4559), 
        .C2(n2385), .ZN(n4567) );
  OAI22_X1 U5140 ( .A1(n4565), .A2(n4564), .B1(n4804), .B2(n4372), .ZN(n4566)
         );
  AOI211_X1 U5141 ( .C1(n4568), .C2(REG3_REG_0__SCAN_IN), .A(n4567), .B(n4566), 
        .ZN(n4787) );
  INV_X1 U5142 ( .A(DATAI_26_), .ZN(n4570) );
  AOI22_X1 U5143 ( .A1(n4835), .A2(keyinput61), .B1(n4570), .B2(keyinput87), 
        .ZN(n4569) );
  OAI221_X1 U5144 ( .B1(n4835), .B2(keyinput61), .C1(n4570), .C2(keyinput87), 
        .A(n4569), .ZN(n4579) );
  INV_X1 U5145 ( .A(DATAI_22_), .ZN(n4572) );
  INV_X1 U5146 ( .A(DATAI_21_), .ZN(n4840) );
  AOI22_X1 U5147 ( .A1(n4572), .A2(keyinput44), .B1(keyinput113), .B2(n4840), 
        .ZN(n4571) );
  OAI221_X1 U5148 ( .B1(n4572), .B2(keyinput44), .C1(n4840), .C2(keyinput113), 
        .A(n4571), .ZN(n4578) );
  INV_X1 U5149 ( .A(DATAI_19_), .ZN(n4574) );
  AOI22_X1 U5150 ( .A1(n4574), .A2(keyinput79), .B1(keyinput2), .B2(n2593), 
        .ZN(n4573) );
  OAI221_X1 U5151 ( .B1(n4574), .B2(keyinput79), .C1(n2593), .C2(keyinput2), 
        .A(n4573), .ZN(n4577) );
  AOI22_X1 U5152 ( .A1(n2547), .A2(keyinput23), .B1(keyinput4), .B2(n4839), 
        .ZN(n4575) );
  OAI221_X1 U5153 ( .B1(n2547), .B2(keyinput23), .C1(n4839), .C2(keyinput4), 
        .A(n4575), .ZN(n4576) );
  NOR4_X1 U5154 ( .A1(n4579), .A2(n4578), .A3(n4577), .A4(n4576), .ZN(n4620)
         );
  AOI22_X1 U5155 ( .A1(n4581), .A2(keyinput15), .B1(keyinput109), .B2(n2382), 
        .ZN(n4580) );
  OAI221_X1 U5156 ( .B1(n4581), .B2(keyinput15), .C1(n2382), .C2(keyinput109), 
        .A(n4580), .ZN(n4590) );
  INV_X1 U5157 ( .A(DATAI_9_), .ZN(n4838) );
  AOI22_X1 U5158 ( .A1(n4838), .A2(keyinput86), .B1(keyinput18), .B2(n4583), 
        .ZN(n4582) );
  OAI221_X1 U5159 ( .B1(n4838), .B2(keyinput86), .C1(n4583), .C2(keyinput18), 
        .A(n4582), .ZN(n4589) );
  XNOR2_X1 U5160 ( .A(DATAI_6_), .B(keyinput101), .ZN(n4587) );
  XNOR2_X1 U5161 ( .A(DATAI_4_), .B(keyinput70), .ZN(n4586) );
  XNOR2_X1 U5162 ( .A(DATAI_3_), .B(keyinput63), .ZN(n4585) );
  XNOR2_X1 U5163 ( .A(keyinput43), .B(DATAI_2_), .ZN(n4584) );
  NAND4_X1 U5164 ( .A1(n4587), .A2(n4586), .A3(n4585), .A4(n4584), .ZN(n4588)
         );
  NOR3_X1 U5165 ( .A1(n4590), .A2(n4589), .A3(n4588), .ZN(n4619) );
  AOI22_X1 U5166 ( .A1(n4805), .A2(keyinput36), .B1(n4592), .B2(keyinput92), 
        .ZN(n4591) );
  OAI221_X1 U5167 ( .B1(n4805), .B2(keyinput36), .C1(n4592), .C2(keyinput92), 
        .A(n4591), .ZN(n4604) );
  AOI22_X1 U5168 ( .A1(n4594), .A2(keyinput39), .B1(keyinput41), .B2(n4810), 
        .ZN(n4593) );
  OAI221_X1 U5169 ( .B1(n4594), .B2(keyinput39), .C1(n4810), .C2(keyinput41), 
        .A(n4593), .ZN(n4603) );
  AOI22_X1 U5170 ( .A1(n4597), .A2(keyinput97), .B1(n4596), .B2(keyinput90), 
        .ZN(n4595) );
  OAI221_X1 U5171 ( .B1(n4597), .B2(keyinput97), .C1(n4596), .C2(keyinput90), 
        .A(n4595), .ZN(n4602) );
  AOI22_X1 U5172 ( .A1(n4600), .A2(keyinput96), .B1(keyinput91), .B2(n4599), 
        .ZN(n4598) );
  OAI221_X1 U5173 ( .B1(n4600), .B2(keyinput96), .C1(n4599), .C2(keyinput91), 
        .A(n4598), .ZN(n4601) );
  NOR4_X1 U5174 ( .A1(n4604), .A2(n4603), .A3(n4602), .A4(n4601), .ZN(n4618)
         );
  AOI22_X1 U5175 ( .A1(n4607), .A2(keyinput27), .B1(keyinput62), .B2(n4606), 
        .ZN(n4605) );
  OAI221_X1 U5176 ( .B1(n4607), .B2(keyinput27), .C1(n4606), .C2(keyinput62), 
        .A(n4605), .ZN(n4616) );
  XNOR2_X1 U5177 ( .A(n4608), .B(keyinput51), .ZN(n4615) );
  XNOR2_X1 U5178 ( .A(REG3_REG_0__SCAN_IN), .B(keyinput58), .ZN(n4612) );
  XNOR2_X1 U5179 ( .A(REG3_REG_4__SCAN_IN), .B(keyinput110), .ZN(n4611) );
  XNOR2_X1 U5180 ( .A(IR_REG_12__SCAN_IN), .B(keyinput22), .ZN(n4610) );
  XNOR2_X1 U5181 ( .A(IR_REG_11__SCAN_IN), .B(keyinput94), .ZN(n4609) );
  NAND4_X1 U5182 ( .A1(n4612), .A2(n4611), .A3(n4610), .A4(n4609), .ZN(n4614)
         );
  XNOR2_X1 U5183 ( .A(keyinput16), .B(n2577), .ZN(n4613) );
  NOR4_X1 U5184 ( .A1(n4616), .A2(n4615), .A3(n4614), .A4(n4613), .ZN(n4617)
         );
  NAND4_X1 U5185 ( .A1(n4620), .A2(n4619), .A3(n4618), .A4(n4617), .ZN(n4785)
         );
  INV_X1 U5186 ( .A(IR_REG_29__SCAN_IN), .ZN(n4621) );
  XOR2_X1 U5187 ( .A(n4621), .B(keyinput24), .Z(n4625) );
  XOR2_X1 U5188 ( .A(n2671), .B(keyinput72), .Z(n4624) );
  XOR2_X1 U5189 ( .A(n4815), .B(keyinput30), .Z(n4623) );
  XNOR2_X1 U5190 ( .A(IR_REG_28__SCAN_IN), .B(keyinput34), .ZN(n4622) );
  NAND4_X1 U5191 ( .A1(n4625), .A2(n4624), .A3(n4623), .A4(n4622), .ZN(n4631)
         );
  XNOR2_X1 U5192 ( .A(IR_REG_22__SCAN_IN), .B(keyinput53), .ZN(n4629) );
  XNOR2_X1 U5193 ( .A(IR_REG_18__SCAN_IN), .B(keyinput25), .ZN(n4628) );
  XNOR2_X1 U5194 ( .A(IR_REG_27__SCAN_IN), .B(keyinput52), .ZN(n4627) );
  XNOR2_X1 U5195 ( .A(IR_REG_26__SCAN_IN), .B(keyinput125), .ZN(n4626) );
  NAND4_X1 U5196 ( .A1(n4629), .A2(n4628), .A3(n4627), .A4(n4626), .ZN(n4630)
         );
  NOR2_X1 U5197 ( .A1(n4631), .A2(n4630), .ZN(n4677) );
  AOI22_X1 U5198 ( .A1(n4634), .A2(keyinput99), .B1(keyinput59), .B2(n4633), 
        .ZN(n4632) );
  OAI221_X1 U5199 ( .B1(n4634), .B2(keyinput99), .C1(n4633), .C2(keyinput59), 
        .A(n4632), .ZN(n4646) );
  AOI22_X1 U5200 ( .A1(n4636), .A2(keyinput102), .B1(keyinput56), .B2(n4836), 
        .ZN(n4635) );
  OAI221_X1 U5201 ( .B1(n4636), .B2(keyinput102), .C1(n4836), .C2(keyinput56), 
        .A(n4635), .ZN(n4645) );
  AOI22_X1 U5202 ( .A1(n4639), .A2(keyinput57), .B1(keyinput106), .B2(n4638), 
        .ZN(n4637) );
  OAI221_X1 U5203 ( .B1(n4639), .B2(keyinput57), .C1(n4638), .C2(keyinput106), 
        .A(n4637), .ZN(n4644) );
  XOR2_X1 U5204 ( .A(n4640), .B(keyinput69), .Z(n4642) );
  XNOR2_X1 U5205 ( .A(IR_REG_31__SCAN_IN), .B(keyinput17), .ZN(n4641) );
  NAND2_X1 U5206 ( .A1(n4642), .A2(n4641), .ZN(n4643) );
  NOR4_X1 U5207 ( .A1(n4646), .A2(n4645), .A3(n4644), .A4(n4643), .ZN(n4676)
         );
  AOI22_X1 U5208 ( .A1(n4649), .A2(keyinput1), .B1(keyinput111), .B2(n4648), 
        .ZN(n4647) );
  OAI221_X1 U5209 ( .B1(n4649), .B2(keyinput1), .C1(n4648), .C2(keyinput111), 
        .A(n4647), .ZN(n4661) );
  AOI22_X1 U5210 ( .A1(n4803), .A2(keyinput10), .B1(keyinput6), .B2(n4651), 
        .ZN(n4650) );
  OAI221_X1 U5211 ( .B1(n4803), .B2(keyinput10), .C1(n4651), .C2(keyinput6), 
        .A(n4650), .ZN(n4660) );
  AOI22_X1 U5212 ( .A1(n4654), .A2(keyinput126), .B1(keyinput103), .B2(n4653), 
        .ZN(n4652) );
  OAI221_X1 U5213 ( .B1(n4654), .B2(keyinput126), .C1(n4653), .C2(keyinput103), 
        .A(n4652), .ZN(n4659) );
  AOI22_X1 U5214 ( .A1(n4657), .A2(keyinput93), .B1(keyinput8), .B2(n4656), 
        .ZN(n4655) );
  OAI221_X1 U5215 ( .B1(n4657), .B2(keyinput93), .C1(n4656), .C2(keyinput8), 
        .A(n4655), .ZN(n4658) );
  NOR4_X1 U5216 ( .A1(n4661), .A2(n4660), .A3(n4659), .A4(n4658), .ZN(n4675)
         );
  AOI22_X1 U5217 ( .A1(n4664), .A2(keyinput66), .B1(keyinput78), .B2(n4663), 
        .ZN(n4662) );
  OAI221_X1 U5218 ( .B1(n4664), .B2(keyinput66), .C1(n4663), .C2(keyinput78), 
        .A(n4662), .ZN(n4673) );
  AOI22_X1 U5219 ( .A1(n4667), .A2(keyinput121), .B1(keyinput75), .B2(n4666), 
        .ZN(n4665) );
  OAI221_X1 U5220 ( .B1(n4667), .B2(keyinput121), .C1(n4666), .C2(keyinput75), 
        .A(n4665), .ZN(n4672) );
  AOI22_X1 U5221 ( .A1(n2436), .A2(keyinput5), .B1(keyinput105), .B2(n4826), 
        .ZN(n4668) );
  OAI221_X1 U5222 ( .B1(n2436), .B2(keyinput5), .C1(n4826), .C2(keyinput105), 
        .A(n4668), .ZN(n4671) );
  AOI22_X1 U5223 ( .A1(n2498), .A2(keyinput124), .B1(n4847), .B2(keyinput55), 
        .ZN(n4669) );
  OAI221_X1 U5224 ( .B1(n2498), .B2(keyinput124), .C1(n4847), .C2(keyinput55), 
        .A(n4669), .ZN(n4670) );
  NOR4_X1 U5225 ( .A1(n4673), .A2(n4672), .A3(n4671), .A4(n4670), .ZN(n4674)
         );
  NAND4_X1 U5226 ( .A1(n4677), .A2(n4676), .A3(n4675), .A4(n4674), .ZN(n4784)
         );
  AOI22_X1 U5227 ( .A1(n4680), .A2(keyinput64), .B1(n4679), .B2(keyinput73), 
        .ZN(n4678) );
  OAI221_X1 U5228 ( .B1(n4680), .B2(keyinput64), .C1(n4679), .C2(keyinput73), 
        .A(n4678), .ZN(n4689) );
  AOI22_X1 U5229 ( .A1(n4848), .A2(keyinput108), .B1(n4682), .B2(keyinput77), 
        .ZN(n4681) );
  OAI221_X1 U5230 ( .B1(n4848), .B2(keyinput108), .C1(n4682), .C2(keyinput77), 
        .A(n4681), .ZN(n4688) );
  AOI22_X1 U5231 ( .A1(n4845), .A2(keyinput120), .B1(n4684), .B2(keyinput45), 
        .ZN(n4683) );
  OAI221_X1 U5232 ( .B1(n4845), .B2(keyinput120), .C1(n4684), .C2(keyinput45), 
        .A(n4683), .ZN(n4687) );
  AOI22_X1 U5233 ( .A1(n4846), .A2(keyinput19), .B1(n4852), .B2(keyinput35), 
        .ZN(n4685) );
  OAI221_X1 U5234 ( .B1(n4846), .B2(keyinput19), .C1(n4852), .C2(keyinput35), 
        .A(n4685), .ZN(n4686) );
  NOR4_X1 U5235 ( .A1(n4689), .A2(n4688), .A3(n4687), .A4(n4686), .ZN(n4726)
         );
  AOI22_X1 U5236 ( .A1(n2448), .A2(keyinput84), .B1(keyinput21), .B2(n4851), 
        .ZN(n4690) );
  OAI221_X1 U5237 ( .B1(n2448), .B2(keyinput84), .C1(n4851), .C2(keyinput21), 
        .A(n4690), .ZN(n4699) );
  AOI22_X1 U5238 ( .A1(n4692), .A2(keyinput117), .B1(keyinput9), .B2(n2475), 
        .ZN(n4691) );
  OAI221_X1 U5239 ( .B1(n4692), .B2(keyinput117), .C1(n2475), .C2(keyinput9), 
        .A(n4691), .ZN(n4698) );
  AOI22_X1 U5240 ( .A1(n4850), .A2(keyinput88), .B1(keyinput100), .B2(n4849), 
        .ZN(n4693) );
  OAI221_X1 U5241 ( .B1(n4850), .B2(keyinput88), .C1(n4849), .C2(keyinput100), 
        .A(n4693), .ZN(n4697) );
  AOI22_X1 U5242 ( .A1(n4695), .A2(keyinput107), .B1(n4858), .B2(keyinput114), 
        .ZN(n4694) );
  OAI221_X1 U5243 ( .B1(n4695), .B2(keyinput107), .C1(n4858), .C2(keyinput114), 
        .A(n4694), .ZN(n4696) );
  NOR4_X1 U5244 ( .A1(n4699), .A2(n4698), .A3(n4697), .A4(n4696), .ZN(n4725)
         );
  AOI22_X1 U5245 ( .A1(n4701), .A2(keyinput0), .B1(keyinput83), .B2(n4857), 
        .ZN(n4700) );
  OAI221_X1 U5246 ( .B1(n4701), .B2(keyinput0), .C1(n4857), .C2(keyinput83), 
        .A(n4700), .ZN(n4712) );
  AOI22_X1 U5247 ( .A1(n4704), .A2(keyinput49), .B1(n4703), .B2(keyinput7), 
        .ZN(n4702) );
  OAI221_X1 U5248 ( .B1(n4704), .B2(keyinput49), .C1(n4703), .C2(keyinput7), 
        .A(n4702), .ZN(n4711) );
  AOI22_X1 U5249 ( .A1(n4859), .A2(keyinput89), .B1(n4706), .B2(keyinput98), 
        .ZN(n4705) );
  OAI221_X1 U5250 ( .B1(n4859), .B2(keyinput89), .C1(n4706), .C2(keyinput98), 
        .A(n4705), .ZN(n4710) );
  XOR2_X1 U5251 ( .A(n4804), .B(keyinput119), .Z(n4708) );
  XNOR2_X1 U5252 ( .A(REG2_REG_1__SCAN_IN), .B(keyinput33), .ZN(n4707) );
  NAND2_X1 U5253 ( .A1(n4708), .A2(n4707), .ZN(n4709) );
  NOR4_X1 U5254 ( .A1(n4712), .A2(n4711), .A3(n4710), .A4(n4709), .ZN(n4724)
         );
  INV_X1 U5255 ( .A(REG2_REG_8__SCAN_IN), .ZN(n4714) );
  AOI22_X1 U5256 ( .A1(n4714), .A2(keyinput127), .B1(n3225), .B2(keyinput40), 
        .ZN(n4713) );
  OAI221_X1 U5257 ( .B1(n4714), .B2(keyinput127), .C1(n3225), .C2(keyinput40), 
        .A(n4713), .ZN(n4722) );
  AOI22_X1 U5258 ( .A1(n4862), .A2(keyinput116), .B1(keyinput122), .B2(n4861), 
        .ZN(n4715) );
  OAI221_X1 U5259 ( .B1(n4862), .B2(keyinput116), .C1(n4861), .C2(keyinput122), 
        .A(n4715), .ZN(n4721) );
  AOI22_X1 U5260 ( .A1(n4154), .A2(keyinput118), .B1(keyinput12), .B2(n4717), 
        .ZN(n4716) );
  OAI221_X1 U5261 ( .B1(n4154), .B2(keyinput118), .C1(n4717), .C2(keyinput12), 
        .A(n4716), .ZN(n4720) );
  INV_X1 U5262 ( .A(REG2_REG_18__SCAN_IN), .ZN(n4860) );
  AOI22_X1 U5263 ( .A1(n4860), .A2(keyinput11), .B1(n4072), .B2(keyinput74), 
        .ZN(n4718) );
  OAI221_X1 U5264 ( .B1(n4860), .B2(keyinput11), .C1(n4072), .C2(keyinput74), 
        .A(n4718), .ZN(n4719) );
  NOR4_X1 U5265 ( .A1(n4722), .A2(n4721), .A3(n4720), .A4(n4719), .ZN(n4723)
         );
  NAND4_X1 U5266 ( .A1(n4726), .A2(n4725), .A3(n4724), .A4(n4723), .ZN(n4783)
         );
  AOI22_X1 U5267 ( .A1(n4013), .A2(keyinput123), .B1(n4052), .B2(keyinput85), 
        .ZN(n4727) );
  OAI221_X1 U5268 ( .B1(n4013), .B2(keyinput123), .C1(n4052), .C2(keyinput85), 
        .A(n4727), .ZN(n4736) );
  AOI22_X1 U5269 ( .A1(n3379), .A2(keyinput95), .B1(keyinput32), .B2(n3980), 
        .ZN(n4728) );
  OAI221_X1 U5270 ( .B1(n3379), .B2(keyinput95), .C1(n3980), .C2(keyinput32), 
        .A(n4728), .ZN(n4735) );
  INV_X1 U5271 ( .A(ADDR_REG_16__SCAN_IN), .ZN(n4730) );
  AOI22_X1 U5272 ( .A1(n4792), .A2(keyinput29), .B1(keyinput76), .B2(n4730), 
        .ZN(n4729) );
  OAI221_X1 U5273 ( .B1(n4792), .B2(keyinput29), .C1(n4730), .C2(keyinput76), 
        .A(n4729), .ZN(n4734) );
  INV_X1 U5274 ( .A(ADDR_REG_11__SCAN_IN), .ZN(n4732) );
  AOI22_X1 U5275 ( .A1(n4732), .A2(keyinput82), .B1(n4791), .B2(keyinput115), 
        .ZN(n4731) );
  OAI221_X1 U5276 ( .B1(n4732), .B2(keyinput82), .C1(n4791), .C2(keyinput115), 
        .A(n4731), .ZN(n4733) );
  NOR4_X1 U5277 ( .A1(n4736), .A2(n4735), .A3(n4734), .A4(n4733), .ZN(n4781)
         );
  INV_X1 U5278 ( .A(ADDR_REG_10__SCAN_IN), .ZN(n4739) );
  INV_X1 U5279 ( .A(ADDR_REG_7__SCAN_IN), .ZN(n4738) );
  AOI22_X1 U5280 ( .A1(n4739), .A2(keyinput81), .B1(keyinput20), .B2(n4738), 
        .ZN(n4737) );
  OAI221_X1 U5281 ( .B1(n4739), .B2(keyinput81), .C1(n4738), .C2(keyinput20), 
        .A(n4737), .ZN(n4749) );
  INV_X1 U5282 ( .A(ADDR_REG_2__SCAN_IN), .ZN(n4742) );
  INV_X1 U5283 ( .A(ADDR_REG_3__SCAN_IN), .ZN(n4741) );
  AOI22_X1 U5284 ( .A1(n4742), .A2(keyinput68), .B1(keyinput26), .B2(n4741), 
        .ZN(n4740) );
  OAI221_X1 U5285 ( .B1(n4742), .B2(keyinput68), .C1(n4741), .C2(keyinput26), 
        .A(n4740), .ZN(n4748) );
  AOI22_X1 U5286 ( .A1(n4795), .A2(keyinput13), .B1(keyinput104), .B2(n4744), 
        .ZN(n4743) );
  OAI221_X1 U5287 ( .B1(n4795), .B2(keyinput13), .C1(n4744), .C2(keyinput104), 
        .A(n4743), .ZN(n4747) );
  AOI22_X1 U5288 ( .A1(n4793), .A2(keyinput46), .B1(keyinput37), .B2(n4794), 
        .ZN(n4745) );
  OAI221_X1 U5289 ( .B1(n4793), .B2(keyinput46), .C1(n4794), .C2(keyinput37), 
        .A(n4745), .ZN(n4746) );
  NOR4_X1 U5290 ( .A1(n4749), .A2(n4748), .A3(n4747), .A4(n4746), .ZN(n4780)
         );
  AOI22_X1 U5291 ( .A1(n4751), .A2(keyinput14), .B1(keyinput60), .B2(n4790), 
        .ZN(n4750) );
  OAI221_X1 U5292 ( .B1(n4751), .B2(keyinput14), .C1(n4790), .C2(keyinput60), 
        .A(n4750), .ZN(n4764) );
  AOI22_X1 U5293 ( .A1(n4754), .A2(keyinput80), .B1(keyinput65), .B2(n4753), 
        .ZN(n4752) );
  OAI221_X1 U5294 ( .B1(n4754), .B2(keyinput80), .C1(n4753), .C2(keyinput65), 
        .A(n4752), .ZN(n4763) );
  AOI22_X1 U5295 ( .A1(n4757), .A2(keyinput42), .B1(keyinput71), .B2(n4756), 
        .ZN(n4755) );
  OAI221_X1 U5296 ( .B1(n4757), .B2(keyinput42), .C1(n4756), .C2(keyinput71), 
        .A(n4755), .ZN(n4762) );
  AOI22_X1 U5297 ( .A1(n4760), .A2(keyinput38), .B1(keyinput50), .B2(n4759), 
        .ZN(n4758) );
  OAI221_X1 U5298 ( .B1(n4760), .B2(keyinput38), .C1(n4759), .C2(keyinput50), 
        .A(n4758), .ZN(n4761) );
  NOR4_X1 U5299 ( .A1(n4764), .A2(n4763), .A3(n4762), .A4(n4761), .ZN(n4779)
         );
  AOI22_X1 U5300 ( .A1(n4789), .A2(keyinput112), .B1(keyinput3), .B2(n4766), 
        .ZN(n4765) );
  OAI221_X1 U5301 ( .B1(n4789), .B2(keyinput112), .C1(n4766), .C2(keyinput3), 
        .A(n4765), .ZN(n4777) );
  AOI22_X1 U5302 ( .A1(n4769), .A2(keyinput67), .B1(n4768), .B2(keyinput48), 
        .ZN(n4767) );
  OAI221_X1 U5303 ( .B1(n4769), .B2(keyinput67), .C1(n4768), .C2(keyinput48), 
        .A(n4767), .ZN(n4776) );
  AOI22_X1 U5304 ( .A1(n4822), .A2(keyinput54), .B1(keyinput47), .B2(n4771), 
        .ZN(n4770) );
  OAI221_X1 U5305 ( .B1(n4822), .B2(keyinput54), .C1(n4771), .C2(keyinput47), 
        .A(n4770), .ZN(n4775) );
  XNOR2_X1 U5306 ( .A(REG3_REG_2__SCAN_IN), .B(keyinput28), .ZN(n4773) );
  XNOR2_X1 U5307 ( .A(REG3_REG_19__SCAN_IN), .B(keyinput31), .ZN(n4772) );
  NAND2_X1 U5308 ( .A1(n4773), .A2(n4772), .ZN(n4774) );
  NOR4_X1 U5309 ( .A1(n4777), .A2(n4776), .A3(n4775), .A4(n4774), .ZN(n4778)
         );
  NAND4_X1 U5310 ( .A1(n4781), .A2(n4780), .A3(n4779), .A4(n4778), .ZN(n4782)
         );
  NOR4_X1 U5311 ( .A1(n4785), .A2(n4784), .A3(n4783), .A4(n4782), .ZN(n4786)
         );
  XNOR2_X1 U5312 ( .A(n4787), .B(n4786), .ZN(n4872) );
  INV_X1 U5313 ( .A(n4788), .ZN(n4834) );
  NOR4_X1 U5314 ( .A1(DATAO_REG_17__SCAN_IN), .A2(DATAO_REG_18__SCAN_IN), .A3(
        DATAO_REG_21__SCAN_IN), .A4(n4789), .ZN(n4802) );
  NOR4_X1 U5315 ( .A1(DATAO_REG_15__SCAN_IN), .A2(DATAO_REG_14__SCAN_IN), .A3(
        DATAO_REG_16__SCAN_IN), .A4(n4790), .ZN(n4801) );
  NAND4_X1 U5316 ( .A1(ADDR_REG_16__SCAN_IN), .A2(ADDR_REG_11__SCAN_IN), .A3(
        ADDR_REG_7__SCAN_IN), .A4(n4791), .ZN(n4799) );
  NAND4_X1 U5317 ( .A1(REG2_REG_26__SCAN_IN), .A2(REG2_REG_22__SCAN_IN), .A3(
        n3379), .A4(n4792), .ZN(n4798) );
  NAND4_X1 U5318 ( .A1(DATAO_REG_5__SCAN_IN), .A2(DATAO_REG_10__SCAN_IN), .A3(
        n4794), .A4(n4793), .ZN(n4797) );
  NAND4_X1 U5319 ( .A1(ADDR_REG_2__SCAN_IN), .A2(ADDR_REG_10__SCAN_IN), .A3(
        ADDR_REG_3__SCAN_IN), .A4(n4795), .ZN(n4796) );
  NOR4_X1 U5320 ( .A1(n4799), .A2(n4798), .A3(n4797), .A4(n4796), .ZN(n4800)
         );
  NAND3_X1 U5321 ( .A1(n4802), .A2(n4801), .A3(n4800), .ZN(n4833) );
  NAND4_X1 U5322 ( .A1(D_REG_23__SCAN_IN), .A2(D_REG_11__SCAN_IN), .A3(
        D_REG_20__SCAN_IN), .A4(n4803), .ZN(n4820) );
  NAND4_X1 U5323 ( .A1(REG3_REG_17__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .A3(
        REG0_REG_10__SCAN_IN), .A4(REG0_REG_5__SCAN_IN), .ZN(n4809) );
  NAND4_X1 U5324 ( .A1(REG3_REG_27__SCAN_IN), .A2(REG3_REG_28__SCAN_IN), .A3(
        n4805), .A4(n2382), .ZN(n4808) );
  NAND4_X1 U5325 ( .A1(IR_REG_30__SCAN_IN), .A2(IR_REG_29__SCAN_IN), .A3(
        REG0_REG_0__SCAN_IN), .A4(REG3_REG_0__SCAN_IN), .ZN(n4807) );
  NAND2_X1 U5326 ( .A1(IR_REG_20__SCAN_IN), .A2(n2577), .ZN(n4806) );
  OR4_X1 U5327 ( .A1(n4809), .A2(n4808), .A3(n4807), .A4(n4806), .ZN(n4812) );
  NAND4_X1 U5328 ( .A1(REG3_REG_24__SCAN_IN), .A2(REG3_REG_21__SCAN_IN), .A3(
        REG3_REG_8__SCAN_IN), .A4(n4810), .ZN(n4811) );
  NOR4_X1 U5329 ( .A1(REG3_REG_7__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .A3(
        n4812), .A4(n4811), .ZN(n4813) );
  NAND4_X1 U5330 ( .A1(n2356), .A2(n4815), .A3(n4814), .A4(n4813), .ZN(n4819)
         );
  INV_X1 U5331 ( .A(DATAI_3_), .ZN(n4816) );
  NAND4_X1 U5332 ( .A1(n4816), .A2(D_REG_14__SCAN_IN), .A3(
        DATAO_REG_26__SCAN_IN), .A4(DATAO_REG_30__SCAN_IN), .ZN(n4818) );
  NOR4_X1 U5333 ( .A1(n4820), .A2(n4819), .A3(n4818), .A4(n4817), .ZN(n4831)
         );
  NAND4_X1 U5334 ( .A1(n4822), .A2(IR_REG_28__SCAN_IN), .A3(IR_REG_14__SCAN_IN), .A4(IR_REG_27__SCAN_IN), .ZN(n4823) );
  NOR2_X1 U5335 ( .A1(n4824), .A2(n4823), .ZN(n4830) );
  NOR4_X1 U5336 ( .A1(n4825), .A2(REG3_REG_9__SCAN_IN), .A3(
        REG3_REG_6__SCAN_IN), .A4(REG3_REG_19__SCAN_IN), .ZN(n4829) );
  NOR4_X1 U5337 ( .A1(n4827), .A2(n4826), .A3(REG2_REG_1__SCAN_IN), .A4(
        REG3_REG_2__SCAN_IN), .ZN(n4828) );
  NAND4_X1 U5338 ( .A1(n4831), .A2(n4830), .A3(n4829), .A4(n4828), .ZN(n4832)
         );
  NOR3_X1 U5339 ( .A1(n4834), .A2(n4833), .A3(n4832), .ZN(n4870) );
  NAND4_X1 U5340 ( .A1(DATAI_22_), .A2(DATAI_26_), .A3(n4836), .A4(n4835), 
        .ZN(n4844) );
  NAND4_X1 U5341 ( .A1(D_REG_0__SCAN_IN), .A2(D_REG_16__SCAN_IN), .A3(
        D_REG_28__SCAN_IN), .A4(D_REG_30__SCAN_IN), .ZN(n4843) );
  INV_X1 U5342 ( .A(DATAI_6_), .ZN(n4837) );
  NAND4_X1 U5343 ( .A1(DATAI_7_), .A2(n4839), .A3(n4838), .A4(n4837), .ZN(
        n4842) );
  NAND4_X1 U5344 ( .A1(DATAI_19_), .A2(DATAI_14_), .A3(n4840), .A4(n2593), 
        .ZN(n4841) );
  NOR4_X1 U5345 ( .A1(n4844), .A2(n4843), .A3(n4842), .A4(n4841), .ZN(n4869)
         );
  NAND4_X1 U5346 ( .A1(REG0_REG_27__SCAN_IN), .A2(REG0_REG_21__SCAN_IN), .A3(
        n4846), .A4(n4845), .ZN(n4856) );
  NAND4_X1 U5347 ( .A1(REG0_REG_16__SCAN_IN), .A2(REG0_REG_14__SCAN_IN), .A3(
        n4848), .A4(n4847), .ZN(n4855) );
  NAND4_X1 U5348 ( .A1(REG1_REG_8__SCAN_IN), .A2(REG1_REG_18__SCAN_IN), .A3(
        n4850), .A4(n4849), .ZN(n4854) );
  NAND4_X1 U5349 ( .A1(REG1_REG_12__SCAN_IN), .A2(n4852), .A3(n2448), .A4(
        n4851), .ZN(n4853) );
  NOR4_X1 U5350 ( .A1(n4856), .A2(n4855), .A3(n4854), .A4(n4853), .ZN(n4868)
         );
  NAND4_X1 U5351 ( .A1(REG1_REG_27__SCAN_IN), .A2(REG1_REG_29__SCAN_IN), .A3(
        REG2_REG_8__SCAN_IN), .A4(n4857), .ZN(n4866) );
  NAND4_X1 U5352 ( .A1(REG1_REG_23__SCAN_IN), .A2(REG1_REG_21__SCAN_IN), .A3(
        n4859), .A4(n4858), .ZN(n4865) );
  NAND4_X1 U5353 ( .A1(REG2_REG_16__SCAN_IN), .A2(REG2_REG_21__SCAN_IN), .A3(
        REG2_REG_24__SCAN_IN), .A4(n4860), .ZN(n4864) );
  NAND4_X1 U5354 ( .A1(REG2_REG_10__SCAN_IN), .A2(n4154), .A3(n4862), .A4(
        n4861), .ZN(n4863) );
  NOR4_X1 U5355 ( .A1(n4866), .A2(n4865), .A3(n4864), .A4(n4863), .ZN(n4867)
         );
  NAND4_X1 U5356 ( .A1(n4870), .A2(n4869), .A3(n4868), .A4(n4867), .ZN(n4871)
         );
  XNOR2_X1 U5357 ( .A(n4872), .B(n4871), .ZN(U3290) );
  XNOR2_X1 U2390 ( .A(n3890), .B(n4500), .ZN(n4403) );
  CLKBUF_X1 U2406 ( .A(n3872), .Z(n2134) );
  INV_X2 U2998 ( .A(n4372), .ZN(n4142) );
endmodule

