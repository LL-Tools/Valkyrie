

module b17_C_SARLock_k_128_1 ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, 
        DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, 
        DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, 
        DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, 
        DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, 
        DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, 
        HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN, 
        P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, 
        P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN, 
        P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, 
        P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN, 
        P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN, 
        P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN, 
        P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN, 
        P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN, 
        P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN, 
        P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN, 
        P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN, 
        P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN, 
        P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN, 
        P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN, 
        P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN, 
        P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN, 
        P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN, 
        P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN, 
        P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN, 
        P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN, 
        P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN, 
        P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN, 
        P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN, 
        P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN, 
        P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN, 
        P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN, 
        P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN, 
        P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN, 
        P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN, 
        P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN, 
        P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN, 
        P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN, 
        P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN, 
        P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN, 
        P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN, 
        P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN, 
        P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN, 
        P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, 
        P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, 
        P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, 
        P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, 
        P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, keyinput65, 
        keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, 
        keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, 
        keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, 
        keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, 
        keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, 
        keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, 
        keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, 
        keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, 
        keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, 
        keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, 
        keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, 
        keyinput126, keyinput127, U355, U356, U357, U358, U359, U360, U361, 
        U362, U363, U364, U366, U367, U368, U369, U370, U371, U372, U373, U374, 
        U375, U347, U348, U349, U350, U351, U352, U353, U354, U365, U376, U247, 
        U246, U245, U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, 
        U234, U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223, 
        U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254, U255, 
        U256, U257, U258, U259, U260, U261, U262, U263, U264, U265, U266, U267, 
        U268, U269, U270, U271, U272, U273, U274, U275, U276, U277, U278, U279, 
        U280, U281, U282, U212, U215, U213, U214, P3_U3274, P3_U3275, P3_U3276, 
        P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058, P3_U3057, P3_U3056, 
        P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051, P3_U3050, P3_U3049, 
        P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044, P3_U3043, P3_U3042, 
        P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037, P3_U3036, P3_U3035, 
        P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030, P3_U3029, P3_U3280, 
        P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025, P3_U3024, P3_U3023, 
        P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018, P3_U3017, P3_U3016, 
        P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011, P3_U3010, P3_U3009, 
        P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004, P3_U3003, P3_U3002, 
        P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998, P3_U2997, P3_U2996, 
        P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991, P3_U2990, P3_U2989, 
        P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984, P3_U2983, P3_U2982, 
        P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977, P3_U2976, P3_U2975, 
        P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970, P3_U2969, P3_U2968, 
        P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963, P3_U2962, P3_U2961, 
        P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956, P3_U2955, P3_U2954, 
        P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949, P3_U2948, P3_U2947, 
        P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942, P3_U2941, P3_U2940, 
        P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935, P3_U2934, P3_U2933, 
        P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928, P3_U2927, P3_U2926, 
        P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921, P3_U2920, P3_U2919, 
        P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914, P3_U2913, P3_U2912, 
        P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907, P3_U2906, P3_U2905, 
        P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900, P3_U2899, P3_U2898, 
        P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893, P3_U2892, P3_U2891, 
        P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886, P3_U2885, P3_U2884, 
        P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879, P3_U2878, P3_U2877, 
        P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872, P3_U2871, P3_U2870, 
        P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288, P3_U3289, P3_U3290, 
        P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863, P3_U2862, P3_U2861, 
        P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856, P3_U2855, P3_U2854, 
        P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849, P3_U2848, P3_U2847, 
        P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842, P3_U2841, P3_U2840, 
        P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835, P3_U2834, P3_U2833, 
        P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828, P3_U2827, P3_U2826, 
        P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821, P3_U2820, P3_U2819, 
        P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814, P3_U2813, P3_U2812, 
        P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807, P3_U2806, P3_U2805, 
        P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800, P3_U2799, P3_U2798, 
        P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793, P3_U2792, P3_U2791, 
        P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786, P3_U2785, P3_U2784, 
        P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779, P3_U2778, P3_U2777, 
        P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772, P3_U2771, P3_U2770, 
        P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765, P3_U2764, P3_U2763, 
        P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758, P3_U2757, P3_U2756, 
        P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751, P3_U2750, P3_U2749, 
        P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744, P3_U2743, P3_U2742, 
        P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737, P3_U2736, P3_U2735, 
        P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730, P3_U2729, P3_U2728, 
        P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723, P3_U2722, P3_U2721, 
        P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716, P3_U2715, P3_U2714, 
        P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709, P3_U2708, P3_U2707, 
        P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702, P3_U2701, P3_U2700, 
        P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695, P3_U2694, P3_U2693, 
        P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688, P3_U2687, P3_U2686, 
        P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681, P3_U2680, P3_U2679, 
        P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674, P3_U2673, P3_U2672, 
        P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667, P3_U2666, P3_U2665, 
        P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660, P3_U2659, P3_U2658, 
        P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653, P3_U2652, P3_U2651, 
        P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646, P3_U2645, P3_U2644, 
        P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639, P3_U3292, P3_U2638, 
        P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636, P3_U3296, P3_U2635, 
        P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299, P2_U3585, P2_U3586, 
        P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, 
        P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, 
        P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, 
        P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, 
        P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, 
        P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593, P2_U3178, P2_U3177, 
        P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, P2_U3170, 
        P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, P2_U3163, 
        P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, P2_U3156, 
        P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151, P2_U3150, P2_U3149, 
        P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144, P2_U3143, P2_U3142, 
        P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137, P2_U3136, P2_U3135, 
        P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130, P2_U3129, P2_U3128, 
        P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123, P2_U3122, P2_U3121, 
        P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116, P2_U3115, P2_U3114, 
        P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109, P2_U3108, P2_U3107, 
        P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102, P2_U3101, P2_U3100, 
        P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095, P2_U3094, P2_U3093, 
        P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088, P2_U3087, P2_U3086, 
        P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081, P2_U3080, P2_U3079, 
        P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074, P2_U3073, P2_U3072, 
        P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067, P2_U3066, P2_U3065, 
        P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060, P2_U3059, P2_U3058, 
        P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053, P2_U3052, P2_U3051, 
        P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596, P2_U3599, P2_U3600, 
        P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604, P2_U3605, P2_U3046, 
        P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041, P2_U3040, P2_U3039, 
        P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034, P2_U3033, P2_U3032, 
        P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027, P2_U3026, P2_U3025, 
        P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020, P2_U3019, P2_U3018, 
        P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013, P2_U3012, P2_U3011, 
        P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006, P2_U3005, P2_U3004, 
        P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999, P2_U2998, P2_U2997, 
        P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992, P2_U2991, P2_U2990, 
        P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985, P2_U2984, P2_U2983, 
        P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978, P2_U2977, P2_U2976, 
        P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971, P2_U2970, P2_U2969, 
        P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964, P2_U2963, P2_U2962, 
        P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957, P2_U2956, P2_U2955, 
        P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950, P2_U2949, P2_U2948, 
        P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943, P2_U2942, P2_U2941, 
        P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936, P2_U2935, P2_U2934, 
        P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929, P2_U2928, P2_U2927, 
        P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922, P2_U2921, P2_U2920, 
        P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915, P2_U2914, P2_U2913, 
        P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908, P2_U2907, P2_U2906, 
        P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901, P2_U2900, P2_U2899, 
        P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894, P2_U2893, P2_U2892, 
        P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887, P2_U2886, P2_U2885, 
        P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880, P2_U2879, P2_U2878, 
        P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873, P2_U2872, P2_U2871, 
        P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866, P2_U2865, P2_U2864, 
        P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859, P2_U2858, P2_U2857, 
        P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852, P2_U2851, P2_U2850, 
        P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845, P2_U2844, P2_U2843, 
        P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838, P2_U2837, P2_U2836, 
        P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831, P2_U2830, P2_U2829, 
        P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824, P2_U2823, P2_U2822, 
        P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609, P2_U2818, P2_U3610, 
        P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612, P2_U2814, P1_U3458, 
        P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225, P1_U3224, P1_U3223, 
        P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, 
        P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3210, P1_U3209, 
        P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204, P1_U3203, P1_U3202, 
        P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197, P1_U3196, P1_U3195, 
        P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192, P1_U3191, P1_U3190, 
        P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185, P1_U3184, P1_U3183, 
        P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178, P1_U3177, P1_U3176, 
        P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171, P1_U3170, P1_U3169, 
        P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164, P1_U3466, P1_U3163, 
        P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158, P1_U3157, P1_U3156, 
        P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151, P1_U3150, P1_U3149, 
        P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144, P1_U3143, P1_U3142, 
        P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137, P1_U3136, P1_U3135, 
        P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130, P1_U3129, P1_U3128, 
        P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123, P1_U3122, P1_U3121, 
        P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116, P1_U3115, P1_U3114, 
        P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109, P1_U3108, P1_U3107, 
        P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102, P1_U3101, P1_U3100, 
        P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095, P1_U3094, P1_U3093, 
        P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088, P1_U3087, P1_U3086, 
        P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081, P1_U3080, P1_U3079, 
        P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074, P1_U3073, P1_U3072, 
        P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067, P1_U3066, P1_U3065, 
        P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060, P1_U3059, P1_U3058, 
        P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053, P1_U3052, P1_U3051, 
        P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046, P1_U3045, P1_U3044, 
        P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039, P1_U3038, P1_U3037, 
        P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468, P1_U3469, P1_U3472, 
        P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476, P1_U3477, P1_U3478, 
        P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027, P1_U3026, P1_U3025, 
        P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020, P1_U3019, P1_U3018, 
        P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013, P1_U3012, P1_U3011, 
        P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006, P1_U3005, P1_U3004, 
        P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999, P1_U2998, P1_U2997, 
        P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992, P1_U2991, P1_U2990, 
        P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985, P1_U2984, P1_U2983, 
        P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978, P1_U2977, P1_U2976, 
        P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971, P1_U2970, P1_U2969, 
        P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964, P1_U2963, P1_U2962, 
        P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957, P1_U2956, P1_U2955, 
        P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950, P1_U2949, P1_U2948, 
        P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943, P1_U2942, P1_U2941, 
        P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936, P1_U2935, P1_U2934, 
        P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929, P1_U2928, P1_U2927, 
        P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922, P1_U2921, P1_U2920, 
        P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915, P1_U2914, P1_U2913, 
        P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908, P1_U2907, P1_U2906, 
        P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901, P1_U2900, P1_U2899, 
        P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894, P1_U2893, P1_U2892, 
        P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887, P1_U2886, P1_U2885, 
        P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880, P1_U2879, P1_U2878, 
        P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873, P1_U2872, P1_U2871, 
        P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866, P1_U2865, P1_U2864, 
        P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859, P1_U2858, P1_U2857, 
        P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852, P1_U2851, P1_U2850, 
        P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845, P1_U2844, P1_U2843, 
        P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838, P1_U2837, P1_U2836, 
        P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831, P1_U2830, P1_U2829, 
        P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824, P1_U2823, P1_U2822, 
        P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817, P1_U2816, P1_U2815, 
        P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810, P1_U2809, P1_U2808, 
        P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806, P1_U3484, P1_U2805, 
        P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802, P1_U3487, P1_U2801
 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput0, keyinput1, keyinput2,
         keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8,
         keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779,
         n9781, n9782, n9783, n9784, n9786, n9787, n9788, n9789, n9790, n9791,
         n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801,
         n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811,
         n9812, n9813, n9814, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9988, n9989, n9990, n9991, n9992, n9993,
         n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002,
         n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010,
         n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018,
         n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026,
         n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034,
         n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042,
         n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050,
         n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058,
         n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066,
         n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074,
         n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082,
         n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090,
         n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098,
         n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106,
         n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114,
         n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122,
         n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130,
         n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138,
         n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146,
         n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154,
         n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162,
         n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170,
         n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178,
         n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186,
         n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194,
         n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202,
         n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210,
         n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218,
         n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226,
         n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234,
         n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242,
         n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250,
         n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258,
         n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266,
         n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274,
         n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282,
         n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290,
         n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298,
         n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306,
         n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314,
         n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322,
         n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330,
         n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338,
         n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346,
         n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354,
         n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362,
         n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370,
         n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378,
         n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386,
         n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394,
         n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402,
         n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410,
         n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418,
         n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426,
         n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434,
         n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442,
         n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450,
         n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458,
         n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466,
         n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474,
         n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482,
         n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490,
         n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498,
         n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506,
         n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514,
         n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522,
         n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530,
         n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538,
         n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546,
         n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554,
         n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562,
         n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570,
         n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578,
         n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586,
         n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594,
         n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602,
         n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610,
         n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618,
         n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626,
         n10627, n10628, n10629, n10630, n10631, n10632, n10633, n10634,
         n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642,
         n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650,
         n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658,
         n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666,
         n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674,
         n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682,
         n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690,
         n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698,
         n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10706,
         n10707, n10708, n10709, n10710, n10711, n10712, n10713, n10714,
         n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722,
         n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730,
         n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738,
         n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746,
         n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754,
         n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762,
         n10763, n10764, n10765, n10766, n10767, n10768, n10769, n10770,
         n10771, n10772, n10773, n10774, n10775, n10776, n10777, n10778,
         n10779, n10780, n10781, n10782, n10783, n10784, n10785, n10786,
         n10787, n10788, n10789, n10790, n10791, n10792, n10793, n10794,
         n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802,
         n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810,
         n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818,
         n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826,
         n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834,
         n10835, n10836, n10837, n10838, n10839, n10840, n10841, n10842,
         n10843, n10844, n10845, n10846, n10847, n10848, n10849, n10850,
         n10851, n10852, n10853, n10854, n10855, n10856, n10857, n10858,
         n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866,
         n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10874,
         n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882,
         n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890,
         n10891, n10892, n10893, n10894, n10895, n10896, n10897, n10898,
         n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906,
         n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914,
         n10915, n10916, n10917, n10918, n10919, n10920, n10921, n10922,
         n10923, n10924, n10925, n10926, n10927, n10928, n10929, n10930,
         n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938,
         n10939, n10940, n10941, n10942, n10943, n10944, n10945, n10946,
         n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954,
         n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962,
         n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970,
         n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978,
         n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986,
         n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994,
         n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002,
         n11003, n11004, n11005, n11006, n11007, n11008, n11009, n11010,
         n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018,
         n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026,
         n11027, n11028, n11029, n11030, n11031, n11032, n11033, n11034,
         n11035, n11036, n11037, n11038, n11039, n11040, n11041, n11042,
         n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050,
         n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058,
         n11059, n11060, n11061, n11062, n11063, n11064, n11065, n11066,
         n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074,
         n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082,
         n11083, n11084, n11085, n11086, n11087, n11088, n11089, n11090,
         n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098,
         n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106,
         n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11114,
         n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122,
         n11123, n11124, n11125, n11126, n11127, n11128, n11129, n11130,
         n11131, n11132, n11133, n11134, n11135, n11136, n11137, n11138,
         n11139, n11140, n11141, n11142, n11143, n11144, n11145, n11146,
         n11147, n11148, n11149, n11150, n11151, n11152, n11153, n11154,
         n11155, n11156, n11157, n11158, n11159, n11160, n11161, n11162,
         n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170,
         n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178,
         n11179, n11180, n11181, n11182, n11183, n11184, n11185, n11186,
         n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194,
         n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202,
         n11203, n11204, n11205, n11206, n11207, n11208, n11209, n11210,
         n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218,
         n11219, n11220, n11221, n11222, n11223, n11224, n11225, n11226,
         n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234,
         n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242,
         n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250,
         n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258,
         n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266,
         n11267, n11268, n11269, n11270, n11271, n11272, n11273, n11274,
         n11275, n11276, n11277, n11278, n11279, n11280, n11281, n11282,
         n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11290,
         n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298,
         n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306,
         n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314,
         n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322,
         n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330,
         n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338,
         n11339, n11340, n11341, n11342, n11343, n11344, n11345, n11346,
         n11347, n11348, n11349, n11350, n11351, n11352, n11353, n11354,
         n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362,
         n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370,
         n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378,
         n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386,
         n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394,
         n11395, n11396, n11397, n11398, n11399, n11400, n11401, n11402,
         n11403, n11404, n11405, n11406, n11407, n11408, n11409, n11410,
         n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418,
         n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426,
         n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434,
         n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442,
         n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450,
         n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458,
         n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466,
         n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474,
         n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482,
         n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490,
         n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498,
         n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506,
         n11507, n11508, n11509, n11510, n11511, n11512, n11513, n11514,
         n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522,
         n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530,
         n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538,
         n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546,
         n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554,
         n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562,
         n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570,
         n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578,
         n11579, n11580, n11581, n11582, n11583, n11584, n11585, n11586,
         n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594,
         n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602,
         n11603, n11604, n11605, n11606, n11607, n11608, n11609, n11610,
         n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618,
         n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626,
         n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634,
         n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642,
         n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650,
         n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658,
         n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666,
         n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674,
         n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11682,
         n11683, n11684, n11685, n11686, n11687, n11688, n11689, n11690,
         n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698,
         n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706,
         n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714,
         n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722,
         n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730,
         n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738,
         n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746,
         n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754,
         n11755, n11756, n11757, n11758, n11759, n11760, n11761, n11762,
         n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11770,
         n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11778,
         n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786,
         n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794,
         n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802,
         n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810,
         n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818,
         n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11826,
         n11827, n11828, n11829, n11830, n11831, n11832, n11833, n11834,
         n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11842,
         n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850,
         n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858,
         n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866,
         n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874,
         n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882,
         n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890,
         n11891, n11892, n11893, n11894, n11895, n11896, n11897, n11898,
         n11899, n11900, n11901, n11902, n11903, n11904, n11905, n11906,
         n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914,
         n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922,
         n11923, n11924, n11925, n11926, n11927, n11928, n11929, n11930,
         n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938,
         n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946,
         n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954,
         n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962,
         n11963, n11964, n11965, n11966, n11967, n11968, n11969, n11970,
         n11971, n11972, n11973, n11974, n11975, n11976, n11977, n11978,
         n11979, n11980, n11981, n11982, n11983, n11984, n11985, n11986,
         n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994,
         n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002,
         n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010,
         n12011, n12012, n12013, n12014, n12015, n12016, n12017, n12018,
         n12019, n12020, n12021, n12022, n12023, n12024, n12025, n12026,
         n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034,
         n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042,
         n12043, n12044, n12045, n12046, n12047, n12048, n12049, n12050,
         n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058,
         n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066,
         n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074,
         n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082,
         n12083, n12084, n12085, n12086, n12087, n12088, n12089, n12090,
         n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098,
         n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106,
         n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114,
         n12115, n12116, n12117, n12118, n12119, n12120, n12121, n12122,
         n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130,
         n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138,
         n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12146,
         n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154,
         n12155, n12156, n12157, n12158, n12159, n12160, n12161, n12162,
         n12163, n12164, n12165, n12166, n12167, n12168, n12169, n12170,
         n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178,
         n12179, n12180, n12181, n12182, n12183, n12184, n12185, n12186,
         n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194,
         n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202,
         n12203, n12204, n12205, n12206, n12207, n12208, n12209, n12210,
         n12211, n12212, n12213, n12214, n12215, n12216, n12217, n12218,
         n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226,
         n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234,
         n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242,
         n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250,
         n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258,
         n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266,
         n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274,
         n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282,
         n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290,
         n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298,
         n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306,
         n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314,
         n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12323,
         n12324, n12325, n12326, n12327, n12328, n12329, n12330, n12331,
         n12332, n12333, n12334, n12335, n12336, n12337, n12338, n12339,
         n12340, n12341, n12342, n12343, n12344, n12345, n12346, n12347,
         n12348, n12349, n12350, n12351, n12352, n12353, n12354, n12355,
         n12356, n12357, n12358, n12359, n12360, n12361, n12362, n12363,
         n12364, n12365, n12366, n12367, n12368, n12369, n12370, n12371,
         n12372, n12373, n12374, n12375, n12376, n12377, n12378, n12379,
         n12380, n12381, n12382, n12383, n12384, n12385, n12386, n12387,
         n12388, n12389, n12390, n12391, n12392, n12393, n12394, n12395,
         n12396, n12397, n12398, n12399, n12400, n12401, n12402, n12403,
         n12404, n12405, n12406, n12407, n12408, n12409, n12410, n12411,
         n12412, n12413, n12414, n12415, n12416, n12417, n12418, n12419,
         n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427,
         n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435,
         n12436, n12437, n12438, n12439, n12440, n12441, n12442, n12443,
         n12444, n12445, n12446, n12447, n12448, n12449, n12450, n12451,
         n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459,
         n12460, n12461, n12462, n12463, n12464, n12465, n12466, n12467,
         n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475,
         n12476, n12477, n12478, n12479, n12480, n12481, n12482, n12483,
         n12484, n12485, n12486, n12487, n12488, n12489, n12490, n12491,
         n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499,
         n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507,
         n12508, n12509, n12510, n12511, n12512, n12513, n12514, n12515,
         n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523,
         n12524, n12525, n12526, n12527, n12528, n12529, n12530, n12531,
         n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12539,
         n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547,
         n12548, n12549, n12550, n12551, n12552, n12553, n12554, n12555,
         n12556, n12557, n12558, n12559, n12560, n12561, n12562, n12563,
         n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571,
         n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579,
         n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12587,
         n12588, n12589, n12590, n12591, n12592, n12593, n12594, n12595,
         n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603,
         n12604, n12605, n12606, n12607, n12608, n12609, n12610, n12611,
         n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619,
         n12620, n12621, n12622, n12623, n12624, n12625, n12626, n12627,
         n12628, n12629, n12630, n12631, n12632, n12633, n12634, n12635,
         n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643,
         n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651,
         n12652, n12653, n12654, n12655, n12656, n12657, n12658, n12659,
         n12660, n12661, n12662, n12663, n12664, n12665, n12666, n12667,
         n12668, n12669, n12670, n12671, n12672, n12673, n12674, n12675,
         n12676, n12677, n12678, n12679, n12680, n12681, n12682, n12683,
         n12684, n12685, n12686, n12687, n12688, n12689, n12690, n12691,
         n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699,
         n12700, n12701, n12702, n12703, n12704, n12705, n12706, n12707,
         n12708, n12709, n12710, n12711, n12712, n12713, n12714, n12715,
         n12716, n12717, n12718, n12719, n12720, n12721, n12722, n12723,
         n12724, n12725, n12726, n12727, n12728, n12729, n12730, n12731,
         n12732, n12733, n12734, n12735, n12736, n12737, n12738, n12739,
         n12740, n12741, n12742, n12743, n12744, n12745, n12746, n12747,
         n12748, n12749, n12750, n12751, n12752, n12753, n12754, n12755,
         n12756, n12757, n12758, n12759, n12760, n12761, n12762, n12763,
         n12764, n12765, n12766, n12767, n12768, n12769, n12770, n12771,
         n12772, n12773, n12774, n12775, n12776, n12777, n12778, n12779,
         n12780, n12781, n12782, n12783, n12784, n12785, n12786, n12787,
         n12788, n12789, n12790, n12791, n12792, n12793, n12794, n12795,
         n12796, n12797, n12798, n12799, n12800, n12801, n12802, n12803,
         n12804, n12805, n12806, n12807, n12808, n12809, n12810, n12811,
         n12812, n12813, n12814, n12815, n12816, n12817, n12818, n12819,
         n12820, n12821, n12822, n12823, n12824, n12825, n12826, n12827,
         n12828, n12829, n12830, n12831, n12832, n12833, n12834, n12835,
         n12836, n12837, n12838, n12839, n12840, n12841, n12842, n12843,
         n12844, n12845, n12846, n12847, n12848, n12849, n12850, n12851,
         n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859,
         n12860, n12861, n12862, n12863, n12864, n12865, n12866, n12867,
         n12868, n12869, n12870, n12871, n12872, n12873, n12874, n12875,
         n12876, n12877, n12878, n12879, n12880, n12881, n12882, n12883,
         n12884, n12885, n12886, n12887, n12888, n12889, n12890, n12891,
         n12892, n12893, n12894, n12895, n12896, n12897, n12898, n12899,
         n12900, n12901, n12902, n12903, n12904, n12905, n12906, n12907,
         n12908, n12909, n12910, n12911, n12912, n12913, n12914, n12915,
         n12916, n12917, n12918, n12919, n12920, n12921, n12922, n12923,
         n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931,
         n12932, n12933, n12934, n12935, n12936, n12937, n12938, n12939,
         n12940, n12941, n12942, n12943, n12944, n12945, n12946, n12947,
         n12948, n12949, n12950, n12951, n12952, n12953, n12954, n12955,
         n12956, n12957, n12958, n12959, n12960, n12961, n12962, n12963,
         n12964, n12965, n12966, n12967, n12968, n12969, n12970, n12971,
         n12972, n12973, n12974, n12975, n12976, n12977, n12978, n12979,
         n12980, n12981, n12982, n12983, n12984, n12985, n12986, n12987,
         n12988, n12989, n12990, n12991, n12992, n12993, n12994, n12995,
         n12996, n12997, n12998, n12999, n13000, n13001, n13002, n13003,
         n13004, n13005, n13006, n13007, n13008, n13009, n13010, n13011,
         n13012, n13013, n13014, n13015, n13016, n13017, n13018, n13019,
         n13020, n13021, n13022, n13023, n13024, n13025, n13026, n13027,
         n13028, n13029, n13030, n13031, n13032, n13033, n13034, n13035,
         n13036, n13037, n13038, n13039, n13040, n13041, n13042, n13043,
         n13044, n13045, n13046, n13047, n13048, n13049, n13050, n13051,
         n13052, n13053, n13054, n13055, n13056, n13057, n13058, n13059,
         n13060, n13061, n13062, n13063, n13064, n13065, n13066, n13067,
         n13068, n13069, n13070, n13071, n13072, n13073, n13074, n13075,
         n13076, n13077, n13078, n13079, n13080, n13081, n13082, n13083,
         n13084, n13085, n13086, n13087, n13088, n13089, n13090, n13091,
         n13092, n13093, n13094, n13095, n13096, n13097, n13098, n13099,
         n13100, n13101, n13102, n13103, n13104, n13105, n13106, n13107,
         n13108, n13109, n13110, n13111, n13112, n13113, n13114, n13115,
         n13116, n13117, n13118, n13119, n13120, n13121, n13122, n13123,
         n13124, n13125, n13126, n13127, n13128, n13129, n13130, n13131,
         n13132, n13133, n13134, n13135, n13136, n13137, n13138, n13139,
         n13140, n13141, n13142, n13143, n13144, n13145, n13146, n13147,
         n13148, n13149, n13150, n13151, n13152, n13153, n13154, n13155,
         n13156, n13157, n13158, n13159, n13160, n13161, n13162, n13163,
         n13164, n13165, n13166, n13167, n13168, n13169, n13170, n13171,
         n13172, n13173, n13174, n13175, n13176, n13177, n13178, n13179,
         n13180, n13181, n13182, n13183, n13184, n13185, n13186, n13187,
         n13188, n13189, n13190, n13191, n13192, n13193, n13194, n13195,
         n13196, n13197, n13198, n13199, n13200, n13201, n13202, n13203,
         n13204, n13205, n13206, n13207, n13208, n13209, n13210, n13211,
         n13212, n13213, n13214, n13215, n13216, n13217, n13218, n13219,
         n13220, n13221, n13222, n13223, n13224, n13225, n13226, n13227,
         n13228, n13229, n13230, n13231, n13232, n13233, n13234, n13235,
         n13236, n13237, n13238, n13239, n13240, n13241, n13242, n13243,
         n13244, n13245, n13246, n13247, n13248, n13249, n13250, n13251,
         n13252, n13253, n13254, n13255, n13256, n13257, n13258, n13259,
         n13260, n13261, n13262, n13263, n13264, n13265, n13266, n13267,
         n13268, n13269, n13270, n13271, n13272, n13273, n13274, n13275,
         n13276, n13277, n13278, n13279, n13280, n13281, n13282, n13283,
         n13284, n13285, n13286, n13287, n13288, n13289, n13290, n13291,
         n13292, n13293, n13294, n13295, n13296, n13297, n13298, n13299,
         n13300, n13301, n13302, n13303, n13304, n13305, n13306, n13307,
         n13308, n13309, n13310, n13311, n13312, n13313, n13314, n13315,
         n13316, n13317, n13318, n13319, n13320, n13321, n13322, n13323,
         n13324, n13325, n13326, n13327, n13328, n13329, n13330, n13331,
         n13332, n13333, n13334, n13335, n13336, n13337, n13338, n13339,
         n13340, n13341, n13342, n13343, n13344, n13345, n13346, n13347,
         n13348, n13349, n13350, n13351, n13352, n13353, n13354, n13355,
         n13356, n13357, n13358, n13359, n13360, n13361, n13362, n13363,
         n13364, n13365, n13366, n13367, n13368, n13369, n13370, n13371,
         n13372, n13373, n13374, n13375, n13376, n13377, n13378, n13379,
         n13380, n13381, n13382, n13383, n13384, n13385, n13386, n13387,
         n13388, n13389, n13390, n13391, n13392, n13393, n13394, n13395,
         n13396, n13397, n13398, n13399, n13400, n13401, n13402, n13403,
         n13404, n13405, n13406, n13407, n13408, n13409, n13410, n13411,
         n13412, n13413, n13414, n13415, n13416, n13417, n13418, n13419,
         n13420, n13421, n13422, n13423, n13424, n13425, n13426, n13427,
         n13428, n13429, n13430, n13431, n13432, n13433, n13434, n13435,
         n13436, n13437, n13438, n13439, n13440, n13441, n13442, n13443,
         n13444, n13445, n13446, n13447, n13448, n13449, n13450, n13451,
         n13452, n13453, n13454, n13455, n13456, n13457, n13458, n13459,
         n13460, n13461, n13462, n13463, n13464, n13465, n13466, n13467,
         n13468, n13469, n13470, n13471, n13472, n13473, n13474, n13475,
         n13476, n13477, n13478, n13479, n13480, n13481, n13482, n13483,
         n13484, n13485, n13486, n13487, n13488, n13489, n13490, n13491,
         n13492, n13493, n13494, n13495, n13496, n13497, n13498, n13499,
         n13500, n13501, n13502, n13503, n13504, n13505, n13506, n13507,
         n13508, n13509, n13510, n13511, n13512, n13513, n13514, n13515,
         n13516, n13517, n13518, n13519, n13520, n13521, n13522, n13523,
         n13524, n13525, n13526, n13527, n13528, n13529, n13530, n13531,
         n13532, n13533, n13534, n13535, n13536, n13537, n13538, n13539,
         n13540, n13541, n13542, n13543, n13544, n13545, n13546, n13547,
         n13548, n13549, n13550, n13551, n13552, n13553, n13554, n13555,
         n13556, n13557, n13558, n13559, n13560, n13561, n13562, n13563,
         n13564, n13565, n13566, n13567, n13568, n13569, n13570, n13571,
         n13572, n13573, n13574, n13575, n13576, n13577, n13578, n13579,
         n13580, n13581, n13582, n13583, n13584, n13585, n13586, n13587,
         n13588, n13589, n13591, n13592, n13593, n13594, n13595, n13596,
         n13597, n13598, n13599, n13600, n13601, n13602, n13603, n13604,
         n13605, n13606, n13607, n13608, n13609, n13610, n13611, n13612,
         n13613, n13614, n13615, n13616, n13617, n13618, n13619, n13620,
         n13621, n13622, n13623, n13624, n13625, n13626, n13627, n13628,
         n13629, n13630, n13631, n13632, n13633, n13634, n13635, n13636,
         n13637, n13638, n13639, n13640, n13641, n13642, n13643, n13644,
         n13645, n13646, n13647, n13648, n13649, n13650, n13651, n13652,
         n13653, n13654, n13655, n13656, n13657, n13658, n13659, n13660,
         n13661, n13662, n13663, n13664, n13665, n13666, n13667, n13668,
         n13669, n13670, n13671, n13672, n13673, n13674, n13675, n13676,
         n13677, n13678, n13679, n13680, n13681, n13682, n13683, n13684,
         n13685, n13686, n13687, n13688, n13689, n13690, n13691, n13692,
         n13693, n13694, n13695, n13696, n13697, n13698, n13699, n13700,
         n13701, n13702, n13703, n13704, n13705, n13706, n13707, n13708,
         n13709, n13710, n13711, n13712, n13713, n13714, n13715, n13716,
         n13717, n13718, n13719, n13720, n13721, n13722, n13723, n13724,
         n13725, n13726, n13727, n13728, n13729, n13730, n13731, n13732,
         n13733, n13734, n13735, n13736, n13737, n13738, n13739, n13740,
         n13741, n13742, n13743, n13744, n13745, n13746, n13747, n13748,
         n13749, n13750, n13751, n13752, n13753, n13754, n13755, n13756,
         n13757, n13758, n13759, n13760, n13761, n13762, n13763, n13764,
         n13765, n13766, n13767, n13768, n13769, n13770, n13771, n13772,
         n13773, n13774, n13775, n13776, n13777, n13778, n13779, n13780,
         n13781, n13782, n13783, n13784, n13785, n13786, n13787, n13788,
         n13789, n13790, n13791, n13792, n13793, n13794, n13795, n13796,
         n13797, n13798, n13799, n13800, n13801, n13802, n13803, n13804,
         n13805, n13806, n13807, n13808, n13809, n13810, n13811, n13812,
         n13813, n13814, n13815, n13816, n13817, n13818, n13819, n13820,
         n13821, n13822, n13823, n13824, n13825, n13826, n13827, n13828,
         n13829, n13830, n13831, n13832, n13833, n13834, n13835, n13836,
         n13837, n13838, n13839, n13840, n13841, n13842, n13843, n13844,
         n13845, n13846, n13847, n13848, n13849, n13850, n13851, n13852,
         n13853, n13854, n13855, n13856, n13857, n13858, n13859, n13860,
         n13861, n13862, n13863, n13864, n13865, n13866, n13867, n13868,
         n13869, n13870, n13871, n13872, n13873, n13874, n13875, n13876,
         n13877, n13878, n13879, n13880, n13881, n13882, n13883, n13884,
         n13885, n13886, n13887, n13888, n13889, n13890, n13891, n13892,
         n13893, n13894, n13895, n13896, n13897, n13898, n13899, n13900,
         n13901, n13902, n13903, n13904, n13905, n13906, n13907, n13908,
         n13909, n13910, n13911, n13912, n13913, n13914, n13915, n13916,
         n13917, n13918, n13919, n13920, n13921, n13922, n13923, n13924,
         n13925, n13926, n13927, n13928, n13929, n13930, n13931, n13932,
         n13933, n13934, n13935, n13936, n13937, n13938, n13939, n13940,
         n13941, n13942, n13943, n13944, n13945, n13946, n13947, n13948,
         n13949, n13950, n13951, n13952, n13953, n13954, n13955, n13956,
         n13957, n13958, n13959, n13960, n13961, n13962, n13963, n13964,
         n13965, n13966, n13967, n13968, n13969, n13970, n13971, n13972,
         n13973, n13974, n13975, n13976, n13977, n13978, n13979, n13980,
         n13981, n13982, n13983, n13984, n13985, n13986, n13987, n13988,
         n13989, n13990, n13991, n13992, n13993, n13994, n13995, n13996,
         n13997, n13998, n13999, n14000, n14001, n14002, n14003, n14004,
         n14005, n14006, n14007, n14008, n14009, n14010, n14011, n14012,
         n14013, n14014, n14015, n14016, n14017, n14018, n14019, n14020,
         n14021, n14022, n14023, n14024, n14025, n14026, n14027, n14028,
         n14029, n14030, n14031, n14032, n14033, n14034, n14035, n14036,
         n14037, n14038, n14039, n14040, n14041, n14042, n14043, n14044,
         n14045, n14046, n14047, n14048, n14049, n14050, n14051, n14052,
         n14053, n14054, n14055, n14056, n14057, n14058, n14059, n14060,
         n14061, n14062, n14063, n14064, n14065, n14066, n14067, n14068,
         n14069, n14070, n14071, n14072, n14073, n14074, n14075, n14076,
         n14077, n14078, n14079, n14080, n14081, n14082, n14083, n14084,
         n14085, n14086, n14087, n14088, n14089, n14090, n14091, n14092,
         n14093, n14094, n14095, n14096, n14097, n14098, n14099, n14100,
         n14101, n14102, n14103, n14104, n14105, n14106, n14107, n14108,
         n14109, n14110, n14111, n14112, n14113, n14114, n14115, n14116,
         n14117, n14118, n14119, n14120, n14121, n14122, n14123, n14124,
         n14125, n14126, n14127, n14128, n14129, n14130, n14131, n14132,
         n14133, n14134, n14135, n14136, n14137, n14138, n14139, n14140,
         n14141, n14142, n14143, n14144, n14145, n14146, n14147, n14148,
         n14149, n14150, n14151, n14152, n14153, n14154, n14155, n14156,
         n14157, n14158, n14159, n14160, n14161, n14162, n14163, n14164,
         n14165, n14166, n14167, n14168, n14169, n14170, n14171, n14172,
         n14173, n14174, n14175, n14176, n14177, n14178, n14179, n14180,
         n14181, n14182, n14183, n14184, n14185, n14186, n14187, n14188,
         n14189, n14190, n14191, n14192, n14193, n14194, n14195, n14196,
         n14197, n14198, n14199, n14200, n14201, n14202, n14203, n14204,
         n14205, n14206, n14207, n14208, n14209, n14210, n14211, n14212,
         n14213, n14214, n14215, n14216, n14217, n14218, n14219, n14220,
         n14221, n14222, n14223, n14224, n14225, n14226, n14227, n14228,
         n14229, n14230, n14231, n14232, n14233, n14234, n14235, n14236,
         n14237, n14238, n14239, n14240, n14241, n14242, n14243, n14244,
         n14245, n14246, n14247, n14248, n14249, n14250, n14251, n14252,
         n14253, n14254, n14255, n14256, n14257, n14258, n14259, n14260,
         n14261, n14262, n14263, n14264, n14265, n14266, n14267, n14268,
         n14269, n14270, n14271, n14272, n14273, n14274, n14275, n14276,
         n14277, n14278, n14279, n14280, n14281, n14282, n14283, n14284,
         n14285, n14286, n14287, n14288, n14289, n14290, n14291, n14292,
         n14293, n14294, n14295, n14296, n14297, n14298, n14299, n14300,
         n14301, n14302, n14303, n14304, n14305, n14306, n14307, n14308,
         n14309, n14310, n14311, n14312, n14313, n14314, n14315, n14316,
         n14317, n14318, n14319, n14320, n14321, n14322, n14323, n14324,
         n14325, n14326, n14327, n14328, n14329, n14330, n14331, n14332,
         n14333, n14334, n14335, n14336, n14337, n14338, n14339, n14340,
         n14341, n14342, n14343, n14344, n14345, n14346, n14347, n14348,
         n14349, n14350, n14351, n14352, n14353, n14354, n14355, n14356,
         n14357, n14358, n14359, n14360, n14361, n14362, n14363, n14364,
         n14365, n14366, n14367, n14368, n14369, n14370, n14371, n14372,
         n14373, n14374, n14375, n14376, n14377, n14378, n14379, n14380,
         n14381, n14382, n14383, n14384, n14385, n14386, n14387, n14388,
         n14389, n14390, n14391, n14392, n14393, n14394, n14395, n14396,
         n14397, n14398, n14399, n14400, n14401, n14402, n14403, n14404,
         n14405, n14406, n14407, n14408, n14409, n14410, n14411, n14412,
         n14413, n14414, n14415, n14416, n14417, n14418, n14419, n14420,
         n14421, n14422, n14423, n14424, n14425, n14426, n14427, n14428,
         n14429, n14430, n14431, n14432, n14433, n14434, n14435, n14436,
         n14437, n14438, n14439, n14440, n14441, n14442, n14443, n14444,
         n14445, n14446, n14447, n14448, n14449, n14450, n14451, n14452,
         n14453, n14454, n14455, n14456, n14457, n14458, n14459, n14460,
         n14461, n14462, n14463, n14464, n14465, n14466, n14467, n14468,
         n14469, n14470, n14471, n14472, n14473, n14474, n14475, n14476,
         n14477, n14478, n14479, n14480, n14481, n14482, n14483, n14484,
         n14485, n14486, n14487, n14488, n14489, n14490, n14491, n14492,
         n14493, n14494, n14495, n14496, n14497, n14498, n14499, n14500,
         n14501, n14502, n14503, n14504, n14505, n14506, n14507, n14508,
         n14509, n14510, n14511, n14512, n14513, n14514, n14515, n14516,
         n14517, n14518, n14519, n14520, n14521, n14522, n14523, n14524,
         n14525, n14526, n14527, n14528, n14529, n14530, n14531, n14532,
         n14533, n14534, n14535, n14536, n14537, n14538, n14539, n14540,
         n14541, n14542, n14543, n14544, n14545, n14546, n14547, n14548,
         n14549, n14550, n14551, n14552, n14553, n14554, n14555, n14556,
         n14557, n14558, n14559, n14560, n14561, n14562, n14563, n14564,
         n14565, n14566, n14567, n14568, n14569, n14570, n14571, n14572,
         n14573, n14574, n14575, n14576, n14577, n14578, n14579, n14580,
         n14581, n14582, n14583, n14584, n14585, n14586, n14587, n14588,
         n14589, n14590, n14591, n14592, n14593, n14594, n14595, n14596,
         n14597, n14598, n14599, n14600, n14601, n14602, n14603, n14604,
         n14605, n14606, n14607, n14608, n14609, n14610, n14611, n14612,
         n14613, n14614, n14615, n14616, n14617, n14618, n14619, n14620,
         n14621, n14622, n14623, n14624, n14625, n14626, n14627, n14628,
         n14629, n14630, n14631, n14632, n14633, n14634, n14635, n14636,
         n14637, n14638, n14639, n14640, n14641, n14642, n14643, n14644,
         n14645, n14646, n14647, n14648, n14649, n14650, n14651, n14652,
         n14653, n14654, n14655, n14656, n14657, n14658, n14659, n14660,
         n14661, n14662, n14663, n14664, n14665, n14666, n14667, n14668,
         n14669, n14670, n14671, n14672, n14673, n14674, n14675, n14676,
         n14677, n14678, n14679, n14680, n14681, n14682, n14683, n14684,
         n14685, n14686, n14687, n14688, n14689, n14690, n14691, n14692,
         n14693, n14694, n14695, n14696, n14697, n14698, n14699, n14700,
         n14701, n14702, n14703, n14704, n14705, n14706, n14707, n14708,
         n14709, n14710, n14711, n14712, n14713, n14714, n14715, n14716,
         n14717, n14718, n14719, n14720, n14721, n14722, n14723, n14724,
         n14725, n14726, n14727, n14728, n14729, n14730, n14731, n14732,
         n14733, n14734, n14735, n14736, n14737, n14738, n14739, n14740,
         n14741, n14742, n14743, n14744, n14745, n14746, n14747, n14748,
         n14749, n14750, n14751, n14752, n14753, n14754, n14755, n14756,
         n14757, n14758, n14759, n14760, n14761, n14762, n14763, n14764,
         n14765, n14766, n14767, n14768, n14769, n14770, n14771, n14772,
         n14773, n14774, n14775, n14776, n14777, n14778, n14779, n14780,
         n14781, n14782, n14783, n14784, n14785, n14786, n14787, n14788,
         n14789, n14790, n14791, n14792, n14793, n14794, n14795, n14796,
         n14797, n14798, n14799, n14800, n14801, n14802, n14803, n14804,
         n14805, n14806, n14807, n14808, n14809, n14810, n14811, n14812,
         n14813, n14814, n14815, n14816, n14817, n14818, n14819, n14820,
         n14821, n14822, n14823, n14824, n14825, n14826, n14827, n14828,
         n14829, n14830, n14831, n14832, n14833, n14834, n14835, n14836,
         n14837, n14838, n14839, n14840, n14841, n14842, n14843, n14844,
         n14845, n14846, n14847, n14848, n14849, n14850, n14851, n14852,
         n14853, n14854, n14855, n14856, n14857, n14858, n14859, n14860,
         n14861, n14862, n14863, n14864, n14865, n14866, n14867, n14868,
         n14869, n14870, n14871, n14872, n14873, n14874, n14875, n14876,
         n14877, n14878, n14879, n14880, n14881, n14882, n14883, n14884,
         n14885, n14886, n14887, n14888, n14889, n14890, n14891, n14892,
         n14893, n14894, n14895, n14896, n14897, n14898, n14899, n14900,
         n14901, n14902, n14903, n14904, n14905, n14906, n14907, n14908,
         n14909, n14910, n14911, n14912, n14913, n14914, n14915, n14916,
         n14917, n14918, n14919, n14920, n14921, n14922, n14923, n14924,
         n14925, n14926, n14927, n14928, n14929, n14930, n14931, n14932,
         n14933, n14934, n14935, n14936, n14937, n14938, n14939, n14940,
         n14941, n14942, n14943, n14944, n14945, n14946, n14947, n14948,
         n14949, n14950, n14951, n14952, n14953, n14954, n14955, n14956,
         n14957, n14958, n14959, n14960, n14961, n14962, n14963, n14964,
         n14965, n14966, n14967, n14968, n14969, n14970, n14971, n14972,
         n14973, n14974, n14975, n14976, n14977, n14978, n14979, n14980,
         n14981, n14982, n14983, n14984, n14985, n14986, n14987, n14988,
         n14989, n14990, n14991, n14992, n14993, n14994, n14995, n14996,
         n14997, n14998, n14999, n15000, n15001, n15002, n15003, n15004,
         n15005, n15006, n15007, n15008, n15009, n15010, n15011, n15012,
         n15013, n15014, n15015, n15016, n15017, n15018, n15019, n15020,
         n15021, n15022, n15023, n15024, n15025, n15026, n15027, n15028,
         n15029, n15030, n15031, n15032, n15033, n15034, n15035, n15036,
         n15037, n15038, n15039, n15040, n15041, n15042, n15043, n15044,
         n15045, n15046, n15047, n15048, n15049, n15050, n15051, n15052,
         n15053, n15054, n15055, n15056, n15057, n15058, n15059, n15060,
         n15061, n15062, n15063, n15064, n15065, n15066, n15067, n15068,
         n15069, n15070, n15071, n15072, n15073, n15074, n15075, n15076,
         n15077, n15078, n15079, n15080, n15081, n15082, n15083, n15084,
         n15085, n15086, n15087, n15088, n15089, n15090, n15091, n15092,
         n15093, n15094, n15095, n15096, n15097, n15098, n15099, n15100,
         n15101, n15102, n15103, n15104, n15105, n15106, n15107, n15108,
         n15109, n15110, n15111, n15112, n15113, n15114, n15115, n15116,
         n15117, n15118, n15119, n15120, n15121, n15122, n15123, n15124,
         n15125, n15126, n15127, n15128, n15129, n15130, n15131, n15132,
         n15133, n15134, n15135, n15136, n15137, n15138, n15139, n15140,
         n15141, n15142, n15143, n15144, n15145, n15146, n15147, n15148,
         n15149, n15150, n15151, n15152, n15153, n15154, n15155, n15156,
         n15157, n15158, n15159, n15160, n15161, n15162, n15163, n15164,
         n15165, n15166, n15167, n15168, n15169, n15170, n15171, n15172,
         n15173, n15174, n15175, n15176, n15177, n15178, n15179, n15180,
         n15181, n15182, n15183, n15184, n15185, n15186, n15187, n15188,
         n15189, n15190, n15191, n15192, n15193, n15194, n15195, n15196,
         n15197, n15198, n15199, n15200, n15201, n15202, n15203, n15204,
         n15205, n15206, n15207, n15208, n15209, n15210, n15211, n15212,
         n15213, n15214, n15215, n15216, n15217, n15218, n15219, n15220,
         n15221, n15222, n15223, n15224, n15225, n15226, n15227, n15228,
         n15229, n15230, n15231, n15232, n15233, n15234, n15235, n15236,
         n15237, n15238, n15239, n15240, n15241, n15242, n15243, n15244,
         n15245, n15246, n15247, n15248, n15249, n15250, n15251, n15252,
         n15253, n15254, n15255, n15256, n15257, n15258, n15259, n15260,
         n15261, n15262, n15263, n15264, n15265, n15266, n15267, n15268,
         n15269, n15270, n15271, n15272, n15273, n15274, n15275, n15276,
         n15277, n15278, n15279, n15280, n15281, n15282, n15283, n15284,
         n15285, n15286, n15287, n15288, n15289, n15290, n15291, n15292,
         n15293, n15294, n15295, n15296, n15297, n15298, n15299, n15300,
         n15301, n15302, n15303, n15304, n15305, n15306, n15307, n15308,
         n15309, n15310, n15311, n15312, n15313, n15314, n15315, n15316,
         n15317, n15318, n15319, n15320, n15321, n15322, n15323, n15324,
         n15325, n15326, n15327, n15328, n15329, n15330, n15331, n15332,
         n15333, n15334, n15335, n15336, n15337, n15338, n15339, n15340,
         n15341, n15342, n15343, n15344, n15345, n15346, n15347, n15348,
         n15349, n15350, n15351, n15352, n15353, n15354, n15355, n15356,
         n15357, n15358, n15359, n15360, n15361, n15362, n15363, n15364,
         n15365, n15366, n15367, n15368, n15369, n15370, n15371, n15372,
         n15373, n15374, n15375, n15376, n15377, n15378, n15379, n15380,
         n15381, n15382, n15383, n15384, n15385, n15386, n15387, n15388,
         n15389, n15390, n15391, n15392, n15393, n15394, n15395, n15396,
         n15397, n15398, n15399, n15400, n15401, n15402, n15403, n15404,
         n15405, n15406, n15407, n15408, n15409, n15410, n15411, n15412,
         n15413, n15414, n15415, n15416, n15417, n15418, n15419, n15420,
         n15421, n15422, n15423, n15424, n15425, n15426, n15427, n15428,
         n15429, n15430, n15431, n15432, n15433, n15434, n15435, n15436,
         n15437, n15438, n15439, n15440, n15441, n15442, n15443, n15444,
         n15445, n15446, n15447, n15448, n15449, n15450, n15451, n15452,
         n15453, n15454, n15455, n15456, n15457, n15458, n15459, n15460,
         n15461, n15462, n15463, n15464, n15465, n15466, n15467, n15468,
         n15469, n15470, n15471, n15472, n15473, n15474, n15475, n15476,
         n15477, n15478, n15479, n15480, n15481, n15482, n15483, n15484,
         n15485, n15486, n15487, n15488, n15489, n15490, n15491, n15492,
         n15493, n15494, n15495, n15496, n15497, n15498, n15499, n15500,
         n15501, n15502, n15503, n15504, n15505, n15506, n15507, n15508,
         n15509, n15510, n15511, n15512, n15513, n15514, n15515, n15516,
         n15517, n15518, n15519, n15520, n15521, n15522, n15523, n15524,
         n15525, n15526, n15527, n15528, n15529, n15530, n15531, n15532,
         n15533, n15534, n15535, n15536, n15537, n15538, n15539, n15540,
         n15541, n15542, n15543, n15544, n15545, n15546, n15547, n15548,
         n15549, n15550, n15551, n15552, n15553, n15554, n15555, n15556,
         n15557, n15558, n15559, n15560, n15561, n15562, n15563, n15564,
         n15565, n15566, n15567, n15568, n15569, n15570, n15571, n15572,
         n15573, n15574, n15575, n15576, n15577, n15578, n15579, n15580,
         n15581, n15582, n15583, n15584, n15585, n15586, n15587, n15588,
         n15589, n15590, n15591, n15592, n15593, n15594, n15595, n15596,
         n15597, n15598, n15599, n15600, n15601, n15602, n15603, n15604,
         n15605, n15606, n15607, n15608, n15609, n15610, n15611, n15612,
         n15613, n15614, n15615, n15616, n15617, n15618, n15619, n15620,
         n15621, n15622, n15623, n15624, n15625, n15626, n15627, n15628,
         n15629, n15630, n15631, n15632, n15633, n15634, n15635, n15636,
         n15637, n15638, n15639, n15640, n15641, n15642, n15643, n15644,
         n15645, n15646, n15647, n15648, n15649, n15650, n15651, n15652,
         n15653, n15654, n15655, n15656, n15657, n15658, n15659, n15660,
         n15661, n15662, n15663, n15664, n15665, n15666, n15667, n15668,
         n15669, n15670, n15671, n15672, n15673, n15674, n15675, n15676,
         n15677, n15678, n15679, n15680, n15681, n15682, n15683, n15684,
         n15685, n15686, n15687, n15688, n15689, n15690, n15691, n15692,
         n15693, n15694, n15695, n15696, n15697, n15698, n15699, n15700,
         n15701, n15702, n15703, n15704, n15705, n15706, n15707, n15708,
         n15709, n15710, n15711, n15712, n15713, n15714, n15715, n15716,
         n15717, n15718, n15719, n15720, n15721, n15722, n15723, n15724,
         n15725, n15726, n15727, n15728, n15729, n15730, n15731, n15732,
         n15733, n15734, n15735, n15736, n15737, n15738, n15739, n15740,
         n15741, n15742, n15743, n15744, n15745, n15746, n15747, n15748,
         n15749, n15750, n15751, n15752, n15753, n15754, n15755, n15756,
         n15757, n15758, n15759, n15760, n15761, n15762, n15763, n15764,
         n15765, n15766, n15767, n15768, n15769, n15770, n15771, n15772,
         n15773, n15774, n15775, n15776, n15777, n15778, n15779, n15780,
         n15781, n15782, n15783, n15784, n15785, n15786, n15787, n15788,
         n15789, n15790, n15791, n15792, n15793, n15794, n15795, n15796,
         n15797, n15798, n15799, n15800, n15801, n15802, n15803, n15804,
         n15805, n15806, n15807, n15808, n15809, n15810, n15811, n15812,
         n15813, n15814, n15815, n15816, n15817, n15818, n15819, n15820,
         n15821, n15822, n15823, n15824, n15825, n15826, n15827, n15828,
         n15829, n15830, n15831, n15832, n15833, n15834, n15835, n15836,
         n15837, n15838, n15839, n15840, n15841, n15842, n15843, n15844,
         n15845, n15846, n15847, n15848, n15849, n15850, n15851, n15852,
         n15853, n15854, n15855, n15856, n15857, n15858, n15859, n15860,
         n15861, n15862, n15863, n15864, n15865, n15866, n15867, n15868,
         n15869, n15870, n15871, n15872, n15873, n15874, n15875, n15876,
         n15877, n15878, n15879, n15880, n15881, n15882, n15883, n15884,
         n15885, n15886, n15887, n15888, n15889, n15890, n15891, n15892,
         n15893, n15894, n15895, n15896, n15897, n15898, n15899, n15900,
         n15901, n15902, n15903, n15904, n15905, n15906, n15907, n15908,
         n15909, n15910, n15911, n15912, n15913, n15914, n15915, n15916,
         n15917, n15918, n15919, n15920, n15921, n15922, n15923, n15924,
         n15925, n15926, n15927, n15928, n15929, n15930, n15931, n15932,
         n15933, n15934, n15935, n15936, n15937, n15938, n15939, n15940,
         n15941, n15942, n15943, n15944, n15945, n15946, n15947, n15948,
         n15949, n15950, n15951, n15952, n15953, n15954, n15955, n15956,
         n15957, n15958, n15959, n15960, n15961, n15962, n15963, n15964,
         n15965, n15966, n15967, n15968, n15969, n15970, n15971, n15972,
         n15973, n15974, n15975, n15976, n15977, n15978, n15979, n15980,
         n15981, n15982, n15983, n15984, n15985, n15986, n15987, n15988,
         n15989, n15990, n15991, n15992, n15993, n15994, n15995, n15996,
         n15997, n15998, n15999, n16000, n16001, n16002, n16003, n16004,
         n16005, n16006, n16007, n16008, n16009, n16010, n16011, n16012,
         n16013, n16014, n16015, n16016, n16017, n16018, n16019, n16020,
         n16021, n16022, n16023, n16024, n16025, n16026, n16027, n16028,
         n16029, n16030, n16031, n16032, n16033, n16034, n16035, n16036,
         n16037, n16038, n16039, n16040, n16041, n16042, n16043, n16044,
         n16045, n16046, n16047, n16048, n16049, n16050, n16051, n16052,
         n16053, n16054, n16055, n16056, n16057, n16058, n16059, n16060,
         n16061, n16062, n16063, n16064, n16065, n16066, n16067, n16068,
         n16069, n16070, n16071, n16072, n16073, n16074, n16075, n16076,
         n16077, n16078, n16079, n16080, n16081, n16082, n16083, n16084,
         n16085, n16086, n16087, n16088, n16089, n16090, n16091, n16092,
         n16093, n16094, n16095, n16096, n16097, n16098, n16099, n16100,
         n16101, n16102, n16103, n16104, n16105, n16106, n16107, n16108,
         n16109, n16110, n16111, n16112, n16113, n16114, n16115, n16116,
         n16117, n16118, n16119, n16120, n16121, n16122, n16123, n16124,
         n16125, n16126, n16127, n16128, n16129, n16130, n16131, n16132,
         n16133, n16134, n16135, n16136, n16137, n16138, n16139, n16140,
         n16141, n16142, n16143, n16144, n16145, n16146, n16147, n16148,
         n16149, n16150, n16151, n16152, n16153, n16154, n16155, n16156,
         n16157, n16158, n16159, n16160, n16161, n16162, n16163, n16164,
         n16165, n16166, n16167, n16168, n16169, n16170, n16171, n16172,
         n16173, n16174, n16175, n16176, n16177, n16178, n16179, n16180,
         n16181, n16182, n16183, n16184, n16185, n16186, n16187, n16188,
         n16189, n16190, n16191, n16192, n16193, n16194, n16195, n16196,
         n16197, n16198, n16199, n16200, n16201, n16202, n16203, n16204,
         n16205, n16206, n16207, n16208, n16209, n16210, n16211, n16212,
         n16213, n16214, n16215, n16216, n16217, n16218, n16219, n16220,
         n16221, n16222, n16223, n16224, n16225, n16226, n16227, n16228,
         n16229, n16230, n16231, n16232, n16233, n16234, n16235, n16236,
         n16237, n16238, n16239, n16240, n16241, n16242, n16243, n16244,
         n16245, n16246, n16247, n16248, n16249, n16250, n16251, n16252,
         n16253, n16254, n16255, n16256, n16257, n16258, n16259, n16260,
         n16261, n16262, n16263, n16264, n16265, n16266, n16267, n16268,
         n16269, n16270, n16271, n16272, n16273, n16274, n16275, n16276,
         n16277, n16278, n16279, n16280, n16281, n16282, n16283, n16284,
         n16285, n16286, n16287, n16288, n16289, n16290, n16291, n16292,
         n16293, n16294, n16295, n16296, n16297, n16298, n16299, n16300,
         n16301, n16302, n16303, n16304, n16305, n16306, n16307, n16308,
         n16309, n16310, n16311, n16312, n16313, n16314, n16315, n16316,
         n16317, n16318, n16319, n16320, n16321, n16322, n16323, n16324,
         n16325, n16326, n16327, n16328, n16329, n16330, n16331, n16332,
         n16333, n16334, n16335, n16336, n16337, n16338, n16339, n16340,
         n16341, n16342, n16343, n16344, n16345, n16346, n16347, n16348,
         n16349, n16350, n16351, n16352, n16353, n16354, n16355, n16356,
         n16357, n16358, n16359, n16360, n16361, n16362, n16363, n16364,
         n16365, n16366, n16367, n16368, n16369, n16370, n16371, n16372,
         n16373, n16374, n16375, n16376, n16377, n16378, n16379, n16380,
         n16381, n16382, n16383, n16384, n16385, n16386, n16387, n16388,
         n16389, n16390, n16391, n16392, n16393, n16394, n16395, n16396,
         n16397, n16398, n16399, n16400, n16401, n16402, n16403, n16404,
         n16405, n16406, n16407, n16408, n16409, n16410, n16411, n16412,
         n16413, n16414, n16415, n16416, n16417, n16418, n16419, n16420,
         n16421, n16422, n16423, n16424, n16425, n16426, n16427, n16428,
         n16429, n16430, n16431, n16432, n16433, n16434, n16435, n16436,
         n16437, n16438, n16439, n16440, n16441, n16442, n16443, n16444,
         n16445, n16446, n16447, n16448, n16449, n16450, n16451, n16452,
         n16453, n16454, n16455, n16456, n16457, n16458, n16459, n16460,
         n16461, n16462, n16463, n16464, n16465, n16466, n16467, n16468,
         n16469, n16470, n16471, n16472, n16473, n16474, n16475, n16476,
         n16477, n16478, n16479, n16480, n16481, n16482, n16483, n16484,
         n16485, n16486, n16487, n16488, n16489, n16490, n16491, n16492,
         n16493, n16494, n16495, n16496, n16497, n16498, n16499, n16500,
         n16501, n16502, n16503, n16504, n16505, n16506, n16507, n16508,
         n16509, n16510, n16511, n16512, n16513, n16514, n16515, n16516,
         n16517, n16518, n16519, n16520, n16521, n16522, n16523, n16524,
         n16525, n16526, n16527, n16528, n16529, n16530, n16531, n16532,
         n16533, n16534, n16535, n16536, n16537, n16538, n16539, n16540,
         n16541, n16542, n16543, n16544, n16545, n16546, n16547, n16548,
         n16549, n16550, n16551, n16552, n16553, n16554, n16555, n16556,
         n16557, n16558, n16559, n16560, n16561, n16562, n16563, n16564,
         n16565, n16566, n16567, n16568, n16569, n16570, n16571, n16572,
         n16573, n16574, n16575, n16576, n16577, n16578, n16579, n16580,
         n16581, n16582, n16583, n16584, n16585, n16586, n16587, n16588,
         n16589, n16590, n16591, n16592, n16593, n16594, n16595, n16596,
         n16597, n16598, n16599, n16600, n16601, n16602, n16603, n16604,
         n16605, n16606, n16607, n16608, n16609, n16610, n16611, n16612,
         n16613, n16614, n16615, n16616, n16617, n16618, n16619, n16620,
         n16621, n16622, n16623, n16624, n16625, n16626, n16627, n16628,
         n16629, n16630, n16631, n16632, n16633, n16634, n16635, n16636,
         n16637, n16638, n16639, n16640, n16641, n16642, n16643, n16644,
         n16645, n16646, n16647, n16648, n16649, n16650, n16651, n16652,
         n16653, n16654, n16655, n16656, n16657, n16658, n16659, n16660,
         n16661, n16662, n16663, n16664, n16665, n16666, n16667, n16668,
         n16669, n16670, n16671, n16672, n16673, n16674, n16675, n16676,
         n16677, n16678, n16679, n16680, n16681, n16682, n16683, n16684,
         n16685, n16686, n16687, n16688, n16689, n16690, n16691, n16692,
         n16693, n16694, n16695, n16696, n16697, n16698, n16699, n16700,
         n16701, n16702, n16703, n16704, n16705, n16706, n16707, n16708,
         n16709, n16710, n16711, n16712, n16713, n16714, n16715, n16716,
         n16717, n16718, n16719, n16720, n16721, n16722, n16723, n16724,
         n16725, n16726, n16727, n16728, n16729, n16730, n16731, n16732,
         n16733, n16734, n16735, n16736, n16737, n16738, n16739, n16740,
         n16741, n16742, n16743, n16744, n16745, n16746, n16747, n16748,
         n16749, n16750, n16751, n16752, n16753, n16754, n16755, n16756,
         n16757, n16758, n16759, n16760, n16761, n16762, n16763, n16764,
         n16765, n16766, n16767, n16768, n16769, n16770, n16771, n16772,
         n16773, n16774, n16775, n16776, n16777, n16778, n16779, n16780,
         n16781, n16782, n16783, n16784, n16785, n16786, n16787, n16788,
         n16789, n16790, n16791, n16792, n16793, n16794, n16795, n16796,
         n16797, n16798, n16799, n16800, n16801, n16802, n16803, n16804,
         n16805, n16806, n16807, n16808, n16809, n16810, n16811, n16812,
         n16813, n16814, n16815, n16816, n16817, n16818, n16819, n16820,
         n16821, n16822, n16823, n16824, n16825, n16826, n16827, n16828,
         n16829, n16830, n16831, n16832, n16833, n16834, n16835, n16836,
         n16837, n16838, n16839, n16840, n16841, n16842, n16843, n16844,
         n16845, n16846, n16847, n16848, n16849, n16850, n16851, n16852,
         n16853, n16854, n16855, n16856, n16857, n16858, n16859, n16860,
         n16861, n16862, n16863, n16864, n16865, n16866, n16867, n16868,
         n16869, n16870, n16871, n16872, n16873, n16874, n16875, n16876,
         n16877, n16878, n16879, n16880, n16881, n16882, n16883, n16884,
         n16885, n16886, n16887, n16888, n16889, n16890, n16891, n16892,
         n16893, n16894, n16895, n16896, n16897, n16898, n16899, n16900,
         n16901, n16902, n16903, n16904, n16905, n16906, n16907, n16908,
         n16909, n16910, n16911, n16912, n16913, n16914, n16915, n16916,
         n16917, n16918, n16919, n16920, n16921, n16922, n16923, n16924,
         n16925, n16926, n16927, n16928, n16929, n16930, n16931, n16932,
         n16933, n16934, n16935, n16936, n16937, n16938, n16939, n16940,
         n16941, n16942, n16943, n16944, n16945, n16946, n16947, n16948,
         n16949, n16950, n16951, n16952, n16953, n16954, n16955, n16956,
         n16957, n16958, n16959, n16960, n16961, n16962, n16963, n16964,
         n16965, n16966, n16967, n16968, n16969, n16970, n16971, n16972,
         n16973, n16974, n16975, n16976, n16977, n16978, n16979, n16980,
         n16981, n16982, n16983, n16984, n16985, n16986, n16987, n16988,
         n16989, n16990, n16991, n16992, n16993, n16994, n16995, n16996,
         n16997, n16998, n16999, n17000, n17001, n17002, n17003, n17004,
         n17005, n17006, n17007, n17008, n17009, n17010, n17011, n17012,
         n17013, n17014, n17015, n17016, n17017, n17018, n17019, n17020,
         n17021, n17022, n17023, n17024, n17025, n17026, n17027, n17028,
         n17029, n17030, n17031, n17032, n17033, n17034, n17035, n17036,
         n17037, n17038, n17039, n17040, n17041, n17042, n17043, n17044,
         n17045, n17046, n17047, n17048, n17049, n17050, n17051, n17052,
         n17053, n17054, n17055, n17056, n17057, n17058, n17059, n17060,
         n17061, n17062, n17063, n17064, n17065, n17066, n17067, n17068,
         n17069, n17070, n17071, n17072, n17073, n17074, n17075, n17076,
         n17077, n17078, n17079, n17080, n17081, n17082, n17083, n17084,
         n17085, n17086, n17087, n17088, n17089, n17090, n17091, n17092,
         n17093, n17094, n17095, n17096, n17097, n17098, n17099, n17100,
         n17101, n17102, n17103, n17104, n17105, n17106, n17107, n17108,
         n17109, n17110, n17111, n17112, n17113, n17114, n17115, n17116,
         n17117, n17118, n17119, n17120, n17121, n17122, n17123, n17124,
         n17125, n17126, n17127, n17128, n17129, n17130, n17131, n17132,
         n17133, n17134, n17135, n17136, n17137, n17138, n17139, n17140,
         n17141, n17142, n17143, n17144, n17145, n17146, n17147, n17148,
         n17149, n17150, n17151, n17152, n17153, n17154, n17155, n17156,
         n17157, n17158, n17159, n17160, n17161, n17162, n17163, n17164,
         n17165, n17166, n17167, n17168, n17169, n17170, n17171, n17172,
         n17173, n17174, n17175, n17176, n17177, n17178, n17179, n17180,
         n17181, n17182, n17183, n17184, n17185, n17186, n17187, n17188,
         n17189, n17190, n17191, n17192, n17193, n17194, n17195, n17196,
         n17197, n17198, n17199, n17200, n17201, n17202, n17203, n17204,
         n17205, n17206, n17207, n17208, n17209, n17210, n17211, n17212,
         n17213, n17214, n17215, n17216, n17217, n17218, n17219, n17220,
         n17221, n17222, n17223, n17224, n17225, n17226, n17227, n17228,
         n17229, n17230, n17231, n17232, n17233, n17234, n17235, n17236,
         n17237, n17238, n17239, n17240, n17241, n17242, n17243, n17244,
         n17245, n17246, n17247, n17248, n17249, n17250, n17251, n17252,
         n17253, n17254, n17255, n17256, n17257, n17258, n17259, n17260,
         n17261, n17262, n17263, n17264, n17265, n17266, n17267, n17268,
         n17269, n17270, n17271, n17272, n17273, n17274, n17275, n17276,
         n17277, n17278, n17279, n17280, n17281, n17282, n17283, n17284,
         n17285, n17286, n17287, n17288, n17289, n17290, n17291, n17292,
         n17293, n17294, n17295, n17296, n17297, n17298, n17299, n17300,
         n17301, n17302, n17303, n17304, n17305, n17306, n17307, n17308,
         n17309, n17310, n17311, n17312, n17313, n17314, n17315, n17316,
         n17317, n17318, n17319, n17320, n17321, n17322, n17323, n17324,
         n17325, n17326, n17327, n17328, n17329, n17330, n17331, n17332,
         n17333, n17334, n17335, n17336, n17337, n17338, n17339, n17340,
         n17341, n17342, n17343, n17344, n17345, n17346, n17347, n17348,
         n17349, n17350, n17351, n17352, n17353, n17354, n17355, n17356,
         n17357, n17358, n17359, n17360, n17361, n17362, n17363, n17364,
         n17365, n17366, n17367, n17368, n17369, n17370, n17371, n17372,
         n17373, n17374, n17375, n17376, n17377, n17378, n17379, n17380,
         n17381, n17382, n17383, n17384, n17385, n17386, n17387, n17388,
         n17389, n17390, n17391, n17392, n17393, n17394, n17395, n17396,
         n17397, n17398, n17399, n17400, n17401, n17402, n17403, n17404,
         n17405, n17406, n17407, n17408, n17409, n17410, n17411, n17412,
         n17413, n17414, n17415, n17416, n17417, n17418, n17419, n17420,
         n17421, n17422, n17423, n17424, n17425, n17426, n17427, n17428,
         n17429, n17430, n17431, n17432, n17433, n17434, n17435, n17436,
         n17437, n17438, n17439, n17440, n17441, n17442, n17443, n17444,
         n17445, n17446, n17447, n17448, n17449, n17450, n17451, n17452,
         n17453, n17454, n17455, n17456, n17457, n17458, n17459, n17460,
         n17461, n17462, n17463, n17464, n17465, n17466, n17467, n17468,
         n17469, n17470, n17471, n17472, n17473, n17474, n17475, n17476,
         n17477, n17478, n17479, n17480, n17481, n17482, n17483, n17484,
         n17485, n17486, n17487, n17488, n17489, n17490, n17491, n17492,
         n17493, n17494, n17495, n17496, n17497, n17498, n17499, n17500,
         n17501, n17502, n17503, n17504, n17505, n17506, n17507, n17508,
         n17509, n17510, n17511, n17512, n17513, n17514, n17515, n17516,
         n17517, n17518, n17519, n17520, n17521, n17522, n17523, n17524,
         n17525, n17526, n17527, n17528, n17529, n17530, n17531, n17532,
         n17533, n17534, n17535, n17536, n17537, n17538, n17539, n17540,
         n17541, n17542, n17543, n17544, n17545, n17546, n17547, n17548,
         n17549, n17550, n17551, n17552, n17553, n17554, n17555, n17556,
         n17557, n17558, n17559, n17560, n17561, n17562, n17563, n17564,
         n17565, n17566, n17567, n17568, n17569, n17570, n17571, n17572,
         n17573, n17574, n17575, n17576, n17577, n17578, n17579, n17580,
         n17581, n17582, n17583, n17584, n17585, n17586, n17587, n17588,
         n17589, n17590, n17591, n17592, n17593, n17594, n17595, n17596,
         n17597, n17598, n17599, n17600, n17601, n17602, n17603, n17604,
         n17605, n17606, n17607, n17608, n17609, n17610, n17611, n17612,
         n17613, n17614, n17615, n17616, n17617, n17618, n17619, n17620,
         n17621, n17622, n17623, n17624, n17625, n17626, n17627, n17628,
         n17629, n17630, n17631, n17632, n17633, n17634, n17635, n17636,
         n17637, n17638, n17639, n17640, n17641, n17642, n17643, n17644,
         n17645, n17646, n17647, n17648, n17649, n17650, n17651, n17652,
         n17653, n17654, n17655, n17656, n17657, n17658, n17659, n17660,
         n17661, n17662, n17663, n17664, n17665, n17666, n17667, n17668,
         n17669, n17670, n17671, n17672, n17673, n17674, n17675, n17676,
         n17677, n17678, n17679, n17680, n17681, n17682, n17683, n17684,
         n17685, n17686, n17687, n17688, n17689, n17690, n17691, n17692,
         n17693, n17694, n17695, n17696, n17697, n17698, n17699, n17700,
         n17701, n17702, n17703, n17704, n17705, n17706, n17707, n17708,
         n17709, n17710, n17711, n17712, n17713, n17714, n17715, n17716,
         n17717, n17718, n17719, n17720, n17721, n17722, n17723, n17724,
         n17725, n17726, n17727, n17728, n17729, n17730, n17731, n17732,
         n17733, n17734, n17735, n17736, n17737, n17738, n17739, n17740,
         n17741, n17742, n17743, n17744, n17745, n17746, n17747, n17748,
         n17749, n17750, n17751, n17752, n17753, n17754, n17755, n17756,
         n17757, n17758, n17759, n17760, n17761, n17762, n17763, n17764,
         n17765, n17766, n17767, n17768, n17769, n17770, n17771, n17772,
         n17773, n17774, n17775, n17776, n17777, n17778, n17779, n17780,
         n17781, n17782, n17783, n17784, n17785, n17786, n17787, n17788,
         n17789, n17790, n17791, n17792, n17793, n17794, n17795, n17796,
         n17797, n17798, n17799, n17800, n17801, n17802, n17803, n17804,
         n17805, n17806, n17807, n17808, n17809, n17810, n17811, n17812,
         n17813, n17814, n17815, n17816, n17817, n17818, n17819, n17820,
         n17821, n17822, n17823, n17824, n17825, n17826, n17827, n17828,
         n17829, n17830, n17831, n17832, n17833, n17834, n17835, n17836,
         n17837, n17838, n17839, n17840, n17841, n17842, n17843, n17844,
         n17845, n17846, n17847, n17848, n17849, n17850, n17851, n17852,
         n17853, n17854, n17855, n17856, n17857, n17858, n17859, n17860,
         n17861, n17862, n17863, n17864, n17865, n17866, n17867, n17868,
         n17869, n17870, n17871, n17872, n17873, n17874, n17875, n17876,
         n17877, n17878, n17879, n17880, n17881, n17882, n17883, n17884,
         n17885, n17886, n17887, n17888, n17889, n17890, n17891, n17892,
         n17893, n17894, n17895, n17896, n17897, n17898, n17899, n17900,
         n17901, n17902, n17903, n17904, n17905, n17906, n17907, n17908,
         n17909, n17910, n17911, n17912, n17913, n17914, n17915, n17916,
         n17917, n17918, n17919, n17920, n17921, n17922, n17923, n17924,
         n17925, n17926, n17927, n17928, n17929, n17930, n17931, n17932,
         n17933, n17934, n17935, n17936, n17937, n17938, n17939, n17940,
         n17941, n17942, n17943, n17944, n17945, n17946, n17947, n17948,
         n17949, n17950, n17951, n17952, n17953, n17954, n17955, n17956,
         n17957, n17958, n17959, n17960, n17961, n17962, n17963, n17964,
         n17965, n17966, n17967, n17968, n17969, n17970, n17971, n17972,
         n17973, n17974, n17975, n17976, n17977, n17978, n17979, n17980,
         n17981, n17982, n17983, n17984, n17985, n17986, n17987, n17988,
         n17989, n17990, n17991, n17992, n17993, n17994, n17995, n17996,
         n17997, n17998, n17999, n18000, n18001, n18002, n18003, n18004,
         n18005, n18006, n18007, n18008, n18009, n18010, n18011, n18012,
         n18013, n18014, n18015, n18016, n18017, n18018, n18019, n18020,
         n18021, n18022, n18023, n18024, n18025, n18026, n18027, n18028,
         n18029, n18030, n18031, n18032, n18033, n18034, n18035, n18036,
         n18037, n18038, n18039, n18040, n18041, n18042, n18043, n18044,
         n18045, n18046, n18047, n18048, n18049, n18050, n18051, n18052,
         n18053, n18054, n18055, n18056, n18057, n18058, n18059, n18060,
         n18061, n18062, n18063, n18064, n18065, n18066, n18067, n18068,
         n18069, n18070, n18071, n18072, n18073, n18074, n18075, n18076,
         n18077, n18078, n18079, n18080, n18081, n18082, n18083, n18084,
         n18085, n18086, n18087, n18088, n18089, n18090, n18091, n18092,
         n18093, n18094, n18095, n18096, n18097, n18098, n18099, n18100,
         n18101, n18102, n18103, n18104, n18105, n18106, n18107, n18108,
         n18109, n18110, n18111, n18112, n18113, n18114, n18115, n18116,
         n18117, n18118, n18119, n18120, n18121, n18122, n18123, n18124,
         n18125, n18126, n18127, n18128, n18129, n18130, n18131, n18132,
         n18133, n18134, n18135, n18136, n18137, n18138, n18139, n18140,
         n18141, n18142, n18143, n18144, n18145, n18146, n18147, n18148,
         n18149, n18150, n18151, n18152, n18153, n18154, n18155, n18156,
         n18157, n18158, n18159, n18160, n18161, n18162, n18163, n18164,
         n18165, n18166, n18167, n18168, n18169, n18170, n18171, n18172,
         n18173, n18174, n18175, n18176, n18177, n18178, n18179, n18180,
         n18181, n18182, n18183, n18184, n18185, n18186, n18187, n18188,
         n18189, n18190, n18191, n18192, n18193, n18194, n18195, n18196,
         n18197, n18198, n18199, n18200, n18201, n18202, n18203, n18204,
         n18205, n18206, n18207, n18208, n18209, n18210, n18211, n18212,
         n18213, n18214, n18215, n18216, n18217, n18218, n18219, n18220,
         n18221, n18222, n18223, n18224, n18225, n18226, n18227, n18228,
         n18229, n18230, n18231, n18232, n18233, n18234, n18235, n18236,
         n18237, n18238, n18239, n18240, n18241, n18242, n18243, n18244,
         n18245, n18246, n18247, n18248, n18249, n18250, n18251, n18252,
         n18253, n18254, n18255, n18256, n18257, n18258, n18259, n18260,
         n18261, n18262, n18263, n18264, n18265, n18266, n18267, n18268,
         n18269, n18270, n18271, n18272, n18273, n18274, n18275, n18276,
         n18277, n18278, n18279, n18280, n18281, n18282, n18283, n18284,
         n18285, n18286, n18287, n18288, n18289, n18290, n18291, n18292,
         n18293, n18294, n18295, n18296, n18297, n18298, n18299, n18300,
         n18301, n18302, n18303, n18304, n18305, n18306, n18307, n18308,
         n18309, n18310, n18311, n18312, n18313, n18314, n18315, n18316,
         n18317, n18318, n18319, n18320, n18321, n18322, n18323, n18324,
         n18325, n18326, n18327, n18328, n18329, n18330, n18331, n18332,
         n18333, n18334, n18335, n18336, n18337, n18338, n18339, n18340,
         n18341, n18342, n18343, n18344, n18345, n18346, n18347, n18348,
         n18349, n18350, n18351, n18352, n18353, n18354, n18355, n18356,
         n18357, n18358, n18359, n18360, n18361, n18362, n18363, n18364,
         n18365, n18366, n18367, n18368, n18369, n18370, n18371, n18372,
         n18373, n18374, n18375, n18376, n18377, n18378, n18379, n18380,
         n18381, n18382, n18383, n18384, n18385, n18386, n18387, n18388,
         n18389, n18390, n18391, n18392, n18393, n18394, n18395, n18396,
         n18397, n18398, n18399, n18400, n18401, n18402, n18403, n18404,
         n18405, n18406, n18407, n18408, n18409, n18410, n18411, n18412,
         n18413, n18414, n18415, n18416, n18417, n18418, n18419, n18420,
         n18421, n18422, n18423, n18424, n18425, n18426, n18427, n18428,
         n18429, n18430, n18431, n18432, n18433, n18434, n18435, n18436,
         n18437, n18438, n18439, n18440, n18441, n18442, n18443, n18444,
         n18445, n18446, n18447, n18448, n18449, n18450, n18451, n18452,
         n18453, n18454, n18455, n18456, n18457, n18458, n18459, n18460,
         n18461, n18462, n18463, n18464, n18465, n18466, n18467, n18468,
         n18469, n18470, n18471, n18472, n18473, n18474, n18475, n18476,
         n18477, n18478, n18479, n18480, n18481, n18482, n18483, n18484,
         n18485, n18486, n18487, n18488, n18489, n18490, n18491, n18492,
         n18493, n18494, n18495, n18496, n18497, n18498, n18499, n18500,
         n18501, n18502, n18503, n18504, n18505, n18506, n18507, n18508,
         n18509, n18510, n18511, n18512, n18513, n18514, n18515, n18516,
         n18517, n18518, n18519, n18520, n18521, n18522, n18523, n18524,
         n18525, n18526, n18527, n18528, n18529, n18530, n18531, n18532,
         n18533, n18534, n18535, n18536, n18537, n18538, n18539, n18540,
         n18541, n18542, n18543, n18544, n18545, n18546, n18547, n18548,
         n18549, n18550, n18551, n18552, n18553, n18554, n18555, n18556,
         n18557, n18558, n18559, n18560, n18561, n18562, n18563, n18564,
         n18565, n18566, n18567, n18568, n18569, n18570, n18571, n18572,
         n18573, n18574, n18575, n18576, n18577, n18578, n18579, n18580,
         n18581, n18582, n18583, n18584, n18585, n18586, n18587, n18588,
         n18589, n18590, n18591, n18592, n18593, n18594, n18595, n18596,
         n18597, n18598, n18599, n18600, n18601, n18602, n18603, n18604,
         n18605, n18606, n18607, n18608, n18609, n18610, n18611, n18612,
         n18613, n18614, n18615, n18616, n18617, n18618, n18619, n18620,
         n18621, n18622, n18623, n18624, n18625, n18626, n18627, n18628,
         n18629, n18630, n18631, n18632, n18633, n18634, n18635, n18636,
         n18637, n18638, n18639, n18640, n18641, n18642, n18643, n18644,
         n18645, n18646, n18647, n18648, n18649, n18650, n18651, n18652,
         n18653, n18654, n18655, n18656, n18657, n18658, n18659, n18660,
         n18661, n18662, n18663, n18664, n18665, n18666, n18667, n18668,
         n18669, n18670, n18671, n18672, n18673, n18674, n18675, n18676,
         n18677, n18678, n18679, n18680, n18681, n18682, n18683, n18684,
         n18685, n18686, n18687, n18688, n18689, n18690, n18691, n18692,
         n18693, n18694, n18695, n18696, n18697, n18698, n18699, n18700,
         n18701, n18702, n18703, n18704, n18705, n18706, n18707, n18708,
         n18709, n18710, n18711, n18712, n18713, n18714, n18715, n18716,
         n18717, n18718, n18719, n18720, n18721, n18722, n18723, n18724,
         n18725, n18726, n18727, n18728, n18729, n18730, n18731, n18732,
         n18733, n18734, n18735, n18736, n18737, n18738, n18739, n18740,
         n18741, n18742, n18743, n18744, n18745, n18746, n18747, n18748,
         n18749, n18750, n18751, n18752, n18753, n18754, n18755, n18756,
         n18757, n18758, n18759, n18760, n18761, n18762, n18763, n18764,
         n18765, n18766, n18767, n18768, n18769, n18770, n18771, n18772,
         n18773, n18774, n18775, n18776, n18777, n18778, n18779, n18780,
         n18781, n18782, n18783, n18784, n18785, n18786, n18787, n18788,
         n18789, n18790, n18791, n18792, n18793, n18794, n18795, n18796,
         n18797, n18798, n18799, n18800, n18801, n18802, n18803, n18804,
         n18805, n18806, n18807, n18808, n18809, n18810, n18811, n18812,
         n18813, n18814, n18815, n18816, n18817, n18818, n18819, n18820,
         n18821, n18822, n18823, n18824, n18825, n18826, n18827, n18828,
         n18829, n18830, n18831, n18832, n18833, n18834, n18835, n18836,
         n18837, n18838, n18839, n18840, n18841, n18842, n18843, n18844,
         n18845, n18846, n18847, n18848, n18849, n18850, n18851, n18852,
         n18853, n18854, n18855, n18856, n18857, n18858, n18859, n18860,
         n18861, n18862, n18863, n18864, n18865, n18866, n18867, n18868,
         n18869, n18870, n18871, n18872, n18873, n18874, n18875, n18876,
         n18877, n18878, n18879, n18880, n18881, n18882, n18883, n18884,
         n18885, n18886, n18887, n18888, n18889, n18890, n18891, n18892,
         n18893, n18894, n18895, n18896, n18897, n18898, n18899, n18900,
         n18901, n18902, n18903, n18904, n18905, n18906, n18907, n18908,
         n18909, n18910, n18911, n18912, n18913, n18914, n18915, n18916,
         n18917, n18918, n18919, n18920, n18921, n18922, n18923, n18924,
         n18925, n18926, n18927, n18928, n18929, n18930, n18931, n18932,
         n18933, n18934, n18935, n18936, n18937, n18938, n18939, n18940,
         n18941, n18942, n18943, n18944, n18945, n18946, n18947, n18948,
         n18949, n18950, n18951, n18952, n18953, n18954, n18955, n18956,
         n18957, n18958, n18959, n18960, n18961, n18962, n18963, n18964,
         n18965, n18966, n18967, n18968, n18969, n18970, n18971, n18972,
         n18973, n18974, n18975, n18976, n18977, n18978, n18979, n18980,
         n18981, n18982, n18983, n18984, n18985, n18986, n18987, n18988,
         n18989, n18990, n18991, n18992, n18993, n18994, n18995, n18996,
         n18997, n18998, n18999, n19000, n19001, n19002, n19003, n19004,
         n19005, n19006, n19007, n19008, n19009, n19010, n19011, n19012,
         n19013, n19014, n19015, n19016, n19017, n19018, n19019, n19020,
         n19021, n19022, n19023, n19024, n19025, n19026, n19027, n19028,
         n19029, n19030, n19031, n19032, n19033, n19034, n19035, n19036,
         n19037, n19038, n19039, n19040, n19041, n19042, n19043, n19044,
         n19045, n19046, n19047, n19048, n19049, n19050, n19051, n19052,
         n19053, n19054, n19055, n19056, n19057, n19058, n19059, n19060,
         n19061, n19062, n19063, n19064, n19065, n19066, n19067, n19068,
         n19069, n19070, n19071, n19072, n19073, n19074, n19075, n19076,
         n19077, n19078, n19079, n19080, n19081, n19082, n19083, n19084,
         n19085, n19086, n19087, n19088, n19089, n19090, n19091, n19092,
         n19093, n19094, n19095, n19096, n19097, n19098, n19099, n19100,
         n19101, n19102, n19103, n19104, n19105, n19106, n19107, n19108,
         n19109, n19110, n19111, n19112, n19113, n19114, n19115, n19116,
         n19117, n19118, n19119, n19120, n19121, n19122, n19123, n19124,
         n19125, n19126, n19127, n19128, n19129, n19130, n19131, n19132,
         n19133, n19134, n19135, n19136, n19137, n19138, n19139, n19140,
         n19141, n19142, n19143, n19144, n19145, n19146, n19147, n19148,
         n19149, n19150, n19151, n19152, n19153, n19154, n19155, n19156,
         n19157, n19158, n19159, n19160, n19161, n19162, n19163, n19164,
         n19165, n19166, n19167, n19168, n19169, n19170, n19171, n19172,
         n19173, n19174, n19175, n19176, n19177, n19178, n19179, n19180,
         n19181, n19182, n19183, n19184, n19185, n19186, n19187, n19188,
         n19189, n19190, n19191, n19192, n19193, n19194, n19195, n19196,
         n19197, n19198, n19199, n19200, n19201, n19202, n19203, n19204,
         n19205, n19206, n19207, n19208, n19209, n19210, n19211, n19212,
         n19213, n19214, n19215, n19216, n19217, n19218, n19219, n19220,
         n19221, n19222, n19223, n19224, n19225, n19226, n19227, n19228,
         n19229, n19230, n19231, n19232, n19233, n19234, n19235, n19236,
         n19237, n19238, n19239, n19240, n19241, n19242, n19243, n19244,
         n19245, n19246, n19247, n19248, n19249, n19250, n19251, n19252,
         n19253, n19254, n19255, n19256, n19257, n19258, n19259, n19260,
         n19261, n19262, n19263, n19264, n19265, n19266, n19267, n19268,
         n19269, n19270, n19271, n19272, n19273, n19274, n19275, n19276,
         n19277, n19278, n19279, n19280, n19281, n19282, n19283, n19284,
         n19285, n19286, n19287, n19288, n19289, n19290, n19291, n19292,
         n19293, n19294, n19295, n19296, n19297, n19298, n19299, n19300,
         n19301, n19302, n19303, n19304, n19305, n19306, n19307, n19308,
         n19309, n19310, n19311, n19312, n19313, n19314, n19315, n19316,
         n19317, n19318, n19319, n19320, n19321, n19322, n19323, n19324,
         n19325, n19326, n19327, n19328, n19329, n19330, n19331, n19332,
         n19333, n19334, n19335, n19336, n19337, n19338, n19339, n19340,
         n19341, n19342, n19343, n19344, n19345, n19346, n19347, n19348,
         n19349, n19350, n19351, n19352, n19353, n19354, n19355, n19356,
         n19357, n19358, n19359, n19360, n19361, n19362, n19363, n19364,
         n19365, n19366, n19367, n19368, n19369, n19370, n19371, n19372,
         n19373, n19374, n19375, n19376, n19377, n19378, n19379, n19380,
         n19381, n19382, n19383, n19384, n19385, n19386, n19387, n19388,
         n19389, n19390, n19391, n19392, n19393, n19394, n19395, n19396,
         n19397, n19398, n19399, n19400, n19401, n19402, n19403, n19404,
         n19405, n19406, n19407, n19408, n19409, n19410, n19411, n19412,
         n19413, n19414, n19415, n19416, n19417, n19418, n19419, n19420,
         n19421, n19422, n19423, n19424, n19425, n19426, n19427, n19428,
         n19429, n19430, n19431, n19432, n19433, n19434, n19435, n19436,
         n19437, n19438, n19439, n19440, n19441, n19442, n19443, n19444,
         n19445, n19446, n19447, n19448, n19449, n19450, n19451, n19452,
         n19453, n19454, n19455, n19456, n19457, n19458, n19459, n19460,
         n19461, n19462, n19463, n19464, n19465, n19466, n19467, n19468,
         n19469, n19470, n19471, n19472, n19473, n19474, n19475, n19476,
         n19477, n19478, n19479, n19480, n19481, n19482, n19483, n19484,
         n19485, n19486, n19487, n19488, n19489, n19490, n19491, n19492,
         n19493, n19494, n19495, n19496, n19497, n19498, n19499, n19500,
         n19501, n19502, n19503, n19504, n19505, n19506, n19507, n19508,
         n19509, n19510, n19511, n19512, n19513, n19514, n19515, n19516,
         n19517, n19518, n19519, n19520, n19521, n19522, n19523, n19524,
         n19525, n19526, n19527, n19528, n19529, n19530, n19531, n19532,
         n19533, n19534, n19535, n19536, n19537, n19538, n19539, n19540,
         n19541, n19542, n19543, n19544, n19545, n19546, n19547, n19548,
         n19549, n19550, n19551, n19552, n19553, n19554, n19555, n19556,
         n19557, n19558, n19559, n19560, n19561, n19562, n19563, n19564,
         n19565, n19566, n19567, n19568, n19569, n19570, n19571, n19572,
         n19573, n19574, n19575, n19576, n19577, n19578, n19579, n19580,
         n19581, n19582, n19583, n19584, n19585, n19586, n19587, n19588,
         n19589, n19590, n19591, n19592, n19593, n19594, n19595, n19596,
         n19597, n19598, n19599, n19600, n19601, n19602, n19603, n19604,
         n19605, n19606, n19607, n19608, n19609, n19610, n19611, n19612,
         n19613, n19614, n19615, n19616, n19617, n19618, n19619, n19620,
         n19621, n19622, n19623, n19624, n19625, n19626, n19627, n19628,
         n19629, n19630, n19631, n19632, n19633, n19634, n19635, n19636,
         n19637, n19638, n19639, n19640, n19641, n19642, n19643, n19644,
         n19645, n19646, n19647, n19648, n19649, n19650, n19651, n19652,
         n19653, n19654, n19655, n19656, n19657, n19658, n19659, n19660,
         n19661, n19662, n19663, n19664, n19665, n19666, n19667, n19668,
         n19669, n19670, n19671, n19672, n19673, n19674, n19675, n19676,
         n19677, n19678, n19679, n19680, n19681, n19682, n19683, n19684,
         n19685, n19686, n19687, n19688, n19689, n19690, n19691, n19692,
         n19693, n19694, n19695, n19696, n19697, n19698, n19699, n19700,
         n19701, n19702, n19703, n19704, n19705, n19706, n19707, n19708,
         n19709, n19710, n19711, n19712, n19713, n19714, n19715, n19716,
         n19717, n19718, n19719, n19720, n19721, n19722, n19723, n19724,
         n19725, n19726, n19727, n19728, n19729, n19730, n19731, n19732,
         n19733, n19734, n19735, n19736, n19737, n19738, n19739, n19740,
         n19741, n19742, n19743, n19744, n19745, n19746, n19747, n19748,
         n19749, n19750, n19751, n19752, n19753, n19754, n19755, n19756,
         n19757, n19758, n19759, n19760, n19761, n19762, n19763, n19764,
         n19765, n19766, n19767, n19768, n19769, n19770, n19771, n19772,
         n19773, n19774, n19775, n19776, n19777, n19778, n19779, n19780,
         n19781, n19782, n19783, n19784, n19785, n19786, n19787, n19788,
         n19789, n19790, n19791, n19792, n19793, n19794, n19795, n19796,
         n19797, n19798, n19799, n19800, n19801, n19802, n19803, n19804,
         n19805, n19806, n19807, n19808, n19809, n19810, n19811, n19812,
         n19813, n19814, n19815, n19816, n19817, n19818, n19819, n19820,
         n19821, n19822, n19823, n19824, n19825, n19826, n19827, n19828,
         n19829, n19830, n19831, n19832, n19833, n19834, n19835, n19836,
         n19837, n19838, n19839, n19840, n19841, n19842, n19843, n19844,
         n19845, n19846, n19847, n19848, n19849, n19850, n19851, n19852,
         n19853, n19854, n19855, n19856, n19857, n19858, n19859, n19860,
         n19861, n19862, n19863, n19864, n19865, n19866, n19867, n19868,
         n19869, n19870, n19871, n19872, n19873, n19874, n19875, n19876,
         n19877, n19878, n19879, n19880, n19881, n19882, n19883, n19884,
         n19885, n19886, n19887, n19888, n19889, n19890, n19891, n19892,
         n19893, n19894, n19895, n19896, n19897, n19898, n19899, n19900,
         n19901, n19902, n19903, n19904, n19905, n19906, n19907, n19908,
         n19909, n19910, n19911, n19912, n19913, n19914, n19915, n19916,
         n19917, n19918, n19919, n19920, n19921, n19922, n19923, n19924,
         n19925, n19926, n19927, n19928, n19929, n19930, n19931, n19932,
         n19933, n19934, n19935, n19936, n19937, n19938, n19939, n19940,
         n19941, n19942, n19943, n19944, n19945, n19946, n19947, n19948,
         n19949, n19950, n19951, n19952, n19953, n19954, n19955, n19956,
         n19957, n19958, n19959, n19960, n19961, n19962, n19963, n19964,
         n19965, n19966, n19967, n19968, n19969, n19970, n19971, n19972,
         n19973, n19974, n19975, n19976, n19977, n19978, n19979, n19980,
         n19981, n19982, n19983, n19984, n19985, n19986, n19987, n19988,
         n19989, n19990, n19991, n19992, n19993, n19994, n19995, n19996,
         n19997, n19998, n19999, n20000, n20001, n20002, n20003, n20004,
         n20005, n20006, n20007, n20008, n20009, n20010, n20011, n20012,
         n20013, n20014, n20015, n20016, n20017, n20018, n20019, n20020,
         n20021, n20022, n20023, n20024, n20025, n20026, n20027, n20028,
         n20029, n20030, n20031, n20032, n20033, n20034, n20035, n20036,
         n20037, n20038, n20039, n20040, n20041, n20042, n20043, n20044,
         n20045, n20046, n20047, n20048, n20049, n20050, n20051, n20052,
         n20053, n20054, n20055, n20056, n20057, n20058, n20059, n20060,
         n20061, n20062, n20063, n20064, n20065, n20066, n20067, n20068,
         n20069, n20070, n20071, n20072, n20073, n20074, n20075, n20076,
         n20077, n20078, n20079, n20080, n20081, n20082, n20083, n20084,
         n20085, n20086, n20087, n20088, n20089, n20090, n20091, n20092,
         n20093, n20094, n20095, n20096, n20097, n20098, n20099, n20100,
         n20101, n20102, n20103, n20104, n20105, n20106, n20107, n20108,
         n20109, n20110, n20111, n20112, n20113, n20114, n20115, n20116,
         n20117, n20118, n20119, n20120, n20121, n20122, n20123, n20124,
         n20125, n20126, n20127, n20128, n20129, n20130, n20131, n20132,
         n20133, n20134, n20135, n20136, n20137, n20138, n20139, n20140,
         n20141, n20142, n20143, n20144, n20145, n20146, n20147, n20148,
         n20149, n20150, n20151, n20152, n20153, n20154, n20155, n20156,
         n20157, n20158, n20159, n20160, n20161, n20162, n20163, n20164,
         n20165, n20166, n20167, n20168, n20169, n20170, n20171, n20172,
         n20173, n20174, n20175, n20176, n20177, n20178, n20179, n20180,
         n20181, n20182, n20183, n20184, n20185, n20186, n20187, n20188,
         n20189, n20190, n20191, n20192, n20193, n20194, n20195, n20196,
         n20197, n20198, n20199, n20200, n20201, n20202, n20203, n20204,
         n20205, n20206, n20207, n20208, n20209, n20210, n20211, n20212,
         n20213, n20214, n20215, n20216, n20217, n20218, n20219, n20220,
         n20221, n20222, n20223, n20224, n20225, n20226, n20227, n20228,
         n20229, n20230, n20231, n20232, n20233, n20234, n20235, n20236,
         n20237, n20238, n20239, n20240, n20241, n20242, n20243, n20244,
         n20245, n20246, n20247, n20248, n20249, n20250, n20251, n20252,
         n20253, n20254, n20255, n20256, n20257, n20258, n20259, n20260,
         n20261, n20262, n20263, n20264, n20265, n20266, n20267, n20268,
         n20269, n20270, n20271, n20272, n20273, n20274, n20275, n20276,
         n20277, n20278, n20279, n20280, n20281, n20282, n20283, n20284,
         n20285, n20286, n20287, n20288, n20289, n20290, n20291, n20292,
         n20293, n20294, n20295, n20296, n20297, n20298, n20299, n20300,
         n20301, n20302, n20303, n20304, n20305, n20306, n20307, n20308,
         n20309, n20310, n20311, n20312, n20313, n20314, n20315, n20316,
         n20317, n20318, n20319, n20320, n20321, n20322, n20323, n20324,
         n20325, n20326, n20327, n20328, n20329, n20330, n20331, n20332,
         n20333, n20334, n20335, n20336, n20337, n20338, n20339, n20340,
         n20341, n20342, n20343, n20344, n20345, n20346, n20347, n20348,
         n20349, n20350, n20351, n20352, n20353, n20354, n20355, n20356,
         n20357, n20358, n20359, n20360, n20361, n20362, n20363, n20364,
         n20365, n20366, n20367, n20368, n20369, n20370, n20371, n20372,
         n20373, n20374, n20375, n20376, n20377, n20378, n20379, n20380,
         n20381, n20382, n20383, n20384, n20385, n20386, n20387, n20388,
         n20389, n20390, n20391, n20392, n20393, n20394, n20395, n20396,
         n20397, n20398, n20399, n20400, n20401, n20402, n20403, n20404,
         n20405, n20406, n20407, n20408, n20409, n20410, n20411, n20412,
         n20413, n20414, n20415, n20416, n20417, n20418, n20419, n20420,
         n20421, n20422, n20423, n20424, n20425, n20426, n20427, n20428,
         n20429, n20430, n20431, n20432, n20433, n20434, n20435, n20436,
         n20437, n20438, n20439, n20440, n20441, n20442, n20443, n20444,
         n20445, n20446, n20447, n20448, n20449, n20450, n20451, n20452,
         n20453, n20454, n20455, n20456, n20457, n20458, n20459, n20460,
         n20461, n20462, n20463, n20464, n20465, n20466, n20467, n20468,
         n20469, n20470, n20471, n20472, n20473, n20474, n20475, n20476,
         n20477, n20478, n20479, n20480, n20481, n20482, n20483, n20484,
         n20485, n20486, n20487, n20488, n20489, n20490, n20491, n20492,
         n20493, n20494, n20495, n20496, n20497, n20498, n20499, n20500,
         n20501, n20502, n20503, n20504, n20505, n20506, n20507, n20508,
         n20509, n20510, n20511, n20512, n20513, n20514, n20515, n20516,
         n20517, n20518, n20519, n20520, n20521, n20522, n20523, n20524,
         n20525, n20526, n20527, n20528, n20529, n20530, n20531, n20532,
         n20533, n20534, n20535, n20536, n20537, n20538, n20539, n20540,
         n20541, n20542, n20543, n20544, n20545, n20546, n20547, n20548,
         n20549, n20550, n20551, n20552, n20553, n20554, n20555, n20556,
         n20557, n20558, n20559, n20560, n20561, n20562, n20563, n20564,
         n20565, n20566, n20567, n20568, n20569, n20570, n20571, n20572,
         n20573, n20574, n20575, n20576, n20577, n20578, n20579, n20580,
         n20581, n20582, n20583, n20584, n20585, n20586, n20587, n20588,
         n20589, n20590, n20591, n20592, n20593, n20594, n20595, n20596,
         n20597, n20598, n20599, n20600, n20601, n20602, n20603, n20604,
         n20605, n20606, n20607, n20608, n20609, n20610, n20611, n20612,
         n20613, n20614, n20615, n20616, n20617, n20618, n20619, n20620,
         n20621, n20622, n20623, n20624, n20625, n20626, n20627, n20628,
         n20629, n20630, n20631, n20632, n20633, n20634, n20635, n20636,
         n20637, n20638, n20639, n20640, n20641, n20642, n20643, n20644,
         n20645, n20646, n20647, n20648, n20649, n20650, n20651, n20652,
         n20653, n20654, n20655, n20656, n20657, n20658, n20659, n20660,
         n20661, n20662, n20663, n20664, n20665, n20666, n20667, n20668,
         n20669, n20670, n20671, n20672, n20673, n20674, n20675, n20676,
         n20677, n20678, n20679, n20680, n20681, n20682, n20683, n20684,
         n20685, n20686, n20687, n20688, n20689, n20690, n20691, n20692,
         n20693, n20694, n20695, n20696, n20697, n20698, n20699, n20700,
         n20701, n20702, n20703, n20704, n20705, n20706, n20707, n20708,
         n20709, n20710, n20711, n20712, n20713, n20714, n20715, n20716,
         n20717, n20718, n20719, n20720, n20721, n20722, n20723, n20724,
         n20725, n20726, n20727, n20728, n20729, n20730, n20731, n20732,
         n20733, n20734, n20735, n20736, n20737, n20738, n20739, n20740,
         n20741, n20742, n20743, n20744, n20745, n20746, n20747, n20748,
         n20749, n20750, n20751, n20752, n20753, n20754, n20755, n20756,
         n20757, n20758, n20759, n20760, n20761, n20762, n20763, n20764,
         n20765, n20766, n20767, n20768, n20769, n20770, n20771, n20772,
         n20773, n20774, n20775, n20776, n20777, n20778, n20779, n20780,
         n20781, n20782, n20783, n20784, n20785, n20786, n20787, n20788,
         n20789, n20790, n20791, n20792, n20793, n20794, n20795, n20796,
         n20797, n20798, n20799, n20800, n20801, n20802, n20803, n20804,
         n20805, n20806, n20807, n20808, n20809, n20810, n20811, n20812,
         n20813, n20814, n20815, n20816, n20817, n20818, n20819, n20820,
         n20821, n20822, n20823, n20824, n20825, n20826, n20827, n20828,
         n20829, n20830, n20831, n20832, n20833, n20834, n20835, n20836,
         n20837, n20838, n20839, n20840, n20841, n20842, n20843, n20844,
         n20845, n20846, n20847, n20848, n20849, n20850, n20851, n20852,
         n20853, n20854, n20855, n20856, n20857, n20858, n20859, n20860,
         n20861, n20862, n20863, n20864, n20865, n20866, n20867, n20868,
         n20869, n20870, n20871, n20872, n20873, n20874, n20875, n20876,
         n20877, n20878, n20879, n20880, n20881, n20882, n20883, n20884,
         n20885, n20886, n20887, n20888, n20889, n20890, n20891, n20892,
         n20893, n20894, n20895, n20896, n20897, n20898, n20899, n20900,
         n20901, n20902, n20903, n20904, n20905, n20906, n20907, n20908,
         n20909, n20910, n20911, n20912, n20913, n20914, n20915, n20916,
         n20917, n20918, n20919, n20920, n20921, n20922, n20923, n20924,
         n20925, n20926, n20927, n20928, n20929, n20930, n20931, n20932,
         n20933, n20934, n20935, n20936, n20937, n20938, n20939, n20940,
         n20941, n20942, n20943, n20944, n20945, n20946, n20947, n20948,
         n20949, n20950, n20951, n20952, n20953, n20954, n20955, n20956,
         n20957, n20958, n20959, n20960, n20961, n20962, n20963, n20964,
         n20965, n20966, n20967, n20968, n20969, n20970, n20971, n20972,
         n20973, n20974, n20975, n20976, n20977, n20978, n20979, n20980,
         n20981, n20982, n20983, n20984, n20985, n20986, n20987, n20988,
         n20989, n20990, n20991, n20992, n20993, n20994, n20995, n20996,
         n20997, n20998, n20999, n21000, n21001, n21002, n21003, n21004,
         n21005, n21006, n21007, n21008, n21009, n21010, n21011, n21012,
         n21013, n21014, n21015, n21016, n21017, n21018, n21019, n21020,
         n21021, n21022, n21023, n21024, n21025, n21026, n21027, n21028,
         n21029, n21030, n21031, n21032, n21033, n21034, n21035, n21036,
         n21037, n21038, n21039, n21040, n21041, n21042, n21043, n21044,
         n21045, n21046, n21047, n21048, n21049, n21050, n21051, n21052,
         n21053, n21054, n21055, n21056, n21057, n21058, n21059, n21060,
         n21061, n21062, n21063, n21064, n21065, n21066, n21067, n21068,
         n21069, n21070, n21071, n21072, n21073, n21074, n21075, n21076,
         n21077, n21078, n21079, n21080, n21081, n21082, n21083, n21084,
         n21085, n21086, n21087, n21088, n21089, n21090, n21091, n21092,
         n21093, n21094, n21095, n21096, n21097, n21098, n21099, n21100,
         n21101, n21102, n21103, n21104, n21105, n21106, n21107, n21108,
         n21109, n21110, n21111, n21112, n21113, n21114, n21115, n21116,
         n21117, n21118, n21119, n21120, n21121, n21122, n21123, n21124,
         n21125, n21126, n21127, n21128, n21129, n21130, n21131, n21132,
         n21133, n21134, n21135, n21136, n21137, n21138, n21139, n21140,
         n21141, n21142, n21143;

  NAND2_X1 U11215 ( .A1(n17591), .A2(n17500), .ZN(n17775) );
  AOI21_X1 U11216 ( .B1(n15637), .B2(n18611), .A(n15636), .ZN(n17155) );
  INV_X2 U11217 ( .A(n14665), .ZN(n18873) );
  NOR3_X1 U11218 ( .A1(n15552), .A2(n15550), .A3(n17156), .ZN(n12024) );
  CLKBUF_X2 U11219 ( .A(n12313), .Z(n9829) );
  OR2_X1 U11220 ( .A1(n11348), .A2(n11349), .ZN(n11350) );
  INV_X2 U11221 ( .A(n17072), .ZN(n17049) );
  AND2_X1 U11222 ( .A1(n9819), .A2(n10330), .ZN(n12443) );
  AND2_X1 U11223 ( .A1(n12622), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10850) );
  AND2_X1 U11224 ( .A1(n10391), .A2(n10330), .ZN(n10789) );
  AND2_X1 U11225 ( .A1(n10271), .A2(n10384), .ZN(n12449) );
  AND2_X1 U11226 ( .A1(n12612), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10754) );
  INV_X1 U11227 ( .A(n16983), .ZN(n17101) );
  INV_X4 U11228 ( .A(n11820), .ZN(n17070) );
  CLKBUF_X3 U11229 ( .A(n14922), .Z(n9775) );
  INV_X1 U11230 ( .A(n10513), .ZN(n10537) );
  BUF_X1 U11231 ( .A(n11210), .Z(n12921) );
  CLKBUF_X2 U11232 ( .A(n11231), .Z(n13090) );
  CLKBUF_X1 U11233 ( .A(n9788), .Z(n20136) );
  CLKBUF_X3 U11234 ( .A(n10534), .Z(n9776) );
  BUF_X1 U11237 ( .A(n10353), .Z(n12305) );
  AND2_X1 U11238 ( .A1(n13541), .A2(n13446), .ZN(n11201) );
  CLKBUF_X1 U11239 ( .A(n18449), .Z(n9770) );
  NOR2_X1 U11240 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18427), .ZN(
        n18449) );
  CLKBUF_X2 U11241 ( .A(n11239), .Z(n13128) );
  NOR2_X1 U11242 ( .A1(n10535), .A2(n9776), .ZN(n10536) );
  NOR2_X2 U11243 ( .A1(n11692), .A2(n13276), .ZN(n11623) );
  NOR2_X1 U11244 ( .A1(n10482), .A2(n10353), .ZN(n10477) );
  NAND2_X1 U11245 ( .A1(n10537), .A2(n10536), .ZN(n14922) );
  AND2_X2 U11246 ( .A1(n12615), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12448) );
  NAND2_X1 U11247 ( .A1(n11084), .A2(n14886), .ZN(n11089) );
  AND2_X1 U11248 ( .A1(n12469), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10653) );
  NOR2_X1 U11249 ( .A1(n18140), .A2(n12020), .ZN(n12045) );
  NAND2_X1 U11250 ( .A1(n20113), .A2(n9823), .ZN(n11624) );
  INV_X2 U11251 ( .A(n16987), .ZN(n17110) );
  INV_X1 U11252 ( .A(n18130), .ZN(n15550) );
  AND2_X1 U11253 ( .A1(n11581), .A2(n11580), .ZN(n13466) );
  NOR3_X1 U11254 ( .A1(n14711), .A2(n14701), .A3(n9895), .ZN(n10065) );
  INV_X1 U11255 ( .A(n11060), .ZN(n10849) );
  INV_X1 U11257 ( .A(n18072), .ZN(n18551) );
  INV_X1 U11258 ( .A(n17847), .ZN(n18589) );
  NAND4_X1 U11259 ( .A1(n12019), .A2(n18135), .A3(n12024), .A4(n17308), .ZN(
        n17346) );
  NAND2_X1 U11260 ( .A1(n14045), .A2(n14047), .ZN(n14046) );
  BUF_X1 U11261 ( .A(n12304), .Z(n13480) );
  AOI22_X1 U11262 ( .A1(n14970), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B1(
        n14959), .B2(n14958), .ZN(n14962) );
  AOI21_X1 U11263 ( .B1(n15260), .B2(n15026), .A(n14850), .ZN(n15016) );
  INV_X1 U11264 ( .A(n16790), .ZN(n16713) );
  INV_X2 U11265 ( .A(n10222), .ZN(n17103) );
  INV_X1 U11266 ( .A(n17780), .ZN(n17768) );
  INV_X1 U11267 ( .A(n18563), .ZN(n18587) );
  INV_X1 U11268 ( .A(n19891), .ZN(n19957) );
  NAND2_X1 U11269 ( .A1(n15016), .A2(n15015), .ZN(n15014) );
  INV_X1 U11270 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n19796) );
  NOR2_X2 U11271 ( .A1(n17155), .A2(n17379), .ZN(n17304) );
  NAND2_X1 U11272 ( .A1(n12048), .A2(n18760), .ZN(n17784) );
  AND2_X1 U11273 ( .A1(n9912), .A2(n9911), .ZN(n9771) );
  AND2_X2 U11274 ( .A1(n9833), .A2(n11219), .ZN(n9772) );
  XOR2_X1 U11275 ( .A(n11275), .B(n11342), .Z(n9773) );
  BUF_X4 U11276 ( .A(n11624), .Z(n13276) );
  XNOR2_X2 U11277 ( .A(n10681), .B(n10682), .ZN(n13851) );
  NAND2_X2 U11278 ( .A1(n11490), .A2(n11489), .ZN(n15781) );
  NOR2_X2 U11279 ( .A1(n13860), .A2(n13862), .ZN(n13861) );
  NAND2_X2 U11280 ( .A1(n16085), .A2(n14846), .ZN(n10101) );
  NAND2_X2 U11281 ( .A1(n12321), .A2(n12320), .ZN(n12327) );
  NAND2_X2 U11282 ( .A1(n11502), .A2(n15782), .ZN(n13923) );
  NAND2_X1 U11283 ( .A1(n11122), .A2(n14886), .ZN(n12129) );
  AND2_X2 U11284 ( .A1(n13439), .A2(n11259), .ZN(n9782) );
  BUF_X1 U11285 ( .A(n14922), .Z(n9774) );
  NOR2_X2 U11287 ( .A1(n17680), .A2(n17895), .ZN(n17587) );
  NAND2_X4 U11288 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n11786), .ZN(
        n16987) );
  INV_X2 U11289 ( .A(n9829), .ZN(n10599) );
  OR2_X4 U11290 ( .A1(n11146), .A2(n11147), .ZN(n11251) );
  NOR2_X2 U11291 ( .A1(n14333), .A2(n14325), .ZN(n10181) );
  NOR2_X2 U11292 ( .A1(n12107), .A2(n16098), .ZN(n12109) );
  AND3_X2 U11293 ( .A1(n11175), .A2(n11173), .A3(n9798), .ZN(n11187) );
  INV_X4 U11294 ( .A(n11821), .ZN(n17092) );
  INV_X2 U11295 ( .A(n9822), .ZN(n11266) );
  NAND4_X4 U11296 ( .A1(n11209), .A2(n11208), .A3(n11207), .A4(n11206), .ZN(
        n9822) );
  AND2_X4 U11297 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15390) );
  INV_X4 U11298 ( .A(n12421), .ZN(n12615) );
  OR2_X4 U11299 ( .A1(n18576), .A2(n11788), .ZN(n10222) );
  NOR2_X4 U11301 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11140) );
  INV_X4 U11303 ( .A(n12424), .ZN(n10392) );
  AOI21_X2 U11304 ( .B1(n15060), .B2(n9957), .A(n9955), .ZN(n15261) );
  NOR2_X1 U11305 ( .A1(n11766), .A2(n11768), .ZN(n12287) );
  NAND2_X1 U11306 ( .A1(n9812), .A2(n14438), .ZN(n11766) );
  AND2_X1 U11307 ( .A1(n9918), .A2(n9916), .ZN(n15291) );
  CLKBUF_X1 U11308 ( .A(n16107), .Z(n9797) );
  NOR2_X1 U11309 ( .A1(n10128), .A2(n14754), .ZN(n15133) );
  OR2_X1 U11310 ( .A1(n14678), .A2(n12215), .ZN(n14926) );
  NOR3_X2 U11311 ( .A1(n14780), .A2(n10126), .A3(n12168), .ZN(n14754) );
  AND2_X1 U11312 ( .A1(n10727), .A2(n11048), .ZN(n13881) );
  INV_X1 U11313 ( .A(n17164), .ZN(n17160) );
  NOR2_X1 U11314 ( .A1(n9809), .A2(n10729), .ZN(n10083) );
  NOR2_X1 U11316 ( .A1(n12255), .A2(n12256), .ZN(n10081) );
  NOR2_X2 U11317 ( .A1(n17369), .A2(n17182), .ZN(n17178) );
  INV_X1 U11318 ( .A(n17775), .ZN(n17765) );
  NAND2_X1 U11320 ( .A1(P3_EAX_REG_25__SCAN_IN), .A2(n17183), .ZN(n17182) );
  AND2_X1 U11321 ( .A1(n10097), .A2(n15229), .ZN(n10096) );
  NAND2_X1 U11322 ( .A1(n17567), .A2(n17628), .ZN(n17536) );
  AND2_X1 U11323 ( .A1(n14189), .A2(n10060), .ZN(n14026) );
  OR2_X1 U11324 ( .A1(n11462), .A2(n10154), .ZN(n11494) );
  NOR2_X1 U11325 ( .A1(n10605), .A2(n10616), .ZN(n10731) );
  NAND2_X1 U11326 ( .A1(n11410), .A2(n11409), .ZN(n20252) );
  NOR2_X2 U11327 ( .A1(n17115), .A2(n15432), .ZN(n17001) );
  NAND2_X1 U11328 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(n17304), .ZN(n17302) );
  NOR2_X2 U11330 ( .A1(n17984), .A2(n18587), .ZN(n18008) );
  NAND2_X1 U11331 ( .A1(n11348), .A2(n11349), .ZN(n11391) );
  NOR2_X1 U11332 ( .A1(n15639), .A2(n17155), .ZN(n17300) );
  AND2_X1 U11333 ( .A1(n11089), .A2(n10106), .ZN(n11119) );
  AND2_X1 U11334 ( .A1(n11089), .A2(n10105), .ZN(n11110) );
  AOI21_X2 U11335 ( .B1(n18570), .B2(n18562), .A(n18569), .ZN(n18563) );
  NOR2_X1 U11336 ( .A1(n18117), .A2(n17409), .ZN(n17402) );
  AND2_X1 U11337 ( .A1(n12096), .A2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12123) );
  XNOR2_X1 U11338 ( .A(n10826), .B(n10825), .ZN(n13382) );
  CLKBUF_X1 U11339 ( .A(n10546), .Z(n15397) );
  OR2_X1 U11340 ( .A1(n13698), .A2(n11624), .ZN(n11259) );
  INV_X2 U11341 ( .A(n10951), .ZN(n10125) );
  NAND2_X1 U11342 ( .A1(n11397), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11577) );
  INV_X1 U11343 ( .A(n10539), .ZN(n13348) );
  CLKBUF_X2 U11345 ( .A(n11013), .Z(n14912) );
  AND2_X2 U11346 ( .A1(n9779), .A2(n19796), .ZN(n10820) );
  CLKBUF_X2 U11347 ( .A(n11288), .Z(n20127) );
  INV_X1 U11348 ( .A(n10814), .ZN(n10124) );
  NAND3_X1 U11350 ( .A1(n10352), .A2(n10477), .A3(n10351), .ZN(n10513) );
  CLKBUF_X3 U11351 ( .A(n10399), .Z(n9779) );
  NAND2_X1 U11352 ( .A1(n10350), .A2(n10349), .ZN(n10399) );
  INV_X2 U11353 ( .A(n20081), .ZN(n11744) );
  CLKBUF_X2 U11354 ( .A(n11234), .Z(n12978) );
  BUF_X2 U11355 ( .A(n11233), .Z(n12867) );
  BUF_X2 U11356 ( .A(n11232), .Z(n12937) );
  INV_X4 U11357 ( .A(n15492), .ZN(n17095) );
  BUF_X2 U11358 ( .A(n11241), .Z(n13050) );
  CLKBUF_X2 U11359 ( .A(n11201), .Z(n12965) );
  CLKBUF_X2 U11360 ( .A(n11441), .Z(n13540) );
  INV_X4 U11361 ( .A(n11799), .ZN(n17074) );
  INV_X1 U11362 ( .A(n12432), .ZN(n9777) );
  BUF_X2 U11363 ( .A(n11237), .Z(n12964) );
  BUF_X2 U11364 ( .A(n11238), .Z(n13134) );
  AND2_X1 U11365 ( .A1(n11133), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11138) );
  INV_X1 U11366 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n19836) );
  INV_X4 U11367 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10330) );
  NAND2_X1 U11369 ( .A1(n10151), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14971) );
  INV_X1 U11370 ( .A(n14980), .ZN(n10151) );
  AOI21_X1 U11371 ( .B1(n13977), .B2(n20038), .A(n13974), .ZN(n13975) );
  AND2_X1 U11372 ( .A1(n13178), .A2(n13177), .ZN(n13179) );
  NAND2_X1 U11373 ( .A1(n14999), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14980) );
  XNOR2_X1 U11374 ( .A(n13964), .B(n13963), .ZN(n13977) );
  OR2_X1 U11375 ( .A1(n15650), .A2(n20094), .ZN(n13178) );
  NOR2_X1 U11376 ( .A1(n15261), .A2(n15262), .ZN(n15260) );
  NOR2_X1 U11377 ( .A1(n14333), .A2(n14476), .ZN(n14344) );
  XNOR2_X1 U11378 ( .A(n13995), .B(n13150), .ZN(n14307) );
  NAND2_X1 U11379 ( .A1(n14006), .A2(n14156), .ZN(n14152) );
  OAI21_X1 U11380 ( .B1(n14996), .B2(n20991), .A(n14997), .ZN(n14877) );
  AND2_X1 U11381 ( .A1(n11102), .A2(n15068), .ZN(n16075) );
  OR2_X1 U11382 ( .A1(n15083), .A2(n10805), .ZN(n16081) );
  AND2_X1 U11383 ( .A1(n12221), .A2(n12220), .ZN(n10025) );
  NAND2_X1 U11384 ( .A1(n10092), .A2(n9977), .ZN(n16085) );
  NAND2_X1 U11385 ( .A1(n11059), .A2(n9837), .ZN(n10092) );
  AOI211_X1 U11386 ( .C1(n15133), .C2(n16181), .A(n15132), .B(n15131), .ZN(
        n15136) );
  OAI21_X1 U11387 ( .B1(n10065), .B2(n12216), .A(n14926), .ZN(n15137) );
  AND2_X1 U11388 ( .A1(n10159), .A2(n9888), .ZN(n14057) );
  AOI21_X1 U11389 ( .B1(n14142), .B2(n20063), .A(n10056), .ZN(n12303) );
  NOR2_X1 U11390 ( .A1(n10069), .A2(n10068), .ZN(n14691) );
  OR2_X1 U11391 ( .A1(n12298), .A2(n10057), .ZN(n10056) );
  AOI211_X1 U11392 ( .C1(n15116), .C2(n16181), .A(n15115), .B(n15114), .ZN(
        n15126) );
  INV_X1 U11393 ( .A(n14774), .ZN(n15159) );
  AOI21_X1 U11394 ( .B1(n10201), .B2(n10196), .A(n10195), .ZN(n10194) );
  AND2_X1 U11395 ( .A1(n16272), .A2(n15564), .ZN(n11920) );
  OR2_X1 U11396 ( .A1(n10801), .A2(n10849), .ZN(n10802) );
  OR2_X1 U11397 ( .A1(n10083), .A2(n10768), .ZN(n10082) );
  NOR2_X1 U11398 ( .A1(n14708), .A2(n14709), .ZN(n12201) );
  NOR2_X1 U11399 ( .A1(n17442), .A2(n11912), .ZN(n11913) );
  INV_X1 U11400 ( .A(n16854), .ZN(n16859) );
  OR2_X1 U11401 ( .A1(n11911), .A2(n10220), .ZN(n11912) );
  AND2_X1 U11402 ( .A1(n14397), .A2(n14406), .ZN(n14511) );
  AND2_X1 U11403 ( .A1(n14420), .A2(n14417), .ZN(n14406) );
  AND2_X2 U11404 ( .A1(n19924), .A2(n13216), .ZN(n19891) );
  NOR2_X1 U11405 ( .A1(n17465), .A2(n16254), .ZN(n17791) );
  AND2_X1 U11406 ( .A1(n11486), .A2(n11485), .ZN(n15788) );
  NOR2_X1 U11407 ( .A1(n14500), .A2(n14379), .ZN(n15803) );
  AND2_X1 U11408 ( .A1(n11752), .A2(n15873), .ZN(n15798) );
  NAND2_X1 U11409 ( .A1(n11524), .A2(n9901), .ZN(n14397) );
  INV_X1 U11410 ( .A(n10669), .ZN(n9912) );
  AND2_X1 U11411 ( .A1(n14352), .A2(n11510), .ZN(n13924) );
  AND2_X1 U11412 ( .A1(n10100), .A2(n10099), .ZN(n10098) );
  NOR2_X1 U11413 ( .A1(n15051), .A2(n9875), .ZN(n15018) );
  XNOR2_X1 U11414 ( .A(n11494), .B(n11493), .ZN(n12720) );
  AND2_X1 U11415 ( .A1(n10726), .A2(n10725), .ZN(n10728) );
  INV_X1 U11416 ( .A(n17189), .ZN(n17183) );
  NAND2_X1 U11417 ( .A1(n17536), .A2(n11909), .ZN(n17476) );
  AND2_X1 U11418 ( .A1(n14862), .A2(n10103), .ZN(n10100) );
  INV_X1 U11419 ( .A(n17608), .ZN(n17974) );
  OR2_X1 U11420 ( .A1(n11462), .A2(n10153), .ZN(n11481) );
  NAND2_X1 U11421 ( .A1(n10206), .A2(n9838), .ZN(n13572) );
  NAND2_X1 U11422 ( .A1(n12084), .A2(n17681), .ZN(n17608) );
  NOR2_X1 U11423 ( .A1(n14748), .A2(n14747), .ZN(n15049) );
  NAND2_X1 U11424 ( .A1(n9948), .A2(n9947), .ZN(n11462) );
  NAND2_X1 U11425 ( .A1(n12336), .A2(n12335), .ZN(n10206) );
  XNOR2_X1 U11426 ( .A(n13476), .B(n14612), .ZN(n19788) );
  XNOR2_X1 U11427 ( .A(n11419), .B(n20252), .ZN(n20763) );
  NOR2_X1 U11428 ( .A1(n14061), .A2(n14048), .ZN(n14187) );
  AND2_X1 U11429 ( .A1(n11742), .A2(n14504), .ZN(n15872) );
  OAI21_X1 U11430 ( .B1(n17639), .B2(n11904), .A(n17628), .ZN(n11905) );
  INV_X1 U11431 ( .A(n19153), .ZN(n10698) );
  NOR2_X2 U11432 ( .A1(n13967), .A2(n20092), .ZN(n13968) );
  NAND2_X1 U11433 ( .A1(n10625), .A2(n14672), .ZN(n10746) );
  NOR2_X1 U11434 ( .A1(n9952), .A2(n10606), .ZN(n10732) );
  OR2_X1 U11435 ( .A1(n9952), .A2(n10616), .ZN(n10687) );
  NOR2_X2 U11436 ( .A1(n9952), .A2(n10618), .ZN(n10733) );
  OR2_X1 U11437 ( .A1(n15573), .A2(n10849), .ZN(n14867) );
  AND2_X1 U11438 ( .A1(n13488), .A2(n10071), .ZN(n15308) );
  NAND2_X1 U11439 ( .A1(n11746), .A2(n13950), .ZN(n14504) );
  NAND2_X1 U11440 ( .A1(n11746), .A2(n13445), .ZN(n20080) );
  OR3_X1 U11441 ( .A1(n10622), .A2(n10599), .A3(n15395), .ZN(n10701) );
  NAND2_X1 U11442 ( .A1(n13480), .A2(n10619), .ZN(n19473) );
  AND2_X1 U11443 ( .A1(n13480), .A2(n10615), .ZN(n19539) );
  AND2_X1 U11444 ( .A1(n20252), .A2(n11440), .ZN(n9947) );
  AND2_X1 U11445 ( .A1(n13480), .A2(n10613), .ZN(n19638) );
  AND2_X1 U11446 ( .A1(n13480), .A2(n10617), .ZN(n19418) );
  NOR2_X1 U11447 ( .A1(n10605), .A2(n10606), .ZN(n19317) );
  NAND2_X1 U11448 ( .A1(n10600), .A2(n10599), .ZN(n9952) );
  NAND2_X1 U11449 ( .A1(n10600), .A2(n9829), .ZN(n10605) );
  NAND2_X1 U11450 ( .A1(n12310), .A2(n12309), .ZN(n13478) );
  NAND2_X1 U11451 ( .A1(n20760), .A2(n20098), .ZN(n11410) );
  INV_X2 U11452 ( .A(n13650), .ZN(n9778) );
  NAND2_X1 U11453 ( .A1(n12078), .A2(n17715), .ZN(n17705) );
  XNOR2_X1 U11454 ( .A(n11391), .B(n20254), .ZN(n20760) );
  XNOR2_X1 U11455 ( .A(n11901), .B(n11900), .ZN(n17700) );
  AND2_X1 U11456 ( .A1(n11104), .A2(n11111), .ZN(n14574) );
  INV_X1 U11457 ( .A(n13466), .ZN(n13423) );
  INV_X1 U11458 ( .A(n15395), .ZN(n14672) );
  NOR2_X2 U11459 ( .A1(n19092), .A2(n19268), .ZN(n13777) );
  NOR2_X2 U11460 ( .A1(n19161), .A2(n19268), .ZN(n19162) );
  NAND2_X1 U11461 ( .A1(n10594), .A2(n10591), .ZN(n15395) );
  AND2_X1 U11462 ( .A1(n13897), .A2(n13896), .ZN(n15884) );
  AOI21_X1 U11463 ( .B1(n11895), .B2(n10013), .A(n10012), .ZN(n10011) );
  AND2_X1 U11464 ( .A1(n10574), .A2(n10573), .ZN(n10587) );
  NOR2_X1 U11465 ( .A1(n13875), .A2(n13874), .ZN(n13897) );
  AND2_X1 U11466 ( .A1(n10971), .A2(n10585), .ZN(n10973) );
  XNOR2_X1 U11467 ( .A(n11302), .B(n11301), .ZN(n12672) );
  OR2_X1 U11468 ( .A1(n10572), .A2(n10571), .ZN(n10574) );
  AOI21_X1 U11469 ( .B1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n20098), .A(
        n11575), .ZN(n11576) );
  OR2_X1 U11470 ( .A1(n10584), .A2(n10583), .ZN(n10971) );
  NOR2_X1 U11471 ( .A1(n11085), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n11090) );
  OAI211_X1 U11472 ( .C1(n10582), .C2(n21127), .A(n10581), .B(n10580), .ZN(
        n10583) );
  NAND3_X1 U11473 ( .A1(n10223), .A2(n10558), .A3(n10221), .ZN(n10595) );
  OR2_X2 U11474 ( .A1(n17345), .A2(n18613), .ZN(n17412) );
  NOR2_X2 U11475 ( .A1(n13736), .A2(n13735), .ZN(n13740) );
  CLKBUF_X1 U11476 ( .A(n10579), .Z(n14924) );
  NOR2_X1 U11477 ( .A1(n15428), .A2(n15427), .ZN(n15536) );
  INV_X2 U11478 ( .A(n10579), .ZN(n10582) );
  NOR2_X2 U11479 ( .A1(n17274), .A2(n11867), .ZN(n17694) );
  AND2_X1 U11480 ( .A1(n10533), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9826) );
  AND2_X1 U11481 ( .A1(n10518), .A2(n10517), .ZN(n10554) );
  NAND2_X1 U11482 ( .A1(n10815), .A2(n10123), .ZN(n13504) );
  AND4_X1 U11483 ( .A1(n10553), .A2(n10552), .A3(n10551), .A4(n10550), .ZN(
        n10223) );
  NOR2_X1 U11484 ( .A1(n9846), .A2(n12091), .ZN(n12120) );
  NAND2_X1 U11485 ( .A1(n17761), .A2(n11883), .ZN(n11885) );
  NAND2_X1 U11486 ( .A1(n10532), .A2(n10953), .ZN(n15416) );
  AND2_X1 U11487 ( .A1(n11025), .A2(n11019), .ZN(n11042) );
  AND2_X1 U11488 ( .A1(n15544), .A2(n10527), .ZN(n10532) );
  NOR2_X1 U11489 ( .A1(n11279), .A2(n13545), .ZN(n11270) );
  NAND2_X1 U11490 ( .A1(n17291), .A2(n12034), .ZN(n12044) );
  NOR2_X1 U11491 ( .A1(n11026), .A2(n11027), .ZN(n11025) );
  NAND2_X1 U11492 ( .A1(n12115), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12117) );
  AND2_X1 U11493 ( .A1(n12114), .A2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n12115) );
  AND2_X1 U11494 ( .A1(n14222), .A2(n11269), .ZN(n13153) );
  NAND2_X1 U11495 ( .A1(n10537), .A2(n16218), .ZN(n10953) );
  AND2_X1 U11496 ( .A1(n11720), .A2(n11721), .ZN(n11268) );
  AND2_X1 U11497 ( .A1(n10555), .A2(n19841), .ZN(n10521) );
  AND2_X1 U11499 ( .A1(n10538), .A2(n10524), .ZN(n12633) );
  MUX2_X1 U11500 ( .A(n11016), .B(P2_EBX_REG_2__SCAN_IN), .S(n14912), .Z(
        n11027) );
  NAND2_X1 U11501 ( .A1(n11722), .A2(n11709), .ZN(n13440) );
  INV_X2 U11502 ( .A(n12167), .ZN(n12156) );
  AND2_X1 U11503 ( .A1(n11724), .A2(n11264), .ZN(n11282) );
  NOR2_X2 U11504 ( .A1(n11397), .A2(n20098), .ZN(n11571) );
  INV_X1 U11505 ( .A(n9795), .ZN(n11722) );
  NOR2_X1 U11506 ( .A1(n12112), .A2(n18882), .ZN(n12114) );
  AOI211_X2 U11507 ( .C1(n17083), .C2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A(
        n11797), .B(n11796), .ZN(n17274) );
  NAND2_X1 U11508 ( .A1(n10479), .A2(n10523), .ZN(n10495) );
  CLKBUF_X1 U11509 ( .A(n11261), .Z(n14548) );
  NAND2_X2 U11510 ( .A1(n10369), .A2(n10368), .ZN(n15544) );
  NAND2_X1 U11511 ( .A1(n10809), .A2(n10822), .ZN(n12167) );
  AOI211_X2 U11512 ( .C1(n17053), .C2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A(
        n12008), .B(n12007), .ZN(n18130) );
  NOR2_X1 U11513 ( .A1(n16218), .A2(n19836), .ZN(n19841) );
  INV_X1 U11514 ( .A(n10535), .ZN(n19845) );
  NAND2_X1 U11515 ( .A1(n10534), .A2(n10476), .ZN(n10523) );
  AND3_X1 U11516 ( .A1(n11879), .A2(n10228), .A3(n11878), .ZN(n10241) );
  NAND2_X1 U11517 ( .A1(n11828), .A2(n10015), .ZN(n17293) );
  NAND2_X1 U11518 ( .A1(n10399), .A2(n10441), .ZN(n10479) );
  CLKBUF_X3 U11519 ( .A(n10482), .Z(n10808) );
  AND4_X1 U11520 ( .A1(n11841), .A2(n11840), .A3(n11839), .A4(n11838), .ZN(
        n10226) );
  INV_X1 U11521 ( .A(n10399), .ZN(n10534) );
  AND2_X1 U11522 ( .A1(n12109), .A2(n10038), .ZN(n12099) );
  INV_X2 U11523 ( .A(n16322), .ZN(n16373) );
  INV_X1 U11524 ( .A(n10371), .ZN(n10496) );
  NAND2_X1 U11525 ( .A1(n10338), .A2(n10337), .ZN(n13807) );
  NAND2_X2 U11526 ( .A1(n10143), .A2(n10141), .ZN(n10482) );
  NAND2_X2 U11527 ( .A1(n10313), .A2(n10312), .ZN(n10480) );
  INV_X2 U11528 ( .A(n18428), .ZN(n18497) );
  NAND2_X1 U11529 ( .A1(n10366), .A2(n10365), .ZN(n10441) );
  NOR2_X1 U11530 ( .A1(n11153), .A2(n11152), .ZN(n11159) );
  BUF_X4 U11531 ( .A(n10417), .Z(n12401) );
  AND4_X1 U11532 ( .A1(n11214), .A2(n11213), .A3(n11212), .A4(n11211), .ZN(
        n9833) );
  AND4_X1 U11533 ( .A1(n11172), .A2(n11171), .A3(n11170), .A4(n11169), .ZN(
        n11188) );
  NAND2_X1 U11534 ( .A1(n10046), .A2(n10045), .ZN(n12107) );
  AND4_X1 U11535 ( .A1(n11200), .A2(n11199), .A3(n11198), .A4(n11197), .ZN(
        n11207) );
  AND4_X1 U11536 ( .A1(n11167), .A2(n11166), .A3(n11165), .A4(n11164), .ZN(
        n11168) );
  AND4_X1 U11537 ( .A1(n11180), .A2(n11179), .A3(n11178), .A4(n11177), .ZN(
        n11186) );
  AND4_X1 U11538 ( .A1(n11196), .A2(n11195), .A3(n11194), .A4(n11193), .ZN(
        n11208) );
  AND4_X1 U11539 ( .A1(n11157), .A2(n11156), .A3(n11155), .A4(n11154), .ZN(
        n11158) );
  AND4_X1 U11540 ( .A1(n11184), .A2(n11183), .A3(n11182), .A4(n11181), .ZN(
        n11185) );
  INV_X1 U11541 ( .A(n16970), .ZN(n17053) );
  AND4_X1 U11542 ( .A1(n11205), .A2(n11204), .A3(n11203), .A4(n11202), .ZN(
        n11206) );
  AND4_X1 U11543 ( .A1(n11192), .A2(n11191), .A3(n11190), .A4(n11189), .ZN(
        n11209) );
  AND2_X2 U11544 ( .A1(n10392), .A2(n10330), .ZN(n12450) );
  AND2_X1 U11545 ( .A1(n10392), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10417) );
  NAND2_X2 U11546 ( .A1(n18772), .A2(n18645), .ZN(n18703) );
  INV_X2 U11547 ( .A(n16405), .ZN(U215) );
  INV_X1 U11548 ( .A(n9847), .ZN(n17094) );
  BUF_X1 U11549 ( .A(n11464), .Z(n11398) );
  NAND2_X1 U11550 ( .A1(n12100), .A2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12104) );
  NAND2_X2 U11551 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n19773), .ZN(n19771) );
  NOR2_X1 U11552 ( .A1(n15147), .A2(n10149), .ZN(n9902) );
  INV_X2 U11553 ( .A(n11781), .ZN(n17114) );
  NOR2_X1 U11554 ( .A1(n12103), .A2(n14628), .ZN(n12100) );
  OR2_X2 U11555 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n11783), .ZN(
        n11799) );
  CLKBUF_X1 U11556 ( .A(n10385), .Z(n12432) );
  AND2_X2 U11557 ( .A1(n11138), .A2(n13446), .ZN(n11441) );
  AND2_X2 U11558 ( .A1(n9821), .A2(n10330), .ZN(n10412) );
  AND2_X2 U11559 ( .A1(n13541), .A2(n11141), .ZN(n11241) );
  OR3_X1 U11560 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(n11787), .ZN(n16966) );
  AND2_X2 U11561 ( .A1(n11139), .A2(n13546), .ZN(n11240) );
  OR2_X2 U11562 ( .A1(n11782), .A2(n16789), .ZN(n15492) );
  AND2_X2 U11563 ( .A1(n10385), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10425) );
  INV_X4 U11564 ( .A(n11811), .ZN(n16967) );
  INV_X2 U11565 ( .A(n16408), .ZN(n16410) );
  AND2_X2 U11566 ( .A1(n11130), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13541) );
  AND2_X2 U11567 ( .A1(n11131), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11141) );
  NAND3_X1 U11568 ( .A1(n15372), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10281) );
  AND2_X1 U11569 ( .A1(n10024), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11786) );
  NOR3_X1 U11570 ( .A1(n18764), .A2(n18775), .A3(P3_STATE2_REG_1__SCAN_IN), 
        .ZN(n18611) );
  NAND2_X1 U11571 ( .A1(n18732), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11789) );
  OR3_X2 U11572 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(n18576), .ZN(n16983) );
  NAND2_X2 U11573 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n18576) );
  NAND3_X1 U11574 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n15540) );
  INV_X1 U11575 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n16194) );
  INV_X1 U11576 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n9816) );
  INV_X1 U11578 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11133) );
  AND2_X2 U11579 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13546) );
  NOR2_X1 U11580 ( .A1(n14956), .A2(n14955), .ZN(n14957) );
  NAND2_X1 U11581 ( .A1(n18865), .A2(n18866), .ZN(n18864) );
  AOI22_X4 U11582 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n12093), .B1(n14927), 
        .B2(n19836), .ZN(n12116) );
  AOI21_X2 U11583 ( .B1(n14692), .B2(n14694), .A(n14693), .ZN(n14778) );
  NAND2_X1 U11584 ( .A1(n13164), .A2(n9781), .ZN(n10235) );
  INV_X1 U11585 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n9781) );
  NAND2_X1 U11586 ( .A1(n13851), .A2(n13850), .ZN(n9783) );
  INV_X1 U11587 ( .A(n12247), .ZN(n9784) );
  NAND2_X1 U11588 ( .A1(n15095), .A2(n15251), .ZN(n12249) );
  NOR2_X1 U11590 ( .A1(n14697), .A2(n14699), .ZN(n14698) );
  AOI21_X2 U11591 ( .B1(n10101), .B2(n9853), .A(n10094), .ZN(n14996) );
  NAND2_X1 U11592 ( .A1(n13439), .A2(n11259), .ZN(n9786) );
  INV_X1 U11593 ( .A(n20113), .ZN(n13529) );
  NAND2_X1 U11594 ( .A1(n9833), .A2(n11219), .ZN(n9788) );
  AND4_X1 U11595 ( .A1(n11218), .A2(n11217), .A3(n11216), .A4(n11215), .ZN(
        n11219) );
  AND4_X2 U11596 ( .A1(n11244), .A2(n11236), .A3(n11242), .A4(n11243), .ZN(
        n9836) );
  NAND2_X1 U11597 ( .A1(n11139), .A2(n11138), .ZN(n9789) );
  INV_X2 U11598 ( .A(n9789), .ZN(n11239) );
  INV_X1 U11599 ( .A(n13965), .ZN(n9790) );
  OR2_X2 U11600 ( .A1(n9799), .A2(n9800), .ZN(n11253) );
  AND2_X2 U11601 ( .A1(n11159), .A2(n11158), .ZN(n9791) );
  INV_X1 U11602 ( .A(n14971), .ZN(n9792) );
  NOR2_X1 U11603 ( .A1(n15005), .A2(n20991), .ZN(n9793) );
  AND2_X1 U11604 ( .A1(n9793), .A2(n9794), .ZN(n15149) );
  AND2_X1 U11605 ( .A1(n9902), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n9794) );
  CLKBUF_X1 U11606 ( .A(n11269), .Z(n13545) );
  NAND2_X1 U11607 ( .A1(n11258), .A2(n11257), .ZN(n13698) );
  NOR2_X2 U11608 ( .A1(n16556), .A2(n16903), .ZN(n16869) );
  NOR3_X4 U11609 ( .A1(n18117), .A2(n18114), .A3(n15635), .ZN(n17146) );
  NOR2_X2 U11610 ( .A1(n17895), .A2(n17974), .ZN(n17918) );
  NAND2_X1 U11611 ( .A1(n11263), .A2(n11251), .ZN(n9795) );
  NAND2_X1 U11612 ( .A1(n11263), .A2(n11251), .ZN(n11540) );
  AOI21_X1 U11613 ( .B1(n14222), .B2(n20136), .A(n13965), .ZN(n11724) );
  AND2_X1 U11614 ( .A1(n11245), .A2(n9791), .ZN(n11258) );
  INV_X1 U11615 ( .A(n13746), .ZN(n9796) );
  OR2_X2 U11616 ( .A1(n12567), .A2(n12566), .ZN(n12570) );
  NOR2_X2 U11617 ( .A1(n14698), .A2(n12538), .ZN(n12567) );
  OAI211_X1 U11618 ( .C1(n12858), .C2(n11282), .A(n11271), .B(n11270), .ZN(
        n11719) );
  AND2_X1 U11619 ( .A1(n11176), .A2(n11174), .ZN(n9798) );
  AND2_X2 U11620 ( .A1(n14831), .A2(n14832), .ZN(n14830) );
  NOR2_X2 U11621 ( .A1(n15268), .A2(n15269), .ZN(n14831) );
  NAND4_X1 U11622 ( .A1(n11223), .A2(n11220), .A3(n11222), .A4(n11221), .ZN(
        n9799) );
  NAND4_X1 U11623 ( .A1(n11227), .A2(n11226), .A3(n11225), .A4(n11224), .ZN(
        n9800) );
  XNOR2_X1 U11624 ( .A(n11275), .B(n11342), .ZN(n9801) );
  AND2_X2 U11625 ( .A1(n10218), .A2(n9802), .ZN(n14679) );
  NOR2_X1 U11626 ( .A1(n12594), .A2(n14680), .ZN(n9802) );
  NAND2_X1 U11627 ( .A1(n10218), .A2(n14684), .ZN(n9803) );
  NAND2_X1 U11628 ( .A1(n9910), .A2(n11344), .ZN(n11348) );
  NAND2_X1 U11629 ( .A1(n9773), .A2(n11286), .ZN(n9910) );
  NAND3_X1 U11630 ( .A1(n14394), .A2(n10202), .A3(n10198), .ZN(n10197) );
  NAND2_X1 U11631 ( .A1(n9912), .A2(n9911), .ZN(n9804) );
  NAND2_X1 U11632 ( .A1(n9912), .A2(n9911), .ZN(n9805) );
  AOI211_X1 U11633 ( .C1(n21130), .C2(n15954), .A(n15152), .B(n15151), .ZN(
        n15153) );
  CLKBUF_X1 U11634 ( .A(n10206), .Z(n9806) );
  NAND2_X1 U11635 ( .A1(n12318), .A2(n12317), .ZN(n12331) );
  NAND2_X1 U11636 ( .A1(n11584), .A2(n11254), .ZN(n11255) );
  AND2_X4 U11637 ( .A1(n13541), .A2(n13594), .ZN(n11210) );
  XNOR2_X2 U11638 ( .A(n11389), .B(n11388), .ZN(n14543) );
  OAI21_X1 U11639 ( .B1(n10237), .B2(n10633), .A(n10632), .ZN(n9807) );
  OR2_X1 U11640 ( .A1(n15154), .A2(n21140), .ZN(n9808) );
  NAND2_X1 U11641 ( .A1(n9808), .A2(n15153), .ZN(P2_U3017) );
  NAND2_X1 U11642 ( .A1(n9771), .A2(n10840), .ZN(n9809) );
  XNOR2_X1 U11643 ( .A(n10559), .B(n10560), .ZN(n9810) );
  OAI21_X1 U11644 ( .B1(n10237), .B2(n10633), .A(n10632), .ZN(n10669) );
  NAND2_X2 U11645 ( .A1(n10529), .A2(n10528), .ZN(n10559) );
  NOR2_X2 U11646 ( .A1(n17373), .A2(n17173), .ZN(n17169) );
  NOR4_X2 U11647 ( .A1(n17361), .A2(n17351), .A3(n17232), .A4(n17204), .ZN(
        n17194) );
  INV_X2 U11648 ( .A(n18145), .ZN(n17291) );
  NAND2_X1 U11649 ( .A1(n10197), .A2(n10194), .ZN(n9811) );
  AND2_X1 U11650 ( .A1(n10181), .A2(n10180), .ZN(n9812) );
  CLKBUF_X1 U11651 ( .A(n13412), .Z(n9813) );
  NAND3_X1 U11652 ( .A1(n9908), .A2(n11255), .A3(n9907), .ZN(n9814) );
  NAND2_X1 U11653 ( .A1(n10197), .A2(n10194), .ZN(n14386) );
  OAI21_X2 U11654 ( .B1(n11540), .B2(n9791), .A(n11250), .ZN(n9908) );
  XNOR2_X2 U11655 ( .A(n9909), .B(n11365), .ZN(n11389) );
  NAND2_X1 U11656 ( .A1(n12663), .A2(n12662), .ZN(n20543) );
  AOI211_X4 U11657 ( .C1(n17065), .C2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A(
        n11958), .B(n11957), .ZN(n18114) );
  NOR2_X2 U11658 ( .A1(n14046), .A2(n10161), .ZN(n14034) );
  AND2_X1 U11659 ( .A1(n10533), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10579) );
  AOI21_X2 U11660 ( .B1(n9826), .B2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n10544), .ZN(n10560) );
  INV_X2 U11661 ( .A(n10441), .ZN(n10476) );
  XNOR2_X1 U11662 ( .A(n10178), .B(n13412), .ZN(n14534) );
  NOR2_X2 U11663 ( .A1(n13616), .A2(n14589), .ZN(n13726) );
  INV_X2 U11665 ( .A(n10353), .ZN(n12311) );
  NAND2_X2 U11666 ( .A1(n10369), .A2(n10352), .ZN(n10512) );
  OR2_X1 U11667 ( .A1(n9810), .A2(n10593), .ZN(n10594) );
  AND2_X1 U11668 ( .A1(n13501), .A2(n12330), .ZN(n13496) );
  NAND2_X2 U11669 ( .A1(n10183), .A2(n10182), .ZN(n14431) );
  AND2_X1 U11670 ( .A1(n11274), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11342) );
  NAND4_X2 U11671 ( .A1(n11209), .A2(n11208), .A3(n11207), .A4(n11206), .ZN(
        n9823) );
  NOR2_X1 U11672 ( .A1(n18576), .A2(n11782), .ZN(n17096) );
  INV_X1 U11673 ( .A(n17096), .ZN(n16970) );
  AND3_X4 U11674 ( .A1(n10267), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n9818) );
  NAND2_X2 U11675 ( .A1(n11380), .A2(n11379), .ZN(n12670) );
  AND2_X4 U11676 ( .A1(n15391), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n9819) );
  AND2_X2 U11677 ( .A1(n15391), .A2(n16194), .ZN(n9820) );
  AND2_X2 U11678 ( .A1(n15391), .A2(n16194), .ZN(n9821) );
  NOR2_X2 U11679 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15401) );
  NOR2_X2 U11680 ( .A1(n15005), .A2(n20991), .ZN(n14999) );
  AOI211_X1 U11681 ( .C1(n16117), .C2(n15954), .A(n14953), .B(n14952), .ZN(
        n14954) );
  NAND2_X2 U11682 ( .A1(n13494), .A2(n12334), .ZN(n13476) );
  AND2_X2 U11683 ( .A1(n10367), .A2(n10511), .ZN(n10538) );
  NAND2_X2 U11684 ( .A1(n11597), .A2(n13529), .ZN(n13439) );
  NAND2_X2 U11685 ( .A1(n10280), .A2(n10279), .ZN(n10371) );
  AND2_X1 U11686 ( .A1(n13546), .A2(n13446), .ZN(n13028) );
  AND2_X2 U11687 ( .A1(n13546), .A2(n13446), .ZN(n9825) );
  AND2_X1 U11688 ( .A1(n13546), .A2(n13446), .ZN(n9824) );
  NAND2_X2 U11689 ( .A1(n20035), .A2(n20034), .ZN(n20033) );
  XNOR2_X2 U11690 ( .A(n11437), .B(n20061), .ZN(n20035) );
  XNOR2_X2 U11691 ( .A(n11417), .B(n20069), .ZN(n13708) );
  NAND2_X2 U11692 ( .A1(n13689), .A2(n11387), .ZN(n11417) );
  XNOR2_X2 U11693 ( .A(n11386), .B(n20090), .ZN(n13691) );
  NAND2_X2 U11694 ( .A1(n14536), .A2(n10176), .ZN(n11386) );
  NOR2_X2 U11695 ( .A1(n13572), .A2(n12339), .ZN(n19029) );
  AND2_X1 U11696 ( .A1(n13594), .A2(n11140), .ZN(n9827) );
  AND2_X1 U11697 ( .A1(n13594), .A2(n11140), .ZN(n11237) );
  NOR2_X4 U11698 ( .A1(n14020), .A2(n13027), .ZN(n14004) );
  NAND2_X2 U11699 ( .A1(n14386), .A2(n14385), .ZN(n14368) );
  AND2_X1 U11700 ( .A1(n15390), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n9828) );
  OAI21_X2 U11701 ( .B1(n14006), .B2(n14156), .A(n14152), .ZN(n15675) );
  AND2_X2 U11702 ( .A1(n14004), .A2(n13049), .ZN(n14006) );
  NAND2_X2 U11703 ( .A1(n13760), .A2(n13762), .ZN(n13761) );
  AND2_X4 U11704 ( .A1(n13594), .A2(n13546), .ZN(n11317) );
  NOR2_X4 U11705 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13594) );
  NAND2_X1 U11706 ( .A1(n10590), .A2(n9919), .ZN(n12313) );
  NOR2_X2 U11707 ( .A1(n13678), .A2(n10212), .ZN(n13760) );
  AND2_X1 U11708 ( .A1(n9779), .A2(n19796), .ZN(n9830) );
  AND2_X1 U11709 ( .A1(n9779), .A2(n19796), .ZN(n9831) );
  NOR2_X2 U11710 ( .A1(n13761), .A2(n10207), .ZN(n13909) );
  NOR2_X2 U11711 ( .A1(n14719), .A2(n14721), .ZN(n14720) );
  AND2_X2 U11713 ( .A1(n14735), .A2(n10215), .ZN(n12458) );
  NOR2_X4 U11714 ( .A1(n14733), .A2(n12385), .ZN(n14735) );
  NOR2_X2 U11715 ( .A1(n14713), .A2(n14714), .ZN(n12512) );
  NOR2_X2 U11716 ( .A1(n14720), .A2(n12460), .ZN(n14713) );
  AND2_X2 U11717 ( .A1(n10386), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10659) );
  INV_X1 U11718 ( .A(n11419), .ZN(n9948) );
  INV_X1 U11719 ( .A(n12338), .ZN(n12564) );
  NAND2_X1 U11720 ( .A1(n10170), .A2(n13049), .ZN(n10169) );
  NOR2_X1 U11721 ( .A1(n14153), .A2(n10171), .ZN(n10170) );
  INV_X1 U11722 ( .A(n14156), .ZN(n10171) );
  NAND2_X1 U11723 ( .A1(n17740), .A2(n11890), .ZN(n11893) );
  NAND2_X1 U11724 ( .A1(n19539), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n9922) );
  NAND2_X1 U11725 ( .A1(n20127), .A2(n9823), .ZN(n11397) );
  NAND2_X1 U11726 ( .A1(n10251), .A2(n10250), .ZN(n10256) );
  XNOR2_X1 U11727 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n10255) );
  AND2_X1 U11728 ( .A1(n9852), .A2(n11075), .ZN(n10115) );
  NAND2_X1 U11729 ( .A1(n12858), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13123) );
  AND2_X1 U11730 ( .A1(n12767), .A2(n13919), .ZN(n10152) );
  INV_X1 U11731 ( .A(n13199), .ZN(n12767) );
  NAND2_X1 U11732 ( .A1(n10180), .A2(n10181), .ZN(n10179) );
  NOR2_X1 U11733 ( .A1(n14099), .A2(n10055), .ZN(n10054) );
  INV_X1 U11734 ( .A(n14123), .ZN(n10055) );
  NAND2_X1 U11735 ( .A1(n13151), .A2(n11507), .ZN(n11503) );
  NAND2_X1 U11736 ( .A1(n11463), .A2(n11476), .ZN(n10154) );
  INV_X1 U11737 ( .A(n11623), .ZN(n11708) );
  AND2_X1 U11738 ( .A1(n11251), .A2(n20113), .ZN(n11541) );
  INV_X1 U11739 ( .A(n11584), .ZN(n13957) );
  AND2_X1 U11740 ( .A1(n9877), .A2(n14731), .ZN(n10111) );
  AND2_X1 U11741 ( .A1(n12537), .A2(n9900), .ZN(n12538) );
  NAND4_X1 U11742 ( .A1(n10371), .A2(n11013), .A3(n12636), .A4(n12305), .ZN(
        n10539) );
  INV_X1 U11743 ( .A(n10670), .ZN(n9911) );
  INV_X1 U11744 ( .A(n14979), .ZN(n14891) );
  INV_X1 U11745 ( .A(n14988), .ZN(n14890) );
  NOR2_X1 U11746 ( .A1(n9779), .A2(n10808), .ZN(n10809) );
  AND2_X1 U11747 ( .A1(n10808), .A2(n19796), .ZN(n10806) );
  AND2_X1 U11748 ( .A1(n11013), .A2(n10525), .ZN(n10526) );
  OR2_X1 U11749 ( .A1(n18722), .A2(n11783), .ZN(n11821) );
  XNOR2_X1 U11750 ( .A(n17293), .B(n12058), .ZN(n11882) );
  AOI21_X2 U11751 ( .B1(n16432), .B2(n10244), .A(n15538), .ZN(n15637) );
  AND2_X1 U11752 ( .A1(n19924), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13747) );
  INV_X1 U11753 ( .A(n12893), .ZN(n13961) );
  NOR2_X1 U11754 ( .A1(n10169), .A2(n10168), .ZN(n10167) );
  INV_X1 U11755 ( .A(n13170), .ZN(n10168) );
  NOR2_X2 U11756 ( .A1(n13171), .A2(n13996), .ZN(n13995) );
  INV_X1 U11757 ( .A(n14511), .ZN(n10195) );
  NOR2_X1 U11758 ( .A1(n13466), .A2(n13168), .ZN(n15598) );
  AND3_X1 U11759 ( .A1(n14148), .A2(n14147), .A3(n11769), .ZN(n12292) );
  INV_X1 U11760 ( .A(n14147), .ZN(n10051) );
  NAND2_X1 U11761 ( .A1(n14552), .A2(n20098), .ZN(n13173) );
  CLKBUF_X1 U11762 ( .A(n14543), .Z(n14544) );
  NOR2_X1 U11763 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(n14878), .ZN(n14893) );
  NAND2_X1 U11764 ( .A1(n12099), .A2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12112) );
  INV_X1 U11765 ( .A(n15092), .ZN(n10091) );
  AND4_X1 U11766 ( .A1(n10793), .A2(n10792), .A3(n10791), .A4(n10790), .ZN(
        n10794) );
  AND4_X1 U11767 ( .A1(n10780), .A2(n10779), .A3(n10778), .A4(n10777), .ZN(
        n10797) );
  AND4_X1 U11768 ( .A1(n10784), .A2(n10783), .A3(n10782), .A4(n10781), .ZN(
        n10796) );
  OR2_X1 U11769 ( .A1(n9964), .A2(n9962), .ZN(n9960) );
  NAND2_X1 U11770 ( .A1(n16790), .A2(n17493), .ZN(n9992) );
  AND2_X1 U11771 ( .A1(n9986), .A2(n16790), .ZN(n16539) );
  INV_X1 U11772 ( .A(n17114), .ZN(n17065) );
  OAI21_X1 U11773 ( .B1(n17728), .B2(n10014), .A(n10011), .ZN(n17712) );
  INV_X1 U11774 ( .A(n17714), .ZN(n10012) );
  INV_X1 U11775 ( .A(n11253), .ZN(n13965) );
  INV_X1 U11776 ( .A(n19539), .ZN(n10705) );
  NAND2_X1 U11777 ( .A1(n19418), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n9923) );
  NOR2_X1 U11778 ( .A1(n10227), .A2(n10645), .ZN(n10650) );
  OAI21_X1 U11779 ( .B1(n11522), .B2(n10200), .A(n10199), .ZN(n10204) );
  NAND2_X1 U11780 ( .A1(n11667), .A2(n10205), .ZN(n10200) );
  OAI21_X1 U11781 ( .B1(n14352), .B2(n11667), .A(n10205), .ZN(n10199) );
  CLKBUF_X1 U11782 ( .A(n13133), .Z(n13112) );
  CLKBUF_X1 U11783 ( .A(n11317), .Z(n12957) );
  AOI22_X1 U11784 ( .A1(n11239), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11238), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11151) );
  AOI22_X1 U11785 ( .A1(n11234), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11231), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11149) );
  INV_X1 U11786 ( .A(n10848), .ZN(n11052) );
  NOR2_X1 U11787 ( .A1(n17288), .A2(n11868), .ZN(n11888) );
  NOR2_X1 U11788 ( .A1(n11288), .A2(n11251), .ZN(n11245) );
  XNOR2_X1 U11789 ( .A(n11462), .B(n11463), .ZN(n12707) );
  INV_X1 U11790 ( .A(n14005), .ZN(n13049) );
  NAND2_X1 U11791 ( .A1(n10165), .A2(n12920), .ZN(n10164) );
  INV_X1 U11792 ( .A(n14178), .ZN(n10165) );
  NAND2_X1 U11793 ( .A1(n10204), .A2(n9951), .ZN(n10198) );
  OAI21_X1 U11794 ( .B1(n11522), .B2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n11524), .ZN(n9951) );
  INV_X1 U11795 ( .A(n13123), .ZN(n13143) );
  INV_X1 U11796 ( .A(n13895), .ZN(n9906) );
  INV_X1 U11797 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n21068) );
  NOR2_X2 U11798 ( .A1(n20136), .A2(n20623), .ZN(n12838) );
  AND2_X1 U11799 ( .A1(n14352), .A2(n14455), .ZN(n13161) );
  AND2_X1 U11800 ( .A1(n10063), .A2(n9898), .ZN(n10062) );
  AND2_X1 U11801 ( .A1(n14181), .A2(n10064), .ZN(n10063) );
  INV_X1 U11802 ( .A(n14491), .ZN(n10064) );
  NAND2_X1 U11803 ( .A1(n9945), .A2(n11518), .ZN(n14396) );
  AND2_X1 U11804 ( .A1(n14422), .A2(n11519), .ZN(n9945) );
  NAND2_X1 U11805 ( .A1(n13696), .A2(n11692), .ZN(n11700) );
  CLKBUF_X1 U11806 ( .A(n11629), .Z(n11696) );
  NAND2_X1 U11807 ( .A1(n11380), .A2(n11333), .ZN(n11337) );
  OAI211_X1 U11808 ( .C1(n11345), .C2(n13447), .A(n11347), .B(n11346), .ZN(
        n11349) );
  OAI22_X1 U11809 ( .A1(n11574), .A2(n11573), .B1(n11592), .B2(n11572), .ZN(
        n11575) );
  NAND2_X1 U11810 ( .A1(n11537), .A2(n11569), .ZN(n11591) );
  OR2_X1 U11811 ( .A1(n11570), .A2(n11536), .ZN(n11537) );
  AND2_X1 U11812 ( .A1(n11571), .A2(n11541), .ZN(n11579) );
  OAI21_X1 U11813 ( .B1(n20791), .B2(n15933), .A(n15613), .ZN(n20097) );
  AND2_X1 U11814 ( .A1(n10258), .A2(n10257), .ZN(n10456) );
  NOR2_X1 U11815 ( .A1(n12131), .A2(n10114), .ZN(n10113) );
  NAND2_X1 U11816 ( .A1(n10108), .A2(n11091), .ZN(n10107) );
  INV_X1 U11817 ( .A(n9893), .ZN(n10108) );
  NAND2_X1 U11818 ( .A1(n11067), .A2(n9860), .ZN(n11085) );
  INV_X1 U11819 ( .A(n10844), .ZN(n11043) );
  AND3_X1 U11820 ( .A1(n10538), .A2(n19845), .A3(n9779), .ZN(n10545) );
  NOR2_X1 U11821 ( .A1(n10074), .A2(n13584), .ZN(n10073) );
  INV_X1 U11822 ( .A(n13570), .ZN(n10074) );
  NAND2_X1 U11823 ( .A1(n14706), .A2(n12515), .ZN(n12537) );
  NAND2_X1 U11824 ( .A1(n12512), .A2(n12514), .ZN(n12515) );
  AND2_X1 U11825 ( .A1(n10216), .A2(n16021), .ZN(n10215) );
  AND2_X1 U11826 ( .A1(n10133), .A2(n10132), .ZN(n10131) );
  INV_X1 U11827 ( .A(n13914), .ZN(n10132) );
  OR2_X1 U11828 ( .A1(n10044), .A2(n12275), .ZN(n10043) );
  NAND2_X1 U11829 ( .A1(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n10044) );
  OR2_X1 U11830 ( .A1(n10048), .A2(n16113), .ZN(n10047) );
  NAND2_X1 U11831 ( .A1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n10048) );
  AND4_X1 U11832 ( .A1(n10788), .A2(n10787), .A3(n10786), .A4(n10785), .ZN(
        n10795) );
  AND2_X1 U11833 ( .A1(n15986), .A2(n11060), .ZN(n14902) );
  INV_X1 U11834 ( .A(n15008), .ZN(n10095) );
  AND2_X1 U11835 ( .A1(n10140), .A2(n10139), .ZN(n10138) );
  INV_X1 U11836 ( .A(n15234), .ZN(n10139) );
  INV_X1 U11837 ( .A(n9961), .ZN(n9959) );
  INV_X1 U11838 ( .A(n14854), .ZN(n9962) );
  NAND2_X1 U11839 ( .A1(n9924), .A2(n10680), .ZN(n10681) );
  INV_X1 U11840 ( .A(n13790), .ZN(n9925) );
  NAND2_X1 U11841 ( .A1(n10125), .A2(n10124), .ZN(n10123) );
  OAI21_X1 U11842 ( .B1(n12167), .B2(n10122), .A(n10819), .ZN(n13503) );
  AND2_X1 U11843 ( .A1(n10480), .A2(n19796), .ZN(n10822) );
  AND2_X1 U11844 ( .A1(n10492), .A2(n10480), .ZN(n10494) );
  AND2_X1 U11845 ( .A1(n10262), .A2(n10261), .ZN(n10460) );
  OR2_X1 U11846 ( .A1(n10260), .A2(n10259), .ZN(n10262) );
  NAND2_X1 U11847 ( .A1(n10142), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10141) );
  NAND2_X1 U11848 ( .A1(n10144), .A2(n10330), .ZN(n10143) );
  NAND2_X1 U11849 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n18745), .ZN(
        n11787) );
  NAND2_X1 U11850 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18722), .ZN(
        n11782) );
  AND2_X1 U11851 ( .A1(n9887), .A2(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n9998) );
  OR2_X1 U11852 ( .A1(n17694), .A2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10022) );
  NAND2_X1 U11853 ( .A1(n16416), .A2(n12026), .ZN(n15528) );
  NAND2_X1 U11854 ( .A1(n15528), .A2(n17346), .ZN(n16433) );
  OAI21_X1 U11855 ( .B1(n12041), .B2(n12043), .A(n12040), .ZN(n15527) );
  NAND2_X1 U11856 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11788) );
  AOI211_X1 U11857 ( .C1(n16967), .C2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A(
        n11996), .B(n11995), .ZN(n11997) );
  NOR2_X1 U11858 ( .A1(n12953), .A2(n14373), .ZN(n13013) );
  NOR2_X1 U11859 ( .A1(n20113), .A2(n9822), .ZN(n13744) );
  OR2_X1 U11860 ( .A1(n20785), .A2(n13204), .ZN(n19924) );
  OR2_X1 U11861 ( .A1(n13625), .A2(n13624), .ZN(n13736) );
  NOR2_X1 U11862 ( .A1(n13104), .A2(n15653), .ZN(n13105) );
  NAND2_X1 U11863 ( .A1(n13105), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13205) );
  OAI21_X1 U11864 ( .B1(n12695), .B2(n15667), .A(n13085), .ZN(n14153) );
  NAND2_X1 U11865 ( .A1(n13044), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n13045) );
  OR2_X1 U11866 ( .A1(n13045), .A2(n14337), .ZN(n13067) );
  OAI21_X1 U11867 ( .B1(n9811), .B2(n9949), .A(n11524), .ZN(n14358) );
  NAND2_X1 U11868 ( .A1(n9903), .A2(n9950), .ZN(n9949) );
  NOR2_X1 U11869 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n9950) );
  AND2_X1 U11870 ( .A1(n12956), .A2(n12955), .ZN(n14260) );
  OR2_X1 U11871 ( .A1(n15753), .A2(n12695), .ZN(n12918) );
  XNOR2_X1 U11872 ( .A(n14352), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14385) );
  INV_X1 U11873 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n14132) );
  INV_X1 U11874 ( .A(n13623), .ZN(n12679) );
  OR2_X1 U11875 ( .A1(n12292), .A2(n11709), .ZN(n12294) );
  AND2_X1 U11876 ( .A1(n11691), .A2(n11690), .ZN(n14024) );
  AND2_X1 U11877 ( .A1(n14205), .A2(n9886), .ZN(n14089) );
  INV_X1 U11878 ( .A(n14090), .ZN(n10053) );
  OR2_X1 U11879 ( .A1(n14217), .A2(n14216), .ZN(n14219) );
  AND2_X1 U11880 ( .A1(n11514), .A2(n9869), .ZN(n10182) );
  OR2_X1 U11881 ( .A1(n15886), .A2(n13213), .ZN(n14217) );
  OR2_X1 U11882 ( .A1(n15921), .A2(n13825), .ZN(n13875) );
  AND2_X1 U11883 ( .A1(n11335), .A2(n11334), .ZN(n12662) );
  NOR2_X1 U11884 ( .A1(n20422), .A2(n20259), .ZN(n20580) );
  OR2_X1 U11885 ( .A1(n20629), .A2(n20548), .ZN(n20575) );
  AND2_X1 U11886 ( .A1(n20543), .A2(n20179), .ZN(n20569) );
  AOI21_X1 U11887 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n20538), .A(n20259), 
        .ZN(n20630) );
  NAND2_X1 U11888 ( .A1(n20098), .A2(n20097), .ZN(n20259) );
  AND2_X1 U11889 ( .A1(n14896), .A2(n14564), .ZN(n14565) );
  NOR2_X1 U11890 ( .A1(n10118), .A2(n14864), .ZN(n10117) );
  NAND2_X1 U11891 ( .A1(n10120), .A2(n10119), .ZN(n10118) );
  NOR2_X1 U11892 ( .A1(P2_EBX_REG_25__SCAN_IN), .A2(P2_EBX_REG_24__SCAN_IN), 
        .ZN(n10119) );
  OR2_X1 U11893 ( .A1(n14893), .A2(n10104), .ZN(n14910) );
  OR2_X1 U11894 ( .A1(n10910), .A2(n10909), .ZN(n19015) );
  NAND2_X1 U11895 ( .A1(n13680), .A2(n12341), .ZN(n10214) );
  OR2_X1 U11896 ( .A1(n10210), .A2(n10208), .ZN(n10207) );
  INV_X1 U11897 ( .A(n13911), .ZN(n10208) );
  AND2_X1 U11898 ( .A1(n14577), .A2(n13812), .ZN(n10133) );
  AND2_X1 U11899 ( .A1(n13373), .A2(n13372), .ZN(n15377) );
  NAND3_X1 U11900 ( .A1(n10032), .A2(n10030), .A3(n10029), .ZN(n14927) );
  NAND2_X1 U11901 ( .A1(n10034), .A2(n10037), .ZN(n10029) );
  NAND2_X1 U11902 ( .A1(n12123), .A2(n10031), .ZN(n10030) );
  OR2_X1 U11903 ( .A1(n12123), .A2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n10032) );
  NAND2_X1 U11904 ( .A1(n12120), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12121) );
  AND2_X1 U11905 ( .A1(n9834), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10038) );
  NAND2_X1 U11906 ( .A1(n10147), .A2(n10145), .ZN(n16107) );
  OAI211_X1 U11907 ( .C1(n9915), .C2(n15349), .A(n9859), .B(n10776), .ZN(
        n10147) );
  INV_X1 U11908 ( .A(n10146), .ZN(n10145) );
  NAND2_X1 U11909 ( .A1(n10586), .A2(n10587), .ZN(n9919) );
  NAND2_X1 U11910 ( .A1(n10086), .A2(n10084), .ZN(n14932) );
  AOI21_X1 U11911 ( .B1(n10087), .B2(n10089), .A(n10085), .ZN(n10084) );
  INV_X1 U11912 ( .A(n14944), .ZN(n10085) );
  NAND2_X1 U11913 ( .A1(n14996), .A2(n20991), .ZN(n14876) );
  OR2_X1 U11914 ( .A1(n10102), .A2(n15230), .ZN(n10097) );
  INV_X1 U11915 ( .A(n15230), .ZN(n10099) );
  OR2_X1 U11916 ( .A1(n14867), .A2(n15241), .ZN(n15229) );
  NAND2_X1 U11917 ( .A1(n12244), .A2(n12237), .ZN(n9974) );
  INV_X1 U11918 ( .A(n12244), .ZN(n9976) );
  NOR2_X1 U11919 ( .A1(n9963), .A2(n9962), .ZN(n9961) );
  INV_X1 U11920 ( .A(n15057), .ZN(n9963) );
  NOR2_X1 U11921 ( .A1(n11117), .A2(n9965), .ZN(n9964) );
  INV_X1 U11922 ( .A(n15047), .ZN(n9965) );
  AND2_X1 U11923 ( .A1(n9835), .A2(n11088), .ZN(n9977) );
  AOI21_X1 U11924 ( .B1(n15395), .B2(n12326), .A(n12325), .ZN(n13498) );
  NAND2_X1 U11925 ( .A1(n13499), .A2(n13498), .ZN(n13501) );
  AND2_X2 U11926 ( .A1(n10485), .A2(n10525), .ZN(n10369) );
  NOR2_X1 U11927 ( .A1(n10605), .A2(n10607), .ZN(n19265) );
  NAND2_X1 U11928 ( .A1(n19788), .A2(n19817), .ZN(n19314) );
  NAND2_X1 U11929 ( .A1(n10610), .A2(n9829), .ZN(n10702) );
  NOR2_X1 U11930 ( .A1(n10622), .A2(n14672), .ZN(n10610) );
  INV_X1 U11931 ( .A(n10702), .ZN(n19605) );
  NAND2_X1 U11932 ( .A1(n10336), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10337) );
  NAND2_X1 U11933 ( .A1(n10331), .A2(n10330), .ZN(n10338) );
  OR2_X1 U11934 ( .A1(n19788), .A2(n19817), .ZN(n19537) );
  OAI21_X2 U11935 ( .B1(n16244), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n13772), 
        .ZN(n19647) );
  NOR2_X1 U11936 ( .A1(n16506), .A2(n16713), .ZN(n16499) );
  OR2_X1 U11937 ( .A1(n16499), .A2(n17449), .ZN(n9981) );
  AND2_X1 U11939 ( .A1(n9991), .A2(n9989), .ZN(n16521) );
  NOR2_X1 U11940 ( .A1(n17480), .A2(n9990), .ZN(n9989) );
  INV_X1 U11941 ( .A(n9992), .ZN(n9990) );
  OR2_X1 U11942 ( .A1(n16539), .A2(n17501), .ZN(n16537) );
  NOR2_X1 U11943 ( .A1(n9984), .A2(n17514), .ZN(n9983) );
  AOI21_X1 U11944 ( .B1(n17498), .B2(n16594), .A(n16713), .ZN(n16563) );
  OR2_X1 U11945 ( .A1(n16563), .A2(n16564), .ZN(n9988) );
  AOI211_X1 U11946 ( .C1(n16967), .C2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A(
        n12016), .B(n12015), .ZN(n12017) );
  NAND2_X1 U11947 ( .A1(n17065), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n9938) );
  NOR2_X1 U11948 ( .A1(n11815), .A2(n9940), .ZN(n9939) );
  AND2_X1 U11949 ( .A1(n11812), .A2(n9937), .ZN(n9936) );
  NAND2_X1 U11950 ( .A1(n17092), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n9937) );
  INV_X1 U11951 ( .A(n11829), .ZN(n10017) );
  AOI21_X1 U11952 ( .B1(n17110), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A(
        n11837), .ZN(n11838) );
  NOR2_X1 U11953 ( .A1(n15492), .A2(n17086), .ZN(n11837) );
  INV_X2 U11954 ( .A(n9847), .ZN(n17083) );
  NAND2_X1 U11955 ( .A1(n16277), .A2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12050) );
  AND2_X1 U11956 ( .A1(n16444), .A2(n10004), .ZN(n16277) );
  AND2_X1 U11957 ( .A1(n10005), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n10004) );
  NAND2_X1 U11958 ( .A1(n17444), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n16443) );
  INV_X1 U11959 ( .A(n16443), .ZN(n16444) );
  NOR2_X1 U11960 ( .A1(n17545), .A2(n17546), .ZN(n17528) );
  AND2_X1 U11961 ( .A1(n9998), .A2(n9997), .ZN(n9996) );
  INV_X1 U11962 ( .A(n17581), .ZN(n9997) );
  AOI21_X1 U11963 ( .B1(n11920), .B2(n17628), .A(n11919), .ZN(n15625) );
  NAND2_X1 U11964 ( .A1(n17951), .A2(n15568), .ZN(n17467) );
  NAND2_X1 U11965 ( .A1(n17520), .A2(n10018), .ZN(n11910) );
  NOR2_X1 U11966 ( .A1(n10020), .A2(n10019), .ZN(n10018) );
  NAND2_X1 U11967 ( .A1(n17536), .A2(n17519), .ZN(n17520) );
  AND2_X1 U11968 ( .A1(n11905), .A2(n9941), .ZN(n17568) );
  AOI21_X1 U11969 ( .B1(n17467), .B2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n9942), .ZN(n9941) );
  NOR2_X1 U11970 ( .A1(n17628), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n9942) );
  NAND2_X1 U11971 ( .A1(n17568), .A2(n17893), .ZN(n17567) );
  INV_X1 U11972 ( .A(n17694), .ZN(n17628) );
  NAND2_X1 U11973 ( .A1(n9928), .A2(n9926), .ZN(n17951) );
  NAND2_X1 U11974 ( .A1(n9929), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n9928) );
  NAND2_X1 U11975 ( .A1(n17700), .A2(n9927), .ZN(n9926) );
  INV_X1 U11976 ( .A(n11902), .ZN(n9929) );
  NAND2_X1 U11977 ( .A1(n11903), .A2(n20862), .ZN(n17691) );
  AND2_X1 U11978 ( .A1(n17699), .A2(n11902), .ZN(n11903) );
  NAND2_X1 U11979 ( .A1(n17700), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17699) );
  XNOR2_X1 U11980 ( .A(n11893), .B(n11892), .ZN(n17728) );
  NAND2_X1 U11981 ( .A1(n17728), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n17727) );
  XNOR2_X1 U11982 ( .A(n11886), .B(n11885), .ZN(n17749) );
  NAND2_X1 U11983 ( .A1(n17770), .A2(n11880), .ZN(n17762) );
  XNOR2_X1 U11984 ( .A(n11882), .B(n11881), .ZN(n17763) );
  NAND2_X1 U11985 ( .A1(n17779), .A2(n17771), .ZN(n17770) );
  AOI21_X1 U11986 ( .B1(n11937), .B2(n11936), .A(n11935), .ZN(n18552) );
  INV_X1 U11987 ( .A(n15527), .ZN(n18555) );
  NAND2_X1 U11988 ( .A1(n19891), .A2(n15651), .ZN(n10174) );
  OR2_X1 U11989 ( .A1(n12292), .A2(n11770), .ZN(n14145) );
  NAND2_X1 U11990 ( .A1(n19966), .A2(n13965), .ZN(n15737) );
  NAND2_X1 U11991 ( .A1(n13172), .A2(n13171), .ZN(n15650) );
  INV_X1 U11992 ( .A(n13959), .ZN(n13150) );
  OR2_X1 U11993 ( .A1(n20046), .A2(n13174), .ZN(n14425) );
  OAI22_X1 U11994 ( .A1(n12292), .A2(n11692), .B1(n11712), .B2(n11711), .ZN(
        n11715) );
  XNOR2_X1 U11995 ( .A(n11529), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14310) );
  NAND2_X1 U11996 ( .A1(n11528), .A2(n11527), .ZN(n11529) );
  OR2_X1 U11997 ( .A1(n11767), .A2(n12284), .ZN(n11527) );
  XNOR2_X1 U11998 ( .A(n12286), .B(n10231), .ZN(n14317) );
  OR2_X1 U11999 ( .A1(n11710), .A2(n14149), .ZN(n15649) );
  OR3_X1 U12000 ( .A1(n14470), .A2(n14455), .A3(n14325), .ZN(n14449) );
  AND2_X1 U12001 ( .A1(n11736), .A2(n11735), .ZN(n14505) );
  AND2_X1 U12002 ( .A1(n11746), .A2(n11717), .ZN(n20063) );
  INV_X1 U12003 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20622) );
  NAND2_X1 U12004 ( .A1(n16223), .A2(n13253), .ZN(n19838) );
  OR2_X1 U12005 ( .A1(n19083), .A2(n12637), .ZN(n14841) );
  NOR2_X1 U12006 ( .A1(n15062), .A2(n15290), .ZN(n15045) );
  NAND2_X1 U12007 ( .A1(n16070), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15062) );
  AND2_X1 U12008 ( .A1(n16125), .A2(n13266), .ZN(n16114) );
  OR2_X1 U12009 ( .A1(n18790), .A2(n9779), .ZN(n16055) );
  INV_X1 U12010 ( .A(n15067), .ZN(n16118) );
  NOR2_X1 U12011 ( .A1(n9971), .A2(n21140), .ZN(n9969) );
  NOR2_X1 U12012 ( .A1(n9975), .A2(n9972), .ZN(n9971) );
  INV_X1 U12013 ( .A(n9974), .ZN(n9972) );
  NAND2_X1 U12014 ( .A1(n9976), .A2(n9974), .ZN(n9973) );
  INV_X1 U12015 ( .A(n15360), .ZN(n21130) );
  INV_X1 U12016 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17137) );
  INV_X1 U12017 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n18775) );
  INV_X1 U12018 ( .A(n18089), .ZN(n18084) );
  NOR2_X1 U12019 ( .A1(n18089), .A2(n18093), .ZN(n18085) );
  NAND2_X1 U12020 ( .A1(n19638), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n9921) );
  NOR2_X1 U12021 ( .A1(n11716), .A2(n11582), .ZN(n11247) );
  AOI21_X1 U12022 ( .B1(n11210), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A(n9905), .ZN(n9904) );
  AND2_X1 U12023 ( .A1(n9827), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n9905)
         );
  INV_X1 U12024 ( .A(n10728), .ZN(n10729) );
  NAND2_X1 U12025 ( .A1(n10484), .A2(n10511), .ZN(n10487) );
  INV_X1 U12026 ( .A(n14548), .ZN(n12858) );
  OR2_X1 U12027 ( .A1(n11577), .A2(n11475), .ZN(n11477) );
  INV_X1 U12028 ( .A(n11463), .ZN(n10153) );
  OR2_X1 U12029 ( .A1(n11451), .A2(n11450), .ZN(n11457) );
  INV_X1 U12030 ( .A(n11363), .ZN(n11411) );
  AND3_X1 U12031 ( .A1(n11604), .A2(n11603), .A3(n11726), .ZN(n11611) );
  NAND2_X1 U12032 ( .A1(n11253), .A2(n11252), .ZN(n11254) );
  NAND2_X1 U12033 ( .A1(n9788), .A2(n11253), .ZN(n11584) );
  AOI21_X1 U12034 ( .B1(n10256), .B2(n10255), .A(n10254), .ZN(n10258) );
  NAND2_X1 U12035 ( .A1(n10668), .A2(n10667), .ZN(n10670) );
  AND2_X1 U12036 ( .A1(n10766), .A2(n10765), .ZN(n10768) );
  AOI22_X1 U12037 ( .A1(n9820), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_14__6__SCAN_IN), .B2(n12612), .ZN(n10293) );
  INV_X1 U12038 ( .A(n18135), .ZN(n12020) );
  AOI21_X1 U12039 ( .B1(n18594), .B2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n11925), .ZN(n11934) );
  NOR2_X1 U12040 ( .A1(n12038), .A2(n12039), .ZN(n11925) );
  OAI211_X1 U12041 ( .C1(n13151), .C2(n11280), .A(n13440), .B(n11268), .ZN(
        n11279) );
  NOR2_X1 U12042 ( .A1(n12912), .A2(n14388), .ZN(n12913) );
  AND2_X1 U12043 ( .A1(n12846), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12866) );
  INV_X1 U12044 ( .A(n14088), .ZN(n10156) );
  NOR2_X1 U12045 ( .A1(n12813), .A2(n10158), .ZN(n10157) );
  INV_X1 U12046 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12666) );
  NAND2_X1 U12047 ( .A1(n10236), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n10185) );
  NAND2_X1 U12048 ( .A1(n11524), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n10184) );
  OR2_X1 U12049 ( .A1(n11312), .A2(n11311), .ZN(n11507) );
  NOR2_X1 U12050 ( .A1(n10193), .A2(n9849), .ZN(n10187) );
  NAND2_X1 U12051 ( .A1(n10192), .A2(n10191), .ZN(n10188) );
  OR2_X1 U12052 ( .A1(n11429), .A2(n11428), .ZN(n11453) );
  NAND2_X1 U12053 ( .A1(n9948), .A2(n20252), .ZN(n11439) );
  OR2_X1 U12054 ( .A1(n11323), .A2(n11322), .ZN(n11382) );
  INV_X1 U12055 ( .A(n11252), .ZN(n11263) );
  INV_X1 U12056 ( .A(n11507), .ZN(n11491) );
  OR2_X1 U12057 ( .A1(n11298), .A2(n11297), .ZN(n11371) );
  NOR2_X1 U12058 ( .A1(n20127), .A2(n20098), .ZN(n11361) );
  OR2_X1 U12059 ( .A1(n11408), .A2(n11407), .ZN(n11454) );
  AND2_X1 U12060 ( .A1(n10511), .A2(n13807), .ZN(n10352) );
  NOR2_X1 U12061 ( .A1(n14951), .A2(n10036), .ZN(n10035) );
  INV_X1 U12062 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n10036) );
  NOR2_X1 U12063 ( .A1(n14896), .A2(n14564), .ZN(n14906) );
  INV_X1 U12064 ( .A(n14869), .ZN(n10120) );
  AND2_X1 U12065 ( .A1(n11067), .A2(n10115), .ZN(n11080) );
  INV_X1 U12066 ( .A(n11063), .ZN(n10116) );
  NAND2_X1 U12067 ( .A1(n10127), .A2(n14761), .ZN(n10126) );
  INV_X1 U12068 ( .A(n14567), .ZN(n10127) );
  AND2_X1 U12069 ( .A1(n12396), .A2(n14730), .ZN(n10216) );
  AND2_X1 U12070 ( .A1(n10033), .A2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n10031) );
  NOR2_X1 U12071 ( .A1(n16092), .A2(n10040), .ZN(n10039) );
  INV_X1 U12072 ( .A(n10770), .ZN(n9913) );
  INV_X1 U12073 ( .A(n10800), .ZN(n10148) );
  AND2_X1 U12074 ( .A1(n15247), .A2(n12254), .ZN(n10140) );
  AND2_X1 U12075 ( .A1(n14830), .A2(n15247), .ZN(n15249) );
  NOR2_X1 U12076 ( .A1(n10077), .A2(n13765), .ZN(n10076) );
  INV_X1 U12077 ( .A(n14592), .ZN(n10077) );
  OR2_X1 U12078 ( .A1(n10724), .A2(n10723), .ZN(n10844) );
  NOR2_X1 U12079 ( .A1(n10665), .A2(n10664), .ZN(n11015) );
  OR2_X1 U12080 ( .A1(n10423), .A2(n10422), .ZN(n10835) );
  NOR2_X1 U12081 ( .A1(n10501), .A2(n10500), .ZN(n15369) );
  INV_X1 U12082 ( .A(n10624), .ZN(n10625) );
  AND2_X1 U12083 ( .A1(n9829), .A2(n10614), .ZN(n10615) );
  AND2_X1 U12084 ( .A1(n10314), .A2(n10330), .ZN(n10318) );
  AOI22_X1 U12085 ( .A1(n10386), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12612), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10278) );
  AND2_X1 U12086 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19599), .ZN(
        n12314) );
  NAND3_X1 U12087 ( .A1(n19786), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n19647), 
        .ZN(n13780) );
  NAND3_X1 U12088 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n18739), .ZN(n11783) );
  NOR2_X1 U12089 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10024) );
  NOR2_X1 U12090 ( .A1(n17072), .A2(n15446), .ZN(n9940) );
  NOR2_X1 U12091 ( .A1(n11789), .A2(n11787), .ZN(n11781) );
  INV_X1 U12092 ( .A(n12044), .ZN(n12019) );
  AND2_X1 U12093 ( .A1(n10007), .A2(n10006), .ZN(n10005) );
  NOR2_X1 U12094 ( .A1(n10009), .A2(n10010), .ZN(n10006) );
  INV_X1 U12095 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n10009) );
  NOR2_X1 U12096 ( .A1(n10008), .A2(n17447), .ZN(n10007) );
  INV_X1 U12097 ( .A(n17456), .ZN(n10008) );
  NOR2_X1 U12098 ( .A1(n20862), .A2(n18024), .ZN(n9927) );
  NOR2_X1 U12099 ( .A1(n17704), .A2(n18024), .ZN(n12079) );
  AOI21_X1 U12100 ( .B1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n20878), .A(
        n11931), .ZN(n12040) );
  INV_X1 U12101 ( .A(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n16922) );
  NAND2_X1 U12102 ( .A1(n12952), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12953) );
  AND2_X1 U12103 ( .A1(n11660), .A2(n11659), .ZN(n14123) );
  INV_X1 U12104 ( .A(n19926), .ZN(n19950) );
  OAI21_X1 U12105 ( .B1(n11345), .B2(n11132), .A(n11276), .ZN(n11302) );
  INV_X1 U12106 ( .A(n11251), .ZN(n14222) );
  AND3_X1 U12107 ( .A1(n9772), .A2(n11253), .A3(n20122), .ZN(n11257) );
  AOI21_X1 U12108 ( .B1(n12707), .B2(n12838), .A(n12706), .ZN(n13755) );
  AND2_X1 U12109 ( .A1(n14306), .A2(n13201), .ZN(n13147) );
  INV_X1 U12110 ( .A(n10169), .ZN(n10166) );
  AOI21_X1 U12111 ( .B1(n12977), .B2(n12976), .A(n12975), .ZN(n14035) );
  AND2_X1 U12112 ( .A1(n14362), .A2(n13201), .ZN(n12975) );
  NAND2_X1 U12113 ( .A1(n14260), .A2(n10162), .ZN(n10161) );
  INV_X1 U12114 ( .A(n10164), .ZN(n10162) );
  AND2_X1 U12115 ( .A1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n12913), .ZN(
        n12952) );
  INV_X1 U12116 ( .A(n14046), .ZN(n10163) );
  AND2_X1 U12117 ( .A1(n12866), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12880) );
  CLKBUF_X1 U12118 ( .A(n14057), .Z(n14058) );
  AND2_X1 U12119 ( .A1(n12829), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12846) );
  AND2_X1 U12120 ( .A1(n12824), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n12829) );
  NOR2_X1 U12121 ( .A1(n12808), .A2(n12809), .ZN(n12824) );
  AND2_X1 U12122 ( .A1(n14210), .A2(n14209), .ZN(n14212) );
  NOR2_X1 U12123 ( .A1(n12779), .A2(n13224), .ZN(n12780) );
  CLKBUF_X1 U12124 ( .A(n13197), .Z(n13198) );
  NAND2_X1 U12125 ( .A1(n12752), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12779) );
  INV_X1 U12126 ( .A(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n13224) );
  AND2_X1 U12127 ( .A1(n12737), .A2(n12736), .ZN(n13895) );
  AND3_X1 U12128 ( .A1(n12735), .A2(n12734), .A3(n12733), .ZN(n12736) );
  INV_X1 U12129 ( .A(n12715), .ZN(n12716) );
  NAND2_X1 U12130 ( .A1(n12716), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12738) );
  NAND2_X1 U12131 ( .A1(n12722), .A2(n12721), .ZN(n13870) );
  INV_X1 U12132 ( .A(n12709), .ZN(n12710) );
  NAND2_X1 U12133 ( .A1(n12710), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12715) );
  AND2_X1 U12134 ( .A1(n13731), .A2(n12708), .ZN(n13757) );
  NAND2_X1 U12135 ( .A1(n12703), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12709) );
  INV_X1 U12136 ( .A(n12702), .ZN(n12703) );
  NOR3_X1 U12137 ( .A1(n21068), .A2(n20044), .A3(n12682), .ZN(n12694) );
  INV_X1 U12138 ( .A(n19861), .ZN(n13703) );
  AND2_X1 U12139 ( .A1(n11695), .A2(n11694), .ZN(n14009) );
  AND2_X1 U12140 ( .A1(n10062), .A2(n10061), .ZN(n10060) );
  INV_X1 U12141 ( .A(n14024), .ZN(n10061) );
  NAND2_X1 U12142 ( .A1(n14189), .A2(n10062), .ZN(n14174) );
  NAND2_X1 U12143 ( .A1(n14189), .A2(n10063), .ZN(n14494) );
  NAND2_X1 U12144 ( .A1(n14189), .A2(n14181), .ZN(n14492) );
  AND2_X1 U12145 ( .A1(n11676), .A2(n11675), .ZN(n14048) );
  NAND2_X1 U12146 ( .A1(n11521), .A2(n9946), .ZN(n14510) );
  NAND2_X1 U12147 ( .A1(n14205), .A2(n14123), .ZN(n14122) );
  NAND2_X1 U12148 ( .A1(n14205), .A2(n10054), .ZN(n14101) );
  AND2_X1 U12149 ( .A1(n11657), .A2(n11656), .ZN(n14206) );
  AND2_X1 U12150 ( .A1(n11651), .A2(n11650), .ZN(n13213) );
  NAND2_X1 U12151 ( .A1(n13923), .A2(n11512), .ZN(n10183) );
  AND2_X1 U12152 ( .A1(n11647), .A2(n11646), .ZN(n15883) );
  NAND2_X1 U12153 ( .A1(n15884), .A2(n15883), .ZN(n15886) );
  NAND2_X1 U12154 ( .A1(n12711), .A2(n9856), .ZN(n11486) );
  INV_X1 U12155 ( .A(n9849), .ZN(n10191) );
  AND2_X1 U12156 ( .A1(n11638), .A2(n11637), .ZN(n13825) );
  AND2_X1 U12157 ( .A1(n13739), .A2(n11635), .ZN(n10050) );
  INV_X1 U12158 ( .A(n15918), .ZN(n11635) );
  NAND2_X1 U12159 ( .A1(n13740), .A2(n13739), .ZN(n15919) );
  NAND2_X1 U12160 ( .A1(n13708), .A2(n13710), .ZN(n13709) );
  AND2_X1 U12161 ( .A1(n15872), .A2(n20080), .ZN(n14519) );
  AND2_X1 U12162 ( .A1(n14504), .A2(n20076), .ZN(n14537) );
  XNOR2_X1 U12163 ( .A(n11338), .B(n11337), .ZN(n11336) );
  CLKBUF_X1 U12164 ( .A(n11597), .Z(n11598) );
  INV_X1 U12165 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13447) );
  INV_X1 U12166 ( .A(n11591), .ZN(n11578) );
  INV_X1 U12167 ( .A(n13596), .ZN(n15591) );
  NOR2_X1 U12168 ( .A1(n20763), .A2(n14544), .ZN(n20219) );
  AND2_X1 U12169 ( .A1(n14544), .A2(n20253), .ZN(n20766) );
  NOR2_X1 U12170 ( .A1(n20543), .A2(n20179), .ZN(n20547) );
  AND2_X1 U12171 ( .A1(n20365), .A2(n20763), .ZN(n20759) );
  AND2_X1 U12172 ( .A1(n20543), .A2(n20095), .ZN(n20450) );
  AND3_X1 U12173 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n20098), .A3(n20097), 
        .ZN(n20143) );
  OR2_X1 U12174 ( .A1(n20543), .A2(n20095), .ZN(n20479) );
  CLKBUF_X1 U12175 ( .A(n20458), .Z(n20765) );
  NOR2_X1 U12176 ( .A1(n13466), .A2(n15630), .ZN(n15609) );
  INV_X1 U12177 ( .A(n20697), .ZN(n15630) );
  NOR2_X1 U12178 ( .A1(n10460), .A2(n10265), .ZN(n16212) );
  NAND2_X1 U12179 ( .A1(n12123), .A2(n10035), .ZN(n12094) );
  NAND2_X1 U12180 ( .A1(n14910), .A2(n14894), .ZN(n14896) );
  NOR3_X1 U12181 ( .A1(n14868), .A2(n14869), .A3(P2_EBX_REG_24__SCAN_IN), .ZN(
        n14889) );
  AND2_X1 U12182 ( .A1(n12129), .A2(n9877), .ZN(n12239) );
  NAND2_X1 U12183 ( .A1(n12129), .A2(n10113), .ZN(n12235) );
  NOR2_X1 U12184 ( .A1(n10109), .A2(n10107), .ZN(n10106) );
  INV_X1 U12185 ( .A(n11109), .ZN(n10109) );
  NAND2_X1 U12186 ( .A1(n11119), .A2(n19006), .ZN(n11122) );
  INV_X1 U12187 ( .A(n10107), .ZN(n10105) );
  NAND2_X1 U12188 ( .A1(n11067), .A2(n9852), .ZN(n11077) );
  OAI22_X1 U12189 ( .A1(n10575), .A2(n10545), .B1(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n10540), .ZN(n10549) );
  AND2_X1 U12190 ( .A1(n9851), .A2(n10072), .ZN(n10071) );
  INV_X1 U12191 ( .A(n13682), .ZN(n10072) );
  AND2_X1 U12192 ( .A1(n13488), .A2(n10073), .ZN(n14603) );
  NAND2_X1 U12193 ( .A1(n13488), .A2(n13570), .ZN(n13583) );
  NAND2_X1 U12194 ( .A1(n13478), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n12335) );
  INV_X1 U12195 ( .A(n14694), .ZN(n10219) );
  AND2_X1 U12196 ( .A1(n16022), .A2(n12459), .ZN(n12460) );
  XNOR2_X1 U12197 ( .A(n12484), .B(n12485), .ZN(n14714) );
  BUF_X1 U12198 ( .A(n12458), .Z(n16022) );
  AND2_X1 U12199 ( .A1(n12142), .A2(n12141), .ZN(n15269) );
  CLKBUF_X1 U12200 ( .A(n14733), .Z(n14734) );
  NAND2_X1 U12201 ( .A1(n10211), .A2(n12343), .ZN(n10210) );
  INV_X1 U12202 ( .A(n14746), .ZN(n10211) );
  AND3_X1 U12203 ( .A1(n10888), .A2(n10887), .A3(n10886), .ZN(n15311) );
  NOR2_X1 U12204 ( .A1(n10137), .A2(n13484), .ZN(n10136) );
  NAND2_X1 U12205 ( .A1(n13536), .A2(n13418), .ZN(n10137) );
  AND3_X1 U12206 ( .A1(n10843), .A2(n10842), .A3(n10841), .ZN(n13862) );
  NAND2_X1 U12207 ( .A1(n12123), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12125) );
  INV_X1 U12208 ( .A(n10081), .ZN(n15236) );
  NAND2_X1 U12209 ( .A1(n10042), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n10041) );
  INV_X1 U12210 ( .A(n10043), .ZN(n10042) );
  NOR2_X1 U12211 ( .A1(n12117), .A2(n10043), .ZN(n12119) );
  NOR2_X1 U12212 ( .A1(n12117), .A2(n18834), .ZN(n12118) );
  NAND2_X1 U12213 ( .A1(n12109), .A2(n9834), .ZN(n12110) );
  NAND2_X1 U12214 ( .A1(n12109), .A2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n12108) );
  NOR2_X1 U12215 ( .A1(n10047), .A2(n10049), .ZN(n10045) );
  INV_X1 U12216 ( .A(n12104), .ZN(n10046) );
  OR2_X1 U12217 ( .A1(n12104), .A2(n10048), .ZN(n12105) );
  NOR2_X1 U12218 ( .A1(n12104), .A2(n16124), .ZN(n12106) );
  NAND2_X1 U12219 ( .A1(n12101), .A2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12103) );
  INV_X1 U12220 ( .A(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n14628) );
  NAND2_X1 U12221 ( .A1(n9804), .A2(n10671), .ZN(n13791) );
  NAND2_X1 U12222 ( .A1(n10591), .A2(n10562), .ZN(n10586) );
  INV_X1 U12223 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n12102) );
  NAND2_X1 U12224 ( .A1(n14561), .A2(n14675), .ZN(n10067) );
  NAND2_X1 U12225 ( .A1(n15149), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14939) );
  OR2_X1 U12226 ( .A1(n14959), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n10232) );
  AOI21_X1 U12227 ( .B1(n14901), .B2(n10088), .A(n14955), .ZN(n10087) );
  INV_X1 U12228 ( .A(n14898), .ZN(n10088) );
  INV_X1 U12229 ( .A(n14901), .ZN(n10089) );
  AND2_X1 U12230 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n15112), .ZN(
        n15156) );
  AND2_X1 U12231 ( .A1(n14688), .A2(n10066), .ZN(n14676) );
  NOR2_X1 U12232 ( .A1(n10068), .A2(n10070), .ZN(n10066) );
  INV_X1 U12233 ( .A(n14688), .ZN(n10069) );
  NOR2_X1 U12234 ( .A1(n14980), .A2(n10149), .ZN(n14963) );
  NOR2_X1 U12235 ( .A1(n14897), .A2(n10849), .ZN(n14960) );
  NOR2_X1 U12236 ( .A1(n15966), .A2(n10849), .ZN(n14959) );
  OR2_X1 U12237 ( .A1(n14903), .A2(n15192), .ZN(n14986) );
  OAI21_X1 U12238 ( .B1(n10096), .B2(n10095), .A(n9864), .ZN(n10094) );
  NAND2_X1 U12239 ( .A1(n10081), .A2(n10080), .ZN(n15238) );
  INV_X1 U12240 ( .A(n15235), .ZN(n10080) );
  NAND2_X1 U12241 ( .A1(n15006), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15005) );
  AND2_X1 U12242 ( .A1(n12150), .A2(n12149), .ZN(n15234) );
  NAND2_X1 U12243 ( .A1(n14830), .A2(n10140), .ZN(n15233) );
  NOR2_X1 U12244 ( .A1(n12244), .A2(n12237), .ZN(n9975) );
  INV_X1 U12245 ( .A(n14738), .ZN(n10078) );
  NOR2_X1 U12246 ( .A1(n9959), .A2(n9958), .ZN(n9957) );
  OAI21_X1 U12247 ( .B1(n9960), .B2(n9958), .A(n9956), .ZN(n9955) );
  INV_X1 U12248 ( .A(n14855), .ZN(n9958) );
  NAND2_X1 U12249 ( .A1(n10092), .A2(n9835), .ZN(n15077) );
  NOR3_X1 U12250 ( .A1(n10135), .A2(n13484), .A3(n10134), .ZN(n13535) );
  INV_X1 U12251 ( .A(n13418), .ZN(n10134) );
  INV_X1 U12252 ( .A(n13419), .ZN(n10135) );
  NAND2_X1 U12253 ( .A1(n13419), .A2(n13418), .ZN(n13483) );
  NAND2_X1 U12254 ( .A1(n9915), .A2(n10770), .ZN(n15344) );
  NAND2_X1 U12255 ( .A1(n15344), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n9920) );
  NAND2_X1 U12256 ( .A1(n13849), .A2(n10684), .ZN(n13884) );
  AND3_X1 U12257 ( .A1(n10507), .A2(n15356), .A3(n13242), .ZN(n21126) );
  NAND2_X1 U12258 ( .A1(n13854), .A2(n13853), .ZN(n13852) );
  NAND2_X1 U12259 ( .A1(n13237), .A2(n10504), .ZN(n16138) );
  NOR2_X1 U12260 ( .A1(n19147), .A2(n19146), .ZN(n19358) );
  INV_X1 U12261 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n15372) );
  AND2_X1 U12262 ( .A1(n19836), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n12326) );
  NAND2_X1 U12263 ( .A1(n12306), .A2(n19796), .ZN(n12323) );
  OR2_X1 U12264 ( .A1(n12327), .A2(n12329), .ZN(n12330) );
  AND2_X1 U12265 ( .A1(n14615), .A2(n13479), .ZN(n14612) );
  AND2_X1 U12266 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10271) );
  AND2_X1 U12267 ( .A1(n15383), .A2(n15382), .ZN(n16232) );
  AND2_X1 U12268 ( .A1(n19788), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19357) );
  NOR2_X1 U12269 ( .A1(n10605), .A2(n10618), .ZN(n19355) );
  INV_X1 U12270 ( .A(n10746), .ZN(n19389) );
  INV_X1 U12271 ( .A(n19418), .ZN(n19415) );
  INV_X1 U12272 ( .A(n19192), .ZN(n19414) );
  AND2_X1 U12273 ( .A1(n19147), .A2(n19807), .ZN(n19787) );
  INV_X1 U12274 ( .A(n19787), .ZN(n19482) );
  OR2_X1 U12275 ( .A1(n19788), .A2(n19381), .ZN(n19598) );
  INV_X1 U12276 ( .A(n19638), .ZN(n19645) );
  INV_X1 U12277 ( .A(n19358), .ZN(n19642) );
  NAND2_X1 U12278 ( .A1(n10311), .A2(n10330), .ZN(n10312) );
  INV_X1 U12279 ( .A(n19167), .ZN(n19179) );
  NOR2_X2 U12280 ( .A1(n13781), .A2(n13780), .ZN(n19177) );
  NOR2_X1 U12281 ( .A1(n17308), .A2(n18117), .ZN(n12026) );
  NOR2_X1 U12282 ( .A1(n18580), .A2(n16433), .ZN(n18554) );
  NAND2_X1 U12283 ( .A1(n10003), .A2(n10002), .ZN(n16464) );
  INV_X1 U12284 ( .A(n17431), .ZN(n9982) );
  NAND4_X1 U12285 ( .A1(n18091), .A2(n18777), .A3(n16793), .A4(n18617), .ZN(
        n16677) );
  NAND4_X1 U12286 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(P3_EBX_REG_3__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .A4(n15431), .ZN(n17122) );
  NOR2_X1 U12287 ( .A1(n17149), .A2(n17131), .ZN(n15431) );
  NOR3_X1 U12288 ( .A1(n17291), .A2(n15550), .A3(n15429), .ZN(n15430) );
  INV_X1 U12289 ( .A(n17051), .ZN(n17100) );
  INV_X1 U12290 ( .A(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n16965) );
  INV_X1 U12291 ( .A(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n20943) );
  INV_X1 U12292 ( .A(n18588), .ZN(n15639) );
  NOR2_X1 U12293 ( .A1(n17345), .A2(n17307), .ZN(n17325) );
  NAND2_X1 U12294 ( .A1(n16444), .A2(n10005), .ZN(n16439) );
  NAND2_X1 U12295 ( .A1(n16444), .A2(n17456), .ZN(n17416) );
  AND2_X1 U12296 ( .A1(n17492), .A2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n17444) );
  INV_X1 U12297 ( .A(n17444), .ZN(n17457) );
  NAND2_X1 U12298 ( .A1(n17528), .A2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n17509) );
  NAND2_X1 U12299 ( .A1(n9994), .A2(n9841), .ZN(n17545) );
  NAND2_X1 U12300 ( .A1(n9994), .A2(n9998), .ZN(n17579) );
  NOR2_X1 U12301 ( .A1(n17711), .A2(n17722), .ZN(n17684) );
  NAND2_X1 U12302 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17734) );
  NOR2_X1 U12303 ( .A1(n18560), .A2(n18619), .ZN(n12048) );
  AND2_X1 U12304 ( .A1(n16309), .A2(n16298), .ZN(n15564) );
  NAND2_X1 U12305 ( .A1(n9934), .A2(n9933), .ZN(n9932) );
  NOR2_X1 U12306 ( .A1(n17628), .A2(n17800), .ZN(n9933) );
  INV_X1 U12307 ( .A(n11912), .ZN(n9934) );
  AOI21_X1 U12308 ( .B1(n17576), .B2(n17827), .A(n11907), .ZN(n11908) );
  NOR2_X1 U12309 ( .A1(n17910), .A2(n17932), .ZN(n15568) );
  OR3_X1 U12310 ( .A1(n10022), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n10021) );
  OR2_X1 U12311 ( .A1(n17691), .A2(n10022), .ZN(n17656) );
  NOR2_X1 U12312 ( .A1(n15429), .A2(n18760), .ZN(n12022) );
  NOR2_X1 U12313 ( .A1(n17706), .A2(n17705), .ZN(n17704) );
  INV_X1 U12314 ( .A(n11899), .ZN(n11900) );
  NAND2_X1 U12315 ( .A1(n17749), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n17748) );
  NAND2_X1 U12316 ( .A1(n17763), .A2(n17762), .ZN(n17761) );
  NOR2_X1 U12317 ( .A1(n15556), .A2(n15533), .ZN(n15566) );
  INV_X1 U12318 ( .A(n18567), .ZN(n18582) );
  NOR2_X1 U12319 ( .A1(n18779), .A2(n15427), .ZN(n18567) );
  NAND2_X1 U12320 ( .A1(n18562), .A2(n18564), .ZN(n16432) );
  INV_X1 U12321 ( .A(n13781), .ZN(n14769) );
  NAND2_X1 U12322 ( .A1(n13528), .A2(n13260), .ZN(n20785) );
  INV_X1 U12323 ( .A(n19942), .ZN(n19909) );
  AND2_X1 U12324 ( .A1(n13747), .A2(n13221), .ZN(n19937) );
  AND2_X1 U12325 ( .A1(n15726), .A2(n13745), .ZN(n19931) );
  INV_X1 U12326 ( .A(n15737), .ZN(n19962) );
  NOR2_X2 U12327 ( .A1(n20025), .A2(n9787), .ZN(n20015) );
  XNOR2_X1 U12328 ( .A(n13207), .B(n13206), .ZN(n13973) );
  OR2_X1 U12329 ( .A1(n13103), .A2(n13069), .ZN(n15667) );
  AND2_X1 U12330 ( .A1(n13067), .A2(n13046), .ZN(n14341) );
  OAI21_X1 U12331 ( .B1(n14368), .B2(n10186), .A(n14352), .ZN(n14359) );
  INV_X1 U12332 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n14373) );
  INV_X1 U12333 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n14388) );
  INV_X1 U12334 ( .A(n20094), .ZN(n20038) );
  INV_X1 U12335 ( .A(n14425), .ZN(n20043) );
  AND2_X1 U12336 ( .A1(n14425), .A2(n13175), .ZN(n20045) );
  AND2_X1 U12337 ( .A1(n15598), .A2(n13703), .ZN(n20046) );
  INV_X1 U12338 ( .A(n20046), .ZN(n19867) );
  OR2_X1 U12339 ( .A1(n15931), .A2(n20544), .ZN(n20094) );
  NAND2_X1 U12340 ( .A1(n12302), .A2(n10058), .ZN(n10057) );
  INV_X1 U12341 ( .A(n13971), .ZN(n10058) );
  XNOR2_X1 U12342 ( .A(n10059), .B(n12296), .ZN(n14142) );
  NAND2_X1 U12343 ( .A1(n12294), .A2(n12293), .ZN(n10059) );
  XNOR2_X1 U12344 ( .A(n13167), .B(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14446) );
  NAND2_X1 U12345 ( .A1(n10235), .A2(n13165), .ZN(n13167) );
  NOR2_X1 U12346 ( .A1(n14320), .A2(n10234), .ZN(n13165) );
  NAND2_X1 U12347 ( .A1(n11524), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n14525) );
  AND2_X1 U12348 ( .A1(n14505), .A2(n11738), .ZN(n15841) );
  NAND2_X1 U12349 ( .A1(n15792), .A2(n15794), .ZN(n15793) );
  INV_X1 U12350 ( .A(n15923), .ZN(n20086) );
  INV_X1 U12351 ( .A(n14519), .ZN(n15897) );
  CLKBUF_X1 U12352 ( .A(n13437), .Z(n13438) );
  INV_X1 U12353 ( .A(n20458), .ZN(n20632) );
  INV_X1 U12354 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n20869) );
  OR2_X1 U12355 ( .A1(n13608), .A2(n13607), .ZN(n20771) );
  INV_X1 U12356 ( .A(n13606), .ZN(n15613) );
  NOR2_X1 U12357 ( .A1(n20493), .A2(n13466), .ZN(n13606) );
  NOR2_X1 U12358 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n14552) );
  OAI211_X1 U12359 ( .C1(n20105), .C2(n20493), .A(n20429), .B(n20104), .ZN(
        n20148) );
  INV_X1 U12360 ( .A(n20371), .ZN(n20391) );
  AND2_X1 U12361 ( .A1(n20759), .A2(n20547), .ZN(n20445) );
  OAI21_X1 U12362 ( .B1(n20546), .B2(n20545), .A(n20630), .ZN(n20565) );
  OAI211_X1 U12363 ( .C1(n20611), .C2(n20581), .A(n20580), .B(n20579), .ZN(
        n20614) );
  INV_X1 U12364 ( .A(n20486), .ZN(n20626) );
  INV_X1 U12365 ( .A(n20499), .ZN(n20640) );
  INV_X1 U12366 ( .A(n20504), .ZN(n20646) );
  INV_X1 U12367 ( .A(n20509), .ZN(n20652) );
  INV_X1 U12368 ( .A(n20514), .ZN(n20658) );
  INV_X1 U12369 ( .A(n20519), .ZN(n20664) );
  INV_X1 U12370 ( .A(n20524), .ZN(n20670) );
  INV_X1 U12371 ( .A(n20634), .ZN(n20680) );
  NAND2_X1 U12372 ( .A1(n20687), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n19861) );
  INV_X1 U12373 ( .A(n15939), .ZN(n15933) );
  INV_X1 U12374 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n15937) );
  AND2_X1 U12375 ( .A1(n15937), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20687) );
  NOR2_X1 U12376 ( .A1(n19836), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n18785) );
  OR2_X1 U12377 ( .A1(n15137), .A2(n18981), .ZN(n12220) );
  NOR2_X1 U12378 ( .A1(n14910), .A2(n14880), .ZN(n15975) );
  NAND2_X1 U12379 ( .A1(n12116), .A2(n10243), .ZN(n18865) );
  OR2_X1 U12380 ( .A1(n19838), .A2(n12173), .ZN(n18960) );
  CLKBUF_X1 U12381 ( .A(n19002), .Z(n18964) );
  INV_X1 U12382 ( .A(n18960), .ZN(n18990) );
  OR2_X1 U12383 ( .A1(n19838), .A2(n12169), .ZN(n18982) );
  INV_X1 U12384 ( .A(n18981), .ZN(n18997) );
  INV_X1 U12385 ( .A(n13761), .ZN(n10209) );
  OR2_X1 U12386 ( .A1(n10923), .A2(n10922), .ZN(n13762) );
  NAND2_X1 U12387 ( .A1(n10213), .A2(n12342), .ZN(n10212) );
  INV_X1 U12388 ( .A(n10214), .ZN(n10213) );
  NOR2_X1 U12389 ( .A1(n10130), .A2(n10129), .ZN(n10128) );
  INV_X1 U12390 ( .A(n14760), .ZN(n10130) );
  INV_X1 U12391 ( .A(n19084), .ZN(n16040) );
  NAND2_X1 U12392 ( .A1(n13724), .A2(n10133), .ZN(n13913) );
  NOR2_X1 U12393 ( .A1(n19086), .A2(n19084), .ZN(n19061) );
  AND2_X1 U12394 ( .A1(n19044), .A2(n12636), .ZN(n19084) );
  NAND2_X1 U12395 ( .A1(n12635), .A2(n19840), .ZN(n19083) );
  INV_X1 U12396 ( .A(n19079), .ZN(n19086) );
  AND2_X1 U12397 ( .A1(n14841), .A2(n13406), .ZN(n19091) );
  NAND2_X1 U12398 ( .A1(n13375), .A2(n13374), .ZN(n19121) );
  AND2_X1 U12399 ( .A1(n13270), .A2(n9779), .ZN(n19139) );
  INV_X1 U12400 ( .A(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n16092) );
  AND2_X1 U12401 ( .A1(n10090), .A2(n9874), .ZN(n15314) );
  INV_X1 U12402 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n16113) );
  NAND2_X1 U12403 ( .A1(n15333), .A2(n10800), .ZN(n16109) );
  INV_X1 U12404 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n10565) );
  NAND2_X1 U12405 ( .A1(n18790), .A2(n12271), .ZN(n16125) );
  INV_X1 U12406 ( .A(n16088), .ZN(n16117) );
  INV_X1 U12407 ( .A(n16114), .ZN(n16068) );
  INV_X1 U12408 ( .A(n12319), .ZN(n15359) );
  INV_X1 U12409 ( .A(n16125), .ZN(n16062) );
  OAI21_X1 U12410 ( .B1(n14932), .B2(n14935), .A(n10238), .ZN(n14917) );
  NAND2_X1 U12411 ( .A1(n10093), .A2(n10096), .ZN(n15007) );
  NAND2_X1 U12412 ( .A1(n10101), .A2(n10098), .ZN(n10093) );
  NAND2_X1 U12413 ( .A1(n9954), .A2(n9960), .ZN(n12222) );
  NAND2_X1 U12414 ( .A1(n15060), .A2(n9961), .ZN(n9954) );
  NOR2_X1 U12415 ( .A1(n15301), .A2(n9917), .ZN(n9916) );
  OR2_X1 U12416 ( .A1(n15045), .A2(n9896), .ZN(n9918) );
  AND2_X1 U12417 ( .A1(n13241), .A2(n11115), .ZN(n9917) );
  NAND2_X1 U12418 ( .A1(n9966), .A2(n9964), .ZN(n15046) );
  NAND2_X1 U12419 ( .A1(n15060), .A2(n15057), .ZN(n9966) );
  AND2_X1 U12420 ( .A1(n10101), .A2(n10103), .ZN(n15071) );
  NAND2_X1 U12421 ( .A1(n10090), .A2(n11074), .ZN(n15093) );
  NAND2_X1 U12422 ( .A1(n15105), .A2(n15104), .ZN(n15333) );
  NAND2_X1 U12423 ( .A1(n11125), .A2(n11007), .ZN(n15360) );
  AND2_X1 U12424 ( .A1(n11125), .A2(n10956), .ZN(n16181) );
  INV_X1 U12425 ( .A(n16157), .ZN(n21137) );
  INV_X1 U12426 ( .A(n16138), .ZN(n15357) );
  OR2_X1 U12427 ( .A1(n12327), .A2(n13346), .ZN(n19817) );
  INV_X1 U12428 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19813) );
  NAND2_X1 U12429 ( .A1(n13501), .A2(n13500), .ZN(n19807) );
  OR2_X1 U12430 ( .A1(n13499), .A2(n13498), .ZN(n13500) );
  INV_X1 U12431 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19804) );
  INV_X1 U12432 ( .A(n19147), .ZN(n19802) );
  INV_X1 U12433 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n21060) );
  INV_X1 U12434 ( .A(n19807), .ZN(n19146) );
  NAND2_X1 U12435 ( .A1(n13494), .A2(n13497), .ZN(n19147) );
  OR2_X1 U12436 ( .A1(n13495), .A2(n13496), .ZN(n13497) );
  AND3_X1 U12437 ( .A1(n10367), .A2(n10476), .A3(n10491), .ZN(n10368) );
  OAI21_X1 U12438 ( .B1(n19272), .B2(n19287), .A(n19271), .ZN(n19290) );
  OR2_X1 U12439 ( .A1(n19314), .A2(n19536), .ZN(n19313) );
  INV_X1 U12440 ( .A(n19468), .ZN(n19449) );
  NOR2_X1 U12441 ( .A1(n19537), .A2(n19414), .ZN(n19468) );
  INV_X1 U12442 ( .A(n19652), .ZN(n19551) );
  INV_X1 U12443 ( .A(n19689), .ZN(n19585) );
  INV_X1 U12444 ( .A(n19675), .ZN(n19620) );
  OAI21_X1 U12445 ( .B1(n19608), .B2(n19607), .A(n19606), .ZN(n19632) );
  AND2_X1 U12446 ( .A1(n16218), .A2(n19179), .ZN(n19640) );
  INV_X1 U12447 ( .A(n19614), .ZN(n19655) );
  AND2_X1 U12448 ( .A1(n9779), .A2(n19179), .ZN(n19653) );
  INV_X1 U12449 ( .A(n19489), .ZN(n19660) );
  AND2_X1 U12450 ( .A1(n13807), .A2(n19179), .ZN(n19664) );
  INV_X1 U12451 ( .A(n19627), .ZN(n19678) );
  AND2_X1 U12452 ( .A1(n10808), .A2(n19179), .ZN(n19676) );
  INV_X1 U12453 ( .A(n19699), .ZN(n19685) );
  OR2_X1 U12454 ( .A1(n19537), .A2(n19642), .ZN(n19699) );
  INV_X1 U12455 ( .A(n19688), .ZN(n19695) );
  INV_X1 U12456 ( .A(n19637), .ZN(n19694) );
  AND2_X1 U12457 ( .A1(n10480), .A2(n19179), .ZN(n19690) );
  AND2_X1 U12458 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n18785), .ZN(n19840) );
  NAND2_X1 U12459 ( .A1(n18783), .A2(n17308), .ZN(n18780) );
  INV_X1 U12460 ( .A(n18783), .ZN(n18777) );
  NAND2_X1 U12461 ( .A1(n18611), .A2(n18555), .ZN(n17345) );
  AND2_X1 U12462 ( .A1(n16461), .A2(n16818), .ZN(n10000) );
  OAI21_X1 U12463 ( .B1(n10003), .B2(n16713), .A(n9999), .ZN(n10001) );
  AOI21_X1 U12464 ( .B1(n9993), .B2(n16467), .A(n9844), .ZN(n9999) );
  OAI21_X1 U12465 ( .B1(n16499), .B2(n9979), .A(n9978), .ZN(n16488) );
  NAND2_X1 U12466 ( .A1(n9982), .A2(n9980), .ZN(n9979) );
  NAND2_X1 U12467 ( .A1(n16713), .A2(n9982), .ZN(n9978) );
  INV_X1 U12468 ( .A(n17449), .ZN(n9980) );
  INV_X1 U12469 ( .A(n9981), .ZN(n16498) );
  NAND2_X1 U12470 ( .A1(n9991), .A2(n9992), .ZN(n16522) );
  AND2_X1 U12471 ( .A1(n16537), .A2(n9993), .ZN(n16527) );
  AND2_X1 U12472 ( .A1(n9988), .A2(n16790), .ZN(n16552) );
  NOR2_X1 U12473 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16575), .ZN(n16560) );
  NOR2_X1 U12474 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n16647), .ZN(n16637) );
  NOR2_X2 U12475 ( .A1(n18780), .A2(n18612), .ZN(n16772) );
  INV_X1 U12476 ( .A(n16772), .ZN(n16794) );
  INV_X1 U12477 ( .A(n16767), .ZN(n16801) );
  INV_X1 U12478 ( .A(n16677), .ZN(n16804) );
  AND2_X1 U12479 ( .A1(P3_EBX_REG_25__SCAN_IN), .A2(n16868), .ZN(n16863) );
  NOR3_X1 U12480 ( .A1(n16813), .A2(n16812), .A3(n16887), .ZN(n16874) );
  INV_X1 U12481 ( .A(n16869), .ZN(n16887) );
  NOR2_X1 U12482 ( .A1(n17291), .A2(n16929), .ZN(n16915) );
  NOR2_X1 U12483 ( .A1(n16945), .A2(n16932), .ZN(n16930) );
  NAND2_X1 U12484 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n16930), .ZN(n16929) );
  NAND2_X1 U12485 ( .A1(n17001), .A2(n16946), .ZN(n16932) );
  AND4_X1 U12486 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(P3_EBX_REG_6__SCAN_IN), 
        .A3(P3_EBX_REG_5__SCAN_IN), .A4(n17127), .ZN(n17118) );
  INV_X1 U12487 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17126) );
  INV_X1 U12488 ( .A(n17122), .ZN(n17127) );
  NAND2_X1 U12489 ( .A1(P3_EAX_REG_27__SCAN_IN), .A2(n17178), .ZN(n17173) );
  NOR2_X1 U12490 ( .A1(n17355), .A2(n17220), .ZN(n17215) );
  NOR2_X1 U12491 ( .A1(n17413), .A2(n17239), .ZN(n17233) );
  NAND2_X1 U12492 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n17233), .ZN(n17232) );
  INV_X1 U12493 ( .A(n17214), .ZN(n17231) );
  NOR2_X1 U12494 ( .A1(n18145), .A2(n17155), .ZN(n17270) );
  NOR3_X1 U12495 ( .A1(n17291), .A2(n17302), .A3(n17237), .ZN(n17276) );
  NOR2_X1 U12496 ( .A1(n11817), .A2(n9935), .ZN(n17288) );
  NOR2_X1 U12497 ( .A1(n10017), .A2(n10016), .ZN(n10015) );
  NOR2_X1 U12498 ( .A1(n16970), .A2(n16934), .ZN(n10016) );
  INV_X1 U12499 ( .A(n17300), .ZN(n17295) );
  AND2_X1 U12500 ( .A1(n17083), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n11843) );
  INV_X1 U12501 ( .A(n17270), .ZN(n17303) );
  NOR2_X1 U12502 ( .A1(n17155), .A2(n15638), .ZN(n17301) );
  NOR2_X1 U12504 ( .A1(n17509), .A2(n17510), .ZN(n17492) );
  NOR2_X1 U12505 ( .A1(n17646), .A2(n9995), .ZN(n17566) );
  INV_X1 U12506 ( .A(n9996), .ZN(n9995) );
  NAND2_X1 U12507 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n17672), .ZN(n17591) );
  INV_X1 U12508 ( .A(n17467), .ZN(n17919) );
  NOR2_X1 U12509 ( .A1(n17768), .A2(n17735), .ZN(n17672) );
  NOR2_X1 U12510 ( .A1(n17702), .A2(n17687), .ZN(n17685) );
  INV_X1 U12511 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17687) );
  NOR2_X2 U12512 ( .A1(n17274), .A2(n17784), .ZN(n17695) );
  INV_X1 U12513 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n17702) );
  NAND2_X1 U12514 ( .A1(n17726), .A2(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n17711) );
  OR2_X1 U12515 ( .A1(n18401), .A2(n18456), .ZN(n18428) );
  INV_X1 U12516 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n17722) );
  NOR2_X1 U12517 ( .A1(n20959), .A2(n17734), .ZN(n17726) );
  OAI21_X2 U12518 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n18766), .A(n16417), 
        .ZN(n17780) );
  INV_X1 U12519 ( .A(n11917), .ZN(n11924) );
  OAI21_X1 U12520 ( .B1(n11921), .B2(n11916), .A(n11915), .ZN(n11917) );
  NAND2_X1 U12521 ( .A1(n9931), .A2(n9930), .ZN(n17433) );
  NOR2_X1 U12522 ( .A1(n11912), .A2(n17800), .ZN(n9930) );
  INV_X1 U12523 ( .A(n17442), .ZN(n9931) );
  NAND2_X1 U12524 ( .A1(n17520), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n17483) );
  NOR2_X1 U12525 ( .A1(n17691), .A2(n17694), .ZN(n17668) );
  NAND2_X1 U12526 ( .A1(n17727), .A2(n11895), .ZN(n17713) );
  NOR2_X1 U12527 ( .A1(n18072), .A2(n18084), .ZN(n18082) );
  AOI221_X1 U12528 ( .B1(n15551), .B2(n18552), .C1(n15550), .C2(n18552), .A(
        n15549), .ZN(n15560) );
  INV_X1 U12529 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18599) );
  INV_X1 U12530 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n20878) );
  INV_X1 U12531 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n18722) );
  AOI211_X1 U12532 ( .C1(n18611), .C2(n18586), .A(n18113), .B(n15539), .ZN(
        n18746) );
  INV_X1 U12533 ( .A(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n20935) );
  INV_X1 U12534 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n18716) );
  AND2_X1 U12535 ( .A1(n13192), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n20092)
         );
  OAI21_X1 U12537 ( .B1(n15650), .B2(n15726), .A(n10172), .ZN(P1_U2812) );
  AOI21_X1 U12538 ( .B1(n10175), .B2(n19948), .A(n10173), .ZN(n10172) );
  INV_X1 U12539 ( .A(n15649), .ZN(n10175) );
  NAND2_X1 U12540 ( .A1(n13160), .A2(n13159), .ZN(P1_U2842) );
  NAND2_X1 U12541 ( .A1(n14307), .A2(n13156), .ZN(n13160) );
  NAND2_X1 U12542 ( .A1(n11762), .A2(n11761), .ZN(n11763) );
  AND2_X1 U12543 ( .A1(n11777), .A2(n11776), .ZN(n11778) );
  OAI21_X1 U12544 ( .B1(n12280), .B2(n16055), .A(n12279), .ZN(n12281) );
  NAND2_X1 U12545 ( .A1(n9973), .A2(n11126), .ZN(n9970) );
  OR4_X1 U12546 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n18623), .A3(n18764), 
        .A4(n18622), .ZN(n18625) );
  NAND2_X1 U12547 ( .A1(n19030), .A2(n13680), .ZN(n13679) );
  INV_X1 U12548 ( .A(n12116), .ZN(n14665) );
  INV_X1 U12549 ( .A(n11820), .ZN(n15498) );
  NOR2_X1 U12550 ( .A1(n16789), .A2(n11788), .ZN(n11832) );
  OR2_X1 U12551 ( .A1(n10873), .A2(n10872), .ZN(n13680) );
  NAND2_X1 U12553 ( .A1(n13894), .A2(n13919), .ZN(n13196) );
  AND2_X1 U12554 ( .A1(n10155), .A2(n9873), .ZN(n14070) );
  NAND2_X1 U12555 ( .A1(n10155), .A2(n10160), .ZN(n9832) );
  AND2_X1 U12556 ( .A1(n14735), .A2(n12396), .ZN(n14729) );
  AND2_X1 U12557 ( .A1(n10039), .A2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n9834) );
  AND2_X1 U12558 ( .A1(n9874), .A2(n15316), .ZN(n9835) );
  AOI21_X1 U12559 ( .B1(n10101), .B2(n10100), .A(n14861), .ZN(n15228) );
  NAND2_X1 U12560 ( .A1(n10163), .A2(n12920), .ZN(n14177) );
  XNOR2_X1 U12561 ( .A(n12512), .B(n12513), .ZN(n14705) );
  XNOR2_X1 U12562 ( .A(n12537), .B(n9900), .ZN(n14697) );
  AND2_X1 U12563 ( .A1(n11058), .A2(n9881), .ZN(n9837) );
  INV_X1 U12564 ( .A(n10482), .ZN(n11013) );
  AND2_X1 U12565 ( .A1(n14616), .A2(n9892), .ZN(n9838) );
  INV_X1 U12566 ( .A(n10383), .ZN(n12424) );
  INV_X1 U12567 ( .A(n16082), .ZN(n10103) );
  AND2_X1 U12568 ( .A1(n12721), .A2(n9906), .ZN(n9839) );
  AND2_X1 U12569 ( .A1(n9966), .A2(n15058), .ZN(n9840) );
  NAND2_X1 U12570 ( .A1(n10209), .A2(n12343), .ZN(n14745) );
  AND2_X1 U12571 ( .A1(n9996), .A2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n9841) );
  AND2_X1 U12572 ( .A1(n10076), .A2(n10075), .ZN(n9842) );
  AND2_X1 U12573 ( .A1(n9981), .A2(n9993), .ZN(n9843) );
  OR3_X1 U12574 ( .A1(n16713), .A2(n16456), .A3(n16793), .ZN(n9844) );
  OR2_X1 U12575 ( .A1(n12251), .A2(n15241), .ZN(n9845) );
  OR2_X1 U12577 ( .A1(n12117), .A2(n10041), .ZN(n9846) );
  OR2_X1 U12578 ( .A1(n11782), .A2(n11787), .ZN(n9847) );
  OR2_X2 U12579 ( .A1(n16789), .A2(n11789), .ZN(n9848) );
  NAND2_X1 U12580 ( .A1(n11059), .A2(n11058), .ZN(n15101) );
  NAND2_X1 U12581 ( .A1(n10155), .A2(n10157), .ZN(n14086) );
  NAND2_X1 U12582 ( .A1(n14026), .A2(n14009), .ZN(n14008) );
  AND2_X1 U12583 ( .A1(n11461), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n9849) );
  NOR2_X1 U12584 ( .A1(n14046), .A2(n10164), .ZN(n14179) );
  AND4_X1 U12585 ( .A1(n11163), .A2(n11162), .A3(n11161), .A4(n11160), .ZN(
        n9850) );
  AND2_X1 U12586 ( .A1(n14057), .A2(n14059), .ZN(n14045) );
  NAND2_X1 U12587 ( .A1(n15095), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15083) );
  NAND2_X1 U12588 ( .A1(n14004), .A2(n10167), .ZN(n13171) );
  NAND2_X1 U12589 ( .A1(n11251), .A2(n9772), .ZN(n11262) );
  AND2_X1 U12590 ( .A1(n10073), .A2(n14604), .ZN(n9851) );
  AND2_X1 U12591 ( .A1(n11065), .A2(n10116), .ZN(n9852) );
  NAND2_X1 U12592 ( .A1(n10183), .A2(n11514), .ZN(n13936) );
  NOR2_X1 U12593 ( .A1(n14711), .A2(n14701), .ZN(n14688) );
  OR2_X1 U12594 ( .A1(n13478), .A2(n13477), .ZN(n13479) );
  OR2_X1 U12595 ( .A1(n9784), .A2(n12251), .ZN(n14918) );
  AND2_X1 U12596 ( .A1(n10098), .A2(n15008), .ZN(n9853) );
  NOR2_X1 U12597 ( .A1(n14692), .A2(n14694), .ZN(n14693) );
  OR2_X1 U12598 ( .A1(n14008), .A2(n14157), .ZN(n9854) );
  AND3_X1 U12599 ( .A1(n11229), .A2(n11235), .A3(n9904), .ZN(n9855) );
  NOR2_X1 U12600 ( .A1(n14817), .A2(n14808), .ZN(n14796) );
  AND2_X1 U12601 ( .A1(n11494), .A2(n11541), .ZN(n9856) );
  NOR2_X1 U12602 ( .A1(n16452), .A2(n10000), .ZN(n9857) );
  OR2_X1 U12603 ( .A1(n12167), .A2(n10543), .ZN(n9858) );
  AND2_X1 U12604 ( .A1(n10800), .A2(n9914), .ZN(n9859) );
  AND2_X1 U12605 ( .A1(n10115), .A2(n18930), .ZN(n9860) );
  INV_X1 U12606 ( .A(n10121), .ZN(n14872) );
  NOR2_X1 U12607 ( .A1(n14868), .A2(n14869), .ZN(n10121) );
  OR2_X1 U12608 ( .A1(n13197), .A2(n14215), .ZN(n9861) );
  AND2_X1 U12609 ( .A1(n10270), .A2(n10330), .ZN(n9862) );
  AND2_X1 U12610 ( .A1(n10275), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9863) );
  INV_X1 U12611 ( .A(n10110), .ZN(n11098) );
  NAND2_X1 U12612 ( .A1(n11089), .A2(n11091), .ZN(n10110) );
  OR2_X1 U12613 ( .A1(n14871), .A2(n10230), .ZN(n9864) );
  INV_X1 U12614 ( .A(n13807), .ZN(n10367) );
  INV_X1 U12615 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n16124) );
  AND3_X1 U12616 ( .A1(n11813), .A2(n9939), .A3(n9938), .ZN(n9865) );
  OR2_X1 U12617 ( .A1(n10496), .A2(n12305), .ZN(n9866) );
  AND2_X1 U12618 ( .A1(n10001), .A2(n9857), .ZN(n9867) );
  AND2_X1 U12619 ( .A1(n10371), .A2(n10482), .ZN(n10485) );
  OR2_X1 U12620 ( .A1(n19473), .A2(n12527), .ZN(n9868) );
  OR2_X1 U12621 ( .A1(n14352), .A2(n13937), .ZN(n9869) );
  INV_X1 U12622 ( .A(n10820), .ZN(n12166) );
  NAND2_X1 U12623 ( .A1(n10806), .A2(n9776), .ZN(n10951) );
  NOR2_X1 U12624 ( .A1(n13678), .A2(n10214), .ZN(n13716) );
  AND2_X1 U12625 ( .A1(n13724), .A2(n10131), .ZN(n9870) );
  AND2_X1 U12626 ( .A1(n14830), .A2(n10138), .ZN(n14816) );
  AND2_X1 U12627 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n12101) );
  NAND2_X1 U12628 ( .A1(n14723), .A2(n14715), .ZN(n14708) );
  INV_X1 U12629 ( .A(n14848), .ZN(n9956) );
  NOR2_X1 U12630 ( .A1(n12104), .A2(n10047), .ZN(n9871) );
  NOR3_X1 U12631 ( .A1(n15051), .A2(n11005), .A3(n15272), .ZN(n14737) );
  AND2_X1 U12632 ( .A1(n15091), .A2(n15315), .ZN(n9872) );
  AND2_X1 U12633 ( .A1(n10157), .A2(n10156), .ZN(n9873) );
  AND2_X1 U12634 ( .A1(n10091), .A2(n11074), .ZN(n9874) );
  OR3_X1 U12635 ( .A1(n10078), .A2(n11005), .A3(n15272), .ZN(n9875) );
  NOR2_X1 U12636 ( .A1(n13732), .A2(n13733), .ZN(n13731) );
  AND2_X1 U12637 ( .A1(n13724), .A2(n14577), .ZN(n9876) );
  XNOR2_X1 U12638 ( .A(n12331), .B(n12332), .ZN(n13495) );
  NOR2_X1 U12639 ( .A1(n13761), .A2(n10210), .ZN(n13910) );
  AND2_X1 U12640 ( .A1(n10113), .A2(n10112), .ZN(n9877) );
  NAND2_X1 U12641 ( .A1(n14735), .A2(n10216), .ZN(n9878) );
  NAND2_X1 U12642 ( .A1(n14705), .A2(n14707), .ZN(n14706) );
  NAND2_X1 U12643 ( .A1(n20033), .A2(n11438), .ZN(n15792) );
  AND2_X1 U12644 ( .A1(n11524), .A2(n11520), .ZN(n9879) );
  NOR2_X1 U12645 ( .A1(n17291), .A2(n17193), .ZN(n17188) );
  AND2_X1 U12646 ( .A1(n12109), .A2(n10039), .ZN(n9880) );
  NAND2_X1 U12647 ( .A1(n10497), .A2(n10496), .ZN(n10492) );
  AND2_X1 U12648 ( .A1(n11069), .A2(n11068), .ZN(n9881) );
  NOR2_X1 U12649 ( .A1(n14081), .A2(n14062), .ZN(n11673) );
  INV_X1 U12650 ( .A(n10079), .ZN(n15273) );
  NOR2_X1 U12651 ( .A1(n15051), .A2(n11005), .ZN(n10079) );
  INV_X1 U12652 ( .A(n12341), .ZN(n19024) );
  OR2_X1 U12653 ( .A1(n10885), .A2(n10884), .ZN(n12341) );
  INV_X1 U12654 ( .A(n11477), .ZN(n11476) );
  INV_X1 U12655 ( .A(n14861), .ZN(n10102) );
  INV_X1 U12656 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n18834) );
  AND2_X1 U12657 ( .A1(n16464), .A2(n16790), .ZN(n9882) );
  AND2_X1 U12658 ( .A1(n10131), .A2(n12140), .ZN(n9883) );
  AND2_X1 U12659 ( .A1(n11518), .A2(n14422), .ZN(n9884) );
  OR2_X1 U12660 ( .A1(n15730), .A2(n15653), .ZN(n9885) );
  AND2_X1 U12661 ( .A1(n10054), .A2(n10053), .ZN(n9886) );
  AND2_X1 U12662 ( .A1(n17622), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n9887) );
  AND2_X1 U12663 ( .A1(n9873), .A2(n12865), .ZN(n9888) );
  INV_X2 U12664 ( .A(n19020), .ZN(n19037) );
  OR2_X2 U12665 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n13256), .ZN(n9889) );
  INV_X1 U12666 ( .A(n16963), .ZN(n17150) );
  INV_X1 U12667 ( .A(n17150), .ZN(n17141) );
  NOR2_X1 U12668 ( .A1(n20760), .A2(n20102), .ZN(n9890) );
  NAND2_X1 U12669 ( .A1(n9806), .A2(n14616), .ZN(n13486) );
  INV_X1 U12670 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10267) );
  NOR2_X1 U12671 ( .A1(n13852), .A2(n13487), .ZN(n13488) );
  NAND2_X1 U12672 ( .A1(n13488), .A2(n9851), .ZN(n13681) );
  NAND2_X1 U12673 ( .A1(n13717), .A2(n10076), .ZN(n13763) );
  NAND2_X1 U12674 ( .A1(n13717), .A2(n14592), .ZN(n13764) );
  AND2_X1 U12675 ( .A1(n16444), .A2(n10007), .ZN(n9891) );
  AND2_X1 U12676 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n9892) );
  NOR2_X1 U12677 ( .A1(n15307), .A2(n13718), .ZN(n13717) );
  AND2_X1 U12678 ( .A1(n12097), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12096) );
  INV_X1 U12679 ( .A(n12128), .ZN(n10114) );
  NAND4_X2 U12680 ( .A1(n10797), .A2(n10796), .A3(n10795), .A4(n10794), .ZN(
        n11060) );
  NOR2_X1 U12681 ( .A1(n12121), .A2(n14990), .ZN(n12097) );
  OR2_X1 U12682 ( .A1(n11079), .A2(n14912), .ZN(n14886) );
  INV_X1 U12683 ( .A(n14886), .ZN(n10104) );
  NAND2_X1 U12684 ( .A1(n17684), .A2(n12049), .ZN(n17646) );
  INV_X1 U12685 ( .A(n17646), .ZN(n9994) );
  AND2_X1 U12686 ( .A1(n14912), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n9893) );
  OR2_X1 U12687 ( .A1(n12117), .A2(n10044), .ZN(n9894) );
  OR2_X1 U12688 ( .A1(n10067), .A2(n10068), .ZN(n9895) );
  INV_X1 U12689 ( .A(n14561), .ZN(n10070) );
  INV_X1 U12690 ( .A(n10034), .ZN(n10033) );
  NAND2_X1 U12691 ( .A1(n10035), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10034) );
  AND2_X1 U12692 ( .A1(n13237), .A2(n16157), .ZN(n9896) );
  NOR2_X1 U12693 ( .A1(n16527), .A2(n17493), .ZN(n9897) );
  AND2_X1 U12694 ( .A1(n14171), .A2(n14041), .ZN(n9898) );
  OR2_X1 U12695 ( .A1(n10435), .A2(n10434), .ZN(n10840) );
  AND2_X1 U12696 ( .A1(n10138), .A2(n14818), .ZN(n9899) );
  INV_X2 U12697 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n20098) );
  INV_X1 U12698 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n10013) );
  NOR2_X1 U12699 ( .A1(n17646), .A2(n16676), .ZN(n16631) );
  INV_X1 U12700 ( .A(n14582), .ZN(n10075) );
  INV_X1 U12701 ( .A(n14097), .ZN(n10158) );
  INV_X1 U12702 ( .A(n16467), .ZN(n10002) );
  NAND2_X1 U12703 ( .A1(n13695), .A2(n13957), .ZN(n11610) );
  AND2_X1 U12704 ( .A1(n12536), .A2(n12564), .ZN(n9900) );
  OR2_X1 U12705 ( .A1(n11520), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n9901) );
  INV_X1 U12706 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n10010) );
  INV_X1 U12707 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n10122) );
  INV_X1 U12708 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n10019) );
  INV_X1 U12709 ( .A(n15122), .ZN(n10150) );
  AND2_X1 U12710 ( .A1(n14370), .A2(n14379), .ZN(n9903) );
  NAND2_X1 U12711 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n10150), .ZN(
        n10149) );
  INV_X1 U12712 ( .A(n10236), .ZN(n10186) );
  INV_X1 U12713 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n10049) );
  INV_X1 U12714 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n10037) );
  INV_X1 U12715 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n10040) );
  INV_X1 U12716 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n10112) );
  NAND3_X2 U12717 ( .A1(n18776), .A2(n18764), .A3(n18775), .ZN(n18091) );
  NOR3_X2 U12718 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18623), .A3(
        n18326), .ZN(n18298) );
  NOR3_X4 U12719 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n18326), .ZN(n18351) );
  NAND3_X2 U12720 ( .A1(n9855), .A2(n11230), .A3(n9836), .ZN(n11252) );
  AND2_X2 U12721 ( .A1(n12722), .A2(n9839), .ZN(n13894) );
  NOR2_X2 U12722 ( .A1(n11265), .A2(n11256), .ZN(n11597) );
  NAND3_X1 U12723 ( .A1(n9908), .A2(n11255), .A3(n9907), .ZN(n11265) );
  NAND2_X1 U12724 ( .A1(n11261), .A2(n20122), .ZN(n9907) );
  NAND3_X1 U12725 ( .A1(n13731), .A2(n12708), .A3(n13823), .ZN(n13822) );
  NAND2_X1 U12726 ( .A1(n14543), .A2(n12838), .ZN(n12660) );
  NAND2_X2 U12727 ( .A1(n12663), .A2(n11340), .ZN(n11388) );
  NAND2_X1 U12728 ( .A1(n11336), .A2(n12662), .ZN(n12663) );
  OAI22_X2 U12729 ( .A1(n13437), .A2(P1_STATE2_REG_0__SCAN_IN), .B1(n11411), 
        .B2(n11362), .ZN(n9909) );
  NAND2_X1 U12730 ( .A1(n9910), .A2(n20151), .ZN(n13609) );
  NAND3_X1 U12731 ( .A1(n20151), .A2(n9910), .A3(n20098), .ZN(n9944) );
  XNOR2_X2 U12732 ( .A(n9805), .B(n10685), .ZN(n10682) );
  NAND2_X1 U12733 ( .A1(n9913), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n9914) );
  NAND2_X1 U12734 ( .A1(n10775), .A2(n10774), .ZN(n10776) );
  OAI21_X1 U12735 ( .B1(n10771), .B2(n10229), .A(n10767), .ZN(n9915) );
  NAND2_X2 U12736 ( .A1(n16107), .A2(n10804), .ZN(n15095) );
  NAND2_X1 U12737 ( .A1(n9920), .A2(n10776), .ZN(n15105) );
  OAI21_X1 U12738 ( .B1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n15344), .A(
        n9920), .ZN(n16115) );
  NAND4_X1 U12739 ( .A1(n9923), .A2(n9922), .A3(n9921), .A4(n9868), .ZN(n10620) );
  NAND3_X1 U12740 ( .A1(n9804), .A2(n10671), .A3(n9925), .ZN(n9924) );
  OAI21_X1 U12741 ( .B1(n13791), .B2(n11060), .A(n14641), .ZN(n11033) );
  OR2_X2 U12742 ( .A1(n12249), .A2(n9845), .ZN(n15227) );
  NAND2_X2 U12743 ( .A1(n18739), .A2(n18745), .ZN(n16789) );
  INV_X2 U12744 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n18745) );
  NOR2_X1 U12745 ( .A1(n17442), .A2(n9932), .ZN(n16299) );
  NOR2_X2 U12746 ( .A1(n17443), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17442) );
  NAND4_X1 U12747 ( .A1(n9865), .A2(n9936), .A3(n11814), .A4(n11816), .ZN(
        n9935) );
  NAND2_X1 U12748 ( .A1(n12286), .A2(n12285), .ZN(n12289) );
  AND2_X2 U12749 ( .A1(n11766), .A2(n9943), .ZN(n12286) );
  NAND2_X1 U12750 ( .A1(n11767), .A2(n11524), .ZN(n9943) );
  NAND3_X1 U12751 ( .A1(n10179), .A2(n14439), .A3(n14318), .ZN(n11767) );
  NAND2_X1 U12752 ( .A1(n9944), .A2(n11299), .ZN(n11370) );
  NAND2_X1 U12753 ( .A1(n14396), .A2(n14397), .ZN(n9946) );
  NAND2_X2 U12754 ( .A1(n11525), .A2(n14358), .ZN(n14354) );
  NAND2_X4 U12755 ( .A1(n11494), .A2(n11505), .ZN(n14352) );
  NOR2_X2 U12756 ( .A1(n9952), .A2(n10607), .ZN(n19153) );
  XNOR2_X2 U12757 ( .A(n9953), .B(n10973), .ZN(n12304) );
  AOI21_X1 U12758 ( .B1(n9953), .B2(n10973), .A(n10972), .ZN(n13854) );
  NAND2_X1 U12759 ( .A1(n15014), .A2(n9975), .ZN(n9967) );
  NAND2_X1 U12760 ( .A1(n15014), .A2(n9969), .ZN(n9968) );
  OAI211_X1 U12761 ( .C1(n15014), .C2(n9976), .A(n9974), .B(n9967), .ZN(n12270) );
  OAI211_X1 U12762 ( .C1(n15014), .C2(n9970), .A(n12266), .B(n9968), .ZN(
        P2_U3025) );
  NOR2_X1 U12763 ( .A1(n16713), .A2(n17533), .ZN(n9984) );
  NAND2_X1 U12764 ( .A1(n9985), .A2(n9983), .ZN(n9986) );
  NAND2_X1 U12765 ( .A1(n16563), .A2(n9993), .ZN(n9985) );
  INV_X1 U12766 ( .A(n16713), .ZN(n9993) );
  INV_X1 U12767 ( .A(n9988), .ZN(n16562) );
  INV_X1 U12768 ( .A(n9986), .ZN(n16551) );
  NAND2_X1 U12769 ( .A1(n16537), .A2(n9993), .ZN(n9991) );
  INV_X1 U12770 ( .A(n16466), .ZN(n10003) );
  INV_X1 U12771 ( .A(n11895), .ZN(n10014) );
  NOR2_X1 U12772 ( .A1(n10241), .A2(n18742), .ZN(n17779) );
  INV_X1 U12773 ( .A(n17471), .ZN(n10020) );
  OR2_X2 U12774 ( .A1(n17691), .A2(n10021), .ZN(n17639) );
  OR2_X1 U12775 ( .A1(n16309), .A2(n10023), .ZN(n17434) );
  INV_X1 U12776 ( .A(n17433), .ZN(n10023) );
  INV_X2 U12777 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18739) );
  INV_X2 U12778 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n18732) );
  NAND2_X1 U12779 ( .A1(n10026), .A2(n10025), .ZN(P2_U2825) );
  NAND3_X1 U12780 ( .A1(n12127), .A2(n18999), .A3(n10027), .ZN(n10026) );
  NAND2_X1 U12781 ( .A1(n10028), .A2(n12126), .ZN(n10027) );
  INV_X1 U12782 ( .A(n15947), .ZN(n10028) );
  NAND2_X1 U12783 ( .A1(n18840), .A2(n18873), .ZN(n18828) );
  NAND2_X1 U12784 ( .A1(n18841), .A2(n18842), .ZN(n18840) );
  NAND2_X1 U12785 ( .A1(n18853), .A2(n12116), .ZN(n18841) );
  NAND2_X1 U12786 ( .A1(n18854), .A2(n18855), .ZN(n18853) );
  AND2_X2 U12787 ( .A1(n20122), .A2(n20113), .ZN(n11709) );
  NAND2_X1 U12788 ( .A1(n13740), .A2(n10050), .ZN(n15921) );
  INV_X1 U12789 ( .A(n14148), .ZN(n10052) );
  NOR3_X2 U12790 ( .A1(n14008), .A2(n14154), .A3(n14157), .ZN(n14148) );
  NOR2_X2 U12791 ( .A1(n10052), .A2(n10051), .ZN(n11710) );
  INV_X1 U12792 ( .A(n10065), .ZN(n14678) );
  INV_X1 U12793 ( .A(n14689), .ZN(n10068) );
  NAND2_X1 U12794 ( .A1(n13717), .A2(n9842), .ZN(n14748) );
  NOR2_X2 U12795 ( .A1(n15238), .A2(n14724), .ZN(n14723) );
  NAND2_X1 U12796 ( .A1(n10801), .A2(n10082), .ZN(n11056) );
  NAND2_X1 U12797 ( .A1(n10083), .A2(n10768), .ZN(n10801) );
  NAND2_X1 U12798 ( .A1(n9771), .A2(n10840), .ZN(n10730) );
  OAI21_X1 U12799 ( .B1(n14899), .B2(n10089), .A(n10087), .ZN(n14946) );
  NAND2_X1 U12800 ( .A1(n14899), .A2(n10087), .ZN(n10086) );
  CLKBUF_X1 U12801 ( .A(n10092), .Z(n10090) );
  NAND2_X1 U12802 ( .A1(n12129), .A2(n10111), .ZN(n14865) );
  NAND2_X1 U12803 ( .A1(n12129), .A2(n12128), .ZN(n12224) );
  NAND2_X1 U12804 ( .A1(n11067), .A2(n11065), .ZN(n11079) );
  NAND2_X1 U12805 ( .A1(n12241), .A2(n10117), .ZN(n14878) );
  NAND2_X1 U12806 ( .A1(n12241), .A2(n14863), .ZN(n14868) );
  NOR2_X4 U12807 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15391) );
  AND2_X2 U12808 ( .A1(n13504), .A2(n13503), .ZN(n10826) );
  NOR2_X1 U12809 ( .A1(n14780), .A2(n14567), .ZN(n14762) );
  OR2_X2 U12810 ( .A1(n14780), .A2(n10126), .ZN(n14760) );
  INV_X1 U12811 ( .A(n12168), .ZN(n10129) );
  NAND2_X1 U12812 ( .A1(n13724), .A2(n9883), .ZN(n15268) );
  NAND2_X2 U12813 ( .A1(n13419), .A2(n10136), .ZN(n15310) );
  NOR2_X2 U12814 ( .A1(n15310), .A2(n15311), .ZN(n13618) );
  NAND2_X1 U12815 ( .A1(n14830), .A2(n9899), .ZN(n14817) );
  NAND4_X1 U12816 ( .A1(n10289), .A2(n10286), .A3(n10287), .A4(n10288), .ZN(
        n10142) );
  NAND4_X1 U12817 ( .A1(n10285), .A2(n10283), .A3(n10282), .A4(n10284), .ZN(
        n10144) );
  OAI21_X1 U12818 ( .B1(n10148), .B2(n15104), .A(n16108), .ZN(n10146) );
  NAND2_X1 U12819 ( .A1(n13894), .A2(n10152), .ZN(n13197) );
  INV_X1 U12820 ( .A(n13197), .ZN(n12785) );
  NAND2_X1 U12821 ( .A1(n9861), .A2(n14117), .ZN(n10159) );
  CLKBUF_X1 U12822 ( .A(n10159), .Z(n10155) );
  INV_X1 U12823 ( .A(n12813), .ZN(n10160) );
  AND2_X1 U12824 ( .A1(n14004), .A2(n10166), .ZN(n13169) );
  NAND3_X1 U12825 ( .A1(n10174), .A2(n15652), .A3(n9885), .ZN(n10173) );
  NAND2_X1 U12826 ( .A1(n10177), .A2(n10178), .ZN(n10176) );
  INV_X1 U12827 ( .A(n9813), .ZN(n10177) );
  NAND2_X1 U12828 ( .A1(n14534), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n14536) );
  NAND2_X2 U12829 ( .A1(n13413), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13412) );
  NAND2_X1 U12830 ( .A1(n11375), .A2(n11374), .ZN(n10178) );
  NAND4_X1 U12831 ( .A1(n11251), .A2(n11253), .A3(n9772), .A4(n11252), .ZN(
        n11261) );
  NAND2_X1 U12832 ( .A1(n14354), .A2(n14455), .ZN(n10180) );
  OAI21_X2 U12833 ( .B1(n14368), .B2(n10185), .A(n10184), .ZN(n11526) );
  INV_X1 U12834 ( .A(n11438), .ZN(n10193) );
  NAND2_X1 U12835 ( .A1(n20033), .A2(n10187), .ZN(n10189) );
  NAND3_X1 U12836 ( .A1(n10189), .A2(n11487), .A3(n10188), .ZN(n11490) );
  OAI211_X1 U12837 ( .C1(n20033), .C2(n10192), .A(n10190), .B(n10191), .ZN(
        n15787) );
  NAND2_X1 U12838 ( .A1(n10193), .A2(n15794), .ZN(n10190) );
  INV_X1 U12839 ( .A(n15794), .ZN(n10192) );
  NOR2_X1 U12840 ( .A1(n10203), .A2(n14352), .ZN(n10196) );
  INV_X1 U12841 ( .A(n10204), .ZN(n10201) );
  INV_X1 U12842 ( .A(n10203), .ZN(n10202) );
  NOR2_X1 U12843 ( .A1(n11522), .A2(n11524), .ZN(n10203) );
  INV_X1 U12844 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n10205) );
  NAND2_X2 U12845 ( .A1(n12311), .A2(n10482), .ZN(n10497) );
  NAND2_X1 U12846 ( .A1(n12568), .A2(n10219), .ZN(n10217) );
  NAND2_X1 U12847 ( .A1(n12570), .A2(n12568), .ZN(n14692) );
  NAND2_X1 U12848 ( .A1(n10217), .A2(n12570), .ZN(n10218) );
  NAND2_X1 U12849 ( .A1(n14034), .A2(n14035), .ZN(n14020) );
  NAND2_X1 U12850 ( .A1(n10771), .A2(n10774), .ZN(n10767) );
  OR2_X1 U12851 ( .A1(n13169), .A2(n13170), .ZN(n13172) );
  NOR2_X1 U12852 ( .A1(n10410), .A2(n10409), .ZN(n10831) );
  INV_X1 U12853 ( .A(n10479), .ZN(n12218) );
  BUF_X1 U12854 ( .A(n11252), .Z(n11288) );
  INV_X1 U12855 ( .A(n13620), .ZN(n12680) );
  NAND2_X1 U12856 ( .A1(n12313), .A2(n12326), .ZN(n12318) );
  XNOR2_X1 U12857 ( .A(n10559), .B(n10560), .ZN(n10592) );
  INV_X2 U12858 ( .A(n10962), .ZN(n10540) );
  NAND2_X2 U12859 ( .A1(n10545), .A2(n13348), .ZN(n10962) );
  AOI22_X1 U12860 ( .A1(n10391), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12622), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10335) );
  AND3_X4 U12861 ( .A1(n10267), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n12469) );
  INV_X2 U12862 ( .A(n14298), .ZN(n14294) );
  AND2_X2 U12863 ( .A1(n13155), .A2(n13703), .ZN(n19966) );
  INV_X1 U12864 ( .A(n14213), .ZN(n13156) );
  AND2_X1 U12865 ( .A1(n17694), .A2(n17788), .ZN(n10220) );
  AND2_X1 U12866 ( .A1(n10554), .A2(n10557), .ZN(n10221) );
  NAND2_X1 U12867 ( .A1(n10441), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10535) );
  INV_X1 U12868 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n15386) );
  INV_X1 U12869 ( .A(n10807), .ZN(n12165) );
  NOR2_X1 U12870 ( .A1(n11844), .A2(n11843), .ZN(n10224) );
  OR2_X1 U12871 ( .A1(n15492), .A2(n16965), .ZN(n10225) );
  AND2_X1 U12872 ( .A1(n10738), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n10227) );
  AND3_X1 U12873 ( .A1(n11875), .A2(n10225), .A3(n11874), .ZN(n10228) );
  OR2_X1 U12874 ( .A1(n13528), .A2(n13527), .ZN(n20025) );
  INV_X1 U12875 ( .A(n12673), .ZN(n12893) );
  NAND2_X2 U12876 ( .A1(n14294), .A2(n13705), .ZN(n14296) );
  AND2_X1 U12877 ( .A1(n10774), .A2(n10772), .ZN(n10229) );
  OR2_X1 U12878 ( .A1(n10849), .A2(n14919), .ZN(n10230) );
  AND2_X1 U12879 ( .A1(n12284), .A2(n11768), .ZN(n10231) );
  AND2_X1 U12880 ( .A1(n10569), .A2(n10568), .ZN(n10233) );
  AND2_X1 U12881 ( .A1(n11524), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n10234) );
  AND3_X1 U12882 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n10236) );
  OR2_X1 U12883 ( .A1(n19718), .A2(P2_STATE_REG_0__SCAN_IN), .ZN(n19856) );
  OR2_X1 U12884 ( .A1(n10604), .A2(n10603), .ZN(n10237) );
  AND2_X1 U12885 ( .A1(n14933), .A2(n14945), .ZN(n10238) );
  AND2_X2 U12886 ( .A1(n19996), .A2(n19970), .ZN(n19993) );
  AND4_X1 U12887 ( .A1(n10649), .A2(n10648), .A3(n10647), .A4(n10646), .ZN(
        n10239) );
  NOR2_X1 U12888 ( .A1(n20485), .A2(n20451), .ZN(n10240) );
  NOR2_X1 U12889 ( .A1(n20485), .A2(n20311), .ZN(n10242) );
  NAND2_X1 U12890 ( .A1(n18117), .A2(n18008), .ZN(n18072) );
  OR2_X1 U12891 ( .A1(n18872), .A2(n18875), .ZN(n10243) );
  OR2_X1 U12892 ( .A1(n17346), .A2(n18117), .ZN(n10244) );
  AND3_X1 U12893 ( .A1(n12089), .A2(n12088), .A3(n12087), .ZN(n10245) );
  NOR2_X1 U12894 ( .A1(n17781), .A2(n17768), .ZN(n17532) );
  INV_X1 U12895 ( .A(n17532), .ZN(n17500) );
  AND2_X1 U12896 ( .A1(n9779), .A2(n10511), .ZN(n10246) );
  OR2_X1 U12897 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n12695) );
  INV_X1 U12898 ( .A(n14070), .ZN(n14087) );
  AND2_X2 U12899 ( .A1(n11138), .A2(n13594), .ZN(n11233) );
  OAI22_X1 U12900 ( .A1(n9775), .A2(n10566), .B1(n15386), .B2(n10565), .ZN(
        n10567) );
  NAND2_X1 U12901 ( .A1(n10634), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n10635) );
  NAND2_X1 U12902 ( .A1(n10539), .A2(n10367), .ZN(n10519) );
  NAND2_X1 U12903 ( .A1(n11533), .A2(n11532), .ZN(n11565) );
  INV_X1 U12904 ( .A(n11538), .ZN(n11546) );
  INV_X1 U12905 ( .A(n12513), .ZN(n12514) );
  AOI22_X1 U12906 ( .A1(n12622), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10382), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10288) );
  AOI22_X1 U12907 ( .A1(n9820), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10391), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10285) );
  NAND2_X1 U12908 ( .A1(n10478), .A2(n10367), .ZN(n10481) );
  AOI22_X1 U12909 ( .A1(n10383), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n9818), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10270) );
  INV_X1 U12910 ( .A(n14118), .ZN(n12784) );
  OR2_X1 U12911 ( .A1(n11577), .A2(n11430), .ZN(n11431) );
  OR2_X1 U12912 ( .A1(n11474), .A2(n11473), .ZN(n11496) );
  AND2_X1 U12913 ( .A1(n10488), .A2(n9866), .ZN(n10489) );
  AOI22_X1 U12914 ( .A1(n10381), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n9819), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10316) );
  OAI21_X1 U12915 ( .B1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n11343), .A(
        n11342), .ZN(n11344) );
  OR2_X1 U12916 ( .A1(n14023), .A2(n14170), .ZN(n13027) );
  INV_X1 U12917 ( .A(n11457), .ZN(n11482) );
  INV_X1 U12918 ( .A(n14184), .ZN(n12920) );
  NAND2_X1 U12919 ( .A1(n11432), .A2(n11431), .ZN(n11440) );
  OR2_X1 U12920 ( .A1(n11360), .A2(n11359), .ZN(n11363) );
  AND2_X1 U12921 ( .A1(n10371), .A2(n10480), .ZN(n10351) );
  XNOR2_X1 U12922 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n10443) );
  INV_X1 U12923 ( .A(n10381), .ZN(n12421) );
  AOI22_X1 U12924 ( .A1(n12622), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10382), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10276) );
  OR2_X1 U12925 ( .A1(n11933), .A2(n11934), .ZN(n11926) );
  NAND2_X1 U12926 ( .A1(n17065), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n11874) );
  OR2_X1 U12927 ( .A1(n11570), .A2(n11569), .ZN(n11592) );
  NAND2_X1 U12928 ( .A1(n11266), .A2(n20113), .ZN(n11720) );
  INV_X1 U12929 ( .A(n13103), .ZN(n13104) );
  NOR2_X1 U12930 ( .A1(n11253), .A2(n20623), .ZN(n12673) );
  NOR2_X1 U12931 ( .A1(n11267), .A2(n20122), .ZN(n11269) );
  NAND2_X1 U12932 ( .A1(n9801), .A2(n11287), .ZN(n20151) );
  NAND2_X1 U12933 ( .A1(n11042), .A2(n11041), .ZN(n11045) );
  OR2_X1 U12934 ( .A1(n12457), .A2(n12456), .ZN(n12488) );
  AND2_X1 U12935 ( .A1(n16217), .A2(n9779), .ZN(n13373) );
  NAND2_X1 U12936 ( .A1(n14900), .A2(n15155), .ZN(n14901) );
  OR2_X1 U12937 ( .A1(n18927), .A2(n10849), .ZN(n11096) );
  INV_X1 U12938 ( .A(n19355), .ZN(n10695) );
  OAI21_X1 U12939 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n18732), .A(
        n11926), .ZN(n11927) );
  INV_X1 U12940 ( .A(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n16969) );
  INV_X1 U12941 ( .A(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17034) );
  INV_X1 U12942 ( .A(n11836), .ZN(n11840) );
  INV_X1 U12943 ( .A(n11908), .ZN(n11909) );
  INV_X1 U12944 ( .A(n9817), .ZN(n12034) );
  NOR2_X1 U12945 ( .A1(n18135), .A2(n15552), .ZN(n15555) );
  INV_X1 U12946 ( .A(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17052) );
  AND2_X1 U12947 ( .A1(n11593), .A2(n11592), .ZN(n13282) );
  NAND2_X1 U12948 ( .A1(n12292), .A2(n12291), .ZN(n12293) );
  OR2_X1 U12949 ( .A1(n13205), .A2(n14303), .ZN(n13207) );
  AND2_X1 U12950 ( .A1(n20623), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n13960) );
  INV_X1 U12951 ( .A(n14394), .ZN(n14395) );
  AND2_X1 U12952 ( .A1(n11746), .A2(n11733), .ZN(n13565) );
  OAI21_X1 U12953 ( .B1(n11591), .B2(n11577), .A(n11576), .ZN(n11581) );
  INV_X1 U12954 ( .A(n20308), .ZN(n20339) );
  INV_X1 U12955 ( .A(n20539), .ZN(n20620) );
  INV_X1 U12956 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20367) );
  OR2_X1 U12957 ( .A1(n10860), .A2(n10859), .ZN(n19028) );
  INV_X1 U12958 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n12091) );
  AND2_X1 U12959 ( .A1(n14867), .A2(n15241), .ZN(n15230) );
  OAI21_X1 U12960 ( .B1(n11056), .B2(n11060), .A(n18961), .ZN(n11057) );
  NOR2_X1 U12961 ( .A1(n10398), .A2(n10397), .ZN(n10814) );
  NAND2_X1 U12962 ( .A1(n12319), .A2(n12326), .ZN(n12321) );
  OAI22_X1 U12963 ( .A1(n18739), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(
        n18594), .B2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12038) );
  INV_X2 U12964 ( .A(n17051), .ZN(n15497) );
  INV_X1 U12965 ( .A(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n16894) );
  NOR2_X1 U12966 ( .A1(n18576), .A2(n11789), .ZN(n11833) );
  XOR2_X1 U12967 ( .A(n17288), .B(n11868), .Z(n11884) );
  NAND2_X1 U12968 ( .A1(n18582), .A2(n18589), .ZN(n17984) );
  INV_X1 U12969 ( .A(n17299), .ZN(n12058) );
  AOI21_X1 U12970 ( .B1(n15528), .B2(n18613), .A(n18758), .ZN(n15529) );
  AOI21_X2 U12971 ( .B1(n12022), .B2(n12021), .A(n16433), .ZN(n18562) );
  NOR2_X1 U12972 ( .A1(n13067), .A2(n15672), .ZN(n13068) );
  AND2_X1 U12973 ( .A1(n13013), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n13022) );
  AND2_X1 U12974 ( .A1(n13973), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13216) );
  OAI21_X1 U12975 ( .B1(n11345), .B2(n13558), .A(n11396), .ZN(n20254) );
  INV_X1 U12976 ( .A(n19937), .ZN(n19899) );
  AND2_X1 U12977 ( .A1(n11678), .A2(n11677), .ZN(n14186) );
  OR2_X1 U12978 ( .A1(n13702), .A2(n13701), .ZN(n13704) );
  NAND2_X1 U12979 ( .A1(n12880), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n12912) );
  INV_X1 U12980 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n12809) );
  NOR2_X1 U12981 ( .A1(n12738), .A2(n14132), .ZN(n12752) );
  INV_X1 U12982 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12682) );
  OR2_X1 U12983 ( .A1(n15813), .A2(n14370), .ZN(n14500) );
  AND2_X1 U12984 ( .A1(n11663), .A2(n11662), .ZN(n14099) );
  OR2_X1 U12985 ( .A1(n13173), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20081) );
  NOR2_X1 U12986 ( .A1(n20484), .A2(n20259), .ZN(n20429) );
  NOR2_X1 U12987 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20458) );
  OR2_X1 U12988 ( .A1(n20629), .A2(n20096), .ZN(n20634) );
  AND2_X1 U12989 ( .A1(n12116), .A2(n14575), .ZN(n18895) );
  INV_X1 U12990 ( .A(n18989), .ZN(n18973) );
  OR2_X1 U12991 ( .A1(n12563), .A2(n12562), .ZN(n14683) );
  INV_X1 U12992 ( .A(n13680), .ZN(n12340) );
  OR2_X1 U12993 ( .A1(n10764), .A2(n10763), .ZN(n10848) );
  OAI21_X1 U12994 ( .B1(n12646), .B2(n12645), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n12647) );
  AND2_X1 U12995 ( .A1(n15336), .A2(n10510), .ZN(n16136) );
  AND3_X1 U12996 ( .A1(n10863), .A2(n10862), .A3(n10861), .ZN(n13484) );
  NAND2_X1 U12997 ( .A1(n10464), .A2(n10461), .ZN(n16217) );
  AND2_X1 U12998 ( .A1(n19147), .A2(n19146), .ZN(n19192) );
  OR2_X1 U12999 ( .A1(n19547), .A2(n19541), .ZN(n19592) );
  INV_X1 U13000 ( .A(n16432), .ZN(n18580) );
  NOR2_X1 U13001 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n16602), .ZN(n16587) );
  NOR2_X1 U13002 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n16672), .ZN(n16656) );
  NOR2_X1 U13003 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n16715), .ZN(n16702) );
  NOR2_X1 U13004 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n16741), .ZN(n16722) );
  INV_X1 U13005 ( .A(n16783), .ZN(n16802) );
  INV_X1 U13006 ( .A(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n21058) );
  NOR3_X1 U13007 ( .A1(n18760), .A2(n17308), .A3(n15635), .ZN(n15636) );
  INV_X1 U13008 ( .A(n16632), .ZN(n17622) );
  INV_X1 U13009 ( .A(n11884), .ZN(n11886) );
  NAND2_X1 U13010 ( .A1(n17712), .A2(n11898), .ZN(n11901) );
  INV_X1 U13011 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n11881) );
  INV_X1 U13012 ( .A(n15529), .ZN(n17307) );
  INV_X1 U13013 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18594) );
  AOI211_X1 U13014 ( .C1(n17053), .C2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A(
        n11978), .B(n11977), .ZN(n18125) );
  AOI22_X1 U13015 ( .A1(n18552), .A2(n18551), .B1(n18556), .B2(n15566), .ZN(
        n18560) );
  INV_X1 U13016 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n20698) );
  AND2_X1 U13017 ( .A1(n13068), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n13103) );
  AND2_X1 U13018 ( .A1(n13022), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n13044) );
  NAND2_X1 U13019 ( .A1(n13747), .A2(n13209), .ZN(n19926) );
  AND2_X1 U13020 ( .A1(n19924), .A2(n13208), .ZN(n19912) );
  AND2_X1 U13021 ( .A1(n19924), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n19940) );
  AND2_X1 U13022 ( .A1(n13747), .A2(n13212), .ZN(n19948) );
  OAI22_X1 U13023 ( .A1(n13994), .A2(n15737), .B1(n19966), .B2(n13157), .ZN(
        n13158) );
  INV_X1 U13024 ( .A(n14265), .ZN(n14285) );
  NAND2_X1 U13025 ( .A1(n13704), .A2(n13703), .ZN(n14298) );
  INV_X1 U13026 ( .A(n13688), .ZN(n20030) );
  INV_X1 U13027 ( .A(n15695), .ZN(n14375) );
  AOI21_X1 U13028 ( .B1(n10158), .B2(n9832), .A(n14098), .ZN(n14414) );
  NAND2_X1 U13029 ( .A1(n12780), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n12808) );
  NAND2_X1 U13030 ( .A1(n12694), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12702) );
  INV_X1 U13031 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n20044) );
  OR2_X1 U13032 ( .A1(n14467), .A2(n11757), .ZN(n14452) );
  NOR2_X1 U13033 ( .A1(n15841), .A2(n11739), .ZN(n15816) );
  AND2_X1 U13034 ( .A1(n11609), .A2(n13703), .ZN(n11746) );
  INV_X1 U13035 ( .A(n15917), .ZN(n15900) );
  INV_X1 U13036 ( .A(n20080), .ZN(n20053) );
  NOR2_X1 U13037 ( .A1(n15872), .A2(n14537), .ZN(n20071) );
  INV_X1 U13038 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13558) );
  OAI22_X1 U13039 ( .A1(n20110), .A2(n20109), .B1(n20370), .B2(n20256), .ZN(
        n20147) );
  INV_X1 U13040 ( .A(n20172), .ZN(n20175) );
  OAI22_X1 U13041 ( .A1(n20186), .A2(n20185), .B1(n20370), .B2(n20309), .ZN(
        n20209) );
  OAI21_X1 U13042 ( .B1(n10242), .B2(n20260), .A(n20580), .ZN(n20278) );
  AND2_X1 U13043 ( .A1(n20766), .A2(n20547), .ZN(n20333) );
  AND2_X1 U13044 ( .A1(n20766), .A2(n20569), .ZN(n20361) );
  OAI211_X1 U13045 ( .C1(n10240), .C2(n20493), .A(n20429), .B(n20375), .ZN(
        n20392) );
  INV_X1 U13046 ( .A(n20479), .ZN(n20366) );
  AND2_X1 U13047 ( .A1(n20759), .A2(n20569), .ZN(n20475) );
  INV_X1 U13048 ( .A(n20495), .ZN(n20532) );
  OAI211_X1 U13049 ( .C1(n20494), .C2(n20493), .A(n20580), .B(n20492), .ZN(
        n20533) );
  INV_X1 U13050 ( .A(n20575), .ZN(n20613) );
  INV_X1 U13051 ( .A(n20530), .ZN(n20678) );
  INV_X1 U13052 ( .A(n20748), .ZN(n20742) );
  INV_X1 U13053 ( .A(n18982), .ZN(n18991) );
  INV_X1 U13054 ( .A(n18994), .ZN(n18950) );
  AND2_X1 U13055 ( .A1(n19838), .A2(n12138), .ZN(n18989) );
  AND2_X1 U13056 ( .A1(n16212), .A2(n19840), .ZN(n13253) );
  NOR2_X1 U13057 ( .A1(n19796), .A2(n18989), .ZN(n19002) );
  OR2_X1 U13058 ( .A1(n10898), .A2(n10897), .ZN(n19016) );
  INV_X1 U13059 ( .A(n19031), .ZN(n19038) );
  OR2_X1 U13060 ( .A1(n12410), .A2(n12409), .ZN(n14730) );
  INV_X1 U13061 ( .A(n14841), .ZN(n16047) );
  INV_X1 U13062 ( .A(n19817), .ZN(n19381) );
  INV_X1 U13063 ( .A(n13344), .ZN(n19136) );
  INV_X1 U13064 ( .A(n12647), .ZN(n13781) );
  INV_X1 U13065 ( .A(n16055), .ZN(n16120) );
  INV_X1 U13066 ( .A(n21140), .ZN(n11126) );
  INV_X1 U13067 ( .A(n9889), .ZN(n18976) );
  NOR2_X1 U13068 ( .A1(n16187), .A2(n15335), .ZN(n15329) );
  INV_X1 U13069 ( .A(n9889), .ZN(n16186) );
  NAND2_X1 U13070 ( .A1(n10475), .A2(n10474), .ZN(n11125) );
  INV_X1 U13071 ( .A(n16181), .ZN(n21133) );
  INV_X1 U13072 ( .A(n19647), .ZN(n19268) );
  NAND2_X1 U13073 ( .A1(n16217), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n16244) );
  NOR2_X2 U13074 ( .A1(n19414), .A2(n19352), .ZN(n19237) );
  INV_X1 U13075 ( .A(n19246), .ZN(n19256) );
  INV_X1 U13076 ( .A(n19261), .ZN(n19289) );
  INV_X1 U13077 ( .A(n19313), .ZN(n19302) );
  NAND2_X1 U13078 ( .A1(n19788), .A2(n19381), .ZN(n19352) );
  INV_X1 U13079 ( .A(n19432), .ZN(n19438) );
  AND2_X1 U13080 ( .A1(n19479), .A2(n19476), .ZN(n19499) );
  NOR2_X2 U13081 ( .A1(n19537), .A2(n19482), .ZN(n19531) );
  INV_X1 U13082 ( .A(n19669), .ZN(n19568) );
  INV_X1 U13083 ( .A(n19636), .ZN(n19619) );
  NAND2_X1 U13084 ( .A1(n19802), .A2(n19146), .ZN(n19536) );
  NOR2_X2 U13085 ( .A1(n14769), .A2(n13780), .ZN(n19178) );
  INV_X1 U13086 ( .A(n19835), .ZN(n19844) );
  NOR2_X1 U13087 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16532), .ZN(n16520) );
  NOR2_X1 U13088 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n16555), .ZN(n16540) );
  NOR2_X1 U13089 ( .A1(n16545), .A2(n16619), .ZN(n16581) );
  NOR2_X1 U13090 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n16626), .ZN(n16607) );
  NOR2_X1 U13091 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n16693), .ZN(n16685) );
  NOR2_X2 U13092 ( .A1(n18716), .A2(n16804), .ZN(n16773) );
  AND3_X2 U13093 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .A3(n16859), .ZN(n16848) );
  NAND2_X1 U13094 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17118), .ZN(n17115) );
  OAI21_X1 U13095 ( .B1(n15536), .B2(n15430), .A(n18611), .ZN(n15635) );
  NOR3_X1 U13096 ( .A1(n17291), .A2(n17351), .A3(n17232), .ZN(n17224) );
  INV_X1 U13097 ( .A(n17205), .ZN(n17230) );
  INV_X1 U13098 ( .A(n16970), .ZN(n17089) );
  INV_X2 U13099 ( .A(n18114), .ZN(n17308) );
  INV_X1 U13100 ( .A(n17591), .ZN(n17638) );
  INV_X1 U13101 ( .A(n18117), .ZN(n18760) );
  NOR3_X1 U13102 ( .A1(n18084), .A2(n17846), .A3(n17812), .ZN(n17872) );
  INV_X1 U13103 ( .A(n17274), .ZN(n15567) );
  INV_X1 U13104 ( .A(n17992), .ZN(n18015) );
  AOI21_X2 U13105 ( .B1(n15560), .B2(n15559), .A(n18619), .ZN(n18089) );
  NAND2_X1 U13106 ( .A1(n18764), .A2(n18112), .ZN(n18401) );
  NOR2_X1 U13107 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18716), .ZN(
        n18740) );
  OAI21_X1 U13108 ( .B1(n15538), .B2(n17307), .A(n15537), .ZN(n18586) );
  INV_X1 U13109 ( .A(n18248), .ZN(n18254) );
  INV_X1 U13110 ( .A(n18156), .ZN(n18486) );
  OR2_X1 U13111 ( .A1(n18760), .A2(n17346), .ZN(n18613) );
  NOR2_X1 U13112 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n13195), .ZN(n16397)
         );
  NAND2_X1 U13113 ( .A1(n13423), .A2(n13200), .ZN(n13528) );
  INV_X1 U13114 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n20574) );
  INV_X1 U13115 ( .A(n19948), .ZN(n19897) );
  INV_X1 U13116 ( .A(n19940), .ZN(n15730) );
  INV_X1 U13117 ( .A(n13158), .ZN(n13159) );
  NAND2_X1 U13118 ( .A1(n19966), .A2(n9790), .ZN(n14213) );
  INV_X1 U13119 ( .A(n14307), .ZN(n14228) );
  OR2_X1 U13120 ( .A1(n14045), .A2(n14060), .ZN(n15754) );
  OR2_X1 U13121 ( .A1(n14212), .A2(n14211), .ZN(n15769) );
  INV_X1 U13122 ( .A(n13723), .ZN(n13846) );
  OR2_X1 U13123 ( .A1(n14298), .A2(n13705), .ZN(n14297) );
  OR2_X1 U13124 ( .A1(n19996), .A2(n11266), .ZN(n19967) );
  NAND2_X1 U13125 ( .A1(n13423), .A2(n13422), .ZN(n19996) );
  INV_X1 U13126 ( .A(n20025), .ZN(n13688) );
  OAI21_X1 U13127 ( .B1(n14212), .B2(n14120), .A(n9832), .ZN(n14430) );
  INV_X1 U13128 ( .A(n20045), .ZN(n20041) );
  AOI21_X1 U13129 ( .B1(n11764), .B2(n20063), .A(n11763), .ZN(n11765) );
  NAND2_X1 U13130 ( .A1(n11746), .A2(n11613), .ZN(n15923) );
  INV_X1 U13131 ( .A(n20063), .ZN(n20083) );
  INV_X1 U13132 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20538) );
  INV_X1 U13133 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n13475) );
  NAND2_X1 U13134 ( .A1(n20219), .A2(n20366), .ZN(n20172) );
  NAND2_X1 U13135 ( .A1(n20219), .A2(n20547), .ZN(n20213) );
  NAND2_X1 U13136 ( .A1(n20219), .A2(n20569), .ZN(n20251) );
  NAND2_X1 U13137 ( .A1(n20219), .A2(n20450), .ZN(n20281) );
  NAND2_X1 U13138 ( .A1(n20766), .A2(n20366), .ZN(n20305) );
  AOI22_X1 U13139 ( .A1(n20315), .A2(n20312), .B1(n20310), .B2(n20484), .ZN(
        n20337) );
  NAND2_X1 U13140 ( .A1(n20766), .A2(n20450), .ZN(n20371) );
  NAND2_X1 U13141 ( .A1(n20759), .A2(n20366), .ZN(n20418) );
  AOI22_X1 U13142 ( .A1(n20427), .A2(n20424), .B1(n20423), .B2(n20422), .ZN(
        n20449) );
  NAND2_X1 U13143 ( .A1(n20759), .A2(n20450), .ZN(n20495) );
  AOI22_X1 U13144 ( .A1(n20491), .A2(n20488), .B1(n20484), .B2(n20483), .ZN(
        n20537) );
  OR2_X1 U13145 ( .A1(n20629), .A2(n20479), .ZN(n20568) );
  NAND2_X1 U13146 ( .A1(n20570), .A2(n20569), .ZN(n20684) );
  INV_X1 U13147 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n20493) );
  INV_X1 U13148 ( .A(n20757), .ZN(n20688) );
  INV_X1 U13149 ( .A(n20740), .ZN(n20796) );
  OR2_X1 U13150 ( .A1(n10953), .A2(n13254), .ZN(n13269) );
  NAND2_X1 U13151 ( .A1(n12269), .A2(n19840), .ZN(n18790) );
  INV_X1 U13152 ( .A(n15116), .ZN(n15951) );
  OR2_X1 U13153 ( .A1(n19838), .A2(n12219), .ZN(n18981) );
  INV_X1 U13154 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n18882) );
  OR2_X1 U13155 ( .A1(n19838), .A2(n12136), .ZN(n18994) );
  AND2_X1 U13156 ( .A1(n13349), .A2(n19840), .ZN(n19020) );
  AND2_X1 U13157 ( .A1(n12654), .A2(n12653), .ZN(n12655) );
  INV_X1 U13158 ( .A(n19083), .ZN(n19044) );
  OR2_X1 U13159 ( .A1(n19083), .A2(n10497), .ZN(n19079) );
  OR2_X1 U13160 ( .A1(n19121), .A2(n19131), .ZN(n19099) );
  INV_X1 U13161 ( .A(n19121), .ZN(n19133) );
  INV_X1 U13162 ( .A(n19143), .ZN(n13344) );
  INV_X1 U13163 ( .A(n12281), .ZN(n12282) );
  INV_X1 U13164 ( .A(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n16078) );
  INV_X1 U13165 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n16098) );
  OR2_X1 U13166 ( .A1(n18790), .A2(n9776), .ZN(n15067) );
  NAND2_X1 U13167 ( .A1(n16125), .A2(n19806), .ZN(n16088) );
  AND2_X1 U13168 ( .A1(n12265), .A2(n12264), .ZN(n12266) );
  NAND2_X1 U13169 ( .A1(n11127), .A2(n11126), .ZN(n11128) );
  NAND2_X1 U13170 ( .A1(n11125), .A2(n19828), .ZN(n16157) );
  NAND2_X1 U13171 ( .A1(n11125), .A2(n19827), .ZN(n21140) );
  INV_X1 U13172 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19821) );
  INV_X1 U13173 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n15547) );
  OR2_X1 U13174 ( .A1(n19414), .A2(n19314), .ZN(n19213) );
  OR2_X1 U13175 ( .A1(n19314), .A2(n19482), .ZN(n19246) );
  OR2_X1 U13176 ( .A1(n19352), .A2(n19482), .ZN(n19261) );
  INV_X1 U13177 ( .A(n19310), .ZN(n19305) );
  AOI211_X2 U13178 ( .C1(n19320), .C2(n19319), .A(n19322), .B(n19318), .ZN(
        n19351) );
  OR2_X1 U13179 ( .A1(n19352), .A2(n19642), .ZN(n19412) );
  OR2_X1 U13180 ( .A1(n19598), .A2(n19414), .ZN(n19432) );
  NAND2_X1 U13181 ( .A1(n19443), .A2(n19787), .ZN(n19503) );
  AOI21_X1 U13182 ( .B1(n19508), .B2(n19509), .A(n19507), .ZN(n19535) );
  OR2_X1 U13183 ( .A1(n19537), .A2(n19536), .ZN(n19636) );
  OR2_X1 U13184 ( .A1(n19598), .A2(n19642), .ZN(n19688) );
  AND2_X1 U13185 ( .A1(n16243), .A2(n16242), .ZN(n19707) );
  INV_X1 U13186 ( .A(n19783), .ZN(n19708) );
  CLKBUF_X1 U13187 ( .A(n19776), .Z(n19770) );
  NOR2_X1 U13188 ( .A1(n18554), .A2(n17345), .ZN(n18783) );
  INV_X1 U13189 ( .A(n12048), .ZN(n16417) );
  INV_X1 U13190 ( .A(n16776), .ZN(n16793) );
  INV_X1 U13191 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16676) );
  INV_X1 U13192 ( .A(n16773), .ZN(n16791) );
  NAND2_X1 U13193 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16863), .ZN(n16854) );
  AND2_X1 U13194 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16874), .ZN(n16868) );
  OR2_X1 U13195 ( .A1(n16950), .A2(n16949), .ZN(n16980) );
  AND3_X1 U13196 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(P3_EBX_REG_9__SCAN_IN), 
        .A3(n17069), .ZN(n17068) );
  INV_X1 U13197 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17133) );
  NOR2_X1 U13198 ( .A1(n17243), .A2(n17273), .ZN(n17266) );
  AOI211_X2 U13199 ( .C1(n17053), .C2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A(
        n11809), .B(n11808), .ZN(n17281) );
  INV_X1 U13200 ( .A(n17301), .ZN(n17298) );
  NAND2_X1 U13201 ( .A1(n17325), .A2(n17308), .ZN(n17324) );
  INV_X1 U13202 ( .A(n17325), .ZN(n17344) );
  INV_X1 U13203 ( .A(n17695), .ZN(n17659) );
  AOI22_X1 U13204 ( .A1(n17773), .A2(n17608), .B1(n17696), .B2(n17951), .ZN(
        n17680) );
  INV_X1 U13205 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n20959) );
  INV_X1 U13206 ( .A(n17773), .ZN(n17785) );
  INV_X1 U13207 ( .A(n18085), .ZN(n18046) );
  INV_X1 U13208 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n18001) );
  INV_X1 U13209 ( .A(n18082), .ZN(n18097) );
  INV_X1 U13210 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18169) );
  INV_X1 U13211 ( .A(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n18333) );
  INV_X1 U13212 ( .A(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n21054) );
  INV_X1 U13213 ( .A(n18527), .ZN(n18477) );
  INV_X1 U13214 ( .A(n18543), .ZN(n18539) );
  INV_X1 U13215 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n18726) );
  INV_X1 U13216 ( .A(n18713), .ZN(n18627) );
  INV_X1 U13217 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n18642) );
  NAND2_X1 U13218 ( .A1(n18642), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n18773) );
  OR4_X1 U13219 ( .A1(n13231), .A2(n13230), .A3(n13229), .A4(n13228), .ZN(
        P1_U2830) );
  OAI21_X1 U13220 ( .B1(n14317), .B2(n15923), .A(n11778), .ZN(P1_U3002) );
  NAND2_X1 U13221 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n19821), .ZN(
        n10263) );
  OAI21_X1 U13222 ( .B1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n19821), .A(
        n10263), .ZN(n10444) );
  INV_X1 U13223 ( .A(n10263), .ZN(n10247) );
  NAND2_X1 U13224 ( .A1(n10443), .A2(n10247), .ZN(n10249) );
  NAND2_X1 U13225 ( .A1(n19813), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10248) );
  NAND2_X1 U13226 ( .A1(n10249), .A2(n10248), .ZN(n10253) );
  XNOR2_X1 U13227 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n10252) );
  NAND2_X1 U13228 ( .A1(n10253), .A2(n10252), .ZN(n10251) );
  NAND2_X1 U13229 ( .A1(n19804), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10250) );
  XNOR2_X1 U13230 ( .A(n10256), .B(n10255), .ZN(n10424) );
  XNOR2_X1 U13231 ( .A(n10253), .B(n10252), .ZN(n10449) );
  NOR2_X1 U13232 ( .A1(n10330), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10254) );
  NOR2_X1 U13233 ( .A1(n21060), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n10257) );
  NOR3_X1 U13234 ( .A1(n10424), .A2(n10449), .A3(n10456), .ZN(n10264) );
  INV_X1 U13235 ( .A(n10264), .ZN(n10266) );
  INV_X1 U13236 ( .A(n10258), .ZN(n10260) );
  AND2_X1 U13237 ( .A1(n21060), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n10259) );
  NAND2_X1 U13238 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n15547), .ZN(
        n10261) );
  XNOR2_X1 U13239 ( .A(n10443), .B(n10263), .ZN(n10445) );
  AND2_X1 U13240 ( .A1(n10445), .A2(n10264), .ZN(n10265) );
  OAI21_X1 U13241 ( .B1(n10444), .B2(n10266), .A(n16212), .ZN(n10268) );
  INV_X1 U13242 ( .A(n10653), .ZN(n12402) );
  INV_X1 U13243 ( .A(n10271), .ZN(n15411) );
  AOI21_X1 U13244 ( .B1(n10271), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n16224) );
  AOI21_X1 U13245 ( .B1(n12402), .B2(n16224), .A(P2_FLUSH_REG_SCAN_IN), .ZN(
        n19816) );
  MUX2_X1 U13246 ( .A(n10268), .B(n19816), .S(P2_STATE2_REG_1__SCAN_IN), .Z(
        n19826) );
  INV_X1 U13247 ( .A(n19826), .ZN(n16249) );
  AND2_X4 U13248 ( .A1(n10269), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10383) );
  AND2_X4 U13249 ( .A1(n15391), .A2(n16194), .ZN(n10386) );
  INV_X2 U13250 ( .A(n10281), .ZN(n12612) );
  AOI22_X1 U13251 ( .A1(n9820), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n12612), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10274) );
  AND2_X4 U13252 ( .A1(n15391), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10385) );
  AND2_X4 U13253 ( .A1(n15401), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10381) );
  AOI22_X1 U13254 ( .A1(n10385), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n10381), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10273) );
  AND2_X4 U13255 ( .A1(n15390), .A2(n9816), .ZN(n12622) );
  AND2_X4 U13256 ( .A1(n15390), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10382) );
  AOI22_X1 U13257 ( .A1(n12622), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n10382), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10272) );
  NAND4_X1 U13258 ( .A1(n9862), .A2(n10274), .A3(n10273), .A4(n10272), .ZN(
        n10280) );
  AOI22_X1 U13259 ( .A1(n10383), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12469), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10275) );
  AOI22_X1 U13260 ( .A1(n10385), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10381), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10277) );
  NAND4_X1 U13261 ( .A1(n9863), .A2(n10278), .A3(n10277), .A4(n10276), .ZN(
        n10279) );
  INV_X2 U13262 ( .A(n10281), .ZN(n10391) );
  AOI22_X1 U13263 ( .A1(n12622), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n10382), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10284) );
  AOI22_X1 U13264 ( .A1(n10383), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n9818), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10283) );
  AOI22_X1 U13265 ( .A1(n10385), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10381), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10282) );
  AOI22_X1 U13266 ( .A1(n9821), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12612), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10289) );
  AOI22_X1 U13267 ( .A1(n10383), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9818), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10287) );
  AOI22_X1 U13268 ( .A1(n9819), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10381), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10286) );
  AOI22_X1 U13269 ( .A1(n10383), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12469), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10292) );
  AOI22_X1 U13270 ( .A1(n10385), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10381), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10291) );
  AOI22_X1 U13271 ( .A1(n12622), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10382), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10290) );
  NAND4_X1 U13272 ( .A1(n10293), .A2(n10292), .A3(n10291), .A4(n10290), .ZN(
        n10294) );
  NAND2_X1 U13273 ( .A1(n10294), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10301) );
  AOI22_X1 U13274 ( .A1(n10386), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12612), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10298) );
  AOI22_X1 U13275 ( .A1(n10385), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n10381), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10297) );
  AOI22_X1 U13276 ( .A1(n12622), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n10382), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10296) );
  AOI22_X1 U13277 ( .A1(n10383), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n9818), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10295) );
  NAND4_X1 U13278 ( .A1(n10298), .A2(n10297), .A3(n10296), .A4(n10295), .ZN(
        n10299) );
  NAND2_X1 U13279 ( .A1(n10299), .A2(n10330), .ZN(n10300) );
  NAND2_X2 U13280 ( .A1(n10301), .A2(n10300), .ZN(n10353) );
  AOI22_X1 U13281 ( .A1(n10386), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10382), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10305) );
  AOI22_X1 U13282 ( .A1(n10391), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12622), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10304) );
  AOI22_X1 U13283 ( .A1(n10383), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12469), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10303) );
  AOI22_X1 U13284 ( .A1(n9819), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10381), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10302) );
  NAND4_X1 U13285 ( .A1(n10305), .A2(n10304), .A3(n10303), .A4(n10302), .ZN(
        n10306) );
  NAND2_X1 U13286 ( .A1(n10306), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10313) );
  AOI22_X1 U13287 ( .A1(n10386), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n10381), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10310) );
  AOI22_X1 U13288 ( .A1(n10391), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12622), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10309) );
  AOI22_X1 U13289 ( .A1(n9819), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n10382), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10308) );
  AOI22_X1 U13290 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n10383), .B1(
        n12469), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10307) );
  NAND4_X1 U13291 ( .A1(n10310), .A2(n10309), .A3(n10308), .A4(n10307), .ZN(
        n10311) );
  AND2_X2 U13292 ( .A1(n10353), .A2(n10480), .ZN(n10525) );
  AOI22_X1 U13293 ( .A1(n10383), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12469), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10314) );
  AOI22_X1 U13294 ( .A1(n12622), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n10382), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10317) );
  AOI22_X1 U13295 ( .A1(n9821), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12612), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10315) );
  NAND4_X1 U13296 ( .A1(n10318), .A2(n10317), .A3(n10316), .A4(n10315), .ZN(
        n10325) );
  AOI22_X1 U13297 ( .A1(n10383), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12469), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10319) );
  AND2_X1 U13298 ( .A1(n10319), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10323) );
  AOI22_X1 U13299 ( .A1(n10386), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10391), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10322) );
  AOI22_X1 U13300 ( .A1(n9819), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10381), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10321) );
  AOI22_X1 U13301 ( .A1(n12622), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10382), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10320) );
  NAND4_X1 U13302 ( .A1(n10323), .A2(n10322), .A3(n10321), .A4(n10320), .ZN(
        n10324) );
  AOI22_X1 U13303 ( .A1(n10385), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n10381), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10329) );
  AOI22_X1 U13304 ( .A1(n10383), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12469), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10328) );
  AOI22_X1 U13305 ( .A1(n9820), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n10382), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10327) );
  AOI22_X1 U13306 ( .A1(n10391), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12622), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10326) );
  NAND4_X1 U13307 ( .A1(n10329), .A2(n10328), .A3(n10327), .A4(n10326), .ZN(
        n10331) );
  AOI22_X1 U13308 ( .A1(n10386), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10382), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10334) );
  AOI22_X1 U13309 ( .A1(n10383), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12469), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10333) );
  AOI22_X1 U13310 ( .A1(n9819), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10381), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10332) );
  NAND4_X1 U13311 ( .A1(n10335), .A2(n10334), .A3(n10333), .A4(n10332), .ZN(
        n10336) );
  AOI22_X1 U13312 ( .A1(n9821), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n12612), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10342) );
  AOI22_X1 U13313 ( .A1(n10383), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12469), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10341) );
  AOI22_X1 U13314 ( .A1(n10385), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n10381), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10340) );
  AOI22_X1 U13315 ( .A1(n12622), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n9828), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10339) );
  NAND4_X1 U13316 ( .A1(n10342), .A2(n10341), .A3(n10340), .A4(n10339), .ZN(
        n10343) );
  NAND2_X1 U13317 ( .A1(n10343), .A2(n10330), .ZN(n10350) );
  AOI22_X1 U13318 ( .A1(n9820), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12612), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10347) );
  AOI22_X1 U13319 ( .A1(n12622), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9828), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10346) );
  AOI22_X1 U13320 ( .A1(n10383), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n9818), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10345) );
  AOI22_X1 U13321 ( .A1(n9819), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10381), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10344) );
  NAND4_X1 U13322 ( .A1(n10347), .A2(n10346), .A3(n10345), .A4(n10344), .ZN(
        n10348) );
  NAND2_X1 U13323 ( .A1(n10348), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10349) );
  NOR2_X1 U13324 ( .A1(n10512), .A2(n9776), .ZN(n10380) );
  NAND2_X1 U13325 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n19835) );
  NOR2_X1 U13326 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(P2_STATE_REG_1__SCAN_IN), 
        .ZN(n19717) );
  AOI211_X1 U13327 ( .C1(P2_STATE_REG_1__SCAN_IN), .C2(P2_STATE_REG_2__SCAN_IN), .A(P2_STATE_REG_0__SCAN_IN), .B(n19717), .ZN(n16220) );
  NAND4_X1 U13328 ( .A1(n10537), .A2(n16212), .A3(n19835), .A4(n16220), .ZN(
        n10379) );
  NAND2_X1 U13329 ( .A1(n11013), .A2(n12305), .ZN(n10354) );
  NAND2_X1 U13330 ( .A1(n10497), .A2(n10354), .ZN(n10372) );
  AOI22_X1 U13331 ( .A1(n9821), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10391), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10358) );
  AOI22_X1 U13332 ( .A1(n12622), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10382), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10357) );
  AOI22_X1 U13333 ( .A1(n10383), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12469), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10356) );
  AOI22_X1 U13334 ( .A1(n9819), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10381), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10355) );
  NAND4_X1 U13335 ( .A1(n10358), .A2(n10357), .A3(n10356), .A4(n10355), .ZN(
        n10359) );
  NAND2_X1 U13336 ( .A1(n10359), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10366) );
  AOI22_X1 U13337 ( .A1(n10391), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12622), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10363) );
  AOI22_X1 U13338 ( .A1(n10386), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n10382), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10362) );
  AOI22_X1 U13339 ( .A1(n10383), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n9818), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10361) );
  AOI22_X1 U13340 ( .A1(n10385), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10381), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10360) );
  NAND4_X1 U13341 ( .A1(n10363), .A2(n10362), .A3(n10361), .A4(n10360), .ZN(
        n10364) );
  NAND2_X1 U13342 ( .A1(n10364), .A2(n10330), .ZN(n10365) );
  AND2_X1 U13343 ( .A1(n9776), .A2(n16218), .ZN(n12172) );
  AOI21_X1 U13344 ( .B1(n10372), .B2(n12172), .A(n10538), .ZN(n10378) );
  INV_X1 U13345 ( .A(n10511), .ZN(n10491) );
  NAND2_X1 U13346 ( .A1(n10492), .A2(n10511), .ZN(n10370) );
  NAND2_X1 U13347 ( .A1(n15544), .A2(n10370), .ZN(n10377) );
  NAND2_X1 U13348 ( .A1(n10372), .A2(n10371), .ZN(n10493) );
  OAI21_X1 U13349 ( .B1(n10371), .B2(n9779), .A(n10476), .ZN(n10373) );
  NAND2_X1 U13350 ( .A1(n10373), .A2(n10480), .ZN(n10374) );
  NAND2_X1 U13351 ( .A1(n10374), .A2(n10511), .ZN(n10375) );
  AND2_X1 U13352 ( .A1(n10493), .A2(n10375), .ZN(n10376) );
  NAND4_X1 U13353 ( .A1(n10379), .A2(n10378), .A3(n10377), .A4(n10376), .ZN(
        n15378) );
  AOI21_X1 U13354 ( .B1(n16249), .B2(n10380), .A(n15378), .ZN(n10469) );
  AND2_X2 U13355 ( .A1(n10382), .A2(n10330), .ZN(n15421) );
  AOI22_X1 U13356 ( .A1(n12448), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n15421), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10390) );
  AND2_X1 U13357 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10384) );
  AOI22_X1 U13358 ( .A1(n12450), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12449), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10389) );
  AND2_X1 U13359 ( .A1(n9818), .A2(n10330), .ZN(n10404) );
  AOI22_X1 U13360 ( .A1(n10425), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10404), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10388) );
  AOI22_X1 U13361 ( .A1(n10659), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10653), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10387) );
  NAND4_X1 U13362 ( .A1(n10390), .A2(n10389), .A3(n10388), .A4(n10387), .ZN(
        n10398) );
  AND2_X2 U13363 ( .A1(n12615), .A2(n10330), .ZN(n12451) );
  AOI22_X1 U13365 ( .A1(n12451), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10658), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10396) );
  AOI22_X1 U13366 ( .A1(n10412), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12443), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10395) );
  AOI22_X1 U13367 ( .A1(n10850), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10789), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10394) );
  AOI22_X1 U13368 ( .A1(n10754), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10417), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10393) );
  NAND4_X1 U13369 ( .A1(n10396), .A2(n10395), .A3(n10394), .A4(n10393), .ZN(
        n10397) );
  MUX2_X1 U13370 ( .A(n10444), .B(n10814), .S(n12218), .Z(n11021) );
  INV_X1 U13371 ( .A(n10443), .ZN(n10411) );
  AOI22_X1 U13372 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n10412), .B1(
        n12443), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10403) );
  AOI22_X1 U13373 ( .A1(n10659), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10658), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10402) );
  AOI22_X1 U13374 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n10789), .B1(
        n10754), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10401) );
  AOI22_X1 U13375 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n10850), .B1(
        n15421), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10400) );
  NAND4_X1 U13376 ( .A1(n10403), .A2(n10402), .A3(n10401), .A4(n10400), .ZN(
        n10410) );
  AOI22_X1 U13377 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n10425), .B1(
        n12448), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10408) );
  AOI22_X1 U13378 ( .A1(n12450), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__2__SCAN_IN), .B2(n12449), .ZN(n10407) );
  AOI22_X1 U13379 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n12401), .B1(
        n10404), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10406) );
  AOI22_X1 U13380 ( .A1(n12451), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n10653), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10405) );
  NAND4_X1 U13381 ( .A1(n10408), .A2(n10407), .A3(n10406), .A4(n10405), .ZN(
        n10409) );
  MUX2_X1 U13382 ( .A(n10831), .B(n10449), .S(n10479), .Z(n11016) );
  OAI21_X1 U13383 ( .B1(n11021), .B2(n10411), .A(n11016), .ZN(n10438) );
  AOI22_X1 U13384 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n10412), .B1(
        n12443), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10416) );
  AOI22_X1 U13385 ( .A1(n10659), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10754), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10415) );
  AOI22_X1 U13386 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n10850), .B1(
        n15421), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10414) );
  AOI22_X1 U13387 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n10658), .B1(
        n10789), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10413) );
  NAND4_X1 U13388 ( .A1(n10416), .A2(n10415), .A3(n10414), .A4(n10413), .ZN(
        n10423) );
  AOI22_X1 U13389 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n10425), .B1(
        n12451), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10421) );
  AOI22_X1 U13390 ( .A1(n12450), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__3__SCAN_IN), .B2(n12449), .ZN(n10420) );
  AOI22_X1 U13391 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n12401), .B1(
        n10404), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10419) );
  AOI22_X1 U13392 ( .A1(n12448), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10653), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10418) );
  NAND4_X1 U13393 ( .A1(n10421), .A2(n10420), .A3(n10419), .A4(n10418), .ZN(
        n10422) );
  INV_X1 U13394 ( .A(n10424), .ZN(n10452) );
  MUX2_X1 U13395 ( .A(n10835), .B(n10452), .S(n10479), .Z(n11018) );
  AOI22_X1 U13396 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n10659), .B1(
        n10425), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10429) );
  AOI22_X1 U13397 ( .A1(n12443), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n10658), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10428) );
  AOI22_X1 U13398 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n10789), .B1(
        n10754), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10427) );
  AOI22_X1 U13399 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n10850), .B1(
        n15421), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10426) );
  NAND4_X1 U13400 ( .A1(n10429), .A2(n10428), .A3(n10427), .A4(n10426), .ZN(
        n10435) );
  AOI22_X1 U13401 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n10412), .B1(
        n12448), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10433) );
  AOI22_X1 U13402 ( .A1(n10404), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__4__SCAN_IN), .B2(n12449), .ZN(n10432) );
  AOI22_X1 U13403 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n12401), .B1(
        n10653), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10431) );
  AOI22_X1 U13404 ( .A1(n12451), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n12450), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10430) );
  NAND4_X1 U13405 ( .A1(n10433), .A2(n10432), .A3(n10431), .A4(n10430), .ZN(
        n10434) );
  INV_X1 U13406 ( .A(n10456), .ZN(n10436) );
  MUX2_X1 U13407 ( .A(n10840), .B(n10436), .S(n10479), .Z(n11036) );
  NAND2_X1 U13408 ( .A1(n11018), .A2(n11036), .ZN(n10440) );
  INV_X1 U13409 ( .A(n10440), .ZN(n10437) );
  AOI21_X1 U13410 ( .B1(n10438), .B2(n10437), .A(n10460), .ZN(n19825) );
  INV_X1 U13411 ( .A(n12172), .ZN(n10439) );
  NOR2_X1 U13412 ( .A1(n10512), .A2(n10439), .ZN(n19828) );
  NAND2_X1 U13413 ( .A1(n19825), .A2(n19828), .ZN(n12267) );
  NAND2_X1 U13414 ( .A1(n10440), .A2(n10479), .ZN(n10455) );
  NAND2_X1 U13415 ( .A1(n10535), .A2(n9779), .ZN(n10442) );
  MUX2_X1 U13416 ( .A(n10479), .B(n10442), .S(n10449), .Z(n10451) );
  OAI21_X1 U13417 ( .B1(n10411), .B2(n10444), .A(n12218), .ZN(n10448) );
  INV_X1 U13418 ( .A(n10444), .ZN(n10446) );
  OAI211_X1 U13419 ( .C1(n9779), .C2(n10446), .A(n10476), .B(n10445), .ZN(
        n10447) );
  OAI211_X1 U13420 ( .C1(n10523), .C2(n10449), .A(n10448), .B(n10447), .ZN(
        n10450) );
  NAND2_X1 U13421 ( .A1(n10451), .A2(n10450), .ZN(n10453) );
  NAND2_X1 U13422 ( .A1(n10453), .A2(n10452), .ZN(n10454) );
  NAND2_X1 U13423 ( .A1(n10455), .A2(n10454), .ZN(n10458) );
  AOI21_X1 U13424 ( .B1(n12218), .B2(n10456), .A(n10460), .ZN(n10457) );
  NAND2_X1 U13425 ( .A1(n10458), .A2(n10457), .ZN(n10459) );
  MUX2_X1 U13426 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B(n10459), .S(
        P2_STATE2_REG_0__SCAN_IN), .Z(n10464) );
  NAND2_X1 U13427 ( .A1(n19845), .A2(n10460), .ZN(n10461) );
  NAND2_X1 U13428 ( .A1(n19835), .A2(n16220), .ZN(n10462) );
  NOR2_X1 U13429 ( .A1(n10511), .A2(n10462), .ZN(n10463) );
  NAND2_X1 U13430 ( .A1(n13373), .A2(n10463), .ZN(n10468) );
  INV_X1 U13431 ( .A(n13373), .ZN(n10466) );
  AOI21_X1 U13432 ( .B1(n10464), .B2(n10476), .A(n10371), .ZN(n10465) );
  NAND2_X1 U13433 ( .A1(n10466), .A2(n10465), .ZN(n10467) );
  NAND4_X1 U13434 ( .A1(n10469), .A2(n12267), .A3(n10468), .A4(n10467), .ZN(
        n10470) );
  NAND2_X1 U13435 ( .A1(n10470), .A2(n19840), .ZN(n10475) );
  NOR2_X1 U13436 ( .A1(n10513), .A2(n19844), .ZN(n10472) );
  NOR2_X1 U13437 ( .A1(n10511), .A2(n19844), .ZN(n10471) );
  MUX2_X1 U13438 ( .A(n10472), .B(n10471), .S(n9776), .Z(n10473) );
  NAND2_X1 U13439 ( .A1(n10473), .A2(n13253), .ZN(n10474) );
  NAND2_X1 U13440 ( .A1(n10477), .A2(n10476), .ZN(n10478) );
  AOI21_X2 U13441 ( .B1(n10497), .B2(n13807), .A(n12636), .ZN(n10488) );
  NAND4_X1 U13442 ( .A1(n10481), .A2(n10496), .A3(n10495), .A4(n10488), .ZN(
        n10530) );
  AND3_X1 U13443 ( .A1(n9776), .A2(n10511), .A3(n10808), .ZN(n10483) );
  AND2_X1 U13444 ( .A1(n10531), .A2(n10483), .ZN(n16211) );
  NAND2_X1 U13445 ( .A1(n11125), .A2(n16211), .ZN(n13237) );
  NAND2_X1 U13446 ( .A1(n10497), .A2(n10808), .ZN(n10484) );
  NAND2_X1 U13447 ( .A1(n10485), .A2(n10491), .ZN(n10486) );
  NAND2_X1 U13448 ( .A1(n10487), .A2(n10486), .ZN(n10490) );
  NAND2_X1 U13449 ( .A1(n10490), .A2(n10489), .ZN(n10516) );
  MUX2_X1 U13450 ( .A(n10516), .B(n10491), .S(n16218), .Z(n10501) );
  NAND2_X1 U13451 ( .A1(n10494), .A2(n10493), .ZN(n15370) );
  NAND2_X1 U13452 ( .A1(n15370), .A2(n13807), .ZN(n10520) );
  INV_X1 U13453 ( .A(n10495), .ZN(n13259) );
  OAI21_X1 U13454 ( .B1(n10538), .B2(n10496), .A(n13259), .ZN(n10499) );
  NAND2_X1 U13455 ( .A1(n10497), .A2(n9776), .ZN(n10555) );
  NAND3_X1 U13456 ( .A1(n10555), .A2(n10538), .A3(n10539), .ZN(n10498) );
  NAND3_X1 U13457 ( .A1(n10520), .A2(n10499), .A3(n10498), .ZN(n10500) );
  NAND2_X1 U13458 ( .A1(n15369), .A2(n10539), .ZN(n10502) );
  NAND2_X1 U13459 ( .A1(n11125), .A2(n10502), .ZN(n10504) );
  INV_X1 U13460 ( .A(n10504), .ZN(n13241) );
  INV_X1 U13461 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n11115) );
  NAND3_X1 U13462 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13240) );
  INV_X1 U13463 ( .A(n13240), .ZN(n10503) );
  OR2_X1 U13464 ( .A1(n10504), .A2(n10503), .ZN(n10507) );
  INV_X1 U13465 ( .A(n11125), .ZN(n10505) );
  NAND2_X1 U13466 ( .A1(n15386), .A2(n19796), .ZN(n15543) );
  INV_X1 U13467 ( .A(n15543), .ZN(n19784) );
  NAND2_X1 U13468 ( .A1(n19784), .A2(n19149), .ZN(n13256) );
  NAND2_X1 U13469 ( .A1(n10505), .A2(n9889), .ZN(n15356) );
  INV_X1 U13470 ( .A(n13237), .ZN(n10506) );
  AOI21_X1 U13471 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13238) );
  NAND2_X1 U13472 ( .A1(n10506), .A2(n13238), .ZN(n13242) );
  INV_X1 U13473 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n21127) );
  INV_X1 U13474 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n15349) );
  NAND2_X1 U13475 ( .A1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n15348) );
  NOR3_X1 U13476 ( .A1(n21127), .A2(n15349), .A3(n15348), .ZN(n10957) );
  INV_X1 U13477 ( .A(n10957), .ZN(n10508) );
  NAND2_X1 U13478 ( .A1(n16138), .A2(n10508), .ZN(n10509) );
  AND2_X1 U13479 ( .A1(n21126), .A2(n10509), .ZN(n15336) );
  NAND2_X1 U13480 ( .A1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16187) );
  NAND2_X1 U13481 ( .A1(n16138), .A2(n16187), .ZN(n10510) );
  AND2_X1 U13482 ( .A1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n16143) );
  NAND2_X1 U13483 ( .A1(n16143), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10958) );
  AND2_X1 U13484 ( .A1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16172) );
  NAND2_X1 U13485 ( .A1(n16172), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16139) );
  NOR2_X1 U13486 ( .A1(n10958), .A2(n16139), .ZN(n12246) );
  AND2_X1 U13487 ( .A1(n21126), .A2(n15357), .ZN(n15304) );
  AOI21_X1 U13488 ( .B1(n16136), .B2(n12246), .A(n15304), .ZN(n15301) );
  NAND2_X1 U13489 ( .A1(n10512), .A2(n10246), .ZN(n10514) );
  NAND2_X1 U13490 ( .A1(n10514), .A2(n10513), .ZN(n10952) );
  INV_X1 U13491 ( .A(n10952), .ZN(n10515) );
  NAND2_X1 U13492 ( .A1(n10515), .A2(n19845), .ZN(n10518) );
  NAND2_X1 U13493 ( .A1(n10516), .A2(n19841), .ZN(n10517) );
  NAND2_X1 U13494 ( .A1(n10520), .A2(n10519), .ZN(n10556) );
  AOI21_X2 U13495 ( .B1(n10556), .B2(n19845), .A(n10521), .ZN(n10522) );
  NAND2_X2 U13496 ( .A1(n10554), .A2(n10522), .ZN(n10575) );
  NAND2_X1 U13497 ( .A1(n10575), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10529) );
  INV_X1 U13498 ( .A(n10523), .ZN(n10524) );
  NAND2_X1 U13499 ( .A1(n12633), .A2(n10526), .ZN(n10527) );
  NOR2_X1 U13500 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n10576) );
  AOI22_X1 U13501 ( .A1(n15416), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n10576), 
        .B2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n10528) );
  INV_X1 U13502 ( .A(n10530), .ZN(n10531) );
  NAND2_X1 U13503 ( .A1(n10531), .A2(n10538), .ZN(n10546) );
  OAI211_X1 U13504 ( .C1(n9779), .C2(n10953), .A(n10546), .B(n10532), .ZN(
        n10533) );
  INV_X1 U13505 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n10543) );
  NAND2_X1 U13506 ( .A1(n10540), .A2(P2_EBX_REG_1__SCAN_IN), .ZN(n10542) );
  NAND2_X1 U13507 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n10541) );
  OAI211_X1 U13508 ( .C1(n9775), .C2(n10543), .A(n10542), .B(n10541), .ZN(
        n10544) );
  INV_X1 U13509 ( .A(n10576), .ZN(n10551) );
  OAI22_X1 U13510 ( .A1(n15397), .A2(n19836), .B1(n10551), .B2(n19821), .ZN(
        n10547) );
  INV_X1 U13511 ( .A(n10547), .ZN(n10548) );
  NAND2_X1 U13512 ( .A1(n10549), .A2(n10548), .ZN(n10597) );
  NAND2_X1 U13513 ( .A1(n12209), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n10553) );
  NAND2_X1 U13514 ( .A1(n10540), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n10552) );
  NAND2_X1 U13515 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n10550) );
  NAND2_X1 U13516 ( .A1(n9826), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10558) );
  OAI211_X1 U13517 ( .C1(n10556), .C2(n10476), .A(P2_STATE2_REG_0__SCAN_IN), 
        .B(n10555), .ZN(n10557) );
  NAND2_X1 U13518 ( .A1(n10597), .A2(n10595), .ZN(n10593) );
  NAND2_X1 U13519 ( .A1(n10592), .A2(n10593), .ZN(n10591) );
  INV_X1 U13520 ( .A(n10559), .ZN(n10561) );
  NAND2_X1 U13521 ( .A1(n10561), .A2(n10560), .ZN(n10562) );
  NAND2_X1 U13522 ( .A1(n10575), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10564) );
  AOI21_X1 U13523 ( .B1(n19836), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n10563) );
  NAND2_X1 U13524 ( .A1(n10564), .A2(n10563), .ZN(n10572) );
  INV_X1 U13525 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13244) );
  NAND2_X1 U13526 ( .A1(n10579), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10570) );
  NAND2_X1 U13527 ( .A1(n10540), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n10569) );
  INV_X1 U13528 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n10566) );
  INV_X1 U13529 ( .A(n10567), .ZN(n10568) );
  NAND2_X1 U13530 ( .A1(n10570), .A2(n10233), .ZN(n10571) );
  NAND2_X1 U13531 ( .A1(n10572), .A2(n10571), .ZN(n10573) );
  NAND2_X1 U13532 ( .A1(n10575), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10578) );
  NAND2_X1 U13533 ( .A1(n10576), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10577) );
  NAND2_X1 U13534 ( .A1(n10578), .A2(n10577), .ZN(n10584) );
  INV_X4 U13535 ( .A(n9774), .ZN(n12209) );
  AOI22_X1 U13536 ( .A1(n12209), .A2(P2_REIP_REG_3__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10581) );
  CLKBUF_X3 U13537 ( .A(n10540), .Z(n10992) );
  NAND2_X1 U13538 ( .A1(n10992), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n10580) );
  NAND2_X1 U13539 ( .A1(n10584), .A2(n10583), .ZN(n10585) );
  INV_X1 U13540 ( .A(n12304), .ZN(n10600) );
  INV_X1 U13541 ( .A(n10586), .ZN(n10589) );
  INV_X1 U13542 ( .A(n10587), .ZN(n10588) );
  NAND2_X1 U13543 ( .A1(n10589), .A2(n10588), .ZN(n10590) );
  INV_X1 U13544 ( .A(n10595), .ZN(n10596) );
  XNOR2_X2 U13545 ( .A(n10597), .B(n10596), .ZN(n12319) );
  NAND2_X1 U13546 ( .A1(n14672), .A2(n15359), .ZN(n10607) );
  INV_X1 U13547 ( .A(n19265), .ZN(n19267) );
  INV_X1 U13548 ( .A(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12517) );
  NAND2_X1 U13549 ( .A1(n15395), .A2(n15359), .ZN(n10606) );
  NAND2_X1 U13550 ( .A1(n19317), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n10598) );
  OAI21_X1 U13551 ( .B1(n19267), .B2(n12517), .A(n10598), .ZN(n10604) );
  NAND2_X1 U13552 ( .A1(n12319), .A2(n9810), .ZN(n10618) );
  INV_X1 U13553 ( .A(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12519) );
  INV_X1 U13554 ( .A(n9810), .ZN(n10601) );
  NAND2_X1 U13555 ( .A1(n12319), .A2(n10601), .ZN(n10616) );
  INV_X1 U13556 ( .A(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10602) );
  OAI22_X1 U13557 ( .A1(n10695), .A2(n12519), .B1(n10687), .B2(n10602), .ZN(
        n10603) );
  INV_X1 U13558 ( .A(n10731), .ZN(n10690) );
  INV_X1 U13559 ( .A(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13811) );
  INV_X1 U13560 ( .A(n10732), .ZN(n10686) );
  INV_X1 U13561 ( .A(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12516) );
  OAI22_X1 U13562 ( .A1(n10690), .A2(n13811), .B1(n10686), .B2(n12516), .ZN(
        n10609) );
  INV_X1 U13563 ( .A(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12518) );
  INV_X1 U13564 ( .A(n10733), .ZN(n10697) );
  INV_X1 U13565 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12312) );
  OAI22_X1 U13566 ( .A1(n12518), .A2(n10697), .B1(n10698), .B2(n12312), .ZN(
        n10608) );
  NOR2_X1 U13567 ( .A1(n10609), .A2(n10608), .ZN(n10630) );
  INV_X1 U13568 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12526) );
  NAND2_X1 U13569 ( .A1(n12304), .A2(n15359), .ZN(n10622) );
  INV_X1 U13570 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10611) );
  OAI22_X1 U13571 ( .A1(n12526), .A2(n10701), .B1(n10702), .B2(n10611), .ZN(
        n10621) );
  INV_X1 U13572 ( .A(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12528) );
  INV_X1 U13573 ( .A(n10618), .ZN(n10612) );
  AND2_X1 U13574 ( .A1(n9829), .A2(n10612), .ZN(n10613) );
  INV_X1 U13575 ( .A(n10616), .ZN(n10614) );
  NOR2_X1 U13576 ( .A1(n9829), .A2(n10616), .ZN(n10617) );
  NOR2_X1 U13577 ( .A1(n9829), .A2(n10618), .ZN(n10619) );
  INV_X1 U13578 ( .A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12527) );
  NOR2_X1 U13579 ( .A1(n10621), .A2(n10620), .ZN(n10629) );
  INV_X1 U13580 ( .A(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12525) );
  INV_X1 U13581 ( .A(n10622), .ZN(n10623) );
  NAND2_X1 U13582 ( .A1(n10623), .A2(n10599), .ZN(n10624) );
  NOR2_X2 U13583 ( .A1(n10624), .A2(n14672), .ZN(n10639) );
  INV_X1 U13584 ( .A(n10639), .ZN(n10747) );
  INV_X1 U13585 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10626) );
  OAI22_X1 U13586 ( .A1(n12525), .A2(n10747), .B1(n10746), .B2(n10626), .ZN(
        n10627) );
  INV_X1 U13587 ( .A(n10627), .ZN(n10628) );
  NAND3_X1 U13588 ( .A1(n10630), .A2(n10629), .A3(n10628), .ZN(n10633) );
  INV_X1 U13589 ( .A(n10835), .ZN(n10631) );
  NAND2_X1 U13590 ( .A1(n10631), .A2(n9776), .ZN(n10632) );
  INV_X1 U13591 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10637) );
  AOI21_X1 U13592 ( .B1(n19418), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A(n9776), .ZN(n10636) );
  INV_X1 U13593 ( .A(n19473), .ZN(n10634) );
  OAI211_X1 U13594 ( .C1(n10687), .C2(n10637), .A(n10636), .B(n10635), .ZN(
        n10638) );
  AOI21_X1 U13595 ( .B1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B2(n19389), .A(
        n10638), .ZN(n10652) );
  AOI22_X1 U13596 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n10732), .B1(
        n19317), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10641) );
  NAND2_X1 U13597 ( .A1(n10639), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n10640) );
  AND2_X1 U13598 ( .A1(n10641), .A2(n10640), .ZN(n10651) );
  INV_X1 U13599 ( .A(n10701), .ZN(n10738) );
  NAND2_X1 U13600 ( .A1(n19153), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n10644) );
  AOI22_X1 U13601 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19638), .B1(
        n19539), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10643) );
  NAND2_X1 U13602 ( .A1(n19605), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n10642) );
  NAND3_X1 U13603 ( .A1(n10644), .A2(n10643), .A3(n10642), .ZN(n10645) );
  NAND2_X1 U13604 ( .A1(n19265), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n10649) );
  NAND2_X1 U13605 ( .A1(n19355), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n10648) );
  NAND2_X1 U13606 ( .A1(n10733), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n10647) );
  NAND2_X1 U13607 ( .A1(n10731), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n10646) );
  NAND4_X1 U13608 ( .A1(n10652), .A2(n10651), .A3(n10650), .A4(n10239), .ZN(
        n10668) );
  AOI22_X1 U13609 ( .A1(n12448), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12401), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10657) );
  AOI22_X1 U13610 ( .A1(n12443), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n10789), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10656) );
  AOI22_X1 U13611 ( .A1(n10404), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12449), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10655) );
  AOI22_X1 U13612 ( .A1(n15421), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n10653), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10654) );
  NAND4_X1 U13613 ( .A1(n10657), .A2(n10656), .A3(n10655), .A4(n10654), .ZN(
        n10665) );
  AOI22_X1 U13614 ( .A1(n12451), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n10658), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10663) );
  AOI22_X1 U13615 ( .A1(n10412), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n10659), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10662) );
  AOI22_X1 U13616 ( .A1(n10425), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12450), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10661) );
  AOI22_X1 U13617 ( .A1(n10850), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10754), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10660) );
  NAND4_X1 U13618 ( .A1(n10663), .A2(n10662), .A3(n10661), .A4(n10660), .ZN(
        n10664) );
  NOR2_X1 U13619 ( .A1(n10814), .A2(n11015), .ZN(n10666) );
  NAND2_X1 U13620 ( .A1(n9776), .A2(n10666), .ZN(n10675) );
  NAND2_X1 U13621 ( .A1(n10675), .A2(n10831), .ZN(n10667) );
  NAND2_X1 U13622 ( .A1(n10670), .A2(n9807), .ZN(n10671) );
  INV_X1 U13623 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13263) );
  NOR2_X1 U13624 ( .A1(n10124), .A2(n13263), .ZN(n13262) );
  INV_X1 U13625 ( .A(n11015), .ZN(n10672) );
  NAND2_X1 U13626 ( .A1(n13262), .A2(n10672), .ZN(n10674) );
  NOR2_X1 U13627 ( .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n10124), .ZN(
        n10673) );
  XOR2_X1 U13628 ( .A(n11015), .B(n10673), .Z(n13333) );
  NAND2_X1 U13629 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n13333), .ZN(
        n13332) );
  NAND2_X1 U13630 ( .A1(n10674), .A2(n13332), .ZN(n10676) );
  XNOR2_X1 U13631 ( .A(n13244), .B(n10676), .ZN(n13248) );
  XNOR2_X1 U13632 ( .A(n10675), .B(n10831), .ZN(n13247) );
  NAND2_X1 U13633 ( .A1(n13248), .A2(n13247), .ZN(n10678) );
  NAND2_X1 U13634 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n10676), .ZN(
        n10677) );
  NAND2_X1 U13635 ( .A1(n10678), .A2(n10677), .ZN(n10679) );
  XNOR2_X1 U13636 ( .A(n10679), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13790) );
  NAND2_X1 U13637 ( .A1(n10679), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10680) );
  INV_X1 U13638 ( .A(n10840), .ZN(n10685) );
  INV_X1 U13639 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n13850) );
  NAND2_X1 U13640 ( .A1(n13851), .A2(n13850), .ZN(n13849) );
  INV_X1 U13641 ( .A(n10681), .ZN(n10683) );
  NAND2_X1 U13642 ( .A1(n10683), .A2(n10682), .ZN(n10684) );
  INV_X1 U13643 ( .A(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12572) );
  INV_X1 U13644 ( .A(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12571) );
  OAI22_X1 U13645 ( .A1(n19267), .A2(n12572), .B1(n10686), .B2(n12571), .ZN(
        n10692) );
  INV_X1 U13646 ( .A(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10689) );
  INV_X1 U13647 ( .A(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10688) );
  OAI22_X1 U13648 ( .A1(n10690), .A2(n10689), .B1(n10687), .B2(n10688), .ZN(
        n10691) );
  NOR2_X1 U13649 ( .A1(n10692), .A2(n10691), .ZN(n10714) );
  INV_X1 U13650 ( .A(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12580) );
  INV_X1 U13651 ( .A(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10693) );
  OAI22_X1 U13652 ( .A1(n12580), .A2(n10747), .B1(n10746), .B2(n10693), .ZN(
        n10694) );
  INV_X1 U13653 ( .A(n10694), .ZN(n10713) );
  INV_X1 U13654 ( .A(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12574) );
  NAND2_X1 U13655 ( .A1(n19317), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n10696) );
  OAI21_X1 U13656 ( .B1(n10695), .B2(n12574), .A(n10696), .ZN(n10700) );
  INV_X1 U13657 ( .A(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12573) );
  INV_X1 U13658 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13571) );
  OAI22_X1 U13659 ( .A1(n12573), .A2(n10697), .B1(n10698), .B2(n13571), .ZN(
        n10699) );
  NOR2_X1 U13660 ( .A1(n10700), .A2(n10699), .ZN(n10712) );
  INV_X1 U13661 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12582) );
  INV_X1 U13662 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10703) );
  OAI22_X1 U13663 ( .A1(n12582), .A2(n10701), .B1(n10702), .B2(n10703), .ZN(
        n10710) );
  INV_X1 U13664 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12584) );
  INV_X1 U13665 ( .A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10704) );
  OAI22_X1 U13666 ( .A1(n12584), .A2(n19473), .B1(n10705), .B2(n10704), .ZN(
        n10708) );
  INV_X1 U13667 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12585) );
  INV_X1 U13668 ( .A(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10706) );
  OAI22_X1 U13669 ( .A1(n12585), .A2(n19645), .B1(n19415), .B2(n10706), .ZN(
        n10707) );
  OR2_X1 U13670 ( .A1(n10708), .A2(n10707), .ZN(n10709) );
  NOR2_X1 U13671 ( .A1(n10710), .A2(n10709), .ZN(n10711) );
  NAND4_X1 U13672 ( .A1(n10714), .A2(n10713), .A3(n10712), .A4(n10711), .ZN(
        n10726) );
  AOI22_X1 U13673 ( .A1(n10412), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12443), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10718) );
  AOI22_X1 U13674 ( .A1(n10659), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10754), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10717) );
  AOI22_X1 U13675 ( .A1(n10850), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n15421), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10716) );
  AOI22_X1 U13676 ( .A1(n10658), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10789), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10715) );
  NAND4_X1 U13677 ( .A1(n10718), .A2(n10717), .A3(n10716), .A4(n10715), .ZN(
        n10724) );
  AOI22_X1 U13678 ( .A1(n10425), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12451), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10722) );
  AOI22_X1 U13679 ( .A1(n12450), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12449), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10721) );
  AOI22_X1 U13680 ( .A1(n12401), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10404), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10720) );
  AOI22_X1 U13681 ( .A1(n12448), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10653), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10719) );
  NAND4_X1 U13682 ( .A1(n10722), .A2(n10721), .A3(n10720), .A4(n10719), .ZN(
        n10723) );
  NAND2_X1 U13683 ( .A1(n11043), .A2(n9776), .ZN(n10725) );
  XNOR2_X2 U13684 ( .A(n10730), .B(n10728), .ZN(n11040) );
  INV_X1 U13685 ( .A(n11040), .ZN(n10727) );
  INV_X1 U13686 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n11048) );
  NOR2_X2 U13687 ( .A1(n13884), .A2(n13881), .ZN(n10771) );
  NAND2_X1 U13688 ( .A1(n10731), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n10737) );
  NAND2_X1 U13689 ( .A1(n10732), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n10736) );
  INV_X1 U13690 ( .A(n10687), .ZN(n19187) );
  NAND2_X1 U13691 ( .A1(n19187), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n10735) );
  NAND2_X1 U13692 ( .A1(n10733), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n10734) );
  NAND4_X1 U13693 ( .A1(n10737), .A2(n10736), .A3(n10735), .A4(n10734), .ZN(
        n10744) );
  AOI22_X1 U13694 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19638), .B1(
        n19539), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10742) );
  AOI22_X1 U13695 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n10634), .B1(
        n19418), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10741) );
  NAND2_X1 U13696 ( .A1(n10738), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n10740) );
  NAND2_X1 U13697 ( .A1(n19605), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n10739) );
  NAND4_X1 U13698 ( .A1(n10742), .A2(n10741), .A3(n10740), .A4(n10739), .ZN(
        n10743) );
  NOR2_X1 U13699 ( .A1(n10744), .A2(n10743), .ZN(n10753) );
  AOI22_X1 U13700 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19265), .B1(
        n19153), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10752) );
  INV_X1 U13701 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10748) );
  INV_X1 U13702 ( .A(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10745) );
  OAI22_X1 U13703 ( .A1(n10748), .A2(n10747), .B1(n10746), .B2(n10745), .ZN(
        n10749) );
  INV_X1 U13704 ( .A(n10749), .ZN(n10751) );
  AOI22_X1 U13705 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19355), .B1(
        n19317), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10750) );
  NAND4_X1 U13706 ( .A1(n10753), .A2(n10752), .A3(n10751), .A4(n10750), .ZN(
        n10766) );
  AOI22_X1 U13707 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n10412), .B1(
        n12443), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10758) );
  AOI22_X1 U13708 ( .A1(n10659), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10754), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10757) );
  AOI22_X1 U13709 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n10850), .B1(
        n15421), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10756) );
  AOI22_X1 U13710 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n10658), .B1(
        n10789), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10755) );
  NAND4_X1 U13711 ( .A1(n10758), .A2(n10757), .A3(n10756), .A4(n10755), .ZN(
        n10764) );
  AOI22_X1 U13712 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n10425), .B1(
        n12451), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10762) );
  AOI22_X1 U13713 ( .A1(n12450), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__6__SCAN_IN), .B2(n12449), .ZN(n10761) );
  AOI22_X1 U13714 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n12401), .B1(
        n10404), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10760) );
  AOI22_X1 U13715 ( .A1(n12448), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10653), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10759) );
  NAND4_X1 U13716 ( .A1(n10762), .A2(n10761), .A3(n10760), .A4(n10759), .ZN(
        n10763) );
  NAND2_X1 U13717 ( .A1(n11052), .A2(n9776), .ZN(n10765) );
  INV_X1 U13718 ( .A(n11056), .ZN(n10774) );
  NAND2_X1 U13719 ( .A1(n11040), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10772) );
  INV_X1 U13720 ( .A(n10772), .ZN(n13882) );
  INV_X1 U13721 ( .A(n10768), .ZN(n10769) );
  NAND2_X1 U13722 ( .A1(n13882), .A2(n10769), .ZN(n10770) );
  INV_X1 U13723 ( .A(n10771), .ZN(n10773) );
  NAND2_X1 U13724 ( .A1(n10773), .A2(n10772), .ZN(n10775) );
  NAND2_X1 U13725 ( .A1(n12443), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n10780) );
  NAND2_X1 U13726 ( .A1(n10412), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n10779) );
  NAND2_X1 U13727 ( .A1(n10659), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n10778) );
  NAND2_X1 U13728 ( .A1(n10754), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n10777) );
  NAND2_X1 U13729 ( .A1(n12448), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n10784) );
  NAND2_X1 U13730 ( .A1(n10425), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n10783) );
  NAND2_X1 U13731 ( .A1(n12451), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n10782) );
  NAND2_X1 U13732 ( .A1(n10653), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n10781) );
  NAND2_X1 U13733 ( .A1(n12450), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n10788) );
  NAND2_X1 U13734 ( .A1(n12401), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n10787) );
  NAND2_X1 U13735 ( .A1(n10404), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n10786) );
  NAND2_X1 U13736 ( .A1(n12449), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n10785) );
  NAND2_X1 U13737 ( .A1(n10850), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n10793) );
  NAND2_X1 U13738 ( .A1(n15421), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n10792) );
  NAND2_X1 U13739 ( .A1(n10658), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n10791) );
  NAND2_X1 U13740 ( .A1(n10789), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n10790) );
  XNOR2_X1 U13741 ( .A(n10801), .B(n10849), .ZN(n10798) );
  XNOR2_X1 U13742 ( .A(n10798), .B(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15104) );
  INV_X1 U13743 ( .A(n10798), .ZN(n10799) );
  NAND2_X1 U13744 ( .A1(n10799), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10800) );
  XNOR2_X1 U13745 ( .A(n10802), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16108) );
  INV_X1 U13746 ( .A(n10802), .ZN(n10803) );
  NAND2_X1 U13747 ( .A1(n10803), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10804) );
  INV_X1 U13748 ( .A(n16172), .ZN(n10805) );
  NOR2_X2 U13749 ( .A1(n16081), .A2(n10958), .ZN(n16070) );
  INV_X1 U13750 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15290) );
  OAI21_X1 U13751 ( .B1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n15357), .A(
        n15291), .ZN(n11011) );
  NOR2_X1 U13752 ( .A1(n10480), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n10807) );
  INV_X2 U13753 ( .A(n12165), .ZN(n12151) );
  AOI22_X1 U13754 ( .A1(n12151), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n10820), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n10811) );
  NAND2_X1 U13755 ( .A1(n12156), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n10810) );
  NAND2_X1 U13756 ( .A1(n10811), .A2(n10810), .ZN(n13232) );
  NOR2_X1 U13757 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19796), .ZN(
        n19818) );
  INV_X1 U13758 ( .A(n10497), .ZN(n10812) );
  NAND2_X1 U13759 ( .A1(n10812), .A2(n9830), .ZN(n10830) );
  OAI21_X1 U13760 ( .B1(n10822), .B2(n19818), .A(n10830), .ZN(n10813) );
  INV_X1 U13761 ( .A(n10813), .ZN(n10815) );
  INV_X1 U13762 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n10817) );
  NAND2_X1 U13763 ( .A1(n9779), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10816) );
  OAI211_X1 U13764 ( .C1(n10480), .C2(n10817), .A(n10816), .B(n19796), .ZN(
        n10818) );
  INV_X1 U13765 ( .A(n10818), .ZN(n10819) );
  INV_X1 U13766 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n15389) );
  AOI22_X1 U13767 ( .A1(n10807), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n9831), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n10821) );
  NAND2_X1 U13768 ( .A1(n10821), .A2(n9858), .ZN(n10825) );
  OR2_X1 U13769 ( .A1(n11015), .A2(n10951), .ZN(n10824) );
  AOI22_X1 U13770 ( .A1(n10497), .A2(n10822), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n10823) );
  NAND2_X1 U13771 ( .A1(n10824), .A2(n10823), .ZN(n13381) );
  NOR2_X1 U13772 ( .A1(n13382), .A2(n13381), .ZN(n10828) );
  NOR2_X1 U13773 ( .A1(n10826), .A2(n10825), .ZN(n10827) );
  NOR2_X2 U13774 ( .A1(n10828), .A2(n10827), .ZN(n10833) );
  NAND2_X1 U13775 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n10829) );
  OAI211_X1 U13776 ( .C1(n10831), .C2(n10951), .A(n10830), .B(n10829), .ZN(
        n10832) );
  XNOR2_X1 U13777 ( .A(n10833), .B(n10832), .ZN(n13233) );
  NOR2_X1 U13778 ( .A1(n13232), .A2(n13233), .ZN(n13234) );
  NOR2_X1 U13779 ( .A1(n10833), .A2(n10832), .ZN(n10834) );
  NOR2_X2 U13780 ( .A1(n13234), .A2(n10834), .ZN(n14638) );
  NAND2_X1 U13781 ( .A1(n12156), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n10839) );
  NAND2_X1 U13782 ( .A1(n10125), .A2(n10835), .ZN(n10838) );
  AOI22_X1 U13783 ( .A1(n10820), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n10837) );
  NAND2_X1 U13784 ( .A1(n12151), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n10836) );
  NAND4_X1 U13785 ( .A1(n10839), .A2(n10838), .A3(n10837), .A4(n10836), .ZN(
        n14637) );
  NAND2_X1 U13786 ( .A1(n14638), .A2(n14637), .ZN(n13860) );
  AOI22_X1 U13787 ( .A1(n12151), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n10820), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n10843) );
  NAND2_X1 U13788 ( .A1(n12156), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n10842) );
  NAND2_X1 U13789 ( .A1(n10125), .A2(n10840), .ZN(n10841) );
  AOI22_X1 U13790 ( .A1(n12156), .A2(P2_REIP_REG_5__SCAN_IN), .B1(n10125), 
        .B2(n10844), .ZN(n10846) );
  AOI22_X1 U13791 ( .A1(n12151), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n10820), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n10845) );
  NAND2_X1 U13792 ( .A1(n10846), .A2(n10845), .ZN(n13886) );
  NAND2_X1 U13793 ( .A1(n13861), .A2(n13886), .ZN(n13885) );
  INV_X1 U13794 ( .A(n13885), .ZN(n10847) );
  AOI21_X1 U13795 ( .B1(n10125), .B2(n10848), .A(n10847), .ZN(n13405) );
  AOI222_X1 U13796 ( .A1(P2_REIP_REG_6__SCAN_IN), .A2(n12156), .B1(n10820), 
        .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .C1(P2_EAX_REG_6__SCAN_IN), 
        .C2(n12151), .ZN(n13404) );
  OAI22_X2 U13797 ( .A1(n13405), .A2(n13404), .B1(n10849), .B2(n10951), .ZN(
        n13419) );
  INV_X1 U13798 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n15340) );
  INV_X1 U13799 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n19116) );
  INV_X1 U13800 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n19733) );
  OAI222_X1 U13801 ( .A1(n15340), .A2(n12166), .B1(n12165), .B2(n19116), .C1(
        n12167), .C2(n19733), .ZN(n13418) );
  AOI22_X1 U13802 ( .A1(n12151), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n10820), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n10863) );
  NAND2_X1 U13803 ( .A1(n12156), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n10862) );
  AOI22_X1 U13804 ( .A1(n10412), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10425), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10854) );
  AOI22_X1 U13805 ( .A1(n10659), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n15421), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10853) );
  AOI22_X1 U13806 ( .A1(n10658), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10789), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10852) );
  AOI22_X1 U13807 ( .A1(n10850), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10754), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10851) );
  NAND4_X1 U13808 ( .A1(n10854), .A2(n10853), .A3(n10852), .A4(n10851), .ZN(
        n10860) );
  AOI22_X1 U13809 ( .A1(n12443), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12448), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10858) );
  AOI22_X1 U13810 ( .A1(n12450), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12449), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10857) );
  AOI22_X1 U13811 ( .A1(n12401), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10404), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10856) );
  AOI22_X1 U13812 ( .A1(n12451), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10653), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10855) );
  NAND4_X1 U13813 ( .A1(n10858), .A2(n10857), .A3(n10856), .A4(n10855), .ZN(
        n10859) );
  NAND2_X1 U13814 ( .A1(n10125), .A2(n19028), .ZN(n10861) );
  AOI22_X1 U13815 ( .A1(n10412), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12443), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10867) );
  AOI22_X1 U13816 ( .A1(n10659), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n10754), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10866) );
  AOI22_X1 U13817 ( .A1(n10850), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n15421), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10865) );
  AOI22_X1 U13818 ( .A1(n10658), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n10789), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10864) );
  NAND4_X1 U13819 ( .A1(n10867), .A2(n10866), .A3(n10865), .A4(n10864), .ZN(
        n10873) );
  AOI22_X1 U13820 ( .A1(n10425), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12451), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10871) );
  AOI22_X1 U13821 ( .A1(n12450), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12449), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10870) );
  AOI22_X1 U13822 ( .A1(n12401), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10404), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10869) );
  AOI22_X1 U13823 ( .A1(n12448), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10653), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10868) );
  NAND4_X1 U13824 ( .A1(n10871), .A2(n10870), .A3(n10869), .A4(n10868), .ZN(
        n10872) );
  AOI22_X1 U13825 ( .A1(n12151), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n10820), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n10875) );
  NAND2_X1 U13826 ( .A1(n12156), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n10874) );
  OAI211_X1 U13827 ( .C1(n12340), .C2(n10951), .A(n10875), .B(n10874), .ZN(
        n13536) );
  AOI22_X1 U13828 ( .A1(n12151), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n10820), 
        .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n10888) );
  NAND2_X1 U13829 ( .A1(n12156), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n10887) );
  AOI22_X1 U13830 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n10412), .B1(
        n12443), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10879) );
  AOI22_X1 U13831 ( .A1(n10659), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10754), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10878) );
  AOI22_X1 U13832 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n10658), .B1(
        n15421), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10877) );
  AOI22_X1 U13833 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n10789), .B1(
        n10850), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10876) );
  NAND4_X1 U13834 ( .A1(n10879), .A2(n10878), .A3(n10877), .A4(n10876), .ZN(
        n10885) );
  AOI22_X1 U13835 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n10425), .B1(
        n12448), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10883) );
  AOI22_X1 U13836 ( .A1(n12450), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__2__SCAN_IN), .B2(n12449), .ZN(n10882) );
  AOI22_X1 U13837 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n12401), .B1(
        n10404), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10881) );
  AOI22_X1 U13838 ( .A1(n12451), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n10653), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10880) );
  NAND4_X1 U13839 ( .A1(n10883), .A2(n10882), .A3(n10881), .A4(n10880), .ZN(
        n10884) );
  NAND2_X1 U13840 ( .A1(n10125), .A2(n12341), .ZN(n10886) );
  AOI22_X1 U13841 ( .A1(n12156), .A2(P2_REIP_REG_11__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n10820), .ZN(n10900) );
  AOI22_X1 U13842 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n10412), .B1(
        n12443), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10892) );
  AOI22_X1 U13843 ( .A1(n10659), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10754), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10891) );
  AOI22_X1 U13844 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n15421), .B1(
        n10850), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10890) );
  AOI22_X1 U13845 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n10658), .B1(
        n10789), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10889) );
  NAND4_X1 U13846 ( .A1(n10892), .A2(n10891), .A3(n10890), .A4(n10889), .ZN(
        n10898) );
  AOI22_X1 U13847 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n10425), .B1(
        n12451), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10896) );
  AOI22_X1 U13848 ( .A1(n12450), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__3__SCAN_IN), .B2(n12449), .ZN(n10895) );
  AOI22_X1 U13849 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n12401), .B1(
        n10404), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10894) );
  AOI22_X1 U13850 ( .A1(n12448), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10653), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10893) );
  NAND4_X1 U13851 ( .A1(n10896), .A2(n10895), .A3(n10894), .A4(n10893), .ZN(
        n10897) );
  AOI22_X1 U13852 ( .A1(n10125), .A2(n19016), .B1(n12151), .B2(
        P2_EAX_REG_11__SCAN_IN), .ZN(n10899) );
  NAND2_X1 U13853 ( .A1(n10900), .A2(n10899), .ZN(n13617) );
  NAND2_X1 U13854 ( .A1(n13618), .A2(n13617), .ZN(n13616) );
  AOI22_X1 U13855 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n10659), .B1(
        n10425), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10904) );
  AOI22_X1 U13856 ( .A1(n12443), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n15421), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10903) );
  AOI22_X1 U13857 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n10754), .B1(
        n10658), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10902) );
  AOI22_X1 U13858 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n10789), .B1(
        n10850), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10901) );
  NAND4_X1 U13859 ( .A1(n10904), .A2(n10903), .A3(n10902), .A4(n10901), .ZN(
        n10910) );
  AOI22_X1 U13860 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n10412), .B1(
        n12448), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10908) );
  AOI22_X1 U13861 ( .A1(n12401), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__4__SCAN_IN), .B2(n12449), .ZN(n10907) );
  AOI22_X1 U13862 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n12450), .B1(
        n10653), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10906) );
  AOI22_X1 U13863 ( .A1(n12451), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n10404), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10905) );
  NAND4_X1 U13864 ( .A1(n10908), .A2(n10907), .A3(n10906), .A4(n10905), .ZN(
        n10909) );
  INV_X1 U13865 ( .A(n19015), .ZN(n10912) );
  AOI22_X1 U13866 ( .A1(n12151), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n10820), 
        .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n10911) );
  OAI21_X1 U13867 ( .B1(n10912), .B2(n10951), .A(n10911), .ZN(n10913) );
  AOI21_X1 U13868 ( .B1(P2_REIP_REG_12__SCAN_IN), .B2(n12156), .A(n10913), 
        .ZN(n14589) );
  AOI22_X1 U13869 ( .A1(n10412), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12443), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10917) );
  AOI22_X1 U13870 ( .A1(n10659), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10754), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10916) );
  AOI22_X1 U13871 ( .A1(n10850), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n15421), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10915) );
  AOI22_X1 U13872 ( .A1(n10658), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10789), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10914) );
  NAND4_X1 U13873 ( .A1(n10917), .A2(n10916), .A3(n10915), .A4(n10914), .ZN(
        n10923) );
  AOI22_X1 U13874 ( .A1(n10425), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12451), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10921) );
  AOI22_X1 U13875 ( .A1(n12450), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12449), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10920) );
  AOI22_X1 U13876 ( .A1(n12401), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10404), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10919) );
  AOI22_X1 U13877 ( .A1(n12448), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10653), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10918) );
  NAND4_X1 U13878 ( .A1(n10921), .A2(n10920), .A3(n10919), .A4(n10918), .ZN(
        n10922) );
  INV_X1 U13879 ( .A(n13762), .ZN(n10926) );
  AOI22_X1 U13880 ( .A1(n12151), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n10820), 
        .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n10925) );
  NAND2_X1 U13881 ( .A1(n12156), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n10924) );
  OAI211_X1 U13882 ( .C1(n10926), .C2(n10951), .A(n10925), .B(n10924), .ZN(
        n13725) );
  AND2_X2 U13883 ( .A1(n13726), .A2(n13725), .ZN(n13724) );
  AOI22_X1 U13884 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n10412), .B1(
        n12443), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10930) );
  AOI22_X1 U13885 ( .A1(n10659), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10850), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10929) );
  AOI22_X1 U13886 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n10754), .B1(
        n10658), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10928) );
  AOI22_X1 U13887 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n15421), .B1(
        n10789), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10927) );
  NAND4_X1 U13888 ( .A1(n10930), .A2(n10929), .A3(n10928), .A4(n10927), .ZN(
        n10936) );
  AOI22_X1 U13889 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n10425), .B1(
        n12448), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10934) );
  AOI22_X1 U13890 ( .A1(n12450), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__6__SCAN_IN), .B2(n12449), .ZN(n10933) );
  AOI22_X1 U13891 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n12401), .B1(
        n10653), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10932) );
  AOI22_X1 U13892 ( .A1(n12451), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n10404), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10931) );
  NAND4_X1 U13893 ( .A1(n10934), .A2(n10933), .A3(n10932), .A4(n10931), .ZN(
        n10935) );
  NOR2_X1 U13894 ( .A1(n10936), .A2(n10935), .ZN(n19011) );
  AOI22_X1 U13895 ( .A1(n12151), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n10820), 
        .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n10938) );
  NAND2_X1 U13896 ( .A1(n12156), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n10937) );
  OAI211_X1 U13897 ( .C1(n19011), .C2(n10951), .A(n10938), .B(n10937), .ZN(
        n14577) );
  AOI22_X1 U13898 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n10412), .B1(
        n12443), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10942) );
  AOI22_X1 U13899 ( .A1(n10659), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10754), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10941) );
  AOI22_X1 U13900 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n15421), .B1(
        n10850), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10940) );
  AOI22_X1 U13901 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n10658), .B1(
        n10789), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10939) );
  NAND4_X1 U13902 ( .A1(n10942), .A2(n10941), .A3(n10940), .A4(n10939), .ZN(
        n10948) );
  AOI22_X1 U13903 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n10425), .B1(
        n12451), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10946) );
  AOI22_X1 U13904 ( .A1(n12450), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__7__SCAN_IN), .B2(n12449), .ZN(n10945) );
  AOI22_X1 U13905 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n12401), .B1(
        n10404), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10944) );
  AOI22_X1 U13906 ( .A1(n12448), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10653), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10943) );
  NAND4_X1 U13907 ( .A1(n10946), .A2(n10945), .A3(n10944), .A4(n10943), .ZN(
        n10947) );
  NOR2_X1 U13908 ( .A1(n10948), .A2(n10947), .ZN(n14746) );
  AOI22_X1 U13909 ( .A1(n12151), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n10820), 
        .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n10950) );
  NAND2_X1 U13910 ( .A1(n12156), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n10949) );
  OAI211_X1 U13911 ( .C1(n14746), .C2(n10951), .A(n10950), .B(n10949), .ZN(
        n13812) );
  AOI222_X1 U13912 ( .A1(P2_REIP_REG_16__SCAN_IN), .A2(n12156), .B1(n12151), 
        .B2(P2_EAX_REG_16__SCAN_IN), .C1(n10820), .C2(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n13914) );
  INV_X1 U13913 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n10961) );
  INV_X1 U13914 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n14840) );
  INV_X1 U13915 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n19748) );
  OAI222_X1 U13916 ( .A1(n12166), .A2(n10961), .B1(n12165), .B2(n14840), .C1(
        n12167), .C2(n19748), .ZN(n12140) );
  XNOR2_X1 U13917 ( .A(n9870), .B(n12140), .ZN(n14839) );
  AND2_X1 U13918 ( .A1(n10952), .A2(n10531), .ZN(n16213) );
  INV_X1 U13919 ( .A(n16213), .ZN(n10955) );
  NAND2_X1 U13920 ( .A1(n10953), .A2(n15544), .ZN(n16223) );
  NAND2_X1 U13921 ( .A1(n16223), .A2(n9779), .ZN(n10954) );
  NAND2_X1 U13922 ( .A1(n10955), .A2(n10954), .ZN(n10956) );
  NAND2_X1 U13923 ( .A1(n16070), .A2(n21137), .ZN(n10960) );
  INV_X1 U13924 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15328) );
  AOI211_X1 U13925 ( .C1(n13237), .C2(n13240), .A(n15357), .B(n13238), .ZN(
        n21128) );
  NAND2_X1 U13926 ( .A1(n10957), .A2(n21128), .ZN(n15335) );
  INV_X1 U13927 ( .A(n15329), .ZN(n15111) );
  NOR2_X1 U13928 ( .A1(n15328), .A2(n15111), .ZN(n16170) );
  NAND2_X1 U13929 ( .A1(n16172), .A2(n16170), .ZN(n16149) );
  INV_X1 U13930 ( .A(n16149), .ZN(n16158) );
  INV_X1 U13931 ( .A(n10958), .ZN(n10959) );
  NAND2_X1 U13932 ( .A1(n16158), .A2(n10959), .ZN(n15294) );
  AOI21_X1 U13933 ( .B1(n10960), .B2(n15294), .A(n11115), .ZN(n15288) );
  NAND3_X1 U13934 ( .A1(n15288), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        n10961), .ZN(n11009) );
  NAND2_X1 U13935 ( .A1(n10992), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n10964) );
  NAND2_X1 U13936 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n10963) );
  OAI211_X1 U13937 ( .C1(n9775), .C2(n19748), .A(n10964), .B(n10963), .ZN(
        n10965) );
  AOI21_X1 U13938 ( .B1(n14924), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n10965), .ZN(n11005) );
  NAND2_X1 U13939 ( .A1(n14924), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n10970) );
  INV_X1 U13940 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n18926) );
  NAND2_X1 U13941 ( .A1(n10992), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n10967) );
  NAND2_X1 U13942 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n10966) );
  OAI211_X1 U13943 ( .C1(n9775), .C2(n18926), .A(n10967), .B(n10966), .ZN(
        n10968) );
  INV_X1 U13944 ( .A(n10968), .ZN(n10969) );
  NAND2_X1 U13945 ( .A1(n10970), .A2(n10969), .ZN(n15309) );
  INV_X1 U13946 ( .A(n10971), .ZN(n10972) );
  AOI22_X1 U13947 ( .A1(n12209), .A2(P2_REIP_REG_4__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10975) );
  NAND2_X1 U13948 ( .A1(n10992), .A2(P2_EBX_REG_4__SCAN_IN), .ZN(n10974) );
  OAI211_X1 U13949 ( .C1(n10582), .C2(n13850), .A(n10975), .B(n10974), .ZN(
        n13853) );
  INV_X1 U13950 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n13900) );
  NAND2_X1 U13951 ( .A1(n10992), .A2(P2_EBX_REG_5__SCAN_IN), .ZN(n10977) );
  NAND2_X1 U13952 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n10976) );
  OAI211_X1 U13953 ( .C1(n13900), .C2(n9775), .A(n10977), .B(n10976), .ZN(
        n10978) );
  AOI21_X1 U13954 ( .B1(n14924), .B2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(
        n10978), .ZN(n13487) );
  AOI22_X1 U13955 ( .A1(n12209), .A2(P2_REIP_REG_6__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10980) );
  NAND2_X1 U13956 ( .A1(n10992), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n10979) );
  OAI211_X1 U13957 ( .C1(n10582), .C2(n15349), .A(n10980), .B(n10979), .ZN(
        n13570) );
  INV_X1 U13958 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n11061) );
  AOI22_X1 U13959 ( .A1(n12209), .A2(P2_REIP_REG_7__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10981) );
  OAI21_X1 U13960 ( .B1(n10962), .B2(n11061), .A(n10981), .ZN(n10982) );
  AOI21_X1 U13961 ( .B1(n14924), .B2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n10982), .ZN(n13584) );
  INV_X1 U13962 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n11062) );
  NAND2_X1 U13963 ( .A1(n14924), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10984) );
  AOI22_X1 U13964 ( .A1(n12209), .A2(P2_REIP_REG_8__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10983) );
  OAI211_X1 U13965 ( .C1(n11062), .C2(n10962), .A(n10984), .B(n10983), .ZN(
        n14604) );
  INV_X1 U13966 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n11075) );
  AOI22_X1 U13967 ( .A1(n12209), .A2(P2_REIP_REG_9__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10985) );
  OAI21_X1 U13968 ( .B1(n10962), .B2(n11075), .A(n10985), .ZN(n10986) );
  AOI21_X1 U13969 ( .B1(n14924), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n10986), .ZN(n13682) );
  NAND2_X1 U13970 ( .A1(n15309), .A2(n15308), .ZN(n15307) );
  INV_X1 U13971 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n15087) );
  NAND2_X1 U13972 ( .A1(n10992), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n10988) );
  NAND2_X1 U13973 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n10987) );
  OAI211_X1 U13974 ( .C1(n9775), .C2(n15087), .A(n10988), .B(n10987), .ZN(
        n10989) );
  AOI21_X1 U13975 ( .B1(n14924), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n10989), .ZN(n13718) );
  INV_X1 U13976 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n16161) );
  AOI22_X1 U13977 ( .A1(n12209), .A2(P2_REIP_REG_12__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), 
        .ZN(n10991) );
  NAND2_X1 U13978 ( .A1(n10992), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n10990) );
  OAI211_X1 U13979 ( .C1(n10582), .C2(n16161), .A(n10991), .B(n10990), .ZN(
        n14592) );
  INV_X1 U13980 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n10995) );
  NAND2_X1 U13981 ( .A1(n10992), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n10994) );
  NAND2_X1 U13982 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n10993) );
  OAI211_X1 U13983 ( .C1(n9775), .C2(n10995), .A(n10994), .B(n10993), .ZN(
        n10996) );
  AOI21_X1 U13984 ( .B1(n14924), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n10996), .ZN(n13765) );
  NAND2_X1 U13985 ( .A1(n12209), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n10998) );
  NAND2_X1 U13986 ( .A1(n10992), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n10997) );
  OAI211_X1 U13987 ( .C1(n15386), .C2(n16078), .A(n10998), .B(n10997), .ZN(
        n10999) );
  AOI21_X1 U13988 ( .B1(n14924), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n10999), .ZN(n14582) );
  INV_X1 U13989 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n19744) );
  NAND2_X1 U13990 ( .A1(n10992), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n11001) );
  NAND2_X1 U13991 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n11000) );
  OAI211_X1 U13992 ( .C1(n9775), .C2(n19744), .A(n11001), .B(n11000), .ZN(
        n11002) );
  AOI21_X1 U13993 ( .B1(n14924), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n11002), .ZN(n14747) );
  AOI22_X1 U13994 ( .A1(n12209), .A2(P2_REIP_REG_16__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), 
        .ZN(n11004) );
  NAND2_X1 U13995 ( .A1(n10992), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n11003) );
  OAI211_X1 U13996 ( .C1(n10582), .C2(n15290), .A(n11004), .B(n11003), .ZN(
        n15048) );
  NAND2_X1 U13997 ( .A1(n15049), .A2(n15048), .ZN(n15051) );
  AOI21_X1 U13998 ( .B1(n11005), .B2(n15051), .A(n10079), .ZN(n18863) );
  NAND2_X1 U13999 ( .A1(n15416), .A2(n9776), .ZN(n11006) );
  NAND2_X1 U14000 ( .A1(n11006), .A2(n15397), .ZN(n11007) );
  AOI22_X1 U14001 ( .A1(n18863), .A2(n21130), .B1(P2_REIP_REG_17__SCAN_IN), 
        .B2(n16186), .ZN(n11008) );
  OAI211_X1 U14002 ( .C1(n14839), .C2(n21133), .A(n11009), .B(n11008), .ZN(
        n11010) );
  AOI21_X1 U14003 ( .B1(n11011), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n11010), .ZN(n11129) );
  INV_X1 U14004 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n11012) );
  INV_X1 U14005 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n13350) );
  NAND2_X1 U14006 ( .A1(n11012), .A2(n13350), .ZN(n11014) );
  MUX2_X1 U14007 ( .A(n11015), .B(n11014), .S(n14912), .Z(n11026) );
  INV_X1 U14008 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n11017) );
  MUX2_X1 U14009 ( .A(n11018), .B(n11017), .S(n14912), .Z(n11019) );
  NOR2_X1 U14010 ( .A1(n11025), .A2(n11019), .ZN(n11020) );
  OR2_X1 U14011 ( .A1(n11042), .A2(n11020), .ZN(n14641) );
  XNOR2_X1 U14012 ( .A(n11033), .B(n21127), .ZN(n13786) );
  MUX2_X1 U14013 ( .A(n11021), .B(n13350), .S(n14912), .Z(n18995) );
  NOR2_X1 U14014 ( .A1(n18995), .A2(n13263), .ZN(n11024) );
  NAND3_X1 U14015 ( .A1(n14912), .A2(P2_EBX_REG_0__SCAN_IN), .A3(
        P2_EBX_REG_1__SCAN_IN), .ZN(n11022) );
  NAND2_X1 U14016 ( .A1(n11026), .A2(n11022), .ZN(n14669) );
  INV_X1 U14017 ( .A(n14669), .ZN(n11023) );
  NOR2_X1 U14018 ( .A1(n11024), .A2(n11023), .ZN(n13331) );
  AND2_X1 U14019 ( .A1(n11024), .A2(n11023), .ZN(n13330) );
  NOR2_X1 U14020 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n13330), .ZN(
        n13329) );
  NOR2_X1 U14021 ( .A1(n13331), .A2(n13329), .ZN(n13246) );
  INV_X1 U14022 ( .A(n11025), .ZN(n11029) );
  NAND2_X1 U14023 ( .A1(n11027), .A2(n11026), .ZN(n11028) );
  NAND2_X1 U14024 ( .A1(n11029), .A2(n11028), .ZN(n14656) );
  XNOR2_X1 U14025 ( .A(n14656), .B(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13245) );
  NAND2_X1 U14026 ( .A1(n13246), .A2(n13245), .ZN(n11032) );
  INV_X1 U14027 ( .A(n14656), .ZN(n11030) );
  NAND2_X1 U14028 ( .A1(n11030), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11031) );
  NAND2_X1 U14029 ( .A1(n11032), .A2(n11031), .ZN(n13787) );
  NAND2_X1 U14030 ( .A1(n13786), .A2(n13787), .ZN(n11035) );
  NAND2_X1 U14031 ( .A1(n11033), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11034) );
  NAND2_X1 U14032 ( .A1(n11035), .A2(n11034), .ZN(n13847) );
  INV_X1 U14033 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n14624) );
  MUX2_X1 U14034 ( .A(n11036), .B(n14624), .S(n14912), .Z(n11041) );
  XNOR2_X1 U14035 ( .A(n11042), .B(n11041), .ZN(n14627) );
  XNOR2_X1 U14036 ( .A(n14627), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13848) );
  NAND2_X1 U14037 ( .A1(n13847), .A2(n13848), .ZN(n11039) );
  INV_X1 U14038 ( .A(n14627), .ZN(n11037) );
  NAND2_X1 U14039 ( .A1(n11037), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11038) );
  NAND2_X1 U14040 ( .A1(n11039), .A2(n11038), .ZN(n13879) );
  NAND2_X1 U14041 ( .A1(n11040), .A2(n10849), .ZN(n11047) );
  MUX2_X1 U14042 ( .A(n11043), .B(P2_EBX_REG_5__SCAN_IN), .S(n14912), .Z(
        n11044) );
  OR2_X2 U14043 ( .A1(n11045), .A2(n11044), .ZN(n11054) );
  NAND2_X1 U14044 ( .A1(n11045), .A2(n11044), .ZN(n11046) );
  NAND2_X1 U14045 ( .A1(n11054), .A2(n11046), .ZN(n18974) );
  NAND2_X1 U14046 ( .A1(n11047), .A2(n18974), .ZN(n11049) );
  XNOR2_X1 U14047 ( .A(n11049), .B(n11048), .ZN(n13880) );
  NAND2_X1 U14048 ( .A1(n13879), .A2(n13880), .ZN(n11051) );
  NAND2_X1 U14049 ( .A1(n11049), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11050) );
  NAND2_X1 U14050 ( .A1(n11051), .A2(n11050), .ZN(n15345) );
  MUX2_X1 U14051 ( .A(n11052), .B(P2_EBX_REG_6__SCAN_IN), .S(n14912), .Z(
        n11053) );
  AND2_X1 U14052 ( .A1(n11054), .A2(n11053), .ZN(n11055) );
  NOR2_X4 U14053 ( .A1(n11054), .A2(n11053), .ZN(n11067) );
  OR2_X1 U14054 ( .A1(n11055), .A2(n11067), .ZN(n18961) );
  XNOR2_X1 U14055 ( .A(n11057), .B(n15349), .ZN(n15346) );
  NAND2_X1 U14056 ( .A1(n15345), .A2(n15346), .ZN(n11059) );
  NAND2_X1 U14057 ( .A1(n11057), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11058) );
  MUX2_X1 U14058 ( .A(n11061), .B(n11060), .S(n10808), .Z(n11065) );
  NOR2_X1 U14059 ( .A1(n10808), .A2(n11062), .ZN(n11063) );
  NAND2_X1 U14060 ( .A1(n11079), .A2(n11063), .ZN(n11064) );
  NAND2_X1 U14061 ( .A1(n11077), .A2(n11064), .ZN(n14611) );
  NOR2_X1 U14062 ( .A1(n14611), .A2(n10849), .ZN(n11070) );
  AND2_X1 U14063 ( .A1(n11070), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16104) );
  INV_X1 U14064 ( .A(n16104), .ZN(n11069) );
  INV_X1 U14065 ( .A(n11065), .ZN(n11066) );
  XNOR2_X1 U14066 ( .A(n11067), .B(n11066), .ZN(n18951) );
  AND2_X1 U14067 ( .A1(n18951), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16100) );
  INV_X1 U14068 ( .A(n16100), .ZN(n11068) );
  INV_X1 U14069 ( .A(n11070), .ZN(n11072) );
  INV_X1 U14070 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n11071) );
  NAND2_X1 U14071 ( .A1(n11072), .A2(n11071), .ZN(n16102) );
  INV_X1 U14072 ( .A(n18951), .ZN(n11073) );
  NAND2_X1 U14073 ( .A1(n11073), .A2(n15340), .ZN(n16101) );
  AND2_X1 U14074 ( .A1(n16102), .A2(n16101), .ZN(n11074) );
  NOR2_X1 U14075 ( .A1(n10808), .A2(n11075), .ZN(n11076) );
  MUX2_X1 U14076 ( .A(n10808), .B(n11076), .S(n11077), .Z(n11078) );
  NOR2_X1 U14077 ( .A1(n11078), .A2(n11080), .ZN(n18935) );
  AOI21_X1 U14078 ( .B1(n18935), .B2(n11060), .A(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15092) );
  INV_X1 U14079 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n18930) );
  NOR2_X1 U14080 ( .A1(n11080), .A2(n18930), .ZN(n11081) );
  NAND2_X1 U14081 ( .A1(n14912), .A2(n11081), .ZN(n11082) );
  AND2_X1 U14082 ( .A1(n14886), .A2(n11082), .ZN(n11083) );
  NAND2_X1 U14083 ( .A1(n11085), .A2(n11083), .ZN(n18927) );
  INV_X1 U14084 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15306) );
  NAND2_X1 U14085 ( .A1(n11096), .A2(n15306), .ZN(n15316) );
  INV_X1 U14086 ( .A(n11090), .ZN(n11084) );
  NAND2_X1 U14087 ( .A1(P2_EBX_REG_11__SCAN_IN), .A2(n11085), .ZN(n11086) );
  NOR2_X1 U14088 ( .A1(n10808), .A2(n11086), .ZN(n11087) );
  NOR2_X1 U14089 ( .A1(n11089), .A2(n11087), .ZN(n18912) );
  AOI21_X1 U14090 ( .B1(n18912), .B2(n11060), .A(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15080) );
  INV_X1 U14091 ( .A(n15080), .ZN(n11088) );
  NAND2_X1 U14092 ( .A1(n14912), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n11091) );
  NOR2_X1 U14093 ( .A1(n11091), .A2(n11090), .ZN(n11092) );
  NOR2_X1 U14094 ( .A1(n11098), .A2(n11092), .ZN(n14597) );
  AOI21_X1 U14095 ( .B1(n14597), .B2(n11060), .A(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n16082) );
  INV_X1 U14096 ( .A(n18912), .ZN(n11094) );
  NAND2_X1 U14097 ( .A1(n11060), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11093) );
  OR2_X1 U14098 ( .A1(n11094), .A2(n11093), .ZN(n15078) );
  AND2_X1 U14099 ( .A1(n11060), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11095) );
  NAND2_X1 U14100 ( .A1(n18935), .A2(n11095), .ZN(n15091) );
  OR2_X1 U14101 ( .A1(n15306), .A2(n11096), .ZN(n15315) );
  AND2_X1 U14102 ( .A1(n15078), .A2(n9872), .ZN(n16084) );
  AND2_X1 U14103 ( .A1(n11060), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n11097) );
  NAND2_X1 U14104 ( .A1(n14597), .A2(n11097), .ZN(n16083) );
  AND2_X1 U14105 ( .A1(n16084), .A2(n16083), .ZN(n14846) );
  INV_X1 U14106 ( .A(n11110), .ZN(n11100) );
  NAND2_X1 U14107 ( .A1(n10110), .A2(n9893), .ZN(n11099) );
  NAND2_X1 U14108 ( .A1(n11100), .A2(n11099), .ZN(n18900) );
  OR2_X1 U14109 ( .A1(n18900), .A2(n10849), .ZN(n11101) );
  INV_X1 U14110 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16148) );
  OR2_X1 U14111 ( .A1(n11101), .A2(n16148), .ZN(n15069) );
  OAI211_X1 U14112 ( .C1(n16085), .C2(n16082), .A(n14846), .B(n15069), .ZN(
        n11102) );
  NAND2_X1 U14113 ( .A1(n11101), .A2(n16148), .ZN(n15068) );
  NAND2_X1 U14114 ( .A1(n14912), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n11103) );
  MUX2_X1 U14115 ( .A(n11103), .B(n14912), .S(n11110), .Z(n11104) );
  INV_X1 U14116 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n14581) );
  NAND2_X1 U14117 ( .A1(n11110), .A2(n14581), .ZN(n11111) );
  NAND2_X1 U14118 ( .A1(n14574), .A2(n11060), .ZN(n11106) );
  INV_X1 U14119 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n11105) );
  NAND2_X1 U14120 ( .A1(n11106), .A2(n11105), .ZN(n16072) );
  INV_X1 U14121 ( .A(n11106), .ZN(n11107) );
  NAND2_X1 U14122 ( .A1(n11107), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n16073) );
  INV_X1 U14123 ( .A(n16073), .ZN(n11108) );
  AOI21_X2 U14124 ( .B1(n16075), .B2(n16072), .A(n11108), .ZN(n15060) );
  OAI21_X1 U14125 ( .B1(P2_EBX_REG_15__SCAN_IN), .B2(P2_EBX_REG_14__SCAN_IN), 
        .A(n14912), .ZN(n11109) );
  INV_X1 U14126 ( .A(n11119), .ZN(n11113) );
  NAND3_X1 U14127 ( .A1(n11111), .A2(P2_EBX_REG_15__SCAN_IN), .A3(n14912), 
        .ZN(n11112) );
  NAND2_X1 U14128 ( .A1(n11113), .A2(n11112), .ZN(n18883) );
  NAND2_X1 U14129 ( .A1(n11060), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11114) );
  OR2_X1 U14130 ( .A1(n18883), .A2(n11114), .ZN(n15057) );
  OR2_X1 U14131 ( .A1(n18883), .A2(n10849), .ZN(n11116) );
  NAND2_X1 U14132 ( .A1(n11116), .A2(n11115), .ZN(n15058) );
  INV_X1 U14133 ( .A(n15058), .ZN(n11117) );
  NAND2_X1 U14134 ( .A1(n14912), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n11118) );
  INV_X1 U14135 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n19006) );
  OAI211_X1 U14136 ( .C1(n11119), .C2(n11118), .A(n14886), .B(n11122), .ZN(
        n18870) );
  OR2_X1 U14137 ( .A1(n18870), .A2(n10849), .ZN(n11120) );
  XNOR2_X1 U14138 ( .A(n11120), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15047) );
  NAND2_X1 U14139 ( .A1(n11060), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11121) );
  OR2_X1 U14140 ( .A1(n18870), .A2(n11121), .ZN(n14854) );
  NAND2_X1 U14141 ( .A1(n14912), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n12128) );
  XNOR2_X1 U14142 ( .A(n12129), .B(n10114), .ZN(n18859) );
  AOI21_X1 U14143 ( .B1(n18859), .B2(n11060), .A(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n14848) );
  AND2_X1 U14144 ( .A1(n11060), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n11123) );
  NAND2_X1 U14145 ( .A1(n18859), .A2(n11123), .ZN(n14855) );
  NAND2_X1 U14146 ( .A1(n9956), .A2(n14855), .ZN(n11124) );
  XNOR2_X1 U14147 ( .A(n12222), .B(n11124), .ZN(n15044) );
  INV_X1 U14148 ( .A(n15044), .ZN(n11127) );
  INV_X1 U14149 ( .A(n10512), .ZN(n16219) );
  NAND2_X1 U14150 ( .A1(n16219), .A2(n12218), .ZN(n12268) );
  INV_X1 U14151 ( .A(n12268), .ZN(n19827) );
  NAND2_X1 U14152 ( .A1(n11129), .A2(n11128), .ZN(P2_U3029) );
  INV_X1 U14153 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11130) );
  INV_X1 U14154 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11131) );
  AOI22_X1 U14155 ( .A1(n11241), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11210), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11137) );
  INV_X2 U14156 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11132) );
  AND2_X2 U14157 ( .A1(n11132), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11139) );
  AND2_X2 U14158 ( .A1(n13541), .A2(n11139), .ZN(n11234) );
  AND2_X4 U14159 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13446) );
  AOI22_X1 U14160 ( .A1(n11234), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11441), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11136) );
  AOI22_X1 U14161 ( .A1(n11239), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n9827), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11135) );
  AND2_X2 U14162 ( .A1(n11141), .A2(n13546), .ZN(n11232) );
  AOI22_X1 U14163 ( .A1(n11232), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13028), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11134) );
  NAND4_X1 U14164 ( .A1(n11137), .A2(n11136), .A3(n11135), .A4(n11134), .ZN(
        n11147) );
  AND2_X2 U14165 ( .A1(n11141), .A2(n11138), .ZN(n11231) );
  AOI22_X1 U14166 ( .A1(n11231), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11201), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11145) );
  AND2_X2 U14167 ( .A1(n11139), .A2(n11140), .ZN(n11464) );
  AOI22_X1 U14168 ( .A1(n11464), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11233), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11144) );
  AND2_X2 U14169 ( .A1(n11140), .A2(n13446), .ZN(n11238) );
  AOI22_X1 U14170 ( .A1(n11240), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11238), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11143) );
  AOI22_X1 U14171 ( .A1(n11228), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11317), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11142) );
  NAND4_X1 U14172 ( .A1(n11145), .A2(n11144), .A3(n11143), .A4(n11142), .ZN(
        n11146) );
  AOI22_X1 U14173 ( .A1(n11210), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11237), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11148) );
  NAND2_X1 U14174 ( .A1(n11149), .A2(n11148), .ZN(n11153) );
  AOI22_X1 U14175 ( .A1(n11317), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n13028), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11150) );
  NAND2_X1 U14176 ( .A1(n11151), .A2(n11150), .ZN(n11152) );
  BUF_X4 U14177 ( .A(n11240), .Z(n13133) );
  AOI22_X1 U14178 ( .A1(n11241), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11240), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11157) );
  AOI22_X1 U14179 ( .A1(n11201), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11228), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11156) );
  AOI22_X1 U14180 ( .A1(n11464), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11441), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11155) );
  AOI22_X1 U14181 ( .A1(n11232), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11233), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11154) );
  NAND2_X1 U14182 ( .A1(n11159), .A2(n11158), .ZN(n11267) );
  AOI22_X1 U14183 ( .A1(n11240), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11239), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11163) );
  AOI22_X1 U14184 ( .A1(n11232), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11201), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11162) );
  AOI22_X1 U14185 ( .A1(n11234), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11441), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11161) );
  AOI22_X1 U14186 ( .A1(n11228), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n13028), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11160) );
  AOI22_X1 U14187 ( .A1(n11464), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11233), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11167) );
  AOI22_X1 U14188 ( .A1(n11241), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11210), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11166) );
  AOI22_X1 U14189 ( .A1(n9827), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11238), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11165) );
  AOI22_X1 U14190 ( .A1(n11231), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11317), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11164) );
  NAND2_X2 U14191 ( .A1(n9850), .A2(n11168), .ZN(n20122) );
  NAND2_X1 U14192 ( .A1(n11464), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11172) );
  NAND2_X1 U14193 ( .A1(n11234), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11171) );
  NAND2_X1 U14194 ( .A1(n11239), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n11170) );
  NAND2_X1 U14195 ( .A1(n11238), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n11169) );
  NAND2_X1 U14196 ( .A1(n11241), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11176) );
  NAND2_X1 U14197 ( .A1(n13133), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n11175) );
  NAND2_X1 U14198 ( .A1(n11210), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11174) );
  NAND2_X1 U14199 ( .A1(n11237), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11173) );
  NAND2_X1 U14200 ( .A1(n11232), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11180) );
  NAND2_X1 U14201 ( .A1(n11228), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11179) );
  NAND2_X1 U14202 ( .A1(n11233), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n11178) );
  NAND2_X1 U14203 ( .A1(n11317), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n11177) );
  NAND2_X1 U14204 ( .A1(n11231), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n11184) );
  NAND2_X1 U14205 ( .A1(n11201), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11183) );
  NAND2_X1 U14206 ( .A1(n11441), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n11182) );
  NAND2_X1 U14207 ( .A1(n13028), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11181) );
  NAND4_X4 U14208 ( .A1(n11188), .A2(n11187), .A3(n11186), .A4(n11185), .ZN(
        n20113) );
  NAND2_X1 U14209 ( .A1(n11241), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11192) );
  NAND2_X1 U14210 ( .A1(n11240), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n11191) );
  NAND2_X1 U14211 ( .A1(n11210), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n11190) );
  NAND2_X1 U14212 ( .A1(n11237), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11189) );
  NAND2_X1 U14213 ( .A1(n11234), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n11196) );
  NAND2_X1 U14214 ( .A1(n11232), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n11195) );
  NAND2_X1 U14215 ( .A1(n11231), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n11194) );
  NAND2_X1 U14216 ( .A1(n11233), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n11193) );
  NAND2_X1 U14217 ( .A1(n11464), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11200) );
  NAND2_X1 U14218 ( .A1(n11239), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n11199) );
  NAND2_X1 U14219 ( .A1(n11441), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n11198) );
  NAND2_X1 U14220 ( .A1(n11238), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n11197) );
  NAND2_X1 U14221 ( .A1(n11201), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n11205) );
  NAND2_X1 U14222 ( .A1(n11228), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n11204) );
  NAND2_X1 U14223 ( .A1(n13028), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n11203) );
  NAND2_X1 U14224 ( .A1(n11317), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n11202) );
  AND2_X2 U14225 ( .A1(n13153), .A2(n13744), .ZN(n13695) );
  AOI22_X1 U14226 ( .A1(n11241), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11240), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11214) );
  AOI22_X1 U14227 ( .A1(n11239), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11441), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11213) );
  AOI22_X1 U14228 ( .A1(n11210), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11237), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11212) );
  AOI22_X1 U14229 ( .A1(n11464), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11238), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11211) );
  AOI22_X1 U14230 ( .A1(n11234), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11233), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11218) );
  AOI22_X1 U14231 ( .A1(n11228), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11317), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11217) );
  AOI22_X1 U14232 ( .A1(n11232), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11231), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11216) );
  AOI22_X1 U14233 ( .A1(n11201), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9824), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11215) );
  AOI22_X1 U14234 ( .A1(n11241), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n13133), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11223) );
  AOI22_X1 U14235 ( .A1(n11239), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11441), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11222) );
  AOI22_X1 U14236 ( .A1(n11210), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11237), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11221) );
  AOI22_X1 U14237 ( .A1(n11464), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11238), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11220) );
  AOI22_X1 U14238 ( .A1(n11234), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11233), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11227) );
  AOI22_X1 U14239 ( .A1(n11232), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11231), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11226) );
  AOI22_X1 U14240 ( .A1(n11201), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n13028), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11225) );
  AOI22_X1 U14241 ( .A1(n11228), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11317), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11224) );
  INV_X1 U14242 ( .A(n11610), .ZN(n11248) );
  AOI22_X1 U14243 ( .A1(n11228), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11317), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11230) );
  AOI22_X1 U14244 ( .A1(n11201), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n13028), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11229) );
  AOI22_X1 U14245 ( .A1(n11232), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11231), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11236) );
  AOI22_X1 U14246 ( .A1(n11234), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11233), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11235) );
  AOI22_X1 U14247 ( .A1(n11464), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n11238), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11244) );
  AOI22_X1 U14248 ( .A1(n11239), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11441), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11243) );
  AOI22_X1 U14249 ( .A1(n11241), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11240), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11242) );
  AND3_X1 U14250 ( .A1(n9772), .A2(n9823), .A3(n20122), .ZN(n11246) );
  NAND2_X1 U14251 ( .A1(n11258), .A2(n11246), .ZN(n13279) );
  OR2_X2 U14252 ( .A1(n13279), .A2(n13965), .ZN(n11716) );
  XNOR2_X1 U14253 ( .A(P1_STATE_REG_1__SCAN_IN), .B(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n11582) );
  NOR2_X1 U14254 ( .A1(n11248), .A2(n11247), .ZN(n11260) );
  NAND2_X1 U14255 ( .A1(n9788), .A2(n11251), .ZN(n11249) );
  NAND2_X1 U14256 ( .A1(n11249), .A2(n9791), .ZN(n11250) );
  NAND2_X1 U14257 ( .A1(n11722), .A2(n11266), .ZN(n11256) );
  NAND2_X1 U14258 ( .A1(n11260), .A2(n9782), .ZN(n11274) );
  AND2_X1 U14259 ( .A1(n11262), .A2(n13151), .ZN(n11264) );
  NAND2_X1 U14260 ( .A1(n9814), .A2(n11266), .ZN(n11271) );
  NAND2_X2 U14261 ( .A1(n13529), .A2(n9822), .ZN(n11280) );
  NAND2_X1 U14262 ( .A1(n11267), .A2(n9823), .ZN(n11721) );
  OAI21_X2 U14263 ( .B1(n11274), .B2(n11719), .A(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n11345) );
  NAND2_X1 U14264 ( .A1(n20622), .A2(n20538), .ZN(n20485) );
  NAND2_X1 U14265 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20618) );
  NAND2_X1 U14266 ( .A1(n20485), .A2(n20618), .ZN(n20421) );
  OR2_X1 U14267 ( .A1(n20687), .A2(n20622), .ZN(n11341) );
  OAI21_X1 U14268 ( .B1(n13173), .B2(n20421), .A(n11341), .ZN(n11272) );
  INV_X1 U14269 ( .A(n11272), .ZN(n11273) );
  OAI21_X2 U14270 ( .B1(n11345), .B2(n12666), .A(n11273), .ZN(n11275) );
  MUX2_X1 U14271 ( .A(n20687), .B(n13173), .S(n20538), .Z(n11276) );
  NAND2_X1 U14272 ( .A1(n9814), .A2(n13744), .ZN(n11731) );
  NAND2_X1 U14273 ( .A1(n13545), .A2(n9772), .ZN(n11732) );
  NAND2_X1 U14274 ( .A1(n14552), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n19864) );
  INV_X1 U14275 ( .A(n19864), .ZN(n11277) );
  NAND2_X1 U14276 ( .A1(n11732), .A2(n11277), .ZN(n11278) );
  NOR2_X1 U14277 ( .A1(n11279), .A2(n11278), .ZN(n11285) );
  INV_X1 U14278 ( .A(n13744), .ZN(n13277) );
  INV_X2 U14279 ( .A(n11709), .ZN(n11692) );
  AND2_X1 U14280 ( .A1(n13277), .A2(n11692), .ZN(n13293) );
  NAND2_X1 U14281 ( .A1(n11262), .A2(n20122), .ZN(n11281) );
  INV_X1 U14282 ( .A(n11724), .ZN(n11602) );
  INV_X1 U14283 ( .A(n11280), .ZN(n11508) );
  AOI22_X1 U14284 ( .A1(n13293), .A2(n11281), .B1(n11602), .B2(n11508), .ZN(
        n11284) );
  INV_X1 U14285 ( .A(n11282), .ZN(n11600) );
  NAND3_X1 U14286 ( .A1(n11600), .A2(n14548), .A3(n20113), .ZN(n11283) );
  NAND4_X1 U14287 ( .A1(n11731), .A2(n11285), .A3(n11284), .A4(n11283), .ZN(
        n11300) );
  NAND2_X1 U14288 ( .A1(n11302), .A2(n11300), .ZN(n11287) );
  INV_X1 U14289 ( .A(n11287), .ZN(n11286) );
  AOI22_X1 U14290 ( .A1(n11232), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12965), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11292) );
  AOI22_X1 U14291 ( .A1(n13050), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n13128), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11291) );
  AOI22_X1 U14292 ( .A1(n13090), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12867), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11290) );
  AOI22_X1 U14293 ( .A1(n12901), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n9825), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11289) );
  NAND4_X1 U14294 ( .A1(n11292), .A2(n11291), .A3(n11290), .A4(n11289), .ZN(
        n11298) );
  AOI22_X1 U14295 ( .A1(n11464), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n11441), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11296) );
  AOI22_X1 U14296 ( .A1(n12978), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12957), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11295) );
  AOI22_X1 U14297 ( .A1(n13112), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12964), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11294) );
  AOI22_X1 U14298 ( .A1(n12921), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n13134), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11293) );
  NAND4_X1 U14299 ( .A1(n11296), .A2(n11295), .A3(n11294), .A4(n11293), .ZN(
        n11297) );
  NAND2_X1 U14300 ( .A1(n11361), .A2(n11371), .ZN(n11299) );
  INV_X1 U14301 ( .A(n11370), .ZN(n11338) );
  INV_X1 U14302 ( .A(n11300), .ZN(n11301) );
  NAND2_X1 U14303 ( .A1(n12672), .A2(n20098), .ZN(n11327) );
  AOI22_X1 U14304 ( .A1(n13050), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n13133), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11306) );
  AOI22_X1 U14305 ( .A1(n13128), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11441), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11305) );
  AOI22_X1 U14306 ( .A1(n12921), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12964), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11304) );
  AOI22_X1 U14307 ( .A1(n11464), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n13134), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11303) );
  NAND4_X1 U14308 ( .A1(n11306), .A2(n11305), .A3(n11304), .A4(n11303), .ZN(
        n11312) );
  AOI22_X1 U14309 ( .A1(n12937), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n13090), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11310) );
  AOI22_X1 U14310 ( .A1(n12978), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12867), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11309) );
  AOI22_X1 U14311 ( .A1(n12965), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9825), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11308) );
  AOI22_X1 U14312 ( .A1(n11228), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11317), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11307) );
  NAND4_X1 U14313 ( .A1(n11310), .A2(n11309), .A3(n11308), .A4(n11307), .ZN(
        n11311) );
  NAND2_X1 U14314 ( .A1(n13151), .A2(n11491), .ZN(n11324) );
  AOI22_X1 U14315 ( .A1(n13050), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n13133), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11316) );
  AOI22_X1 U14316 ( .A1(n12978), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n13090), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11315) );
  AOI22_X1 U14317 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n11441), .B1(
        n13134), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11314) );
  AOI22_X1 U14318 ( .A1(n12901), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n9825), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11313) );
  NAND4_X1 U14319 ( .A1(n11316), .A2(n11315), .A3(n11314), .A4(n11313), .ZN(
        n11323) );
  AOI22_X1 U14320 ( .A1(n11464), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n13128), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11321) );
  AOI22_X1 U14321 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n12937), .B1(
        n12867), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11320) );
  AOI22_X1 U14322 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n12921), .B1(
        n12964), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11319) );
  AOI22_X1 U14323 ( .A1(n12965), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11317), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11318) );
  NAND4_X1 U14324 ( .A1(n11321), .A2(n11320), .A3(n11319), .A4(n11318), .ZN(
        n11322) );
  MUX2_X1 U14325 ( .A(n11503), .B(n11324), .S(n11382), .Z(n11325) );
  INV_X1 U14326 ( .A(n11325), .ZN(n11326) );
  NAND2_X1 U14327 ( .A1(n11326), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11377) );
  NAND2_X1 U14328 ( .A1(n11327), .A2(n11377), .ZN(n11331) );
  NAND2_X1 U14329 ( .A1(n11571), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11330) );
  AOI21_X1 U14330 ( .B1(n11266), .B2(n11382), .A(n20098), .ZN(n11328) );
  AND2_X1 U14331 ( .A1(n11328), .A2(n11503), .ZN(n11329) );
  NAND2_X1 U14332 ( .A1(n11330), .A2(n11329), .ZN(n11376) );
  NAND2_X1 U14333 ( .A1(n11331), .A2(n11376), .ZN(n11380) );
  INV_X1 U14334 ( .A(n11503), .ZN(n11332) );
  NAND2_X1 U14335 ( .A1(n11332), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11333) );
  NOR2_X1 U14336 ( .A1(n9823), .A2(n20098), .ZN(n11364) );
  AOI22_X1 U14337 ( .A1(n11361), .A2(n11491), .B1(n11364), .B2(n11371), .ZN(
        n11335) );
  NAND2_X1 U14338 ( .A1(n11571), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11334) );
  INV_X1 U14339 ( .A(n11337), .ZN(n11339) );
  NAND2_X1 U14340 ( .A1(n11339), .A2(n11338), .ZN(n11340) );
  INV_X1 U14341 ( .A(n11341), .ZN(n11343) );
  INV_X1 U14342 ( .A(n13173), .ZN(n11395) );
  XNOR2_X1 U14343 ( .A(n20618), .B(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n20108) );
  NAND2_X1 U14344 ( .A1(n11395), .A2(n20108), .ZN(n11347) );
  INV_X1 U14345 ( .A(n20687), .ZN(n11394) );
  NAND2_X1 U14346 ( .A1(n11394), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11346) );
  NAND2_X1 U14347 ( .A1(n11391), .A2(n11350), .ZN(n13437) );
  AOI22_X1 U14348 ( .A1(n13050), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n13133), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11354) );
  AOI22_X1 U14349 ( .A1(n13128), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11441), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11353) );
  AOI22_X1 U14350 ( .A1(n11210), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12964), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11352) );
  AOI22_X1 U14351 ( .A1(n11464), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n13134), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11351) );
  NAND4_X1 U14352 ( .A1(n11354), .A2(n11353), .A3(n11352), .A4(n11351), .ZN(
        n11360) );
  AOI22_X1 U14353 ( .A1(n11232), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n13090), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11358) );
  AOI22_X1 U14354 ( .A1(n12978), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12867), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11357) );
  AOI22_X1 U14355 ( .A1(n12965), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9825), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11356) );
  AOI22_X1 U14356 ( .A1(n12901), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12957), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11355) );
  NAND4_X1 U14357 ( .A1(n11358), .A2(n11357), .A3(n11356), .A4(n11355), .ZN(
        n11359) );
  INV_X1 U14358 ( .A(n11361), .ZN(n11362) );
  AOI22_X1 U14359 ( .A1(n11571), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11364), .B2(n11363), .ZN(n11365) );
  NAND2_X1 U14360 ( .A1(n14543), .A2(n11541), .ZN(n11369) );
  NAND2_X1 U14361 ( .A1(n11371), .A2(n11382), .ZN(n11412) );
  XNOR2_X1 U14362 ( .A(n11412), .B(n11411), .ZN(n11367) );
  NAND2_X1 U14363 ( .A1(n11266), .A2(n20122), .ZN(n11381) );
  INV_X1 U14364 ( .A(n11381), .ZN(n11366) );
  AOI21_X1 U14365 ( .B1(n11367), .B2(n11508), .A(n11366), .ZN(n11368) );
  NAND2_X1 U14366 ( .A1(n11369), .A2(n11368), .ZN(n13690) );
  OR2_X1 U14367 ( .A1(n11370), .A2(n9787), .ZN(n11375) );
  OAI21_X1 U14368 ( .B1(n11371), .B2(n11382), .A(n11412), .ZN(n11372) );
  OAI211_X1 U14369 ( .C1(n11372), .C2(n11280), .A(n9791), .B(n11251), .ZN(
        n11373) );
  INV_X1 U14370 ( .A(n11373), .ZN(n11374) );
  INV_X1 U14371 ( .A(n11376), .ZN(n11378) );
  NAND2_X1 U14372 ( .A1(n11378), .A2(n11377), .ZN(n11379) );
  INV_X1 U14373 ( .A(n11541), .ZN(n11385) );
  OAI21_X1 U14374 ( .B1(n11280), .B2(n11382), .A(n11381), .ZN(n11383) );
  INV_X1 U14375 ( .A(n11383), .ZN(n11384) );
  OAI21_X2 U14376 ( .B1(n12670), .B2(n11385), .A(n11384), .ZN(n13413) );
  INV_X1 U14377 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n20090) );
  NAND2_X1 U14378 ( .A1(n13690), .A2(n13691), .ZN(n13689) );
  NAND2_X1 U14379 ( .A1(n11386), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11387) );
  INV_X1 U14380 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n20069) );
  INV_X1 U14381 ( .A(n11388), .ZN(n11390) );
  NAND2_X1 U14382 ( .A1(n11390), .A2(n11389), .ZN(n11419) );
  OAI21_X1 U14383 ( .B1(n20618), .B2(n20367), .A(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n11393) );
  INV_X1 U14384 ( .A(n20618), .ZN(n20215) );
  INV_X1 U14385 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20773) );
  NAND2_X1 U14386 ( .A1(n20773), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n20311) );
  INV_X1 U14387 ( .A(n20311), .ZN(n11392) );
  NAND2_X1 U14388 ( .A1(n20215), .A2(n11392), .ZN(n20338) );
  NAND2_X1 U14389 ( .A1(n11393), .A2(n20338), .ZN(n20103) );
  AOI22_X1 U14390 ( .A1(n11395), .A2(n20103), .B1(n11394), .B2(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n11396) );
  INV_X1 U14391 ( .A(n11577), .ZN(n11560) );
  AOI22_X1 U14392 ( .A1(n13050), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n13133), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11402) );
  AOI22_X1 U14393 ( .A1(n13128), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n13540), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11401) );
  AOI22_X1 U14394 ( .A1(n11210), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12964), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11400) );
  AOI22_X1 U14395 ( .A1(n11398), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n13134), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11399) );
  NAND4_X1 U14396 ( .A1(n11402), .A2(n11401), .A3(n11400), .A4(n11399), .ZN(
        n11408) );
  AOI22_X1 U14397 ( .A1(n12937), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n13090), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11406) );
  AOI22_X1 U14398 ( .A1(n12978), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12867), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11405) );
  AOI22_X1 U14399 ( .A1(n12965), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9825), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11404) );
  AOI22_X1 U14400 ( .A1(n12901), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11317), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11403) );
  NAND4_X1 U14401 ( .A1(n11406), .A2(n11405), .A3(n11404), .A4(n11403), .ZN(
        n11407) );
  AOI22_X1 U14402 ( .A1(n11560), .A2(n11454), .B1(n11571), .B2(
        P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11409) );
  NAND2_X1 U14403 ( .A1(n20763), .A2(n11541), .ZN(n11416) );
  NAND2_X1 U14404 ( .A1(n11412), .A2(n11411), .ZN(n11456) );
  INV_X1 U14405 ( .A(n11454), .ZN(n11413) );
  XNOR2_X1 U14406 ( .A(n11456), .B(n11413), .ZN(n11414) );
  NAND2_X1 U14407 ( .A1(n11414), .A2(n11508), .ZN(n11415) );
  NAND2_X1 U14408 ( .A1(n11416), .A2(n11415), .ZN(n13710) );
  NAND2_X1 U14409 ( .A1(n11417), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11418) );
  NAND2_X2 U14410 ( .A1(n13709), .A2(n11418), .ZN(n11437) );
  INV_X1 U14411 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n20061) );
  NAND2_X1 U14412 ( .A1(n11571), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11432) );
  AOI22_X1 U14413 ( .A1(n13050), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n13133), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11423) );
  AOI22_X1 U14414 ( .A1(n13128), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n13540), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11422) );
  AOI22_X1 U14415 ( .A1(n11210), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12964), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11421) );
  AOI22_X1 U14416 ( .A1(n11398), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n13134), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11420) );
  NAND4_X1 U14417 ( .A1(n11423), .A2(n11422), .A3(n11421), .A4(n11420), .ZN(
        n11429) );
  AOI22_X1 U14418 ( .A1(n12937), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n13090), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11427) );
  AOI22_X1 U14419 ( .A1(n12978), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12867), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11426) );
  INV_X1 U14420 ( .A(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n20936) );
  AOI22_X1 U14421 ( .A1(n12965), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n9825), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11425) );
  AOI22_X1 U14422 ( .A1(n12901), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n11317), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11424) );
  NAND4_X1 U14423 ( .A1(n11427), .A2(n11426), .A3(n11425), .A4(n11424), .ZN(
        n11428) );
  INV_X1 U14424 ( .A(n11453), .ZN(n11430) );
  XNOR2_X1 U14425 ( .A(n11439), .B(n11440), .ZN(n12700) );
  NAND2_X1 U14426 ( .A1(n12700), .A2(n11541), .ZN(n11436) );
  NAND2_X1 U14427 ( .A1(n11456), .A2(n11454), .ZN(n11433) );
  XNOR2_X1 U14428 ( .A(n11433), .B(n11453), .ZN(n11434) );
  NAND2_X1 U14429 ( .A1(n11434), .A2(n11508), .ZN(n11435) );
  NAND2_X1 U14430 ( .A1(n11436), .A2(n11435), .ZN(n20034) );
  NAND2_X1 U14431 ( .A1(n11437), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11438) );
  INV_X1 U14432 ( .A(n11571), .ZN(n11566) );
  INV_X1 U14433 ( .A(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11452) );
  AOI22_X1 U14434 ( .A1(n13050), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13133), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11445) );
  AOI22_X1 U14435 ( .A1(n13128), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n13540), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11444) );
  AOI22_X1 U14436 ( .A1(n11210), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12964), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11443) );
  AOI22_X1 U14437 ( .A1(n11398), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n13134), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11442) );
  NAND4_X1 U14438 ( .A1(n11445), .A2(n11444), .A3(n11443), .A4(n11442), .ZN(
        n11451) );
  AOI22_X1 U14439 ( .A1(n12937), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n13090), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11449) );
  AOI22_X1 U14440 ( .A1(n12978), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12867), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11448) );
  AOI22_X1 U14441 ( .A1(n12965), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9825), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11447) );
  AOI22_X1 U14442 ( .A1(n12901), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11317), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11446) );
  NAND4_X1 U14443 ( .A1(n11449), .A2(n11448), .A3(n11447), .A4(n11446), .ZN(
        n11450) );
  OAI22_X1 U14444 ( .A1(n11566), .A2(n11452), .B1(n11577), .B2(n11482), .ZN(
        n11463) );
  NAND2_X1 U14445 ( .A1(n12707), .A2(n11541), .ZN(n11460) );
  AND2_X1 U14446 ( .A1(n11454), .A2(n11453), .ZN(n11455) );
  NAND2_X1 U14447 ( .A1(n11456), .A2(n11455), .ZN(n11483) );
  XNOR2_X1 U14448 ( .A(n11483), .B(n11457), .ZN(n11458) );
  NAND2_X1 U14449 ( .A1(n11458), .A2(n11508), .ZN(n11459) );
  NAND2_X1 U14450 ( .A1(n11460), .A2(n11459), .ZN(n11461) );
  INV_X1 U14451 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n20974) );
  XNOR2_X1 U14452 ( .A(n11461), .B(n20974), .ZN(n15794) );
  AOI22_X1 U14453 ( .A1(n13050), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n13112), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11468) );
  AOI22_X1 U14454 ( .A1(n13128), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n13540), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11467) );
  AOI22_X1 U14455 ( .A1(n12921), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12964), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11466) );
  AOI22_X1 U14456 ( .A1(n11398), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n13134), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11465) );
  NAND4_X1 U14457 ( .A1(n11468), .A2(n11467), .A3(n11466), .A4(n11465), .ZN(
        n11474) );
  AOI22_X1 U14458 ( .A1(n12937), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n13090), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11472) );
  AOI22_X1 U14459 ( .A1(n12978), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12867), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11471) );
  AOI22_X1 U14460 ( .A1(n12965), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9825), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11470) );
  AOI22_X1 U14461 ( .A1(n12901), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11317), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11469) );
  NAND4_X1 U14462 ( .A1(n11472), .A2(n11471), .A3(n11470), .A4(n11469), .ZN(
        n11473) );
  INV_X1 U14463 ( .A(n11496), .ZN(n11475) );
  INV_X1 U14464 ( .A(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11478) );
  OAI21_X1 U14465 ( .B1(n11566), .B2(n11478), .A(n11477), .ZN(n11479) );
  INV_X1 U14466 ( .A(n11479), .ZN(n11480) );
  NAND2_X1 U14467 ( .A1(n11481), .A2(n11480), .ZN(n12711) );
  OR2_X1 U14468 ( .A1(n11483), .A2(n11482), .ZN(n11495) );
  XNOR2_X1 U14469 ( .A(n11495), .B(n11496), .ZN(n11484) );
  NAND2_X1 U14470 ( .A1(n11484), .A2(n11508), .ZN(n11485) );
  NAND2_X1 U14471 ( .A1(n15788), .A2(n15898), .ZN(n11487) );
  INV_X1 U14472 ( .A(n15788), .ZN(n11488) );
  NAND2_X1 U14473 ( .A1(n11488), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11489) );
  INV_X1 U14474 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11492) );
  OAI22_X1 U14475 ( .A1(n11566), .A2(n11492), .B1(n11577), .B2(n11491), .ZN(
        n11493) );
  INV_X1 U14476 ( .A(n11495), .ZN(n11497) );
  NAND2_X1 U14477 ( .A1(n11497), .A2(n11496), .ZN(n11506) );
  XNOR2_X1 U14478 ( .A(n11506), .B(n11507), .ZN(n11498) );
  AND2_X1 U14479 ( .A1(n11498), .A2(n11508), .ZN(n11499) );
  AOI21_X1 U14480 ( .B1(n12720), .B2(n11541), .A(n11499), .ZN(n11500) );
  INV_X1 U14481 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n15911) );
  NAND2_X1 U14482 ( .A1(n11500), .A2(n15911), .ZN(n15783) );
  NAND2_X1 U14483 ( .A1(n15781), .A2(n15783), .ZN(n11502) );
  INV_X1 U14484 ( .A(n11500), .ZN(n11501) );
  NAND2_X1 U14485 ( .A1(n11501), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15782) );
  NAND2_X1 U14486 ( .A1(n11541), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11504) );
  NOR2_X1 U14487 ( .A1(n11504), .A2(n11503), .ZN(n11505) );
  INV_X1 U14488 ( .A(n11506), .ZN(n11509) );
  NAND3_X1 U14489 ( .A1(n11509), .A2(n11508), .A3(n11507), .ZN(n11510) );
  INV_X1 U14490 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n11511) );
  NAND2_X1 U14491 ( .A1(n13924), .A2(n11511), .ZN(n11512) );
  INV_X1 U14492 ( .A(n13924), .ZN(n11513) );
  NAND2_X1 U14493 ( .A1(n11513), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11514) );
  INV_X1 U14494 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n13937) );
  NAND2_X1 U14495 ( .A1(n14352), .A2(n13937), .ZN(n11515) );
  AND2_X2 U14496 ( .A1(n14431), .A2(n11515), .ZN(n14394) );
  INV_X1 U14497 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n11516) );
  NAND2_X1 U14498 ( .A1(n14352), .A2(n11516), .ZN(n14421) );
  NAND2_X1 U14499 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n11517) );
  NAND2_X1 U14500 ( .A1(n14352), .A2(n11517), .ZN(n14419) );
  AND2_X1 U14501 ( .A1(n14421), .A2(n14419), .ZN(n11518) );
  XNOR2_X1 U14502 ( .A(n14352), .B(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n14422) );
  INV_X1 U14503 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n14408) );
  NAND2_X1 U14504 ( .A1(n14352), .A2(n14408), .ZN(n11519) );
  INV_X1 U14505 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15847) );
  NAND2_X1 U14506 ( .A1(n15847), .A2(n14408), .ZN(n11520) );
  XNOR2_X1 U14507 ( .A(n14352), .B(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14400) );
  NAND2_X1 U14508 ( .A1(n14352), .A2(n15824), .ZN(n14524) );
  AND2_X1 U14509 ( .A1(n14400), .A2(n14524), .ZN(n11521) );
  INV_X1 U14510 ( .A(n14510), .ZN(n11522) );
  INV_X1 U14511 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n11667) );
  NAND2_X1 U14512 ( .A1(n11524), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n14420) );
  INV_X1 U14513 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n11648) );
  NAND2_X1 U14514 ( .A1(n11648), .A2(n15868), .ZN(n11523) );
  NAND2_X1 U14515 ( .A1(n11524), .A2(n11523), .ZN(n14417) );
  INV_X1 U14516 ( .A(n11526), .ZN(n11525) );
  INV_X1 U14517 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n14370) );
  INV_X1 U14518 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14379) );
  AND2_X1 U14519 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n11754) );
  NAND2_X1 U14520 ( .A1(n11754), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14455) );
  INV_X1 U14521 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14325) );
  NOR2_X1 U14522 ( .A1(n11526), .A2(n11524), .ZN(n14333) );
  AND2_X1 U14523 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14438) );
  NAND2_X1 U14524 ( .A1(n14352), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11768) );
  INV_X1 U14525 ( .A(n12287), .ZN(n11528) );
  NOR2_X1 U14526 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14439) );
  OR3_X1 U14527 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n13162) );
  OAI21_X1 U14528 ( .B1(n14354), .B2(n13162), .A(n11524), .ZN(n14318) );
  INV_X1 U14529 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n11774) );
  NAND2_X1 U14530 ( .A1(n11524), .A2(n11774), .ZN(n12284) );
  NAND2_X1 U14531 ( .A1(n20538), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11538) );
  XNOR2_X1 U14532 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11545) );
  NAND2_X1 U14533 ( .A1(n11546), .A2(n11545), .ZN(n11531) );
  NAND2_X1 U14534 ( .A1(n20622), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11530) );
  NAND2_X1 U14535 ( .A1(n11531), .A2(n11530), .ZN(n11557) );
  XNOR2_X1 U14536 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n11556) );
  NAND2_X1 U14537 ( .A1(n11557), .A2(n11556), .ZN(n11533) );
  NAND2_X1 U14538 ( .A1(n20367), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11532) );
  MUX2_X1 U14539 ( .A(n20773), .B(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .S(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n11564) );
  NAND2_X1 U14540 ( .A1(n11565), .A2(n11564), .ZN(n11535) );
  NAND2_X1 U14541 ( .A1(n20773), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11534) );
  NAND2_X1 U14542 ( .A1(n11535), .A2(n11534), .ZN(n11570) );
  AND2_X1 U14543 ( .A1(n20869), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n11536) );
  NAND2_X1 U14544 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n13475), .ZN(
        n11569) );
  OAI21_X1 U14545 ( .B1(n20538), .B2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n11538), .ZN(n11542) );
  INV_X1 U14546 ( .A(n11542), .ZN(n11539) );
  AOI21_X1 U14547 ( .B1(n9795), .B2(n11539), .A(n11266), .ZN(n11544) );
  AOI21_X1 U14548 ( .B1(n14222), .B2(n9822), .A(n20113), .ZN(n11559) );
  NOR2_X1 U14549 ( .A1(n11577), .A2(n11542), .ZN(n11543) );
  OAI22_X1 U14550 ( .A1(n11544), .A2(n11559), .B1(n11579), .B2(n11543), .ZN(
        n11551) );
  INV_X1 U14551 ( .A(n11551), .ZN(n11555) );
  XNOR2_X1 U14552 ( .A(n11546), .B(n11545), .ZN(n11589) );
  NOR2_X1 U14553 ( .A1(n11251), .A2(n20098), .ZN(n11548) );
  NOR2_X1 U14554 ( .A1(n11577), .A2(n9787), .ZN(n11547) );
  AOI211_X1 U14555 ( .C1(n11571), .C2(n11589), .A(n11548), .B(n11547), .ZN(
        n11552) );
  INV_X1 U14556 ( .A(n11552), .ZN(n11554) );
  INV_X1 U14557 ( .A(n11548), .ZN(n11549) );
  NAND3_X1 U14558 ( .A1(n11577), .A2(n20113), .A3(n11549), .ZN(n11550) );
  AOI22_X1 U14559 ( .A1(n11552), .A2(n11551), .B1(n11589), .B2(n11550), .ZN(
        n11553) );
  AOI21_X1 U14560 ( .B1(n11555), .B2(n11554), .A(n11553), .ZN(n11563) );
  XNOR2_X1 U14561 ( .A(n11557), .B(n11556), .ZN(n11588) );
  NOR2_X1 U14562 ( .A1(n11577), .A2(n11588), .ZN(n11558) );
  AOI211_X1 U14563 ( .C1(n11571), .C2(n11588), .A(n11559), .B(n11558), .ZN(
        n11562) );
  NAND2_X1 U14564 ( .A1(n11560), .A2(n11559), .ZN(n11561) );
  OAI22_X1 U14565 ( .A1(n11563), .A2(n11562), .B1(n11588), .B2(n11561), .ZN(
        n11568) );
  XNOR2_X1 U14566 ( .A(n11565), .B(n11564), .ZN(n11587) );
  NAND2_X1 U14567 ( .A1(n11566), .A2(n11587), .ZN(n11567) );
  AOI22_X1 U14568 ( .A1(n11568), .A2(n11567), .B1(n11579), .B2(n11587), .ZN(
        n11574) );
  NOR2_X1 U14569 ( .A1(n11571), .A2(n11592), .ZN(n11573) );
  INV_X1 U14570 ( .A(n11579), .ZN(n11572) );
  NAND2_X1 U14571 ( .A1(n11579), .A2(n11578), .ZN(n11580) );
  INV_X1 U14572 ( .A(n11582), .ZN(n11583) );
  NAND2_X1 U14573 ( .A1(n11583), .A2(n20698), .ZN(n15631) );
  INV_X1 U14574 ( .A(n15631), .ZN(n13459) );
  OR2_X1 U14575 ( .A1(n20113), .A2(n13459), .ZN(n13218) );
  NAND2_X1 U14576 ( .A1(READY11_REG_SCAN_IN), .A2(READY1), .ZN(n20697) );
  NAND2_X1 U14577 ( .A1(n13218), .A2(n20697), .ZN(n11585) );
  OAI211_X1 U14578 ( .C1(n13698), .C2(n11585), .A(n9823), .B(n11584), .ZN(
        n11586) );
  NAND2_X1 U14579 ( .A1(n13423), .A2(n11586), .ZN(n11596) );
  NAND2_X1 U14580 ( .A1(n20113), .A2(n15631), .ZN(n11594) );
  OR3_X1 U14581 ( .A1(n11589), .A2(n11588), .A3(n11587), .ZN(n11590) );
  NAND2_X1 U14582 ( .A1(n11591), .A2(n11590), .ZN(n11593) );
  NOR2_X1 U14583 ( .A1(n15630), .A2(n13282), .ZN(n13463) );
  NAND2_X1 U14584 ( .A1(n11594), .A2(n13463), .ZN(n11595) );
  MUX2_X1 U14585 ( .A(n11596), .B(n11595), .S(n11267), .Z(n11608) );
  OR2_X1 U14586 ( .A1(n11262), .A2(n9787), .ZN(n11718) );
  INV_X1 U14587 ( .A(n11718), .ZN(n11606) );
  AND2_X1 U14588 ( .A1(n11718), .A2(n9823), .ZN(n11599) );
  NAND2_X1 U14589 ( .A1(n11600), .A2(n11599), .ZN(n11730) );
  NAND2_X1 U14590 ( .A1(n9791), .A2(n20122), .ZN(n11601) );
  NOR2_X1 U14591 ( .A1(n11602), .A2(n11601), .ZN(n11604) );
  NAND2_X1 U14592 ( .A1(n14548), .A2(n11266), .ZN(n11603) );
  OR2_X1 U14593 ( .A1(n11262), .A2(n20127), .ZN(n11726) );
  AND2_X1 U14594 ( .A1(n11730), .A2(n11611), .ZN(n11605) );
  NOR2_X1 U14595 ( .A1(n11598), .A2(n11605), .ZN(n13456) );
  AOI21_X1 U14596 ( .B1(n13466), .B2(n11606), .A(n13456), .ZN(n11607) );
  NAND2_X1 U14597 ( .A1(n11608), .A2(n11607), .ZN(n11609) );
  NAND2_X1 U14598 ( .A1(n11611), .A2(n13744), .ZN(n13465) );
  NAND2_X1 U14599 ( .A1(n11611), .A2(n11722), .ZN(n13168) );
  AND2_X1 U14600 ( .A1(n13465), .A2(n13168), .ZN(n13280) );
  OAI21_X1 U14601 ( .B1(n13151), .B2(n11610), .A(n13280), .ZN(n11612) );
  OR2_X1 U14602 ( .A1(n11612), .A2(n9786), .ZN(n11613) );
  INV_X1 U14603 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n13578) );
  NAND2_X1 U14604 ( .A1(n11623), .A2(n13578), .ZN(n11617) );
  INV_X1 U14605 ( .A(n20122), .ZN(n11614) );
  NAND2_X1 U14606 ( .A1(n11614), .A2(n9823), .ZN(n11629) );
  INV_X1 U14607 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20075) );
  NAND2_X1 U14608 ( .A1(n11629), .A2(n20075), .ZN(n11615) );
  OAI211_X1 U14609 ( .C1(n13276), .C2(P1_EBX_REG_1__SCAN_IN), .A(n11615), .B(
        n11692), .ZN(n11616) );
  NAND2_X1 U14610 ( .A1(n11617), .A2(n11616), .ZN(n11621) );
  NAND2_X1 U14611 ( .A1(n11629), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n11620) );
  INV_X1 U14612 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n11618) );
  NAND2_X1 U14613 ( .A1(n11692), .A2(n11618), .ZN(n11619) );
  NAND2_X1 U14614 ( .A1(n11620), .A2(n11619), .ZN(n13561) );
  XNOR2_X1 U14615 ( .A(n11621), .B(n13561), .ZN(n13749) );
  INV_X1 U14616 ( .A(n11624), .ZN(n13696) );
  NAND2_X1 U14617 ( .A1(n13749), .A2(n13696), .ZN(n11622) );
  NAND2_X1 U14618 ( .A1(n11622), .A2(n11621), .ZN(n13625) );
  INV_X1 U14619 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n13627) );
  NAND2_X1 U14620 ( .A1(n11623), .A2(n13627), .ZN(n11627) );
  NAND2_X1 U14621 ( .A1(n11696), .A2(n20090), .ZN(n11625) );
  OAI211_X1 U14622 ( .C1(n13276), .C2(P1_EBX_REG_2__SCAN_IN), .A(n11625), .B(
        n11692), .ZN(n11626) );
  AND2_X1 U14623 ( .A1(n11627), .A2(n11626), .ZN(n13624) );
  NAND2_X1 U14624 ( .A1(n11696), .A2(n11692), .ZN(n13560) );
  MUX2_X1 U14625 ( .A(n11700), .B(n11692), .S(P1_EBX_REG_3__SCAN_IN), .Z(
        n11628) );
  OAI21_X1 U14626 ( .B1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n13560), .A(
        n11628), .ZN(n13735) );
  MUX2_X1 U14627 ( .A(n11708), .B(n11696), .S(P1_EBX_REG_4__SCAN_IN), .Z(
        n11631) );
  INV_X1 U14628 ( .A(n11629), .ZN(n11630) );
  NAND2_X1 U14629 ( .A1(n11630), .A2(n13276), .ZN(n11686) );
  OAI211_X1 U14630 ( .C1(n13696), .C2(n20061), .A(n11631), .B(n11686), .ZN(
        n13739) );
  OR2_X1 U14631 ( .A1(n11700), .A2(P1_EBX_REG_5__SCAN_IN), .ZN(n11634) );
  NAND2_X1 U14632 ( .A1(n11692), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11632) );
  OAI211_X1 U14633 ( .C1(n13276), .C2(P1_EBX_REG_5__SCAN_IN), .A(n11696), .B(
        n11632), .ZN(n11633) );
  NAND2_X1 U14634 ( .A1(n11634), .A2(n11633), .ZN(n15918) );
  MUX2_X1 U14635 ( .A(n11708), .B(n11696), .S(P1_EBX_REG_6__SCAN_IN), .Z(
        n11638) );
  NAND2_X1 U14636 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n13276), .ZN(
        n11636) );
  AND2_X1 U14637 ( .A1(n11686), .A2(n11636), .ZN(n11637) );
  OR2_X1 U14638 ( .A1(n11700), .A2(P1_EBX_REG_7__SCAN_IN), .ZN(n11641) );
  NAND2_X1 U14639 ( .A1(n11692), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11639) );
  OAI211_X1 U14640 ( .C1(n13276), .C2(P1_EBX_REG_7__SCAN_IN), .A(n11696), .B(
        n11639), .ZN(n11640) );
  NAND2_X1 U14641 ( .A1(n11641), .A2(n11640), .ZN(n13874) );
  MUX2_X1 U14642 ( .A(n11708), .B(n11696), .S(P1_EBX_REG_8__SCAN_IN), .Z(
        n11644) );
  NAND2_X1 U14643 ( .A1(n13276), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11642) );
  AND2_X1 U14644 ( .A1(n11686), .A2(n11642), .ZN(n11643) );
  NAND2_X1 U14645 ( .A1(n11644), .A2(n11643), .ZN(n13896) );
  OR2_X1 U14646 ( .A1(n11700), .A2(P1_EBX_REG_9__SCAN_IN), .ZN(n11647) );
  NAND2_X1 U14647 ( .A1(n11692), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11645) );
  OAI211_X1 U14648 ( .C1(n13276), .C2(P1_EBX_REG_9__SCAN_IN), .A(n11696), .B(
        n11645), .ZN(n11646) );
  INV_X1 U14649 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n13930) );
  NAND2_X1 U14650 ( .A1(n11623), .A2(n13930), .ZN(n11651) );
  NAND2_X1 U14651 ( .A1(n11696), .A2(n11648), .ZN(n11649) );
  OAI211_X1 U14652 ( .C1(n13276), .C2(P1_EBX_REG_10__SCAN_IN), .A(n11649), .B(
        n11692), .ZN(n11650) );
  OR2_X1 U14653 ( .A1(n11700), .A2(P1_EBX_REG_11__SCAN_IN), .ZN(n11654) );
  NAND2_X1 U14654 ( .A1(n11692), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11652) );
  OAI211_X1 U14655 ( .C1(n13276), .C2(P1_EBX_REG_11__SCAN_IN), .A(n11696), .B(
        n11652), .ZN(n11653) );
  NAND2_X1 U14656 ( .A1(n11654), .A2(n11653), .ZN(n14216) );
  MUX2_X1 U14657 ( .A(n11708), .B(n11696), .S(P1_EBX_REG_12__SCAN_IN), .Z(
        n11657) );
  NAND2_X1 U14658 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n13276), .ZN(
        n11655) );
  AND2_X1 U14659 ( .A1(n11686), .A2(n11655), .ZN(n11656) );
  NOR2_X2 U14660 ( .A1(n14219), .A2(n14206), .ZN(n14205) );
  OR2_X1 U14661 ( .A1(n11700), .A2(P1_EBX_REG_13__SCAN_IN), .ZN(n11660) );
  NAND2_X1 U14662 ( .A1(n11692), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n11658) );
  OAI211_X1 U14663 ( .C1(n13276), .C2(P1_EBX_REG_13__SCAN_IN), .A(n11696), .B(
        n11658), .ZN(n11659) );
  INV_X1 U14664 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n14199) );
  NAND2_X1 U14665 ( .A1(n11623), .A2(n14199), .ZN(n11663) );
  NAND2_X1 U14666 ( .A1(n11696), .A2(n14408), .ZN(n11661) );
  OAI211_X1 U14667 ( .C1(n13276), .C2(P1_EBX_REG_14__SCAN_IN), .A(n11661), .B(
        n11692), .ZN(n11662) );
  OR2_X1 U14668 ( .A1(n11700), .A2(P1_EBX_REG_15__SCAN_IN), .ZN(n11666) );
  NAND2_X1 U14669 ( .A1(n11692), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11664) );
  OAI211_X1 U14670 ( .C1(n13276), .C2(P1_EBX_REG_15__SCAN_IN), .A(n11629), .B(
        n11664), .ZN(n11665) );
  NAND2_X1 U14671 ( .A1(n11666), .A2(n11665), .ZN(n14090) );
  INV_X1 U14672 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n14195) );
  NAND2_X1 U14673 ( .A1(n11623), .A2(n14195), .ZN(n11670) );
  NAND2_X1 U14674 ( .A1(n11629), .A2(n11667), .ZN(n11668) );
  OAI211_X1 U14675 ( .C1(n13276), .C2(P1_EBX_REG_16__SCAN_IN), .A(n11668), .B(
        n11692), .ZN(n11669) );
  NAND2_X1 U14676 ( .A1(n11670), .A2(n11669), .ZN(n14079) );
  NAND2_X1 U14677 ( .A1(n14089), .A2(n14079), .ZN(n14081) );
  MUX2_X1 U14678 ( .A(n11700), .B(n11692), .S(P1_EBX_REG_17__SCAN_IN), .Z(
        n11672) );
  OR2_X1 U14679 ( .A1(n13560), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n11671) );
  NAND2_X1 U14680 ( .A1(n11672), .A2(n11671), .ZN(n14062) );
  INV_X1 U14681 ( .A(n11673), .ZN(n14061) );
  INV_X1 U14682 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n14191) );
  NAND2_X1 U14683 ( .A1(n11623), .A2(n14191), .ZN(n11676) );
  INV_X1 U14684 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n14369) );
  NAND2_X1 U14685 ( .A1(n11696), .A2(n14369), .ZN(n11674) );
  OAI211_X1 U14686 ( .C1(n13276), .C2(P1_EBX_REG_18__SCAN_IN), .A(n11674), .B(
        n11692), .ZN(n11675) );
  MUX2_X1 U14687 ( .A(n11700), .B(n11692), .S(P1_EBX_REG_19__SCAN_IN), .Z(
        n11678) );
  OR2_X1 U14688 ( .A1(n13560), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11677) );
  AND2_X2 U14689 ( .A1(n14187), .A2(n14186), .ZN(n14189) );
  MUX2_X1 U14690 ( .A(n11708), .B(n11629), .S(P1_EBX_REG_20__SCAN_IN), .Z(
        n11679) );
  OAI211_X1 U14691 ( .C1(n13696), .C2(n14379), .A(n11679), .B(n11686), .ZN(
        n14181) );
  OR2_X1 U14692 ( .A1(n11700), .A2(P1_EBX_REG_21__SCAN_IN), .ZN(n11682) );
  NAND2_X1 U14693 ( .A1(n11692), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11680) );
  OAI211_X1 U14694 ( .C1(n13276), .C2(P1_EBX_REG_21__SCAN_IN), .A(n11629), .B(
        n11680), .ZN(n11681) );
  NAND2_X1 U14695 ( .A1(n11682), .A2(n11681), .ZN(n14491) );
  MUX2_X1 U14696 ( .A(n11700), .B(n11692), .S(P1_EBX_REG_23__SCAN_IN), .Z(
        n11684) );
  OR2_X1 U14697 ( .A1(n13560), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11683) );
  AND2_X1 U14698 ( .A1(n11684), .A2(n11683), .ZN(n14171) );
  MUX2_X1 U14699 ( .A(n11708), .B(n11629), .S(P1_EBX_REG_22__SCAN_IN), .Z(
        n11688) );
  NAND2_X1 U14700 ( .A1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n13276), .ZN(
        n11685) );
  AND2_X1 U14701 ( .A1(n11686), .A2(n11685), .ZN(n11687) );
  NAND2_X1 U14702 ( .A1(n11688), .A2(n11687), .ZN(n14041) );
  INV_X1 U14703 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n14165) );
  NAND2_X1 U14704 ( .A1(n11623), .A2(n14165), .ZN(n11691) );
  INV_X1 U14705 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14331) );
  NAND2_X1 U14706 ( .A1(n11629), .A2(n14331), .ZN(n11689) );
  OAI211_X1 U14707 ( .C1(n13276), .C2(P1_EBX_REG_24__SCAN_IN), .A(n11689), .B(
        n11692), .ZN(n11690) );
  OR2_X1 U14708 ( .A1(n11700), .A2(P1_EBX_REG_25__SCAN_IN), .ZN(n11695) );
  NAND2_X1 U14709 ( .A1(n11692), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11693) );
  OAI211_X1 U14710 ( .C1(n13276), .C2(P1_EBX_REG_25__SCAN_IN), .A(n11696), .B(
        n11693), .ZN(n11694) );
  INV_X1 U14711 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n14159) );
  NAND2_X1 U14712 ( .A1(n11623), .A2(n14159), .ZN(n11699) );
  NAND2_X1 U14713 ( .A1(n11696), .A2(n14325), .ZN(n11697) );
  OAI211_X1 U14714 ( .C1(n13276), .C2(P1_EBX_REG_26__SCAN_IN), .A(n11697), .B(
        n11692), .ZN(n11698) );
  AND2_X1 U14715 ( .A1(n11699), .A2(n11698), .ZN(n14157) );
  MUX2_X1 U14716 ( .A(n11700), .B(n11692), .S(P1_EBX_REG_27__SCAN_IN), .Z(
        n11702) );
  OR2_X1 U14717 ( .A1(n13560), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11701) );
  NAND2_X1 U14718 ( .A1(n11702), .A2(n11701), .ZN(n14154) );
  INV_X1 U14719 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n15644) );
  NAND2_X1 U14720 ( .A1(n11623), .A2(n15644), .ZN(n11705) );
  INV_X1 U14721 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n13166) );
  NAND2_X1 U14722 ( .A1(n11629), .A2(n13166), .ZN(n11703) );
  OAI211_X1 U14723 ( .C1(n13276), .C2(P1_EBX_REG_28__SCAN_IN), .A(n11703), .B(
        n11692), .ZN(n11704) );
  NAND2_X1 U14724 ( .A1(n11705), .A2(n11704), .ZN(n14147) );
  OR2_X1 U14725 ( .A1(n13560), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11707) );
  INV_X1 U14726 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n14146) );
  NAND2_X1 U14727 ( .A1(n13696), .A2(n14146), .ZN(n11706) );
  NAND2_X1 U14728 ( .A1(n11707), .A2(n11706), .ZN(n11711) );
  OAI22_X1 U14729 ( .A1(n11711), .A2(n11709), .B1(P1_EBX_REG_29__SCAN_IN), 
        .B2(n11708), .ZN(n11769) );
  INV_X1 U14730 ( .A(n11710), .ZN(n11712) );
  AND2_X1 U14731 ( .A1(n13276), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11713) );
  AOI21_X1 U14732 ( .B1(n13560), .B2(P1_EBX_REG_30__SCAN_IN), .A(n11713), .ZN(
        n12291) );
  INV_X1 U14733 ( .A(n12291), .ZN(n11714) );
  XNOR2_X1 U14734 ( .A(n11715), .B(n11714), .ZN(n13994) );
  INV_X1 U14735 ( .A(n13994), .ZN(n11764) );
  OAI22_X1 U14736 ( .A1(n11610), .A2(n20127), .B1(n20113), .B2(n11716), .ZN(
        n11717) );
  NOR2_X1 U14737 ( .A1(n11719), .A2(n11718), .ZN(n13445) );
  INV_X1 U14738 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n20076) );
  OAI21_X1 U14739 ( .B1(n20076), .B2(n20075), .A(n20090), .ZN(n20051) );
  NOR2_X1 U14740 ( .A1(n20061), .A2(n20069), .ZN(n20054) );
  INV_X1 U14741 ( .A(n20054), .ZN(n15895) );
  NOR2_X1 U14742 ( .A1(n20974), .A2(n15895), .ZN(n15834) );
  NAND2_X1 U14743 ( .A1(n20051), .A2(n15834), .ZN(n15849) );
  INV_X1 U14744 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15868) );
  INV_X1 U14745 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n15898) );
  NOR3_X1 U14746 ( .A1(n11511), .A2(n15911), .A3(n15898), .ZN(n15876) );
  NAND3_X1 U14747 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(n15876), .ZN(n15852) );
  NOR2_X1 U14748 ( .A1(n15868), .A2(n15852), .ZN(n15855) );
  NAND2_X1 U14749 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n15855), .ZN(
        n11734) );
  NOR2_X1 U14750 ( .A1(n15849), .A2(n11734), .ZN(n11741) );
  NAND2_X1 U14751 ( .A1(n20053), .A2(n11741), .ZN(n11736) );
  OAI211_X1 U14752 ( .C1(n11722), .C2(n9796), .A(n11696), .B(n11721), .ZN(
        n11723) );
  INV_X1 U14753 ( .A(n11723), .ZN(n11729) );
  INV_X1 U14754 ( .A(n13545), .ZN(n11725) );
  NAND3_X1 U14755 ( .A1(n11726), .A2(n11725), .A3(n11724), .ZN(n11727) );
  NAND2_X1 U14756 ( .A1(n11727), .A2(n20113), .ZN(n11728) );
  AND4_X1 U14757 ( .A1(n11731), .A2(n11730), .A3(n11729), .A4(n11728), .ZN(
        n13443) );
  OAI211_X1 U14758 ( .C1(n13440), .C2(n9823), .A(n13443), .B(n11732), .ZN(
        n11733) );
  NOR2_X1 U14759 ( .A1(n20090), .A2(n20075), .ZN(n15871) );
  NAND2_X1 U14760 ( .A1(n15834), .A2(n15871), .ZN(n15851) );
  NOR2_X1 U14761 ( .A1(n11734), .A2(n15851), .ZN(n11743) );
  NAND3_X1 U14762 ( .A1(n13565), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A3(
        n11743), .ZN(n11735) );
  AND2_X1 U14763 ( .A1(n11598), .A2(n20113), .ZN(n13950) );
  INV_X1 U14764 ( .A(n14504), .ZN(n11737) );
  NAND2_X1 U14765 ( .A1(n11737), .A2(n11743), .ZN(n11738) );
  NAND2_X1 U14766 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n11739) );
  NAND3_X1 U14767 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15814) );
  NOR2_X1 U14768 ( .A1(n14369), .A2(n15814), .ZN(n11749) );
  NAND2_X1 U14769 ( .A1(n15816), .A2(n11749), .ZN(n15813) );
  AND2_X1 U14770 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15800) );
  NAND2_X1 U14771 ( .A1(n15803), .A2(n15800), .ZN(n14470) );
  NAND2_X1 U14772 ( .A1(n14438), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11740) );
  NOR2_X1 U14773 ( .A1(n14449), .A2(n11740), .ZN(n12297) );
  AOI21_X1 U14774 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n11741), .A(
        n20080), .ZN(n11748) );
  INV_X1 U14775 ( .A(n13565), .ZN(n11742) );
  AOI21_X1 U14776 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n11743), .A(
        n15872), .ZN(n11747) );
  NAND2_X1 U14777 ( .A1(n13565), .A2(n20076), .ZN(n11745) );
  OAI21_X1 U14778 ( .B1(n11744), .B2(n11746), .A(n11745), .ZN(n20072) );
  NOR3_X1 U14779 ( .A1(n11748), .A2(n11747), .A3(n20072), .ZN(n15848) );
  NAND2_X1 U14780 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n11749), .ZN(
        n14475) );
  NAND2_X1 U14781 ( .A1(n15897), .A2(n14475), .ZN(n11750) );
  NAND2_X1 U14782 ( .A1(n15848), .A2(n11750), .ZN(n15808) );
  AND3_X1 U14783 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n14478) );
  INV_X1 U14784 ( .A(n14478), .ZN(n11751) );
  OR2_X1 U14785 ( .A1(n15808), .A2(n11751), .ZN(n11752) );
  INV_X1 U14786 ( .A(n20072), .ZN(n15870) );
  NAND2_X1 U14787 ( .A1(n15870), .A2(n14519), .ZN(n15873) );
  NOR2_X1 U14788 ( .A1(n14519), .A2(n15800), .ZN(n11753) );
  NOR2_X1 U14789 ( .A1(n15798), .A2(n11753), .ZN(n14474) );
  INV_X1 U14790 ( .A(n11754), .ZN(n14458) );
  NAND2_X1 U14791 ( .A1(n15897), .A2(n14458), .ZN(n11755) );
  NAND2_X1 U14792 ( .A1(n14474), .A2(n11755), .ZN(n14467) );
  AND2_X1 U14793 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n11756) );
  NOR2_X1 U14794 ( .A1(n14519), .A2(n11756), .ZN(n11757) );
  NOR2_X1 U14795 ( .A1(n15798), .A2(n15897), .ZN(n12299) );
  NOR2_X1 U14796 ( .A1(n12299), .A2(n14438), .ZN(n11758) );
  NOR2_X1 U14797 ( .A1(n14452), .A2(n11758), .ZN(n11775) );
  OAI21_X1 U14798 ( .B1(n14519), .B2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n11759) );
  INV_X1 U14799 ( .A(n11759), .ZN(n11760) );
  NAND2_X1 U14800 ( .A1(n11775), .A2(n11760), .ZN(n12301) );
  OAI21_X1 U14801 ( .B1(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n12297), .A(
        n12301), .ZN(n11762) );
  INV_X1 U14802 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n13988) );
  NOR2_X1 U14803 ( .A1(n20081), .A2(n13988), .ZN(n14305) );
  INV_X1 U14804 ( .A(n14305), .ZN(n11761) );
  OAI21_X1 U14805 ( .B1(n14310), .B2(n15923), .A(n11765), .ZN(P1_U3001) );
  NOR2_X1 U14806 ( .A1(n11710), .A2(n11769), .ZN(n11770) );
  INV_X1 U14807 ( .A(n14145), .ZN(n11773) );
  INV_X1 U14808 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n20745) );
  NOR2_X1 U14809 ( .A1(n20081), .A2(n20745), .ZN(n14311) );
  INV_X1 U14810 ( .A(n14438), .ZN(n11771) );
  NOR3_X1 U14811 ( .A1(n14449), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n11771), .ZN(n11772) );
  AOI211_X1 U14812 ( .C1(n11773), .C2(n20063), .A(n14311), .B(n11772), .ZN(
        n11777) );
  OR2_X1 U14813 ( .A1(n11775), .A2(n11774), .ZN(n11776) );
  NOR3_X2 U14814 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(n16789), .ZN(n11779) );
  INV_X2 U14815 ( .A(n11779), .ZN(n17072) );
  AOI22_X1 U14816 ( .A1(n17101), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17049), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11780) );
  OAI21_X1 U14817 ( .B1(n15492), .B2(n21058), .A(n11780), .ZN(n11797) );
  INV_X1 U14818 ( .A(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n16986) );
  INV_X2 U14819 ( .A(n9848), .ZN(n17093) );
  AOI22_X1 U14820 ( .A1(n17092), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17093), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11795) );
  OR2_X2 U14821 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n15540), .ZN(
        n11811) );
  NAND2_X4 U14822 ( .A1(n11786), .A2(n18722), .ZN(n16933) );
  INV_X1 U14823 ( .A(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11785) );
  AOI22_X1 U14824 ( .A1(n17053), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17074), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11784) );
  OAI21_X1 U14825 ( .B1(n16933), .B2(n11785), .A(n11784), .ZN(n11793) );
  INV_X2 U14826 ( .A(n11832), .ZN(n11820) );
  INV_X2 U14827 ( .A(n16966), .ZN(n17036) );
  AOI22_X1 U14828 ( .A1(n15498), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11791) );
  INV_X2 U14829 ( .A(n11833), .ZN(n17051) );
  AOI22_X1 U14830 ( .A1(n17103), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n17100), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11790) );
  OAI211_X1 U14831 ( .C1(n16987), .C2(n20943), .A(n11791), .B(n11790), .ZN(
        n11792) );
  AOI211_X1 U14832 ( .C1(n16967), .C2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A(
        n11793), .B(n11792), .ZN(n11794) );
  OAI211_X1 U14833 ( .C1(n17114), .C2(n16986), .A(n11795), .B(n11794), .ZN(
        n11796) );
  INV_X1 U14834 ( .A(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n15514) );
  AOI22_X1 U14835 ( .A1(n17094), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17054), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11798) );
  OAI21_X1 U14836 ( .B1(n15492), .B2(n15514), .A(n11798), .ZN(n11809) );
  INV_X1 U14837 ( .A(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11807) );
  INV_X2 U14838 ( .A(n9848), .ZN(n17076) );
  AOI22_X1 U14839 ( .A1(n17076), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17100), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11806) );
  INV_X1 U14840 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17128) );
  INV_X2 U14841 ( .A(n16933), .ZN(n17077) );
  AOI22_X1 U14842 ( .A1(n17074), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17077), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11800) );
  OAI21_X1 U14843 ( .B1(n10222), .B2(n17128), .A(n11800), .ZN(n11804) );
  INV_X1 U14844 ( .A(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n21003) );
  AOI22_X1 U14845 ( .A1(n17002), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17070), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11802) );
  AOI22_X1 U14846 ( .A1(n17036), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17049), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11801) );
  OAI211_X1 U14847 ( .C1(n11811), .C2(n21003), .A(n11802), .B(n11801), .ZN(
        n11803) );
  AOI211_X1 U14848 ( .C1(n17110), .C2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A(
        n11804), .B(n11803), .ZN(n11805) );
  OAI211_X1 U14849 ( .C1(n17027), .C2(n11807), .A(n11806), .B(n11805), .ZN(
        n11808) );
  AOI22_X1 U14850 ( .A1(n17094), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11810) );
  OAI21_X1 U14851 ( .B1(n10222), .B2(n17137), .A(n11810), .ZN(n11817) );
  INV_X1 U14852 ( .A(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n15446) );
  AOI22_X1 U14853 ( .A1(n17053), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17074), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11816) );
  INV_X1 U14854 ( .A(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17033) );
  OAI22_X1 U14855 ( .A1(n16983), .A2(n16922), .B1(n16987), .B2(n17033), .ZN(
        n11815) );
  AOI22_X1 U14856 ( .A1(n17095), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17093), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11814) );
  AOI22_X1 U14857 ( .A1(n15498), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17100), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11813) );
  AOI22_X1 U14858 ( .A1(n16967), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17077), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11812) );
  INV_X1 U14859 ( .A(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n16934) );
  AOI22_X1 U14860 ( .A1(n17074), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17100), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11829) );
  AOI22_X1 U14861 ( .A1(n11781), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17095), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11819) );
  AOI22_X1 U14862 ( .A1(n17101), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17103), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11818) );
  OAI211_X1 U14863 ( .C1(n16987), .C2(n17052), .A(n11819), .B(n11818), .ZN(
        n11827) );
  AOI22_X1 U14864 ( .A1(n17070), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17093), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11825) );
  INV_X2 U14865 ( .A(n16966), .ZN(n17102) );
  AOI22_X1 U14866 ( .A1(n17083), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17102), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11824) );
  AOI22_X1 U14867 ( .A1(n17092), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11779), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11823) );
  NAND2_X1 U14868 ( .A1(n16967), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n11822) );
  NAND4_X1 U14869 ( .A1(n11825), .A2(n11824), .A3(n11823), .A4(n11822), .ZN(
        n11826) );
  AOI211_X1 U14870 ( .C1(n17077), .C2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A(
        n11827), .B(n11826), .ZN(n11828) );
  INV_X1 U14871 ( .A(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n16955) );
  AOI22_X1 U14872 ( .A1(n17092), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n16967), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11830) );
  OAI21_X1 U14873 ( .B1(n16955), .B2(n17072), .A(n11830), .ZN(n11831) );
  INV_X1 U14874 ( .A(n11831), .ZN(n11841) );
  INV_X1 U14875 ( .A(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n17073) );
  AOI22_X1 U14876 ( .A1(n11781), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_13__1__SCAN_IN), .B2(n11832), .ZN(n11835) );
  AOI22_X1 U14877 ( .A1(n17096), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_12__1__SCAN_IN), .B2(n11833), .ZN(n11834) );
  OAI211_X1 U14878 ( .C1(n16933), .C2(n17073), .A(n11835), .B(n11834), .ZN(
        n11836) );
  AOI22_X1 U14879 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n17074), .B1(
        P3_INSTQUEUE_REG_9__1__SCAN_IN), .B2(n17076), .ZN(n11839) );
  INV_X1 U14880 ( .A(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n17086) );
  INV_X1 U14881 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17145) );
  AOI22_X1 U14882 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n17054), .B1(
        P3_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n17102), .ZN(n11842) );
  OAI21_X1 U14883 ( .B1(n10222), .B2(n17145), .A(n11842), .ZN(n11844) );
  NAND2_X2 U14884 ( .A1(n10226), .A2(n10224), .ZN(n17299) );
  NAND2_X1 U14885 ( .A1(n17293), .A2(n17299), .ZN(n11868) );
  AOI22_X1 U14886 ( .A1(n17092), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17102), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11855) );
  INV_X1 U14887 ( .A(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11847) );
  AOI22_X1 U14888 ( .A1(n17049), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17093), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11846) );
  AOI22_X1 U14889 ( .A1(n17053), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17095), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11845) );
  OAI211_X1 U14890 ( .C1(n16987), .C2(n11847), .A(n11846), .B(n11845), .ZN(
        n11853) );
  AOI22_X1 U14891 ( .A1(n17103), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n17100), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11851) );
  AOI22_X1 U14892 ( .A1(n17094), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17054), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11850) );
  AOI22_X1 U14893 ( .A1(n17002), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17074), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11849) );
  NAND2_X1 U14894 ( .A1(n16967), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n11848) );
  NAND4_X1 U14895 ( .A1(n11851), .A2(n11850), .A3(n11849), .A4(n11848), .ZN(
        n11852) );
  AOI211_X1 U14896 ( .C1(n17077), .C2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A(
        n11853), .B(n11852), .ZN(n11854) );
  OAI211_X1 U14897 ( .C1(n11820), .C2(n20935), .A(n11855), .B(n11854), .ZN(
        n12064) );
  NAND2_X1 U14898 ( .A1(n11888), .A2(n12064), .ZN(n11891) );
  NOR2_X1 U14899 ( .A1(n17281), .A2(n11891), .ZN(n11896) );
  AOI22_X1 U14900 ( .A1(n17074), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17100), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11866) );
  INV_X1 U14901 ( .A(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11858) );
  AOI22_X1 U14902 ( .A1(n17053), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17095), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11857) );
  AOI22_X1 U14903 ( .A1(n17070), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11856) );
  OAI211_X1 U14904 ( .C1(n16987), .C2(n11858), .A(n11857), .B(n11856), .ZN(
        n11864) );
  AOI22_X1 U14905 ( .A1(n17002), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17083), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11862) );
  AOI22_X1 U14906 ( .A1(n17049), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17093), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11861) );
  AOI22_X1 U14907 ( .A1(n17092), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17054), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11860) );
  NAND2_X1 U14908 ( .A1(n16967), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n11859) );
  NAND4_X1 U14909 ( .A1(n11862), .A2(n11861), .A3(n11860), .A4(n11859), .ZN(
        n11863) );
  AOI211_X1 U14910 ( .C1(n17077), .C2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A(
        n11864), .B(n11863), .ZN(n11865) );
  OAI211_X1 U14911 ( .C1(n10222), .C2(n17126), .A(n11866), .B(n11865), .ZN(
        n12059) );
  NAND2_X1 U14912 ( .A1(n11896), .A2(n12059), .ZN(n11867) );
  INV_X1 U14913 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16272) );
  INV_X1 U14914 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17810) );
  AOI21_X1 U14915 ( .B1(n17274), .B2(n11867), .A(n17694), .ZN(n11899) );
  NAND2_X1 U14916 ( .A1(n12058), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n11880) );
  OAI22_X1 U14917 ( .A1(n16987), .A2(n16969), .B1(n9848), .B2(n18333), .ZN(
        n11873) );
  AOI22_X1 U14918 ( .A1(n17094), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17054), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11871) );
  AOI22_X1 U14919 ( .A1(n17096), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17103), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11870) );
  AOI22_X1 U14920 ( .A1(n16967), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17077), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11869) );
  NAND3_X1 U14921 ( .A1(n11871), .A2(n11870), .A3(n11869), .ZN(n11872) );
  AOI211_X1 U14922 ( .C1(n17092), .C2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A(
        n11873), .B(n11872), .ZN(n11879) );
  AOI22_X1 U14923 ( .A1(n17074), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11779), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11875) );
  AOI22_X1 U14924 ( .A1(n17036), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17100), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11876) );
  OAI21_X1 U14925 ( .B1(n11820), .B2(n21054), .A(n11876), .ZN(n11877) );
  INV_X1 U14926 ( .A(n11877), .ZN(n11878) );
  INV_X1 U14927 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18742) );
  INV_X1 U14928 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18727) );
  XOR2_X1 U14929 ( .A(n18727), .B(n17299), .Z(n17771) );
  NAND2_X1 U14930 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n11882), .ZN(
        n11883) );
  NAND2_X1 U14931 ( .A1(n11884), .A2(n11885), .ZN(n11887) );
  NAND2_X1 U14932 ( .A1(n11887), .A2(n17748), .ZN(n17741) );
  INV_X1 U14933 ( .A(n12064), .ZN(n17285) );
  XNOR2_X1 U14934 ( .A(n17285), .B(n11888), .ZN(n11889) );
  XOR2_X1 U14935 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B(n11889), .Z(
        n17742) );
  NAND2_X1 U14936 ( .A1(n17741), .A2(n17742), .ZN(n17740) );
  NAND2_X1 U14937 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n11889), .ZN(
        n11890) );
  XOR2_X1 U14938 ( .A(n17281), .B(n11891), .Z(n11894) );
  INV_X1 U14939 ( .A(n11894), .ZN(n11892) );
  NAND2_X1 U14940 ( .A1(n11894), .A2(n11893), .ZN(n11895) );
  INV_X1 U14941 ( .A(n12059), .ZN(n17278) );
  XNOR2_X1 U14942 ( .A(n17278), .B(n11896), .ZN(n11897) );
  XOR2_X1 U14943 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n11897), .Z(
        n17714) );
  NAND2_X1 U14944 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n11897), .ZN(
        n11898) );
  NAND2_X1 U14945 ( .A1(n11899), .A2(n11901), .ZN(n11902) );
  INV_X1 U14946 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n20862) );
  INV_X1 U14947 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17986) );
  NOR2_X1 U14948 ( .A1(n18001), .A2(n17986), .ZN(n17651) );
  INV_X1 U14949 ( .A(n17651), .ZN(n17978) );
  INV_X1 U14950 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17645) );
  NOR2_X1 U14951 ( .A1(n17978), .A2(n17645), .ZN(n17966) );
  NAND2_X1 U14952 ( .A1(n17966), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n17607) );
  INV_X1 U14953 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17938) );
  NOR2_X1 U14954 ( .A1(n17607), .A2(n17938), .ZN(n17934) );
  NAND2_X1 U14955 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n17934), .ZN(
        n17910) );
  INV_X1 U14956 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n17932) );
  INV_X1 U14957 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n17912) );
  INV_X1 U14958 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n20946) );
  INV_X1 U14959 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n17962) );
  NAND4_X1 U14960 ( .A1(n20946), .A2(n17962), .A3(n17938), .A4(n17932), .ZN(
        n11904) );
  INV_X1 U14961 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17893) );
  NOR2_X1 U14962 ( .A1(n17912), .A2(n17893), .ZN(n17555) );
  NAND2_X1 U14963 ( .A1(n11905), .A2(n17467), .ZN(n17576) );
  NAND2_X1 U14964 ( .A1(n17555), .A2(n17576), .ZN(n17519) );
  INV_X1 U14965 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17832) );
  INV_X1 U14966 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n17553) );
  INV_X1 U14967 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17541) );
  NOR2_X1 U14968 ( .A1(n17553), .A2(n17541), .ZN(n17865) );
  NAND2_X1 U14969 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17865), .ZN(
        n17505) );
  INV_X1 U14970 ( .A(n17505), .ZN(n17856) );
  NAND2_X1 U14971 ( .A1(n17856), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n17482) );
  NOR2_X1 U14972 ( .A1(n17832), .A2(n17482), .ZN(n17471) );
  NAND2_X1 U14973 ( .A1(n17555), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n17812) );
  INV_X1 U14974 ( .A(n17812), .ZN(n17863) );
  NAND2_X1 U14975 ( .A1(n17863), .A2(n17856), .ZN(n17845) );
  INV_X1 U14976 ( .A(n17845), .ZN(n17851) );
  NAND2_X1 U14977 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17851), .ZN(
        n17854) );
  NOR2_X1 U14978 ( .A1(n17832), .A2(n17854), .ZN(n17827) );
  NOR2_X1 U14979 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17694), .ZN(
        n17561) );
  NAND2_X1 U14980 ( .A1(n17561), .A2(n17553), .ZN(n11906) );
  NOR2_X1 U14981 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n11906), .ZN(
        n17521) );
  INV_X1 U14982 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n17525) );
  NAND2_X1 U14983 ( .A1(n17521), .A2(n17525), .ZN(n17502) );
  NOR3_X1 U14984 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(n17502), .ZN(n11907) );
  NOR2_X2 U14985 ( .A1(n17476), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n17475) );
  NOR2_X1 U14986 ( .A1(n11910), .A2(n17475), .ZN(n17454) );
  OR2_X1 U14987 ( .A1(n17694), .A2(n17475), .ZN(n17453) );
  OAI221_X1 U14988 ( .B1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n17628), 
        .C1(n17810), .C2(n17454), .A(n17453), .ZN(n17443) );
  NOR2_X1 U14989 ( .A1(n17454), .A2(n17628), .ZN(n11911) );
  NAND2_X1 U14990 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17788) );
  NOR2_X2 U14991 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n11913), .ZN(
        n16309) );
  NOR2_X1 U14992 ( .A1(n17694), .A2(n11920), .ZN(n11921) );
  INV_X1 U14993 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n17800) );
  INV_X1 U14994 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16298) );
  NOR2_X1 U14995 ( .A1(n17800), .A2(n16298), .ZN(n16270) );
  NAND2_X1 U14996 ( .A1(n16270), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16284) );
  INV_X1 U14997 ( .A(n16284), .ZN(n15623) );
  NAND2_X1 U14998 ( .A1(n15623), .A2(n16299), .ZN(n11918) );
  INV_X1 U14999 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18728) );
  NAND2_X1 U15000 ( .A1(n18728), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11914) );
  NAND2_X1 U15001 ( .A1(n11918), .A2(n11914), .ZN(n11916) );
  NOR2_X1 U15002 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n18728), .ZN(
        n16292) );
  INV_X1 U15003 ( .A(n16292), .ZN(n11915) );
  AOI22_X1 U15004 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n17694), .B1(
        n17628), .B2(n18728), .ZN(n11923) );
  INV_X1 U15005 ( .A(n11918), .ZN(n11919) );
  INV_X1 U15006 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n20896) );
  NOR2_X1 U15007 ( .A1(n15625), .A2(n20896), .ZN(n15624) );
  OAI21_X1 U15008 ( .B1(n11921), .B2(n15624), .A(n11923), .ZN(n11922) );
  OAI21_X1 U15009 ( .B1(n11924), .B2(n11923), .A(n11922), .ZN(n16293) );
  NAND2_X1 U15010 ( .A1(n18169), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12039) );
  OAI21_X1 U15011 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n18169), .A(
        n12039), .ZN(n12042) );
  NOR2_X1 U15012 ( .A1(n12042), .A2(n12038), .ZN(n11937) );
  OAI22_X1 U15013 ( .A1(n18732), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(
        n18599), .B2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11933) );
  OAI22_X1 U15014 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n11927), .B1(
        P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n20878), .ZN(n11929) );
  NOR2_X1 U15015 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n20878), .ZN(
        n11928) );
  NAND2_X1 U15016 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n11927), .ZN(
        n11930) );
  AOI22_X1 U15017 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n11929), .B1(
        n11928), .B2(n11930), .ZN(n11936) );
  AOI21_X1 U15018 ( .B1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n11930), .A(
        n11929), .ZN(n11931) );
  NAND2_X1 U15019 ( .A1(n11934), .A2(n11933), .ZN(n11932) );
  OAI211_X1 U15020 ( .C1(n11934), .C2(n11933), .A(n11936), .B(n11932), .ZN(
        n12043) );
  NAND2_X1 U15021 ( .A1(n12040), .A2(n12043), .ZN(n11935) );
  INV_X1 U15022 ( .A(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n18336) );
  AOI22_X1 U15023 ( .A1(n17036), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n17049), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11939) );
  AOI22_X1 U15024 ( .A1(n17076), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n15497), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11938) );
  OAI211_X1 U15025 ( .C1(n16987), .C2(n18336), .A(n11939), .B(n11938), .ZN(
        n11948) );
  AOI22_X1 U15026 ( .A1(n17095), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n17083), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11946) );
  AOI22_X1 U15027 ( .A1(n17053), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17065), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11945) );
  INV_X2 U15028 ( .A(n16983), .ZN(n17054) );
  AOI22_X1 U15029 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n17092), .B1(
        n17054), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11940) );
  INV_X1 U15030 ( .A(n11940), .ZN(n11943) );
  INV_X1 U15031 ( .A(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n17075) );
  AOI22_X1 U15032 ( .A1(n16967), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n17074), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11941) );
  OAI21_X1 U15033 ( .B1(n10222), .B2(n17075), .A(n11941), .ZN(n11942) );
  AOI211_X1 U15034 ( .C1(n17070), .C2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A(
        n11943), .B(n11942), .ZN(n11944) );
  NAND3_X1 U15035 ( .A1(n11946), .A2(n11945), .A3(n11944), .ZN(n11947) );
  AOI211_X4 U15036 ( .C1(n17077), .C2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A(
        n11948), .B(n11947), .ZN(n18117) );
  INV_X1 U15037 ( .A(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n16968) );
  AOI22_X1 U15038 ( .A1(n17103), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17076), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11949) );
  OAI21_X1 U15039 ( .B1(n9847), .B2(n16968), .A(n11949), .ZN(n11958) );
  AOI22_X1 U15040 ( .A1(n17095), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17054), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11956) );
  OAI22_X1 U15041 ( .A1(n11799), .A2(n16965), .B1(n16987), .B2(n18333), .ZN(
        n11954) );
  AOI22_X1 U15042 ( .A1(n15498), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11779), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11952) );
  AOI22_X1 U15043 ( .A1(n17036), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n15497), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11951) );
  AOI22_X1 U15044 ( .A1(n16967), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17077), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11950) );
  NAND3_X1 U15045 ( .A1(n11952), .A2(n11951), .A3(n11950), .ZN(n11953) );
  AOI211_X1 U15046 ( .C1(n17053), .C2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A(
        n11954), .B(n11953), .ZN(n11955) );
  OAI211_X1 U15047 ( .C1(n17027), .C2(n21054), .A(n11956), .B(n11955), .ZN(
        n11957) );
  NOR2_X1 U15048 ( .A1(n18760), .A2(n18114), .ZN(n12023) );
  OR2_X1 U15049 ( .A1(n12026), .A2(n12023), .ZN(n18779) );
  INV_X1 U15050 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n16991) );
  AOI22_X1 U15051 ( .A1(n15498), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n15497), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11959) );
  OAI21_X1 U15052 ( .B1(n17072), .B2(n16991), .A(n11959), .ZN(n11968) );
  INV_X1 U15053 ( .A(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n15477) );
  AOI22_X1 U15054 ( .A1(n17092), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n17077), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11966) );
  OAI22_X1 U15055 ( .A1(n17114), .A2(n20943), .B1(n11799), .B2(n21058), .ZN(
        n11964) );
  AOI22_X1 U15056 ( .A1(n17096), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11962) );
  AOI22_X1 U15057 ( .A1(n17101), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17103), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11961) );
  AOI22_X1 U15058 ( .A1(n16967), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17110), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11960) );
  NAND3_X1 U15059 ( .A1(n11962), .A2(n11961), .A3(n11960), .ZN(n11963) );
  AOI211_X1 U15060 ( .C1(n17093), .C2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A(
        n11964), .B(n11963), .ZN(n11965) );
  OAI211_X1 U15061 ( .C1(n15492), .C2(n15477), .A(n11966), .B(n11965), .ZN(
        n11967) );
  AOI211_X4 U15062 ( .C1(n17083), .C2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A(
        n11968), .B(n11967), .ZN(n18145) );
  AOI22_X1 U15063 ( .A1(n17083), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17103), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11969) );
  OAI21_X1 U15064 ( .B1(n15492), .B2(n16922), .A(n11969), .ZN(n11978) );
  INV_X1 U15065 ( .A(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n18342) );
  AOI22_X1 U15066 ( .A1(n17074), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11976) );
  OAI22_X1 U15067 ( .A1(n17072), .A2(n17137), .B1(n9848), .B2(n17034), .ZN(
        n11974) );
  AOI22_X1 U15068 ( .A1(n15498), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17054), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11972) );
  INV_X2 U15069 ( .A(n17114), .ZN(n17002) );
  AOI22_X1 U15070 ( .A1(n17002), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n15497), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11971) );
  AOI22_X1 U15071 ( .A1(n16967), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17077), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11970) );
  NAND3_X1 U15072 ( .A1(n11972), .A2(n11971), .A3(n11970), .ZN(n11973) );
  AOI211_X1 U15073 ( .C1(n17092), .C2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A(
        n11974), .B(n11973), .ZN(n11975) );
  OAI211_X1 U15074 ( .C1(n16987), .C2(n18342), .A(n11976), .B(n11975), .ZN(
        n11977) );
  AOI22_X1 U15075 ( .A1(n17095), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n15497), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11979) );
  OAI21_X1 U15076 ( .B1(n11820), .B2(n16894), .A(n11979), .ZN(n11988) );
  INV_X1 U15077 ( .A(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n15519) );
  AOI22_X1 U15078 ( .A1(n17074), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17076), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11986) );
  INV_X1 U15079 ( .A(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n15516) );
  AOI22_X1 U15080 ( .A1(n17083), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17092), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11980) );
  OAI21_X1 U15081 ( .B1(n16933), .B2(n15516), .A(n11980), .ZN(n11984) );
  INV_X1 U15082 ( .A(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n15433) );
  AOI22_X1 U15083 ( .A1(n17096), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17103), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11982) );
  AOI22_X1 U15084 ( .A1(n17036), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11779), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11981) );
  OAI211_X1 U15085 ( .C1(n16987), .C2(n15433), .A(n11982), .B(n11981), .ZN(
        n11983) );
  AOI211_X1 U15086 ( .C1(n16967), .C2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A(
        n11984), .B(n11983), .ZN(n11985) );
  OAI211_X1 U15087 ( .C1(n16983), .C2(n15519), .A(n11986), .B(n11985), .ZN(
        n11987) );
  AOI211_X4 U15088 ( .C1(n17065), .C2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A(
        n11988), .B(n11987), .ZN(n18135) );
  AOI22_X1 U15089 ( .A1(n17074), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17102), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11998) );
  INV_X1 U15090 ( .A(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17062) );
  AOI22_X1 U15091 ( .A1(n17049), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17093), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11990) );
  AOI22_X1 U15092 ( .A1(n17083), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17103), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11989) );
  OAI211_X1 U15093 ( .C1(n16933), .C2(n17062), .A(n11990), .B(n11989), .ZN(
        n11996) );
  AOI22_X1 U15094 ( .A1(n17053), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17095), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11994) );
  AOI22_X1 U15095 ( .A1(n15498), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n15497), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11993) );
  AOI22_X1 U15096 ( .A1(n17092), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17054), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11992) );
  NAND2_X1 U15097 ( .A1(n17110), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n11991) );
  NAND4_X1 U15098 ( .A1(n11994), .A2(n11993), .A3(n11992), .A4(n11991), .ZN(
        n11995) );
  OAI211_X1 U15099 ( .C1(n17114), .C2(n17052), .A(n11998), .B(n11997), .ZN(
        n15552) );
  AOI22_X1 U15100 ( .A1(n17002), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17103), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11999) );
  OAI21_X1 U15101 ( .B1(n17072), .B2(n17133), .A(n11999), .ZN(n12008) );
  AOI22_X1 U15102 ( .A1(n15498), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17102), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12006) );
  INV_X1 U15103 ( .A(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17018) );
  AOI22_X1 U15104 ( .A1(n17074), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n15497), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12000) );
  OAI21_X1 U15105 ( .B1(n16933), .B2(n17018), .A(n12000), .ZN(n12004) );
  INV_X1 U15106 ( .A(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n15509) );
  AOI22_X1 U15107 ( .A1(n17083), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17054), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12002) );
  AOI22_X1 U15108 ( .A1(n17095), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17076), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12001) );
  OAI211_X1 U15109 ( .C1(n16987), .C2(n15509), .A(n12002), .B(n12001), .ZN(
        n12003) );
  AOI211_X1 U15110 ( .C1(n16967), .C2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A(
        n12004), .B(n12003), .ZN(n12005) );
  OAI211_X1 U15111 ( .C1(n17027), .C2(n20935), .A(n12006), .B(n12005), .ZN(
        n12007) );
  AOI22_X1 U15112 ( .A1(n17092), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17103), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12018) );
  INV_X1 U15113 ( .A(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17013) );
  AOI22_X1 U15114 ( .A1(n17002), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12010) );
  AOI22_X1 U15115 ( .A1(n17083), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n15497), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12009) );
  OAI211_X1 U15116 ( .C1(n16933), .C2(n17013), .A(n12010), .B(n12009), .ZN(
        n12016) );
  AOI22_X1 U15117 ( .A1(n17053), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17054), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12014) );
  AOI22_X1 U15118 ( .A1(n17095), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17070), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12013) );
  AOI22_X1 U15119 ( .A1(n17074), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17093), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12012) );
  NAND2_X1 U15120 ( .A1(n17110), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n12011) );
  NAND4_X1 U15121 ( .A1(n12014), .A2(n12013), .A3(n12012), .A4(n12011), .ZN(
        n12015) );
  OAI211_X1 U15122 ( .C1(n17072), .C2(n17126), .A(n12018), .B(n12017), .ZN(
        n17156) );
  NOR2_X1 U15123 ( .A1(n18130), .A2(n17156), .ZN(n18571) );
  NAND3_X1 U15124 ( .A1(n12019), .A2(n15555), .A3(n18571), .ZN(n15427) );
  NOR2_X2 U15125 ( .A1(n12034), .A2(n15552), .ZN(n18570) );
  INV_X1 U15126 ( .A(n17156), .ZN(n18140) );
  NAND2_X1 U15127 ( .A1(n18570), .A2(n12045), .ZN(n15429) );
  NOR2_X2 U15128 ( .A1(n17308), .A2(n18145), .ZN(n12021) );
  INV_X1 U15129 ( .A(n12021), .ZN(n12025) );
  NAND2_X1 U15130 ( .A1(n12020), .A2(n17156), .ZN(n12027) );
  NOR4_X2 U15131 ( .A1(n12034), .A2(n15550), .A3(n12025), .A4(n12027), .ZN(
        n12035) );
  NAND2_X1 U15132 ( .A1(n12035), .A2(n15552), .ZN(n15531) );
  NAND2_X1 U15133 ( .A1(n17346), .A2(n15531), .ZN(n16416) );
  NOR2_X1 U15134 ( .A1(n17156), .A2(n18135), .ZN(n18588) );
  NAND2_X1 U15135 ( .A1(n17291), .A2(n15639), .ZN(n15638) );
  NAND2_X1 U15136 ( .A1(n12023), .A2(n15638), .ZN(n15534) );
  OAI21_X1 U15137 ( .B1(n15555), .B2(n12024), .A(n15534), .ZN(n12033) );
  NOR2_X1 U15138 ( .A1(n15552), .A2(n12027), .ZN(n15551) );
  NOR2_X1 U15139 ( .A1(n12024), .A2(n15551), .ZN(n12032) );
  AOI22_X1 U15140 ( .A1(n9817), .A2(n12025), .B1(n18130), .B2(n18588), .ZN(
        n12031) );
  NAND2_X1 U15141 ( .A1(n17291), .A2(n12027), .ZN(n12029) );
  NOR2_X1 U15142 ( .A1(n15552), .A2(n12026), .ZN(n12047) );
  INV_X1 U15143 ( .A(n12047), .ZN(n12028) );
  AOI22_X1 U15144 ( .A1(n12029), .A2(n15550), .B1(n12028), .B2(n12027), .ZN(
        n12030) );
  OAI211_X1 U15145 ( .C1(n12032), .C2(n17308), .A(n12031), .B(n12030), .ZN(
        n15532) );
  AOI21_X1 U15146 ( .B1(n12034), .B2(n12033), .A(n15532), .ZN(n12036) );
  NAND2_X1 U15147 ( .A1(n12035), .A2(n12036), .ZN(n15530) );
  NAND2_X1 U15148 ( .A1(n18562), .A2(n15530), .ZN(n17847) );
  NAND3_X1 U15149 ( .A1(n12044), .A2(n15528), .A3(n18760), .ZN(n12037) );
  NAND2_X1 U15150 ( .A1(n12037), .A2(n12036), .ZN(n18569) );
  XNOR2_X1 U15151 ( .A(n12039), .B(n12038), .ZN(n12041) );
  NOR2_X1 U15152 ( .A1(n12043), .A2(n12042), .ZN(n15557) );
  NOR2_X1 U15153 ( .A1(n15527), .A2(n15557), .ZN(n18556) );
  NOR2_X1 U15154 ( .A1(n18117), .A2(n15552), .ZN(n15554) );
  NAND2_X1 U15155 ( .A1(n15554), .A2(n17156), .ZN(n15556) );
  AOI211_X1 U15156 ( .C1(n15550), .C2(n15639), .A(n12045), .B(n12044), .ZN(
        n12046) );
  NAND2_X1 U15157 ( .A1(n12047), .A2(n12046), .ZN(n15533) );
  INV_X1 U15158 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n18764) );
  INV_X1 U15159 ( .A(n18611), .ZN(n18619) );
  NAND2_X1 U15160 ( .A1(n16293), .A2(n17695), .ZN(n12090) );
  NAND2_X1 U15161 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n18099) );
  NAND2_X1 U15162 ( .A1(n18716), .A2(n18099), .ZN(n18766) );
  INV_X1 U15163 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n18621) );
  NOR2_X1 U15164 ( .A1(n18726), .A2(n18621), .ZN(n17735) );
  INV_X1 U15165 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n16454) );
  NAND3_X1 U15166 ( .A1(n17685), .A2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n16667) );
  INV_X1 U15167 ( .A(n16667), .ZN(n12049) );
  NAND2_X1 U15168 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16632) );
  NAND2_X1 U15169 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17581) );
  NAND2_X1 U15170 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17546) );
  NAND2_X1 U15171 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17510) );
  INV_X1 U15172 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17473) );
  INV_X1 U15173 ( .A(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17462) );
  NOR2_X1 U15174 ( .A1(n17473), .A2(n17462), .ZN(n17456) );
  INV_X1 U15175 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17447) );
  INV_X1 U15176 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n16278) );
  XOR2_X2 U15177 ( .A(n16454), .B(n12050), .Z(n16790) );
  INV_X1 U15178 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n18704) );
  NOR2_X1 U15179 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18776) );
  NOR2_X1 U15180 ( .A1(n18704), .A2(n18091), .ZN(n16290) );
  NAND2_X1 U15181 ( .A1(n17456), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17420) );
  NOR2_X1 U15182 ( .A1(n17457), .A2(n17420), .ZN(n17414) );
  NAND3_X1 U15183 ( .A1(n17414), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n16266) );
  NOR2_X1 U15184 ( .A1(n16278), .A2(n16266), .ZN(n12052) );
  NAND2_X1 U15185 ( .A1(n18764), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n17781) );
  NOR2_X1 U15186 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18609) );
  INV_X1 U15187 ( .A(n18609), .ZN(n18763) );
  AOI21_X1 U15188 ( .B1(n18099), .B2(n18763), .A(n18740), .ZN(n12051) );
  INV_X1 U15189 ( .A(n12051), .ZN(n18112) );
  NAND3_X1 U15190 ( .A1(n18775), .A2(n18716), .A3(P3_STATEBS16_REG_SCAN_IN), 
        .ZN(n18456) );
  AOI21_X1 U15191 ( .B1(n17532), .B2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n18497), .ZN(n17580) );
  INV_X1 U15192 ( .A(n17580), .ZN(n17632) );
  NAND2_X1 U15193 ( .A1(n12052), .A2(n17632), .ZN(n16257) );
  XNOR2_X1 U15194 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(
        P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n12055) );
  NOR2_X1 U15195 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n17500), .ZN(
        n16279) );
  INV_X1 U15196 ( .A(n16439), .ZN(n12054) );
  OR2_X1 U15197 ( .A1(n18428), .A2(n12052), .ZN(n12053) );
  OAI211_X1 U15198 ( .C1(n12054), .C2(n17781), .A(n12053), .B(n17780), .ZN(
        n16269) );
  NOR2_X1 U15199 ( .A1(n16279), .A2(n16269), .ZN(n16256) );
  OAI22_X1 U15200 ( .A1(n16257), .A2(n12055), .B1(n16256), .B2(n16454), .ZN(
        n12056) );
  AOI211_X1 U15201 ( .C1(n17638), .C2(n16790), .A(n16290), .B(n12056), .ZN(
        n12089) );
  NAND2_X1 U15202 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17471), .ZN(
        n17811) );
  NOR2_X1 U15203 ( .A1(n17811), .A2(n17788), .ZN(n15569) );
  NAND2_X1 U15204 ( .A1(n17863), .A2(n15569), .ZN(n16254) );
  NOR2_X1 U15205 ( .A1(n16254), .A2(n17467), .ZN(n17427) );
  INV_X1 U15206 ( .A(n17427), .ZN(n17793) );
  NOR2_X1 U15207 ( .A1(n16284), .A2(n17793), .ZN(n16260) );
  NAND2_X1 U15208 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16260), .ZN(
        n12057) );
  XOR2_X1 U15209 ( .A(n18728), .B(n12057), .Z(n16294) );
  NOR2_X2 U15210 ( .A1(n15567), .A2(n17784), .ZN(n17696) );
  NAND2_X1 U15211 ( .A1(n16294), .A2(n17696), .ZN(n12088) );
  INV_X1 U15212 ( .A(n15568), .ZN(n17895) );
  NOR2_X1 U15213 ( .A1(n10241), .A2(n12058), .ZN(n12068) );
  NOR2_X1 U15214 ( .A1(n12068), .A2(n17293), .ZN(n12066) );
  NOR2_X1 U15215 ( .A1(n12066), .A2(n17288), .ZN(n12065) );
  NAND2_X1 U15216 ( .A1(n12065), .A2(n12064), .ZN(n12062) );
  NOR2_X1 U15217 ( .A1(n17281), .A2(n12062), .ZN(n12061) );
  NAND2_X1 U15218 ( .A1(n12061), .A2(n12059), .ZN(n12060) );
  NOR2_X1 U15219 ( .A1(n17274), .A2(n12060), .ZN(n12083) );
  XOR2_X1 U15220 ( .A(n12060), .B(n17274), .Z(n17706) );
  XNOR2_X1 U15221 ( .A(n12061), .B(n17278), .ZN(n12076) );
  XOR2_X1 U15222 ( .A(n12062), .B(n17281), .Z(n12063) );
  NAND2_X1 U15223 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n12063), .ZN(
        n12075) );
  XOR2_X1 U15224 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B(n12063), .Z(
        n17725) );
  INV_X1 U15225 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n18004) );
  XOR2_X1 U15226 ( .A(n12065), .B(n12064), .Z(n17737) );
  XOR2_X1 U15227 ( .A(n12066), .B(n17288), .Z(n12067) );
  NAND2_X1 U15228 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n12067), .ZN(
        n12073) );
  XOR2_X1 U15229 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n12067), .Z(
        n17752) );
  XNOR2_X1 U15230 ( .A(n17293), .B(n12068), .ZN(n12069) );
  NAND2_X1 U15231 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n12069), .ZN(
        n12072) );
  XOR2_X1 U15232 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n12069), .Z(
        n17760) );
  INV_X1 U15233 ( .A(n10241), .ZN(n15640) );
  AOI21_X1 U15234 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n17299), .A(
        n15640), .ZN(n12071) );
  NOR2_X1 U15235 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n17299), .ZN(
        n12070) );
  AOI221_X1 U15236 ( .B1(n15640), .B2(n17299), .C1(n12071), .C2(n18742), .A(
        n12070), .ZN(n17759) );
  NAND2_X1 U15237 ( .A1(n17760), .A2(n17759), .ZN(n17758) );
  NAND2_X1 U15238 ( .A1(n12072), .A2(n17758), .ZN(n17751) );
  NAND2_X1 U15239 ( .A1(n17752), .A2(n17751), .ZN(n17750) );
  NAND2_X1 U15240 ( .A1(n12073), .A2(n17750), .ZN(n17738) );
  NAND2_X1 U15241 ( .A1(n17737), .A2(n17738), .ZN(n17736) );
  NOR2_X1 U15242 ( .A1(n17737), .A2(n17738), .ZN(n12074) );
  AOI21_X1 U15243 ( .B1(n18004), .B2(n17736), .A(n12074), .ZN(n17724) );
  NAND2_X1 U15244 ( .A1(n17725), .A2(n17724), .ZN(n17723) );
  NAND2_X1 U15245 ( .A1(n12075), .A2(n17723), .ZN(n12077) );
  NAND2_X1 U15246 ( .A1(n12076), .A2(n12077), .ZN(n12078) );
  XOR2_X1 U15247 ( .A(n12077), .B(n12076), .Z(n17716) );
  NAND2_X1 U15248 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n17716), .ZN(
        n17715) );
  INV_X1 U15249 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18024) );
  NAND2_X1 U15250 ( .A1(n12083), .A2(n12079), .ZN(n12084) );
  INV_X1 U15251 ( .A(n12079), .ZN(n12082) );
  NAND2_X1 U15252 ( .A1(n17706), .A2(n17705), .ZN(n12081) );
  NAND2_X1 U15253 ( .A1(n12083), .A2(n12082), .ZN(n12080) );
  OAI211_X1 U15254 ( .C1(n12083), .C2(n12082), .A(n12081), .B(n12080), .ZN(
        n17682) );
  NAND2_X1 U15255 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n17682), .ZN(
        n17681) );
  INV_X1 U15256 ( .A(n17918), .ZN(n17465) );
  NAND3_X1 U15257 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n15623), .A3(
        n17791), .ZN(n12085) );
  XNOR2_X1 U15258 ( .A(n18728), .B(n12085), .ZN(n16297) );
  INV_X1 U15259 ( .A(n16297), .ZN(n12086) );
  NOR2_X2 U15260 ( .A1(n18760), .A2(n16417), .ZN(n17773) );
  NAND2_X1 U15261 ( .A1(n12086), .A2(n17773), .ZN(n12087) );
  NAND2_X1 U15262 ( .A1(n12090), .A2(n10245), .ZN(P3_U2799) );
  INV_X1 U15263 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n12275) );
  INV_X1 U15264 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n14990) );
  INV_X1 U15265 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n14951) );
  INV_X1 U15266 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n12092) );
  XNOR2_X1 U15267 ( .A(n12094), .B(n12092), .ZN(n15948) );
  INV_X1 U15268 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12093) );
  INV_X1 U15269 ( .A(n12094), .ZN(n12095) );
  AOI21_X1 U15270 ( .B1(n14951), .B2(n12125), .A(n12095), .ZN(n14949) );
  INV_X1 U15271 ( .A(n14949), .ZN(n15957) );
  NOR2_X1 U15272 ( .A1(n12097), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12098) );
  OR2_X1 U15273 ( .A1(n12096), .A2(n12098), .ZN(n15981) );
  AOI21_X1 U15274 ( .B1(n16078), .B2(n12110), .A(n12099), .ZN(n16069) );
  AOI21_X1 U15275 ( .B1(n16092), .B2(n12108), .A(n9880), .ZN(n16079) );
  AOI21_X1 U15276 ( .B1(n16098), .B2(n12107), .A(n12109), .ZN(n18924) );
  AOI21_X1 U15277 ( .B1(n16113), .B2(n12105), .A(n9871), .ZN(n16099) );
  AOI21_X1 U15278 ( .B1(n16124), .B2(n12104), .A(n12106), .ZN(n18967) );
  AOI21_X1 U15279 ( .B1(n14628), .B2(n12103), .A(n12100), .ZN(n14623) );
  AOI21_X1 U15280 ( .B1(n10565), .B2(n12102), .A(n12101), .ZN(n14651) );
  AOI22_X1 U15281 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n19836), .ZN(n15368) );
  AOI22_X1 U15282 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n12102), .B2(n19836), .ZN(
        n14664) );
  NAND2_X1 U15283 ( .A1(n15368), .A2(n14664), .ZN(n14663) );
  NOR2_X1 U15284 ( .A1(n14651), .A2(n14663), .ZN(n14634) );
  OAI21_X1 U15285 ( .B1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n12101), .A(
        n12103), .ZN(n14635) );
  NAND2_X1 U15286 ( .A1(n14634), .A2(n14635), .ZN(n14620) );
  NOR2_X1 U15287 ( .A1(n14623), .A2(n14620), .ZN(n18977) );
  OAI21_X1 U15288 ( .B1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n12100), .A(
        n12104), .ZN(n18979) );
  NAND2_X1 U15289 ( .A1(n18977), .A2(n18979), .ZN(n18965) );
  NOR2_X1 U15290 ( .A1(n18967), .A2(n18965), .ZN(n18947) );
  OAI21_X1 U15291 ( .B1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n12106), .A(
        n12105), .ZN(n18949) );
  NAND2_X1 U15292 ( .A1(n18947), .A2(n18949), .ZN(n14600) );
  NOR2_X1 U15293 ( .A1(n16099), .A2(n14600), .ZN(n18938) );
  OAI21_X1 U15294 ( .B1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n9871), .A(
        n12107), .ZN(n18940) );
  NAND2_X1 U15295 ( .A1(n18938), .A2(n18940), .ZN(n18923) );
  NOR2_X1 U15296 ( .A1(n18924), .A2(n18923), .ZN(n18918) );
  OAI21_X1 U15297 ( .B1(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n12109), .A(
        n12108), .ZN(n18921) );
  NAND2_X1 U15298 ( .A1(n18918), .A2(n18921), .ZN(n18916) );
  NOR2_X1 U15299 ( .A1(n16079), .A2(n18916), .ZN(n18897) );
  OAI21_X1 U15300 ( .B1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n9880), .A(
        n12110), .ZN(n18896) );
  NAND2_X1 U15301 ( .A1(n18897), .A2(n18896), .ZN(n14575) );
  NOR2_X1 U15302 ( .A1(n16069), .A2(n14575), .ZN(n18885) );
  OR2_X1 U15303 ( .A1(n12099), .A2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12111) );
  NAND2_X1 U15304 ( .A1(n12112), .A2(n12111), .ZN(n18887) );
  NAND2_X1 U15305 ( .A1(n18885), .A2(n18887), .ZN(n18872) );
  AOI21_X1 U15306 ( .B1(n12112), .B2(n18882), .A(n12114), .ZN(n18875) );
  INV_X1 U15307 ( .A(n12115), .ZN(n12113) );
  OAI21_X1 U15308 ( .B1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n12114), .A(
        n12113), .ZN(n18866) );
  NAND2_X1 U15309 ( .A1(n12116), .A2(n18864), .ZN(n18854) );
  OAI21_X1 U15310 ( .B1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n12115), .A(
        n12117), .ZN(n18855) );
  AOI21_X1 U15311 ( .B1(n18834), .B2(n12117), .A(n12118), .ZN(n15033) );
  INV_X1 U15312 ( .A(n15033), .ZN(n18842) );
  OAI21_X1 U15313 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n12118), .A(
        n9894), .ZN(n18829) );
  NAND2_X1 U15314 ( .A1(n18828), .A2(n18829), .ZN(n18827) );
  NAND2_X1 U15315 ( .A1(n18827), .A2(n18873), .ZN(n18817) );
  AOI21_X1 U15316 ( .B1(n9894), .B2(n12275), .A(n12119), .ZN(n12278) );
  INV_X1 U15317 ( .A(n12278), .ZN(n18818) );
  NAND2_X1 U15318 ( .A1(n18817), .A2(n18818), .ZN(n18816) );
  NAND2_X1 U15319 ( .A1(n18873), .A2(n18816), .ZN(n15578) );
  OAI21_X1 U15320 ( .B1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n12119), .A(
        n9846), .ZN(n16061) );
  NAND2_X1 U15321 ( .A1(n15578), .A2(n16061), .ZN(n15577) );
  NAND2_X1 U15322 ( .A1(n15577), .A2(n18873), .ZN(n16014) );
  AOI21_X1 U15323 ( .B1(n9846), .B2(n12091), .A(n12120), .ZN(n15011) );
  INV_X1 U15324 ( .A(n15011), .ZN(n16015) );
  NAND2_X1 U15325 ( .A1(n16014), .A2(n16015), .ZN(n16013) );
  NAND2_X1 U15326 ( .A1(n18873), .A2(n16013), .ZN(n16001) );
  OAI21_X1 U15327 ( .B1(n12120), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n12121), .ZN(n16002) );
  NAND2_X1 U15328 ( .A1(n16001), .A2(n16002), .ZN(n16000) );
  NAND2_X1 U15329 ( .A1(n16000), .A2(n18873), .ZN(n15991) );
  AOI21_X1 U15330 ( .B1(n14990), .B2(n12121), .A(n12097), .ZN(n14993) );
  INV_X1 U15331 ( .A(n14993), .ZN(n15992) );
  NAND2_X1 U15332 ( .A1(n15991), .A2(n15992), .ZN(n15990) );
  NAND2_X1 U15333 ( .A1(n18873), .A2(n15990), .ZN(n15980) );
  NAND2_X1 U15334 ( .A1(n15981), .A2(n15980), .ZN(n15979) );
  NAND2_X1 U15335 ( .A1(n15979), .A2(n12116), .ZN(n15970) );
  INV_X1 U15336 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n15962) );
  INV_X1 U15337 ( .A(n12096), .ZN(n12122) );
  AOI21_X1 U15338 ( .B1(n15962), .B2(n12122), .A(n12123), .ZN(n14972) );
  INV_X1 U15339 ( .A(n14972), .ZN(n15971) );
  NAND2_X1 U15340 ( .A1(n15970), .A2(n15971), .ZN(n15969) );
  NAND2_X1 U15341 ( .A1(n12116), .A2(n15969), .ZN(n14563) );
  OR2_X1 U15342 ( .A1(n12123), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12124) );
  NAND2_X1 U15343 ( .A1(n12125), .A2(n12124), .ZN(n14966) );
  NAND2_X1 U15344 ( .A1(n14563), .A2(n14966), .ZN(n14562) );
  NAND2_X1 U15345 ( .A1(n14562), .A2(n18873), .ZN(n15956) );
  NAND2_X1 U15346 ( .A1(n15957), .A2(n15956), .ZN(n15955) );
  NAND2_X1 U15347 ( .A1(n18873), .A2(n15955), .ZN(n15947) );
  NAND2_X1 U15348 ( .A1(n15948), .A2(n15947), .ZN(n12127) );
  OR4_X1 U15349 ( .A1(n15386), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(
        P2_STATE2_REG_2__SCAN_IN), .A4(P2_STATEBS16_REG_SCAN_IN), .ZN(n19705)
         );
  INV_X2 U15350 ( .A(n19705), .ZN(n18999) );
  INV_X1 U15351 ( .A(n15948), .ZN(n12126) );
  NOR2_X1 U15352 ( .A1(P2_EBX_REG_19__SCAN_IN), .A2(P2_EBX_REG_18__SCAN_IN), 
        .ZN(n12130) );
  NOR2_X1 U15353 ( .A1(n10808), .A2(n12130), .ZN(n12131) );
  INV_X1 U15354 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n14731) );
  NAND2_X1 U15355 ( .A1(n14865), .A2(n14886), .ZN(n12241) );
  NAND2_X1 U15356 ( .A1(n14912), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n14863) );
  INV_X1 U15357 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n12132) );
  NOR2_X1 U15358 ( .A1(n10808), .A2(n12132), .ZN(n14869) );
  INV_X1 U15359 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n14888) );
  NAND2_X1 U15360 ( .A1(n14912), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n14894) );
  INV_X1 U15361 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n12133) );
  NOR2_X1 U15362 ( .A1(n10808), .A2(n12133), .ZN(n14564) );
  NAND2_X1 U15363 ( .A1(n14912), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n14905) );
  NAND2_X1 U15364 ( .A1(n14906), .A2(n14905), .ZN(n14911) );
  NAND2_X1 U15365 ( .A1(n14912), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n12134) );
  XNOR2_X1 U15366 ( .A(n14911), .B(n12134), .ZN(n14908) );
  NOR2_X1 U15367 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n19844), .ZN(n12217) );
  INV_X1 U15368 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n16019) );
  NOR2_X1 U15369 ( .A1(n12217), .A2(n16019), .ZN(n12135) );
  NAND2_X1 U15370 ( .A1(n12218), .A2(n12135), .ZN(n12136) );
  NAND3_X1 U15371 ( .A1(n18785), .A2(P2_STATE2_REG_3__SCAN_IN), .A3(n19149), 
        .ZN(n16250) );
  NAND2_X1 U15372 ( .A1(n16250), .A2(n19705), .ZN(n12137) );
  NOR2_X1 U15373 ( .A1(n16186), .A2(n12137), .ZN(n12138) );
  AOI22_X1 U15374 ( .A1(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n18964), .B1(
        P2_REIP_REG_30__SCAN_IN), .B2(n18989), .ZN(n12139) );
  INV_X1 U15375 ( .A(n12139), .ZN(n12177) );
  AOI222_X1 U15376 ( .A1(P2_REIP_REG_30__SCAN_IN), .A2(n12156), .B1(n12151), 
        .B2(P2_EAX_REG_30__SCAN_IN), .C1(n10820), .C2(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12168) );
  AOI22_X1 U15377 ( .A1(n12151), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n10820), 
        .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n12142) );
  NAND2_X1 U15378 ( .A1(n12156), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n12141) );
  AOI22_X1 U15379 ( .A1(n12151), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n10820), 
        .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n12144) );
  NAND2_X1 U15380 ( .A1(n12156), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n12143) );
  NAND2_X1 U15381 ( .A1(n12144), .A2(n12143), .ZN(n14832) );
  AOI22_X1 U15382 ( .A1(n12151), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n10820), 
        .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n12146) );
  NAND2_X1 U15383 ( .A1(n12156), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n12145) );
  NAND2_X1 U15384 ( .A1(n12146), .A2(n12145), .ZN(n15247) );
  AOI22_X1 U15385 ( .A1(n12151), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n10820), 
        .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n12148) );
  NAND2_X1 U15386 ( .A1(n12156), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n12147) );
  NAND2_X1 U15387 ( .A1(n12148), .A2(n12147), .ZN(n12254) );
  AOI22_X1 U15388 ( .A1(n12151), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n10820), 
        .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n12150) );
  NAND2_X1 U15389 ( .A1(n12156), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n12149) );
  AOI22_X1 U15390 ( .A1(n12151), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n10820), 
        .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n12153) );
  NAND2_X1 U15391 ( .A1(n12156), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n12152) );
  NAND2_X1 U15392 ( .A1(n12153), .A2(n12152), .ZN(n14818) );
  AOI22_X1 U15393 ( .A1(n12151), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n10820), 
        .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n12155) );
  NAND2_X1 U15394 ( .A1(n12156), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n12154) );
  AND2_X1 U15395 ( .A1(n12155), .A2(n12154), .ZN(n14808) );
  AOI22_X1 U15396 ( .A1(n12151), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n10820), 
        .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n12158) );
  NAND2_X1 U15397 ( .A1(n12156), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n12157) );
  NAND2_X1 U15398 ( .A1(n12158), .A2(n12157), .ZN(n14797) );
  NAND2_X1 U15399 ( .A1(n14796), .A2(n14797), .ZN(n14799) );
  AOI22_X1 U15400 ( .A1(n12151), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n10820), 
        .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n12160) );
  NAND2_X1 U15401 ( .A1(n12156), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n12159) );
  AND2_X1 U15402 ( .A1(n12160), .A2(n12159), .ZN(n14789) );
  OR2_X2 U15403 ( .A1(n14799), .A2(n14789), .ZN(n14791) );
  AOI22_X1 U15404 ( .A1(n12151), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n10820), 
        .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n12162) );
  NAND2_X1 U15405 ( .A1(n12156), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n12161) );
  AND2_X1 U15406 ( .A1(n12162), .A2(n12161), .ZN(n14779) );
  OR2_X2 U15407 ( .A1(n14791), .A2(n14779), .ZN(n14780) );
  AOI22_X1 U15408 ( .A1(n12151), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n10820), 
        .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n12164) );
  NAND2_X1 U15409 ( .A1(n12156), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n12163) );
  AND2_X1 U15410 ( .A1(n12164), .A2(n12163), .ZN(n14567) );
  INV_X1 U15411 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n19768) );
  INV_X1 U15412 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15147) );
  INV_X1 U15413 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n14763) );
  OAI222_X1 U15414 ( .A1(n19768), .A2(n12167), .B1(n12166), .B2(n15147), .C1(
        n12165), .C2(n14763), .ZN(n14761) );
  INV_X1 U15415 ( .A(n15133), .ZN(n12175) );
  AND2_X1 U15416 ( .A1(n16220), .A2(n12217), .ZN(n16238) );
  NAND2_X1 U15417 ( .A1(n12172), .A2(n16238), .ZN(n12169) );
  INV_X1 U15418 ( .A(P2_EBX_REG_30__SCAN_IN), .ZN(n12174) );
  INV_X1 U15419 ( .A(n16238), .ZN(n12171) );
  NOR2_X1 U15420 ( .A1(P2_EBX_REG_31__SCAN_IN), .A2(n12217), .ZN(n12170) );
  AOI22_X1 U15421 ( .A1(n12172), .A2(n12171), .B1(n12170), .B2(n16218), .ZN(
        n12173) );
  OAI22_X1 U15422 ( .A1(n12175), .A2(n18982), .B1(n12174), .B2(n18960), .ZN(
        n12176) );
  AOI211_X1 U15423 ( .C1(n14908), .C2(n18950), .A(n12177), .B(n12176), .ZN(
        n12221) );
  INV_X1 U15424 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n12180) );
  NAND2_X1 U15425 ( .A1(n10992), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n12179) );
  NAND2_X1 U15426 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n12178) );
  OAI211_X1 U15427 ( .C1(n9775), .C2(n12180), .A(n12179), .B(n12178), .ZN(
        n12181) );
  AOI21_X1 U15428 ( .B1(n14924), .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n12181), .ZN(n15272) );
  INV_X1 U15429 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n16129) );
  AOI22_X1 U15430 ( .A1(n12209), .A2(P2_REIP_REG_19__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), 
        .ZN(n12183) );
  NAND2_X1 U15431 ( .A1(n10992), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n12182) );
  OAI211_X1 U15432 ( .C1(n10582), .C2(n16129), .A(n12183), .B(n12182), .ZN(
        n14738) );
  INV_X1 U15433 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n12248) );
  AOI22_X1 U15434 ( .A1(n12209), .A2(P2_REIP_REG_20__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), 
        .ZN(n12185) );
  NAND2_X1 U15435 ( .A1(n10992), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n12184) );
  OAI211_X1 U15436 ( .C1(n10582), .C2(n12248), .A(n12185), .B(n12184), .ZN(
        n15017) );
  NAND2_X1 U15437 ( .A1(n15018), .A2(n15017), .ZN(n12255) );
  INV_X1 U15438 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n19753) );
  NAND2_X1 U15439 ( .A1(n10992), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n12187) );
  NAND2_X1 U15440 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n12186) );
  OAI211_X1 U15441 ( .C1(n9775), .C2(n19753), .A(n12187), .B(n12186), .ZN(
        n12188) );
  AOI21_X1 U15442 ( .B1(n14924), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n12188), .ZN(n12256) );
  INV_X1 U15443 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n12191) );
  NAND2_X1 U15444 ( .A1(n10992), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n12190) );
  NAND2_X1 U15445 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n12189) );
  OAI211_X1 U15446 ( .C1(n9775), .C2(n12191), .A(n12190), .B(n12189), .ZN(
        n12192) );
  AOI21_X1 U15447 ( .B1(n14924), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n12192), .ZN(n15235) );
  INV_X1 U15448 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n19756) );
  NAND2_X1 U15449 ( .A1(n10992), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n12194) );
  NAND2_X1 U15450 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n12193) );
  OAI211_X1 U15451 ( .C1(n9775), .C2(n19756), .A(n12194), .B(n12193), .ZN(
        n12195) );
  AOI21_X1 U15452 ( .B1(n14924), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n12195), .ZN(n14724) );
  INV_X1 U15453 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n20991) );
  AOI22_X1 U15454 ( .A1(n12209), .A2(P2_REIP_REG_24__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), 
        .ZN(n12197) );
  NAND2_X1 U15455 ( .A1(n10992), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n12196) );
  OAI211_X1 U15456 ( .C1(n10582), .C2(n20991), .A(n12197), .B(n12196), .ZN(
        n14715) );
  INV_X1 U15457 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n19760) );
  NAND2_X1 U15458 ( .A1(n10992), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n12199) );
  NAND2_X1 U15459 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n12198) );
  OAI211_X1 U15460 ( .C1(n9775), .C2(n19760), .A(n12199), .B(n12198), .ZN(
        n12200) );
  AOI21_X1 U15461 ( .B1(n14924), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n12200), .ZN(n14709) );
  INV_X1 U15462 ( .A(n12201), .ZN(n14711) );
  INV_X1 U15463 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n19762) );
  NAND2_X1 U15464 ( .A1(n10992), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n12203) );
  NAND2_X1 U15465 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n12202) );
  OAI211_X1 U15466 ( .C1(n9775), .C2(n19762), .A(n12203), .B(n12202), .ZN(
        n12204) );
  AOI21_X1 U15467 ( .B1(n14924), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n12204), .ZN(n14701) );
  INV_X1 U15468 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15169) );
  AOI22_X1 U15469 ( .A1(n12209), .A2(P2_REIP_REG_27__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), 
        .ZN(n12206) );
  NAND2_X1 U15470 ( .A1(n10992), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n12205) );
  OAI211_X1 U15471 ( .C1(n10582), .C2(n15169), .A(n12206), .B(n12205), .ZN(
        n14689) );
  INV_X1 U15472 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15155) );
  AOI22_X1 U15473 ( .A1(n12209), .A2(P2_REIP_REG_28__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), 
        .ZN(n12208) );
  NAND2_X1 U15474 ( .A1(n10992), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n12207) );
  OAI211_X1 U15475 ( .C1(n10582), .C2(n15155), .A(n12208), .B(n12207), .ZN(
        n14561) );
  AOI22_X1 U15476 ( .A1(n12209), .A2(P2_REIP_REG_29__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n12211) );
  NAND2_X1 U15477 ( .A1(n10992), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n12210) );
  OAI211_X1 U15478 ( .C1(n10582), .C2(n15147), .A(n12211), .B(n12210), .ZN(
        n14675) );
  INV_X1 U15479 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n19772) );
  NAND2_X1 U15480 ( .A1(n10992), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n12213) );
  NAND2_X1 U15481 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n12212) );
  OAI211_X1 U15482 ( .C1(n9775), .C2(n19772), .A(n12213), .B(n12212), .ZN(
        n12214) );
  AOI21_X1 U15483 ( .B1(n14924), .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n12214), .ZN(n12215) );
  INV_X1 U15484 ( .A(n12215), .ZN(n12216) );
  NAND2_X1 U15485 ( .A1(n12218), .A2(n12217), .ZN(n12219) );
  NAND2_X1 U15486 ( .A1(n14912), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n12223) );
  MUX2_X1 U15487 ( .A(n14912), .B(n12223), .S(n12224), .Z(n12225) );
  OR2_X1 U15488 ( .A1(n12224), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n12229) );
  NAND2_X1 U15489 ( .A1(n12225), .A2(n12229), .ZN(n18847) );
  NAND2_X1 U15490 ( .A1(n11060), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12226) );
  OR2_X1 U15491 ( .A1(n18847), .A2(n12226), .ZN(n14857) );
  INV_X1 U15492 ( .A(n14857), .ZN(n15262) );
  INV_X1 U15493 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n12227) );
  NOR2_X1 U15494 ( .A1(n10808), .A2(n12227), .ZN(n12228) );
  NAND2_X1 U15495 ( .A1(n12229), .A2(n12228), .ZN(n12230) );
  NAND2_X1 U15496 ( .A1(n12230), .A2(n12235), .ZN(n18835) );
  INV_X1 U15497 ( .A(n18835), .ZN(n12232) );
  AND2_X1 U15498 ( .A1(n11060), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12231) );
  NAND2_X1 U15499 ( .A1(n12232), .A2(n12231), .ZN(n15026) );
  OR2_X1 U15500 ( .A1(n18847), .A2(n10849), .ZN(n12233) );
  INV_X1 U15501 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15278) );
  NAND2_X1 U15502 ( .A1(n12233), .A2(n15278), .ZN(n15028) );
  OAI21_X1 U15503 ( .B1(n18835), .B2(n10849), .A(n16129), .ZN(n15027) );
  NAND2_X1 U15504 ( .A1(n15028), .A2(n15027), .ZN(n14850) );
  NAND2_X1 U15505 ( .A1(n14912), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n12234) );
  XNOR2_X1 U15506 ( .A(n12235), .B(n12234), .ZN(n18823) );
  AOI21_X1 U15507 ( .B1(n18823), .B2(n11060), .A(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14849) );
  AND2_X1 U15508 ( .A1(n11060), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12236) );
  NAND2_X1 U15509 ( .A1(n18823), .A2(n12236), .ZN(n14858) );
  INV_X1 U15510 ( .A(n14858), .ZN(n12237) );
  NOR2_X1 U15511 ( .A1(n14849), .A2(n12237), .ZN(n15015) );
  NAND2_X1 U15512 ( .A1(n14912), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n12238) );
  NOR2_X1 U15513 ( .A1(n12239), .A2(n12238), .ZN(n12240) );
  OR2_X1 U15514 ( .A1(n12241), .A2(n12240), .ZN(n18811) );
  OR2_X1 U15515 ( .A1(n18811), .A2(n10849), .ZN(n12242) );
  INV_X1 U15516 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n12260) );
  NAND2_X1 U15517 ( .A1(n12242), .A2(n12260), .ZN(n14853) );
  NAND2_X1 U15518 ( .A1(n11060), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12243) );
  OR2_X1 U15519 ( .A1(n18811), .A2(n12243), .ZN(n14860) );
  NAND2_X1 U15520 ( .A1(n14853), .A2(n14860), .ZN(n12244) );
  AND3_X1 U15521 ( .A1(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n12245) );
  NAND2_X1 U15522 ( .A1(n12246), .A2(n12245), .ZN(n15271) );
  NOR2_X1 U15523 ( .A1(n15271), .A2(n15278), .ZN(n15251) );
  INV_X1 U15524 ( .A(n12249), .ZN(n12247) );
  NAND2_X1 U15525 ( .A1(n12247), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15034) );
  OAI21_X1 U15526 ( .B1(n15034), .B2(n12248), .A(n12260), .ZN(n12250) );
  AND2_X1 U15527 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n12261) );
  NAND2_X1 U15528 ( .A1(n12261), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12251) );
  NAND2_X1 U15529 ( .A1(n12250), .A2(n14918), .ZN(n12280) );
  OR2_X1 U15530 ( .A1(n12280), .A2(n16157), .ZN(n12265) );
  NOR3_X1 U15531 ( .A1(n15278), .A2(n15271), .A3(n12251), .ZN(n15215) );
  INV_X1 U15532 ( .A(n15215), .ZN(n12252) );
  NAND2_X1 U15533 ( .A1(n16138), .A2(n12252), .ZN(n12253) );
  AND2_X1 U15534 ( .A1(n16136), .A2(n12253), .ZN(n15240) );
  INV_X1 U15535 ( .A(n15240), .ZN(n15222) );
  OAI21_X1 U15536 ( .B1(n15249), .B2(n12254), .A(n15233), .ZN(n18813) );
  NAND2_X1 U15537 ( .A1(n12255), .A2(n12256), .ZN(n12257) );
  NAND2_X1 U15538 ( .A1(n15236), .A2(n12257), .ZN(n18814) );
  INV_X1 U15539 ( .A(n18814), .ZN(n12258) );
  NAND2_X1 U15540 ( .A1(n12258), .A2(n21130), .ZN(n12259) );
  NAND2_X1 U15541 ( .A1(n16186), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n12274) );
  OAI211_X1 U15542 ( .C1(n21133), .C2(n18813), .A(n12259), .B(n12274), .ZN(
        n12263) );
  AND2_X1 U15543 ( .A1(n15329), .A2(n15251), .ZN(n16130) );
  AND3_X1 U15544 ( .A1(n16130), .A2(n12261), .A3(n12260), .ZN(n12262) );
  AOI211_X1 U15545 ( .C1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n15222), .A(
        n12263), .B(n12262), .ZN(n12264) );
  OAI21_X1 U15546 ( .B1(n19826), .B2(n12268), .A(n12267), .ZN(n12269) );
  NAND2_X1 U15547 ( .A1(n12270), .A2(n16118), .ZN(n12283) );
  NOR2_X2 U15548 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19786) );
  OR2_X1 U15549 ( .A1(n19786), .A2(n19784), .ZN(n19805) );
  NAND2_X1 U15550 ( .A1(n19805), .A2(n19836), .ZN(n12271) );
  INV_X1 U15551 ( .A(n12326), .ZN(n12273) );
  INV_X1 U15552 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n19846) );
  NAND2_X1 U15553 ( .A1(n19846), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n12272) );
  NAND2_X1 U15554 ( .A1(n12273), .A2(n12272), .ZN(n13266) );
  OAI21_X1 U15555 ( .B1(n16125), .B2(n12275), .A(n12274), .ZN(n12277) );
  NOR2_X1 U15556 ( .A1(n15386), .A2(n19846), .ZN(n19806) );
  NOR2_X1 U15557 ( .A1(n18814), .A2(n16088), .ZN(n12276) );
  AOI211_X1 U15558 ( .C1(n16114), .C2(n12278), .A(n12277), .B(n12276), .ZN(
        n12279) );
  NAND2_X1 U15559 ( .A1(n12283), .A2(n12282), .ZN(P2_U2993) );
  NOR2_X1 U15560 ( .A1(n12284), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12285) );
  NAND2_X1 U15561 ( .A1(n12287), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12288) );
  NAND2_X1 U15562 ( .A1(n12289), .A2(n12288), .ZN(n12290) );
  XNOR2_X1 U15563 ( .A(n12290), .B(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n13976) );
  AOI22_X1 U15564 ( .A1(n13560), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n13276), .ZN(n12295) );
  INV_X1 U15565 ( .A(n12295), .ZN(n12296) );
  INV_X1 U15566 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n20749) );
  NOR2_X1 U15567 ( .A1(n20081), .A2(n20749), .ZN(n13971) );
  INV_X1 U15568 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n13452) );
  AND3_X1 U15569 ( .A1(n12297), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n13452), .ZN(n12298) );
  INV_X1 U15570 ( .A(n12299), .ZN(n12300) );
  NAND3_X1 U15571 ( .A1(n12301), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n12300), .ZN(n12302) );
  OAI21_X1 U15572 ( .B1(n13976), .B2(n15923), .A(n12303), .ZN(P1_U3000) );
  NAND2_X1 U15573 ( .A1(n12304), .A2(n12326), .ZN(n12310) );
  NAND2_X1 U15574 ( .A1(n12305), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12306) );
  NOR2_X1 U15575 ( .A1(n19804), .A2(n19813), .ZN(n19599) );
  NAND2_X1 U15576 ( .A1(n12314), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19644) );
  OAI211_X1 U15577 ( .C1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n12314), .A(
        n19644), .B(n19786), .ZN(n12307) );
  INV_X1 U15578 ( .A(n12307), .ZN(n12308) );
  AOI21_X1 U15579 ( .B1(n12323), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n12308), .ZN(n12309) );
  NAND3_X1 U15580 ( .A1(n12311), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n9779), 
        .ZN(n12338) );
  NOR2_X1 U15581 ( .A1(n12338), .A2(n12312), .ZN(n13477) );
  NAND2_X1 U15582 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19353) );
  NAND2_X1 U15583 ( .A1(n19353), .A2(n19804), .ZN(n12316) );
  INV_X1 U15584 ( .A(n12314), .ZN(n12315) );
  AND2_X1 U15585 ( .A1(n12316), .A2(n12315), .ZN(n19262) );
  AOI22_X1 U15586 ( .A1(n12323), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n19786), .B2(n19262), .ZN(n12317) );
  NAND2_X1 U15587 ( .A1(n12564), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n12332) );
  AOI22_X1 U15588 ( .A1(n12323), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n19786), .B2(n19821), .ZN(n12320) );
  NAND2_X1 U15589 ( .A1(n12564), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12328) );
  XNOR2_X1 U15590 ( .A(n12327), .B(n12328), .ZN(n13499) );
  NAND2_X1 U15591 ( .A1(n12323), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12324) );
  NAND2_X1 U15592 ( .A1(n19813), .A2(n19821), .ZN(n19382) );
  AND2_X1 U15593 ( .A1(n19353), .A2(n19382), .ZN(n19321) );
  NAND2_X1 U15594 ( .A1(n19321), .A2(n19786), .ZN(n19445) );
  NAND2_X1 U15595 ( .A1(n12324), .A2(n19445), .ZN(n12325) );
  INV_X1 U15596 ( .A(n12328), .ZN(n12329) );
  NAND2_X1 U15597 ( .A1(n13495), .A2(n13496), .ZN(n13494) );
  INV_X1 U15598 ( .A(n12332), .ZN(n12333) );
  NAND2_X1 U15599 ( .A1(n12331), .A2(n12333), .ZN(n12334) );
  NAND2_X1 U15600 ( .A1(n13479), .A2(n13476), .ZN(n12336) );
  INV_X1 U15601 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12337) );
  NOR2_X1 U15602 ( .A1(n12338), .A2(n12337), .ZN(n14616) );
  INV_X1 U15603 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12339) );
  NAND2_X1 U15604 ( .A1(n19029), .A2(n19028), .ZN(n13678) );
  AND2_X1 U15605 ( .A1(n19016), .A2(n19015), .ZN(n12342) );
  INV_X1 U15606 ( .A(n19011), .ZN(n12343) );
  AOI22_X1 U15607 ( .A1(n10412), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12443), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12347) );
  AOI22_X1 U15608 ( .A1(n10659), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10754), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12346) );
  AOI22_X1 U15609 ( .A1(n10850), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n15421), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12345) );
  AOI22_X1 U15610 ( .A1(n10658), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10789), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12344) );
  NAND4_X1 U15611 ( .A1(n12347), .A2(n12346), .A3(n12345), .A4(n12344), .ZN(
        n12353) );
  AOI22_X1 U15612 ( .A1(n10425), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12451), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12351) );
  AOI22_X1 U15613 ( .A1(n12450), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12449), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12350) );
  AOI22_X1 U15614 ( .A1(n12401), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10404), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12349) );
  AOI22_X1 U15615 ( .A1(n12448), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10653), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12348) );
  NAND4_X1 U15616 ( .A1(n12351), .A2(n12350), .A3(n12349), .A4(n12348), .ZN(
        n12352) );
  OR2_X1 U15617 ( .A1(n12353), .A2(n12352), .ZN(n13911) );
  AOI22_X1 U15618 ( .A1(n10412), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n12443), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12357) );
  AOI22_X1 U15619 ( .A1(n10659), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10754), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12356) );
  AOI22_X1 U15620 ( .A1(n10850), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n15421), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12355) );
  AOI22_X1 U15621 ( .A1(n10658), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n10789), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12354) );
  NAND4_X1 U15622 ( .A1(n12357), .A2(n12356), .A3(n12355), .A4(n12354), .ZN(
        n12363) );
  AOI22_X1 U15623 ( .A1(n10425), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12451), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12361) );
  AOI22_X1 U15624 ( .A1(n12450), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12449), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12360) );
  AOI22_X1 U15625 ( .A1(n12401), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n10404), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12359) );
  AOI22_X1 U15626 ( .A1(n12448), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10653), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12358) );
  NAND4_X1 U15627 ( .A1(n12361), .A2(n12360), .A3(n12359), .A4(n12358), .ZN(
        n12362) );
  OR2_X1 U15628 ( .A1(n12363), .A2(n12362), .ZN(n14742) );
  NAND2_X1 U15629 ( .A1(n13909), .A2(n14742), .ZN(n14733) );
  AOI22_X1 U15630 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n10412), .B1(
        n12443), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12367) );
  AOI22_X1 U15631 ( .A1(n10659), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10754), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12366) );
  AOI22_X1 U15632 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n15421), .B1(
        n10850), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12365) );
  AOI22_X1 U15633 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n10658), .B1(
        n10789), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12364) );
  NAND4_X1 U15634 ( .A1(n12367), .A2(n12366), .A3(n12365), .A4(n12364), .ZN(
        n12373) );
  AOI22_X1 U15635 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n10425), .B1(
        n12451), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12371) );
  AOI22_X1 U15636 ( .A1(n12450), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__3__SCAN_IN), .B2(n12449), .ZN(n12370) );
  AOI22_X1 U15637 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n12401), .B1(
        n10404), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12369) );
  AOI22_X1 U15638 ( .A1(n12448), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10653), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12368) );
  NAND4_X1 U15639 ( .A1(n12371), .A2(n12370), .A3(n12369), .A4(n12368), .ZN(
        n12372) );
  OR2_X1 U15640 ( .A1(n12373), .A2(n12372), .ZN(n14736) );
  INV_X1 U15641 ( .A(n14736), .ZN(n12384) );
  AOI22_X1 U15642 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n10412), .B1(
        n12443), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12377) );
  AOI22_X1 U15643 ( .A1(n10659), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10754), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12376) );
  AOI22_X1 U15644 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n15421), .B1(
        n10850), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12375) );
  AOI22_X1 U15645 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n10658), .B1(
        n10789), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12374) );
  NAND4_X1 U15646 ( .A1(n12377), .A2(n12376), .A3(n12375), .A4(n12374), .ZN(
        n12383) );
  AOI22_X1 U15647 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n10425), .B1(
        n12451), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12381) );
  AOI22_X1 U15648 ( .A1(n12450), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__2__SCAN_IN), .B2(n12449), .ZN(n12380) );
  AOI22_X1 U15649 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n12401), .B1(
        n10404), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12379) );
  AOI22_X1 U15650 ( .A1(n12448), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10653), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12378) );
  NAND4_X1 U15651 ( .A1(n12381), .A2(n12380), .A3(n12379), .A4(n12378), .ZN(
        n12382) );
  NOR2_X1 U15652 ( .A1(n12383), .A2(n12382), .ZN(n16031) );
  OR2_X1 U15653 ( .A1(n12384), .A2(n16031), .ZN(n12385) );
  AOI22_X1 U15654 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n10412), .B1(
        n12443), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12389) );
  AOI22_X1 U15655 ( .A1(n10659), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10754), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12388) );
  AOI22_X1 U15656 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n15421), .B1(
        n10850), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12387) );
  AOI22_X1 U15657 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n10658), .B1(
        n10789), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12386) );
  NAND4_X1 U15658 ( .A1(n12389), .A2(n12388), .A3(n12387), .A4(n12386), .ZN(
        n12395) );
  AOI22_X1 U15659 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n10425), .B1(
        n12451), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12393) );
  AOI22_X1 U15660 ( .A1(n12450), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__4__SCAN_IN), .B2(n12449), .ZN(n12392) );
  AOI22_X1 U15661 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n12401), .B1(
        n10404), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12391) );
  AOI22_X1 U15662 ( .A1(n12448), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10653), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12390) );
  NAND4_X1 U15663 ( .A1(n12393), .A2(n12392), .A3(n12391), .A4(n12390), .ZN(
        n12394) );
  NOR2_X1 U15664 ( .A1(n12395), .A2(n12394), .ZN(n16025) );
  INV_X1 U15665 ( .A(n16025), .ZN(n12396) );
  AOI22_X1 U15666 ( .A1(n10412), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12443), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12400) );
  AOI22_X1 U15667 ( .A1(n10659), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10754), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12399) );
  AOI22_X1 U15668 ( .A1(n10850), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n15421), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12398) );
  AOI22_X1 U15669 ( .A1(n10658), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10789), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12397) );
  NAND4_X1 U15670 ( .A1(n12400), .A2(n12399), .A3(n12398), .A4(n12397), .ZN(
        n12410) );
  AOI22_X1 U15671 ( .A1(n10425), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12451), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12408) );
  AOI22_X1 U15672 ( .A1(n12450), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12449), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12407) );
  AOI22_X1 U15673 ( .A1(n12401), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10404), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12406) );
  INV_X1 U15674 ( .A(n12448), .ZN(n12403) );
  OAI22_X1 U15675 ( .A1(n12403), .A2(n12582), .B1(n12402), .B2(n13571), .ZN(
        n12404) );
  INV_X1 U15676 ( .A(n12404), .ZN(n12405) );
  NAND4_X1 U15677 ( .A1(n12408), .A2(n12407), .A3(n12406), .A4(n12405), .ZN(
        n12409) );
  AOI22_X1 U15678 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n10412), .B1(
        n12443), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12414) );
  AOI22_X1 U15679 ( .A1(n10659), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10754), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12413) );
  AOI22_X1 U15680 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n15421), .B1(
        n10850), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12412) );
  AOI22_X1 U15681 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n10658), .B1(
        n10789), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12411) );
  NAND4_X1 U15682 ( .A1(n12414), .A2(n12413), .A3(n12412), .A4(n12411), .ZN(
        n12420) );
  AOI22_X1 U15683 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n10425), .B1(
        n12451), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12418) );
  AOI22_X1 U15684 ( .A1(n12450), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__6__SCAN_IN), .B2(n12449), .ZN(n12417) );
  AOI22_X1 U15685 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n10417), .B1(
        n10404), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12416) );
  AOI22_X1 U15686 ( .A1(n12448), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10653), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12415) );
  NAND4_X1 U15687 ( .A1(n12418), .A2(n12417), .A3(n12416), .A4(n12415), .ZN(
        n12419) );
  OR2_X1 U15688 ( .A1(n12420), .A2(n12419), .ZN(n16021) );
  INV_X1 U15689 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12422) );
  INV_X1 U15690 ( .A(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13806) );
  OAI22_X1 U15691 ( .A1(n9777), .A2(n12422), .B1(n12421), .B2(n13806), .ZN(
        n12426) );
  INV_X1 U15692 ( .A(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n19326) );
  INV_X1 U15693 ( .A(n12469), .ZN(n12437) );
  INV_X1 U15694 ( .A(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12423) );
  OAI22_X1 U15695 ( .A1(n19326), .A2(n12424), .B1(n12437), .B2(n12423), .ZN(
        n12425) );
  NOR2_X1 U15696 ( .A1(n12426), .A2(n12425), .ZN(n12429) );
  INV_X1 U15697 ( .A(n10386), .ZN(n12583) );
  AOI22_X1 U15698 ( .A1(n10386), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12622), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12428) );
  AOI22_X1 U15699 ( .A1(n10391), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10382), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12427) );
  XNOR2_X1 U15700 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12616) );
  NAND4_X1 U15701 ( .A1(n12429), .A2(n12428), .A3(n12427), .A4(n12616), .ZN(
        n12442) );
  INV_X1 U15702 ( .A(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12431) );
  INV_X1 U15703 ( .A(n10382), .ZN(n15414) );
  INV_X1 U15704 ( .A(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12430) );
  OAI22_X1 U15705 ( .A1(n9777), .A2(n12431), .B1(n15414), .B2(n12430), .ZN(
        n12436) );
  INV_X1 U15706 ( .A(n12612), .ZN(n12581) );
  INV_X1 U15707 ( .A(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12434) );
  INV_X1 U15708 ( .A(n12622), .ZN(n12586) );
  INV_X1 U15709 ( .A(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12433) );
  OAI22_X1 U15710 ( .A1(n12581), .A2(n12434), .B1(n12586), .B2(n12433), .ZN(
        n12435) );
  NOR2_X1 U15711 ( .A1(n12436), .A2(n12435), .ZN(n12440) );
  INV_X1 U15712 ( .A(n12616), .ZN(n12620) );
  AOI22_X1 U15713 ( .A1(n10392), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9818), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12439) );
  AOI22_X1 U15714 ( .A1(n9821), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12615), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12438) );
  NAND4_X1 U15715 ( .A1(n12440), .A2(n12620), .A3(n12439), .A4(n12438), .ZN(
        n12441) );
  AND2_X1 U15716 ( .A1(n12442), .A2(n12441), .ZN(n12486) );
  NAND2_X1 U15717 ( .A1(n9779), .A2(n12486), .ZN(n12461) );
  AOI22_X1 U15718 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n12443), .B1(
        n10425), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12447) );
  AOI22_X1 U15719 ( .A1(n10659), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10658), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12446) );
  AOI22_X1 U15720 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n10754), .B1(
        n10850), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12445) );
  AOI22_X1 U15721 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n15421), .B1(
        n10789), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12444) );
  NAND4_X1 U15722 ( .A1(n12447), .A2(n12446), .A3(n12445), .A4(n12444), .ZN(
        n12457) );
  AOI22_X1 U15723 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n10412), .B1(
        n12448), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12455) );
  AOI22_X1 U15724 ( .A1(n12450), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__7__SCAN_IN), .B2(n12449), .ZN(n12454) );
  AOI22_X1 U15725 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n10653), .B1(
        n10404), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12453) );
  AOI22_X1 U15726 ( .A1(n12451), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12401), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12452) );
  NAND4_X1 U15727 ( .A1(n12455), .A2(n12454), .A3(n12453), .A4(n12452), .ZN(
        n12456) );
  XNOR2_X1 U15728 ( .A(n12461), .B(n12488), .ZN(n12459) );
  NAND2_X1 U15729 ( .A1(n9776), .A2(n12486), .ZN(n14721) );
  INV_X1 U15730 ( .A(n12461), .ZN(n12462) );
  NAND2_X1 U15731 ( .A1(n12462), .A2(n12488), .ZN(n12484) );
  INV_X1 U15732 ( .A(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12464) );
  INV_X1 U15733 ( .A(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12463) );
  OAI22_X1 U15734 ( .A1(n12583), .A2(n12464), .B1(n12581), .B2(n12463), .ZN(
        n12468) );
  INV_X1 U15735 ( .A(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12466) );
  INV_X1 U15736 ( .A(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12465) );
  OAI22_X1 U15737 ( .A1(n12586), .A2(n12466), .B1(n15414), .B2(n12465), .ZN(
        n12467) );
  NOR2_X1 U15738 ( .A1(n12468), .A2(n12467), .ZN(n12472) );
  AOI22_X1 U15739 ( .A1(n10392), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n9818), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12471) );
  AOI22_X1 U15740 ( .A1(n12432), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n12615), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12470) );
  NAND4_X1 U15741 ( .A1(n12472), .A2(n12471), .A3(n12470), .A4(n12616), .ZN(
        n12483) );
  INV_X1 U15742 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12474) );
  INV_X1 U15743 ( .A(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12473) );
  OAI22_X1 U15744 ( .A1(n12583), .A2(n12474), .B1(n12581), .B2(n12473), .ZN(
        n12478) );
  INV_X1 U15745 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12476) );
  INV_X1 U15746 ( .A(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12475) );
  OAI22_X1 U15747 ( .A1(n12586), .A2(n12476), .B1(n15414), .B2(n12475), .ZN(
        n12477) );
  NOR2_X1 U15748 ( .A1(n12478), .A2(n12477), .ZN(n12481) );
  AOI22_X1 U15749 ( .A1(n10392), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n9818), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12480) );
  AOI22_X1 U15750 ( .A1(n12432), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12615), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12479) );
  NAND4_X1 U15751 ( .A1(n12481), .A2(n12620), .A3(n12480), .A4(n12479), .ZN(
        n12482) );
  NAND2_X1 U15752 ( .A1(n12483), .A2(n12482), .ZN(n12485) );
  INV_X1 U15753 ( .A(n12485), .ZN(n12487) );
  AND3_X1 U15754 ( .A1(n12488), .A2(n12487), .A3(n12486), .ZN(n12509) );
  INV_X1 U15755 ( .A(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12490) );
  INV_X1 U15756 ( .A(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12489) );
  OAI22_X1 U15757 ( .A1(n12583), .A2(n12490), .B1(n12581), .B2(n12489), .ZN(
        n12494) );
  INV_X1 U15758 ( .A(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12492) );
  INV_X1 U15759 ( .A(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12491) );
  OAI22_X1 U15760 ( .A1(n12586), .A2(n12492), .B1(n15414), .B2(n12491), .ZN(
        n12493) );
  NOR2_X1 U15761 ( .A1(n12494), .A2(n12493), .ZN(n12497) );
  AOI22_X1 U15762 ( .A1(n10392), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12469), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12496) );
  AOI22_X1 U15763 ( .A1(n12432), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12615), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12495) );
  NAND4_X1 U15764 ( .A1(n12497), .A2(n12496), .A3(n12495), .A4(n12616), .ZN(
        n12508) );
  INV_X1 U15765 ( .A(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12499) );
  INV_X1 U15766 ( .A(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12498) );
  OAI22_X1 U15767 ( .A1(n12583), .A2(n12499), .B1(n12581), .B2(n12498), .ZN(
        n12503) );
  INV_X1 U15768 ( .A(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12501) );
  INV_X1 U15769 ( .A(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12500) );
  OAI22_X1 U15770 ( .A1(n12586), .A2(n12501), .B1(n15414), .B2(n12500), .ZN(
        n12502) );
  NOR2_X1 U15771 ( .A1(n12503), .A2(n12502), .ZN(n12506) );
  AOI22_X1 U15772 ( .A1(n10392), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9818), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12505) );
  AOI22_X1 U15773 ( .A1(n12432), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12615), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12504) );
  NAND4_X1 U15774 ( .A1(n12506), .A2(n12620), .A3(n12505), .A4(n12504), .ZN(
        n12507) );
  AND2_X1 U15775 ( .A1(n12508), .A2(n12507), .ZN(n12510) );
  NAND2_X1 U15776 ( .A1(n12509), .A2(n12510), .ZN(n12559) );
  OAI211_X1 U15777 ( .C1(n12509), .C2(n12510), .A(n12564), .B(n12559), .ZN(
        n12513) );
  INV_X1 U15778 ( .A(n12510), .ZN(n12511) );
  NOR2_X1 U15779 ( .A1(n9779), .A2(n12511), .ZN(n14707) );
  INV_X1 U15780 ( .A(n12512), .ZN(n14807) );
  OAI22_X1 U15781 ( .A1(n12583), .A2(n12517), .B1(n12581), .B2(n12516), .ZN(
        n12521) );
  OAI22_X1 U15782 ( .A1(n12586), .A2(n12519), .B1(n15414), .B2(n12518), .ZN(
        n12520) );
  NOR2_X1 U15783 ( .A1(n12521), .A2(n12520), .ZN(n12524) );
  AOI22_X1 U15784 ( .A1(n10392), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12469), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12523) );
  AOI22_X1 U15785 ( .A1(n12432), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12615), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12522) );
  NAND4_X1 U15786 ( .A1(n12524), .A2(n12523), .A3(n12522), .A4(n12616), .ZN(
        n12535) );
  OAI22_X1 U15787 ( .A1(n12583), .A2(n12526), .B1(n12581), .B2(n12525), .ZN(
        n12530) );
  OAI22_X1 U15788 ( .A1(n12586), .A2(n12528), .B1(n15414), .B2(n12527), .ZN(
        n12529) );
  NOR2_X1 U15789 ( .A1(n12530), .A2(n12529), .ZN(n12533) );
  AOI22_X1 U15790 ( .A1(n10392), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9818), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12532) );
  AOI22_X1 U15791 ( .A1(n12432), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12615), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12531) );
  NAND4_X1 U15792 ( .A1(n12533), .A2(n12620), .A3(n12532), .A4(n12531), .ZN(
        n12534) );
  AND2_X1 U15793 ( .A1(n12535), .A2(n12534), .ZN(n12560) );
  XNOR2_X1 U15794 ( .A(n12559), .B(n12560), .ZN(n12536) );
  NAND2_X1 U15795 ( .A1(n9776), .A2(n12560), .ZN(n14699) );
  INV_X1 U15796 ( .A(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12540) );
  INV_X1 U15797 ( .A(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12539) );
  OAI22_X1 U15798 ( .A1(n12583), .A2(n12540), .B1(n12581), .B2(n12539), .ZN(
        n12544) );
  INV_X1 U15799 ( .A(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12542) );
  INV_X1 U15800 ( .A(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12541) );
  OAI22_X1 U15801 ( .A1(n12586), .A2(n12542), .B1(n15414), .B2(n12541), .ZN(
        n12543) );
  NOR2_X1 U15802 ( .A1(n12544), .A2(n12543), .ZN(n12547) );
  AOI22_X1 U15803 ( .A1(n10392), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12469), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12546) );
  AOI22_X1 U15804 ( .A1(n12432), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n12615), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12545) );
  NAND4_X1 U15805 ( .A1(n12547), .A2(n12546), .A3(n12545), .A4(n12616), .ZN(
        n12558) );
  INV_X1 U15806 ( .A(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12549) );
  INV_X1 U15807 ( .A(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12548) );
  OAI22_X1 U15808 ( .A1(n12583), .A2(n12549), .B1(n12581), .B2(n12548), .ZN(
        n12553) );
  INV_X1 U15809 ( .A(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12551) );
  INV_X1 U15810 ( .A(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12550) );
  OAI22_X1 U15811 ( .A1(n12586), .A2(n12551), .B1(n15414), .B2(n12550), .ZN(
        n12552) );
  NOR2_X1 U15812 ( .A1(n12553), .A2(n12552), .ZN(n12556) );
  AOI22_X1 U15813 ( .A1(n10392), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n9818), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12555) );
  AOI22_X1 U15814 ( .A1(n12432), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12615), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12554) );
  NAND4_X1 U15815 ( .A1(n12556), .A2(n12620), .A3(n12555), .A4(n12554), .ZN(
        n12557) );
  NAND2_X1 U15816 ( .A1(n12558), .A2(n12557), .ZN(n12562) );
  INV_X1 U15817 ( .A(n12562), .ZN(n12569) );
  INV_X1 U15818 ( .A(n12559), .ZN(n12561) );
  NAND2_X1 U15819 ( .A1(n12561), .A2(n12560), .ZN(n12563) );
  INV_X1 U15820 ( .A(n12563), .ZN(n12565) );
  OAI211_X1 U15821 ( .C1(n12569), .C2(n12565), .A(n14683), .B(n12564), .ZN(
        n12566) );
  NAND2_X1 U15822 ( .A1(n12567), .A2(n12566), .ZN(n12568) );
  NAND2_X1 U15823 ( .A1(n9776), .A2(n12569), .ZN(n14694) );
  OAI22_X1 U15824 ( .A1(n12583), .A2(n12572), .B1(n12581), .B2(n12571), .ZN(
        n12576) );
  OAI22_X1 U15825 ( .A1(n12586), .A2(n12574), .B1(n15414), .B2(n12573), .ZN(
        n12575) );
  NOR2_X1 U15826 ( .A1(n12576), .A2(n12575), .ZN(n12579) );
  AOI22_X1 U15827 ( .A1(n10392), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12469), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12578) );
  AOI22_X1 U15828 ( .A1(n12432), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12615), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12577) );
  NAND4_X1 U15829 ( .A1(n12579), .A2(n12578), .A3(n12577), .A4(n12616), .ZN(
        n12593) );
  OAI22_X1 U15830 ( .A1(n12583), .A2(n12582), .B1(n12581), .B2(n12580), .ZN(
        n12588) );
  OAI22_X1 U15831 ( .A1(n12586), .A2(n12585), .B1(n15414), .B2(n12584), .ZN(
        n12587) );
  NOR2_X1 U15832 ( .A1(n12588), .A2(n12587), .ZN(n12591) );
  AOI22_X1 U15833 ( .A1(n10392), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n9818), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12590) );
  AOI22_X1 U15834 ( .A1(n12432), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12615), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12589) );
  NAND4_X1 U15835 ( .A1(n12591), .A2(n12620), .A3(n12590), .A4(n12589), .ZN(
        n12592) );
  AND2_X1 U15836 ( .A1(n12593), .A2(n12592), .ZN(n14684) );
  INV_X1 U15837 ( .A(n14684), .ZN(n12594) );
  NOR3_X1 U15838 ( .A1(n14683), .A2(n9776), .A3(n12594), .ZN(n12609) );
  AOI22_X1 U15839 ( .A1(n10386), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n10382), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12596) );
  AOI22_X1 U15840 ( .A1(n10391), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12622), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12595) );
  NAND2_X1 U15841 ( .A1(n12596), .A2(n12595), .ZN(n12606) );
  AOI22_X1 U15842 ( .A1(n12432), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12615), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12598) );
  AOI22_X1 U15843 ( .A1(n10392), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n9818), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12597) );
  NAND3_X1 U15844 ( .A1(n12598), .A2(n12597), .A3(n12616), .ZN(n12605) );
  AOI22_X1 U15845 ( .A1(n12432), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12615), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12600) );
  AOI22_X1 U15846 ( .A1(n10392), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12469), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12599) );
  NAND3_X1 U15847 ( .A1(n12600), .A2(n12620), .A3(n12599), .ZN(n12604) );
  AOI22_X1 U15848 ( .A1(n9820), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10382), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12602) );
  AOI22_X1 U15849 ( .A1(n10391), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12622), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12601) );
  NAND2_X1 U15850 ( .A1(n12602), .A2(n12601), .ZN(n12603) );
  OAI22_X1 U15851 ( .A1(n12606), .A2(n12605), .B1(n12604), .B2(n12603), .ZN(
        n12607) );
  INV_X1 U15852 ( .A(n12607), .ZN(n12608) );
  NAND2_X1 U15853 ( .A1(n12609), .A2(n12608), .ZN(n12610) );
  OAI21_X1 U15854 ( .B1(n12609), .B2(n12608), .A(n12610), .ZN(n14680) );
  INV_X1 U15855 ( .A(n12610), .ZN(n12611) );
  NOR2_X1 U15856 ( .A1(n14679), .A2(n12611), .ZN(n12630) );
  INV_X1 U15857 ( .A(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n21056) );
  AOI22_X1 U15858 ( .A1(n9821), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12612), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12614) );
  NAND2_X1 U15859 ( .A1(n12622), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n12613) );
  OAI211_X1 U15860 ( .C1(n15414), .C2(n21056), .A(n12614), .B(n12613), .ZN(
        n12628) );
  AOI22_X1 U15861 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n12432), .B1(
        n12615), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12618) );
  AOI22_X1 U15862 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n10392), .B1(
        n9818), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12617) );
  NAND3_X1 U15863 ( .A1(n12618), .A2(n12617), .A3(n12616), .ZN(n12627) );
  AOI22_X1 U15864 ( .A1(n12432), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12615), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12621) );
  AOI22_X1 U15865 ( .A1(n10392), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12469), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12619) );
  NAND3_X1 U15866 ( .A1(n12621), .A2(n12620), .A3(n12619), .ZN(n12626) );
  AOI22_X1 U15867 ( .A1(n9820), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10391), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12624) );
  AOI22_X1 U15868 ( .A1(n12622), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n10382), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12623) );
  NAND2_X1 U15869 ( .A1(n12624), .A2(n12623), .ZN(n12625) );
  OAI22_X1 U15870 ( .A1(n12628), .A2(n12627), .B1(n12626), .B2(n12625), .ZN(
        n12629) );
  XNOR2_X1 U15871 ( .A(n12630), .B(n12629), .ZN(n13956) );
  AND3_X1 U15872 ( .A1(n16212), .A2(n10495), .A3(n19835), .ZN(n12631) );
  AND2_X1 U15873 ( .A1(n16223), .A2(n12631), .ZN(n12632) );
  AOI21_X1 U15874 ( .B1(n16217), .B2(n16211), .A(n12632), .ZN(n15381) );
  NAND2_X1 U15875 ( .A1(n12633), .A2(n13348), .ZN(n12634) );
  NAND2_X1 U15876 ( .A1(n15381), .A2(n12634), .ZN(n12635) );
  NAND2_X1 U15877 ( .A1(n14912), .A2(n10480), .ZN(n12637) );
  NOR4_X1 U15878 ( .A1(P2_ADDRESS_REG_17__SCAN_IN), .A2(
        P2_ADDRESS_REG_16__SCAN_IN), .A3(P2_ADDRESS_REG_15__SCAN_IN), .A4(
        P2_ADDRESS_REG_14__SCAN_IN), .ZN(n12641) );
  NOR4_X1 U15879 ( .A1(P2_ADDRESS_REG_21__SCAN_IN), .A2(
        P2_ADDRESS_REG_20__SCAN_IN), .A3(P2_ADDRESS_REG_19__SCAN_IN), .A4(
        P2_ADDRESS_REG_18__SCAN_IN), .ZN(n12640) );
  NOR4_X1 U15880 ( .A1(P2_ADDRESS_REG_8__SCAN_IN), .A2(
        P2_ADDRESS_REG_7__SCAN_IN), .A3(P2_ADDRESS_REG_6__SCAN_IN), .A4(
        P2_ADDRESS_REG_4__SCAN_IN), .ZN(n12639) );
  NOR4_X1 U15881 ( .A1(P2_ADDRESS_REG_13__SCAN_IN), .A2(
        P2_ADDRESS_REG_12__SCAN_IN), .A3(P2_ADDRESS_REG_10__SCAN_IN), .A4(
        P2_ADDRESS_REG_9__SCAN_IN), .ZN(n12638) );
  NAND4_X1 U15882 ( .A1(n12641), .A2(n12640), .A3(n12639), .A4(n12638), .ZN(
        n12646) );
  NOR4_X1 U15883 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_11__SCAN_IN), .A4(
        P2_ADDRESS_REG_5__SCAN_IN), .ZN(n12644) );
  NOR4_X1 U15884 ( .A1(P2_ADDRESS_REG_25__SCAN_IN), .A2(
        P2_ADDRESS_REG_24__SCAN_IN), .A3(P2_ADDRESS_REG_23__SCAN_IN), .A4(
        P2_ADDRESS_REG_22__SCAN_IN), .ZN(n12643) );
  NOR4_X1 U15885 ( .A1(P2_ADDRESS_REG_2__SCAN_IN), .A2(
        P2_ADDRESS_REG_28__SCAN_IN), .A3(P2_ADDRESS_REG_27__SCAN_IN), .A4(
        P2_ADDRESS_REG_26__SCAN_IN), .ZN(n12642) );
  INV_X1 U15886 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n19730) );
  NAND4_X1 U15887 ( .A1(n12644), .A2(n12643), .A3(n12642), .A4(n19730), .ZN(
        n12645) );
  INV_X1 U15888 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n14223) );
  OR2_X1 U15889 ( .A1(n14769), .A2(n14223), .ZN(n12649) );
  NAND2_X1 U15890 ( .A1(n14769), .A2(BUF2_REG_14__SCAN_IN), .ZN(n12648) );
  AND2_X1 U15891 ( .A1(n12649), .A2(n12648), .ZN(n19137) );
  INV_X1 U15892 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n12650) );
  OAI22_X1 U15893 ( .A1(n14841), .A2(n19137), .B1(n19044), .B2(n12650), .ZN(
        n12651) );
  AOI21_X1 U15894 ( .B1(n15133), .B2(n19084), .A(n12651), .ZN(n12654) );
  INV_X1 U15895 ( .A(n10525), .ZN(n12652) );
  OR2_X1 U15896 ( .A1(n19083), .A2(n12652), .ZN(n13406) );
  NOR2_X2 U15897 ( .A1(n13406), .A2(n13781), .ZN(n16048) );
  NOR2_X2 U15898 ( .A1(n13406), .A2(n14769), .ZN(n16049) );
  AOI22_X1 U15899 ( .A1(n16048), .A2(BUF2_REG_30__SCAN_IN), .B1(n16049), .B2(
        BUF1_REG_30__SCAN_IN), .ZN(n12653) );
  OAI21_X1 U15900 ( .B1(n13956), .B2(n19079), .A(n12655), .ZN(P2_U2889) );
  NAND2_X1 U15901 ( .A1(n13957), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12690) );
  XNOR2_X1 U15902 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13828) );
  AOI21_X1 U15903 ( .B1(n13201), .B2(n13828), .A(n13960), .ZN(n12657) );
  INV_X2 U15904 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n20623) );
  NAND2_X1 U15905 ( .A1(n13961), .A2(P1_EAX_REG_2__SCAN_IN), .ZN(n12656) );
  OAI211_X1 U15906 ( .C1(n12690), .C2(n13447), .A(n12657), .B(n12656), .ZN(
        n12658) );
  INV_X1 U15907 ( .A(n12658), .ZN(n12659) );
  NAND2_X1 U15908 ( .A1(n12660), .A2(n12659), .ZN(n12661) );
  NAND2_X1 U15909 ( .A1(n13960), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12681) );
  NAND2_X1 U15910 ( .A1(n12661), .A2(n12681), .ZN(n13620) );
  NAND2_X1 U15911 ( .A1(n20543), .A2(n12838), .ZN(n12669) );
  NAND2_X1 U15912 ( .A1(n13961), .A2(P1_EAX_REG_1__SCAN_IN), .ZN(n12665) );
  NAND2_X1 U15913 ( .A1(n20623), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12664) );
  OAI211_X1 U15914 ( .C1(n12690), .C2(n12666), .A(n12665), .B(n12664), .ZN(
        n12667) );
  INV_X1 U15915 ( .A(n12667), .ZN(n12668) );
  NAND2_X1 U15916 ( .A1(n12669), .A2(n12668), .ZN(n13577) );
  NAND2_X1 U15917 ( .A1(n20179), .A2(n9772), .ZN(n12671) );
  NAND2_X1 U15918 ( .A1(n12671), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13408) );
  NAND2_X1 U15919 ( .A1(n12673), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n12675) );
  NAND2_X1 U15920 ( .A1(n20623), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12674) );
  OAI211_X1 U15921 ( .C1(n12690), .C2(n11132), .A(n12675), .B(n12674), .ZN(
        n12676) );
  AOI21_X1 U15922 ( .B1(n12672), .B2(n12838), .A(n12676), .ZN(n13407) );
  OR2_X1 U15923 ( .A1(n13408), .A2(n13407), .ZN(n13410) );
  INV_X1 U15924 ( .A(n13407), .ZN(n12677) );
  OR2_X1 U15925 ( .A1(n12677), .A2(n12695), .ZN(n12678) );
  NAND2_X1 U15926 ( .A1(n13410), .A2(n12678), .ZN(n13576) );
  NAND2_X1 U15927 ( .A1(n13577), .A2(n13576), .ZN(n13623) );
  NAND2_X1 U15928 ( .A1(n12680), .A2(n12679), .ZN(n13621) );
  NAND2_X1 U15929 ( .A1(n13621), .A2(n12681), .ZN(n13711) );
  NAND2_X1 U15930 ( .A1(n20763), .A2(n12838), .ZN(n12689) );
  AND2_X1 U15931 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12684) );
  INV_X1 U15932 ( .A(n12694), .ZN(n12683) );
  OAI21_X1 U15933 ( .B1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n12684), .A(
        n12683), .ZN(n13842) );
  AOI22_X1 U15934 ( .A1(n13201), .A2(n13842), .B1(n13960), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n12686) );
  NAND2_X1 U15935 ( .A1(n13961), .A2(P1_EAX_REG_3__SCAN_IN), .ZN(n12685) );
  OAI211_X1 U15936 ( .C1(n12690), .C2(n13558), .A(n12686), .B(n12685), .ZN(
        n12687) );
  INV_X1 U15937 ( .A(n12687), .ZN(n12688) );
  NAND2_X1 U15938 ( .A1(n12689), .A2(n12688), .ZN(n13712) );
  NAND2_X1 U15939 ( .A1(n13711), .A2(n13712), .ZN(n13732) );
  INV_X1 U15940 ( .A(n12690), .ZN(n12691) );
  NAND2_X1 U15941 ( .A1(n12691), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n12698) );
  INV_X1 U15942 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n12692) );
  AOI21_X1 U15943 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n12692), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12693) );
  AOI21_X1 U15944 ( .B1(n13961), .B2(P1_EAX_REG_4__SCAN_IN), .A(n12693), .ZN(
        n12697) );
  OAI21_X1 U15945 ( .B1(n12694), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n12702), .ZN(n20042) );
  NOR2_X1 U15946 ( .A1(n20042), .A2(n12695), .ZN(n12696) );
  AOI21_X1 U15947 ( .B1(n12698), .B2(n12697), .A(n12696), .ZN(n12699) );
  AOI21_X1 U15948 ( .B1(n12700), .B2(n12838), .A(n12699), .ZN(n13733) );
  INV_X1 U15949 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n13759) );
  INV_X1 U15950 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n12701) );
  NAND2_X1 U15951 ( .A1(n12702), .A2(n12701), .ZN(n12704) );
  NAND2_X1 U15952 ( .A1(n12704), .A2(n12709), .ZN(n19936) );
  INV_X2 U15953 ( .A(n12695), .ZN(n13201) );
  AOI22_X1 U15954 ( .A1(n19936), .A2(n13201), .B1(n13960), .B2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n12705) );
  OAI21_X1 U15955 ( .B1(n12893), .B2(n13759), .A(n12705), .ZN(n12706) );
  INV_X1 U15956 ( .A(n13755), .ZN(n12708) );
  OAI21_X1 U15957 ( .B1(n12710), .B2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n12715), .ZN(n19916) );
  INV_X1 U15958 ( .A(n19916), .ZN(n12714) );
  NAND2_X1 U15959 ( .A1(n12711), .A2(n12838), .ZN(n12713) );
  AOI22_X1 U15960 ( .A1(n13961), .A2(P1_EAX_REG_6__SCAN_IN), .B1(n13960), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n12712) );
  OAI211_X1 U15961 ( .C1(n12695), .C2(n12714), .A(n12713), .B(n12712), .ZN(
        n13823) );
  INV_X1 U15962 ( .A(n13822), .ZN(n12722) );
  OAI21_X1 U15963 ( .B1(n12716), .B2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n12738), .ZN(n19904) );
  NAND2_X1 U15964 ( .A1(n19904), .A2(n13201), .ZN(n12718) );
  AOI22_X1 U15965 ( .A1(n13961), .A2(P1_EAX_REG_7__SCAN_IN), .B1(n13960), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n12717) );
  NAND2_X1 U15966 ( .A1(n12718), .A2(n12717), .ZN(n12719) );
  AOI21_X1 U15967 ( .B1(n12720), .B2(n12838), .A(n12719), .ZN(n13871) );
  INV_X1 U15968 ( .A(n13871), .ZN(n12721) );
  XNOR2_X1 U15969 ( .A(n12738), .B(n14132), .ZN(n14133) );
  NAND2_X1 U15970 ( .A1(n14133), .A2(n13201), .ZN(n12737) );
  AOI22_X1 U15971 ( .A1(n13050), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n13112), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12726) );
  AOI22_X1 U15972 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n13128), .B1(
        n11398), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12725) );
  AOI22_X1 U15973 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n12901), .B1(
        n12965), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12724) );
  AOI22_X1 U15974 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n13090), .B1(
        n13540), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12723) );
  NAND4_X1 U15975 ( .A1(n12726), .A2(n12725), .A3(n12724), .A4(n12723), .ZN(
        n12732) );
  AOI22_X1 U15976 ( .A1(n12937), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12867), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12730) );
  AOI22_X1 U15977 ( .A1(n12921), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12964), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12729) );
  AOI22_X1 U15978 ( .A1(n12978), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n13134), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12728) );
  AOI22_X1 U15979 ( .A1(n12957), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9825), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12727) );
  NAND4_X1 U15980 ( .A1(n12730), .A2(n12729), .A3(n12728), .A4(n12727), .ZN(
        n12731) );
  OAI21_X1 U15981 ( .B1(n12732), .B2(n12731), .A(n12838), .ZN(n12735) );
  NAND2_X1 U15982 ( .A1(n13961), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n12734) );
  NAND2_X1 U15983 ( .A1(n13960), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12733) );
  XOR2_X1 U15984 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B(n12752), .Z(n19890) );
  AOI22_X1 U15985 ( .A1(n12978), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n13540), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12742) );
  AOI22_X1 U15986 ( .A1(n12937), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12965), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12741) );
  AOI22_X1 U15987 ( .A1(n13090), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12867), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12740) );
  AOI22_X1 U15988 ( .A1(n13112), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n13134), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12739) );
  NAND4_X1 U15989 ( .A1(n12742), .A2(n12741), .A3(n12740), .A4(n12739), .ZN(
        n12748) );
  AOI22_X1 U15990 ( .A1(n13050), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12921), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12746) );
  AOI22_X1 U15991 ( .A1(n11398), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12964), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12745) );
  AOI22_X1 U15992 ( .A1(n12901), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n11317), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12744) );
  AOI22_X1 U15993 ( .A1(n13128), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n9825), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12743) );
  NAND4_X1 U15994 ( .A1(n12746), .A2(n12745), .A3(n12744), .A4(n12743), .ZN(
        n12747) );
  OR2_X1 U15995 ( .A1(n12748), .A2(n12747), .ZN(n12749) );
  AOI22_X1 U15996 ( .A1(n12838), .A2(n12749), .B1(n13960), .B2(
        P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n12751) );
  NAND2_X1 U15997 ( .A1(n13961), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n12750) );
  OAI211_X1 U15998 ( .C1(n19890), .C2(n12695), .A(n12751), .B(n12750), .ZN(
        n13919) );
  XNOR2_X1 U15999 ( .A(n12779), .B(n13224), .ZN(n14434) );
  AOI22_X1 U16000 ( .A1(n13128), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13540), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12756) );
  AOI22_X1 U16001 ( .A1(n12937), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12867), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12755) );
  AOI22_X1 U16002 ( .A1(n11398), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n13134), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12754) );
  AOI22_X1 U16003 ( .A1(n12901), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n11317), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12753) );
  NAND4_X1 U16004 ( .A1(n12756), .A2(n12755), .A3(n12754), .A4(n12753), .ZN(
        n12762) );
  AOI22_X1 U16005 ( .A1(n13050), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n13112), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12760) );
  AOI22_X1 U16006 ( .A1(n12978), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n13090), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12759) );
  AOI22_X1 U16007 ( .A1(n12921), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12964), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12758) );
  AOI22_X1 U16008 ( .A1(n12965), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9825), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12757) );
  NAND4_X1 U16009 ( .A1(n12760), .A2(n12759), .A3(n12758), .A4(n12757), .ZN(
        n12761) );
  OAI21_X1 U16010 ( .B1(n12762), .B2(n12761), .A(n12838), .ZN(n12765) );
  NAND2_X1 U16011 ( .A1(n13961), .A2(P1_EAX_REG_10__SCAN_IN), .ZN(n12764) );
  NAND2_X1 U16012 ( .A1(n13960), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12763) );
  NAND3_X1 U16013 ( .A1(n12765), .A2(n12764), .A3(n12763), .ZN(n12766) );
  AOI21_X1 U16014 ( .B1(n14434), .B2(n13201), .A(n12766), .ZN(n13199) );
  AOI22_X1 U16015 ( .A1(n13050), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13112), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12771) );
  AOI22_X1 U16016 ( .A1(n12921), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11398), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12770) );
  AOI22_X1 U16017 ( .A1(n12978), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13540), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12769) );
  AOI22_X1 U16018 ( .A1(n12937), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n9825), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12768) );
  NAND4_X1 U16019 ( .A1(n12771), .A2(n12770), .A3(n12769), .A4(n12768), .ZN(
        n12777) );
  AOI22_X1 U16020 ( .A1(n13090), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12965), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12775) );
  AOI22_X1 U16021 ( .A1(n13128), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12867), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12774) );
  AOI22_X1 U16022 ( .A1(n12964), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n13134), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12773) );
  AOI22_X1 U16023 ( .A1(n12901), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12957), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12772) );
  NAND4_X1 U16024 ( .A1(n12775), .A2(n12774), .A3(n12773), .A4(n12772), .ZN(
        n12776) );
  OR2_X1 U16025 ( .A1(n12777), .A2(n12776), .ZN(n12778) );
  NAND2_X1 U16026 ( .A1(n12838), .A2(n12778), .ZN(n14215) );
  INV_X1 U16027 ( .A(n13960), .ZN(n12782) );
  INV_X1 U16028 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n15729) );
  OAI21_X1 U16029 ( .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n12780), .A(
        n12808), .ZN(n15780) );
  NAND2_X1 U16030 ( .A1(n15780), .A2(n13201), .ZN(n12781) );
  OAI21_X1 U16031 ( .B1(n12782), .B2(n15729), .A(n12781), .ZN(n12783) );
  AOI21_X1 U16032 ( .B1(n13961), .B2(P1_EAX_REG_11__SCAN_IN), .A(n12783), .ZN(
        n14118) );
  NAND2_X1 U16033 ( .A1(n12785), .A2(n12784), .ZN(n14117) );
  XOR2_X1 U16034 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B(n12824), .Z(
        n14427) );
  AOI22_X1 U16035 ( .A1(n13961), .A2(P1_EAX_REG_13__SCAN_IN), .B1(n13960), 
        .B2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n12797) );
  AOI22_X1 U16036 ( .A1(n13112), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11398), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12789) );
  AOI22_X1 U16037 ( .A1(n12978), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n13128), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12788) );
  AOI22_X1 U16038 ( .A1(n12937), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12965), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12787) );
  AOI22_X1 U16039 ( .A1(n12901), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n9825), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12786) );
  NAND4_X1 U16040 ( .A1(n12789), .A2(n12788), .A3(n12787), .A4(n12786), .ZN(
        n12795) );
  AOI22_X1 U16041 ( .A1(n13050), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12921), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12793) );
  AOI22_X1 U16042 ( .A1(n13540), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12867), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12792) );
  AOI22_X1 U16043 ( .A1(n12964), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n13134), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12791) );
  AOI22_X1 U16044 ( .A1(n13090), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12957), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12790) );
  NAND4_X1 U16045 ( .A1(n12793), .A2(n12792), .A3(n12791), .A4(n12790), .ZN(
        n12794) );
  OAI21_X1 U16046 ( .B1(n12795), .B2(n12794), .A(n12838), .ZN(n12796) );
  OAI211_X1 U16047 ( .C1(n14427), .C2(n12695), .A(n12797), .B(n12796), .ZN(
        n14120) );
  INV_X1 U16048 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n14295) );
  AOI22_X1 U16049 ( .A1(n13050), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12921), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12801) );
  AOI22_X1 U16050 ( .A1(n13540), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12867), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12800) );
  AOI22_X1 U16051 ( .A1(n13090), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n9825), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12799) );
  AOI22_X1 U16052 ( .A1(n12901), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n11317), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12798) );
  NAND4_X1 U16053 ( .A1(n12801), .A2(n12800), .A3(n12799), .A4(n12798), .ZN(
        n12807) );
  AOI22_X1 U16054 ( .A1(n12978), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n13128), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12805) );
  AOI22_X1 U16055 ( .A1(n12937), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12965), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12804) );
  AOI22_X1 U16056 ( .A1(n13112), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n12964), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12803) );
  AOI22_X1 U16057 ( .A1(n11398), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n13134), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12802) );
  NAND4_X1 U16058 ( .A1(n12805), .A2(n12804), .A3(n12803), .A4(n12802), .ZN(
        n12806) );
  OAI21_X1 U16059 ( .B1(n12807), .B2(n12806), .A(n12838), .ZN(n12812) );
  XOR2_X1 U16060 ( .A(n12809), .B(n12808), .Z(n15770) );
  INV_X1 U16061 ( .A(n15770), .ZN(n12810) );
  AOI22_X1 U16062 ( .A1(n13960), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n13201), .B2(n12810), .ZN(n12811) );
  OAI211_X1 U16063 ( .C1(n12893), .C2(n14295), .A(n12812), .B(n12811), .ZN(
        n14209) );
  NAND2_X1 U16064 ( .A1(n14120), .A2(n14209), .ZN(n12813) );
  AOI22_X1 U16065 ( .A1(n13050), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n13112), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12817) );
  AOI22_X1 U16066 ( .A1(n13090), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12965), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12816) );
  AOI22_X1 U16067 ( .A1(n12978), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12964), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12815) );
  AOI22_X1 U16068 ( .A1(n12901), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n12957), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12814) );
  NAND4_X1 U16069 ( .A1(n12817), .A2(n12816), .A3(n12815), .A4(n12814), .ZN(
        n12823) );
  AOI22_X1 U16070 ( .A1(n11398), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n13128), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12821) );
  AOI22_X1 U16071 ( .A1(n13540), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12867), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12820) );
  AOI22_X1 U16072 ( .A1(n12921), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n13134), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12819) );
  AOI22_X1 U16073 ( .A1(n12937), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n9825), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12818) );
  NAND4_X1 U16074 ( .A1(n12821), .A2(n12820), .A3(n12819), .A4(n12818), .ZN(
        n12822) );
  NOR2_X1 U16075 ( .A1(n12823), .A2(n12822), .ZN(n12828) );
  INV_X1 U16076 ( .A(n12838), .ZN(n12827) );
  XNOR2_X1 U16077 ( .A(n12829), .B(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n14412) );
  NAND2_X1 U16078 ( .A1(n14412), .A2(n13201), .ZN(n12826) );
  AOI22_X1 U16079 ( .A1(n13961), .A2(P1_EAX_REG_14__SCAN_IN), .B1(n13960), 
        .B2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n12825) );
  OAI211_X1 U16080 ( .C1(n12828), .C2(n12827), .A(n12826), .B(n12825), .ZN(
        n14097) );
  XOR2_X1 U16081 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B(n12846), .Z(
        n15760) );
  INV_X1 U16082 ( .A(n15760), .ZN(n12845) );
  AOI22_X1 U16083 ( .A1(n13112), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12921), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12833) );
  AOI22_X1 U16084 ( .A1(n12937), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12901), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12832) );
  AOI22_X1 U16085 ( .A1(n13090), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12867), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12831) );
  AOI22_X1 U16086 ( .A1(n12978), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12964), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12830) );
  NAND4_X1 U16087 ( .A1(n12833), .A2(n12832), .A3(n12831), .A4(n12830), .ZN(
        n12840) );
  AOI22_X1 U16088 ( .A1(n11398), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n13128), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12837) );
  AOI22_X1 U16089 ( .A1(n12965), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13540), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12836) );
  AOI22_X1 U16090 ( .A1(n13050), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n13134), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12835) );
  AOI22_X1 U16091 ( .A1(n12957), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n9825), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12834) );
  NAND4_X1 U16092 ( .A1(n12837), .A2(n12836), .A3(n12835), .A4(n12834), .ZN(
        n12839) );
  OAI21_X1 U16093 ( .B1(n12840), .B2(n12839), .A(n12838), .ZN(n12843) );
  NAND2_X1 U16094 ( .A1(n13961), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n12842) );
  NAND2_X1 U16095 ( .A1(n13960), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12841) );
  NAND3_X1 U16096 ( .A1(n12843), .A2(n12842), .A3(n12841), .ZN(n12844) );
  AOI21_X1 U16097 ( .B1(n12845), .B2(n13201), .A(n12844), .ZN(n14088) );
  INV_X1 U16098 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n12847) );
  XNOR2_X1 U16099 ( .A(n12866), .B(n12847), .ZN(n14077) );
  NAND2_X1 U16100 ( .A1(n14077), .A2(n13201), .ZN(n12864) );
  AOI22_X1 U16101 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n13128), .B1(
        n13090), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12851) );
  AOI22_X1 U16102 ( .A1(n13050), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n13540), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12850) );
  AOI22_X1 U16103 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n12867), .B1(
        n12957), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12849) );
  AOI22_X1 U16104 ( .A1(n12921), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9825), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12848) );
  NAND4_X1 U16105 ( .A1(n12851), .A2(n12850), .A3(n12849), .A4(n12848), .ZN(
        n12860) );
  AOI22_X1 U16106 ( .A1(n13112), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11398), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12857) );
  AOI21_X1 U16107 ( .B1(n12964), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A(
        n13201), .ZN(n12853) );
  NAND2_X1 U16108 ( .A1(n12901), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n12852) );
  AND2_X1 U16109 ( .A1(n12853), .A2(n12852), .ZN(n12856) );
  AOI22_X1 U16110 ( .A1(n12978), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12965), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12855) );
  AOI22_X1 U16111 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n12937), .B1(
        n13134), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12854) );
  NAND4_X1 U16112 ( .A1(n12857), .A2(n12856), .A3(n12855), .A4(n12854), .ZN(
        n12859) );
  NAND2_X1 U16113 ( .A1(n13123), .A2(n12695), .ZN(n12973) );
  OAI21_X1 U16114 ( .B1(n12860), .B2(n12859), .A(n12973), .ZN(n12862) );
  AOI22_X1 U16115 ( .A1(n13961), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n20623), .ZN(n12861) );
  NAND2_X1 U16116 ( .A1(n12862), .A2(n12861), .ZN(n12863) );
  NAND2_X1 U16117 ( .A1(n12864), .A2(n12863), .ZN(n14071) );
  INV_X1 U16118 ( .A(n14071), .ZN(n12865) );
  XOR2_X1 U16119 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B(n12880), .Z(
        n15755) );
  AOI22_X1 U16120 ( .A1(n13961), .A2(P1_EAX_REG_17__SCAN_IN), .B1(n13960), 
        .B2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n12879) );
  AOI22_X1 U16121 ( .A1(n13050), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n13112), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12871) );
  AOI22_X1 U16122 ( .A1(n13540), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12867), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12870) );
  AOI22_X1 U16123 ( .A1(n11398), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n13134), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12869) );
  AOI22_X1 U16124 ( .A1(n12937), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n12957), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12868) );
  NAND4_X1 U16125 ( .A1(n12871), .A2(n12870), .A3(n12869), .A4(n12868), .ZN(
        n12877) );
  AOI22_X1 U16126 ( .A1(n12978), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n13128), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12875) );
  AOI22_X1 U16127 ( .A1(n13090), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12965), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12874) );
  AOI22_X1 U16128 ( .A1(n12921), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12964), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12873) );
  AOI22_X1 U16129 ( .A1(n12901), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n9825), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12872) );
  NAND4_X1 U16130 ( .A1(n12875), .A2(n12874), .A3(n12873), .A4(n12872), .ZN(
        n12876) );
  OAI21_X1 U16131 ( .B1(n12877), .B2(n12876), .A(n13143), .ZN(n12878) );
  OAI211_X1 U16132 ( .C1(n15755), .C2(n12695), .A(n12879), .B(n12878), .ZN(
        n14059) );
  XNOR2_X1 U16133 ( .A(n12912), .B(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14392) );
  AOI22_X1 U16134 ( .A1(n13128), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12937), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12886) );
  NAND2_X1 U16135 ( .A1(n12901), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n12882) );
  NAND2_X1 U16136 ( .A1(n11398), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n12881) );
  AND3_X1 U16137 ( .A1(n12882), .A2(n12881), .A3(n12695), .ZN(n12885) );
  AOI22_X1 U16138 ( .A1(n13112), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n13134), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12884) );
  AOI22_X1 U16139 ( .A1(n13090), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12964), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12883) );
  NAND4_X1 U16140 ( .A1(n12886), .A2(n12885), .A3(n12884), .A4(n12883), .ZN(
        n12892) );
  AOI22_X1 U16141 ( .A1(n12978), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12921), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12890) );
  AOI22_X1 U16142 ( .A1(n12965), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n13540), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12889) );
  AOI22_X1 U16143 ( .A1(n12867), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12957), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12888) );
  AOI22_X1 U16144 ( .A1(n13050), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9825), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12887) );
  NAND4_X1 U16145 ( .A1(n12890), .A2(n12889), .A3(n12888), .A4(n12887), .ZN(
        n12891) );
  OR2_X1 U16146 ( .A1(n12892), .A2(n12891), .ZN(n12895) );
  INV_X1 U16147 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n14276) );
  OAI22_X1 U16148 ( .A1(n12893), .A2(n14276), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n14388), .ZN(n12894) );
  AOI21_X1 U16149 ( .B1(n12973), .B2(n12895), .A(n12894), .ZN(n12896) );
  AOI21_X1 U16150 ( .B1(n14392), .B2(n13201), .A(n12896), .ZN(n14047) );
  AOI22_X1 U16151 ( .A1(n13050), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13112), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12900) );
  AOI22_X1 U16152 ( .A1(n12978), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n13128), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12899) );
  AOI22_X1 U16153 ( .A1(n11398), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n13134), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12898) );
  AOI22_X1 U16154 ( .A1(n12965), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9825), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12897) );
  NAND4_X1 U16155 ( .A1(n12900), .A2(n12899), .A3(n12898), .A4(n12897), .ZN(
        n12907) );
  AOI22_X1 U16156 ( .A1(n12937), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n13090), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12905) );
  AOI22_X1 U16157 ( .A1(n13540), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12867), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12904) );
  AOI22_X1 U16158 ( .A1(n12921), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12964), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12903) );
  AOI22_X1 U16159 ( .A1(n12901), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12957), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12902) );
  NAND4_X1 U16160 ( .A1(n12905), .A2(n12904), .A3(n12903), .A4(n12902), .ZN(
        n12906) );
  NOR2_X1 U16161 ( .A1(n12907), .A2(n12906), .ZN(n12911) );
  OAI21_X1 U16162 ( .B1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n20574), .A(
        n20623), .ZN(n12908) );
  INV_X1 U16163 ( .A(n12908), .ZN(n12909) );
  AOI21_X1 U16164 ( .B1(n13961), .B2(P1_EAX_REG_19__SCAN_IN), .A(n12909), .ZN(
        n12910) );
  OAI21_X1 U16165 ( .B1(n13123), .B2(n12911), .A(n12910), .ZN(n12919) );
  INV_X1 U16166 ( .A(n12952), .ZN(n12917) );
  INV_X1 U16167 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n12915) );
  INV_X1 U16168 ( .A(n12913), .ZN(n12914) );
  NAND2_X1 U16169 ( .A1(n12915), .A2(n12914), .ZN(n12916) );
  NAND2_X1 U16170 ( .A1(n12917), .A2(n12916), .ZN(n15753) );
  NAND2_X1 U16171 ( .A1(n12919), .A2(n12918), .ZN(n14184) );
  AOI22_X1 U16172 ( .A1(n11398), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n13128), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12925) );
  AOI22_X1 U16173 ( .A1(n12978), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n13090), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12924) );
  AOI22_X1 U16174 ( .A1(n12921), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n13134), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12923) );
  AOI22_X1 U16175 ( .A1(n12965), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12957), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12922) );
  NAND4_X1 U16176 ( .A1(n12925), .A2(n12924), .A3(n12923), .A4(n12922), .ZN(
        n12931) );
  AOI22_X1 U16177 ( .A1(n13050), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n13112), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12929) );
  AOI22_X1 U16178 ( .A1(n12937), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n12867), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12928) );
  AOI22_X1 U16179 ( .A1(n13540), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12964), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12927) );
  AOI22_X1 U16180 ( .A1(n12901), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n9825), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12926) );
  NAND4_X1 U16181 ( .A1(n12929), .A2(n12928), .A3(n12927), .A4(n12926), .ZN(
        n12930) );
  NOR2_X1 U16182 ( .A1(n12931), .A2(n12930), .ZN(n12934) );
  INV_X1 U16183 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n15706) );
  AOI21_X1 U16184 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n15706), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12932) );
  AOI21_X1 U16185 ( .B1(n13961), .B2(P1_EAX_REG_20__SCAN_IN), .A(n12932), .ZN(
        n12933) );
  OAI21_X1 U16186 ( .B1(n13123), .B2(n12934), .A(n12933), .ZN(n12936) );
  XNOR2_X1 U16187 ( .A(n12952), .B(n15706), .ZN(n15703) );
  NAND2_X1 U16188 ( .A1(n15703), .A2(n13201), .ZN(n12935) );
  NAND2_X1 U16189 ( .A1(n12936), .A2(n12935), .ZN(n14178) );
  AOI22_X1 U16190 ( .A1(n13112), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n13128), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12941) );
  AOI22_X1 U16191 ( .A1(n12937), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12965), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12940) );
  AOI22_X1 U16192 ( .A1(n13090), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13540), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12939) );
  AOI22_X1 U16193 ( .A1(n12957), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n9825), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12938) );
  NAND4_X1 U16194 ( .A1(n12941), .A2(n12940), .A3(n12939), .A4(n12938), .ZN(
        n12947) );
  AOI22_X1 U16195 ( .A1(n13050), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12921), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12945) );
  AOI22_X1 U16196 ( .A1(n12978), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11398), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12944) );
  AOI22_X1 U16197 ( .A1(n12901), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12867), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12943) );
  AOI22_X1 U16198 ( .A1(n12964), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n13134), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12942) );
  NAND4_X1 U16199 ( .A1(n12945), .A2(n12944), .A3(n12943), .A4(n12942), .ZN(
        n12946) );
  NOR2_X1 U16200 ( .A1(n12947), .A2(n12946), .ZN(n12951) );
  OAI21_X1 U16201 ( .B1(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n20574), .A(
        n20623), .ZN(n12948) );
  INV_X1 U16202 ( .A(n12948), .ZN(n12949) );
  AOI21_X1 U16203 ( .B1(n13961), .B2(P1_EAX_REG_21__SCAN_IN), .A(n12949), .ZN(
        n12950) );
  OAI21_X1 U16204 ( .B1(n13123), .B2(n12951), .A(n12950), .ZN(n12956) );
  AND2_X1 U16205 ( .A1(n12953), .A2(n14373), .ZN(n12954) );
  OR2_X1 U16206 ( .A1(n12954), .A2(n13013), .ZN(n15695) );
  NAND2_X1 U16207 ( .A1(n14375), .A2(n13201), .ZN(n12955) );
  AOI22_X1 U16208 ( .A1(n13112), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n13128), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12963) );
  AOI22_X1 U16209 ( .A1(n11464), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12937), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12962) );
  AOI22_X1 U16210 ( .A1(n13090), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11228), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12961) );
  NAND2_X1 U16211 ( .A1(n11210), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n12959) );
  NAND2_X1 U16212 ( .A1(n12957), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n12958) );
  AND3_X1 U16213 ( .A1(n12959), .A2(n12695), .A3(n12958), .ZN(n12960) );
  NAND4_X1 U16214 ( .A1(n12963), .A2(n12962), .A3(n12961), .A4(n12960), .ZN(
        n12971) );
  AOI22_X1 U16215 ( .A1(n13050), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n13540), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12969) );
  AOI22_X1 U16216 ( .A1(n12867), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12964), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12968) );
  AOI22_X1 U16217 ( .A1(n12965), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n13134), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12967) );
  AOI22_X1 U16218 ( .A1(n12978), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n9825), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12966) );
  NAND4_X1 U16219 ( .A1(n12969), .A2(n12968), .A3(n12967), .A4(n12966), .ZN(
        n12970) );
  OR2_X1 U16220 ( .A1(n12971), .A2(n12970), .ZN(n12972) );
  NAND2_X1 U16221 ( .A1(n12973), .A2(n12972), .ZN(n12977) );
  AOI22_X1 U16222 ( .A1(n13961), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n20623), .ZN(n12976) );
  INV_X1 U16223 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n12974) );
  XNOR2_X1 U16224 ( .A(n13013), .B(n12974), .ZN(n14362) );
  AOI22_X1 U16225 ( .A1(n13050), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n13112), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12982) );
  AOI22_X1 U16226 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n13090), .B1(
        n12937), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12981) );
  AOI22_X1 U16227 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n12978), .B1(
        n13540), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12980) );
  AOI22_X1 U16228 ( .A1(n13128), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11238), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12979) );
  NAND4_X1 U16229 ( .A1(n12982), .A2(n12981), .A3(n12980), .A4(n12979), .ZN(
        n12988) );
  AOI22_X1 U16230 ( .A1(n11398), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12867), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12986) );
  AOI22_X1 U16231 ( .A1(n12921), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12964), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12985) );
  AOI22_X1 U16232 ( .A1(n12901), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11317), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12984) );
  AOI22_X1 U16233 ( .A1(n12965), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n9825), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12983) );
  NAND4_X1 U16234 ( .A1(n12986), .A2(n12985), .A3(n12984), .A4(n12983), .ZN(
        n12987) );
  NOR2_X1 U16235 ( .A1(n12988), .A2(n12987), .ZN(n13017) );
  AOI22_X1 U16236 ( .A1(n11241), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n13112), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12992) );
  AOI22_X1 U16237 ( .A1(n12921), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n13128), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12991) );
  AOI22_X1 U16238 ( .A1(n12937), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12965), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12990) );
  AOI22_X1 U16239 ( .A1(n13090), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n13540), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12989) );
  NAND4_X1 U16240 ( .A1(n12992), .A2(n12991), .A3(n12990), .A4(n12989), .ZN(
        n12998) );
  AOI22_X1 U16241 ( .A1(n11234), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11398), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12996) );
  AOI22_X1 U16242 ( .A1(n12964), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n13134), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12995) );
  AOI22_X1 U16243 ( .A1(n12901), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11317), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12994) );
  AOI22_X1 U16244 ( .A1(n12867), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n9825), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12993) );
  NAND4_X1 U16245 ( .A1(n12996), .A2(n12995), .A3(n12994), .A4(n12993), .ZN(
        n12997) );
  NOR2_X1 U16246 ( .A1(n12998), .A2(n12997), .ZN(n13016) );
  NOR2_X1 U16247 ( .A1(n13017), .A2(n13016), .ZN(n13040) );
  AOI22_X1 U16248 ( .A1(n11241), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n13112), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13002) );
  AOI22_X1 U16249 ( .A1(n13128), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n13540), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n13001) );
  AOI22_X1 U16250 ( .A1(n12921), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12964), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13000) );
  AOI22_X1 U16251 ( .A1(n11398), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n13134), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12999) );
  NAND4_X1 U16252 ( .A1(n13002), .A2(n13001), .A3(n13000), .A4(n12999), .ZN(
        n13008) );
  AOI22_X1 U16253 ( .A1(n12937), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n13090), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13006) );
  AOI22_X1 U16254 ( .A1(n11234), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12867), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13005) );
  AOI22_X1 U16255 ( .A1(n12965), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n9825), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13004) );
  AOI22_X1 U16256 ( .A1(n11228), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12957), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13003) );
  NAND4_X1 U16257 ( .A1(n13006), .A2(n13005), .A3(n13004), .A4(n13003), .ZN(
        n13007) );
  OR2_X1 U16258 ( .A1(n13008), .A2(n13007), .ZN(n13039) );
  XNOR2_X1 U16259 ( .A(n13040), .B(n13039), .ZN(n13012) );
  NAND2_X1 U16260 ( .A1(n20623), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n13009) );
  NAND2_X1 U16261 ( .A1(n12695), .A2(n13009), .ZN(n13010) );
  AOI21_X1 U16262 ( .B1(n13961), .B2(P1_EAX_REG_24__SCAN_IN), .A(n13010), .ZN(
        n13011) );
  OAI21_X1 U16263 ( .B1(n13012), .B2(n13123), .A(n13011), .ZN(n13015) );
  INV_X1 U16264 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n14346) );
  XNOR2_X1 U16265 ( .A(n13044), .B(n14346), .ZN(n14348) );
  NAND2_X1 U16266 ( .A1(n14348), .A2(n13201), .ZN(n13014) );
  NAND2_X1 U16267 ( .A1(n13015), .A2(n13014), .ZN(n14023) );
  XNOR2_X1 U16268 ( .A(n13017), .B(n13016), .ZN(n13021) );
  INV_X1 U16269 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n13018) );
  AOI21_X1 U16270 ( .B1(n13018), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n13019) );
  AOI21_X1 U16271 ( .B1(n12673), .B2(P1_EAX_REG_23__SCAN_IN), .A(n13019), .ZN(
        n13020) );
  OAI21_X1 U16272 ( .B1(n13123), .B2(n13021), .A(n13020), .ZN(n13026) );
  NOR2_X1 U16273 ( .A1(n13022), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n13023) );
  OR2_X1 U16274 ( .A1(n13044), .A2(n13023), .ZN(n15688) );
  INV_X1 U16275 ( .A(n15688), .ZN(n13024) );
  NAND2_X1 U16276 ( .A1(n13024), .A2(n13201), .ZN(n13025) );
  NAND2_X1 U16277 ( .A1(n13026), .A2(n13025), .ZN(n14170) );
  AOI22_X1 U16278 ( .A1(n11398), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n13128), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13032) );
  AOI22_X1 U16279 ( .A1(n12937), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12867), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n13031) );
  AOI22_X1 U16280 ( .A1(n13112), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11238), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13030) );
  AOI22_X1 U16281 ( .A1(n12965), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n9825), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13029) );
  NAND4_X1 U16282 ( .A1(n13032), .A2(n13031), .A3(n13030), .A4(n13029), .ZN(
        n13038) );
  AOI22_X1 U16283 ( .A1(n11241), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12921), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n13036) );
  AOI22_X1 U16284 ( .A1(n11234), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n13090), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n13035) );
  AOI22_X1 U16285 ( .A1(n13540), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12964), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13034) );
  AOI22_X1 U16286 ( .A1(n11228), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11317), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13033) );
  NAND4_X1 U16287 ( .A1(n13036), .A2(n13035), .A3(n13034), .A4(n13033), .ZN(
        n13037) );
  NOR2_X1 U16288 ( .A1(n13038), .A2(n13037), .ZN(n13062) );
  NAND2_X1 U16289 ( .A1(n13040), .A2(n13039), .ZN(n13061) );
  XNOR2_X1 U16290 ( .A(n13062), .B(n13061), .ZN(n13043) );
  INV_X1 U16291 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n14337) );
  OAI21_X1 U16292 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n14337), .A(n12695), 
        .ZN(n13041) );
  AOI21_X1 U16293 ( .B1(n12673), .B2(P1_EAX_REG_25__SCAN_IN), .A(n13041), .ZN(
        n13042) );
  OAI21_X1 U16294 ( .B1(n13043), .B2(n13123), .A(n13042), .ZN(n13048) );
  NAND2_X1 U16295 ( .A1(n13045), .A2(n14337), .ZN(n13046) );
  NAND2_X1 U16296 ( .A1(n14341), .A2(n13201), .ZN(n13047) );
  NAND2_X1 U16297 ( .A1(n13048), .A2(n13047), .ZN(n14005) );
  AOI22_X1 U16298 ( .A1(n13050), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n13112), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13054) );
  AOI22_X1 U16299 ( .A1(n13128), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n13540), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n13053) );
  AOI22_X1 U16300 ( .A1(n12921), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12964), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13052) );
  AOI22_X1 U16301 ( .A1(n11398), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n13134), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13051) );
  NAND4_X1 U16302 ( .A1(n13054), .A2(n13053), .A3(n13052), .A4(n13051), .ZN(
        n13060) );
  AOI22_X1 U16303 ( .A1(n11232), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n13090), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13058) );
  AOI22_X1 U16304 ( .A1(n11234), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12867), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13057) );
  AOI22_X1 U16305 ( .A1(n12965), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n9825), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13056) );
  AOI22_X1 U16306 ( .A1(n11228), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12957), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13055) );
  NAND4_X1 U16307 ( .A1(n13058), .A2(n13057), .A3(n13056), .A4(n13055), .ZN(
        n13059) );
  OR2_X1 U16308 ( .A1(n13060), .A2(n13059), .ZN(n13080) );
  NOR2_X1 U16309 ( .A1(n13062), .A2(n13061), .ZN(n13081) );
  XOR2_X1 U16310 ( .A(n13080), .B(n13081), .Z(n13063) );
  NAND2_X1 U16311 ( .A1(n13063), .A2(n13143), .ZN(n13066) );
  INV_X1 U16312 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n15672) );
  NOR2_X1 U16313 ( .A1(n15672), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13064) );
  AOI211_X1 U16314 ( .C1(n12673), .C2(P1_EAX_REG_26__SCAN_IN), .A(n13201), .B(
        n13064), .ZN(n13065) );
  XNOR2_X1 U16315 ( .A(n13067), .B(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15678) );
  AOI22_X1 U16316 ( .A1(n13066), .A2(n13065), .B1(n13201), .B2(n15678), .ZN(
        n14156) );
  NOR2_X1 U16317 ( .A1(n13068), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n13069) );
  AOI22_X1 U16318 ( .A1(n11241), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12921), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n13073) );
  AOI22_X1 U16319 ( .A1(n13128), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n13540), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n13072) );
  AOI22_X1 U16320 ( .A1(n11398), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12964), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13071) );
  AOI22_X1 U16321 ( .A1(n11228), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12957), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13070) );
  NAND4_X1 U16322 ( .A1(n13073), .A2(n13072), .A3(n13071), .A4(n13070), .ZN(
        n13079) );
  AOI22_X1 U16323 ( .A1(n12937), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n13090), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n13077) );
  AOI22_X1 U16324 ( .A1(n11234), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12867), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n13076) );
  AOI22_X1 U16325 ( .A1(n13112), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n13134), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13075) );
  AOI22_X1 U16326 ( .A1(n12965), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n9825), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13074) );
  NAND4_X1 U16327 ( .A1(n13077), .A2(n13076), .A3(n13075), .A4(n13074), .ZN(
        n13078) );
  NOR2_X1 U16328 ( .A1(n13079), .A2(n13078), .ZN(n13098) );
  NAND2_X1 U16329 ( .A1(n13081), .A2(n13080), .ZN(n13097) );
  XNOR2_X1 U16330 ( .A(n13098), .B(n13097), .ZN(n13084) );
  AOI21_X1 U16331 ( .B1(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n20623), .A(
        n13201), .ZN(n13083) );
  NAND2_X1 U16332 ( .A1(n13961), .A2(P1_EAX_REG_27__SCAN_IN), .ZN(n13082) );
  OAI211_X1 U16333 ( .C1(n13084), .C2(n13123), .A(n13083), .B(n13082), .ZN(
        n13085) );
  AOI22_X1 U16334 ( .A1(n11241), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13133), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13089) );
  AOI22_X1 U16335 ( .A1(n13128), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13540), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13088) );
  INV_X1 U16336 ( .A(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n20952) );
  AOI22_X1 U16337 ( .A1(n11210), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12964), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13087) );
  AOI22_X1 U16338 ( .A1(n11464), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n13134), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13086) );
  NAND4_X1 U16339 ( .A1(n13089), .A2(n13088), .A3(n13087), .A4(n13086), .ZN(
        n13096) );
  AOI22_X1 U16340 ( .A1(n11232), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n13090), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13094) );
  AOI22_X1 U16341 ( .A1(n11234), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12867), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13093) );
  AOI22_X1 U16342 ( .A1(n12965), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n9825), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13092) );
  AOI22_X1 U16343 ( .A1(n11228), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12957), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13091) );
  NAND4_X1 U16344 ( .A1(n13094), .A2(n13093), .A3(n13092), .A4(n13091), .ZN(
        n13095) );
  OR2_X1 U16345 ( .A1(n13096), .A2(n13095), .ZN(n13119) );
  NOR2_X1 U16346 ( .A1(n13098), .A2(n13097), .ZN(n13120) );
  XOR2_X1 U16347 ( .A(n13119), .B(n13120), .Z(n13099) );
  NAND2_X1 U16348 ( .A1(n13099), .A2(n13143), .ZN(n13102) );
  INV_X1 U16349 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n15653) );
  NOR2_X1 U16350 ( .A1(n15653), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13100) );
  AOI211_X1 U16351 ( .C1(n12673), .C2(P1_EAX_REG_28__SCAN_IN), .A(n13201), .B(
        n13100), .ZN(n13101) );
  XOR2_X1 U16352 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B(n13103), .Z(
        n15651) );
  AOI22_X1 U16353 ( .A1(n13102), .A2(n13101), .B1(n13201), .B2(n15651), .ZN(
        n13170) );
  INV_X1 U16354 ( .A(n13105), .ZN(n13106) );
  INV_X1 U16355 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n21083) );
  NAND2_X1 U16356 ( .A1(n13106), .A2(n21083), .ZN(n13107) );
  NAND2_X1 U16357 ( .A1(n13205), .A2(n13107), .ZN(n14313) );
  AOI22_X1 U16358 ( .A1(n11464), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n13128), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13111) );
  AOI22_X1 U16359 ( .A1(n11234), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12965), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13110) );
  AOI22_X1 U16360 ( .A1(n11210), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n13134), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13109) );
  AOI22_X1 U16361 ( .A1(n11228), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n9825), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13108) );
  NAND4_X1 U16362 ( .A1(n13111), .A2(n13110), .A3(n13109), .A4(n13108), .ZN(
        n13118) );
  AOI22_X1 U16363 ( .A1(n11241), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n13112), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13116) );
  AOI22_X1 U16364 ( .A1(n13090), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12867), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n13115) );
  AOI22_X1 U16365 ( .A1(n13540), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12964), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13114) );
  AOI22_X1 U16366 ( .A1(n11232), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12957), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13113) );
  NAND4_X1 U16367 ( .A1(n13116), .A2(n13115), .A3(n13114), .A4(n13113), .ZN(
        n13117) );
  NOR2_X1 U16368 ( .A1(n13118), .A2(n13117), .ZN(n13127) );
  NAND2_X1 U16369 ( .A1(n13120), .A2(n13119), .ZN(n13126) );
  XNOR2_X1 U16370 ( .A(n13127), .B(n13126), .ZN(n13124) );
  NOR2_X1 U16371 ( .A1(n21083), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13121) );
  AOI211_X1 U16372 ( .C1(n12673), .C2(P1_EAX_REG_29__SCAN_IN), .A(n13201), .B(
        n13121), .ZN(n13122) );
  OAI21_X1 U16373 ( .B1(n13124), .B2(n13123), .A(n13122), .ZN(n13125) );
  OAI21_X1 U16374 ( .B1(n12695), .B2(n14313), .A(n13125), .ZN(n13996) );
  NOR2_X1 U16375 ( .A1(n13127), .A2(n13126), .ZN(n13142) );
  AOI22_X1 U16376 ( .A1(n13128), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n13540), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n13132) );
  AOI22_X1 U16377 ( .A1(n11464), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12964), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13131) );
  AOI22_X1 U16378 ( .A1(n11228), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12957), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13130) );
  AOI22_X1 U16379 ( .A1(n13090), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n9825), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13129) );
  NAND4_X1 U16380 ( .A1(n13132), .A2(n13131), .A3(n13130), .A4(n13129), .ZN(
        n13140) );
  AOI22_X1 U16381 ( .A1(n11241), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13133), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13138) );
  AOI22_X1 U16382 ( .A1(n11232), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12965), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13137) );
  AOI22_X1 U16383 ( .A1(n12978), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12867), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n13136) );
  AOI22_X1 U16384 ( .A1(n11210), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n13134), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13135) );
  NAND4_X1 U16385 ( .A1(n13138), .A2(n13137), .A3(n13136), .A4(n13135), .ZN(
        n13139) );
  NOR2_X1 U16386 ( .A1(n13140), .A2(n13139), .ZN(n13141) );
  XNOR2_X1 U16387 ( .A(n13142), .B(n13141), .ZN(n13144) );
  NAND2_X1 U16388 ( .A1(n13144), .A2(n13143), .ZN(n13149) );
  NAND2_X1 U16389 ( .A1(n20623), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13145) );
  NAND2_X1 U16390 ( .A1(n12695), .A2(n13145), .ZN(n13146) );
  AOI21_X1 U16391 ( .B1(n12673), .B2(P1_EAX_REG_30__SCAN_IN), .A(n13146), .ZN(
        n13148) );
  XNOR2_X1 U16392 ( .A(n13205), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14306) );
  AOI21_X1 U16393 ( .B1(n13149), .B2(n13148), .A(n13147), .ZN(n13959) );
  NAND2_X1 U16394 ( .A1(n13466), .A2(n13445), .ZN(n13462) );
  NAND3_X1 U16395 ( .A1(n13151), .A2(n13965), .A3(n20136), .ZN(n13699) );
  INV_X1 U16396 ( .A(n13699), .ZN(n13152) );
  NAND3_X1 U16397 ( .A1(n13153), .A2(n13696), .A3(n13152), .ZN(n13154) );
  NAND2_X1 U16398 ( .A1(n13462), .A2(n13154), .ZN(n13155) );
  INV_X1 U16399 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n13157) );
  INV_X1 U16400 ( .A(n14354), .ZN(n14332) );
  NOR2_X2 U16401 ( .A1(n14332), .A2(n13161), .ZN(n13164) );
  NOR3_X1 U16402 ( .A1(n14352), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n13162), .ZN(n13163) );
  AOI21_X1 U16403 ( .B1(n13164), .B2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n13163), .ZN(n14320) );
  NAND2_X1 U16404 ( .A1(n14446), .A2(n20046), .ZN(n13180) );
  NAND2_X1 U16405 ( .A1(n20098), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n15931) );
  NAND2_X1 U16406 ( .A1(P1_STATEBS16_REG_SCAN_IN), .A2(n20765), .ZN(n20544) );
  NAND2_X1 U16407 ( .A1(n13173), .A2(n20632), .ZN(n20786) );
  AND2_X1 U16408 ( .A1(n20786), .A2(n20098), .ZN(n13174) );
  NOR2_X1 U16409 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n20623), .ZN(n20788) );
  AOI21_X1 U16410 ( .B1(n20574), .B2(P1_STATE2_REG_1__SCAN_IN), .A(n20788), 
        .ZN(n13411) );
  INV_X1 U16411 ( .A(n13411), .ZN(n13175) );
  NOR2_X1 U16412 ( .A1(n20081), .A2(n15645), .ZN(n14440) );
  NOR2_X1 U16413 ( .A1(n14425), .A2(n15653), .ZN(n13176) );
  AOI211_X1 U16414 ( .C1(n20045), .C2(n15651), .A(n14440), .B(n13176), .ZN(
        n13177) );
  NAND2_X1 U16415 ( .A1(n13180), .A2(n13179), .ZN(P1_U2971) );
  NOR2_X1 U16416 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(P2_BE_N_REG_1__SCAN_IN), 
        .ZN(n13182) );
  NOR4_X1 U16417 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n13181) );
  NAND4_X1 U16418 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(P2_W_R_N_REG_SCAN_IN), 
        .A3(n13182), .A4(n13181), .ZN(n13195) );
  NOR4_X1 U16419 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(
        P1_ADDRESS_REG_14__SCAN_IN), .A3(P1_ADDRESS_REG_13__SCAN_IN), .A4(
        P1_ADDRESS_REG_12__SCAN_IN), .ZN(n13186) );
  NOR4_X1 U16420 ( .A1(P1_ADDRESS_REG_21__SCAN_IN), .A2(
        P1_ADDRESS_REG_19__SCAN_IN), .A3(P1_ADDRESS_REG_18__SCAN_IN), .A4(
        P1_ADDRESS_REG_16__SCAN_IN), .ZN(n13185) );
  NOR4_X1 U16421 ( .A1(P1_ADDRESS_REG_7__SCAN_IN), .A2(
        P1_ADDRESS_REG_6__SCAN_IN), .A3(P1_ADDRESS_REG_5__SCAN_IN), .A4(
        P1_ADDRESS_REG_4__SCAN_IN), .ZN(n13184) );
  NOR4_X1 U16422 ( .A1(P1_ADDRESS_REG_11__SCAN_IN), .A2(
        P1_ADDRESS_REG_10__SCAN_IN), .A3(P1_ADDRESS_REG_9__SCAN_IN), .A4(
        P1_ADDRESS_REG_8__SCAN_IN), .ZN(n13183) );
  AND4_X1 U16423 ( .A1(n13186), .A2(n13185), .A3(n13184), .A4(n13183), .ZN(
        n13191) );
  NOR4_X1 U16424 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(
        P1_ADDRESS_REG_0__SCAN_IN), .A3(P1_ADDRESS_REG_20__SCAN_IN), .A4(
        P1_ADDRESS_REG_17__SCAN_IN), .ZN(n13189) );
  NOR4_X1 U16425 ( .A1(P1_ADDRESS_REG_25__SCAN_IN), .A2(
        P1_ADDRESS_REG_24__SCAN_IN), .A3(P1_ADDRESS_REG_23__SCAN_IN), .A4(
        P1_ADDRESS_REG_22__SCAN_IN), .ZN(n13188) );
  NOR4_X1 U16426 ( .A1(P1_ADDRESS_REG_2__SCAN_IN), .A2(
        P1_ADDRESS_REG_28__SCAN_IN), .A3(P1_ADDRESS_REG_27__SCAN_IN), .A4(
        P1_ADDRESS_REG_26__SCAN_IN), .ZN(n13187) );
  INV_X1 U16427 ( .A(P1_ADDRESS_REG_3__SCAN_IN), .ZN(n20711) );
  AND4_X1 U16428 ( .A1(n13189), .A2(n13188), .A3(n13187), .A4(n20711), .ZN(
        n13190) );
  NAND2_X1 U16429 ( .A1(n13191), .A2(n13190), .ZN(n13192) );
  NOR3_X1 U16430 ( .A1(P1_BE_N_REG_3__SCAN_IN), .A2(P1_ADS_N_REG_SCAN_IN), 
        .A3(P1_BE_N_REG_1__SCAN_IN), .ZN(n13194) );
  INV_X1 U16431 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n20784) );
  NOR4_X1 U16432 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_0__SCAN_IN), 
        .A3(P1_D_C_N_REG_SCAN_IN), .A4(n20784), .ZN(n13193) );
  NAND4_X1 U16433 ( .A1(n20092), .A2(P1_M_IO_N_REG_SCAN_IN), .A3(n13194), .A4(
        n13193), .ZN(U214) );
  NOR2_X1 U16434 ( .A1(n14769), .A2(n13195), .ZN(n16317) );
  NAND2_X1 U16435 ( .A1(n16317), .A2(U214), .ZN(U212) );
  AOI21_X1 U16436 ( .B1(n13199), .B2(n13196), .A(n12785), .ZN(n14436) );
  INV_X1 U16437 ( .A(n14436), .ZN(n13935) );
  NOR2_X1 U16438 ( .A1(n11716), .A2(n19861), .ZN(n13200) );
  INV_X1 U16439 ( .A(n13282), .ZN(n13274) );
  NAND3_X1 U16440 ( .A1(n11598), .A2(n13703), .A3(n13274), .ZN(n13260) );
  NAND2_X1 U16441 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n20623), .ZN(n15930) );
  NAND2_X1 U16442 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n15937), .ZN(n15615) );
  INV_X1 U16443 ( .A(n15931), .ZN(n13202) );
  NAND2_X1 U16444 ( .A1(n13202), .A2(n13201), .ZN(n13203) );
  OAI211_X1 U16445 ( .C1(n15930), .C2(n15615), .A(n20081), .B(n13203), .ZN(
        n13204) );
  INV_X1 U16446 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n14303) );
  INV_X1 U16447 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n13206) );
  NOR2_X1 U16448 ( .A1(n13973), .A2(n15937), .ZN(n13208) );
  NOR2_X1 U16449 ( .A1(n13935), .A2(n15726), .ZN(n13231) );
  NAND2_X1 U16450 ( .A1(n20697), .A2(n20574), .ZN(n13210) );
  INV_X1 U16451 ( .A(n13210), .ZN(n13217) );
  AND3_X1 U16452 ( .A1(n13218), .A2(n13217), .A3(n9823), .ZN(n13209) );
  INV_X1 U16453 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n15901) );
  NAND4_X1 U16454 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(P1_REIP_REG_3__SCAN_IN), 
        .A3(P1_REIP_REG_1__SCAN_IN), .A4(P1_REIP_REG_2__SCAN_IN), .ZN(n19923)
         );
  NAND3_X1 U16455 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(P1_REIP_REG_6__SCAN_IN), 
        .A3(P1_REIP_REG_5__SCAN_IN), .ZN(n14131) );
  NOR3_X1 U16456 ( .A1(n15901), .A2(n19923), .A3(n14131), .ZN(n19885) );
  NAND2_X1 U16457 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(n19885), .ZN(n13222) );
  NOR3_X1 U16458 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(n19926), .A3(n13222), 
        .ZN(n13230) );
  NAND2_X1 U16459 ( .A1(n13210), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n13211) );
  NOR2_X1 U16460 ( .A1(n13276), .A2(n13211), .ZN(n13212) );
  NAND2_X1 U16461 ( .A1(n15886), .A2(n13213), .ZN(n13214) );
  NAND2_X1 U16462 ( .A1(n14217), .A2(n13214), .ZN(n15879) );
  INV_X1 U16463 ( .A(n15879), .ZN(n13215) );
  AND2_X1 U16464 ( .A1(n19948), .A2(n13215), .ZN(n13229) );
  INV_X1 U16465 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n14143) );
  NAND2_X1 U16466 ( .A1(n13218), .A2(n13217), .ZN(n13219) );
  OAI211_X1 U16467 ( .C1(n9787), .C2(n14143), .A(n13219), .B(n9823), .ZN(
        n13220) );
  INV_X1 U16468 ( .A(n13220), .ZN(n13221) );
  NAND2_X1 U16469 ( .A1(n19937), .A2(P1_EBX_REG_10__SCAN_IN), .ZN(n13227) );
  INV_X1 U16470 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n13223) );
  NOR2_X1 U16471 ( .A1(n13223), .A2(n13222), .ZN(n15720) );
  OAI21_X1 U16472 ( .B1(n15720), .B2(n19926), .A(n19924), .ZN(n15732) );
  NOR2_X1 U16473 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20632), .ZN(n13290) );
  NAND2_X1 U16474 ( .A1(n19924), .A2(n13290), .ZN(n19942) );
  OAI21_X1 U16475 ( .B1(n15730), .B2(n13224), .A(n19942), .ZN(n13225) );
  AOI21_X1 U16476 ( .B1(P1_REIP_REG_10__SCAN_IN), .B2(n15732), .A(n13225), 
        .ZN(n13226) );
  OAI211_X1 U16477 ( .C1(n14434), .C2(n19957), .A(n13227), .B(n13226), .ZN(
        n13228) );
  NAND2_X1 U16478 ( .A1(n13233), .A2(n13232), .ZN(n13236) );
  INV_X1 U16479 ( .A(n13234), .ZN(n13235) );
  AND2_X1 U16480 ( .A1(n13236), .A2(n13235), .ZN(n19797) );
  OAI22_X1 U16481 ( .A1(n19797), .A2(n21133), .B1(n13240), .B2(n13237), .ZN(
        n13252) );
  INV_X1 U16482 ( .A(n13238), .ZN(n13239) );
  NAND3_X1 U16483 ( .A1(n13241), .A2(n13240), .A3(n13239), .ZN(n13243) );
  NAND2_X1 U16484 ( .A1(n18976), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n13321) );
  NAND3_X1 U16485 ( .A1(n13243), .A2(n13242), .A3(n13321), .ZN(n13251) );
  OAI22_X1 U16486 ( .A1(n10599), .A2(n15360), .B1(n15356), .B2(n13244), .ZN(
        n13250) );
  XNOR2_X1 U16487 ( .A(n13246), .B(n13245), .ZN(n13327) );
  XNOR2_X1 U16488 ( .A(n13248), .B(n13247), .ZN(n13322) );
  OAI22_X1 U16489 ( .A1(n13327), .A2(n21140), .B1(n16157), .B2(n13322), .ZN(
        n13249) );
  OR4_X1 U16490 ( .A1(n13252), .A2(n13251), .A3(n13250), .A4(n13249), .ZN(
        P2_U3044) );
  INV_X1 U16491 ( .A(n15544), .ZN(n16226) );
  NAND2_X1 U16492 ( .A1(n16226), .A2(n13253), .ZN(n14652) );
  INV_X1 U16493 ( .A(n14652), .ZN(n18998) );
  INV_X1 U16494 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n13255) );
  INV_X1 U16495 ( .A(n13253), .ZN(n13254) );
  OAI211_X1 U16496 ( .C1(n18998), .C2(n13255), .A(n13256), .B(n13269), .ZN(
        P2_U2814) );
  INV_X1 U16497 ( .A(n13256), .ZN(n13257) );
  OAI21_X1 U16498 ( .B1(P2_READREQUEST_REG_SCAN_IN), .B2(n13257), .A(n19838), 
        .ZN(n13258) );
  OAI21_X1 U16499 ( .B1(n13259), .B2(n19838), .A(n13258), .ZN(P2_U3612) );
  AOI21_X1 U16500 ( .B1(n13260), .B2(P1_MEMORYFETCH_REG_SCAN_IN), .A(n13290), 
        .ZN(n13261) );
  NAND2_X1 U16501 ( .A1(n13528), .A2(n13261), .ZN(P1_U2801) );
  XNOR2_X1 U16502 ( .A(n18995), .B(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n15362) );
  AOI21_X1 U16503 ( .B1(n10124), .B2(n13263), .A(n13262), .ZN(n15364) );
  INV_X1 U16504 ( .A(n15364), .ZN(n13264) );
  NAND2_X1 U16505 ( .A1(n18976), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n15358) );
  OAI21_X1 U16506 ( .B1(n16055), .B2(n13264), .A(n15358), .ZN(n13265) );
  AOI21_X1 U16507 ( .B1(n16118), .B2(n15362), .A(n13265), .ZN(n13268) );
  OAI21_X1 U16508 ( .B1(n16062), .B2(n13266), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13267) );
  OAI211_X1 U16509 ( .C1(n16088), .C2(n15359), .A(n13268), .B(n13267), .ZN(
        P2_U3014) );
  INV_X1 U16510 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n13273) );
  NOR2_X2 U16511 ( .A1(n13269), .A2(n9779), .ZN(n19143) );
  NOR2_X1 U16512 ( .A1(n13269), .A2(n19844), .ZN(n13270) );
  OR2_X1 U16513 ( .A1(n19143), .A2(n13270), .ZN(n13294) );
  INV_X1 U16514 ( .A(n19139), .ZN(n13272) );
  AOI22_X1 U16515 ( .A1(n13781), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n14769), .ZN(n13814) );
  INV_X1 U16516 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n13271) );
  OAI222_X1 U16517 ( .A1(n13273), .A2(n13294), .B1(n13272), .B2(n13814), .C1(
        n13271), .C2(n13344), .ZN(P2_U2982) );
  INV_X1 U16518 ( .A(n11716), .ZN(n13421) );
  AOI21_X1 U16519 ( .B1(n11598), .B2(n13274), .A(n13421), .ZN(n13275) );
  AOI21_X1 U16520 ( .B1(n13466), .B2(n13277), .A(n13275), .ZN(n19860) );
  NAND3_X1 U16521 ( .A1(n13277), .A2(n13276), .A3(n15631), .ZN(n13278) );
  NAND2_X1 U16522 ( .A1(n13278), .A2(n20697), .ZN(n20789) );
  NAND2_X1 U16523 ( .A1(n19860), .A2(n20789), .ZN(n15603) );
  AND2_X1 U16524 ( .A1(n15603), .A2(n13703), .ZN(n19869) );
  INV_X1 U16525 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n13289) );
  INV_X1 U16526 ( .A(n13445), .ZN(n13285) );
  NAND2_X1 U16527 ( .A1(n13280), .A2(n13279), .ZN(n13281) );
  NAND2_X1 U16528 ( .A1(n13466), .A2(n13281), .ZN(n13284) );
  NAND2_X1 U16529 ( .A1(n11598), .A2(n13282), .ZN(n13283) );
  OAI211_X1 U16530 ( .C1(n13466), .C2(n13285), .A(n13284), .B(n13283), .ZN(
        n13286) );
  NAND2_X1 U16531 ( .A1(n13286), .A2(n11253), .ZN(n15599) );
  INV_X1 U16532 ( .A(n15599), .ZN(n13287) );
  NAND2_X1 U16533 ( .A1(n19869), .A2(n13287), .ZN(n13288) );
  OAI21_X1 U16534 ( .B1(n19869), .B2(n13289), .A(n13288), .ZN(P1_U3484) );
  INV_X1 U16535 ( .A(n20785), .ZN(n13292) );
  OAI21_X1 U16536 ( .B1(n13290), .B2(P1_READREQUEST_REG_SCAN_IN), .A(n13292), 
        .ZN(n13291) );
  OAI21_X1 U16537 ( .B1(n13293), .B2(n13292), .A(n13291), .ZN(P1_U3487) );
  INV_X2 U16538 ( .A(n13294), .ZN(n13338) );
  AOI22_X1 U16539 ( .A1(n13338), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(
        P2_EAX_REG_27__SCAN_IN), .B2(n19143), .ZN(n13298) );
  INV_X1 U16540 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n13295) );
  OR2_X1 U16541 ( .A1(n14769), .A2(n13295), .ZN(n13297) );
  NAND2_X1 U16542 ( .A1(n14769), .A2(BUF2_REG_11__SCAN_IN), .ZN(n13296) );
  NAND2_X1 U16543 ( .A1(n13297), .A2(n13296), .ZN(n14785) );
  NAND2_X1 U16544 ( .A1(n19139), .A2(n14785), .ZN(n13366) );
  NAND2_X1 U16545 ( .A1(n13298), .A2(n13366), .ZN(P2_U2963) );
  AOI22_X1 U16546 ( .A1(n13338), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(
        P2_EAX_REG_0__SCAN_IN), .B2(n19143), .ZN(n13300) );
  AOI22_X1 U16547 ( .A1(n13781), .A2(BUF1_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n14769), .ZN(n19092) );
  INV_X1 U16548 ( .A(n19092), .ZN(n13299) );
  NAND2_X1 U16549 ( .A1(n19139), .A2(n13299), .ZN(n13362) );
  NAND2_X1 U16550 ( .A1(n13300), .A2(n13362), .ZN(P2_U2967) );
  AOI22_X1 U16551 ( .A1(n13338), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19136), 
        .B2(P2_EAX_REG_21__SCAN_IN), .ZN(n13301) );
  AOI22_X1 U16552 ( .A1(n13781), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n14769), .ZN(n19171) );
  INV_X1 U16553 ( .A(n19171), .ZN(n19054) );
  NAND2_X1 U16554 ( .A1(n19139), .A2(n19054), .ZN(n13370) );
  NAND2_X1 U16555 ( .A1(n13301), .A2(n13370), .ZN(P2_U2957) );
  AOI22_X1 U16556 ( .A1(n13338), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(
        P2_EAX_REG_20__SCAN_IN), .B2(n19143), .ZN(n13302) );
  INV_X1 U16557 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n16363) );
  INV_X1 U16558 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n18129) );
  AOI22_X1 U16559 ( .A1(n13781), .A2(n16363), .B1(n18129), .B2(n14769), .ZN(
        n19062) );
  NAND2_X1 U16560 ( .A1(n19139), .A2(n19062), .ZN(n13308) );
  NAND2_X1 U16561 ( .A1(n13302), .A2(n13308), .ZN(P2_U2956) );
  AOI22_X1 U16562 ( .A1(n13338), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19136), 
        .B2(P2_EAX_REG_1__SCAN_IN), .ZN(n13304) );
  AOI22_X1 U16563 ( .A1(n13781), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n14769), .ZN(n19158) );
  INV_X1 U16564 ( .A(n19158), .ZN(n13303) );
  NAND2_X1 U16565 ( .A1(n19139), .A2(n13303), .ZN(n13368) );
  NAND2_X1 U16566 ( .A1(n13304), .A2(n13368), .ZN(P2_U2968) );
  AOI22_X1 U16567 ( .A1(n13338), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(
        P2_EAX_REG_25__SCAN_IN), .B2(n19143), .ZN(n13305) );
  MUX2_X1 U16568 ( .A(BUF1_REG_9__SCAN_IN), .B(BUF2_REG_9__SCAN_IN), .S(n14769), .Z(n14802) );
  NAND2_X1 U16569 ( .A1(n19139), .A2(n14802), .ZN(n13358) );
  NAND2_X1 U16570 ( .A1(n13305), .A2(n13358), .ZN(P2_U2961) );
  AOI22_X1 U16571 ( .A1(n13338), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(
        P2_EAX_REG_24__SCAN_IN), .B2(n19143), .ZN(n13307) );
  AOI22_X1 U16572 ( .A1(n13781), .A2(BUF1_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n14769), .ZN(n14811) );
  INV_X1 U16573 ( .A(n14811), .ZN(n13306) );
  NAND2_X1 U16574 ( .A1(n19139), .A2(n13306), .ZN(n13364) );
  NAND2_X1 U16575 ( .A1(n13307), .A2(n13364), .ZN(P2_U2960) );
  AOI22_X1 U16576 ( .A1(n13338), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(
        P2_EAX_REG_4__SCAN_IN), .B2(n19143), .ZN(n13309) );
  NAND2_X1 U16577 ( .A1(n13309), .A2(n13308), .ZN(P2_U2971) );
  AOI22_X1 U16578 ( .A1(n13338), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(
        P2_EAX_REG_29__SCAN_IN), .B2(n19143), .ZN(n13312) );
  INV_X1 U16579 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n14229) );
  OR2_X1 U16580 ( .A1(n14769), .A2(n14229), .ZN(n13311) );
  NAND2_X1 U16581 ( .A1(n14769), .A2(BUF2_REG_13__SCAN_IN), .ZN(n13310) );
  NAND2_X1 U16582 ( .A1(n13311), .A2(n13310), .ZN(n14765) );
  NAND2_X1 U16583 ( .A1(n19139), .A2(n14765), .ZN(n13316) );
  NAND2_X1 U16584 ( .A1(n13312), .A2(n13316), .ZN(P2_U2965) );
  AOI22_X1 U16585 ( .A1(n13338), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19143), 
        .B2(P2_EAX_REG_23__SCAN_IN), .ZN(n13314) );
  AOI22_X1 U16586 ( .A1(n13781), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n14769), .ZN(n19181) );
  INV_X1 U16587 ( .A(n19181), .ZN(n13313) );
  NAND2_X1 U16588 ( .A1(n19139), .A2(n13313), .ZN(n13356) );
  NAND2_X1 U16589 ( .A1(n13314), .A2(n13356), .ZN(P2_U2959) );
  AOI22_X1 U16590 ( .A1(n13338), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(
        P2_EAX_REG_22__SCAN_IN), .B2(n19136), .ZN(n13315) );
  INV_X1 U16591 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n16359) );
  INV_X1 U16592 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n18139) );
  AOI22_X1 U16593 ( .A1(n13781), .A2(n16359), .B1(n18139), .B2(n14769), .ZN(
        n16033) );
  NAND2_X1 U16594 ( .A1(n19139), .A2(n16033), .ZN(n13352) );
  NAND2_X1 U16595 ( .A1(n13315), .A2(n13352), .ZN(P2_U2958) );
  AOI22_X1 U16596 ( .A1(n13338), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(
        P2_EAX_REG_13__SCAN_IN), .B2(n19143), .ZN(n13317) );
  NAND2_X1 U16597 ( .A1(n13317), .A2(n13316), .ZN(P2_U2980) );
  AOI22_X1 U16598 ( .A1(n13338), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(
        P2_EAX_REG_2__SCAN_IN), .B2(n19143), .ZN(n13318) );
  OAI22_X1 U16599 ( .A1(n14769), .A2(BUF1_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n13781), .ZN(n19161) );
  INV_X1 U16600 ( .A(n19161), .ZN(n16046) );
  NAND2_X1 U16601 ( .A1(n19139), .A2(n16046), .ZN(n13360) );
  NAND2_X1 U16602 ( .A1(n13318), .A2(n13360), .ZN(P2_U2969) );
  AOI22_X1 U16603 ( .A1(n13338), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(
        P2_EAX_REG_3__SCAN_IN), .B2(n19143), .ZN(n13320) );
  AOI22_X1 U16604 ( .A1(n13781), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n14769), .ZN(n19076) );
  INV_X1 U16605 ( .A(n19076), .ZN(n13319) );
  NAND2_X1 U16606 ( .A1(n19139), .A2(n13319), .ZN(n13354) );
  NAND2_X1 U16607 ( .A1(n13320), .A2(n13354), .ZN(P2_U2970) );
  OAI21_X1 U16608 ( .B1(n16125), .B2(n10565), .A(n13321), .ZN(n13324) );
  NOR2_X1 U16609 ( .A1(n13322), .A2(n16055), .ZN(n13323) );
  AOI211_X1 U16610 ( .C1(n14651), .C2(n16114), .A(n13324), .B(n13323), .ZN(
        n13326) );
  NAND2_X1 U16611 ( .A1(n9829), .A2(n16117), .ZN(n13325) );
  OAI211_X1 U16612 ( .C1(n13327), .C2(n15067), .A(n13326), .B(n13325), .ZN(
        P2_U3012) );
  INV_X1 U16613 ( .A(n13331), .ZN(n13328) );
  AOI222_X1 U16614 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n13331), .B1(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n13330), .C1(n13329), .C2(
        n13328), .ZN(n13378) );
  OAI21_X1 U16615 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n13333), .A(
        n13332), .ZN(n13383) );
  AND2_X1 U16616 ( .A1(n18976), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n13385) );
  INV_X1 U16617 ( .A(n13385), .ZN(n13334) );
  OAI21_X1 U16618 ( .B1(n16055), .B2(n13383), .A(n13334), .ZN(n13336) );
  OAI22_X1 U16619 ( .A1(n16068), .A2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B1(
        n14672), .B2(n16088), .ZN(n13335) );
  AOI211_X1 U16620 ( .C1(n16062), .C2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n13336), .B(n13335), .ZN(n13337) );
  OAI21_X1 U16621 ( .B1(n13378), .B2(n15067), .A(n13337), .ZN(P2_U3013) );
  INV_X1 U16622 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n13398) );
  NAND2_X1 U16623 ( .A1(n13338), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n13341) );
  INV_X1 U16624 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n16353) );
  OR2_X1 U16625 ( .A1(n14769), .A2(n16353), .ZN(n13340) );
  NAND2_X1 U16626 ( .A1(n14769), .A2(BUF2_REG_10__SCAN_IN), .ZN(n13339) );
  NAND2_X1 U16627 ( .A1(n13340), .A2(n13339), .ZN(n19051) );
  NAND2_X1 U16628 ( .A1(n19139), .A2(n19051), .ZN(n13342) );
  OAI211_X1 U16629 ( .C1(n13398), .C2(n13344), .A(n13341), .B(n13342), .ZN(
        P2_U2962) );
  INV_X1 U16630 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n19110) );
  NAND2_X1 U16631 ( .A1(n13338), .A2(P2_LWORD_REG_10__SCAN_IN), .ZN(n13343) );
  OAI211_X1 U16632 ( .C1(n19110), .C2(n13344), .A(n13343), .B(n13342), .ZN(
        P2_U2977) );
  NAND2_X1 U16633 ( .A1(n9779), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n13345) );
  AND4_X1 U16634 ( .A1(n12311), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n13345), 
        .A4(n19796), .ZN(n13346) );
  INV_X1 U16635 ( .A(n16217), .ZN(n13347) );
  NAND2_X1 U16636 ( .A1(n13347), .A2(n16213), .ZN(n15380) );
  NAND2_X1 U16637 ( .A1(n15369), .A2(n13348), .ZN(n15398) );
  NAND2_X1 U16638 ( .A1(n15380), .A2(n15398), .ZN(n13349) );
  NAND2_X1 U16639 ( .A1(n19020), .A2(n10480), .ZN(n19031) );
  MUX2_X1 U16640 ( .A(n13350), .B(n15359), .S(n19020), .Z(n13351) );
  OAI21_X1 U16641 ( .B1(n19817), .B2(n19031), .A(n13351), .ZN(P2_U2887) );
  AOI22_X1 U16642 ( .A1(n13338), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19136), 
        .B2(P2_EAX_REG_6__SCAN_IN), .ZN(n13353) );
  NAND2_X1 U16643 ( .A1(n13353), .A2(n13352), .ZN(P2_U2973) );
  AOI22_X1 U16644 ( .A1(n13338), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19136), 
        .B2(P2_EAX_REG_19__SCAN_IN), .ZN(n13355) );
  NAND2_X1 U16645 ( .A1(n13355), .A2(n13354), .ZN(P2_U2955) );
  AOI22_X1 U16646 ( .A1(n13338), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19136), 
        .B2(P2_EAX_REG_7__SCAN_IN), .ZN(n13357) );
  NAND2_X1 U16647 ( .A1(n13357), .A2(n13356), .ZN(P2_U2974) );
  AOI22_X1 U16648 ( .A1(n13338), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(
        P2_EAX_REG_9__SCAN_IN), .B2(n19143), .ZN(n13359) );
  NAND2_X1 U16649 ( .A1(n13359), .A2(n13358), .ZN(P2_U2976) );
  AOI22_X1 U16650 ( .A1(n13338), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(
        P2_EAX_REG_18__SCAN_IN), .B2(n19143), .ZN(n13361) );
  NAND2_X1 U16651 ( .A1(n13361), .A2(n13360), .ZN(P2_U2954) );
  AOI22_X1 U16652 ( .A1(n13338), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(
        P2_EAX_REG_16__SCAN_IN), .B2(n19143), .ZN(n13363) );
  NAND2_X1 U16653 ( .A1(n13363), .A2(n13362), .ZN(P2_U2952) );
  AOI22_X1 U16654 ( .A1(n13338), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(
        P2_EAX_REG_8__SCAN_IN), .B2(n19136), .ZN(n13365) );
  NAND2_X1 U16655 ( .A1(n13365), .A2(n13364), .ZN(P2_U2975) );
  AOI22_X1 U16656 ( .A1(n13338), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n19136), 
        .B2(P2_EAX_REG_11__SCAN_IN), .ZN(n13367) );
  NAND2_X1 U16657 ( .A1(n13367), .A2(n13366), .ZN(P2_U2978) );
  AOI22_X1 U16658 ( .A1(n13338), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19136), 
        .B2(P2_EAX_REG_17__SCAN_IN), .ZN(n13369) );
  NAND2_X1 U16659 ( .A1(n13369), .A2(n13368), .ZN(P2_U2953) );
  AOI22_X1 U16660 ( .A1(n13338), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19136), 
        .B2(P2_EAX_REG_5__SCAN_IN), .ZN(n13371) );
  NAND2_X1 U16661 ( .A1(n13371), .A2(n13370), .ZN(P2_U2972) );
  INV_X1 U16662 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n14783) );
  INV_X1 U16663 ( .A(n16220), .ZN(n19847) );
  NOR2_X1 U16664 ( .A1(n15544), .A2(n19847), .ZN(n13372) );
  NAND2_X1 U16665 ( .A1(n15377), .A2(n19840), .ZN(n13375) );
  NAND2_X1 U16666 ( .A1(n19136), .A2(n16220), .ZN(n13374) );
  NAND2_X1 U16667 ( .A1(n19121), .A2(n19845), .ZN(n19094) );
  NAND2_X1 U16668 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_STATE2_REG_2__SCAN_IN), .ZN(n19815) );
  OR2_X1 U16669 ( .A1(n19815), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n19123) );
  INV_X2 U16670 ( .A(n19123), .ZN(n19131) );
  INV_X2 U16671 ( .A(n19099), .ZN(n19128) );
  AOI22_X1 U16672 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(n19128), .B1(n19131), 
        .B2(P2_UWORD_REG_11__SCAN_IN), .ZN(n13376) );
  OAI21_X1 U16673 ( .B1(n14783), .B2(n19094), .A(n13376), .ZN(P2_U2924) );
  INV_X1 U16674 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n14819) );
  AOI22_X1 U16675 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(n19128), .B1(n19131), 
        .B2(P2_UWORD_REG_7__SCAN_IN), .ZN(n13377) );
  OAI21_X1 U16676 ( .B1(n14819), .B2(n19094), .A(n13377), .ZN(P2_U2928) );
  MUX2_X1 U16677 ( .A(n15389), .B(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .S(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .Z(n13388) );
  INV_X1 U16678 ( .A(n13378), .ZN(n13380) );
  OAI22_X1 U16679 ( .A1(n15356), .A2(n15389), .B1(n14672), .B2(n15360), .ZN(
        n13379) );
  AOI21_X1 U16680 ( .B1(n13380), .B2(n11126), .A(n13379), .ZN(n13387) );
  XNOR2_X1 U16681 ( .A(n13382), .B(n13381), .ZN(n19811) );
  NOR2_X1 U16682 ( .A1(n16157), .A2(n13383), .ZN(n13384) );
  AOI211_X1 U16683 ( .C1(n19811), .C2(n16181), .A(n13385), .B(n13384), .ZN(
        n13386) );
  OAI211_X1 U16684 ( .C1(n15357), .C2(n13388), .A(n13387), .B(n13386), .ZN(
        P2_U3045) );
  INV_X1 U16685 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n13390) );
  AOI22_X1 U16686 ( .A1(n19131), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n19128), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n13389) );
  OAI21_X1 U16687 ( .B1(n13390), .B2(n19094), .A(n13389), .ZN(P2_U2931) );
  INV_X1 U16688 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n14824) );
  AOI22_X1 U16689 ( .A1(n19131), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19128), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n13391) );
  OAI21_X1 U16690 ( .B1(n14824), .B2(n19094), .A(n13391), .ZN(P2_U2930) );
  INV_X1 U16691 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n14834) );
  AOI22_X1 U16692 ( .A1(n19131), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19128), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n13392) );
  OAI21_X1 U16693 ( .B1(n14834), .B2(n19094), .A(n13392), .ZN(P2_U2932) );
  INV_X1 U16694 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n13394) );
  AOI22_X1 U16695 ( .A1(n19131), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n19128), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n13393) );
  OAI21_X1 U16696 ( .B1(n13394), .B2(n19094), .A(n13393), .ZN(P2_U2933) );
  INV_X1 U16697 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n13915) );
  AOI22_X1 U16698 ( .A1(n19131), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n19128), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n13395) );
  OAI21_X1 U16699 ( .B1(n13915), .B2(n19094), .A(n13395), .ZN(P2_U2935) );
  AOI22_X1 U16700 ( .A1(n19131), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19128), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n13396) );
  OAI21_X1 U16701 ( .B1(n14840), .B2(n19094), .A(n13396), .ZN(P2_U2934) );
  AOI22_X1 U16702 ( .A1(n19131), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n19128), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n13397) );
  OAI21_X1 U16703 ( .B1(n13398), .B2(n19094), .A(n13397), .ZN(P2_U2925) );
  INV_X1 U16704 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n13400) );
  AOI22_X1 U16705 ( .A1(P2_UWORD_REG_6__SCAN_IN), .A2(n19131), .B1(n19128), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n13399) );
  OAI21_X1 U16706 ( .B1(n13400), .B2(n19094), .A(n13399), .ZN(P2_U2929) );
  AOI22_X1 U16707 ( .A1(n19131), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n19128), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n13401) );
  OAI21_X1 U16708 ( .B1(n14763), .B2(n19094), .A(n13401), .ZN(P2_U2922) );
  INV_X1 U16709 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n14800) );
  AOI22_X1 U16710 ( .A1(n19131), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n19128), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n13402) );
  OAI21_X1 U16711 ( .B1(n14800), .B2(n19094), .A(n13402), .ZN(P2_U2926) );
  INV_X1 U16712 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n14810) );
  AOI22_X1 U16713 ( .A1(n19131), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n19128), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n13403) );
  OAI21_X1 U16714 ( .B1(n14810), .B2(n19094), .A(n13403), .ZN(P2_U2927) );
  XNOR2_X1 U16715 ( .A(n13405), .B(n13404), .ZN(n18972) );
  INV_X1 U16716 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n19118) );
  INV_X1 U16717 ( .A(n16033), .ZN(n19174) );
  OAI222_X1 U16718 ( .A1(n18972), .A2(n19061), .B1(n19044), .B2(n19118), .C1(
        n19174), .C2(n19091), .ZN(P2_U2913) );
  NAND2_X1 U16719 ( .A1(n13408), .A2(n13407), .ZN(n13409) );
  AND2_X1 U16720 ( .A1(n13410), .A2(n13409), .ZN(n13817) );
  INV_X1 U16721 ( .A(n13817), .ZN(n13706) );
  NAND2_X1 U16722 ( .A1(n13411), .A2(n14425), .ZN(n13416) );
  NAND2_X1 U16723 ( .A1(n11744), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n13563) );
  INV_X1 U16724 ( .A(n13563), .ZN(n13415) );
  OAI21_X1 U16725 ( .B1(n13413), .B2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n9813), .ZN(n13564) );
  NOR2_X1 U16726 ( .A1(n13564), .A2(n19867), .ZN(n13414) );
  AOI211_X1 U16727 ( .C1(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .C2(n13416), .A(
        n13415), .B(n13414), .ZN(n13417) );
  OAI21_X1 U16728 ( .B1(n20094), .B2(n13706), .A(n13417), .ZN(P1_U2999) );
  OAI21_X1 U16729 ( .B1(n13419), .B2(n13418), .A(n13483), .ZN(n18954) );
  OAI222_X1 U16730 ( .A1(n18954), .A2(n19061), .B1(n19181), .B2(n19091), .C1(
        n19116), .C2(n19044), .ZN(P2_U2912) );
  INV_X1 U16731 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n14271) );
  NAND2_X1 U16732 ( .A1(n13950), .A2(n13459), .ZN(n13457) );
  NOR2_X1 U16733 ( .A1(n20113), .A2(n15631), .ZN(n13420) );
  NAND2_X1 U16734 ( .A1(n13421), .A2(n13420), .ZN(n15608) );
  AOI21_X1 U16735 ( .B1(n13457), .B2(n15608), .A(n19861), .ZN(n13422) );
  NAND2_X1 U16736 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n15939) );
  NAND2_X1 U16737 ( .A1(n20098), .A2(n15933), .ZN(n19970) );
  INV_X2 U16738 ( .A(n19970), .ZN(n19994) );
  AOI22_X1 U16739 ( .A1(P1_UWORD_REG_3__SCAN_IN), .A2(n19994), .B1(n19993), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n13424) );
  OAI21_X1 U16740 ( .B1(n14271), .B2(n19967), .A(n13424), .ZN(P1_U2917) );
  INV_X1 U16741 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n13426) );
  AOI22_X1 U16742 ( .A1(P1_UWORD_REG_0__SCAN_IN), .A2(n19994), .B1(n19993), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n13425) );
  OAI21_X1 U16743 ( .B1(n13426), .B2(n19967), .A(n13425), .ZN(P1_U2920) );
  INV_X1 U16744 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n13428) );
  AOI22_X1 U16745 ( .A1(P1_UWORD_REG_1__SCAN_IN), .A2(n19994), .B1(n19993), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n13427) );
  OAI21_X1 U16746 ( .B1(n13428), .B2(n19967), .A(n13427), .ZN(P1_U2919) );
  INV_X1 U16747 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n13430) );
  AOI22_X1 U16748 ( .A1(P1_UWORD_REG_10__SCAN_IN), .A2(n19994), .B1(n19993), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n13429) );
  OAI21_X1 U16749 ( .B1(n13430), .B2(n19967), .A(n13429), .ZN(P1_U2910) );
  INV_X1 U16750 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n13432) );
  AOI22_X1 U16751 ( .A1(P1_UWORD_REG_4__SCAN_IN), .A2(n19994), .B1(n19993), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n13431) );
  OAI21_X1 U16752 ( .B1(n13432), .B2(n19967), .A(n13431), .ZN(P1_U2916) );
  INV_X1 U16753 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n13434) );
  AOI22_X1 U16754 ( .A1(P1_UWORD_REG_5__SCAN_IN), .A2(n19994), .B1(n19993), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n13433) );
  OAI21_X1 U16755 ( .B1(n13434), .B2(n19967), .A(n13433), .ZN(P1_U2915) );
  INV_X1 U16756 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n13436) );
  AOI22_X1 U16757 ( .A1(P1_UWORD_REG_9__SCAN_IN), .A2(n19994), .B1(n19993), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n13435) );
  OAI21_X1 U16758 ( .B1(n13436), .B2(n19967), .A(n13435), .ZN(P1_U2911) );
  NAND2_X1 U16759 ( .A1(n13698), .A2(n13440), .ZN(n13441) );
  NOR2_X1 U16760 ( .A1(n13695), .A2(n13441), .ZN(n13442) );
  NAND3_X1 U16761 ( .A1(n13443), .A2(n13439), .A3(n13442), .ZN(n14551) );
  INV_X1 U16762 ( .A(n14551), .ZN(n13948) );
  INV_X1 U16763 ( .A(n13465), .ZN(n13444) );
  OR2_X1 U16764 ( .A1(n13445), .A2(n13444), .ZN(n13549) );
  XNOR2_X1 U16765 ( .A(n13446), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13449) );
  XNOR2_X1 U16766 ( .A(n13447), .B(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13448) );
  AOI22_X1 U16767 ( .A1(n13549), .A2(n13449), .B1(n13950), .B2(n13448), .ZN(
        n13451) );
  INV_X1 U16768 ( .A(n13449), .ZN(n13453) );
  NAND3_X1 U16769 ( .A1(n13948), .A2(n13545), .A3(n13453), .ZN(n13450) );
  OAI211_X1 U16770 ( .C1(n13438), .C2(n13948), .A(n13451), .B(n13450), .ZN(
        n13589) );
  NOR2_X1 U16771 ( .A1(n15937), .A2(n20076), .ZN(n14554) );
  OAI22_X1 U16772 ( .A1(n13452), .A2(n20075), .B1(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14555) );
  INV_X1 U16773 ( .A(n14555), .ZN(n13454) );
  AOI222_X1 U16774 ( .A1(n13589), .A2(n14552), .B1(n14554), .B2(n13454), .C1(
        n13453), .C2(n13606), .ZN(n13470) );
  NOR2_X1 U16775 ( .A1(n9796), .A2(n11267), .ZN(n13455) );
  NOR2_X1 U16776 ( .A1(n13456), .A2(n13455), .ZN(n13461) );
  NAND2_X1 U16777 ( .A1(n13457), .A2(n13698), .ZN(n13458) );
  OAI211_X1 U16778 ( .C1(n13696), .C2(n13459), .A(n13458), .B(n15609), .ZN(
        n13460) );
  NAND3_X1 U16779 ( .A1(n13462), .A2(n13461), .A3(n13460), .ZN(n13467) );
  INV_X1 U16780 ( .A(n13463), .ZN(n13464) );
  OAI22_X1 U16781 ( .A1(n13466), .A2(n13465), .B1(n13439), .B2(n13464), .ZN(
        n13702) );
  OR2_X1 U16782 ( .A1(n13467), .A2(n13702), .ZN(n13596) );
  INV_X1 U16783 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n19868) );
  NAND2_X1 U16784 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n15933), .ZN(n13604) );
  OR2_X1 U16785 ( .A1(n19868), .A2(n13604), .ZN(n13468) );
  OAI21_X1 U16786 ( .B1(n15591), .B2(n19861), .A(n13468), .ZN(n13473) );
  AOI21_X1 U16787 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n20098), .A(n13473), 
        .ZN(n13952) );
  NAND2_X1 U16788 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n13952), .ZN(
        n13469) );
  OAI21_X1 U16789 ( .B1(n13470), .B2(n13952), .A(n13469), .ZN(P1_U3472) );
  INV_X1 U16790 ( .A(n13952), .ZN(n14558) );
  INV_X1 U16791 ( .A(n13439), .ZN(n13472) );
  INV_X1 U16792 ( .A(n20254), .ZN(n20482) );
  OR2_X1 U16793 ( .A1(n11391), .A2(n20482), .ZN(n13471) );
  XNOR2_X1 U16794 ( .A(n13471), .B(n13475), .ZN(n13597) );
  INV_X1 U16795 ( .A(n13597), .ZN(n19938) );
  NAND4_X1 U16796 ( .A1(n13473), .A2(n13472), .A3(n14552), .A4(n19938), .ZN(
        n13474) );
  OAI21_X1 U16797 ( .B1(n13475), .B2(n14558), .A(n13474), .ZN(P1_U3468) );
  NAND2_X1 U16798 ( .A1(n13478), .A2(n13477), .ZN(n14615) );
  NOR2_X1 U16799 ( .A1(n19020), .A2(n11017), .ZN(n13481) );
  AOI21_X1 U16800 ( .B1(n13480), .B2(n19020), .A(n13481), .ZN(n13482) );
  OAI21_X1 U16801 ( .B1(n19788), .B2(n19031), .A(n13482), .ZN(P2_U2884) );
  AOI21_X1 U16802 ( .B1(n13484), .B2(n13483), .A(n13535), .ZN(n16180) );
  INV_X1 U16803 ( .A(n16180), .ZN(n13485) );
  INV_X1 U16804 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n19114) );
  OAI222_X1 U16805 ( .A1(n13485), .A2(n19061), .B1(n14811), .B2(n19091), .C1(
        n19114), .C2(n19044), .ZN(P2_U2911) );
  XOR2_X1 U16806 ( .A(n13486), .B(P2_INSTQUEUE_REG_0__5__SCAN_IN), .Z(n13493)
         );
  NAND2_X1 U16807 ( .A1(n13487), .A2(n13852), .ZN(n13490) );
  INV_X1 U16808 ( .A(n13488), .ZN(n13489) );
  NAND2_X1 U16809 ( .A1(n13490), .A2(n13489), .ZN(n18980) );
  NOR2_X1 U16810 ( .A1(n19037), .A2(n18980), .ZN(n13491) );
  AOI21_X1 U16811 ( .B1(P2_EBX_REG_5__SCAN_IN), .B2(n19037), .A(n13491), .ZN(
        n13492) );
  OAI21_X1 U16812 ( .B1(n13493), .B2(n19031), .A(n13492), .ZN(P2_U2882) );
  XNOR2_X1 U16813 ( .A(n19147), .B(n19797), .ZN(n13508) );
  INV_X1 U16814 ( .A(n19811), .ZN(n13502) );
  NAND2_X1 U16815 ( .A1(n19146), .A2(n13502), .ZN(n13505) );
  OAI21_X1 U16816 ( .B1(n19146), .B2(n13502), .A(n13505), .ZN(n19078) );
  XNOR2_X1 U16817 ( .A(n13504), .B(n13503), .ZN(n15363) );
  NOR2_X1 U16818 ( .A1(n19817), .A2(n15363), .ZN(n19085) );
  NOR2_X1 U16819 ( .A1(n19078), .A2(n19085), .ZN(n19077) );
  INV_X1 U16820 ( .A(n13505), .ZN(n13506) );
  NOR2_X1 U16821 ( .A1(n19077), .A2(n13506), .ZN(n13507) );
  NOR2_X1 U16822 ( .A1(n13507), .A2(n13508), .ZN(n19056) );
  AOI21_X1 U16823 ( .B1(n13508), .B2(n13507), .A(n19056), .ZN(n13512) );
  INV_X1 U16824 ( .A(n19091), .ZN(n19055) );
  AOI22_X1 U16825 ( .A1(n19055), .A2(n16046), .B1(P2_EAX_REG_2__SCAN_IN), .B2(
        n19083), .ZN(n13511) );
  INV_X1 U16826 ( .A(n19797), .ZN(n13509) );
  NAND2_X1 U16827 ( .A1(n13509), .A2(n19084), .ZN(n13510) );
  OAI211_X1 U16828 ( .C1(n13512), .C2(n19079), .A(n13511), .B(n13510), .ZN(
        P2_U2917) );
  MUX2_X1 U16829 ( .A(n14672), .B(n11012), .S(n19037), .Z(n13513) );
  OAI21_X1 U16830 ( .B1(n19146), .B2(n19031), .A(n13513), .ZN(P2_U2886) );
  INV_X1 U16831 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n14653) );
  MUX2_X1 U16832 ( .A(n10599), .B(n14653), .S(n19037), .Z(n13514) );
  OAI21_X1 U16833 ( .B1(n19147), .B2(n19031), .A(n13514), .ZN(P2_U2885) );
  INV_X1 U16834 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n13516) );
  AOI22_X1 U16835 ( .A1(P1_UWORD_REG_14__SCAN_IN), .A2(n19994), .B1(n19993), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n13515) );
  OAI21_X1 U16836 ( .B1(n13516), .B2(n19967), .A(n13515), .ZN(P1_U2906) );
  INV_X1 U16837 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n13518) );
  AOI22_X1 U16838 ( .A1(P1_UWORD_REG_6__SCAN_IN), .A2(n19994), .B1(n19993), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n13517) );
  OAI21_X1 U16839 ( .B1(n13518), .B2(n19967), .A(n13517), .ZN(P1_U2914) );
  INV_X1 U16840 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n13520) );
  AOI22_X1 U16841 ( .A1(P1_UWORD_REG_8__SCAN_IN), .A2(n19994), .B1(n19993), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n13519) );
  OAI21_X1 U16842 ( .B1(n13520), .B2(n19967), .A(n13519), .ZN(P1_U2912) );
  INV_X1 U16843 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n13522) );
  AOI22_X1 U16844 ( .A1(P1_UWORD_REG_12__SCAN_IN), .A2(n19994), .B1(n19993), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n13521) );
  OAI21_X1 U16845 ( .B1(n13522), .B2(n19967), .A(n13521), .ZN(P1_U2908) );
  INV_X1 U16846 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n13524) );
  AOI22_X1 U16847 ( .A1(P1_UWORD_REG_13__SCAN_IN), .A2(n19994), .B1(n19993), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n13523) );
  OAI21_X1 U16848 ( .B1(n13524), .B2(n19967), .A(n13523), .ZN(P1_U2907) );
  AOI22_X1 U16849 ( .A1(P1_UWORD_REG_2__SCAN_IN), .A2(n19994), .B1(n19993), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n13525) );
  OAI21_X1 U16850 ( .B1(n14276), .B2(n19967), .A(n13525), .ZN(P1_U2918) );
  INV_X1 U16851 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n20976) );
  AOI22_X1 U16852 ( .A1(P1_UWORD_REG_7__SCAN_IN), .A2(n19994), .B1(n19993), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n13526) );
  OAI21_X1 U16853 ( .B1(n20976), .B2(n19967), .A(n13526), .ZN(P1_U2913) );
  AND2_X1 U16854 ( .A1(n11280), .A2(n15630), .ZN(n13527) );
  OR2_X1 U16855 ( .A1(n20025), .A2(n20113), .ZN(n13650) );
  INV_X1 U16856 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n13534) );
  INV_X1 U16857 ( .A(n20015), .ZN(n13533) );
  INV_X1 U16858 ( .A(n20092), .ZN(n20093) );
  INV_X1 U16859 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n13530) );
  NOR2_X1 U16860 ( .A1(n20093), .A2(n13530), .ZN(n13531) );
  AOI21_X1 U16861 ( .B1(DATAI_15_), .B2(n20093), .A(n13531), .ZN(n14289) );
  INV_X1 U16862 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n13532) );
  OAI222_X1 U16863 ( .A1(n13650), .A2(n13534), .B1(n13533), .B2(n14289), .C1(
        n13532), .C2(n13688), .ZN(P1_U2967) );
  OAI21_X1 U16864 ( .B1(n13536), .B2(n13535), .A(n15310), .ZN(n18941) );
  INV_X1 U16865 ( .A(n14802), .ZN(n13537) );
  INV_X1 U16866 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n19112) );
  OAI222_X1 U16867 ( .A1(n18941), .A2(n19061), .B1(n13537), .B2(n19091), .C1(
        n19112), .C2(n19044), .ZN(P2_U2910) );
  NAND2_X1 U16868 ( .A1(n20760), .A2(n14551), .ZN(n13555) );
  NAND2_X1 U16869 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13539) );
  INV_X1 U16870 ( .A(n13539), .ZN(n13538) );
  MUX2_X1 U16871 ( .A(n13539), .B(n13538), .S(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n13552) );
  INV_X1 U16872 ( .A(n13950), .ZN(n15585) );
  INV_X1 U16873 ( .A(n13540), .ZN(n13544) );
  NOR2_X1 U16874 ( .A1(n13446), .A2(n13558), .ZN(n13542) );
  NOR2_X1 U16875 ( .A1(n13542), .A2(n13541), .ZN(n13543) );
  NAND2_X1 U16876 ( .A1(n13544), .A2(n13543), .ZN(n13556) );
  NAND3_X1 U16877 ( .A1(n13948), .A2(n13545), .A3(n13556), .ZN(n13551) );
  MUX2_X1 U16878 ( .A(n11140), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n13446), .Z(n13547) );
  NOR2_X1 U16879 ( .A1(n13547), .A2(n13546), .ZN(n13548) );
  NAND2_X1 U16880 ( .A1(n13549), .A2(n13548), .ZN(n13550) );
  OAI211_X1 U16881 ( .C1(n13552), .C2(n15585), .A(n13551), .B(n13550), .ZN(
        n13553) );
  INV_X1 U16882 ( .A(n13553), .ZN(n13554) );
  NAND2_X1 U16883 ( .A1(n13555), .A2(n13554), .ZN(n13588) );
  AOI22_X1 U16884 ( .A1(n13588), .A2(n14552), .B1(n13606), .B2(n13556), .ZN(
        n13557) );
  MUX2_X1 U16885 ( .A(n13558), .B(n13557), .S(n14558), .Z(n13559) );
  INV_X1 U16886 ( .A(n13559), .ZN(P1_U3469) );
  OR2_X1 U16887 ( .A1(n13560), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13562) );
  AND2_X1 U16888 ( .A1(n13562), .A2(n13561), .ZN(n13818) );
  OAI21_X1 U16889 ( .B1(n15923), .B2(n13564), .A(n13563), .ZN(n13568) );
  AOI21_X1 U16890 ( .B1(n20053), .B2(n20076), .A(n20072), .ZN(n14532) );
  NOR3_X1 U16891 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n20053), .A3(
        n13565), .ZN(n13566) );
  AOI21_X1 U16892 ( .B1(n14532), .B2(n14504), .A(n13566), .ZN(n13567) );
  AOI211_X1 U16893 ( .C1(n20063), .C2(n13818), .A(n13568), .B(n13567), .ZN(
        n13569) );
  INV_X1 U16894 ( .A(n13569), .ZN(P1_U3031) );
  OAI21_X1 U16895 ( .B1(n13570), .B2(n13488), .A(n13583), .ZN(n16116) );
  NOR2_X1 U16896 ( .A1(n13486), .A2(n13571), .ZN(n13573) );
  OAI211_X1 U16897 ( .C1(n13573), .C2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A(
        n19038), .B(n13572), .ZN(n13575) );
  NAND2_X1 U16898 ( .A1(n19037), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n13574) );
  OAI211_X1 U16899 ( .C1(n16116), .C2(n19037), .A(n13575), .B(n13574), .ZN(
        P2_U2881) );
  OAI21_X1 U16900 ( .B1(n13577), .B2(n13576), .A(n13623), .ZN(n20050) );
  XNOR2_X1 U16901 ( .A(n13749), .B(n13696), .ZN(n14533) );
  INV_X1 U16902 ( .A(n14533), .ZN(n13579) );
  OAI22_X1 U16903 ( .A1(n15737), .A2(n13579), .B1(n13578), .B2(n19966), .ZN(
        n13580) );
  INV_X1 U16904 ( .A(n13580), .ZN(n13581) );
  OAI21_X1 U16905 ( .B1(n20050), .B2(n14213), .A(n13581), .ZN(P1_U2871) );
  INV_X1 U16906 ( .A(n13818), .ZN(n13582) );
  OAI222_X1 U16907 ( .A1(n13706), .A2(n14213), .B1(n11618), .B2(n19966), .C1(
        n13582), .C2(n15737), .ZN(P1_U2872) );
  XOR2_X1 U16908 ( .A(n13572), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .Z(n13587)
         );
  AOI21_X1 U16909 ( .B1(n13584), .B2(n13583), .A(n14603), .ZN(n13585) );
  INV_X1 U16910 ( .A(n13585), .ZN(n18953) );
  MUX2_X1 U16911 ( .A(n11061), .B(n18953), .S(n19020), .Z(n13586) );
  OAI21_X1 U16912 ( .B1(n13587), .B2(n19031), .A(n13586), .ZN(P2_U2880) );
  MUX2_X1 U16913 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n13588), .S(
        n13596), .Z(n15595) );
  NAND2_X1 U16914 ( .A1(n15595), .A2(n15937), .ZN(n13593) );
  NOR2_X1 U16915 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n15937), .ZN(n13599) );
  NAND2_X1 U16916 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n13599), .ZN(
        n13592) );
  MUX2_X1 U16917 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n13589), .S(
        n13596), .Z(n15592) );
  AOI22_X1 U16918 ( .A1(n13599), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n15592), .B2(n15937), .ZN(n13591) );
  AOI21_X1 U16919 ( .B1(n13593), .B2(n13592), .A(n13591), .ZN(n15606) );
  INV_X1 U16920 ( .A(n13594), .ZN(n13595) );
  NAND2_X1 U16921 ( .A1(n15606), .A2(n13595), .ZN(n13613) );
  OAI21_X1 U16922 ( .B1(n13439), .B2(n13597), .A(n13596), .ZN(n13598) );
  NAND2_X1 U16923 ( .A1(n13598), .A2(n15937), .ZN(n13601) );
  NAND2_X1 U16924 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n13599), .ZN(
        n13600) );
  NAND2_X1 U16925 ( .A1(n13601), .A2(n13600), .ZN(n13603) );
  NAND2_X1 U16926 ( .A1(n15591), .A2(n13475), .ZN(n13602) );
  NAND2_X1 U16927 ( .A1(n13603), .A2(n13602), .ZN(n15602) );
  AND2_X1 U16928 ( .A1(n15602), .A2(n19868), .ZN(n13605) );
  AOI21_X1 U16929 ( .B1(n13613), .B2(n13605), .A(n13604), .ZN(n13608) );
  NAND2_X1 U16930 ( .A1(n20623), .A2(n15937), .ZN(n15935) );
  INV_X1 U16931 ( .A(n15935), .ZN(n20791) );
  INV_X1 U16932 ( .A(n20259), .ZN(n13607) );
  NAND2_X1 U16933 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20493), .ZN(n20761) );
  INV_X1 U16934 ( .A(n20761), .ZN(n14545) );
  NOR2_X1 U16935 ( .A1(n13609), .A2(n14545), .ZN(n13611) );
  INV_X1 U16936 ( .A(n20544), .ZN(n20758) );
  NOR2_X1 U16937 ( .A1(P1_STATEBS16_REG_SCAN_IN), .A2(n20632), .ZN(n20762) );
  MUX2_X1 U16938 ( .A(n20758), .B(n20762), .S(n20543), .Z(n13610) );
  OAI21_X1 U16939 ( .B1(n13611), .B2(n13610), .A(n20771), .ZN(n13612) );
  OAI21_X1 U16940 ( .B1(n20771), .B2(n20622), .A(n13612), .ZN(P1_U3477) );
  AND3_X1 U16941 ( .A1(n13613), .A2(n15933), .A3(n15602), .ZN(n15617) );
  INV_X1 U16942 ( .A(n12672), .ZN(n20217) );
  OAI22_X1 U16943 ( .A1(n20179), .A2(n20632), .B1(n20217), .B2(n14545), .ZN(
        n13614) );
  OAI21_X1 U16944 ( .B1(n15617), .B2(n13614), .A(n20771), .ZN(n13615) );
  OAI21_X1 U16945 ( .B1(n20771), .B2(n20538), .A(n13615), .ZN(P1_U3478) );
  INV_X1 U16946 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n19108) );
  INV_X1 U16947 ( .A(n14785), .ZN(n13619) );
  OAI21_X1 U16948 ( .B1(n13618), .B2(n13617), .A(n13616), .ZN(n18914) );
  OAI222_X1 U16949 ( .A1(n19044), .A2(n19108), .B1(n13619), .B2(n19091), .C1(
        n18914), .C2(n19061), .ZN(P2_U2908) );
  INV_X1 U16950 ( .A(n13621), .ZN(n13622) );
  AOI21_X1 U16951 ( .B1(n13620), .B2(n13623), .A(n13622), .ZN(n13707) );
  NAND2_X1 U16952 ( .A1(n13625), .A2(n13624), .ZN(n13626) );
  NAND2_X1 U16953 ( .A1(n13736), .A2(n13626), .ZN(n20082) );
  OAI22_X1 U16954 ( .A1(n15737), .A2(n20082), .B1(n13627), .B2(n19966), .ZN(
        n13628) );
  AOI21_X1 U16955 ( .B1(n13707), .B2(n13156), .A(n13628), .ZN(n13629) );
  INV_X1 U16956 ( .A(n13629), .ZN(P1_U2870) );
  AOI22_X1 U16957 ( .A1(n9778), .A2(P1_EAX_REG_17__SCAN_IN), .B1(
        P1_UWORD_REG_1__SCAN_IN), .B2(n20030), .ZN(n13633) );
  NAND2_X1 U16958 ( .A1(n20093), .A2(DATAI_1_), .ZN(n13631) );
  NAND2_X1 U16959 ( .A1(n20092), .A2(BUF1_REG_1__SCAN_IN), .ZN(n13630) );
  AND2_X1 U16960 ( .A1(n13631), .A2(n13630), .ZN(n20115) );
  INV_X1 U16961 ( .A(n20115), .ZN(n13632) );
  NAND2_X1 U16962 ( .A1(n20015), .A2(n13632), .ZN(n13658) );
  NAND2_X1 U16963 ( .A1(n13633), .A2(n13658), .ZN(P1_U2938) );
  AOI22_X1 U16964 ( .A1(n9778), .A2(P1_EAX_REG_7__SCAN_IN), .B1(
        P1_LWORD_REG_7__SCAN_IN), .B2(n20030), .ZN(n13637) );
  NAND2_X1 U16965 ( .A1(n20093), .A2(DATAI_7_), .ZN(n13635) );
  NAND2_X1 U16966 ( .A1(n20092), .A2(BUF1_REG_7__SCAN_IN), .ZN(n13634) );
  AND2_X1 U16967 ( .A1(n13635), .A2(n13634), .ZN(n20146) );
  INV_X1 U16968 ( .A(n20146), .ZN(n13636) );
  NAND2_X1 U16969 ( .A1(n20015), .A2(n13636), .ZN(n13664) );
  NAND2_X1 U16970 ( .A1(n13637), .A2(n13664), .ZN(P1_U2959) );
  AOI22_X1 U16971 ( .A1(n9778), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_UWORD_REG_0__SCAN_IN), .B2(n20030), .ZN(n13641) );
  NAND2_X1 U16972 ( .A1(n20093), .A2(DATAI_0_), .ZN(n13639) );
  NAND2_X1 U16973 ( .A1(n20092), .A2(BUF1_REG_0__SCAN_IN), .ZN(n13638) );
  AND2_X1 U16974 ( .A1(n13639), .A2(n13638), .ZN(n20106) );
  INV_X1 U16975 ( .A(n20106), .ZN(n13640) );
  NAND2_X1 U16976 ( .A1(n20015), .A2(n13640), .ZN(n13674) );
  NAND2_X1 U16977 ( .A1(n13641), .A2(n13674), .ZN(P1_U2937) );
  AOI22_X1 U16978 ( .A1(n9778), .A2(P1_EAX_REG_19__SCAN_IN), .B1(
        P1_UWORD_REG_3__SCAN_IN), .B2(n20030), .ZN(n13645) );
  NAND2_X1 U16979 ( .A1(n20093), .A2(DATAI_3_), .ZN(n13643) );
  NAND2_X1 U16980 ( .A1(n20092), .A2(BUF1_REG_3__SCAN_IN), .ZN(n13642) );
  AND2_X1 U16981 ( .A1(n13643), .A2(n13642), .ZN(n20124) );
  INV_X1 U16982 ( .A(n20124), .ZN(n13644) );
  NAND2_X1 U16983 ( .A1(n20015), .A2(n13644), .ZN(n13666) );
  NAND2_X1 U16984 ( .A1(n13645), .A2(n13666), .ZN(P1_U2940) );
  AOI22_X1 U16985 ( .A1(n9778), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_UWORD_REG_2__SCAN_IN), .B2(n20030), .ZN(n13649) );
  NAND2_X1 U16986 ( .A1(n20093), .A2(DATAI_2_), .ZN(n13647) );
  NAND2_X1 U16987 ( .A1(n20092), .A2(BUF1_REG_2__SCAN_IN), .ZN(n13646) );
  AND2_X1 U16988 ( .A1(n13647), .A2(n13646), .ZN(n20119) );
  INV_X1 U16989 ( .A(n20119), .ZN(n13648) );
  NAND2_X1 U16990 ( .A1(n20015), .A2(n13648), .ZN(n13676) );
  NAND2_X1 U16991 ( .A1(n13649), .A2(n13676), .ZN(P1_U2939) );
  AOI22_X1 U16992 ( .A1(n9778), .A2(P1_EAX_REG_20__SCAN_IN), .B1(
        P1_UWORD_REG_4__SCAN_IN), .B2(n20030), .ZN(n13654) );
  NAND2_X1 U16993 ( .A1(n20093), .A2(DATAI_4_), .ZN(n13652) );
  NAND2_X1 U16994 ( .A1(n20092), .A2(BUF1_REG_4__SCAN_IN), .ZN(n13651) );
  AND2_X1 U16995 ( .A1(n13652), .A2(n13651), .ZN(n20129) );
  INV_X1 U16996 ( .A(n20129), .ZN(n13653) );
  NAND2_X1 U16997 ( .A1(n20015), .A2(n13653), .ZN(n13662) );
  NAND2_X1 U16998 ( .A1(n13654), .A2(n13662), .ZN(P1_U2941) );
  AOI22_X1 U16999 ( .A1(n9778), .A2(P1_EAX_REG_5__SCAN_IN), .B1(
        P1_LWORD_REG_5__SCAN_IN), .B2(n20025), .ZN(n13657) );
  NAND2_X1 U17000 ( .A1(n20093), .A2(DATAI_5_), .ZN(n13656) );
  NAND2_X1 U17001 ( .A1(n20092), .A2(BUF1_REG_5__SCAN_IN), .ZN(n13655) );
  AND2_X1 U17002 ( .A1(n13656), .A2(n13655), .ZN(n20133) );
  INV_X1 U17003 ( .A(n20133), .ZN(n14262) );
  NAND2_X1 U17004 ( .A1(n20015), .A2(n14262), .ZN(n13660) );
  NAND2_X1 U17005 ( .A1(n13657), .A2(n13660), .ZN(P1_U2957) );
  AOI22_X1 U17006 ( .A1(n9778), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_LWORD_REG_1__SCAN_IN), .B2(n20025), .ZN(n13659) );
  NAND2_X1 U17007 ( .A1(n13659), .A2(n13658), .ZN(P1_U2953) );
  AOI22_X1 U17008 ( .A1(n9778), .A2(P1_EAX_REG_21__SCAN_IN), .B1(
        P1_UWORD_REG_5__SCAN_IN), .B2(n20030), .ZN(n13661) );
  NAND2_X1 U17009 ( .A1(n13661), .A2(n13660), .ZN(P1_U2942) );
  AOI22_X1 U17010 ( .A1(n9778), .A2(P1_EAX_REG_4__SCAN_IN), .B1(
        P1_LWORD_REG_4__SCAN_IN), .B2(n20025), .ZN(n13663) );
  NAND2_X1 U17011 ( .A1(n13663), .A2(n13662), .ZN(P1_U2956) );
  AOI22_X1 U17012 ( .A1(n9778), .A2(P1_EAX_REG_23__SCAN_IN), .B1(
        P1_UWORD_REG_7__SCAN_IN), .B2(n20030), .ZN(n13665) );
  NAND2_X1 U17013 ( .A1(n13665), .A2(n13664), .ZN(P1_U2944) );
  AOI22_X1 U17014 ( .A1(n9778), .A2(P1_EAX_REG_3__SCAN_IN), .B1(
        P1_LWORD_REG_3__SCAN_IN), .B2(n20025), .ZN(n13667) );
  NAND2_X1 U17015 ( .A1(n13667), .A2(n13666), .ZN(P1_U2955) );
  AOI22_X1 U17016 ( .A1(n9778), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_UWORD_REG_6__SCAN_IN), .B2(n20030), .ZN(n13671) );
  NAND2_X1 U17017 ( .A1(n20093), .A2(DATAI_6_), .ZN(n13669) );
  NAND2_X1 U17018 ( .A1(n20092), .A2(BUF1_REG_6__SCAN_IN), .ZN(n13668) );
  AND2_X1 U17019 ( .A1(n13669), .A2(n13668), .ZN(n20138) );
  INV_X1 U17020 ( .A(n20138), .ZN(n13670) );
  NAND2_X1 U17021 ( .A1(n20015), .A2(n13670), .ZN(n13672) );
  NAND2_X1 U17022 ( .A1(n13671), .A2(n13672), .ZN(P1_U2943) );
  AOI22_X1 U17023 ( .A1(n9778), .A2(P1_EAX_REG_6__SCAN_IN), .B1(
        P1_LWORD_REG_6__SCAN_IN), .B2(n20025), .ZN(n13673) );
  NAND2_X1 U17024 ( .A1(n13673), .A2(n13672), .ZN(P1_U2958) );
  AOI22_X1 U17025 ( .A1(n9778), .A2(P1_EAX_REG_0__SCAN_IN), .B1(
        P1_LWORD_REG_0__SCAN_IN), .B2(n20030), .ZN(n13675) );
  NAND2_X1 U17026 ( .A1(n13675), .A2(n13674), .ZN(P1_U2952) );
  AOI22_X1 U17027 ( .A1(n9778), .A2(P1_EAX_REG_2__SCAN_IN), .B1(
        P1_LWORD_REG_2__SCAN_IN), .B2(n20025), .ZN(n13677) );
  NAND2_X1 U17028 ( .A1(n13677), .A2(n13676), .ZN(P1_U2954) );
  INV_X1 U17029 ( .A(n13678), .ZN(n19030) );
  OAI211_X1 U17030 ( .C1(n19030), .C2(n13680), .A(n19038), .B(n13679), .ZN(
        n13684) );
  AOI21_X1 U17031 ( .B1(n13682), .B2(n13681), .A(n15308), .ZN(n15325) );
  NAND2_X1 U17032 ( .A1(n19020), .A2(n15325), .ZN(n13683) );
  OAI211_X1 U17033 ( .C1(n19020), .C2(n11075), .A(n13684), .B(n13683), .ZN(
        P2_U2878) );
  INV_X1 U17034 ( .A(P1_UWORD_REG_11__SCAN_IN), .ZN(n20997) );
  INV_X1 U17035 ( .A(DATAI_11_), .ZN(n13686) );
  NAND2_X1 U17036 ( .A1(n20092), .A2(BUF1_REG_11__SCAN_IN), .ZN(n13685) );
  OAI21_X1 U17037 ( .B1(n20092), .B2(n13686), .A(n13685), .ZN(n14299) );
  NAND2_X1 U17038 ( .A1(n20015), .A2(n14299), .ZN(n20023) );
  NAND2_X1 U17039 ( .A1(n9778), .A2(P1_EAX_REG_27__SCAN_IN), .ZN(n13687) );
  OAI211_X1 U17040 ( .C1(n13688), .C2(n20997), .A(n20023), .B(n13687), .ZN(
        P1_U2948) );
  OAI21_X1 U17041 ( .B1(n13691), .B2(n13690), .A(n13689), .ZN(n20074) );
  AOI22_X1 U17042 ( .A1(n20043), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n11744), .B2(P1_REIP_REG_2__SCAN_IN), .ZN(n13692) );
  OAI21_X1 U17043 ( .B1(n20041), .B2(n13828), .A(n13692), .ZN(n13693) );
  AOI21_X1 U17044 ( .B1(n13707), .B2(n20038), .A(n13693), .ZN(n13694) );
  OAI21_X1 U17045 ( .B1(n19867), .B2(n20074), .A(n13694), .ZN(P1_U2997) );
  INV_X1 U17046 ( .A(n13695), .ZN(n13700) );
  NAND2_X1 U17047 ( .A1(n13696), .A2(n15609), .ZN(n13697) );
  OAI22_X1 U17048 ( .A1(n13700), .A2(n13699), .B1(n13698), .B2(n13697), .ZN(
        n13701) );
  NAND2_X1 U17049 ( .A1(n11262), .A2(n9790), .ZN(n13705) );
  INV_X1 U17050 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n19997) );
  OAI222_X1 U17051 ( .A1(n14296), .A2(n13706), .B1(n14294), .B2(n19997), .C1(
        n14297), .C2(n20106), .ZN(P1_U2904) );
  INV_X1 U17052 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n19992) );
  OAI222_X1 U17053 ( .A1(n14296), .A2(n20050), .B1(n14294), .B2(n19992), .C1(
        n14297), .C2(n20115), .ZN(P1_U2903) );
  INV_X1 U17054 ( .A(n13707), .ZN(n13835) );
  INV_X1 U17055 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n19990) );
  OAI222_X1 U17056 ( .A1(n14296), .A2(n13835), .B1(n14294), .B2(n19990), .C1(
        n14297), .C2(n20119), .ZN(P1_U2902) );
  OAI21_X1 U17057 ( .B1(n13708), .B2(n13710), .A(n13709), .ZN(n20064) );
  XOR2_X1 U17058 ( .A(n13711), .B(n13712), .Z(n13723) );
  AOI22_X1 U17059 ( .A1(n20043), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B1(
        n11744), .B2(P1_REIP_REG_3__SCAN_IN), .ZN(n13713) );
  OAI21_X1 U17060 ( .B1(n20041), .B2(n13842), .A(n13713), .ZN(n13714) );
  AOI21_X1 U17061 ( .B1(n13723), .B2(n20038), .A(n13714), .ZN(n13715) );
  OAI21_X1 U17062 ( .B1(n20064), .B2(n19867), .A(n13715), .ZN(P1_U2996) );
  XNOR2_X1 U17063 ( .A(n13716), .B(n19016), .ZN(n13722) );
  NAND2_X1 U17064 ( .A1(n19037), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n13721) );
  AND2_X1 U17065 ( .A1(n15307), .A2(n13718), .ZN(n13719) );
  NOR2_X1 U17066 ( .A1(n13717), .A2(n13719), .ZN(n18907) );
  NAND2_X1 U17067 ( .A1(n18907), .A2(n19020), .ZN(n13720) );
  OAI211_X1 U17068 ( .C1(n13722), .C2(n19031), .A(n13721), .B(n13720), .ZN(
        P2_U2876) );
  INV_X1 U17069 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n19988) );
  OAI222_X1 U17070 ( .A1(n14296), .A2(n13846), .B1(n14294), .B2(n19988), .C1(
        n14297), .C2(n20124), .ZN(P1_U2901) );
  INV_X1 U17071 ( .A(n13724), .ZN(n14578) );
  INV_X1 U17072 ( .A(n13725), .ZN(n13728) );
  INV_X1 U17073 ( .A(n13726), .ZN(n13727) );
  NAND2_X1 U17074 ( .A1(n13728), .A2(n13727), .ZN(n13729) );
  NAND2_X1 U17075 ( .A1(n14578), .A2(n13729), .ZN(n18906) );
  INV_X1 U17076 ( .A(n14765), .ZN(n13730) );
  INV_X1 U17077 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n19104) );
  OAI222_X1 U17078 ( .A1(n18906), .A2(n19061), .B1(n13730), .B2(n19091), .C1(
        n19104), .C2(n19044), .ZN(P2_U2906) );
  INV_X1 U17079 ( .A(n13731), .ZN(n13756) );
  NAND2_X1 U17080 ( .A1(n13732), .A2(n13733), .ZN(n13734) );
  AND2_X1 U17081 ( .A1(n13756), .A2(n13734), .ZN(n20037) );
  INV_X1 U17082 ( .A(n20037), .ZN(n13742) );
  INV_X1 U17083 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n19986) );
  OAI222_X1 U17084 ( .A1(n14296), .A2(n13742), .B1(n19986), .B2(n14294), .C1(
        n14297), .C2(n20129), .ZN(P1_U2900) );
  AND2_X1 U17085 ( .A1(n13736), .A2(n13735), .ZN(n13737) );
  OR2_X1 U17086 ( .A1(n13740), .A2(n13737), .ZN(n13838) );
  INV_X1 U17087 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n13738) );
  OAI222_X1 U17088 ( .A1(n13838), .A2(n15737), .B1(n19966), .B2(n13738), .C1(
        n13846), .C2(n14213), .ZN(P1_U2869) );
  OR2_X1 U17089 ( .A1(n13740), .A2(n13739), .ZN(n13741) );
  NAND2_X1 U17090 ( .A1(n15919), .A2(n13741), .ZN(n20056) );
  INV_X1 U17091 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n13743) );
  OAI222_X1 U17092 ( .A1(n20056), .A2(n15737), .B1(n19966), .B2(n13743), .C1(
        n13742), .C2(n14213), .ZN(P1_U2868) );
  NAND2_X1 U17093 ( .A1(n13747), .A2(n13744), .ZN(n13745) );
  INV_X1 U17094 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n13748) );
  INV_X1 U17095 ( .A(n11720), .ZN(n13746) );
  AND2_X1 U17096 ( .A1(n13747), .A2(n13746), .ZN(n19939) );
  INV_X1 U17097 ( .A(n13609), .ZN(n20577) );
  AOI22_X1 U17098 ( .A1(n19950), .A2(n13748), .B1(n19939), .B2(n20577), .ZN(
        n13753) );
  AOI22_X1 U17099 ( .A1(n19948), .A2(n13749), .B1(n19937), .B2(
        P1_EBX_REG_1__SCAN_IN), .ZN(n13752) );
  INV_X1 U17100 ( .A(n19924), .ZN(n19895) );
  AOI22_X1 U17101 ( .A1(n19891), .A2(n20044), .B1(n19895), .B2(
        P1_REIP_REG_1__SCAN_IN), .ZN(n13751) );
  NAND2_X1 U17102 ( .A1(n19940), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13750) );
  AND4_X1 U17103 ( .A1(n13753), .A2(n13752), .A3(n13751), .A4(n13750), .ZN(
        n13754) );
  OAI21_X1 U17104 ( .B1(n19931), .B2(n20050), .A(n13754), .ZN(P1_U2839) );
  AND2_X1 U17105 ( .A1(n13756), .A2(n13755), .ZN(n13758) );
  OR2_X1 U17106 ( .A1(n13758), .A2(n13757), .ZN(n19932) );
  OAI222_X1 U17107 ( .A1(n19932), .A2(n14296), .B1(n13759), .B2(n14294), .C1(
        n14297), .C2(n20133), .ZN(P1_U2899) );
  INV_X1 U17108 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n13769) );
  OAI211_X1 U17109 ( .C1(n13760), .C2(n13762), .A(n13761), .B(n19038), .ZN(
        n13768) );
  NAND2_X1 U17110 ( .A1(n13764), .A2(n13765), .ZN(n13766) );
  NAND2_X1 U17111 ( .A1(n13763), .A2(n13766), .ZN(n15074) );
  INV_X1 U17112 ( .A(n15074), .ZN(n18903) );
  NAND2_X1 U17113 ( .A1(n18903), .A2(n19020), .ZN(n13767) );
  OAI211_X1 U17114 ( .C1(n19020), .C2(n13769), .A(n13768), .B(n13767), .ZN(
        P2_U2874) );
  NAND2_X1 U17115 ( .A1(n19357), .A2(n19787), .ZN(n13770) );
  NAND2_X1 U17116 ( .A1(n13770), .A2(n19786), .ZN(n13779) );
  INV_X1 U17117 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19794) );
  NAND2_X1 U17118 ( .A1(n19794), .A2(n19804), .ZN(n19215) );
  INV_X1 U17119 ( .A(n19215), .ZN(n16208) );
  NAND2_X1 U17120 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n16208), .ZN(
        n19214) );
  INV_X1 U17121 ( .A(n19214), .ZN(n13771) );
  OR2_X1 U17122 ( .A1(n13779), .A2(n13771), .ZN(n13776) );
  NAND2_X1 U17123 ( .A1(n10733), .A2(n19796), .ZN(n13774) );
  NOR2_X1 U17124 ( .A1(n19353), .A2(n19215), .ZN(n19255) );
  NOR2_X1 U17125 ( .A1(n19255), .A2(n19786), .ZN(n13773) );
  AOI21_X1 U17126 ( .B1(n15386), .B2(n19149), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n19849) );
  NAND2_X1 U17127 ( .A1(n19849), .A2(n19815), .ZN(n13772) );
  AOI21_X1 U17128 ( .B1(n13774), .B2(n13773), .A(n19268), .ZN(n13775) );
  NAND2_X1 U17129 ( .A1(n13776), .A2(n13775), .ZN(n19258) );
  INV_X1 U17130 ( .A(n19258), .ZN(n19243) );
  INV_X1 U17131 ( .A(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13785) );
  OAI21_X1 U17132 ( .B1(n10733), .B2(n19255), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n13778) );
  OAI21_X1 U17133 ( .B1(n13779), .B2(n19214), .A(n13778), .ZN(n19257) );
  AOI22_X1 U17134 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n19178), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n19177), .ZN(n19652) );
  AOI22_X1 U17135 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n19178), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19177), .ZN(n19554) );
  INV_X1 U17136 ( .A(n19554), .ZN(n19649) );
  NAND2_X1 U17137 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19647), .ZN(n19167) );
  AOI22_X1 U17138 ( .A1(n19649), .A2(n19289), .B1(n19255), .B2(n19640), .ZN(
        n13782) );
  OAI21_X1 U17139 ( .B1(n19652), .B2(n19246), .A(n13782), .ZN(n13783) );
  AOI21_X1 U17140 ( .B1(n13777), .B2(n19257), .A(n13783), .ZN(n13784) );
  OAI21_X1 U17141 ( .B1(n19243), .B2(n13785), .A(n13784), .ZN(P2_U3072) );
  XNOR2_X1 U17142 ( .A(n13786), .B(n13787), .ZN(n21141) );
  INV_X1 U17143 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n14640) );
  NAND2_X1 U17144 ( .A1(n16186), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n21132) );
  OAI21_X1 U17145 ( .B1(n16125), .B2(n14640), .A(n21132), .ZN(n13789) );
  NOR2_X1 U17146 ( .A1(n16068), .A2(n14635), .ZN(n13788) );
  AOI211_X1 U17147 ( .C1(n16117), .C2(n13480), .A(n13789), .B(n13788), .ZN(
        n13793) );
  XOR2_X1 U17148 ( .A(n13791), .B(n13790), .Z(n21138) );
  NAND2_X1 U17149 ( .A1(n21138), .A2(n16120), .ZN(n13792) );
  OAI211_X1 U17150 ( .C1(n21141), .C2(n15067), .A(n13793), .B(n13792), .ZN(
        P2_U3011) );
  INV_X1 U17151 ( .A(n19536), .ZN(n19545) );
  NAND2_X1 U17152 ( .A1(n19357), .A2(n19545), .ZN(n13794) );
  NAND2_X1 U17153 ( .A1(n13794), .A2(n19786), .ZN(n13802) );
  NAND2_X1 U17154 ( .A1(n19794), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n19264) );
  INV_X1 U17155 ( .A(n19264), .ZN(n19354) );
  NAND2_X1 U17156 ( .A1(n19354), .A2(n19813), .ZN(n13801) );
  INV_X1 U17157 ( .A(n13801), .ZN(n13795) );
  OR2_X1 U17158 ( .A1(n13802), .A2(n13795), .ZN(n13799) );
  INV_X1 U17159 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n19149) );
  OAI21_X1 U17160 ( .B1(n10731), .B2(n19149), .A(n19796), .ZN(n13797) );
  NOR2_X1 U17161 ( .A1(n19821), .A2(n13801), .ZN(n19308) );
  INV_X1 U17162 ( .A(n19308), .ZN(n13796) );
  AOI21_X1 U17163 ( .B1(n13797), .B2(n13796), .A(n19268), .ZN(n13798) );
  NAND2_X1 U17164 ( .A1(n13799), .A2(n13798), .ZN(n19310) );
  OAI21_X1 U17165 ( .B1(n10731), .B2(n19308), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n13800) );
  OAI21_X1 U17166 ( .B1(n13802), .B2(n13801), .A(n13800), .ZN(n19309) );
  NOR2_X2 U17167 ( .A1(n19352), .A2(n19536), .ZN(n19347) );
  AOI22_X1 U17168 ( .A1(n19649), .A2(n19347), .B1(n19640), .B2(n19308), .ZN(
        n13803) );
  OAI21_X1 U17169 ( .B1(n19652), .B2(n19313), .A(n13803), .ZN(n13804) );
  AOI21_X1 U17170 ( .B1(n13777), .B2(n19309), .A(n13804), .ZN(n13805) );
  OAI21_X1 U17171 ( .B1(n19305), .B2(n13806), .A(n13805), .ZN(P2_U3088) );
  NOR2_X2 U17172 ( .A1(n19076), .A2(n19268), .ZN(n19665) );
  AOI22_X1 U17173 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n19177), .B1(
        BUF1_REG_27__SCAN_IN), .B2(n19178), .ZN(n19669) );
  AOI22_X1 U17174 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n19178), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19177), .ZN(n19571) );
  INV_X1 U17175 ( .A(n19571), .ZN(n19666) );
  AOI22_X1 U17176 ( .A1(n19666), .A2(n19347), .B1(n19308), .B2(n19664), .ZN(
        n13808) );
  OAI21_X1 U17177 ( .B1(n19313), .B2(n19669), .A(n13808), .ZN(n13809) );
  AOI21_X1 U17178 ( .B1(n19665), .B2(n19309), .A(n13809), .ZN(n13810) );
  OAI21_X1 U17179 ( .B1(n19305), .B2(n13811), .A(n13810), .ZN(P2_U3091) );
  INV_X1 U17180 ( .A(n13812), .ZN(n13813) );
  XNOR2_X1 U17181 ( .A(n9876), .B(n13813), .ZN(n15296) );
  INV_X1 U17182 ( .A(n15296), .ZN(n18888) );
  OAI222_X1 U17183 ( .A1(n19044), .A2(n13271), .B1(n18888), .B2(n19061), .C1(
        n19091), .C2(n13814), .ZN(P2_U2904) );
  NAND2_X1 U17184 ( .A1(n19926), .A2(n19924), .ZN(n14074) );
  INV_X1 U17185 ( .A(n14074), .ZN(n13821) );
  INV_X1 U17186 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n20780) );
  INV_X1 U17187 ( .A(n19931), .ZN(n19954) );
  OAI21_X1 U17188 ( .B1(n19940), .B2(n19891), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13815) );
  OAI21_X1 U17189 ( .B1(n19899), .B2(n11618), .A(n13815), .ZN(n13816) );
  AOI21_X1 U17190 ( .B1(n13817), .B2(n19954), .A(n13816), .ZN(n13820) );
  AOI22_X1 U17191 ( .A1(n12672), .A2(n19939), .B1(n19948), .B2(n13818), .ZN(
        n13819) );
  OAI211_X1 U17192 ( .C1(n13821), .C2(n20780), .A(n13820), .B(n13819), .ZN(
        P1_U2840) );
  OR2_X1 U17193 ( .A1(n13757), .A2(n13823), .ZN(n13824) );
  AND2_X1 U17194 ( .A1(n13822), .A2(n13824), .ZN(n19913) );
  INV_X1 U17195 ( .A(n19913), .ZN(n13836) );
  XOR2_X1 U17196 ( .A(n13825), .B(n15921), .Z(n19910) );
  INV_X1 U17197 ( .A(n19966), .ZN(n14203) );
  AOI22_X1 U17198 ( .A1(n19962), .A2(n19910), .B1(P1_EBX_REG_6__SCAN_IN), .B2(
        n14203), .ZN(n13826) );
  OAI21_X1 U17199 ( .B1(n13836), .B2(n14213), .A(n13826), .ZN(P1_U2866) );
  INV_X1 U17200 ( .A(n20082), .ZN(n13833) );
  NAND2_X1 U17201 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_2__SCAN_IN), 
        .ZN(n13837) );
  NAND2_X1 U17202 ( .A1(n19950), .A2(n13837), .ZN(n13830) );
  NAND2_X1 U17203 ( .A1(n19924), .A2(n13830), .ZN(n13839) );
  AOI22_X1 U17204 ( .A1(n19940), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n13839), .B2(P1_REIP_REG_2__SCAN_IN), .ZN(n13827) );
  OAI21_X1 U17205 ( .B1(n19957), .B2(n13828), .A(n13827), .ZN(n13832) );
  INV_X1 U17206 ( .A(n13438), .ZN(n20102) );
  AOI22_X1 U17207 ( .A1(n20102), .A2(n19939), .B1(n19937), .B2(
        P1_EBX_REG_2__SCAN_IN), .ZN(n13829) );
  OAI21_X1 U17208 ( .B1(n13830), .B2(n13748), .A(n13829), .ZN(n13831) );
  AOI211_X1 U17209 ( .C1(n19948), .C2(n13833), .A(n13832), .B(n13831), .ZN(
        n13834) );
  OAI21_X1 U17210 ( .B1(n13835), .B2(n19931), .A(n13834), .ZN(P1_U2838) );
  INV_X1 U17211 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n19983) );
  OAI222_X1 U17212 ( .A1(n14296), .A2(n13836), .B1(n14294), .B2(n19983), .C1(
        n14297), .C2(n20138), .ZN(P1_U2898) );
  NOR3_X1 U17213 ( .A1(n19926), .A2(P1_REIP_REG_3__SCAN_IN), .A3(n13837), .ZN(
        n13844) );
  INV_X1 U17214 ( .A(n13838), .ZN(n20062) );
  AOI22_X1 U17215 ( .A1(n19948), .A2(n20062), .B1(n19937), .B2(
        P1_EBX_REG_3__SCAN_IN), .ZN(n13841) );
  AOI22_X1 U17216 ( .A1(n19940), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B1(
        P1_REIP_REG_3__SCAN_IN), .B2(n13839), .ZN(n13840) );
  OAI211_X1 U17217 ( .C1(n13842), .C2(n19957), .A(n13841), .B(n13840), .ZN(
        n13843) );
  AOI211_X1 U17218 ( .C1(n19939), .C2(n20760), .A(n13844), .B(n13843), .ZN(
        n13845) );
  OAI21_X1 U17219 ( .B1(n13846), .B2(n19931), .A(n13845), .ZN(P1_U2837) );
  XNOR2_X1 U17220 ( .A(n13847), .B(n13848), .ZN(n13869) );
  OAI21_X1 U17221 ( .B1(n13851), .B2(n13850), .A(n9783), .ZN(n13866) );
  OAI21_X1 U17222 ( .B1(n13854), .B2(n13853), .A(n13852), .ZN(n19041) );
  INV_X1 U17223 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n19729) );
  OAI22_X1 U17224 ( .A1(n16125), .A2(n14628), .B1(n19729), .B2(n9889), .ZN(
        n13855) );
  AOI21_X1 U17225 ( .B1(n16114), .B2(n14623), .A(n13855), .ZN(n13856) );
  OAI21_X1 U17226 ( .B1(n19041), .B2(n16088), .A(n13856), .ZN(n13857) );
  AOI21_X1 U17227 ( .B1(n13866), .B2(n16120), .A(n13857), .ZN(n13858) );
  OAI21_X1 U17228 ( .B1(n13869), .B2(n15067), .A(n13858), .ZN(P2_U3010) );
  OAI21_X1 U17229 ( .B1(n15357), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n21126), .ZN(n13890) );
  NAND2_X1 U17230 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n21128), .ZN(
        n15347) );
  INV_X1 U17231 ( .A(n15347), .ZN(n13859) );
  AOI22_X1 U17232 ( .A1(n16186), .A2(P2_REIP_REG_4__SCAN_IN), .B1(n13850), 
        .B2(n13859), .ZN(n13864) );
  AOI21_X1 U17233 ( .B1(n13862), .B2(n13860), .A(n13861), .ZN(n19063) );
  NAND2_X1 U17234 ( .A1(n16181), .A2(n19063), .ZN(n13863) );
  OAI211_X1 U17235 ( .C1(n19041), .C2(n15360), .A(n13864), .B(n13863), .ZN(
        n13865) );
  AOI21_X1 U17236 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n13890), .A(
        n13865), .ZN(n13868) );
  NAND2_X1 U17237 ( .A1(n13866), .A2(n21137), .ZN(n13867) );
  OAI211_X1 U17238 ( .C1(n13869), .C2(n21140), .A(n13868), .B(n13867), .ZN(
        P2_U3042) );
  NAND2_X1 U17239 ( .A1(n13822), .A2(n13871), .ZN(n13872) );
  AND2_X1 U17240 ( .A1(n13870), .A2(n13872), .ZN(n19906) );
  INV_X1 U17241 ( .A(n19906), .ZN(n13873) );
  INV_X1 U17242 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n19981) );
  OAI222_X1 U17243 ( .A1(n14296), .A2(n13873), .B1(n14294), .B2(n19981), .C1(
        n14297), .C2(n20146), .ZN(P1_U2897) );
  AND2_X1 U17244 ( .A1(n13875), .A2(n13874), .ZN(n13876) );
  NOR2_X1 U17245 ( .A1(n13897), .A2(n13876), .ZN(n15907) );
  INV_X1 U17246 ( .A(n15907), .ZN(n19898) );
  INV_X1 U17247 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n19900) );
  OAI22_X1 U17248 ( .A1(n15737), .A2(n19898), .B1(n19900), .B2(n19966), .ZN(
        n13877) );
  AOI21_X1 U17249 ( .B1(n19906), .B2(n13156), .A(n13877), .ZN(n13878) );
  INV_X1 U17250 ( .A(n13878), .ZN(P1_U2865) );
  XNOR2_X1 U17251 ( .A(n13879), .B(n13880), .ZN(n13905) );
  NOR2_X1 U17252 ( .A1(n13882), .A2(n13881), .ZN(n13883) );
  XNOR2_X1 U17253 ( .A(n13884), .B(n13883), .ZN(n13903) );
  OAI21_X1 U17254 ( .B1(n13861), .B2(n13886), .A(n13885), .ZN(n19060) );
  NOR2_X1 U17255 ( .A1(n15360), .A2(n18980), .ZN(n13889) );
  OAI21_X1 U17256 ( .B1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A(n15348), .ZN(n13887) );
  OAI22_X1 U17257 ( .A1(n13887), .A2(n15347), .B1(n9889), .B2(n13900), .ZN(
        n13888) );
  AOI211_X1 U17258 ( .C1(n13890), .C2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(
        n13889), .B(n13888), .ZN(n13891) );
  OAI21_X1 U17259 ( .B1(n19060), .B2(n21133), .A(n13891), .ZN(n13892) );
  AOI21_X1 U17260 ( .B1(n13903), .B2(n21137), .A(n13892), .ZN(n13893) );
  OAI21_X1 U17261 ( .B1(n13905), .B2(n21140), .A(n13893), .ZN(P2_U3041) );
  AOI21_X1 U17262 ( .B1(n13895), .B2(n13870), .A(n13894), .ZN(n13928) );
  INV_X1 U17263 ( .A(n13928), .ZN(n14141) );
  INV_X1 U17264 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n13899) );
  NOR2_X1 U17265 ( .A1(n13897), .A2(n13896), .ZN(n13898) );
  OR2_X1 U17266 ( .A1(n15884), .A2(n13898), .ZN(n15902) );
  OAI222_X1 U17267 ( .A1(n14141), .A2(n14213), .B1(n19966), .B2(n13899), .C1(
        n15902), .C2(n15737), .ZN(P1_U2864) );
  INV_X1 U17268 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n18988) );
  OAI22_X1 U17269 ( .A1(n16125), .A2(n18988), .B1(n16068), .B2(n18979), .ZN(
        n13902) );
  OAI22_X1 U17270 ( .A1(n16088), .A2(n18980), .B1(n9889), .B2(n13900), .ZN(
        n13901) );
  AOI211_X1 U17271 ( .C1(n13903), .C2(n16120), .A(n13902), .B(n13901), .ZN(
        n13904) );
  OAI21_X1 U17272 ( .B1(n15067), .B2(n13905), .A(n13904), .ZN(P2_U3009) );
  INV_X1 U17273 ( .A(DATAI_8_), .ZN(n13907) );
  INV_X1 U17274 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n13906) );
  MUX2_X1 U17275 ( .A(n13907), .B(n13906), .S(n20092), .Z(n19998) );
  INV_X1 U17276 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n13908) );
  OAI222_X1 U17277 ( .A1(n14296), .A2(n14141), .B1(n14297), .B2(n19998), .C1(
        n13908), .C2(n14294), .ZN(P1_U2896) );
  NOR2_X1 U17278 ( .A1(n13910), .A2(n13911), .ZN(n13912) );
  OR2_X1 U17279 ( .A1(n13909), .A2(n13912), .ZN(n19007) );
  AOI21_X1 U17280 ( .B1(n13914), .B2(n13913), .A(n9870), .ZN(n18876) );
  OAI22_X1 U17281 ( .A1(n19092), .A2(n14841), .B1(n19044), .B2(n13915), .ZN(
        n13916) );
  AOI21_X1 U17282 ( .B1(n19084), .B2(n18876), .A(n13916), .ZN(n13918) );
  AOI22_X1 U17283 ( .A1(n16048), .A2(BUF2_REG_16__SCAN_IN), .B1(n16049), .B2(
        BUF1_REG_16__SCAN_IN), .ZN(n13917) );
  OAI211_X1 U17284 ( .C1(n19007), .C2(n19079), .A(n13918), .B(n13917), .ZN(
        P2_U2903) );
  OAI21_X1 U17285 ( .B1(n13894), .B2(n13919), .A(n13196), .ZN(n19889) );
  INV_X1 U17286 ( .A(DATAI_9_), .ZN(n13921) );
  INV_X1 U17287 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n13920) );
  MUX2_X1 U17288 ( .A(n13921), .B(n13920), .S(n20092), .Z(n20001) );
  INV_X1 U17289 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n13922) );
  OAI222_X1 U17290 ( .A1(n14296), .A2(n19889), .B1(n14297), .B2(n20001), .C1(
        n13922), .C2(n14294), .ZN(P1_U2895) );
  XNOR2_X1 U17291 ( .A(n13924), .B(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13925) );
  XNOR2_X1 U17292 ( .A(n13923), .B(n13925), .ZN(n15899) );
  AOI22_X1 U17293 ( .A1(n20043), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        n11744), .B2(P1_REIP_REG_8__SCAN_IN), .ZN(n13926) );
  OAI21_X1 U17294 ( .B1(n20041), .B2(n14133), .A(n13926), .ZN(n13927) );
  AOI21_X1 U17295 ( .B1(n13928), .B2(n20038), .A(n13927), .ZN(n13929) );
  OAI21_X1 U17296 ( .B1(n15899), .B2(n19867), .A(n13929), .ZN(P1_U2991) );
  OAI22_X1 U17297 ( .A1(n15737), .A2(n15879), .B1(n13930), .B2(n19966), .ZN(
        n13931) );
  AOI21_X1 U17298 ( .B1(n14436), .B2(n13156), .A(n13931), .ZN(n13932) );
  INV_X1 U17299 ( .A(n13932), .ZN(P1_U2862) );
  INV_X1 U17300 ( .A(DATAI_10_), .ZN(n13933) );
  MUX2_X1 U17301 ( .A(n13933), .B(n16353), .S(n20092), .Z(n20004) );
  INV_X1 U17302 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n13934) );
  OAI222_X1 U17303 ( .A1(n14296), .A2(n13935), .B1(n14297), .B2(n20004), .C1(
        n13934), .C2(n14294), .ZN(P1_U2894) );
  MUX2_X1 U17304 ( .A(n13937), .B(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .S(
        n14352), .Z(n13938) );
  XNOR2_X1 U17305 ( .A(n13936), .B(n13938), .ZN(n15888) );
  INV_X1 U17306 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n13940) );
  INV_X1 U17307 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n13939) );
  OAI22_X1 U17308 ( .A1(n14425), .A2(n13940), .B1(n20081), .B2(n13939), .ZN(
        n13942) );
  NOR2_X1 U17309 ( .A1(n19889), .A2(n20094), .ZN(n13941) );
  AOI211_X1 U17310 ( .C1(n20045), .C2(n19890), .A(n13942), .B(n13941), .ZN(
        n13943) );
  OAI21_X1 U17311 ( .B1(n15888), .B2(n19867), .A(n13943), .ZN(P1_U2990) );
  INV_X1 U17312 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n18561) );
  NAND3_X1 U17313 ( .A1(n17027), .A2(n15540), .A3(n18561), .ZN(n18100) );
  NOR2_X1 U17314 ( .A1(P3_FLUSH_REG_SCAN_IN), .A2(n18100), .ZN(n13944) );
  NAND3_X1 U17315 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_0__SCAN_IN), .A3(P3_STATE2_REG_2__SCAN_IN), .ZN(n18714)
         );
  OAI21_X1 U17316 ( .B1(n13944), .B2(n18714), .A(n18401), .ZN(n18110) );
  INV_X1 U17317 ( .A(n18110), .ZN(n13945) );
  NOR2_X1 U17318 ( .A1(n17735), .A2(n18766), .ZN(n18104) );
  AOI21_X1 U17319 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n18104), .ZN(n18105) );
  NOR2_X1 U17320 ( .A1(n13945), .A2(n18105), .ZN(n13947) );
  INV_X1 U17321 ( .A(n18456), .ZN(n18191) );
  NOR2_X1 U17322 ( .A1(n18716), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18149) );
  OR2_X1 U17323 ( .A1(n18149), .A2(n13945), .ZN(n18103) );
  OR2_X1 U17324 ( .A1(n18191), .A2(n18103), .ZN(n13946) );
  MUX2_X1 U17325 ( .A(n13947), .B(n13946), .S(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .Z(P3_U2864) );
  OAI22_X1 U17326 ( .A1(n20217), .A2(n13948), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n14548), .ZN(n15583) );
  OAI22_X1 U17327 ( .A1(n15937), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n15613), .ZN(n13949) );
  AOI21_X1 U17328 ( .B1(n15583), .B2(n14552), .A(n13949), .ZN(n13953) );
  AOI21_X1 U17329 ( .B1(n13950), .B2(n14552), .A(n13952), .ZN(n13951) );
  OAI22_X1 U17330 ( .A1(n13953), .A2(n13952), .B1(n13951), .B2(n11132), .ZN(
        P1_U3474) );
  NOR2_X1 U17331 ( .A1(n15137), .A2(n19037), .ZN(n13954) );
  AOI21_X1 U17332 ( .B1(P2_EBX_REG_30__SCAN_IN), .B2(n19037), .A(n13954), .ZN(
        n13955) );
  OAI21_X1 U17333 ( .B1(n13956), .B2(n19031), .A(n13955), .ZN(P2_U2857) );
  NAND2_X1 U17334 ( .A1(n14294), .A2(n13957), .ZN(n13967) );
  INV_X1 U17335 ( .A(n13967), .ZN(n13958) );
  NAND2_X1 U17336 ( .A1(n13958), .A2(n20092), .ZN(n14265) );
  INV_X1 U17337 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n16318) );
  NAND2_X1 U17338 ( .A1(n13995), .A2(n13959), .ZN(n13964) );
  AOI22_X1 U17339 ( .A1(n13961), .A2(P1_EAX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n13960), .ZN(n13962) );
  INV_X1 U17340 ( .A(n13962), .ZN(n13963) );
  AND2_X1 U17341 ( .A1(n14294), .A2(n13965), .ZN(n13966) );
  NAND2_X1 U17342 ( .A1(n13977), .A2(n13966), .ZN(n13970) );
  AOI22_X1 U17343 ( .A1(n13968), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n14298), .ZN(n13969) );
  OAI211_X1 U17344 ( .C1(n14265), .C2(n16318), .A(n13970), .B(n13969), .ZN(
        P1_U2873) );
  AOI21_X1 U17345 ( .B1(n20043), .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n13971), .ZN(n13972) );
  OAI21_X1 U17346 ( .B1(n20041), .B2(n13973), .A(n13972), .ZN(n13974) );
  OAI21_X1 U17347 ( .B1(n13976), .B2(n19867), .A(n13975), .ZN(P1_U2968) );
  INV_X1 U17348 ( .A(n13977), .ZN(n13984) );
  INV_X1 U17349 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n15654) );
  INV_X1 U17350 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n14012) );
  INV_X1 U17351 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n13978) );
  INV_X1 U17352 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n20732) );
  INV_X1 U17353 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n20728) );
  INV_X1 U17354 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n20722) );
  NAND3_X1 U17355 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(P1_REIP_REG_12__SCAN_IN), 
        .A3(n15720), .ZN(n14121) );
  NOR2_X1 U17356 ( .A1(n20722), .A2(n14121), .ZN(n14103) );
  NAND2_X1 U17357 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(n14103), .ZN(n14072) );
  NAND2_X1 U17358 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(P1_REIP_REG_15__SCAN_IN), 
        .ZN(n14075) );
  NOR3_X1 U17359 ( .A1(n20728), .A2(n14072), .A3(n14075), .ZN(n14051) );
  NAND3_X1 U17360 ( .A1(n14051), .A2(P1_REIP_REG_19__SCAN_IN), .A3(
        P1_REIP_REG_18__SCAN_IN), .ZN(n14037) );
  NAND2_X1 U17361 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(P1_REIP_REG_20__SCAN_IN), 
        .ZN(n14036) );
  NOR4_X1 U17362 ( .A1(n13978), .A2(n20732), .A3(n14037), .A4(n14036), .ZN(
        n14011) );
  NAND2_X1 U17363 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(n14011), .ZN(n14013) );
  NOR2_X1 U17364 ( .A1(n14012), .A2(n14013), .ZN(n15669) );
  NAND2_X1 U17365 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(n15669), .ZN(n15668) );
  NOR2_X1 U17366 ( .A1(n15654), .A2(n15668), .ZN(n15655) );
  NAND2_X1 U17367 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(n15655), .ZN(n15642) );
  INV_X1 U17368 ( .A(n15642), .ZN(n13997) );
  NAND4_X1 U17369 ( .A1(n19924), .A2(P1_REIP_REG_30__SCAN_IN), .A3(
        P1_REIP_REG_29__SCAN_IN), .A4(n13997), .ZN(n13979) );
  NAND2_X1 U17370 ( .A1(n14074), .A2(n13979), .ZN(n13987) );
  NOR3_X1 U17371 ( .A1(n19926), .A2(n15642), .A3(n20745), .ZN(n13986) );
  NAND3_X1 U17372 ( .A1(n13986), .A2(P1_REIP_REG_30__SCAN_IN), .A3(n20749), 
        .ZN(n13981) );
  AOI22_X1 U17373 ( .A1(n19937), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n19940), .ZN(n13980) );
  OAI211_X1 U17374 ( .C1(n13987), .C2(n20749), .A(n13981), .B(n13980), .ZN(
        n13982) );
  AOI21_X1 U17375 ( .B1(n14142), .B2(n19948), .A(n13982), .ZN(n13983) );
  OAI21_X1 U17376 ( .B1(n13984), .B2(n15726), .A(n13983), .ZN(P1_U2809) );
  NAND2_X1 U17377 ( .A1(n14307), .A2(n19912), .ZN(n13993) );
  INV_X1 U17378 ( .A(n14306), .ZN(n13985) );
  OAI22_X1 U17379 ( .A1(n14303), .A2(n15730), .B1(n19957), .B2(n13985), .ZN(
        n13991) );
  INV_X1 U17380 ( .A(n13986), .ZN(n13989) );
  AOI21_X1 U17381 ( .B1(n13989), .B2(n13988), .A(n13987), .ZN(n13990) );
  AOI211_X1 U17382 ( .C1(n19937), .C2(P1_EBX_REG_30__SCAN_IN), .A(n13991), .B(
        n13990), .ZN(n13992) );
  OAI211_X1 U17383 ( .C1(n19897), .C2(n13994), .A(n13993), .B(n13992), .ZN(
        P1_U2810) );
  AOI21_X1 U17384 ( .B1(n13996), .B2(n13171), .A(n13995), .ZN(n14315) );
  NAND2_X1 U17385 ( .A1(n14315), .A2(n19912), .ZN(n14003) );
  OAI21_X1 U17386 ( .B1(n19926), .B2(n13997), .A(n19924), .ZN(n15643) );
  NOR3_X1 U17387 ( .A1(n19926), .A2(P1_REIP_REG_29__SCAN_IN), .A3(n15642), 
        .ZN(n14001) );
  INV_X1 U17388 ( .A(n14313), .ZN(n13998) );
  AOI22_X1 U17389 ( .A1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n19940), .B1(
        n19891), .B2(n13998), .ZN(n13999) );
  OAI21_X1 U17390 ( .B1(n19899), .B2(n14146), .A(n13999), .ZN(n14000) );
  AOI211_X1 U17391 ( .C1(P1_REIP_REG_29__SCAN_IN), .C2(n15643), .A(n14001), 
        .B(n14000), .ZN(n14002) );
  OAI211_X1 U17392 ( .C1(n19897), .C2(n14145), .A(n14003), .B(n14002), .ZN(
        P1_U2811) );
  INV_X1 U17393 ( .A(n14004), .ZN(n14022) );
  AND2_X1 U17394 ( .A1(n14022), .A2(n14005), .ZN(n14007) );
  OR2_X1 U17395 ( .A1(n14007), .A2(n14006), .ZN(n14338) );
  OR2_X1 U17396 ( .A1(n14026), .A2(n14009), .ZN(n14010) );
  NAND2_X1 U17397 ( .A1(n14008), .A2(n14010), .ZN(n14465) );
  NOR2_X1 U17398 ( .A1(n14465), .A2(n19897), .ZN(n14018) );
  INV_X1 U17399 ( .A(n14011), .ZN(n14028) );
  OAI21_X1 U17400 ( .B1(n19895), .B2(n14028), .A(n14074), .ZN(n15681) );
  INV_X1 U17401 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n14029) );
  NAND2_X1 U17402 ( .A1(n19950), .A2(n14029), .ZN(n14027) );
  AOI21_X1 U17403 ( .B1(n15681), .B2(n14027), .A(n14012), .ZN(n14017) );
  NOR3_X1 U17404 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(n19926), .A3(n14013), 
        .ZN(n14016) );
  INV_X1 U17405 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n14162) );
  AOI22_X1 U17406 ( .A1(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n19940), .B1(
        n19891), .B2(n14341), .ZN(n14014) );
  OAI21_X1 U17407 ( .B1(n19899), .B2(n14162), .A(n14014), .ZN(n14015) );
  NOR4_X1 U17408 ( .A1(n14018), .A2(n14017), .A3(n14016), .A4(n14015), .ZN(
        n14019) );
  OAI21_X1 U17409 ( .B1(n14338), .B2(n15726), .A(n14019), .ZN(P1_U2815) );
  BUF_X1 U17410 ( .A(n14020), .Z(n14021) );
  OR2_X1 U17411 ( .A1(n14021), .A2(n14170), .ZN(n14168) );
  AOI21_X1 U17412 ( .B1(n14023), .B2(n14168), .A(n14004), .ZN(n14349) );
  INV_X1 U17413 ( .A(n14349), .ZN(n14252) );
  AND2_X1 U17414 ( .A1(n14174), .A2(n14024), .ZN(n14025) );
  NOR2_X1 U17415 ( .A1(n14026), .A2(n14025), .ZN(n14473) );
  OAI22_X1 U17416 ( .A1(n15681), .A2(n14029), .B1(n14028), .B2(n14027), .ZN(
        n14032) );
  AOI22_X1 U17417 ( .A1(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n19940), .B1(
        n19891), .B2(n14348), .ZN(n14030) );
  OAI21_X1 U17418 ( .B1(n19899), .B2(n14165), .A(n14030), .ZN(n14031) );
  AOI211_X1 U17419 ( .C1(n14473), .C2(n19948), .A(n14032), .B(n14031), .ZN(
        n14033) );
  OAI21_X1 U17420 ( .B1(n14252), .B2(n15726), .A(n14033), .ZN(P1_U2816) );
  OAI21_X1 U17421 ( .B1(n14034), .B2(n14035), .A(n14021), .ZN(n14361) );
  NAND4_X1 U17422 ( .A1(n19950), .A2(n14051), .A3(P1_REIP_REG_19__SCAN_IN), 
        .A4(P1_REIP_REG_18__SCAN_IN), .ZN(n15697) );
  NOR2_X1 U17423 ( .A1(n14036), .A2(n15697), .ZN(n15680) );
  INV_X1 U17424 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n21011) );
  INV_X1 U17425 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n15698) );
  OR2_X1 U17426 ( .A1(n14037), .A2(n15698), .ZN(n15689) );
  OAI21_X1 U17427 ( .B1(n19895), .B2(n15689), .A(n14074), .ZN(n15696) );
  OAI21_X1 U17428 ( .B1(P1_REIP_REG_21__SCAN_IN), .B2(n19926), .A(n15696), 
        .ZN(n14038) );
  AOI22_X1 U17429 ( .A1(n19940), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B1(
        P1_REIP_REG_22__SCAN_IN), .B2(n14038), .ZN(n14040) );
  NAND2_X1 U17430 ( .A1(n19891), .A2(n14362), .ZN(n14039) );
  OAI211_X1 U17431 ( .C1(n19899), .C2(n21011), .A(n14040), .B(n14039), .ZN(
        n14043) );
  INV_X1 U17432 ( .A(n14041), .ZN(n14173) );
  XNOR2_X1 U17433 ( .A(n14494), .B(n14173), .ZN(n15807) );
  NOR2_X1 U17434 ( .A1(n15807), .A2(n19897), .ZN(n14042) );
  AOI211_X1 U17435 ( .C1(n20732), .C2(n15680), .A(n14043), .B(n14042), .ZN(
        n14044) );
  OAI21_X1 U17436 ( .B1(n14361), .B2(n15726), .A(n14044), .ZN(P1_U2818) );
  OAI21_X1 U17437 ( .B1(n14045), .B2(n14047), .A(n14046), .ZN(n14389) );
  AND2_X1 U17438 ( .A1(n14061), .A2(n14048), .ZN(n14049) );
  OR2_X1 U17439 ( .A1(n14049), .A2(n14187), .ZN(n15822) );
  INV_X1 U17440 ( .A(n15822), .ZN(n14055) );
  AOI21_X1 U17441 ( .B1(n19891), .B2(n14392), .A(n19909), .ZN(n14050) );
  OAI21_X1 U17442 ( .B1(n14388), .B2(n15730), .A(n14050), .ZN(n14054) );
  NAND2_X1 U17443 ( .A1(n19950), .A2(n14051), .ZN(n15711) );
  OAI21_X1 U17444 ( .B1(n19926), .B2(n14051), .A(n19924), .ZN(n15708) );
  AOI22_X1 U17445 ( .A1(n15708), .A2(P1_REIP_REG_18__SCAN_IN), .B1(n19937), 
        .B2(P1_EBX_REG_18__SCAN_IN), .ZN(n14052) );
  OAI21_X1 U17446 ( .B1(P1_REIP_REG_18__SCAN_IN), .B2(n15711), .A(n14052), 
        .ZN(n14053) );
  AOI211_X1 U17447 ( .C1(n14055), .C2(n19948), .A(n14054), .B(n14053), .ZN(
        n14056) );
  OAI21_X1 U17448 ( .B1(n14389), .B2(n15726), .A(n14056), .ZN(P1_U2822) );
  NOR2_X1 U17449 ( .A1(n14058), .A2(n14059), .ZN(n14060) );
  AOI21_X1 U17450 ( .B1(n14062), .B2(n14081), .A(n11673), .ZN(n14515) );
  INV_X1 U17451 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n14065) );
  AOI21_X1 U17452 ( .B1(n19891), .B2(n15755), .A(n19909), .ZN(n14064) );
  NAND2_X1 U17453 ( .A1(n19937), .A2(P1_EBX_REG_17__SCAN_IN), .ZN(n14063) );
  OAI211_X1 U17454 ( .C1(n15730), .C2(n14065), .A(n14064), .B(n14063), .ZN(
        n14066) );
  AOI21_X1 U17455 ( .B1(n14515), .B2(n19948), .A(n14066), .ZN(n14069) );
  OR2_X1 U17456 ( .A1(n19926), .A2(n14072), .ZN(n14093) );
  OAI21_X1 U17457 ( .B1(n14075), .B2(n14093), .A(n20728), .ZN(n14067) );
  NAND2_X1 U17458 ( .A1(n14067), .A2(n15708), .ZN(n14068) );
  OAI211_X1 U17459 ( .C1(n15754), .C2(n15726), .A(n14069), .B(n14068), .ZN(
        P1_U2823) );
  AOI21_X1 U17460 ( .B1(n14071), .B2(n14087), .A(n14058), .ZN(n14404) );
  INV_X1 U17461 ( .A(n14404), .ZN(n14288) );
  INV_X1 U17462 ( .A(n14072), .ZN(n14073) );
  NAND2_X1 U17463 ( .A1(n19924), .A2(n14073), .ZN(n14104) );
  NAND2_X1 U17464 ( .A1(n14074), .A2(n14104), .ZN(n14114) );
  INV_X1 U17465 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n21103) );
  OAI21_X1 U17466 ( .B1(P1_REIP_REG_16__SCAN_IN), .B2(P1_REIP_REG_15__SCAN_IN), 
        .A(n14075), .ZN(n14076) );
  OAI22_X1 U17467 ( .A1(n14114), .A2(n21103), .B1(n14093), .B2(n14076), .ZN(
        n14084) );
  INV_X1 U17468 ( .A(n14077), .ZN(n14402) );
  AOI21_X1 U17469 ( .B1(n19940), .B2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n19909), .ZN(n14078) );
  OAI21_X1 U17470 ( .B1(n14402), .B2(n19957), .A(n14078), .ZN(n14083) );
  OR2_X1 U17471 ( .A1(n14089), .A2(n14079), .ZN(n14080) );
  NAND2_X1 U17472 ( .A1(n14081), .A2(n14080), .ZN(n15832) );
  OAI22_X1 U17473 ( .A1(n15832), .A2(n19897), .B1(n14195), .B2(n19899), .ZN(
        n14082) );
  NOR3_X1 U17474 ( .A1(n14084), .A2(n14083), .A3(n14082), .ZN(n14085) );
  OAI21_X1 U17475 ( .B1(n14288), .B2(n15726), .A(n14085), .ZN(P1_U2824) );
  AOI21_X1 U17476 ( .B1(n14088), .B2(n14086), .A(n14070), .ZN(n15761) );
  INV_X1 U17477 ( .A(n15761), .ZN(n14290) );
  AOI21_X1 U17478 ( .B1(n14090), .B2(n14101), .A(n14089), .ZN(n14530) );
  AOI22_X1 U17479 ( .A1(n19937), .A2(P1_EBX_REG_15__SCAN_IN), .B1(n19891), 
        .B2(n15760), .ZN(n14091) );
  INV_X1 U17480 ( .A(n14091), .ZN(n14095) );
  INV_X1 U17481 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n20724) );
  AOI21_X1 U17482 ( .B1(n19940), .B2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n19909), .ZN(n14092) );
  OAI221_X1 U17483 ( .B1(P1_REIP_REG_15__SCAN_IN), .B2(n14093), .C1(n20724), 
        .C2(n14114), .A(n14092), .ZN(n14094) );
  AOI211_X1 U17484 ( .C1(n14530), .C2(n19948), .A(n14095), .B(n14094), .ZN(
        n14096) );
  OAI21_X1 U17485 ( .B1(n14290), .B2(n15726), .A(n14096), .ZN(P1_U2825) );
  INV_X1 U17486 ( .A(n14086), .ZN(n14098) );
  INV_X1 U17487 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n14113) );
  NAND2_X1 U17488 ( .A1(n14122), .A2(n14099), .ZN(n14100) );
  NAND2_X1 U17489 ( .A1(n14101), .A2(n14100), .ZN(n15840) );
  INV_X1 U17490 ( .A(n15840), .ZN(n14102) );
  AOI22_X1 U17491 ( .A1(n14102), .A2(n19948), .B1(n19937), .B2(
        P1_EBX_REG_14__SCAN_IN), .ZN(n14112) );
  NAND2_X1 U17492 ( .A1(n14104), .A2(n14103), .ZN(n14109) );
  NAND2_X1 U17493 ( .A1(n19940), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n14105) );
  AND2_X1 U17494 ( .A1(n14105), .A2(n19942), .ZN(n14108) );
  INV_X1 U17495 ( .A(n14412), .ZN(n14106) );
  NAND2_X1 U17496 ( .A1(n19891), .A2(n14106), .ZN(n14107) );
  OAI211_X1 U17497 ( .C1(n19926), .C2(n14109), .A(n14108), .B(n14107), .ZN(
        n14110) );
  INV_X1 U17498 ( .A(n14110), .ZN(n14111) );
  OAI211_X1 U17499 ( .C1(n14114), .C2(n14113), .A(n14112), .B(n14111), .ZN(
        n14115) );
  AOI21_X1 U17500 ( .B1(n14414), .B2(n19912), .A(n14115), .ZN(n14116) );
  INV_X1 U17501 ( .A(n14116), .ZN(P1_U2826) );
  NAND2_X1 U17502 ( .A1(n13198), .A2(n14118), .ZN(n14119) );
  NAND2_X1 U17503 ( .A1(n14117), .A2(n14119), .ZN(n14214) );
  OAI21_X1 U17504 ( .B1(n14214), .B2(n14215), .A(n14117), .ZN(n14210) );
  INV_X1 U17505 ( .A(n14121), .ZN(n14124) );
  OAI21_X1 U17506 ( .B1(n19926), .B2(n14124), .A(n19924), .ZN(n15723) );
  OAI21_X1 U17507 ( .B1(n14205), .B2(n14123), .A(n14122), .ZN(n14202) );
  AOI22_X1 U17508 ( .A1(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n19940), .B1(
        n19937), .B2(P1_EBX_REG_13__SCAN_IN), .ZN(n14126) );
  NAND3_X1 U17509 ( .A1(n19950), .A2(n20722), .A3(n14124), .ZN(n14125) );
  NAND2_X1 U17510 ( .A1(n14126), .A2(n14125), .ZN(n14127) );
  AOI211_X1 U17511 ( .C1(n14427), .C2(n19891), .A(n14127), .B(n19909), .ZN(
        n14128) );
  OAI21_X1 U17512 ( .B1(n19897), .B2(n14202), .A(n14128), .ZN(n14129) );
  AOI21_X1 U17513 ( .B1(P1_REIP_REG_13__SCAN_IN), .B2(n15723), .A(n14129), 
        .ZN(n14130) );
  OAI21_X1 U17514 ( .B1(n14430), .B2(n15726), .A(n14130), .ZN(P1_U2827) );
  NOR2_X1 U17515 ( .A1(n19926), .A2(n19923), .ZN(n19922) );
  NOR2_X1 U17516 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n14131), .ZN(n14139) );
  OAI22_X1 U17517 ( .A1(n14133), .A2(n19957), .B1(n15730), .B2(n14132), .ZN(
        n14134) );
  AOI21_X1 U17518 ( .B1(P1_EBX_REG_8__SCAN_IN), .B2(n19937), .A(n14134), .ZN(
        n14135) );
  OAI21_X1 U17519 ( .B1(n19897), .B2(n15902), .A(n14135), .ZN(n14138) );
  OAI21_X1 U17520 ( .B1(n19926), .B2(n19885), .A(n19924), .ZN(n14136) );
  INV_X1 U17521 ( .A(n14136), .ZN(n19894) );
  OAI21_X1 U17522 ( .B1(n19894), .B2(n15901), .A(n19942), .ZN(n14137) );
  AOI211_X1 U17523 ( .C1(n19922), .C2(n14139), .A(n14138), .B(n14137), .ZN(
        n14140) );
  OAI21_X1 U17524 ( .B1(n14141), .B2(n15726), .A(n14140), .ZN(P1_U2832) );
  INV_X1 U17525 ( .A(n14142), .ZN(n14144) );
  OAI22_X1 U17526 ( .A1(n14144), .A2(n15737), .B1(n19966), .B2(n14143), .ZN(
        P1_U2841) );
  INV_X1 U17527 ( .A(n14315), .ZN(n14234) );
  OAI222_X1 U17528 ( .A1(n14213), .A2(n14234), .B1(n14146), .B2(n19966), .C1(
        n14145), .C2(n15737), .ZN(P1_U2843) );
  NOR2_X1 U17529 ( .A1(n14148), .A2(n14147), .ZN(n14149) );
  OAI22_X1 U17530 ( .A1(n15649), .A2(n15737), .B1(n15644), .B2(n19966), .ZN(
        n14150) );
  INV_X1 U17531 ( .A(n14150), .ZN(n14151) );
  OAI21_X1 U17532 ( .B1(n15650), .B2(n14213), .A(n14151), .ZN(P1_U2844) );
  AOI21_X1 U17533 ( .B1(n14153), .B2(n14152), .A(n13169), .ZN(n15664) );
  INV_X1 U17534 ( .A(n15664), .ZN(n14242) );
  INV_X1 U17535 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n14155) );
  XNOR2_X1 U17536 ( .A(n9854), .B(n14154), .ZN(n15662) );
  OAI222_X1 U17537 ( .A1(n14213), .A2(n14242), .B1(n14155), .B2(n19966), .C1(
        n15662), .C2(n15737), .ZN(P1_U2845) );
  NAND2_X1 U17538 ( .A1(n14008), .A2(n14157), .ZN(n14158) );
  AND2_X1 U17539 ( .A1(n9854), .A2(n14158), .ZN(n15673) );
  NOR2_X1 U17540 ( .A1(n19966), .A2(n14159), .ZN(n14160) );
  AOI21_X1 U17541 ( .B1(n15673), .B2(n19962), .A(n14160), .ZN(n14161) );
  OAI21_X1 U17542 ( .B1(n15675), .B2(n14213), .A(n14161), .ZN(P1_U2846) );
  OAI22_X1 U17543 ( .A1(n14465), .A2(n15737), .B1(n14162), .B2(n19966), .ZN(
        n14163) );
  INV_X1 U17544 ( .A(n14163), .ZN(n14164) );
  OAI21_X1 U17545 ( .B1(n14338), .B2(n14213), .A(n14164), .ZN(P1_U2847) );
  NOR2_X1 U17546 ( .A1(n19966), .A2(n14165), .ZN(n14166) );
  AOI21_X1 U17547 ( .B1(n14473), .B2(n19962), .A(n14166), .ZN(n14167) );
  OAI21_X1 U17548 ( .B1(n14252), .B2(n14213), .A(n14167), .ZN(P1_U2848) );
  INV_X1 U17549 ( .A(n14168), .ZN(n14169) );
  AOI21_X1 U17550 ( .B1(n14170), .B2(n14021), .A(n14169), .ZN(n15685) );
  INV_X1 U17551 ( .A(n15685), .ZN(n14256) );
  INV_X1 U17552 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n14176) );
  INV_X1 U17553 ( .A(n14171), .ZN(n14172) );
  OAI21_X1 U17554 ( .B1(n14494), .B2(n14173), .A(n14172), .ZN(n14175) );
  NAND2_X1 U17555 ( .A1(n14175), .A2(n14174), .ZN(n15683) );
  OAI222_X1 U17556 ( .A1(n14213), .A2(n14256), .B1(n14176), .B2(n19966), .C1(
        n15683), .C2(n15737), .ZN(P1_U2849) );
  OAI222_X1 U17557 ( .A1(n14213), .A2(n14361), .B1(n19966), .B2(n21011), .C1(
        n15737), .C2(n15807), .ZN(P1_U2850) );
  AND2_X1 U17558 ( .A1(n14177), .A2(n14178), .ZN(n14180) );
  OR2_X1 U17559 ( .A1(n14180), .A2(n14179), .ZN(n15701) );
  INV_X1 U17560 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n14183) );
  OR2_X1 U17561 ( .A1(n14189), .A2(n14181), .ZN(n14182) );
  AND2_X1 U17562 ( .A1(n14492), .A2(n14182), .ZN(n14503) );
  INV_X1 U17563 ( .A(n14503), .ZN(n15700) );
  OAI222_X1 U17564 ( .A1(n14213), .A2(n15701), .B1(n19966), .B2(n14183), .C1(
        n15700), .C2(n15737), .ZN(P1_U2852) );
  NAND2_X1 U17565 ( .A1(n14046), .A2(n14184), .ZN(n14185) );
  AND2_X1 U17566 ( .A1(n14177), .A2(n14185), .ZN(n15750) );
  INV_X1 U17567 ( .A(n15750), .ZN(n14275) );
  INV_X1 U17568 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n14190) );
  NOR2_X1 U17569 ( .A1(n14187), .A2(n14186), .ZN(n14188) );
  OR2_X1 U17570 ( .A1(n14189), .A2(n14188), .ZN(n15713) );
  OAI222_X1 U17571 ( .A1(n14213), .A2(n14275), .B1(n14190), .B2(n19966), .C1(
        n15713), .C2(n15737), .ZN(P1_U2853) );
  OAI22_X1 U17572 ( .A1(n15822), .A2(n15737), .B1(n14191), .B2(n19966), .ZN(
        n14192) );
  INV_X1 U17573 ( .A(n14192), .ZN(n14193) );
  OAI21_X1 U17574 ( .B1(n14389), .B2(n14213), .A(n14193), .ZN(P1_U2854) );
  AOI22_X1 U17575 ( .A1(n14515), .A2(n19962), .B1(P1_EBX_REG_17__SCAN_IN), 
        .B2(n14203), .ZN(n14194) );
  OAI21_X1 U17576 ( .B1(n15754), .B2(n14213), .A(n14194), .ZN(P1_U2855) );
  OAI22_X1 U17577 ( .A1(n15832), .A2(n15737), .B1(n14195), .B2(n19966), .ZN(
        n14196) );
  INV_X1 U17578 ( .A(n14196), .ZN(n14197) );
  OAI21_X1 U17579 ( .B1(n14288), .B2(n14213), .A(n14197), .ZN(P1_U2856) );
  AOI22_X1 U17580 ( .A1(n14530), .A2(n19962), .B1(P1_EBX_REG_15__SCAN_IN), 
        .B2(n14203), .ZN(n14198) );
  OAI21_X1 U17581 ( .B1(n14290), .B2(n14213), .A(n14198), .ZN(P1_U2857) );
  OAI22_X1 U17582 ( .A1(n15840), .A2(n15737), .B1(n14199), .B2(n19966), .ZN(
        n14200) );
  AOI21_X1 U17583 ( .B1(n14414), .B2(n13156), .A(n14200), .ZN(n14201) );
  INV_X1 U17584 ( .A(n14201), .ZN(P1_U2858) );
  INV_X1 U17585 ( .A(n14202), .ZN(n15843) );
  AOI22_X1 U17586 ( .A1(n15843), .A2(n19962), .B1(P1_EBX_REG_13__SCAN_IN), 
        .B2(n14203), .ZN(n14204) );
  OAI21_X1 U17587 ( .B1(n14430), .B2(n14213), .A(n14204), .ZN(P1_U2859) );
  INV_X1 U17588 ( .A(n14205), .ZN(n14208) );
  NAND2_X1 U17589 ( .A1(n14219), .A2(n14206), .ZN(n14207) );
  NAND2_X1 U17590 ( .A1(n14208), .A2(n14207), .ZN(n15862) );
  INV_X1 U17591 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n20973) );
  NOR2_X1 U17592 ( .A1(n14210), .A2(n14209), .ZN(n14211) );
  OAI222_X1 U17593 ( .A1(n15862), .A2(n15737), .B1(n19966), .B2(n20973), .C1(
        n15769), .C2(n14213), .ZN(P1_U2860) );
  INV_X1 U17594 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n21031) );
  XOR2_X1 U17595 ( .A(n14215), .B(n14214), .Z(n15777) );
  NAND2_X1 U17596 ( .A1(n15777), .A2(n13156), .ZN(n14221) );
  NAND2_X1 U17597 ( .A1(n14217), .A2(n14216), .ZN(n14218) );
  AND2_X1 U17598 ( .A1(n14219), .A2(n14218), .ZN(n15863) );
  NAND2_X1 U17599 ( .A1(n19962), .A2(n15863), .ZN(n14220) );
  OAI211_X1 U17600 ( .C1(n21031), .C2(n19966), .A(n14221), .B(n14220), .ZN(
        P1_U2861) );
  NAND3_X1 U17601 ( .A1(n14294), .A2(n14222), .A3(n9790), .ZN(n14283) );
  INV_X1 U17602 ( .A(DATAI_14_), .ZN(n14224) );
  MUX2_X1 U17603 ( .A(n14224), .B(n14223), .S(n20092), .Z(n20013) );
  OAI22_X1 U17604 ( .A1(n14283), .A2(n20013), .B1(n14294), .B2(n13516), .ZN(
        n14225) );
  AOI21_X1 U17605 ( .B1(BUF1_REG_30__SCAN_IN), .B2(n14285), .A(n14225), .ZN(
        n14227) );
  NAND2_X1 U17606 ( .A1(n13968), .A2(DATAI_30_), .ZN(n14226) );
  OAI211_X1 U17607 ( .C1(n14228), .C2(n14296), .A(n14227), .B(n14226), .ZN(
        P1_U2874) );
  INV_X1 U17608 ( .A(DATAI_13_), .ZN(n14230) );
  MUX2_X1 U17609 ( .A(n14230), .B(n14229), .S(n20092), .Z(n20010) );
  OAI22_X1 U17610 ( .A1(n14283), .A2(n20010), .B1(n14294), .B2(n13524), .ZN(
        n14231) );
  AOI21_X1 U17611 ( .B1(BUF1_REG_29__SCAN_IN), .B2(n14285), .A(n14231), .ZN(
        n14233) );
  NAND2_X1 U17612 ( .A1(n13968), .A2(DATAI_29_), .ZN(n14232) );
  OAI211_X1 U17613 ( .C1(n14234), .C2(n14296), .A(n14233), .B(n14232), .ZN(
        P1_U2875) );
  INV_X1 U17614 ( .A(DATAI_12_), .ZN(n14235) );
  INV_X1 U17615 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n21043) );
  MUX2_X1 U17616 ( .A(n14235), .B(n21043), .S(n20092), .Z(n20007) );
  OAI22_X1 U17617 ( .A1(n14283), .A2(n20007), .B1(n14294), .B2(n13522), .ZN(
        n14236) );
  AOI21_X1 U17618 ( .B1(BUF1_REG_28__SCAN_IN), .B2(n14285), .A(n14236), .ZN(
        n14238) );
  NAND2_X1 U17619 ( .A1(n13968), .A2(DATAI_28_), .ZN(n14237) );
  OAI211_X1 U17620 ( .C1(n15650), .C2(n14296), .A(n14238), .B(n14237), .ZN(
        P1_U2876) );
  INV_X1 U17621 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n16325) );
  INV_X1 U17622 ( .A(n14283), .ZN(n14263) );
  AOI22_X1 U17623 ( .A1(n14263), .A2(n14299), .B1(P1_EAX_REG_27__SCAN_IN), 
        .B2(n14298), .ZN(n14239) );
  OAI21_X1 U17624 ( .B1(n16325), .B2(n14265), .A(n14239), .ZN(n14240) );
  AOI21_X1 U17625 ( .B1(n13968), .B2(DATAI_27_), .A(n14240), .ZN(n14241) );
  OAI21_X1 U17626 ( .B1(n14242), .B2(n14296), .A(n14241), .ZN(P1_U2877) );
  OAI22_X1 U17627 ( .A1(n14283), .A2(n20004), .B1(n14294), .B2(n13430), .ZN(
        n14243) );
  AOI21_X1 U17628 ( .B1(BUF1_REG_26__SCAN_IN), .B2(n14285), .A(n14243), .ZN(
        n14245) );
  NAND2_X1 U17629 ( .A1(n13968), .A2(DATAI_26_), .ZN(n14244) );
  OAI211_X1 U17630 ( .C1(n15675), .C2(n14296), .A(n14245), .B(n14244), .ZN(
        P1_U2878) );
  OAI22_X1 U17631 ( .A1(n14283), .A2(n20001), .B1(n14294), .B2(n13436), .ZN(
        n14246) );
  AOI21_X1 U17632 ( .B1(n14285), .B2(BUF1_REG_25__SCAN_IN), .A(n14246), .ZN(
        n14248) );
  NAND2_X1 U17633 ( .A1(n13968), .A2(DATAI_25_), .ZN(n14247) );
  OAI211_X1 U17634 ( .C1(n14338), .C2(n14296), .A(n14248), .B(n14247), .ZN(
        P1_U2879) );
  OAI22_X1 U17635 ( .A1(n14283), .A2(n19998), .B1(n14294), .B2(n13520), .ZN(
        n14249) );
  AOI21_X1 U17636 ( .B1(n14285), .B2(BUF1_REG_24__SCAN_IN), .A(n14249), .ZN(
        n14251) );
  NAND2_X1 U17637 ( .A1(n13968), .A2(DATAI_24_), .ZN(n14250) );
  OAI211_X1 U17638 ( .C1(n14252), .C2(n14296), .A(n14251), .B(n14250), .ZN(
        P1_U2880) );
  OAI22_X1 U17639 ( .A1(n14283), .A2(n20146), .B1(n14294), .B2(n20976), .ZN(
        n14254) );
  INV_X1 U17640 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n16332) );
  NOR2_X1 U17641 ( .A1(n14265), .A2(n16332), .ZN(n14253) );
  AOI211_X1 U17642 ( .C1(DATAI_23_), .C2(n13968), .A(n14254), .B(n14253), .ZN(
        n14255) );
  OAI21_X1 U17643 ( .B1(n14256), .B2(n14296), .A(n14255), .ZN(P1_U2881) );
  OAI22_X1 U17644 ( .A1(n14283), .A2(n20138), .B1(n14294), .B2(n13518), .ZN(
        n14257) );
  AOI21_X1 U17645 ( .B1(n14285), .B2(BUF1_REG_22__SCAN_IN), .A(n14257), .ZN(
        n14259) );
  NAND2_X1 U17646 ( .A1(n13968), .A2(DATAI_22_), .ZN(n14258) );
  OAI211_X1 U17647 ( .C1(n14361), .C2(n14296), .A(n14259), .B(n14258), .ZN(
        P1_U2882) );
  NOR2_X1 U17648 ( .A1(n14179), .A2(n14260), .ZN(n14261) );
  OR2_X1 U17649 ( .A1(n14034), .A2(n14261), .ZN(n15739) );
  INV_X1 U17650 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n16336) );
  AOI22_X1 U17651 ( .A1(n14263), .A2(n14262), .B1(P1_EAX_REG_21__SCAN_IN), 
        .B2(n14298), .ZN(n14264) );
  OAI21_X1 U17652 ( .B1(n16336), .B2(n14265), .A(n14264), .ZN(n14266) );
  AOI21_X1 U17653 ( .B1(n13968), .B2(DATAI_21_), .A(n14266), .ZN(n14267) );
  OAI21_X1 U17654 ( .B1(n15739), .B2(n14296), .A(n14267), .ZN(P1_U2883) );
  OAI22_X1 U17655 ( .A1(n14283), .A2(n20129), .B1(n14294), .B2(n13432), .ZN(
        n14268) );
  AOI21_X1 U17656 ( .B1(n14285), .B2(BUF1_REG_20__SCAN_IN), .A(n14268), .ZN(
        n14270) );
  NAND2_X1 U17657 ( .A1(n13968), .A2(DATAI_20_), .ZN(n14269) );
  OAI211_X1 U17658 ( .C1(n15701), .C2(n14296), .A(n14270), .B(n14269), .ZN(
        P1_U2884) );
  OAI22_X1 U17659 ( .A1(n14283), .A2(n20124), .B1(n14294), .B2(n14271), .ZN(
        n14272) );
  AOI21_X1 U17660 ( .B1(n14285), .B2(BUF1_REG_19__SCAN_IN), .A(n14272), .ZN(
        n14274) );
  NAND2_X1 U17661 ( .A1(n13968), .A2(DATAI_19_), .ZN(n14273) );
  OAI211_X1 U17662 ( .C1(n14275), .C2(n14296), .A(n14274), .B(n14273), .ZN(
        P1_U2885) );
  OAI22_X1 U17663 ( .A1(n14283), .A2(n20119), .B1(n14294), .B2(n14276), .ZN(
        n14277) );
  AOI21_X1 U17664 ( .B1(n14285), .B2(BUF1_REG_18__SCAN_IN), .A(n14277), .ZN(
        n14279) );
  NAND2_X1 U17665 ( .A1(n13968), .A2(DATAI_18_), .ZN(n14278) );
  OAI211_X1 U17666 ( .C1(n14389), .C2(n14296), .A(n14279), .B(n14278), .ZN(
        P1_U2886) );
  OAI22_X1 U17667 ( .A1(n14283), .A2(n20115), .B1(n14294), .B2(n13428), .ZN(
        n14280) );
  AOI21_X1 U17668 ( .B1(n14285), .B2(BUF1_REG_17__SCAN_IN), .A(n14280), .ZN(
        n14282) );
  NAND2_X1 U17669 ( .A1(n13968), .A2(DATAI_17_), .ZN(n14281) );
  OAI211_X1 U17670 ( .C1(n15754), .C2(n14296), .A(n14282), .B(n14281), .ZN(
        P1_U2887) );
  OAI22_X1 U17671 ( .A1(n14283), .A2(n20106), .B1(n14294), .B2(n13426), .ZN(
        n14284) );
  AOI21_X1 U17672 ( .B1(n14285), .B2(BUF1_REG_16__SCAN_IN), .A(n14284), .ZN(
        n14287) );
  NAND2_X1 U17673 ( .A1(n13968), .A2(DATAI_16_), .ZN(n14286) );
  OAI211_X1 U17674 ( .C1(n14288), .C2(n14296), .A(n14287), .B(n14286), .ZN(
        P1_U2888) );
  OAI222_X1 U17675 ( .A1(n14296), .A2(n14290), .B1(n14294), .B2(n13534), .C1(
        n14297), .C2(n14289), .ZN(P1_U2889) );
  INV_X1 U17676 ( .A(n14414), .ZN(n14292) );
  INV_X1 U17677 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n14291) );
  OAI222_X1 U17678 ( .A1(n14292), .A2(n14296), .B1(n14291), .B2(n14294), .C1(
        n14297), .C2(n20013), .ZN(P1_U2890) );
  INV_X1 U17679 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n14293) );
  OAI222_X1 U17680 ( .A1(n14296), .A2(n14430), .B1(n14297), .B2(n20010), .C1(
        n14293), .C2(n14294), .ZN(P1_U2891) );
  OAI222_X1 U17681 ( .A1(n15769), .A2(n14296), .B1(n14295), .B2(n14294), .C1(
        n14297), .C2(n20007), .ZN(P1_U2892) );
  INV_X1 U17682 ( .A(n15777), .ZN(n14302) );
  INV_X1 U17683 ( .A(n14297), .ZN(n14300) );
  AOI22_X1 U17684 ( .A1(n14300), .A2(n14299), .B1(P1_EAX_REG_11__SCAN_IN), 
        .B2(n14298), .ZN(n14301) );
  OAI21_X1 U17685 ( .B1(n14302), .B2(n14296), .A(n14301), .ZN(P1_U2893) );
  NOR2_X1 U17686 ( .A1(n14425), .A2(n14303), .ZN(n14304) );
  AOI211_X1 U17687 ( .C1(n20045), .C2(n14306), .A(n14305), .B(n14304), .ZN(
        n14309) );
  NAND2_X1 U17688 ( .A1(n14307), .A2(n20038), .ZN(n14308) );
  OAI211_X1 U17689 ( .C1(n14310), .C2(n19867), .A(n14309), .B(n14308), .ZN(
        P1_U2969) );
  AOI21_X1 U17690 ( .B1(n20043), .B2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n14311), .ZN(n14312) );
  OAI21_X1 U17691 ( .B1(n20041), .B2(n14313), .A(n14312), .ZN(n14314) );
  AOI21_X1 U17692 ( .B1(n14315), .B2(n20038), .A(n14314), .ZN(n14316) );
  OAI21_X1 U17693 ( .B1(n14317), .B2(n19867), .A(n14316), .ZN(P1_U2970) );
  OAI21_X1 U17694 ( .B1(n14332), .B2(n14455), .A(n14352), .ZN(n14319) );
  NAND2_X1 U17695 ( .A1(n14319), .A2(n14318), .ZN(n14326) );
  NOR2_X1 U17696 ( .A1(n14320), .A2(n14326), .ZN(n14321) );
  XNOR2_X1 U17697 ( .A(n14321), .B(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14454) );
  NAND2_X1 U17698 ( .A1(n11744), .A2(P1_REIP_REG_27__SCAN_IN), .ZN(n14448) );
  NAND2_X1 U17699 ( .A1(n20043), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14322) );
  OAI211_X1 U17700 ( .C1(n20041), .C2(n15667), .A(n14448), .B(n14322), .ZN(
        n14323) );
  AOI21_X1 U17701 ( .B1(n15664), .B2(n20038), .A(n14323), .ZN(n14324) );
  OAI21_X1 U17702 ( .B1(n14454), .B2(n19867), .A(n14324), .ZN(P1_U2972) );
  XNOR2_X1 U17703 ( .A(n14326), .B(n14325), .ZN(n14462) );
  AND2_X1 U17704 ( .A1(n11744), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n14457) );
  NOR2_X1 U17705 ( .A1(n14425), .A2(n15672), .ZN(n14327) );
  AOI211_X1 U17706 ( .C1(n20045), .C2(n15678), .A(n14457), .B(n14327), .ZN(
        n14330) );
  INV_X1 U17707 ( .A(n15675), .ZN(n14328) );
  NAND2_X1 U17708 ( .A1(n14328), .A2(n20038), .ZN(n14329) );
  OAI211_X1 U17709 ( .C1(n14462), .C2(n19867), .A(n14330), .B(n14329), .ZN(
        P1_U2973) );
  INV_X1 U17710 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n14476) );
  NAND3_X1 U17711 ( .A1(n14332), .A2(n14331), .A3(n14476), .ZN(n14335) );
  NAND2_X1 U17712 ( .A1(n14344), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14334) );
  MUX2_X1 U17713 ( .A(n14335), .B(n14334), .S(n14352), .Z(n14336) );
  XOR2_X1 U17714 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .B(n14336), .Z(
        n14469) );
  NAND2_X1 U17715 ( .A1(n11744), .A2(P1_REIP_REG_25__SCAN_IN), .ZN(n14464) );
  OAI21_X1 U17716 ( .B1(n14425), .B2(n14337), .A(n14464), .ZN(n14340) );
  NOR2_X1 U17717 ( .A1(n14338), .A2(n20094), .ZN(n14339) );
  AOI211_X1 U17718 ( .C1(n20045), .C2(n14341), .A(n14340), .B(n14339), .ZN(
        n14342) );
  OAI21_X1 U17719 ( .B1(n14469), .B2(n19867), .A(n14342), .ZN(P1_U2974) );
  NOR2_X1 U17720 ( .A1(n14344), .A2(n14354), .ZN(n14343) );
  MUX2_X1 U17721 ( .A(n14344), .B(n14343), .S(n11524), .Z(n14345) );
  XNOR2_X1 U17722 ( .A(n14345), .B(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14482) );
  NOR2_X1 U17723 ( .A1(n20081), .A2(n14029), .ZN(n14472) );
  NOR2_X1 U17724 ( .A1(n14425), .A2(n14346), .ZN(n14347) );
  AOI211_X1 U17725 ( .C1(n20045), .C2(n14348), .A(n14472), .B(n14347), .ZN(
        n14351) );
  NAND2_X1 U17726 ( .A1(n14349), .A2(n20038), .ZN(n14350) );
  OAI211_X1 U17727 ( .C1(n14482), .C2(n19867), .A(n14351), .B(n14350), .ZN(
        P1_U2975) );
  XNOR2_X1 U17728 ( .A(n14352), .B(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14353) );
  XNOR2_X1 U17729 ( .A(n14354), .B(n14353), .ZN(n14489) );
  NAND2_X1 U17730 ( .A1(n11744), .A2(P1_REIP_REG_23__SCAN_IN), .ZN(n14483) );
  NAND2_X1 U17731 ( .A1(n20043), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14355) );
  OAI211_X1 U17732 ( .C1(n20041), .C2(n15688), .A(n14483), .B(n14355), .ZN(
        n14356) );
  AOI21_X1 U17733 ( .B1(n15685), .B2(n20038), .A(n14356), .ZN(n14357) );
  OAI21_X1 U17734 ( .B1(n14489), .B2(n19867), .A(n14357), .ZN(P1_U2976) );
  NAND2_X1 U17735 ( .A1(n14359), .A2(n14358), .ZN(n14360) );
  XOR2_X1 U17736 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n14360), .Z(
        n15799) );
  INV_X1 U17737 ( .A(n14361), .ZN(n14366) );
  INV_X1 U17738 ( .A(n14362), .ZN(n14364) );
  AOI22_X1 U17739 ( .A1(n20043), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B1(
        n11744), .B2(P1_REIP_REG_22__SCAN_IN), .ZN(n14363) );
  OAI21_X1 U17740 ( .B1(n20041), .B2(n14364), .A(n14363), .ZN(n14365) );
  AOI21_X1 U17741 ( .B1(n14366), .B2(n20038), .A(n14365), .ZN(n14367) );
  OAI21_X1 U17742 ( .B1(n15799), .B2(n19867), .A(n14367), .ZN(P1_U2977) );
  NAND2_X1 U17743 ( .A1(n14352), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15745) );
  NOR2_X1 U17744 ( .A1(n14368), .A2(n15745), .ZN(n14378) );
  OAI21_X1 U17745 ( .B1(n14352), .B2(n14369), .A(n14368), .ZN(n15747) );
  NAND2_X1 U17746 ( .A1(n11524), .A2(n14370), .ZN(n15744) );
  NOR2_X1 U17747 ( .A1(n15747), .A2(n15744), .ZN(n15743) );
  MUX2_X1 U17748 ( .A(n14378), .B(n15743), .S(n14379), .Z(n14371) );
  XOR2_X1 U17749 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n14371), .Z(
        n14490) );
  NAND2_X1 U17750 ( .A1(n14490), .A2(n20046), .ZN(n14377) );
  INV_X1 U17751 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n14372) );
  NOR2_X1 U17752 ( .A1(n20081), .A2(n14372), .ZN(n14496) );
  NOR2_X1 U17753 ( .A1(n14425), .A2(n14373), .ZN(n14374) );
  AOI211_X1 U17754 ( .C1(n20045), .C2(n14375), .A(n14496), .B(n14374), .ZN(
        n14376) );
  OAI211_X1 U17755 ( .C1(n20094), .C2(n15739), .A(n14377), .B(n14376), .ZN(
        P1_U2978) );
  NOR2_X1 U17756 ( .A1(n15743), .A2(n14378), .ZN(n14380) );
  XNOR2_X1 U17757 ( .A(n14380), .B(n14379), .ZN(n14509) );
  NOR2_X1 U17758 ( .A1(n20081), .A2(n15698), .ZN(n14502) );
  NOR2_X1 U17759 ( .A1(n14425), .A2(n15706), .ZN(n14381) );
  AOI211_X1 U17760 ( .C1(n20045), .C2(n15703), .A(n14502), .B(n14381), .ZN(
        n14384) );
  INV_X1 U17761 ( .A(n15701), .ZN(n14382) );
  NAND2_X1 U17762 ( .A1(n14382), .A2(n20038), .ZN(n14383) );
  OAI211_X1 U17763 ( .C1(n14509), .C2(n19867), .A(n14384), .B(n14383), .ZN(
        P1_U2979) );
  OAI21_X1 U17764 ( .B1(n9811), .B2(n14385), .A(n14368), .ZN(n15817) );
  INV_X1 U17765 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n14387) );
  OAI22_X1 U17766 ( .A1(n14425), .A2(n14388), .B1(n20081), .B2(n14387), .ZN(
        n14391) );
  NOR2_X1 U17767 ( .A1(n14389), .A2(n20094), .ZN(n14390) );
  AOI211_X1 U17768 ( .C1(n20045), .C2(n14392), .A(n14391), .B(n14390), .ZN(
        n14393) );
  OAI21_X1 U17769 ( .B1(n19867), .B2(n15817), .A(n14393), .ZN(P1_U2981) );
  OAI21_X1 U17770 ( .B1(n14395), .B2(n14396), .A(n14406), .ZN(n14523) );
  INV_X1 U17771 ( .A(n14397), .ZN(n14398) );
  OAI21_X1 U17772 ( .B1(n14523), .B2(n14398), .A(n14524), .ZN(n14399) );
  XOR2_X1 U17773 ( .A(n14400), .B(n14399), .Z(n15825) );
  AOI22_X1 U17774 ( .A1(n20043), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B1(
        n11744), .B2(P1_REIP_REG_16__SCAN_IN), .ZN(n14401) );
  OAI21_X1 U17775 ( .B1(n20041), .B2(n14402), .A(n14401), .ZN(n14403) );
  AOI21_X1 U17776 ( .B1(n14404), .B2(n20038), .A(n14403), .ZN(n14405) );
  OAI21_X1 U17777 ( .B1(n15825), .B2(n19867), .A(n14405), .ZN(P1_U2983) );
  NAND2_X1 U17778 ( .A1(n14395), .A2(n14406), .ZN(n14407) );
  AOI22_X1 U17779 ( .A1(n14407), .A2(n9884), .B1(n11524), .B2(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n14410) );
  MUX2_X1 U17780 ( .A(n14408), .B(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .S(
        n14352), .Z(n14409) );
  XNOR2_X1 U17781 ( .A(n14410), .B(n14409), .ZN(n15838) );
  INV_X1 U17782 ( .A(n15838), .ZN(n14416) );
  AOI22_X1 U17783 ( .A1(n20043), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        n11744), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n14411) );
  OAI21_X1 U17784 ( .B1(n20041), .B2(n14412), .A(n14411), .ZN(n14413) );
  AOI21_X1 U17785 ( .B1(n14414), .B2(n20038), .A(n14413), .ZN(n14415) );
  OAI21_X1 U17786 ( .B1(n14416), .B2(n19867), .A(n14415), .ZN(P1_U2985) );
  INV_X1 U17787 ( .A(n14417), .ZN(n14418) );
  AOI21_X1 U17788 ( .B1(n14394), .B2(n14419), .A(n14418), .ZN(n15767) );
  AND2_X1 U17789 ( .A1(n14420), .A2(n14421), .ZN(n15766) );
  NAND2_X1 U17790 ( .A1(n15767), .A2(n15766), .ZN(n15765) );
  NAND2_X1 U17791 ( .A1(n15765), .A2(n14421), .ZN(n14423) );
  XNOR2_X1 U17792 ( .A(n14423), .B(n14422), .ZN(n15844) );
  NAND2_X1 U17793 ( .A1(n15844), .A2(n20046), .ZN(n14429) );
  INV_X1 U17794 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n14424) );
  OAI22_X1 U17795 ( .A1(n14425), .A2(n14424), .B1(n20081), .B2(n20722), .ZN(
        n14426) );
  AOI21_X1 U17796 ( .B1(n20045), .B2(n14427), .A(n14426), .ZN(n14428) );
  OAI211_X1 U17797 ( .C1(n20094), .C2(n14430), .A(n14429), .B(n14428), .ZN(
        P1_U2986) );
  MUX2_X1 U17798 ( .A(n14431), .B(n14395), .S(n14352), .Z(n14432) );
  XNOR2_X1 U17799 ( .A(n14432), .B(n11648), .ZN(n15875) );
  AOI22_X1 U17800 ( .A1(n20043), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        n11744), .B2(P1_REIP_REG_10__SCAN_IN), .ZN(n14433) );
  OAI21_X1 U17801 ( .B1(n20041), .B2(n14434), .A(n14433), .ZN(n14435) );
  AOI21_X1 U17802 ( .B1(n14436), .B2(n20038), .A(n14435), .ZN(n14437) );
  OAI21_X1 U17803 ( .B1(n15875), .B2(n19867), .A(n14437), .ZN(P1_U2989) );
  NAND2_X1 U17804 ( .A1(n14452), .A2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14444) );
  INV_X1 U17805 ( .A(n14449), .ZN(n14442) );
  NOR2_X1 U17806 ( .A1(n14439), .A2(n14438), .ZN(n14441) );
  AOI21_X1 U17807 ( .B1(n14442), .B2(n14441), .A(n14440), .ZN(n14443) );
  OAI211_X1 U17808 ( .C1(n20083), .C2(n15649), .A(n14444), .B(n14443), .ZN(
        n14445) );
  AOI21_X1 U17809 ( .B1(n14446), .B2(n20086), .A(n14445), .ZN(n14447) );
  INV_X1 U17810 ( .A(n14447), .ZN(P1_U3003) );
  OAI21_X1 U17811 ( .B1(n14449), .B2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n14448), .ZN(n14451) );
  NOR2_X1 U17812 ( .A1(n15662), .A2(n20083), .ZN(n14450) );
  AOI211_X1 U17813 ( .C1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n14452), .A(
        n14451), .B(n14450), .ZN(n14453) );
  OAI21_X1 U17814 ( .B1(n14454), .B2(n15923), .A(n14453), .ZN(P1_U3004) );
  NOR3_X1 U17815 ( .A1(n14470), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n14455), .ZN(n14456) );
  AOI211_X1 U17816 ( .C1(n20063), .C2(n15673), .A(n14457), .B(n14456), .ZN(
        n14461) );
  OR3_X1 U17817 ( .A1(n14470), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(
        n14458), .ZN(n14463) );
  INV_X1 U17818 ( .A(n14463), .ZN(n14459) );
  OAI21_X1 U17819 ( .B1(n14467), .B2(n14459), .A(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14460) );
  OAI211_X1 U17820 ( .C1(n14462), .C2(n15923), .A(n14461), .B(n14460), .ZN(
        P1_U3005) );
  OAI211_X1 U17821 ( .C1(n14465), .C2(n20083), .A(n14464), .B(n14463), .ZN(
        n14466) );
  AOI21_X1 U17822 ( .B1(n14467), .B2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n14466), .ZN(n14468) );
  OAI21_X1 U17823 ( .B1(n14469), .B2(n15923), .A(n14468), .ZN(P1_U3006) );
  NOR3_X1 U17824 ( .A1(n14470), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        n14476), .ZN(n14471) );
  AOI211_X1 U17825 ( .C1(n20063), .C2(n14473), .A(n14472), .B(n14471), .ZN(
        n14481) );
  INV_X1 U17826 ( .A(n14474), .ZN(n14487) );
  INV_X1 U17827 ( .A(n20071), .ZN(n15854) );
  INV_X1 U17828 ( .A(n14475), .ZN(n14477) );
  NAND4_X1 U17829 ( .A1(n14478), .A2(n14477), .A3(n15800), .A4(n14476), .ZN(
        n14484) );
  OAI22_X1 U17830 ( .A1(n15854), .A2(n14484), .B1(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n20080), .ZN(n14479) );
  OAI21_X1 U17831 ( .B1(n14487), .B2(n14479), .A(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14480) );
  OAI211_X1 U17832 ( .C1(n14482), .C2(n15923), .A(n14481), .B(n14480), .ZN(
        P1_U3007) );
  NOR2_X1 U17833 ( .A1(n15683), .A2(n20083), .ZN(n14486) );
  OAI21_X1 U17834 ( .B1(n15841), .B2(n14484), .A(n14483), .ZN(n14485) );
  AOI211_X1 U17835 ( .C1(n14487), .C2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n14486), .B(n14485), .ZN(n14488) );
  OAI21_X1 U17836 ( .B1(n14489), .B2(n15923), .A(n14488), .ZN(P1_U3008) );
  INV_X1 U17837 ( .A(n15798), .ZN(n14499) );
  INV_X1 U17838 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n20949) );
  NAND2_X1 U17839 ( .A1(n14490), .A2(n20086), .ZN(n14498) );
  NAND2_X1 U17840 ( .A1(n14492), .A2(n14491), .ZN(n14493) );
  NAND2_X1 U17841 ( .A1(n14494), .A2(n14493), .ZN(n15738) );
  NOR2_X1 U17842 ( .A1(n15738), .A2(n20083), .ZN(n14495) );
  AOI211_X1 U17843 ( .C1(n15803), .C2(n20949), .A(n14496), .B(n14495), .ZN(
        n14497) );
  OAI211_X1 U17844 ( .C1(n14499), .C2(n20949), .A(n14498), .B(n14497), .ZN(
        P1_U3010) );
  NOR2_X1 U17845 ( .A1(n14500), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n14501) );
  AOI211_X1 U17846 ( .C1(n20063), .C2(n14503), .A(n14502), .B(n14501), .ZN(
        n14508) );
  AOI21_X1 U17847 ( .B1(n14505), .B2(n14504), .A(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n14506) );
  OAI21_X1 U17848 ( .B1(n15808), .B2(n14506), .A(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14507) );
  OAI211_X1 U17849 ( .C1(n14509), .C2(n15923), .A(n14508), .B(n14507), .ZN(
        P1_U3011) );
  AOI21_X1 U17850 ( .B1(n14395), .B2(n14511), .A(n14510), .ZN(n14513) );
  NOR2_X1 U17851 ( .A1(n14513), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14512) );
  MUX2_X1 U17852 ( .A(n14513), .B(n14512), .S(n11524), .Z(n14514) );
  XNOR2_X1 U17853 ( .A(n14514), .B(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15759) );
  AOI22_X1 U17854 ( .A1(n14515), .A2(n20063), .B1(n11744), .B2(
        P1_REIP_REG_17__SCAN_IN), .ZN(n14522) );
  NAND2_X1 U17855 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n14516) );
  INV_X1 U17856 ( .A(n15816), .ZN(n15823) );
  OAI21_X1 U17857 ( .B1(n14516), .B2(n15823), .A(n10205), .ZN(n14520) );
  INV_X1 U17858 ( .A(n15814), .ZN(n14518) );
  OAI21_X1 U17859 ( .B1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n14519), .A(
        n15848), .ZN(n15828) );
  INV_X1 U17860 ( .A(n15828), .ZN(n14517) );
  OAI21_X1 U17861 ( .B1(n14519), .B2(n14518), .A(n14517), .ZN(n15818) );
  NAND2_X1 U17862 ( .A1(n14520), .A2(n15818), .ZN(n14521) );
  OAI211_X1 U17863 ( .C1(n15759), .C2(n15923), .A(n14522), .B(n14521), .ZN(
        P1_U3014) );
  NOR2_X1 U17864 ( .A1(n14523), .A2(n9879), .ZN(n14527) );
  NAND2_X1 U17865 ( .A1(n14525), .A2(n14524), .ZN(n14526) );
  XNOR2_X1 U17866 ( .A(n14527), .B(n14526), .ZN(n15764) );
  NOR2_X1 U17867 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n15823), .ZN(
        n15829) );
  AOI21_X1 U17868 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n15828), .A(
        n15829), .ZN(n14528) );
  OAI21_X1 U17869 ( .B1(n20081), .B2(n20724), .A(n14528), .ZN(n14529) );
  AOI21_X1 U17870 ( .B1(n14530), .B2(n20063), .A(n14529), .ZN(n14531) );
  OAI21_X1 U17871 ( .B1(n15764), .B2(n15923), .A(n14531), .ZN(P1_U3016) );
  OR2_X1 U17872 ( .A1(n14532), .A2(n20075), .ZN(n14542) );
  AOI22_X1 U17873 ( .A1(n20063), .A2(n14533), .B1(n11744), .B2(
        P1_REIP_REG_1__SCAN_IN), .ZN(n14541) );
  OR2_X1 U17874 ( .A1(n14534), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n14535) );
  AND2_X1 U17875 ( .A1(n14536), .A2(n14535), .ZN(n20047) );
  NAND2_X1 U17876 ( .A1(n20047), .A2(n20086), .ZN(n14540) );
  NOR2_X1 U17877 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n14537), .ZN(
        n14538) );
  NAND2_X1 U17878 ( .A1(n15897), .A2(n14538), .ZN(n14539) );
  NAND4_X1 U17879 ( .A1(n14542), .A2(n14541), .A3(n14540), .A4(n14539), .ZN(
        P1_U3030) );
  INV_X1 U17880 ( .A(n14544), .ZN(n20365) );
  NAND2_X1 U17881 ( .A1(n20543), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n20628) );
  XNOR2_X1 U17882 ( .A(n20365), .B(n20628), .ZN(n14546) );
  OAI22_X1 U17883 ( .A1(n14546), .A2(n20632), .B1(n13438), .B2(n14545), .ZN(
        n14547) );
  MUX2_X1 U17884 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n14547), .S(
        n20771), .Z(P1_U3476) );
  NOR2_X1 U17885 ( .A1(n15585), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n14550) );
  NOR3_X1 U17886 ( .A1(n14548), .A2(n13594), .A3(n13446), .ZN(n14549) );
  AOI211_X1 U17887 ( .C1(n20577), .C2(n14551), .A(n14550), .B(n14549), .ZN(
        n15586) );
  INV_X1 U17888 ( .A(n14552), .ZN(n14557) );
  NOR3_X1 U17889 ( .A1(n13594), .A2(n13446), .A3(n15613), .ZN(n14553) );
  AOI21_X1 U17890 ( .B1(n14555), .B2(n14554), .A(n14553), .ZN(n14556) );
  OAI21_X1 U17891 ( .B1(n15586), .B2(n14557), .A(n14556), .ZN(n14559) );
  MUX2_X1 U17892 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n14559), .S(
        n14558), .Z(P1_U3473) );
  INV_X1 U17893 ( .A(n14676), .ZN(n14560) );
  OAI21_X1 U17894 ( .B1(n14691), .B2(n14561), .A(n14560), .ZN(n15163) );
  OAI211_X1 U17895 ( .C1(n14563), .C2(n14966), .A(n18999), .B(n14562), .ZN(
        n14573) );
  OR2_X1 U17896 ( .A1(n14906), .A2(n14565), .ZN(n14897) );
  INV_X1 U17897 ( .A(n14897), .ZN(n14571) );
  AOI22_X1 U17898 ( .A1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n18964), .B1(
        P2_REIP_REG_28__SCAN_IN), .B2(n18989), .ZN(n14566) );
  INV_X1 U17899 ( .A(n14566), .ZN(n14570) );
  AND2_X1 U17900 ( .A1(n14780), .A2(n14567), .ZN(n14568) );
  NOR2_X1 U17901 ( .A1(n14762), .A2(n14568), .ZN(n14774) );
  OAI22_X1 U17902 ( .A1(n15159), .A2(n18982), .B1(n12133), .B2(n18960), .ZN(
        n14569) );
  AOI211_X1 U17903 ( .C1(n14571), .C2(n18950), .A(n14570), .B(n14569), .ZN(
        n14572) );
  OAI211_X1 U17904 ( .C1(n18981), .C2(n15163), .A(n14573), .B(n14572), .ZN(
        P2_U2827) );
  INV_X1 U17905 ( .A(n14574), .ZN(n14588) );
  XOR2_X1 U17906 ( .A(n16069), .B(n18895), .Z(n14576) );
  NAND2_X1 U17907 ( .A1(n14576), .A2(n18999), .ZN(n14587) );
  INV_X1 U17908 ( .A(n14577), .ZN(n14579) );
  AOI21_X1 U17909 ( .B1(n14579), .B2(n14578), .A(n9876), .ZN(n19042) );
  AOI22_X1 U17910 ( .A1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n18964), .B1(
        P2_REIP_REG_14__SCAN_IN), .B2(n18989), .ZN(n14580) );
  OAI211_X1 U17911 ( .C1(n18960), .C2(n14581), .A(n14580), .B(n9889), .ZN(
        n14585) );
  INV_X1 U17912 ( .A(n13763), .ZN(n14583) );
  OAI21_X1 U17913 ( .B1(n14583), .B2(n10075), .A(n14748), .ZN(n19014) );
  NOR2_X1 U17914 ( .A1(n19014), .A2(n18981), .ZN(n14584) );
  AOI211_X1 U17915 ( .C1(n18991), .C2(n19042), .A(n14585), .B(n14584), .ZN(
        n14586) );
  OAI211_X1 U17916 ( .C1(n18994), .C2(n14588), .A(n14587), .B(n14586), .ZN(
        P2_U2841) );
  AOI21_X1 U17917 ( .B1(n13616), .B2(n14589), .A(n13726), .ZN(n16164) );
  INV_X1 U17918 ( .A(n16164), .ZN(n19050) );
  NAND2_X1 U17919 ( .A1(n18873), .A2(n18916), .ZN(n14590) );
  XNOR2_X1 U17920 ( .A(n16079), .B(n14590), .ZN(n14591) );
  NAND2_X1 U17921 ( .A1(n14591), .A2(n18999), .ZN(n14599) );
  OR2_X1 U17922 ( .A1(n13717), .A2(n14592), .ZN(n14593) );
  NAND2_X1 U17923 ( .A1(n13764), .A2(n14593), .ZN(n19023) );
  NOR2_X1 U17924 ( .A1(n19023), .A2(n18981), .ZN(n14596) );
  INV_X1 U17925 ( .A(P2_EBX_REG_12__SCAN_IN), .ZN(n19019) );
  AOI22_X1 U17926 ( .A1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n18964), .B1(
        P2_REIP_REG_12__SCAN_IN), .B2(n18989), .ZN(n14594) );
  OAI211_X1 U17927 ( .C1(n18960), .C2(n19019), .A(n14594), .B(n9889), .ZN(
        n14595) );
  AOI211_X1 U17928 ( .C1(n14597), .C2(n18950), .A(n14596), .B(n14595), .ZN(
        n14598) );
  OAI211_X1 U17929 ( .C1(n18982), .C2(n19050), .A(n14599), .B(n14598), .ZN(
        P2_U2843) );
  NAND2_X1 U17930 ( .A1(n12116), .A2(n14600), .ZN(n14601) );
  XNOR2_X1 U17931 ( .A(n16099), .B(n14601), .ZN(n14602) );
  NAND2_X1 U17932 ( .A1(n14602), .A2(n18999), .ZN(n14610) );
  OAI21_X1 U17933 ( .B1(n14604), .B2(n14603), .A(n13681), .ZN(n19036) );
  INV_X1 U17934 ( .A(n19036), .ZN(n16184) );
  INV_X1 U17935 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n14607) );
  AOI22_X1 U17936 ( .A1(P2_EBX_REG_8__SCAN_IN), .A2(n18990), .B1(n18991), .B2(
        n16180), .ZN(n14606) );
  AOI21_X1 U17937 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n18964), .A(
        n16186), .ZN(n14605) );
  OAI211_X1 U17938 ( .C1(n14607), .C2(n18973), .A(n14606), .B(n14605), .ZN(
        n14608) );
  AOI21_X1 U17939 ( .B1(n16184), .B2(n18997), .A(n14608), .ZN(n14609) );
  OAI211_X1 U17940 ( .C1(n18994), .C2(n14611), .A(n14610), .B(n14609), .ZN(
        P2_U2847) );
  NAND2_X1 U17941 ( .A1(n14612), .A2(n13476), .ZN(n14614) );
  NAND2_X1 U17942 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n12305), .ZN(
        n14613) );
  NAND2_X1 U17943 ( .A1(n14614), .A2(n14613), .ZN(n14618) );
  INV_X1 U17944 ( .A(n14615), .ZN(n14617) );
  OR3_X1 U17945 ( .A1(n14618), .A2(n14617), .A3(n14616), .ZN(n14619) );
  NAND2_X1 U17946 ( .A1(n13486), .A2(n14619), .ZN(n19065) );
  AND2_X1 U17947 ( .A1(n18873), .A2(n14620), .ZN(n14622) );
  AOI21_X1 U17948 ( .B1(n14623), .B2(n14622), .A(n19705), .ZN(n14621) );
  OAI21_X1 U17949 ( .B1(n14623), .B2(n14622), .A(n14621), .ZN(n14633) );
  INV_X1 U17950 ( .A(n19041), .ZN(n14631) );
  OAI21_X1 U17951 ( .B1(n18960), .B2(n14624), .A(n9889), .ZN(n14625) );
  AOI21_X1 U17952 ( .B1(n18991), .B2(n19063), .A(n14625), .ZN(n14626) );
  OAI21_X1 U17953 ( .B1(n14627), .B2(n18994), .A(n14626), .ZN(n14630) );
  INV_X1 U17954 ( .A(n19002), .ZN(n18987) );
  OAI22_X1 U17955 ( .A1(n14628), .A2(n18987), .B1(n19729), .B2(n18973), .ZN(
        n14629) );
  AOI211_X1 U17956 ( .C1(n14631), .C2(n18997), .A(n14630), .B(n14629), .ZN(
        n14632) );
  OAI211_X1 U17957 ( .C1(n19065), .C2(n14652), .A(n14633), .B(n14632), .ZN(
        P2_U2851) );
  NOR2_X1 U17958 ( .A1(n14665), .A2(n14634), .ZN(n14636) );
  XNOR2_X1 U17959 ( .A(n14636), .B(n14635), .ZN(n14648) );
  NOR2_X1 U17960 ( .A1(n19788), .A2(n14652), .ZN(n14647) );
  OR2_X1 U17961 ( .A1(n14638), .A2(n14637), .ZN(n14639) );
  NAND2_X1 U17962 ( .A1(n14639), .A2(n13860), .ZN(n21134) );
  INV_X1 U17963 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n19728) );
  OAI22_X1 U17964 ( .A1(n11017), .A2(n18960), .B1(n19728), .B2(n18973), .ZN(
        n14643) );
  OAI22_X1 U17965 ( .A1(n14641), .A2(n18994), .B1(n14640), .B2(n18987), .ZN(
        n14642) );
  OR2_X1 U17966 ( .A1(n14643), .A2(n14642), .ZN(n14644) );
  AOI21_X1 U17967 ( .B1(n12304), .B2(n18997), .A(n14644), .ZN(n14645) );
  OAI21_X1 U17968 ( .B1(n21134), .B2(n18982), .A(n14645), .ZN(n14646) );
  AOI211_X1 U17969 ( .C1(n14648), .C2(n18999), .A(n14647), .B(n14646), .ZN(
        n14649) );
  INV_X1 U17970 ( .A(n14649), .ZN(P2_U2852) );
  NAND2_X1 U17971 ( .A1(n12116), .A2(n14663), .ZN(n14650) );
  XNOR2_X1 U17972 ( .A(n14651), .B(n14650), .ZN(n14661) );
  NOR2_X1 U17973 ( .A1(n19147), .A2(n14652), .ZN(n14660) );
  OAI22_X1 U17974 ( .A1(n14653), .A2(n18960), .B1(n10566), .B2(n18973), .ZN(
        n14654) );
  AOI21_X1 U17975 ( .B1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n18964), .A(
        n14654), .ZN(n14655) );
  OAI21_X1 U17976 ( .B1(n14656), .B2(n18994), .A(n14655), .ZN(n14657) );
  AOI21_X1 U17977 ( .B1(n9829), .B2(n18997), .A(n14657), .ZN(n14658) );
  OAI21_X1 U17978 ( .B1(n19797), .B2(n18982), .A(n14658), .ZN(n14659) );
  AOI211_X1 U17979 ( .C1(n14661), .C2(n18999), .A(n14660), .B(n14659), .ZN(
        n14662) );
  INV_X1 U17980 ( .A(n14662), .ZN(P2_U2853) );
  OAI211_X1 U17981 ( .C1(n15368), .C2(n14664), .A(n12116), .B(n14663), .ZN(
        n15388) );
  NAND2_X1 U17982 ( .A1(n18999), .A2(n14665), .ZN(n18922) );
  AOI22_X1 U17983 ( .A1(P2_EBX_REG_1__SCAN_IN), .A2(n18990), .B1(
        P2_REIP_REG_1__SCAN_IN), .B2(n18989), .ZN(n14666) );
  OAI21_X1 U17984 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n18922), .A(
        n14666), .ZN(n14667) );
  AOI21_X1 U17985 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n18964), .A(
        n14667), .ZN(n14668) );
  OAI21_X1 U17986 ( .B1(n14669), .B2(n18994), .A(n14668), .ZN(n14670) );
  AOI21_X1 U17987 ( .B1(n19811), .B2(n18991), .A(n14670), .ZN(n14671) );
  OAI21_X1 U17988 ( .B1(n14672), .B2(n18981), .A(n14671), .ZN(n14673) );
  AOI21_X1 U17989 ( .B1(n19807), .B2(n18998), .A(n14673), .ZN(n14674) );
  OAI21_X1 U17990 ( .B1(n15388), .B2(n19705), .A(n14674), .ZN(P2_U2854) );
  OR2_X1 U17991 ( .A1(n14676), .A2(n14675), .ZN(n14677) );
  NAND2_X1 U17992 ( .A1(n14678), .A2(n14677), .ZN(n14948) );
  INV_X1 U17993 ( .A(n14679), .ZN(n14759) );
  NAND2_X1 U17994 ( .A1(n9803), .A2(n14680), .ZN(n14758) );
  NAND3_X1 U17995 ( .A1(n14759), .A2(n19038), .A3(n14758), .ZN(n14682) );
  NAND2_X1 U17996 ( .A1(n19037), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n14681) );
  OAI211_X1 U17997 ( .C1(n19037), .C2(n14948), .A(n14682), .B(n14681), .ZN(
        P2_U2858) );
  NAND2_X1 U17998 ( .A1(n12570), .A2(n14683), .ZN(n14685) );
  XNOR2_X1 U17999 ( .A(n14685), .B(n14684), .ZN(n14777) );
  NOR2_X1 U18000 ( .A1(n15163), .A2(n19037), .ZN(n14686) );
  AOI21_X1 U18001 ( .B1(P2_EBX_REG_28__SCAN_IN), .B2(n19037), .A(n14686), .ZN(
        n14687) );
  OAI21_X1 U18002 ( .B1(n14777), .B2(n19031), .A(n14687), .ZN(P2_U2859) );
  NOR2_X1 U18003 ( .A1(n14688), .A2(n14689), .ZN(n14690) );
  OR2_X1 U18004 ( .A1(n14691), .A2(n14690), .ZN(n15168) );
  NAND2_X1 U18005 ( .A1(n14778), .A2(n19038), .ZN(n14696) );
  NAND2_X1 U18006 ( .A1(n19037), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n14695) );
  OAI211_X1 U18007 ( .C1(n15168), .C2(n19037), .A(n14696), .B(n14695), .ZN(
        P2_U2860) );
  AOI21_X1 U18008 ( .B1(n14697), .B2(n14699), .A(n14698), .ZN(n14700) );
  INV_X1 U18009 ( .A(n14700), .ZN(n14795) );
  AND2_X1 U18010 ( .A1(n14711), .A2(n14701), .ZN(n14702) );
  OR2_X1 U18011 ( .A1(n14702), .A2(n14688), .ZN(n15977) );
  NOR2_X1 U18012 ( .A1(n15977), .A2(n19037), .ZN(n14703) );
  AOI21_X1 U18013 ( .B1(P2_EBX_REG_26__SCAN_IN), .B2(n19037), .A(n14703), .ZN(
        n14704) );
  OAI21_X1 U18014 ( .B1(n14795), .B2(n19031), .A(n14704), .ZN(P2_U2861) );
  OAI21_X1 U18015 ( .B1(n14705), .B2(n14707), .A(n14706), .ZN(n14805) );
  NAND2_X1 U18016 ( .A1(n14708), .A2(n14709), .ZN(n14710) );
  NAND2_X1 U18017 ( .A1(n14711), .A2(n14710), .ZN(n15988) );
  MUX2_X1 U18018 ( .A(n15988), .B(n14888), .S(n19037), .Z(n14712) );
  OAI21_X1 U18019 ( .B1(n14805), .B2(n19031), .A(n14712), .ZN(P2_U2862) );
  INV_X1 U18020 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n14874) );
  NAND2_X1 U18021 ( .A1(n14713), .A2(n14714), .ZN(n14806) );
  NAND3_X1 U18022 ( .A1(n14807), .A2(n19038), .A3(n14806), .ZN(n14718) );
  OR2_X1 U18023 ( .A1(n14723), .A2(n14715), .ZN(n14716) );
  NAND2_X1 U18024 ( .A1(n14708), .A2(n14716), .ZN(n15209) );
  INV_X1 U18025 ( .A(n15209), .ZN(n15999) );
  NAND2_X1 U18026 ( .A1(n15999), .A2(n19020), .ZN(n14717) );
  OAI211_X1 U18027 ( .C1(n19020), .C2(n14874), .A(n14718), .B(n14717), .ZN(
        P2_U2863) );
  AOI21_X1 U18028 ( .B1(n14719), .B2(n14721), .A(n14720), .ZN(n14722) );
  INV_X1 U18029 ( .A(n14722), .ZN(n14823) );
  INV_X1 U18030 ( .A(n14723), .ZN(n14726) );
  NAND2_X1 U18031 ( .A1(n15238), .A2(n14724), .ZN(n14725) );
  NAND2_X1 U18032 ( .A1(n14726), .A2(n14725), .ZN(n16010) );
  NOR2_X1 U18033 ( .A1(n16010), .A2(n19037), .ZN(n14727) );
  AOI21_X1 U18034 ( .B1(P2_EBX_REG_23__SCAN_IN), .B2(n19037), .A(n14727), .ZN(
        n14728) );
  OAI21_X1 U18035 ( .B1(n14823), .B2(n19031), .A(n14728), .ZN(P2_U2864) );
  OAI21_X1 U18036 ( .B1(n14729), .B2(n14730), .A(n9878), .ZN(n14829) );
  MUX2_X1 U18037 ( .A(n18814), .B(n14731), .S(n19037), .Z(n14732) );
  OAI21_X1 U18038 ( .B1(n14829), .B2(n19031), .A(n14732), .ZN(P2_U2866) );
  NOR2_X1 U18039 ( .A1(n14734), .A2(n16031), .ZN(n16030) );
  INV_X1 U18040 ( .A(n14735), .ZN(n16026) );
  OAI21_X1 U18041 ( .B1(n16030), .B2(n14736), .A(n16026), .ZN(n14838) );
  NOR2_X1 U18042 ( .A1(n14737), .A2(n14738), .ZN(n14739) );
  OR2_X1 U18043 ( .A1(n15018), .A2(n14739), .ZN(n16131) );
  NOR2_X1 U18044 ( .A1(n16131), .A2(n19037), .ZN(n14740) );
  AOI21_X1 U18045 ( .B1(P2_EBX_REG_19__SCAN_IN), .B2(n19037), .A(n14740), .ZN(
        n14741) );
  OAI21_X1 U18046 ( .B1(n14838), .B2(n19031), .A(n14741), .ZN(P2_U2868) );
  OAI21_X1 U18047 ( .B1(n13909), .B2(n14742), .A(n14734), .ZN(n14845) );
  NAND2_X1 U18048 ( .A1(n19037), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n14744) );
  NAND2_X1 U18049 ( .A1(n18863), .A2(n19020), .ZN(n14743) );
  OAI211_X1 U18050 ( .C1(n14845), .C2(n19031), .A(n14744), .B(n14743), .ZN(
        P2_U2870) );
  XNOR2_X1 U18051 ( .A(n14745), .B(n14746), .ZN(n14752) );
  AND2_X1 U18052 ( .A1(n14748), .A2(n14747), .ZN(n14749) );
  OR2_X1 U18053 ( .A1(n14749), .A2(n15049), .ZN(n18889) );
  INV_X1 U18054 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n14750) );
  MUX2_X1 U18055 ( .A(n18889), .B(n14750), .S(n19037), .Z(n14751) );
  OAI21_X1 U18056 ( .B1(n14752), .B2(n19031), .A(n14751), .ZN(P2_U2872) );
  INV_X1 U18057 ( .A(n16049), .ZN(n14757) );
  AOI222_X1 U18058 ( .A1(n12156), .A2(P2_REIP_REG_31__SCAN_IN), .B1(n12151), 
        .B2(P2_EAX_REG_31__SCAN_IN), .C1(n10820), .C2(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14753) );
  XNOR2_X1 U18059 ( .A(n14754), .B(n14753), .ZN(n15116) );
  AOI22_X1 U18060 ( .A1(n15116), .A2(n19084), .B1(P2_EAX_REG_31__SCAN_IN), 
        .B2(n19083), .ZN(n14756) );
  NAND2_X1 U18061 ( .A1(n16048), .A2(BUF2_REG_31__SCAN_IN), .ZN(n14755) );
  OAI211_X1 U18062 ( .C1(n16318), .C2(n14757), .A(n14756), .B(n14755), .ZN(
        P2_U2888) );
  NAND3_X1 U18063 ( .A1(n14759), .A2(n19086), .A3(n14758), .ZN(n14768) );
  OAI21_X1 U18064 ( .B1(n14762), .B2(n14761), .A(n14760), .ZN(n15142) );
  OAI22_X1 U18065 ( .A1(n16040), .A2(n15142), .B1(n19044), .B2(n14763), .ZN(
        n14764) );
  AOI21_X1 U18066 ( .B1(n16047), .B2(n14765), .A(n14764), .ZN(n14767) );
  AOI22_X1 U18067 ( .A1(n16048), .A2(BUF2_REG_29__SCAN_IN), .B1(n16049), .B2(
        BUF1_REG_29__SCAN_IN), .ZN(n14766) );
  NAND3_X1 U18068 ( .A1(n14768), .A2(n14767), .A3(n14766), .ZN(P2_U2890) );
  OR2_X1 U18069 ( .A1(n14769), .A2(n21043), .ZN(n14771) );
  NAND2_X1 U18070 ( .A1(n14769), .A2(BUF2_REG_12__SCAN_IN), .ZN(n14770) );
  AND2_X1 U18071 ( .A1(n14771), .A2(n14770), .ZN(n19048) );
  INV_X1 U18072 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n14772) );
  OAI22_X1 U18073 ( .A1(n19048), .A2(n14841), .B1(n19044), .B2(n14772), .ZN(
        n14773) );
  AOI21_X1 U18074 ( .B1(n19084), .B2(n14774), .A(n14773), .ZN(n14776) );
  AOI22_X1 U18075 ( .A1(n16048), .A2(BUF2_REG_28__SCAN_IN), .B1(n16049), .B2(
        BUF1_REG_28__SCAN_IN), .ZN(n14775) );
  OAI211_X1 U18076 ( .C1(n14777), .C2(n19079), .A(n14776), .B(n14775), .ZN(
        P2_U2891) );
  INV_X1 U18077 ( .A(n14778), .ZN(n14788) );
  INV_X1 U18078 ( .A(n14791), .ZN(n14782) );
  INV_X1 U18079 ( .A(n14779), .ZN(n14781) );
  OAI21_X1 U18080 ( .B1(n14782), .B2(n14781), .A(n14780), .ZN(n15974) );
  OAI22_X1 U18081 ( .A1(n16040), .A2(n15974), .B1(n19044), .B2(n14783), .ZN(
        n14784) );
  AOI21_X1 U18082 ( .B1(n16047), .B2(n14785), .A(n14784), .ZN(n14787) );
  AOI22_X1 U18083 ( .A1(n16048), .A2(BUF2_REG_27__SCAN_IN), .B1(n16049), .B2(
        BUF1_REG_27__SCAN_IN), .ZN(n14786) );
  OAI211_X1 U18084 ( .C1(n14788), .C2(n19079), .A(n14787), .B(n14786), .ZN(
        P2_U2892) );
  NAND2_X1 U18085 ( .A1(n14799), .A2(n14789), .ZN(n14790) );
  NAND2_X1 U18086 ( .A1(n14791), .A2(n14790), .ZN(n15976) );
  OAI22_X1 U18087 ( .A1(n16040), .A2(n15976), .B1(n19044), .B2(n13398), .ZN(
        n14792) );
  AOI21_X1 U18088 ( .B1(n16047), .B2(n19051), .A(n14792), .ZN(n14794) );
  AOI22_X1 U18089 ( .A1(n16048), .A2(BUF2_REG_26__SCAN_IN), .B1(n16049), .B2(
        BUF1_REG_26__SCAN_IN), .ZN(n14793) );
  OAI211_X1 U18090 ( .C1(n14795), .C2(n19079), .A(n14794), .B(n14793), .ZN(
        P2_U2893) );
  OR2_X1 U18091 ( .A1(n14796), .A2(n14797), .ZN(n14798) );
  AND2_X1 U18092 ( .A1(n14799), .A2(n14798), .ZN(n15194) );
  INV_X1 U18093 ( .A(n15194), .ZN(n15987) );
  OAI22_X1 U18094 ( .A1(n16040), .A2(n15987), .B1(n19044), .B2(n14800), .ZN(
        n14801) );
  AOI21_X1 U18095 ( .B1(n16047), .B2(n14802), .A(n14801), .ZN(n14804) );
  AOI22_X1 U18096 ( .A1(n16048), .A2(BUF2_REG_25__SCAN_IN), .B1(n16049), .B2(
        BUF1_REG_25__SCAN_IN), .ZN(n14803) );
  OAI211_X1 U18097 ( .C1(n14805), .C2(n19079), .A(n14804), .B(n14803), .ZN(
        P2_U2894) );
  NAND3_X1 U18098 ( .A1(n14807), .A2(n19086), .A3(n14806), .ZN(n14815) );
  AND2_X1 U18099 ( .A1(n14817), .A2(n14808), .ZN(n14809) );
  NOR2_X1 U18100 ( .A1(n14796), .A2(n14809), .ZN(n15998) );
  OAI22_X1 U18101 ( .A1(n14811), .A2(n14841), .B1(n19044), .B2(n14810), .ZN(
        n14812) );
  AOI21_X1 U18102 ( .B1(n19084), .B2(n15998), .A(n14812), .ZN(n14814) );
  AOI22_X1 U18103 ( .A1(n16048), .A2(BUF2_REG_24__SCAN_IN), .B1(n16049), .B2(
        BUF1_REG_24__SCAN_IN), .ZN(n14813) );
  NAND3_X1 U18104 ( .A1(n14815), .A2(n14814), .A3(n14813), .ZN(P2_U2895) );
  OAI21_X1 U18105 ( .B1(n14818), .B2(n14816), .A(n14817), .ZN(n16018) );
  INV_X1 U18106 ( .A(n16018), .ZN(n15219) );
  OAI22_X1 U18107 ( .A1(n19181), .A2(n14841), .B1(n19044), .B2(n14819), .ZN(
        n14820) );
  AOI21_X1 U18108 ( .B1(n19084), .B2(n15219), .A(n14820), .ZN(n14822) );
  AOI22_X1 U18109 ( .A1(n16048), .A2(BUF2_REG_23__SCAN_IN), .B1(n16049), .B2(
        BUF1_REG_23__SCAN_IN), .ZN(n14821) );
  OAI211_X1 U18110 ( .C1(n14823), .C2(n19079), .A(n14822), .B(n14821), .ZN(
        P2_U2896) );
  NOR2_X1 U18111 ( .A1(n16040), .A2(n18813), .ZN(n14826) );
  OAI22_X1 U18112 ( .A1(n19171), .A2(n14841), .B1(n19044), .B2(n14824), .ZN(
        n14825) );
  NOR2_X1 U18113 ( .A1(n14826), .A2(n14825), .ZN(n14828) );
  AOI22_X1 U18114 ( .A1(n16048), .A2(BUF2_REG_21__SCAN_IN), .B1(n16049), .B2(
        BUF1_REG_21__SCAN_IN), .ZN(n14827) );
  OAI211_X1 U18115 ( .C1(n14829), .C2(n19079), .A(n14828), .B(n14827), .ZN(
        P2_U2898) );
  NOR2_X1 U18116 ( .A1(n14832), .A2(n14831), .ZN(n14833) );
  NOR2_X1 U18117 ( .A1(n14830), .A2(n14833), .ZN(n18838) );
  OAI22_X1 U18118 ( .A1(n19076), .A2(n14841), .B1(n19044), .B2(n14834), .ZN(
        n14835) );
  AOI21_X1 U18119 ( .B1(n19084), .B2(n18838), .A(n14835), .ZN(n14837) );
  AOI22_X1 U18120 ( .A1(n16048), .A2(BUF2_REG_19__SCAN_IN), .B1(n16049), .B2(
        BUF1_REG_19__SCAN_IN), .ZN(n14836) );
  OAI211_X1 U18121 ( .C1(n14838), .C2(n19079), .A(n14837), .B(n14836), .ZN(
        P2_U2900) );
  INV_X1 U18122 ( .A(n14839), .ZN(n18862) );
  OAI22_X1 U18123 ( .A1(n19158), .A2(n14841), .B1(n19044), .B2(n14840), .ZN(
        n14842) );
  AOI21_X1 U18124 ( .B1(n19084), .B2(n18862), .A(n14842), .ZN(n14844) );
  AOI22_X1 U18125 ( .A1(n16048), .A2(BUF2_REG_17__SCAN_IN), .B1(n16049), .B2(
        BUF1_REG_17__SCAN_IN), .ZN(n14843) );
  OAI211_X1 U18126 ( .C1(n14845), .C2(n19079), .A(n14844), .B(n14843), .ZN(
        P2_U2902) );
  NAND4_X1 U18127 ( .A1(n15047), .A2(n15068), .A3(n16072), .A4(n15058), .ZN(
        n14847) );
  NOR2_X1 U18128 ( .A1(n14848), .A2(n14847), .ZN(n14852) );
  NOR2_X1 U18129 ( .A1(n14850), .A2(n14849), .ZN(n14851) );
  AND3_X1 U18130 ( .A1(n14853), .A2(n14852), .A3(n14851), .ZN(n14862) );
  AND4_X1 U18131 ( .A1(n16073), .A2(n14854), .A3(n15057), .A4(n15069), .ZN(
        n14856) );
  AND4_X1 U18132 ( .A1(n14857), .A2(n14856), .A3(n14855), .A4(n15026), .ZN(
        n14859) );
  NAND3_X1 U18133 ( .A1(n14860), .A2(n14859), .A3(n14858), .ZN(n14861) );
  INV_X1 U18134 ( .A(n14863), .ZN(n14864) );
  NAND2_X1 U18135 ( .A1(n14865), .A2(n14864), .ZN(n14866) );
  NAND2_X1 U18136 ( .A1(n14868), .A2(n14866), .ZN(n15573) );
  INV_X1 U18137 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15241) );
  AOI21_X1 U18138 ( .B1(n14869), .B2(n14868), .A(n10121), .ZN(n16012) );
  NAND2_X1 U18139 ( .A1(n16012), .A2(n11060), .ZN(n14870) );
  XNOR2_X1 U18140 ( .A(n14870), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15008) );
  INV_X1 U18141 ( .A(n16012), .ZN(n14871) );
  INV_X1 U18142 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n14919) );
  NOR2_X1 U18143 ( .A1(n10808), .A2(n14874), .ZN(n14873) );
  MUX2_X1 U18144 ( .A(n14874), .B(n14873), .S(n14872), .Z(n14875) );
  NOR2_X1 U18145 ( .A1(n14875), .A2(n10104), .ZN(n15997) );
  NAND2_X1 U18146 ( .A1(n15997), .A2(n11060), .ZN(n14997) );
  NAND2_X1 U18147 ( .A1(n14877), .A2(n14876), .ZN(n14977) );
  NAND2_X1 U18148 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(n14878), .ZN(n14879) );
  NOR2_X1 U18149 ( .A1(n10808), .A2(n14879), .ZN(n14880) );
  AND2_X1 U18150 ( .A1(n11060), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14881) );
  NAND2_X1 U18151 ( .A1(n15975), .A2(n14881), .ZN(n14904) );
  INV_X1 U18152 ( .A(n15975), .ZN(n14882) );
  INV_X1 U18153 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15185) );
  OAI21_X1 U18154 ( .B1(n14882), .B2(n10849), .A(n15185), .ZN(n14883) );
  NAND2_X1 U18155 ( .A1(n14904), .A2(n14883), .ZN(n14979) );
  NOR2_X1 U18156 ( .A1(n14889), .A2(n14888), .ZN(n14884) );
  NAND2_X1 U18157 ( .A1(n14912), .A2(n14884), .ZN(n14885) );
  NAND2_X1 U18158 ( .A1(n14886), .A2(n14885), .ZN(n14887) );
  AOI21_X1 U18159 ( .B1(n14889), .B2(n14888), .A(n14887), .ZN(n15986) );
  NOR2_X1 U18160 ( .A1(n14902), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14988) );
  NAND2_X1 U18161 ( .A1(n14891), .A2(n14890), .ZN(n14892) );
  NOR2_X2 U18162 ( .A1(n14977), .A2(n14892), .ZN(n14956) );
  OR2_X1 U18163 ( .A1(n14894), .A2(n14893), .ZN(n14895) );
  NAND2_X1 U18164 ( .A1(n14896), .A2(n14895), .ZN(n15966) );
  NAND2_X1 U18165 ( .A1(n14956), .A2(n10232), .ZN(n14899) );
  OAI21_X1 U18166 ( .B1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(n14960), .ZN(n14898) );
  INV_X1 U18167 ( .A(n14960), .ZN(n14900) );
  INV_X1 U18168 ( .A(n14902), .ZN(n14903) );
  INV_X1 U18169 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15192) );
  NAND2_X1 U18170 ( .A1(n14986), .A2(n14904), .ZN(n14955) );
  XNOR2_X1 U18171 ( .A(n14906), .B(n14905), .ZN(n14909) );
  OAI21_X1 U18172 ( .B1(n14909), .B2(n10849), .A(n15147), .ZN(n14944) );
  AOI21_X1 U18173 ( .B1(n14908), .B2(n11060), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14935) );
  AND2_X1 U18174 ( .A1(n11060), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14907) );
  NAND2_X1 U18175 ( .A1(n14908), .A2(n14907), .ZN(n14933) );
  INV_X1 U18176 ( .A(n14909), .ZN(n15952) );
  NAND3_X1 U18177 ( .A1(n15952), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n11060), .ZN(n14945) );
  INV_X1 U18178 ( .A(n14910), .ZN(n14914) );
  NOR2_X1 U18179 ( .A1(n14911), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n14913) );
  MUX2_X1 U18180 ( .A(n14914), .B(n14913), .S(n14912), .Z(n15941) );
  NAND2_X1 U18181 ( .A1(n15941), .A2(n11060), .ZN(n14915) );
  XNOR2_X1 U18182 ( .A(n14915), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14916) );
  XNOR2_X1 U18183 ( .A(n14917), .B(n14916), .ZN(n15130) );
  NAND2_X1 U18184 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15122) );
  XNOR2_X1 U18185 ( .A(n14939), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n15128) );
  INV_X1 U18186 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n19775) );
  NAND2_X1 U18187 ( .A1(n10992), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n14921) );
  NAND2_X1 U18188 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n14920) );
  OAI211_X1 U18189 ( .C1(n9775), .C2(n19775), .A(n14921), .B(n14920), .ZN(
        n14923) );
  AOI21_X1 U18190 ( .B1(n14924), .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A(
        n14923), .ZN(n14925) );
  XNOR2_X2 U18191 ( .A(n14926), .B(n14925), .ZN(n16020) );
  NOR2_X1 U18192 ( .A1(n9889), .A2(n19775), .ZN(n15115) );
  NOR2_X1 U18193 ( .A1(n16068), .A2(n14927), .ZN(n14928) );
  AOI211_X1 U18194 ( .C1(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .C2(n16062), .A(
        n15115), .B(n14928), .ZN(n14929) );
  OAI21_X1 U18195 ( .B1(n16020), .B2(n16088), .A(n14929), .ZN(n14930) );
  AOI21_X1 U18196 ( .B1(n15128), .B2(n16120), .A(n14930), .ZN(n14931) );
  OAI21_X1 U18197 ( .B1(n15130), .B2(n15067), .A(n14931), .ZN(P2_U2983) );
  NAND2_X1 U18198 ( .A1(n14932), .A2(n14945), .ZN(n14937) );
  INV_X1 U18199 ( .A(n14933), .ZN(n14934) );
  NOR2_X1 U18200 ( .A1(n14935), .A2(n14934), .ZN(n14936) );
  XNOR2_X1 U18201 ( .A(n14937), .B(n14936), .ZN(n15141) );
  OR2_X1 U18202 ( .A1(n15149), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14938) );
  AND2_X1 U18203 ( .A1(n14939), .A2(n14938), .ZN(n15139) );
  NOR2_X1 U18204 ( .A1(n9889), .A2(n19772), .ZN(n15132) );
  NOR2_X1 U18205 ( .A1(n16068), .A2(n15948), .ZN(n14940) );
  AOI211_X1 U18206 ( .C1(n16062), .C2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n15132), .B(n14940), .ZN(n14941) );
  OAI21_X1 U18207 ( .B1(n15137), .B2(n16088), .A(n14941), .ZN(n14942) );
  AOI21_X1 U18208 ( .B1(n15139), .B2(n16120), .A(n14942), .ZN(n14943) );
  OAI21_X1 U18209 ( .B1(n15141), .B2(n15067), .A(n14943), .ZN(P2_U2984) );
  NAND2_X1 U18210 ( .A1(n14945), .A2(n14944), .ZN(n14947) );
  XOR2_X1 U18211 ( .A(n14947), .B(n14946), .Z(n15154) );
  INV_X1 U18212 ( .A(n14948), .ZN(n15954) );
  NAND2_X1 U18213 ( .A1(n16114), .A2(n14949), .ZN(n14950) );
  NAND2_X1 U18214 ( .A1(n16186), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n15143) );
  OAI211_X1 U18215 ( .C1(n16125), .C2(n14951), .A(n14950), .B(n15143), .ZN(
        n14953) );
  NOR2_X1 U18216 ( .A1(n14963), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15150) );
  NOR3_X1 U18217 ( .A1(n15149), .A2(n15150), .A3(n16055), .ZN(n14952) );
  OAI21_X1 U18218 ( .B1(n15154), .B2(n15067), .A(n14954), .ZN(P2_U2985) );
  INV_X1 U18219 ( .A(n14957), .ZN(n14958) );
  XNOR2_X1 U18220 ( .A(n14960), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14961) );
  XNOR2_X1 U18221 ( .A(n14962), .B(n14961), .ZN(n15167) );
  AOI21_X1 U18222 ( .B1(n9792), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14964) );
  NOR2_X1 U18223 ( .A1(n14964), .A2(n14963), .ZN(n15165) );
  NOR2_X1 U18224 ( .A1(n15163), .A2(n16088), .ZN(n14968) );
  NAND2_X1 U18225 ( .A1(n16186), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n15158) );
  NAND2_X1 U18226 ( .A1(n16062), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14965) );
  OAI211_X1 U18227 ( .C1(n16068), .C2(n14966), .A(n15158), .B(n14965), .ZN(
        n14967) );
  AOI211_X1 U18228 ( .C1(n15165), .C2(n16120), .A(n14968), .B(n14967), .ZN(
        n14969) );
  OAI21_X1 U18229 ( .B1(n15167), .B2(n15067), .A(n14969), .ZN(P2_U2986) );
  XNOR2_X1 U18230 ( .A(n14970), .B(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15179) );
  XNOR2_X1 U18231 ( .A(n14971), .B(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15176) );
  INV_X1 U18232 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n19765) );
  NOR2_X1 U18233 ( .A1(n9889), .A2(n19765), .ZN(n15171) );
  AOI21_X1 U18234 ( .B1(n16062), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n15171), .ZN(n14974) );
  NAND2_X1 U18235 ( .A1(n16114), .A2(n14972), .ZN(n14973) );
  OAI211_X1 U18236 ( .C1(n15168), .C2(n16088), .A(n14974), .B(n14973), .ZN(
        n14975) );
  AOI21_X1 U18237 ( .B1(n15176), .B2(n16120), .A(n14975), .ZN(n14976) );
  OAI21_X1 U18238 ( .B1(n15179), .B2(n15067), .A(n14976), .ZN(P2_U2987) );
  AOI21_X1 U18239 ( .B1(n14977), .B2(n14986), .A(n14988), .ZN(n14978) );
  XOR2_X1 U18240 ( .A(n14979), .B(n14978), .Z(n15190) );
  AOI21_X1 U18241 ( .B1(n15185), .B2(n14980), .A(n9792), .ZN(n15188) );
  NOR2_X1 U18242 ( .A1(n9889), .A2(n19762), .ZN(n15182) );
  NOR2_X1 U18243 ( .A1(n16068), .A2(n15981), .ZN(n14981) );
  AOI211_X1 U18244 ( .C1(n16062), .C2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n15182), .B(n14981), .ZN(n14982) );
  OAI21_X1 U18245 ( .B1(n15977), .B2(n16088), .A(n14982), .ZN(n14983) );
  AOI21_X1 U18246 ( .B1(n15188), .B2(n16120), .A(n14983), .ZN(n14984) );
  OAI21_X1 U18247 ( .B1(n15190), .B2(n15067), .A(n14984), .ZN(P2_U2988) );
  OR2_X1 U18248 ( .A1(n14999), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14985) );
  NAND2_X1 U18249 ( .A1(n14980), .A2(n14985), .ZN(n15203) );
  INV_X1 U18250 ( .A(n14986), .ZN(n14987) );
  NOR2_X1 U18251 ( .A1(n14988), .A2(n14987), .ZN(n14989) );
  XNOR2_X1 U18252 ( .A(n14977), .B(n14989), .ZN(n15191) );
  NAND2_X1 U18253 ( .A1(n15191), .A2(n16118), .ZN(n14995) );
  NAND2_X1 U18254 ( .A1(n16186), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n15195) );
  OAI21_X1 U18255 ( .B1(n16125), .B2(n14990), .A(n15195), .ZN(n14992) );
  NOR2_X1 U18256 ( .A1(n15988), .A2(n16088), .ZN(n14991) );
  AOI211_X1 U18257 ( .C1(n16114), .C2(n14993), .A(n14992), .B(n14991), .ZN(
        n14994) );
  OAI211_X1 U18258 ( .C1(n16055), .C2(n15203), .A(n14995), .B(n14994), .ZN(
        P2_U2989) );
  XOR2_X1 U18259 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n14997), .Z(
        n14998) );
  XNOR2_X1 U18260 ( .A(n14996), .B(n14998), .ZN(n15213) );
  AOI21_X1 U18261 ( .B1(n20991), .B2(n15005), .A(n14999), .ZN(n15211) );
  AND2_X1 U18262 ( .A1(n18976), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n15204) );
  AOI21_X1 U18263 ( .B1(n16062), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n15204), .ZN(n15002) );
  INV_X1 U18264 ( .A(n16002), .ZN(n15000) );
  NAND2_X1 U18265 ( .A1(n16114), .A2(n15000), .ZN(n15001) );
  OAI211_X1 U18266 ( .C1(n15209), .C2(n16088), .A(n15002), .B(n15001), .ZN(
        n15003) );
  AOI21_X1 U18267 ( .B1(n15211), .B2(n16120), .A(n15003), .ZN(n15004) );
  OAI21_X1 U18268 ( .B1(n15213), .B2(n15067), .A(n15004), .ZN(P2_U2990) );
  INV_X1 U18269 ( .A(n15227), .ZN(n15006) );
  OAI21_X1 U18270 ( .B1(n15006), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n15005), .ZN(n15225) );
  XOR2_X1 U18271 ( .A(n15008), .B(n15007), .Z(n15214) );
  NAND2_X1 U18272 ( .A1(n15214), .A2(n16118), .ZN(n15013) );
  NAND2_X1 U18273 ( .A1(n16186), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n15216) );
  OAI21_X1 U18274 ( .B1(n16125), .B2(n12091), .A(n15216), .ZN(n15010) );
  NOR2_X1 U18275 ( .A1(n16010), .A2(n16088), .ZN(n15009) );
  AOI211_X1 U18276 ( .C1(n16114), .C2(n15011), .A(n15010), .B(n15009), .ZN(
        n15012) );
  OAI211_X1 U18277 ( .C1(n16055), .C2(n15225), .A(n15013), .B(n15012), .ZN(
        P2_U2991) );
  OAI21_X1 U18278 ( .B1(n15016), .B2(n15015), .A(n15014), .ZN(n15259) );
  OR2_X1 U18279 ( .A1(n15018), .A2(n15017), .ZN(n15019) );
  NAND2_X1 U18280 ( .A1(n12255), .A2(n15019), .ZN(n18825) );
  INV_X1 U18281 ( .A(n18825), .ZN(n15024) );
  INV_X1 U18282 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n15020) );
  NOR2_X1 U18283 ( .A1(n9889), .A2(n15020), .ZN(n15250) );
  AOI21_X1 U18284 ( .B1(n16062), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n15250), .ZN(n15021) );
  OAI21_X1 U18285 ( .B1(n18829), .B2(n16068), .A(n15021), .ZN(n15023) );
  XOR2_X1 U18286 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .B(n15034), .Z(
        n15254) );
  NOR2_X1 U18287 ( .A1(n15254), .A2(n16055), .ZN(n15022) );
  AOI211_X1 U18288 ( .C1(n16117), .C2(n15024), .A(n15023), .B(n15022), .ZN(
        n15025) );
  OAI21_X1 U18289 ( .B1(n15259), .B2(n15067), .A(n15025), .ZN(P2_U2994) );
  NAND2_X1 U18290 ( .A1(n15027), .A2(n15026), .ZN(n15030) );
  INV_X1 U18291 ( .A(n15028), .ZN(n15264) );
  NOR2_X1 U18292 ( .A1(n15260), .A2(n15264), .ZN(n15029) );
  XOR2_X1 U18293 ( .A(n15030), .B(n15029), .Z(n16135) );
  INV_X1 U18294 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n21044) );
  OAI22_X1 U18295 ( .A1(n16125), .A2(n18834), .B1(n21044), .B2(n9889), .ZN(
        n15032) );
  NOR2_X1 U18296 ( .A1(n16131), .A2(n16088), .ZN(n15031) );
  AOI211_X1 U18297 ( .C1(n15033), .C2(n16114), .A(n15032), .B(n15031), .ZN(
        n15037) );
  INV_X1 U18298 ( .A(n15034), .ZN(n15035) );
  AOI21_X1 U18299 ( .B1(n16129), .B2(n9784), .A(n15035), .ZN(n16132) );
  NAND2_X1 U18300 ( .A1(n16132), .A2(n16120), .ZN(n15036) );
  OAI211_X1 U18301 ( .C1(n16135), .C2(n15067), .A(n15037), .B(n15036), .ZN(
        P2_U2995) );
  NOR2_X1 U18302 ( .A1(n19748), .A2(n9889), .ZN(n15040) );
  INV_X1 U18303 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n15038) );
  OAI22_X1 U18304 ( .A1(n16125), .A2(n15038), .B1(n16068), .B2(n18866), .ZN(
        n15039) );
  AOI211_X1 U18305 ( .C1(n16117), .C2(n18863), .A(n15040), .B(n15039), .ZN(
        n15043) );
  INV_X1 U18306 ( .A(n15271), .ZN(n15041) );
  NAND2_X1 U18307 ( .A1(n15095), .A2(n15041), .ZN(n15266) );
  OAI211_X1 U18308 ( .C1(n15045), .C2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n16120), .B(n15266), .ZN(n15042) );
  OAI211_X1 U18309 ( .C1(n15044), .C2(n15067), .A(n15043), .B(n15042), .ZN(
        P2_U2997) );
  AOI211_X1 U18310 ( .C1(n15290), .C2(n15062), .A(n16055), .B(n15045), .ZN(
        n15056) );
  OAI21_X1 U18311 ( .B1(n9840), .B2(n15047), .A(n15046), .ZN(n15285) );
  NOR2_X1 U18312 ( .A1(n15285), .A2(n15067), .ZN(n15055) );
  OR2_X1 U18313 ( .A1(n15049), .A2(n15048), .ZN(n15050) );
  NAND2_X1 U18314 ( .A1(n15051), .A2(n15050), .ZN(n19010) );
  NAND2_X1 U18315 ( .A1(n18976), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n15284) );
  OAI21_X1 U18316 ( .B1(n16125), .B2(n18882), .A(n15284), .ZN(n15052) );
  AOI21_X1 U18317 ( .B1(n16114), .B2(n18875), .A(n15052), .ZN(n15053) );
  OAI21_X1 U18318 ( .B1(n19010), .B2(n16088), .A(n15053), .ZN(n15054) );
  OR3_X1 U18319 ( .A1(n15056), .A2(n15055), .A3(n15054), .ZN(P2_U2998) );
  NAND2_X1 U18320 ( .A1(n15058), .A2(n15057), .ZN(n15059) );
  XNOR2_X1 U18321 ( .A(n15060), .B(n15059), .ZN(n15303) );
  INV_X1 U18322 ( .A(n18887), .ZN(n15065) );
  AND2_X1 U18323 ( .A1(n18976), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n15292) );
  AOI21_X1 U18324 ( .B1(n16062), .B2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n15292), .ZN(n15061) );
  OAI21_X1 U18325 ( .B1(n18889), .B2(n16088), .A(n15061), .ZN(n15064) );
  OAI21_X1 U18326 ( .B1(n16070), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n15062), .ZN(n15298) );
  NOR2_X1 U18327 ( .A1(n15298), .A2(n16055), .ZN(n15063) );
  AOI211_X1 U18328 ( .C1(n16114), .C2(n15065), .A(n15064), .B(n15063), .ZN(
        n15066) );
  OAI21_X1 U18329 ( .B1(n15303), .B2(n15067), .A(n15066), .ZN(P2_U2999) );
  NOR2_X1 U18330 ( .A1(n16081), .A2(n16161), .ZN(n16080) );
  INV_X1 U18331 ( .A(n16081), .ZN(n15085) );
  NAND2_X1 U18332 ( .A1(n15085), .A2(n16143), .ZN(n16071) );
  OAI21_X1 U18333 ( .B1(n16080), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n16071), .ZN(n16156) );
  NAND2_X1 U18334 ( .A1(n15069), .A2(n15068), .ZN(n15070) );
  XNOR2_X1 U18335 ( .A(n15071), .B(n15070), .ZN(n16153) );
  INV_X1 U18336 ( .A(n18896), .ZN(n18902) );
  AOI22_X1 U18337 ( .A1(n16062), .A2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .B1(
        n16114), .B2(n18902), .ZN(n15073) );
  NAND2_X1 U18338 ( .A1(n18976), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n15072) );
  OAI211_X1 U18339 ( .C1(n15074), .C2(n16088), .A(n15073), .B(n15072), .ZN(
        n15075) );
  AOI21_X1 U18340 ( .B1(n16153), .B2(n16118), .A(n15075), .ZN(n15076) );
  OAI21_X1 U18341 ( .B1(n16156), .B2(n16055), .A(n15076), .ZN(P2_U3001) );
  NAND2_X1 U18342 ( .A1(n15077), .A2(n9872), .ZN(n15082) );
  INV_X1 U18343 ( .A(n15078), .ZN(n15079) );
  NOR2_X1 U18344 ( .A1(n15080), .A2(n15079), .ZN(n15081) );
  XNOR2_X1 U18345 ( .A(n15082), .B(n15081), .ZN(n16179) );
  INV_X1 U18346 ( .A(n15083), .ZN(n15084) );
  AOI21_X1 U18347 ( .B1(n15084), .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15086) );
  NOR2_X1 U18348 ( .A1(n15086), .A2(n15085), .ZN(n16176) );
  NAND2_X1 U18349 ( .A1(n16176), .A2(n16120), .ZN(n15090) );
  NOR2_X1 U18350 ( .A1(n9889), .A2(n15087), .ZN(n16174) );
  OAI22_X1 U18351 ( .A1(n16125), .A2(n10040), .B1(n16068), .B2(n18921), .ZN(
        n15088) );
  AOI211_X1 U18352 ( .C1(n18907), .C2(n16117), .A(n16174), .B(n15088), .ZN(
        n15089) );
  OAI211_X1 U18353 ( .C1(n16179), .C2(n15067), .A(n15090), .B(n15089), .ZN(
        P2_U3003) );
  INV_X1 U18354 ( .A(n15091), .ZN(n15313) );
  NOR2_X1 U18355 ( .A1(n15092), .A2(n15313), .ZN(n15094) );
  XOR2_X1 U18356 ( .A(n15094), .B(n15093), .Z(n15332) );
  INV_X1 U18357 ( .A(n15095), .ZN(n15096) );
  NAND2_X1 U18358 ( .A1(n15096), .A2(n15328), .ZN(n15323) );
  NAND3_X1 U18359 ( .A1(n15323), .A2(n16120), .A3(n15083), .ZN(n15100) );
  INV_X1 U18360 ( .A(n15325), .ZN(n18942) );
  NOR2_X1 U18361 ( .A1(n16088), .A2(n18942), .ZN(n15098) );
  OAI22_X1 U18362 ( .A1(n16125), .A2(n10049), .B1(n16068), .B2(n18940), .ZN(
        n15097) );
  AOI211_X1 U18363 ( .C1(n18976), .C2(P2_REIP_REG_9__SCAN_IN), .A(n15098), .B(
        n15097), .ZN(n15099) );
  OAI211_X1 U18364 ( .C1(n15067), .C2(n15332), .A(n15100), .B(n15099), .ZN(
        P2_U3005) );
  INV_X1 U18365 ( .A(n16101), .ZN(n15102) );
  NOR2_X1 U18366 ( .A1(n15102), .A2(n16100), .ZN(n15103) );
  XNOR2_X1 U18367 ( .A(n15101), .B(n15103), .ZN(n15343) );
  OR2_X1 U18368 ( .A1(n15105), .A2(n15104), .ZN(n15334) );
  NAND3_X1 U18369 ( .A1(n15334), .A2(n15333), .A3(n16120), .ZN(n15110) );
  NOR2_X1 U18370 ( .A1(n16088), .A2(n18953), .ZN(n15108) );
  INV_X1 U18371 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n15106) );
  OAI22_X1 U18372 ( .A1(n16125), .A2(n15106), .B1(n16068), .B2(n18949), .ZN(
        n15107) );
  AOI211_X1 U18373 ( .C1(n18976), .C2(P2_REIP_REG_7__SCAN_IN), .A(n15108), .B(
        n15107), .ZN(n15109) );
  OAI211_X1 U18374 ( .C1(n15343), .C2(n15067), .A(n15110), .B(n15109), .ZN(
        P2_U3007) );
  NAND3_X1 U18375 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(n15215), .ZN(n15117) );
  NOR2_X1 U18376 ( .A1(n15117), .A2(n15111), .ZN(n15206) );
  NOR2_X1 U18377 ( .A1(n15185), .A2(n15192), .ZN(n15180) );
  AND2_X1 U18378 ( .A1(n15206), .A2(n15180), .ZN(n15112) );
  NAND2_X1 U18379 ( .A1(n10150), .A2(n15156), .ZN(n15144) );
  INV_X1 U18380 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15113) );
  NOR4_X1 U18381 ( .A1(n15144), .A2(n15147), .A3(n15113), .A4(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n15114) );
  AOI21_X1 U18382 ( .B1(n16138), .B2(n15117), .A(n20991), .ZN(n15118) );
  NAND2_X1 U18383 ( .A1(n16136), .A2(n15118), .ZN(n15205) );
  INV_X1 U18384 ( .A(n15304), .ZN(n15120) );
  NAND2_X1 U18385 ( .A1(n15205), .A2(n15120), .ZN(n15193) );
  INV_X1 U18386 ( .A(n15180), .ZN(n15119) );
  NAND2_X1 U18387 ( .A1(n15120), .A2(n15119), .ZN(n15121) );
  AND2_X1 U18388 ( .A1(n15193), .A2(n15121), .ZN(n15170) );
  OAI21_X1 U18389 ( .B1(n15122), .B2(n15147), .A(n16138), .ZN(n15123) );
  NAND2_X1 U18390 ( .A1(n15170), .A2(n15123), .ZN(n15134) );
  NOR2_X1 U18391 ( .A1(n15357), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15124) );
  OAI21_X1 U18392 ( .B1(n15134), .B2(n15124), .A(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n15125) );
  OAI211_X1 U18393 ( .C1(n16020), .C2(n15360), .A(n15126), .B(n15125), .ZN(
        n15127) );
  AOI21_X1 U18394 ( .B1(n15128), .B2(n21137), .A(n15127), .ZN(n15129) );
  OAI21_X1 U18395 ( .B1(n15130), .B2(n21140), .A(n15129), .ZN(P2_U3015) );
  NOR3_X1 U18396 ( .A1(n15144), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n15147), .ZN(n15131) );
  NAND2_X1 U18397 ( .A1(n15134), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15135) );
  OAI211_X1 U18398 ( .C1(n15137), .C2(n15360), .A(n15136), .B(n15135), .ZN(
        n15138) );
  AOI21_X1 U18399 ( .B1(n15139), .B2(n21137), .A(n15138), .ZN(n15140) );
  OAI21_X1 U18400 ( .B1(n15141), .B2(n21140), .A(n15140), .ZN(P2_U3016) );
  NAND2_X1 U18401 ( .A1(n15156), .A2(n15169), .ZN(n15173) );
  NAND2_X1 U18402 ( .A1(n15170), .A2(n15173), .ZN(n15161) );
  AOI21_X1 U18403 ( .B1(n15156), .B2(n15155), .A(n15161), .ZN(n15148) );
  INV_X1 U18404 ( .A(n15142), .ZN(n15953) );
  OAI21_X1 U18405 ( .B1(n15144), .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n15143), .ZN(n15145) );
  AOI21_X1 U18406 ( .B1(n16181), .B2(n15953), .A(n15145), .ZN(n15146) );
  OAI21_X1 U18407 ( .B1(n15148), .B2(n15147), .A(n15146), .ZN(n15152) );
  NOR3_X1 U18408 ( .A1(n15150), .A2(n15149), .A3(n16157), .ZN(n15151) );
  NAND3_X1 U18409 ( .A1(n15156), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        n15155), .ZN(n15157) );
  OAI211_X1 U18410 ( .C1(n21133), .C2(n15159), .A(n15158), .B(n15157), .ZN(
        n15160) );
  AOI21_X1 U18411 ( .B1(n15161), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n15160), .ZN(n15162) );
  OAI21_X1 U18412 ( .B1(n15163), .B2(n15360), .A(n15162), .ZN(n15164) );
  AOI21_X1 U18413 ( .B1(n15165), .B2(n21137), .A(n15164), .ZN(n15166) );
  OAI21_X1 U18414 ( .B1(n15167), .B2(n21140), .A(n15166), .ZN(P2_U3018) );
  INV_X1 U18415 ( .A(n15168), .ZN(n15968) );
  NOR2_X1 U18416 ( .A1(n15170), .A2(n15169), .ZN(n15175) );
  INV_X1 U18417 ( .A(n15171), .ZN(n15172) );
  OAI211_X1 U18418 ( .C1(n21133), .C2(n15974), .A(n15173), .B(n15172), .ZN(
        n15174) );
  AOI211_X1 U18419 ( .C1(n15968), .C2(n21130), .A(n15175), .B(n15174), .ZN(
        n15178) );
  NAND2_X1 U18420 ( .A1(n15176), .A2(n21137), .ZN(n15177) );
  OAI211_X1 U18421 ( .C1(n15179), .C2(n21140), .A(n15178), .B(n15177), .ZN(
        P2_U3019) );
  NOR2_X1 U18422 ( .A1(n15977), .A2(n15360), .ZN(n15187) );
  INV_X1 U18423 ( .A(n15976), .ZN(n15183) );
  NAND2_X1 U18424 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n15206), .ZN(
        n15197) );
  AOI211_X1 U18425 ( .C1(n15185), .C2(n15192), .A(n15180), .B(n15197), .ZN(
        n15181) );
  AOI211_X1 U18426 ( .C1(n16181), .C2(n15183), .A(n15182), .B(n15181), .ZN(
        n15184) );
  OAI21_X1 U18427 ( .B1(n15193), .B2(n15185), .A(n15184), .ZN(n15186) );
  AOI211_X1 U18428 ( .C1(n15188), .C2(n21137), .A(n15187), .B(n15186), .ZN(
        n15189) );
  OAI21_X1 U18429 ( .B1(n15190), .B2(n21140), .A(n15189), .ZN(P2_U3020) );
  NAND2_X1 U18430 ( .A1(n15191), .A2(n11126), .ZN(n15202) );
  INV_X1 U18431 ( .A(n15988), .ZN(n15200) );
  NOR2_X1 U18432 ( .A1(n15193), .A2(n15192), .ZN(n15199) );
  NAND2_X1 U18433 ( .A1(n16181), .A2(n15194), .ZN(n15196) );
  OAI211_X1 U18434 ( .C1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .C2(n15197), .A(
        n15196), .B(n15195), .ZN(n15198) );
  AOI211_X1 U18435 ( .C1(n15200), .C2(n21130), .A(n15199), .B(n15198), .ZN(
        n15201) );
  OAI211_X1 U18436 ( .C1(n15203), .C2(n16157), .A(n15202), .B(n15201), .ZN(
        P2_U3021) );
  AOI21_X1 U18437 ( .B1(n16181), .B2(n15998), .A(n15204), .ZN(n15208) );
  OAI21_X1 U18438 ( .B1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n15206), .A(
        n15205), .ZN(n15207) );
  OAI211_X1 U18439 ( .C1(n15209), .C2(n15360), .A(n15208), .B(n15207), .ZN(
        n15210) );
  AOI21_X1 U18440 ( .B1(n15211), .B2(n21137), .A(n15210), .ZN(n15212) );
  OAI21_X1 U18441 ( .B1(n15213), .B2(n21140), .A(n15212), .ZN(P2_U3022) );
  NAND2_X1 U18442 ( .A1(n15214), .A2(n11126), .ZN(n15224) );
  NAND2_X1 U18443 ( .A1(n15215), .A2(n15329), .ZN(n15242) );
  XNOR2_X1 U18444 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15217) );
  OAI21_X1 U18445 ( .B1(n15242), .B2(n15217), .A(n15216), .ZN(n15218) );
  AOI21_X1 U18446 ( .B1(n16181), .B2(n15219), .A(n15218), .ZN(n15220) );
  OAI21_X1 U18447 ( .B1(n16010), .B2(n15360), .A(n15220), .ZN(n15221) );
  AOI21_X1 U18448 ( .B1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n15222), .A(
        n15221), .ZN(n15223) );
  OAI211_X1 U18449 ( .C1(n15225), .C2(n16157), .A(n15224), .B(n15223), .ZN(
        P2_U3023) );
  NAND2_X1 U18450 ( .A1(n14918), .A2(n15241), .ZN(n15226) );
  NAND2_X1 U18451 ( .A1(n15227), .A2(n15226), .ZN(n16056) );
  INV_X1 U18452 ( .A(n15229), .ZN(n15231) );
  NOR2_X1 U18453 ( .A1(n15231), .A2(n15230), .ZN(n15232) );
  XNOR2_X1 U18454 ( .A(n15228), .B(n15232), .ZN(n16058) );
  NAND2_X1 U18455 ( .A1(n16058), .A2(n11126), .ZN(n15246) );
  AOI21_X1 U18456 ( .B1(n15234), .B2(n15233), .A(n14816), .ZN(n16034) );
  NAND2_X1 U18457 ( .A1(n15236), .A2(n15235), .ZN(n15237) );
  NAND2_X1 U18458 ( .A1(n15238), .A2(n15237), .ZN(n16054) );
  NOR2_X1 U18459 ( .A1(n16054), .A2(n15360), .ZN(n15244) );
  NAND2_X1 U18460 ( .A1(P2_REIP_REG_22__SCAN_IN), .A2(n18976), .ZN(n15239) );
  OAI221_X1 U18461 ( .B1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n15242), 
        .C1(n15241), .C2(n15240), .A(n15239), .ZN(n15243) );
  AOI211_X1 U18462 ( .C1(n16181), .C2(n16034), .A(n15244), .B(n15243), .ZN(
        n15245) );
  OAI211_X1 U18463 ( .C1(n16056), .C2(n16157), .A(n15246), .B(n15245), .ZN(
        P2_U3024) );
  XNOR2_X1 U18464 ( .A(n16129), .B(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15257) );
  NOR2_X1 U18465 ( .A1(n14830), .A2(n15247), .ZN(n15248) );
  NOR2_X1 U18466 ( .A1(n15249), .A2(n15248), .ZN(n16039) );
  AOI21_X1 U18467 ( .B1(n16181), .B2(n16039), .A(n15250), .ZN(n15253) );
  OAI21_X1 U18468 ( .B1(n15251), .B2(n15357), .A(n16136), .ZN(n16128) );
  NAND2_X1 U18469 ( .A1(n16128), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15252) );
  OAI211_X1 U18470 ( .C1(n18825), .C2(n15360), .A(n15253), .B(n15252), .ZN(
        n15256) );
  NOR2_X1 U18471 ( .A1(n15254), .A2(n16157), .ZN(n15255) );
  AOI211_X1 U18472 ( .C1(n16130), .C2(n15257), .A(n15256), .B(n15255), .ZN(
        n15258) );
  OAI21_X1 U18473 ( .B1(n15259), .B2(n21140), .A(n15258), .ZN(P2_U3026) );
  INV_X1 U18474 ( .A(n15260), .ZN(n15265) );
  OAI21_X1 U18475 ( .B1(n15264), .B2(n15262), .A(n15261), .ZN(n15263) );
  OAI21_X1 U18476 ( .B1(n15265), .B2(n15264), .A(n15263), .ZN(n16065) );
  INV_X1 U18477 ( .A(n16065), .ZN(n15282) );
  NAND2_X1 U18478 ( .A1(n15266), .A2(n15278), .ZN(n15267) );
  AND2_X1 U18479 ( .A1(n15267), .A2(n12249), .ZN(n16063) );
  INV_X1 U18480 ( .A(n16128), .ZN(n15279) );
  AOI21_X1 U18481 ( .B1(n15269), .B2(n15268), .A(n14831), .ZN(n18849) );
  NAND2_X1 U18482 ( .A1(n15278), .A2(n15329), .ZN(n15270) );
  OAI22_X1 U18483 ( .A1(n15271), .A2(n15270), .B1(n12180), .B2(n9889), .ZN(
        n15276) );
  AND2_X1 U18484 ( .A1(n15273), .A2(n15272), .ZN(n15274) );
  OR2_X1 U18485 ( .A1(n15274), .A2(n14737), .ZN(n18851) );
  NOR2_X1 U18486 ( .A1(n18851), .A2(n15360), .ZN(n15275) );
  AOI211_X1 U18487 ( .C1(n18849), .C2(n16181), .A(n15276), .B(n15275), .ZN(
        n15277) );
  OAI21_X1 U18488 ( .B1(n15279), .B2(n15278), .A(n15277), .ZN(n15280) );
  AOI21_X1 U18489 ( .B1(n16063), .B2(n21137), .A(n15280), .ZN(n15281) );
  OAI21_X1 U18490 ( .B1(n15282), .B2(n21140), .A(n15281), .ZN(P2_U3028) );
  NAND2_X1 U18491 ( .A1(n16181), .A2(n18876), .ZN(n15283) );
  OAI211_X1 U18492 ( .C1(n19010), .C2(n15360), .A(n15284), .B(n15283), .ZN(
        n15287) );
  NOR2_X1 U18493 ( .A1(n15285), .A2(n21140), .ZN(n15286) );
  AOI211_X1 U18494 ( .C1(n15288), .C2(n15290), .A(n15287), .B(n15286), .ZN(
        n15289) );
  OAI21_X1 U18495 ( .B1(n15291), .B2(n15290), .A(n15289), .ZN(P2_U3030) );
  INV_X1 U18496 ( .A(n15292), .ZN(n15293) );
  OAI21_X1 U18497 ( .B1(n15294), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n15293), .ZN(n15295) );
  AOI21_X1 U18498 ( .B1(n16181), .B2(n15296), .A(n15295), .ZN(n15297) );
  OAI21_X1 U18499 ( .B1(n18889), .B2(n15360), .A(n15297), .ZN(n15300) );
  NOR2_X1 U18500 ( .A1(n15298), .A2(n16157), .ZN(n15299) );
  AOI211_X1 U18501 ( .C1(n15301), .C2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n15300), .B(n15299), .ZN(n15302) );
  OAI21_X1 U18502 ( .B1(n15303), .B2(n21140), .A(n15302), .ZN(P2_U3031) );
  XNOR2_X1 U18503 ( .A(n15083), .B(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n16093) );
  NAND2_X1 U18504 ( .A1(n16093), .A2(n21137), .ZN(n15322) );
  AOI21_X1 U18505 ( .B1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n16136), .A(
        n15304), .ZN(n16175) );
  NOR2_X1 U18506 ( .A1(n18926), .A2(n9889), .ZN(n15305) );
  AOI221_X1 U18507 ( .B1(n16175), .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), 
        .C1(n16170), .C2(n15306), .A(n15305), .ZN(n15321) );
  OAI21_X1 U18508 ( .B1(n15309), .B2(n15308), .A(n15307), .ZN(n19027) );
  INV_X1 U18509 ( .A(n19027), .ZN(n16094) );
  XNOR2_X1 U18510 ( .A(n15311), .B(n15310), .ZN(n19053) );
  INV_X1 U18511 ( .A(n19053), .ZN(n15312) );
  AOI22_X1 U18512 ( .A1(n21130), .A2(n16094), .B1(n16181), .B2(n15312), .ZN(
        n15320) );
  OR2_X1 U18513 ( .A1(n15314), .A2(n15313), .ZN(n15318) );
  NAND2_X1 U18514 ( .A1(n15316), .A2(n15315), .ZN(n15317) );
  XNOR2_X1 U18515 ( .A(n15318), .B(n15317), .ZN(n16095) );
  NAND2_X1 U18516 ( .A1(n16095), .A2(n11126), .ZN(n15319) );
  NAND4_X1 U18517 ( .A1(n15322), .A2(n15321), .A3(n15320), .A4(n15319), .ZN(
        P2_U3036) );
  NAND3_X1 U18518 ( .A1(n15323), .A2(n21137), .A3(n15083), .ZN(n15331) );
  INV_X1 U18519 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n19736) );
  OAI22_X1 U18520 ( .A1(n21133), .A2(n18941), .B1(n19736), .B2(n9889), .ZN(
        n15324) );
  AOI21_X1 U18521 ( .B1(n21130), .B2(n15325), .A(n15324), .ZN(n15326) );
  OAI21_X1 U18522 ( .B1(n16136), .B2(n15328), .A(n15326), .ZN(n15327) );
  AOI21_X1 U18523 ( .B1(n15329), .B2(n15328), .A(n15327), .ZN(n15330) );
  OAI211_X1 U18524 ( .C1(n15332), .C2(n21140), .A(n15331), .B(n15330), .ZN(
        P2_U3037) );
  NAND3_X1 U18525 ( .A1(n15334), .A2(n15333), .A3(n21137), .ZN(n15342) );
  INV_X1 U18526 ( .A(n15335), .ZN(n16188) );
  INV_X1 U18527 ( .A(n15336), .ZN(n16182) );
  OAI22_X1 U18528 ( .A1(n15360), .A2(n18953), .B1(n19733), .B2(n9889), .ZN(
        n15337) );
  AOI21_X1 U18529 ( .B1(n16182), .B2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n15337), .ZN(n15338) );
  OAI21_X1 U18530 ( .B1(n18954), .B2(n21133), .A(n15338), .ZN(n15339) );
  AOI21_X1 U18531 ( .B1(n16188), .B2(n15340), .A(n15339), .ZN(n15341) );
  OAI211_X1 U18532 ( .C1(n15343), .C2(n21140), .A(n15342), .B(n15341), .ZN(
        P2_U3039) );
  XOR2_X1 U18533 ( .A(n15345), .B(n15346), .Z(n16119) );
  NOR2_X1 U18534 ( .A1(n15348), .A2(n15347), .ZN(n15350) );
  NAND2_X1 U18535 ( .A1(n15350), .A2(n15349), .ZN(n15353) );
  INV_X1 U18536 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n19732) );
  OAI22_X1 U18537 ( .A1(n15360), .A2(n16116), .B1(n19732), .B2(n9889), .ZN(
        n15351) );
  AOI21_X1 U18538 ( .B1(n16182), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n15351), .ZN(n15352) );
  OAI211_X1 U18539 ( .C1(n21133), .C2(n18972), .A(n15353), .B(n15352), .ZN(
        n15354) );
  AOI21_X1 U18540 ( .B1(n16119), .B2(n11126), .A(n15354), .ZN(n15355) );
  OAI21_X1 U18541 ( .B1(n16115), .B2(n16157), .A(n15355), .ZN(P2_U3040) );
  MUX2_X1 U18542 ( .A(n15357), .B(n15356), .S(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .Z(n15367) );
  OAI21_X1 U18543 ( .B1(n15360), .B2(n15359), .A(n15358), .ZN(n15361) );
  AOI21_X1 U18544 ( .B1(n11126), .B2(n15362), .A(n15361), .ZN(n15366) );
  INV_X1 U18545 ( .A(n15363), .ZN(n19088) );
  AOI22_X1 U18546 ( .A1(n21137), .A2(n15364), .B1(n16181), .B2(n19088), .ZN(
        n15365) );
  NAND3_X1 U18547 ( .A1(n15367), .A2(n15366), .A3(n15365), .ZN(P2_U3046) );
  NOR2_X1 U18548 ( .A1(n14665), .A2(n15368), .ZN(n19000) );
  AOI21_X1 U18549 ( .B1(n14665), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n19000), .ZN(n15387) );
  NAND2_X1 U18550 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n15387), .ZN(n15376) );
  INV_X1 U18551 ( .A(n15369), .ZN(n15425) );
  NAND2_X1 U18552 ( .A1(n12319), .A2(n15425), .ZN(n15374) );
  INV_X1 U18553 ( .A(n15416), .ZN(n15392) );
  AND2_X1 U18554 ( .A1(n15370), .A2(n9779), .ZN(n15371) );
  NOR2_X1 U18555 ( .A1(n10531), .A2(n15371), .ZN(n15393) );
  MUX2_X1 U18556 ( .A(n15392), .B(n15393), .S(n15372), .Z(n15373) );
  NAND2_X1 U18557 ( .A1(n15374), .A2(n15373), .ZN(n16198) );
  NAND2_X1 U18558 ( .A1(n16198), .A2(n19784), .ZN(n15375) );
  OAI211_X1 U18559 ( .C1(n12327), .C2(n16244), .A(n15376), .B(n15375), .ZN(
        n15385) );
  NAND2_X1 U18560 ( .A1(n15377), .A2(n19835), .ZN(n15383) );
  INV_X1 U18561 ( .A(n15378), .ZN(n15379) );
  AND3_X1 U18562 ( .A1(n15381), .A2(n15380), .A3(n15379), .ZN(n15382) );
  INV_X1 U18563 ( .A(n19840), .ZN(n18788) );
  INV_X1 U18564 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n21000) );
  NOR2_X1 U18565 ( .A1(n19836), .A2(n19815), .ZN(n16248) );
  INV_X1 U18566 ( .A(n16248), .ZN(n16252) );
  OAI22_X1 U18567 ( .A1(n16232), .A2(n18788), .B1(n21000), .B2(n16252), .ZN(
        n15384) );
  AOI21_X1 U18568 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19836), .A(n15384), 
        .ZN(n15542) );
  MUX2_X1 U18569 ( .A(n15385), .B(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .S(
        n15542), .Z(P2_U3601) );
  OR2_X1 U18570 ( .A1(n15387), .A2(n15386), .ZN(n15408) );
  OAI21_X1 U18571 ( .B1(n12116), .B2(n15389), .A(n15388), .ZN(n15407) );
  INV_X1 U18572 ( .A(n15390), .ZN(n15399) );
  OAI22_X1 U18573 ( .A1(n15393), .A2(n15391), .B1(n15392), .B2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15394) );
  AOI22_X1 U18574 ( .A1(n15395), .A2(n15425), .B1(n15399), .B2(n15394), .ZN(
        n16197) );
  OAI222_X1 U18575 ( .A1(n15408), .A2(n15407), .B1(n15543), .B2(n16197), .C1(
        n16244), .C2(n19146), .ZN(n15396) );
  MUX2_X1 U18576 ( .A(n15396), .B(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .S(
        n15542), .Z(P2_U3600) );
  NAND2_X1 U18577 ( .A1(n15398), .A2(n15397), .ZN(n15415) );
  NAND2_X1 U18578 ( .A1(n15399), .A2(n16194), .ZN(n15417) );
  AND2_X1 U18579 ( .A1(n15414), .A2(n15417), .ZN(n15400) );
  NAND2_X1 U18580 ( .A1(n15415), .A2(n15400), .ZN(n15405) );
  OR2_X1 U18581 ( .A1(n16213), .A2(n16211), .ZN(n15418) );
  INV_X1 U18582 ( .A(n15400), .ZN(n15403) );
  NOR2_X1 U18583 ( .A1(n15401), .A2(n10271), .ZN(n15402) );
  AOI22_X1 U18584 ( .A1(n15418), .A2(n15403), .B1(n15402), .B2(n15416), .ZN(
        n15404) );
  NAND2_X1 U18585 ( .A1(n15405), .A2(n15404), .ZN(n15406) );
  AOI21_X1 U18586 ( .B1(n9829), .B2(n15425), .A(n15406), .ZN(n16193) );
  INV_X1 U18587 ( .A(n15407), .ZN(n15409) );
  OAI222_X1 U18588 ( .A1(n19147), .A2(n16244), .B1(n16193), .B2(n15543), .C1(
        n15409), .C2(n15408), .ZN(n15410) );
  MUX2_X1 U18589 ( .A(n15410), .B(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(
        n15542), .Z(P2_U3599) );
  NAND2_X1 U18590 ( .A1(n15416), .A2(n15411), .ZN(n15412) );
  NAND2_X1 U18591 ( .A1(n15412), .A2(n15417), .ZN(n15413) );
  AOI21_X1 U18592 ( .B1(n15415), .B2(n15414), .A(n15413), .ZN(n15420) );
  AOI22_X1 U18593 ( .A1(n15418), .A2(n15417), .B1(n10271), .B2(n15416), .ZN(
        n15419) );
  MUX2_X1 U18594 ( .A(n15420), .B(n15419), .S(n10330), .Z(n15423) );
  INV_X1 U18595 ( .A(n15421), .ZN(n15422) );
  NAND2_X1 U18596 ( .A1(n15423), .A2(n15422), .ZN(n15424) );
  AOI21_X1 U18597 ( .B1(n13480), .B2(n15425), .A(n15424), .ZN(n16201) );
  OAI22_X1 U18598 ( .A1(n19788), .A2(n16244), .B1(n16201), .B2(n15543), .ZN(
        n15426) );
  MUX2_X1 U18599 ( .A(n15426), .B(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n15542), .Z(P2_U3596) );
  INV_X1 U18600 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n16813) );
  INV_X1 U18601 ( .A(P3_EBX_REG_22__SCAN_IN), .ZN(n16812) );
  INV_X1 U18602 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n16556) );
  INV_X1 U18603 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n16945) );
  INV_X1 U18604 ( .A(n18552), .ZN(n15428) );
  INV_X1 U18605 ( .A(n17146), .ZN(n17149) );
  NAND2_X1 U18606 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n17131) );
  NAND4_X1 U18607 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(P3_EBX_REG_11__SCAN_IN), 
        .A3(P3_EBX_REG_10__SCAN_IN), .A4(P3_EBX_REG_9__SCAN_IN), .ZN(n15432)
         );
  INV_X1 U18608 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n16603) );
  NAND4_X1 U18609 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(P3_EBX_REG_15__SCAN_IN), 
        .A3(P3_EBX_REG_14__SCAN_IN), .A4(P3_EBX_REG_13__SCAN_IN), .ZN(n16950)
         );
  NOR2_X1 U18610 ( .A1(n16603), .A2(n16950), .ZN(n16946) );
  NAND2_X1 U18611 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16915), .ZN(n16903) );
  NAND2_X1 U18612 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n16859), .ZN(n15512) );
  NAND2_X1 U18613 ( .A1(n17291), .A2(n17146), .ZN(n16963) );
  NOR2_X1 U18614 ( .A1(n17150), .A2(n16848), .ZN(n16849) );
  OAI22_X1 U18615 ( .A1(n11799), .A2(n15433), .B1(n9848), .B2(n16894), .ZN(
        n15443) );
  AOI22_X1 U18616 ( .A1(n17054), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17049), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n15441) );
  AOI22_X1 U18617 ( .A1(n17095), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17083), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n15440) );
  AOI22_X1 U18618 ( .A1(n17089), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17110), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n15434) );
  OAI21_X1 U18619 ( .B1(n17027), .B2(n15516), .A(n15434), .ZN(n15438) );
  AOI22_X1 U18620 ( .A1(n17036), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n15497), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n15436) );
  AOI22_X1 U18621 ( .A1(n17002), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17070), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n15435) );
  OAI211_X1 U18622 ( .C1(n16933), .C2(n15514), .A(n15436), .B(n15435), .ZN(
        n15437) );
  AOI211_X1 U18623 ( .C1(n16967), .C2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A(
        n15438), .B(n15437), .ZN(n15439) );
  NAND3_X1 U18624 ( .A1(n15441), .A2(n15440), .A3(n15439), .ZN(n15442) );
  AOI211_X1 U18625 ( .C1(n17103), .C2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A(
        n15443), .B(n15442), .ZN(n15510) );
  AOI22_X1 U18626 ( .A1(n17076), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n15497), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n15444) );
  OAI21_X1 U18627 ( .B1(n15492), .B2(n17034), .A(n15444), .ZN(n15454) );
  AOI22_X1 U18628 ( .A1(n17101), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17103), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n15452) );
  AOI22_X1 U18629 ( .A1(n16967), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17102), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n15445) );
  OAI21_X1 U18630 ( .B1(n17027), .B2(n15446), .A(n15445), .ZN(n15450) );
  INV_X1 U18631 ( .A(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n18443) );
  AOI22_X1 U18632 ( .A1(n15498), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n17049), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n15448) );
  AOI22_X1 U18633 ( .A1(n17002), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17083), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n15447) );
  OAI211_X1 U18634 ( .C1(n16987), .C2(n18443), .A(n15448), .B(n15447), .ZN(
        n15449) );
  AOI211_X1 U18635 ( .C1(n17077), .C2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A(
        n15450), .B(n15449), .ZN(n15451) );
  OAI211_X1 U18636 ( .C1(n11799), .C2(n18342), .A(n15452), .B(n15451), .ZN(
        n15453) );
  AOI211_X1 U18637 ( .C1(n17089), .C2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A(
        n15454), .B(n15453), .ZN(n16856) );
  OAI22_X1 U18638 ( .A1(n11799), .A2(n18336), .B1(n17086), .B2(n16933), .ZN(
        n15464) );
  AOI22_X1 U18639 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n17083), .B1(
        P3_INSTQUEUE_REG_15__1__SCAN_IN), .B2(n15497), .ZN(n15462) );
  AOI22_X1 U18640 ( .A1(n17089), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n17095), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n15461) );
  AOI22_X1 U18641 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n17101), .B1(
        P3_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n17049), .ZN(n15455) );
  OAI21_X1 U18642 ( .B1(n17027), .B2(n16955), .A(n15455), .ZN(n15459) );
  AOI22_X1 U18643 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n17102), .B1(
        n17070), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n15457) );
  AOI22_X1 U18644 ( .A1(n17002), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_12__1__SCAN_IN), .B2(n17076), .ZN(n15456) );
  OAI211_X1 U18645 ( .C1(n11811), .C2(n17073), .A(n15457), .B(n15456), .ZN(
        n15458) );
  AOI211_X1 U18646 ( .C1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .C2(n17110), .A(
        n15459), .B(n15458), .ZN(n15460) );
  NAND3_X1 U18647 ( .A1(n15462), .A2(n15461), .A3(n15460), .ZN(n15463) );
  AOI211_X1 U18648 ( .C1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .C2(n17103), .A(
        n15464), .B(n15463), .ZN(n16865) );
  AOI22_X1 U18649 ( .A1(n17002), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17102), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n15474) );
  AOI22_X1 U18650 ( .A1(n17103), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n15497), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n15465) );
  OAI21_X1 U18651 ( .B1(n9847), .B2(n16969), .A(n15465), .ZN(n15472) );
  AOI22_X1 U18652 ( .A1(n17092), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17049), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n15470) );
  AOI22_X1 U18653 ( .A1(n17089), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17070), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n15467) );
  AOI22_X1 U18654 ( .A1(n17095), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17093), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n15466) );
  OAI211_X1 U18655 ( .C1(n16933), .C2(n16965), .A(n15467), .B(n15466), .ZN(
        n15468) );
  AOI21_X1 U18656 ( .B1(n16967), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A(
        n15468), .ZN(n15469) );
  OAI211_X1 U18657 ( .C1(n16987), .C2(n21054), .A(n15470), .B(n15469), .ZN(
        n15471) );
  AOI211_X1 U18658 ( .C1(n17054), .C2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A(
        n15472), .B(n15471), .ZN(n15473) );
  OAI211_X1 U18659 ( .C1(n11799), .C2(n18333), .A(n15474), .B(n15473), .ZN(
        n16871) );
  AOI22_X1 U18660 ( .A1(n15498), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n16967), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n15485) );
  AOI22_X1 U18661 ( .A1(n17036), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17049), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n15476) );
  AOI22_X1 U18662 ( .A1(n17083), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17093), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n15475) );
  OAI211_X1 U18663 ( .C1(n16933), .C2(n15477), .A(n15476), .B(n15475), .ZN(
        n15483) );
  AOI22_X1 U18664 ( .A1(n17089), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17103), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n15481) );
  AOI22_X1 U18665 ( .A1(n17002), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n17095), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n15480) );
  AOI22_X1 U18666 ( .A1(n17054), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n15497), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n15479) );
  NAND2_X1 U18667 ( .A1(n17074), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n15478) );
  NAND4_X1 U18668 ( .A1(n15481), .A2(n15480), .A3(n15479), .A4(n15478), .ZN(
        n15482) );
  AOI211_X1 U18669 ( .C1(n17110), .C2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A(
        n15483), .B(n15482), .ZN(n15484) );
  OAI211_X1 U18670 ( .C1(n17027), .C2(n16991), .A(n15485), .B(n15484), .ZN(
        n16872) );
  NAND2_X1 U18671 ( .A1(n16871), .A2(n16872), .ZN(n16870) );
  NOR2_X1 U18672 ( .A1(n16865), .A2(n16870), .ZN(n16864) );
  AOI22_X1 U18673 ( .A1(n17036), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17093), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n15496) );
  INV_X1 U18674 ( .A(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n21070) );
  AOI22_X1 U18675 ( .A1(n15498), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n15497), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n15486) );
  OAI21_X1 U18676 ( .B1(n16983), .B2(n21070), .A(n15486), .ZN(n15494) );
  AOI22_X1 U18677 ( .A1(n16967), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17074), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n15491) );
  INV_X1 U18678 ( .A(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n18439) );
  AOI22_X1 U18679 ( .A1(n17089), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17002), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n15488) );
  AOI22_X1 U18680 ( .A1(n17103), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17049), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n15487) );
  OAI211_X1 U18681 ( .C1(n16987), .C2(n18439), .A(n15488), .B(n15487), .ZN(
        n15489) );
  AOI21_X1 U18682 ( .B1(n17077), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A(
        n15489), .ZN(n15490) );
  OAI211_X1 U18683 ( .C1(n15492), .C2(n16934), .A(n15491), .B(n15490), .ZN(
        n15493) );
  AOI211_X1 U18684 ( .C1(n17083), .C2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A(
        n15494), .B(n15493), .ZN(n15495) );
  OAI211_X1 U18685 ( .C1(n17027), .C2(n17062), .A(n15496), .B(n15495), .ZN(
        n16861) );
  NAND2_X1 U18686 ( .A1(n16864), .A2(n16861), .ZN(n16860) );
  NOR2_X1 U18687 ( .A1(n16856), .A2(n16860), .ZN(n16855) );
  AOI22_X1 U18688 ( .A1(n17002), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n15497), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n15508) );
  AOI22_X1 U18689 ( .A1(n15498), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n17049), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n15500) );
  AOI22_X1 U18690 ( .A1(n17089), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17083), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n15499) );
  OAI211_X1 U18691 ( .C1(n16987), .C2(n20935), .A(n15500), .B(n15499), .ZN(
        n15506) );
  AOI22_X1 U18692 ( .A1(n17101), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17093), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n15504) );
  AOI22_X1 U18693 ( .A1(n17095), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17103), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n15503) );
  AOI22_X1 U18694 ( .A1(n17092), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17102), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n15502) );
  NAND2_X1 U18695 ( .A1(n16967), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n15501) );
  NAND4_X1 U18696 ( .A1(n15504), .A2(n15503), .A3(n15502), .A4(n15501), .ZN(
        n15505) );
  AOI211_X1 U18697 ( .C1(n17077), .C2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A(
        n15506), .B(n15505), .ZN(n15507) );
  OAI211_X1 U18698 ( .C1(n11799), .C2(n15509), .A(n15508), .B(n15507), .ZN(
        n16852) );
  NAND2_X1 U18699 ( .A1(n16855), .A2(n16852), .ZN(n16851) );
  NOR2_X1 U18700 ( .A1(n15510), .A2(n16851), .ZN(n16846) );
  AOI21_X1 U18701 ( .B1(n15510), .B2(n16851), .A(n16846), .ZN(n17168) );
  AOI22_X1 U18702 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16849), .B1(n17168), 
        .B2(n17150), .ZN(n15511) );
  OAI21_X1 U18703 ( .B1(P3_EBX_REG_28__SCAN_IN), .B2(n15512), .A(n15511), .ZN(
        P3_U2675) );
  AOI22_X1 U18704 ( .A1(n17049), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17093), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n15513) );
  OAI21_X1 U18705 ( .B1(n16983), .B2(n15514), .A(n15513), .ZN(n15525) );
  AOI22_X1 U18706 ( .A1(n17095), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17083), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n15523) );
  AOI22_X1 U18707 ( .A1(n17074), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17110), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n15515) );
  OAI21_X1 U18708 ( .B1(n10222), .B2(n15516), .A(n15515), .ZN(n15521) );
  AOI22_X1 U18709 ( .A1(n17002), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17070), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n15518) );
  AOI22_X1 U18710 ( .A1(n17102), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17100), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n15517) );
  OAI211_X1 U18711 ( .C1(n16933), .C2(n15519), .A(n15518), .B(n15517), .ZN(
        n15520) );
  AOI211_X1 U18712 ( .C1(n16967), .C2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A(
        n15521), .B(n15520), .ZN(n15522) );
  OAI211_X1 U18713 ( .C1(n17027), .C2(n21003), .A(n15523), .B(n15522), .ZN(
        n15524) );
  AOI211_X1 U18714 ( .C1(n17089), .C2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A(
        n15525), .B(n15524), .ZN(n17249) );
  NOR2_X1 U18715 ( .A1(n17150), .A2(n17001), .ZN(n17030) );
  INV_X1 U18716 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n16648) );
  OAI222_X1 U18717 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n18145), .B1(
        P3_EBX_REG_13__SCAN_IN), .B2(n17001), .C1(n17030), .C2(n16648), .ZN(
        n15526) );
  OAI21_X1 U18718 ( .B1(n17249), .B2(n17141), .A(n15526), .ZN(P3_U2690) );
  NAND2_X1 U18719 ( .A1(READY22_REG_SCAN_IN), .A2(READY2), .ZN(n18768) );
  NAND2_X1 U18720 ( .A1(n18555), .A2(n18768), .ZN(n15538) );
  INV_X2 U18721 ( .A(n18773), .ZN(n18772) );
  NAND2_X2 U18722 ( .A1(n18772), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n18707) );
  OAI211_X1 U18723 ( .C1(P3_STATE_REG_1__SCAN_IN), .C2(P3_STATE_REG_2__SCAN_IN), .A(n18642), .B(n18707), .ZN(n18758) );
  INV_X1 U18724 ( .A(n15530), .ZN(n18564) );
  OAI21_X1 U18725 ( .B1(n15533), .B2(n15532), .A(n15531), .ZN(n15535) );
  NAND2_X1 U18726 ( .A1(n15535), .A2(n15534), .ZN(n15549) );
  NOR3_X1 U18727 ( .A1(n15637), .A2(n15536), .A3(n15549), .ZN(n15537) );
  NOR2_X1 U18728 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18716), .ZN(n18113) );
  INV_X1 U18729 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n18101) );
  NOR2_X1 U18730 ( .A1(n18101), .A2(n18714), .ZN(n15539) );
  INV_X1 U18731 ( .A(n18746), .ZN(n18743) );
  AOI21_X1 U18732 ( .B1(n15540), .B2(n18561), .A(n16432), .ZN(n18608) );
  NAND3_X1 U18733 ( .A1(n18743), .A2(n18776), .A3(n18608), .ZN(n15541) );
  OAI21_X1 U18734 ( .B1(n18743), .B2(n18561), .A(n15541), .ZN(P3_U3284) );
  INV_X1 U18735 ( .A(n15542), .ZN(n15548) );
  NOR4_X1 U18736 ( .A1(n15544), .A2(n16224), .A3(n9779), .A4(n15543), .ZN(
        n15545) );
  NAND2_X1 U18737 ( .A1(n15548), .A2(n15545), .ZN(n15546) );
  OAI21_X1 U18738 ( .B1(n15548), .B2(n15547), .A(n15546), .ZN(P2_U3595) );
  INV_X1 U18739 ( .A(n15552), .ZN(n18121) );
  OAI21_X1 U18740 ( .B1(n18121), .B2(n18760), .A(n18758), .ZN(n15553) );
  OAI21_X1 U18741 ( .B1(n15554), .B2(n15553), .A(n18768), .ZN(n16415) );
  OAI22_X1 U18742 ( .A1(n15557), .A2(n15556), .B1(n15555), .B2(n16415), .ZN(
        n15558) );
  NAND2_X1 U18743 ( .A1(n15558), .A2(n18555), .ZN(n15559) );
  NAND2_X1 U18744 ( .A1(n15566), .A2(n18089), .ZN(n18095) );
  NOR2_X1 U18745 ( .A1(n15567), .A2(n18095), .ZN(n18017) );
  INV_X1 U18746 ( .A(n16260), .ZN(n16276) );
  NAND2_X1 U18747 ( .A1(n17791), .A2(n15623), .ZN(n16259) );
  AOI22_X1 U18748 ( .A1(n18017), .A2(n16276), .B1(n18082), .B2(n16259), .ZN(
        n15627) );
  INV_X1 U18749 ( .A(n18008), .ZN(n18010) );
  NAND2_X1 U18750 ( .A1(n18010), .A2(n18089), .ZN(n18078) );
  INV_X1 U18751 ( .A(n18078), .ZN(n16291) );
  INV_X1 U18752 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17477) );
  NOR2_X1 U18753 ( .A1(n17477), .A2(n17832), .ZN(n17787) );
  AOI21_X1 U18754 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18005) );
  INV_X1 U18755 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n18054) );
  NOR3_X1 U18756 ( .A1(n10013), .A2(n18054), .A3(n18004), .ZN(n18007) );
  NAND4_X1 U18757 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A4(n18007), .ZN(n17933) );
  NOR2_X1 U18758 ( .A1(n18005), .A2(n17933), .ZN(n17950) );
  NAND2_X1 U18759 ( .A1(n15568), .A2(n17950), .ZN(n17848) );
  OAI21_X1 U18760 ( .B1(n17854), .B2(n17848), .A(n18567), .ZN(n17833) );
  OAI21_X1 U18761 ( .B1(n17787), .B2(n18582), .A(n17833), .ZN(n17809) );
  AOI21_X1 U18762 ( .B1(n18567), .B2(n17788), .A(n17809), .ZN(n17790) );
  OAI21_X1 U18763 ( .B1(n18742), .B2(n17800), .A(n18587), .ZN(n15562) );
  NAND2_X1 U18764 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18006) );
  NOR2_X1 U18765 ( .A1(n17933), .A2(n18006), .ZN(n17908) );
  NAND2_X1 U18766 ( .A1(n15568), .A2(n17908), .ZN(n17887) );
  NOR2_X1 U18767 ( .A1(n17847), .A2(n18587), .ZN(n17892) );
  INV_X1 U18768 ( .A(n17892), .ZN(n18068) );
  OAI21_X1 U18769 ( .B1(n16254), .B2(n17887), .A(n18068), .ZN(n15561) );
  NAND4_X1 U18770 ( .A1(n17790), .A2(n18046), .A3(n15562), .A4(n15561), .ZN(
        n15626) );
  AOI21_X1 U18771 ( .B1(n17984), .B2(n17800), .A(n15626), .ZN(n15563) );
  INV_X1 U18772 ( .A(n15563), .ZN(n16302) );
  AOI22_X1 U18773 ( .A1(n16291), .A2(n16298), .B1(n18091), .B2(n16302), .ZN(
        n15572) );
  NAND3_X1 U18774 ( .A1(n15567), .A2(n18089), .A3(n15566), .ZN(n17992) );
  NAND2_X1 U18775 ( .A1(n17694), .A2(n16298), .ZN(n16310) );
  OAI21_X1 U18776 ( .B1(n15564), .B2(n16299), .A(n16310), .ZN(n15565) );
  XOR2_X1 U18777 ( .A(n15565), .B(n16272), .Z(n16274) );
  INV_X1 U18778 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n18701) );
  NOR2_X1 U18779 ( .A1(n18091), .A2(n18701), .ZN(n16267) );
  INV_X1 U18780 ( .A(n16270), .ZN(n16275) );
  INV_X1 U18781 ( .A(n17951), .ZN(n17692) );
  INV_X1 U18782 ( .A(n15566), .ZN(n18557) );
  NOR2_X1 U18783 ( .A1(n18557), .A2(n15567), .ZN(n17850) );
  INV_X1 U18784 ( .A(n17850), .ZN(n17954) );
  OAI22_X1 U18785 ( .A1(n17974), .A2(n18072), .B1(n17692), .B2(n17954), .ZN(
        n17894) );
  AOI21_X1 U18786 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n18587), .A(
        n17847), .ZN(n18064) );
  OAI22_X1 U18787 ( .A1(n18582), .A2(n17848), .B1(n18064), .B2(n17887), .ZN(
        n17813) );
  AOI21_X1 U18788 ( .B1(n15568), .B2(n17894), .A(n17813), .ZN(n17846) );
  NAND2_X1 U18789 ( .A1(n15569), .A2(n17872), .ZN(n17794) );
  NOR3_X1 U18790 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n16275), .A3(
        n17794), .ZN(n15570) );
  AOI211_X1 U18791 ( .C1(n18015), .C2(n16274), .A(n16267), .B(n15570), .ZN(
        n15571) );
  OAI221_X1 U18792 ( .B1(n16272), .B2(n15627), .C1(n16272), .C2(n15572), .A(
        n15571), .ZN(P3_U2833) );
  OAI22_X1 U18793 ( .A1(n15573), .A2(n18994), .B1(n12191), .B2(n18973), .ZN(
        n15574) );
  INV_X1 U18794 ( .A(n15574), .ZN(n15582) );
  AOI22_X1 U18795 ( .A1(P2_EBX_REG_22__SCAN_IN), .A2(n18990), .B1(
        P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n18964), .ZN(n15581) );
  INV_X1 U18796 ( .A(n16034), .ZN(n15575) );
  OAI22_X1 U18797 ( .A1(n16054), .A2(n18981), .B1(n18982), .B2(n15575), .ZN(
        n15576) );
  INV_X1 U18798 ( .A(n15576), .ZN(n15580) );
  OAI211_X1 U18799 ( .C1(n16061), .C2(n15578), .A(n18999), .B(n15577), .ZN(
        n15579) );
  NAND4_X1 U18800 ( .A1(n15582), .A2(n15581), .A3(n15580), .A4(n15579), .ZN(
        P2_U2833) );
  INV_X1 U18801 ( .A(n15595), .ZN(n15597) );
  INV_X1 U18802 ( .A(n15583), .ZN(n15584) );
  OAI211_X1 U18803 ( .C1(n11132), .C2(n15585), .A(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n15584), .ZN(n15588) );
  INV_X1 U18804 ( .A(n15586), .ZN(n15587) );
  OAI21_X1 U18805 ( .B1(n20622), .B2(n15588), .A(n15587), .ZN(n15590) );
  NAND2_X1 U18806 ( .A1(n20622), .A2(n15588), .ZN(n15589) );
  OAI21_X1 U18807 ( .B1(n15591), .B2(n15590), .A(n15589), .ZN(n15594) );
  AND2_X1 U18808 ( .A1(n20367), .A2(n15594), .ZN(n15593) );
  OAI222_X1 U18809 ( .A1(n20773), .A2(n15595), .B1(n20367), .B2(n15594), .C1(
        n15593), .C2(n15592), .ZN(n15596) );
  OAI21_X1 U18810 ( .B1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n15597), .A(
        n15596), .ZN(n15607) );
  NOR2_X1 U18811 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(P1_MORE_REG_SCAN_IN), .ZN(
        n15604) );
  INV_X1 U18812 ( .A(n15598), .ZN(n15600) );
  AND2_X1 U18813 ( .A1(n15600), .A2(n15599), .ZN(n15601) );
  OAI211_X1 U18814 ( .C1(n15604), .C2(n15603), .A(n15602), .B(n15601), .ZN(
        n15605) );
  AOI211_X1 U18815 ( .C1(n15607), .C2(n20869), .A(n15606), .B(n15605), .ZN(
        n15622) );
  INV_X1 U18816 ( .A(n15622), .ZN(n15612) );
  INV_X1 U18817 ( .A(n15608), .ZN(n15610) );
  NAND3_X1 U18818 ( .A1(n15610), .A2(n15609), .A3(n20574), .ZN(n15611) );
  NOR2_X1 U18819 ( .A1(n15937), .A2(n15630), .ZN(n20787) );
  INV_X1 U18820 ( .A(n20787), .ZN(n15929) );
  OAI211_X1 U18821 ( .C1(n20687), .C2(n20788), .A(n15611), .B(n15929), .ZN(
        n15932) );
  AOI221_X1 U18822 ( .B1(n20098), .B2(n15937), .C1(n15612), .C2(n15937), .A(
        n15932), .ZN(n15938) );
  NOR2_X1 U18823 ( .A1(n15613), .A2(n15935), .ZN(n15614) );
  NOR2_X1 U18824 ( .A1(n15938), .A2(n15614), .ZN(n15620) );
  AOI21_X1 U18825 ( .B1(n15615), .B2(n20697), .A(P1_STATE2_REG_2__SCAN_IN), 
        .ZN(n15616) );
  NOR2_X1 U18826 ( .A1(n15617), .A2(n15616), .ZN(n15618) );
  NAND2_X1 U18827 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n15618), .ZN(n15619) );
  OAI22_X1 U18828 ( .A1(n15620), .A2(P1_STATE2_REG_0__SCAN_IN), .B1(n15938), 
        .B2(n15619), .ZN(n15621) );
  OAI21_X1 U18829 ( .B1(n15622), .B2(n19861), .A(n15621), .ZN(P1_U3161) );
  NAND2_X1 U18830 ( .A1(n15623), .A2(n20896), .ZN(n16265) );
  AOI21_X1 U18831 ( .B1(n15625), .B2(n20896), .A(n15624), .ZN(n16261) );
  AOI22_X1 U18832 ( .A1(n16291), .A2(n16284), .B1(n18091), .B2(n15626), .ZN(
        n16287) );
  AOI21_X1 U18833 ( .B1(n16287), .B2(n15627), .A(n20896), .ZN(n15628) );
  AOI21_X1 U18834 ( .B1(n18015), .B2(n16261), .A(n15628), .ZN(n15629) );
  INV_X2 U18835 ( .A(n18091), .ZN(n18093) );
  NAND2_X1 U18836 ( .A1(n18093), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n16255) );
  OAI211_X1 U18837 ( .C1(n17794), .C2(n16265), .A(n15629), .B(n16255), .ZN(
        P3_U2832) );
  INV_X1 U18838 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n19858) );
  INV_X1 U18839 ( .A(HOLD), .ZN(n20703) );
  NOR2_X1 U18840 ( .A1(n19858), .A2(n20703), .ZN(n20692) );
  AOI22_X1 U18841 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(HOLD), .B1(
        P1_STATE_REG_0__SCAN_IN), .B2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n15632) );
  NAND2_X1 U18842 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n15630), .ZN(n20695) );
  OAI211_X1 U18843 ( .C1(n20692), .C2(n15632), .A(n15631), .B(n20695), .ZN(
        P1_U3195) );
  INV_X1 U18844 ( .A(n19993), .ZN(n15633) );
  INV_X1 U18845 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n16406) );
  NOR2_X1 U18846 ( .A1(n15633), .A2(n16406), .ZN(P1_U2905) );
  NOR2_X1 U18847 ( .A1(n19844), .A2(n19836), .ZN(n19701) );
  OAI221_X1 U18848 ( .B1(n19701), .B2(P2_STATEBS16_REG_SCAN_IN), .C1(n19701), 
        .C2(n19836), .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n15634) );
  AOI21_X1 U18849 ( .B1(n19149), .B2(n15634), .A(n16248), .ZN(P2_U3178) );
  OAI221_X1 U18850 ( .B1(n21000), .B2(n16252), .C1(n16249), .C2(n16252), .A(
        n19268), .ZN(n19822) );
  NOR2_X1 U18851 ( .A1(n21060), .A2(n19822), .ZN(P2_U3047) );
  INV_X1 U18852 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n17379) );
  OR2_X1 U18853 ( .A1(n17291), .A2(n17155), .ZN(n17199) );
  AOI22_X1 U18854 ( .A1(n17301), .A2(BUF2_REG_0__SCAN_IN), .B1(n17300), .B2(
        n15640), .ZN(n15641) );
  OAI221_X1 U18855 ( .B1(n17304), .B2(n17379), .C1(n17304), .C2(n17199), .A(
        n15641), .ZN(P3_U2735) );
  AND2_X1 U18856 ( .A1(n15642), .A2(n19950), .ZN(n15648) );
  INV_X1 U18857 ( .A(n15643), .ZN(n15646) );
  INV_X1 U18858 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n15645) );
  OAI22_X1 U18859 ( .A1(n15646), .A2(n15645), .B1(n15644), .B2(n19899), .ZN(
        n15647) );
  AOI21_X1 U18860 ( .B1(n15655), .B2(n15648), .A(n15647), .ZN(n15652) );
  NAND2_X1 U18861 ( .A1(n15668), .A2(n15654), .ZN(n15657) );
  INV_X1 U18862 ( .A(n15655), .ZN(n15656) );
  NAND2_X1 U18863 ( .A1(n15657), .A2(n15656), .ZN(n15660) );
  NAND2_X1 U18864 ( .A1(n19937), .A2(P1_EBX_REG_27__SCAN_IN), .ZN(n15659) );
  AOI22_X1 U18865 ( .A1(n19940), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .B1(
        n19895), .B2(P1_REIP_REG_27__SCAN_IN), .ZN(n15658) );
  OAI211_X1 U18866 ( .C1(n15660), .C2(n19926), .A(n15659), .B(n15658), .ZN(
        n15661) );
  INV_X1 U18867 ( .A(n15661), .ZN(n15666) );
  INV_X1 U18868 ( .A(n15662), .ZN(n15663) );
  AOI22_X1 U18869 ( .A1(n15664), .A2(n19912), .B1(n15663), .B2(n19948), .ZN(
        n15665) );
  OAI211_X1 U18870 ( .C1(n15667), .C2(n19957), .A(n15666), .B(n15665), .ZN(
        P1_U2813) );
  AOI22_X1 U18871 ( .A1(n19937), .A2(P1_EBX_REG_26__SCAN_IN), .B1(
        P1_REIP_REG_26__SCAN_IN), .B2(n19895), .ZN(n15671) );
  OAI211_X1 U18872 ( .C1(P1_REIP_REG_26__SCAN_IN), .C2(n15669), .A(n19950), 
        .B(n15668), .ZN(n15670) );
  OAI211_X1 U18873 ( .C1(n15730), .C2(n15672), .A(n15671), .B(n15670), .ZN(
        n15677) );
  INV_X1 U18874 ( .A(n15673), .ZN(n15674) );
  OAI22_X1 U18875 ( .A1(n15675), .A2(n15726), .B1(n15674), .B2(n19897), .ZN(
        n15676) );
  AOI211_X1 U18876 ( .C1(n15678), .C2(n19891), .A(n15677), .B(n15676), .ZN(
        n15679) );
  INV_X1 U18877 ( .A(n15679), .ZN(P1_U2814) );
  AOI22_X1 U18878 ( .A1(n19937), .A2(P1_EBX_REG_23__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n19940), .ZN(n15687) );
  AOI21_X1 U18879 ( .B1(P1_REIP_REG_22__SCAN_IN), .B2(n15680), .A(
        P1_REIP_REG_23__SCAN_IN), .ZN(n15682) );
  OAI22_X1 U18880 ( .A1(n15683), .A2(n19897), .B1(n15682), .B2(n15681), .ZN(
        n15684) );
  AOI21_X1 U18881 ( .B1(n15685), .B2(n19912), .A(n15684), .ZN(n15686) );
  OAI211_X1 U18882 ( .C1(n15688), .C2(n19957), .A(n15687), .B(n15686), .ZN(
        P1_U2817) );
  NOR3_X1 U18883 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(n19926), .A3(n15689), 
        .ZN(n15691) );
  INV_X1 U18884 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n15742) );
  OAI22_X1 U18885 ( .A1(n15696), .A2(n14372), .B1(n15742), .B2(n19899), .ZN(
        n15690) );
  AOI211_X1 U18886 ( .C1(n19940), .C2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n15691), .B(n15690), .ZN(n15694) );
  OAI22_X1 U18887 ( .A1(n15739), .A2(n15726), .B1(n15738), .B2(n19897), .ZN(
        n15692) );
  INV_X1 U18888 ( .A(n15692), .ZN(n15693) );
  OAI211_X1 U18889 ( .C1(n15695), .C2(n19957), .A(n15694), .B(n15693), .ZN(
        P1_U2819) );
  AOI21_X1 U18890 ( .B1(n15698), .B2(n15697), .A(n15696), .ZN(n15699) );
  AOI21_X1 U18891 ( .B1(n19937), .B2(P1_EBX_REG_20__SCAN_IN), .A(n15699), .ZN(
        n15705) );
  OAI22_X1 U18892 ( .A1(n15701), .A2(n15726), .B1(n15700), .B2(n19897), .ZN(
        n15702) );
  AOI21_X1 U18893 ( .B1(n15703), .B2(n19891), .A(n15702), .ZN(n15704) );
  OAI211_X1 U18894 ( .C1(n15706), .C2(n15730), .A(n15705), .B(n15704), .ZN(
        P1_U2820) );
  NAND2_X1 U18895 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(P1_REIP_REG_18__SCAN_IN), 
        .ZN(n15707) );
  OAI21_X1 U18896 ( .B1(P1_REIP_REG_19__SCAN_IN), .B2(P1_REIP_REG_18__SCAN_IN), 
        .A(n15707), .ZN(n15710) );
  AOI22_X1 U18897 ( .A1(n15708), .A2(P1_REIP_REG_19__SCAN_IN), .B1(n19937), 
        .B2(P1_EBX_REG_19__SCAN_IN), .ZN(n15709) );
  OAI21_X1 U18898 ( .B1(n15711), .B2(n15710), .A(n15709), .ZN(n15712) );
  AOI211_X1 U18899 ( .C1(n19940), .C2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n19909), .B(n15712), .ZN(n15715) );
  INV_X1 U18900 ( .A(n15713), .ZN(n15809) );
  AOI22_X1 U18901 ( .A1(n15750), .A2(n19912), .B1(n15809), .B2(n19948), .ZN(
        n15714) );
  OAI211_X1 U18902 ( .C1(n15753), .C2(n19957), .A(n15715), .B(n15714), .ZN(
        P1_U2821) );
  INV_X1 U18903 ( .A(n15862), .ZN(n15716) );
  NAND2_X1 U18904 ( .A1(n19948), .A2(n15716), .ZN(n15719) );
  NAND2_X1 U18905 ( .A1(n19937), .A2(P1_EBX_REG_12__SCAN_IN), .ZN(n15718) );
  NAND2_X1 U18906 ( .A1(n19940), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15717) );
  AND4_X1 U18907 ( .A1(n15719), .A2(n15718), .A3(n19942), .A4(n15717), .ZN(
        n15725) );
  INV_X1 U18908 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n20958) );
  NAND2_X1 U18909 ( .A1(n19950), .A2(n15720), .ZN(n15728) );
  INV_X1 U18910 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n15721) );
  OAI21_X1 U18911 ( .B1(n20958), .B2(n15728), .A(n15721), .ZN(n15722) );
  AOI22_X1 U18912 ( .A1(n15770), .A2(n19891), .B1(n15723), .B2(n15722), .ZN(
        n15724) );
  OAI211_X1 U18913 ( .C1(n15726), .C2(n15769), .A(n15725), .B(n15724), .ZN(
        P1_U2828) );
  INV_X1 U18914 ( .A(n15863), .ZN(n15727) );
  OAI22_X1 U18915 ( .A1(n15728), .A2(P1_REIP_REG_11__SCAN_IN), .B1(n19897), 
        .B2(n15727), .ZN(n15735) );
  NOR2_X1 U18916 ( .A1(n15730), .A2(n15729), .ZN(n15731) );
  AOI211_X1 U18917 ( .C1(n15732), .C2(P1_REIP_REG_11__SCAN_IN), .A(n19909), 
        .B(n15731), .ZN(n15733) );
  OAI21_X1 U18918 ( .B1(n21031), .B2(n19899), .A(n15733), .ZN(n15734) );
  AOI211_X1 U18919 ( .C1(n19912), .C2(n15777), .A(n15735), .B(n15734), .ZN(
        n15736) );
  OAI21_X1 U18920 ( .B1(n15780), .B2(n19957), .A(n15736), .ZN(P1_U2829) );
  OAI22_X1 U18921 ( .A1(n15739), .A2(n14213), .B1(n15738), .B2(n15737), .ZN(
        n15740) );
  INV_X1 U18922 ( .A(n15740), .ZN(n15741) );
  OAI21_X1 U18923 ( .B1(n19966), .B2(n15742), .A(n15741), .ZN(P1_U2851) );
  AOI22_X1 U18924 ( .A1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n20043), .B1(
        n11744), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n15752) );
  INV_X1 U18925 ( .A(n15743), .ZN(n15749) );
  NAND2_X1 U18926 ( .A1(n15747), .A2(n15744), .ZN(n15746) );
  MUX2_X1 U18927 ( .A(n15747), .B(n15746), .S(n15745), .Z(n15748) );
  NAND2_X1 U18928 ( .A1(n15749), .A2(n15748), .ZN(n15810) );
  AOI22_X1 U18929 ( .A1(n15810), .A2(n20046), .B1(n20038), .B2(n15750), .ZN(
        n15751) );
  OAI211_X1 U18930 ( .C1(n15753), .C2(n20041), .A(n15752), .B(n15751), .ZN(
        P1_U2980) );
  AOI22_X1 U18931 ( .A1(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n20043), .B1(
        n11744), .B2(P1_REIP_REG_17__SCAN_IN), .ZN(n15758) );
  INV_X1 U18932 ( .A(n15754), .ZN(n15756) );
  AOI22_X1 U18933 ( .A1(n15756), .A2(n20038), .B1(n20045), .B2(n15755), .ZN(
        n15757) );
  OAI211_X1 U18934 ( .C1(n19867), .C2(n15759), .A(n15758), .B(n15757), .ZN(
        P1_U2982) );
  AOI22_X1 U18935 ( .A1(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n20043), .B1(
        n11744), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n15763) );
  AOI22_X1 U18936 ( .A1(n15761), .A2(n20038), .B1(n20045), .B2(n15760), .ZN(
        n15762) );
  OAI211_X1 U18937 ( .C1(n15764), .C2(n19867), .A(n15763), .B(n15762), .ZN(
        P1_U2984) );
  OAI21_X1 U18938 ( .B1(n15767), .B2(n15766), .A(n15765), .ZN(n15768) );
  INV_X1 U18939 ( .A(n15768), .ZN(n15857) );
  AOI22_X1 U18940 ( .A1(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n20043), .B1(
        n11744), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n15773) );
  INV_X1 U18941 ( .A(n15769), .ZN(n15771) );
  AOI22_X1 U18942 ( .A1(n20038), .A2(n15771), .B1(n15770), .B2(n20045), .ZN(
        n15772) );
  OAI211_X1 U18943 ( .C1(n15857), .C2(n19867), .A(n15773), .B(n15772), .ZN(
        P1_U2987) );
  AOI22_X1 U18944 ( .A1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n20043), .B1(
        n11744), .B2(P1_REIP_REG_11__SCAN_IN), .ZN(n15779) );
  NOR2_X1 U18945 ( .A1(n14431), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15775) );
  NOR2_X1 U18946 ( .A1(n14395), .A2(n11648), .ZN(n15774) );
  MUX2_X1 U18947 ( .A(n15775), .B(n15774), .S(n14352), .Z(n15776) );
  XNOR2_X1 U18948 ( .A(n15776), .B(n15868), .ZN(n15865) );
  AOI22_X1 U18949 ( .A1(n20038), .A2(n15777), .B1(n20046), .B2(n15865), .ZN(
        n15778) );
  OAI211_X1 U18950 ( .C1(n15780), .C2(n20041), .A(n15779), .B(n15778), .ZN(
        P1_U2988) );
  AOI22_X1 U18951 ( .A1(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n20043), .B1(
        n11744), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n15786) );
  NAND2_X1 U18952 ( .A1(n15783), .A2(n15782), .ZN(n15784) );
  XNOR2_X1 U18953 ( .A(n15781), .B(n15784), .ZN(n15908) );
  AOI22_X1 U18954 ( .A1(n15908), .A2(n20046), .B1(n20038), .B2(n19906), .ZN(
        n15785) );
  OAI211_X1 U18955 ( .C1(n19904), .C2(n20041), .A(n15786), .B(n15785), .ZN(
        P1_U2992) );
  AOI22_X1 U18956 ( .A1(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n20043), .B1(
        n11744), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n15791) );
  XNOR2_X1 U18957 ( .A(n15788), .B(n15898), .ZN(n15789) );
  XNOR2_X1 U18958 ( .A(n15787), .B(n15789), .ZN(n15914) );
  AOI22_X1 U18959 ( .A1(n15914), .A2(n20046), .B1(n20038), .B2(n19913), .ZN(
        n15790) );
  OAI211_X1 U18960 ( .C1(n19916), .C2(n20041), .A(n15791), .B(n15790), .ZN(
        P1_U2993) );
  AOI22_X1 U18961 ( .A1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n20043), .B1(
        n11744), .B2(P1_REIP_REG_5__SCAN_IN), .ZN(n15797) );
  OAI21_X1 U18962 ( .B1(n15792), .B2(n15794), .A(n15793), .ZN(n15924) );
  INV_X1 U18963 ( .A(n15924), .ZN(n15795) );
  INV_X1 U18964 ( .A(n19932), .ZN(n19963) );
  AOI22_X1 U18965 ( .A1(n15795), .A2(n20046), .B1(n20038), .B2(n19963), .ZN(
        n15796) );
  OAI211_X1 U18966 ( .C1(n19936), .C2(n20041), .A(n15797), .B(n15796), .ZN(
        P1_U2994) );
  AOI22_X1 U18967 ( .A1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n15798), .B1(
        n11744), .B2(P1_REIP_REG_22__SCAN_IN), .ZN(n15806) );
  INV_X1 U18968 ( .A(n15799), .ZN(n15804) );
  INV_X1 U18969 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15801) );
  AOI21_X1 U18970 ( .B1(n15801), .B2(n20949), .A(n15800), .ZN(n15802) );
  AOI22_X1 U18971 ( .A1(n15804), .A2(n20086), .B1(n15803), .B2(n15802), .ZN(
        n15805) );
  OAI211_X1 U18972 ( .C1(n20083), .C2(n15807), .A(n15806), .B(n15805), .ZN(
        P1_U3009) );
  AOI22_X1 U18973 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n15808), .B1(
        n11744), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n15812) );
  AOI22_X1 U18974 ( .A1(n15810), .A2(n20086), .B1(n20063), .B2(n15809), .ZN(
        n15811) );
  OAI211_X1 U18975 ( .C1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n15813), .A(
        n15812), .B(n15811), .ZN(P1_U3012) );
  NOR2_X1 U18976 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n15814), .ZN(
        n15815) );
  AOI22_X1 U18977 ( .A1(n11744), .A2(P1_REIP_REG_18__SCAN_IN), .B1(n15816), 
        .B2(n15815), .ZN(n15821) );
  INV_X1 U18978 ( .A(n15817), .ZN(n15819) );
  AOI22_X1 U18979 ( .A1(n15819), .A2(n20086), .B1(
        P1_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n15818), .ZN(n15820) );
  OAI211_X1 U18980 ( .C1(n20083), .C2(n15822), .A(n15821), .B(n15820), .ZN(
        P1_U3013) );
  INV_X1 U18981 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15824) );
  NOR3_X1 U18982 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n15824), .A3(
        n15823), .ZN(n15827) );
  NOR2_X1 U18983 ( .A1(n15825), .A2(n15923), .ZN(n15826) );
  AOI211_X1 U18984 ( .C1(n11744), .C2(P1_REIP_REG_16__SCAN_IN), .A(n15827), 
        .B(n15826), .ZN(n15831) );
  OAI21_X1 U18985 ( .B1(n15829), .B2(n15828), .A(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15830) );
  OAI211_X1 U18986 ( .C1(n20083), .C2(n15832), .A(n15831), .B(n15830), .ZN(
        P1_U3015) );
  NAND2_X1 U18987 ( .A1(n20071), .A2(n15871), .ZN(n15896) );
  NAND2_X1 U18988 ( .A1(n20053), .A2(n20051), .ZN(n15833) );
  NAND2_X1 U18989 ( .A1(n15896), .A2(n15833), .ZN(n20065) );
  NAND2_X1 U18990 ( .A1(n20065), .A2(n15834), .ZN(n15917) );
  NAND4_X1 U18991 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(n15855), .A4(n15900), .ZN(
        n15836) );
  NAND2_X1 U18992 ( .A1(n11744), .A2(P1_REIP_REG_14__SCAN_IN), .ZN(n15835) );
  OAI221_X1 U18993 ( .B1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n15836), 
        .C1(n14408), .C2(n15848), .A(n15835), .ZN(n15837) );
  AOI21_X1 U18994 ( .B1(n15838), .B2(n20086), .A(n15837), .ZN(n15839) );
  OAI21_X1 U18995 ( .B1(n20083), .B2(n15840), .A(n15839), .ZN(P1_U3017) );
  INV_X1 U18996 ( .A(n15841), .ZN(n15842) );
  AOI22_X1 U18997 ( .A1(P1_REIP_REG_13__SCAN_IN), .A2(n11744), .B1(n15847), 
        .B2(n15842), .ZN(n15846) );
  AOI22_X1 U18998 ( .A1(n15844), .A2(n20086), .B1(n20063), .B2(n15843), .ZN(
        n15845) );
  OAI211_X1 U18999 ( .C1(n15848), .C2(n15847), .A(n15846), .B(n15845), .ZN(
        P1_U3018) );
  NOR2_X1 U19000 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n15852), .ZN(
        n15864) );
  INV_X1 U19001 ( .A(n15864), .ZN(n15853) );
  INV_X1 U19002 ( .A(n15872), .ZN(n20073) );
  INV_X1 U19003 ( .A(n15849), .ZN(n15893) );
  OAI221_X1 U19004 ( .B1(n20080), .B2(n15893), .C1(n20080), .C2(n15855), .A(
        n15870), .ZN(n15850) );
  AOI221_X1 U19005 ( .B1(n15852), .B2(n20073), .C1(n15851), .C2(n20073), .A(
        n15850), .ZN(n15869) );
  OAI21_X1 U19006 ( .B1(n15854), .B2(n15853), .A(n15869), .ZN(n15859) );
  NAND2_X1 U19007 ( .A1(n15855), .A2(n15900), .ZN(n15856) );
  OAI22_X1 U19008 ( .A1(n15857), .A2(n15923), .B1(
        P1_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n15856), .ZN(n15858) );
  AOI21_X1 U19009 ( .B1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n15859), .A(
        n15858), .ZN(n15861) );
  NAND2_X1 U19010 ( .A1(n11744), .A2(P1_REIP_REG_12__SCAN_IN), .ZN(n15860) );
  OAI211_X1 U19011 ( .C1(n20083), .C2(n15862), .A(n15861), .B(n15860), .ZN(
        P1_U3019) );
  AOI22_X1 U19012 ( .A1(n11744), .A2(P1_REIP_REG_11__SCAN_IN), .B1(n20063), 
        .B2(n15863), .ZN(n15867) );
  AOI22_X1 U19013 ( .A1(n15865), .A2(n20086), .B1(n15864), .B2(n15900), .ZN(
        n15866) );
  OAI211_X1 U19014 ( .C1(n15869), .C2(n15868), .A(n15867), .B(n15866), .ZN(
        P1_U3020) );
  OAI21_X1 U19015 ( .B1(n15872), .B2(n15871), .A(n15870), .ZN(n20052) );
  NAND2_X1 U19016 ( .A1(n15876), .A2(n15893), .ZN(n15874) );
  OAI21_X1 U19017 ( .B1(n20052), .B2(n15874), .A(n15873), .ZN(n15892) );
  INV_X1 U19018 ( .A(n15875), .ZN(n15881) );
  NAND2_X1 U19019 ( .A1(n15876), .A2(n15900), .ZN(n15887) );
  AOI221_X1 U19020 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .C1(n11648), .C2(n13937), .A(
        n15887), .ZN(n15877) );
  AOI21_X1 U19021 ( .B1(n11744), .B2(P1_REIP_REG_10__SCAN_IN), .A(n15877), 
        .ZN(n15878) );
  OAI21_X1 U19022 ( .B1(n20083), .B2(n15879), .A(n15878), .ZN(n15880) );
  AOI21_X1 U19023 ( .B1(n15881), .B2(n20086), .A(n15880), .ZN(n15882) );
  OAI21_X1 U19024 ( .B1(n11648), .B2(n15892), .A(n15882), .ZN(P1_U3021) );
  OR2_X1 U19025 ( .A1(n15884), .A2(n15883), .ZN(n15885) );
  AND2_X1 U19026 ( .A1(n15886), .A2(n15885), .ZN(n19958) );
  NOR2_X1 U19027 ( .A1(n20081), .A2(n13939), .ZN(n15890) );
  OAI22_X1 U19028 ( .A1(n15888), .A2(n15923), .B1(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n15887), .ZN(n15889) );
  AOI211_X1 U19029 ( .C1(n20063), .C2(n19958), .A(n15890), .B(n15889), .ZN(
        n15891) );
  OAI21_X1 U19030 ( .B1(n13937), .B2(n15892), .A(n15891), .ZN(P1_U3022) );
  NAND2_X1 U19031 ( .A1(n20054), .A2(n20974), .ZN(n15928) );
  NOR2_X1 U19032 ( .A1(n15893), .A2(n20080), .ZN(n15894) );
  AOI211_X1 U19033 ( .C1(n20073), .C2(n15895), .A(n15894), .B(n20052), .ZN(
        n15922) );
  OAI21_X1 U19034 ( .B1(n15896), .B2(n15928), .A(n15922), .ZN(n15913) );
  AOI21_X1 U19035 ( .B1(n15898), .B2(n15897), .A(n15913), .ZN(n15910) );
  INV_X1 U19036 ( .A(n15899), .ZN(n15905) );
  NAND2_X1 U19037 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n15900), .ZN(
        n15912) );
  AOI221_X1 U19038 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(n11511), .C2(n15911), .A(
        n15912), .ZN(n15904) );
  OAI22_X1 U19039 ( .A1(n20083), .A2(n15902), .B1(n15901), .B2(n20081), .ZN(
        n15903) );
  AOI211_X1 U19040 ( .C1(n15905), .C2(n20086), .A(n15904), .B(n15903), .ZN(
        n15906) );
  OAI21_X1 U19041 ( .B1(n15910), .B2(n11511), .A(n15906), .ZN(P1_U3023) );
  AOI222_X1 U19042 ( .A1(n15908), .A2(n20086), .B1(n20063), .B2(n15907), .C1(
        P1_REIP_REG_7__SCAN_IN), .C2(n11744), .ZN(n15909) );
  OAI221_X1 U19043 ( .B1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n15912), .C1(
        n15911), .C2(n15910), .A(n15909), .ZN(P1_U3024) );
  AOI22_X1 U19044 ( .A1(n11744), .A2(P1_REIP_REG_6__SCAN_IN), .B1(n20063), 
        .B2(n19910), .ZN(n15916) );
  AOI22_X1 U19045 ( .A1(n15914), .A2(n20086), .B1(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n15913), .ZN(n15915) );
  OAI211_X1 U19046 ( .C1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n15917), .A(
        n15916), .B(n15915), .ZN(P1_U3025) );
  INV_X1 U19047 ( .A(n20065), .ZN(n20055) );
  NAND2_X1 U19048 ( .A1(n15919), .A2(n15918), .ZN(n15920) );
  AND2_X1 U19049 ( .A1(n15921), .A2(n15920), .ZN(n19961) );
  AOI22_X1 U19050 ( .A1(n11744), .A2(P1_REIP_REG_5__SCAN_IN), .B1(n20063), 
        .B2(n19961), .ZN(n15927) );
  OAI22_X1 U19051 ( .A1(n15924), .A2(n15923), .B1(n15922), .B2(n20974), .ZN(
        n15925) );
  INV_X1 U19052 ( .A(n15925), .ZN(n15926) );
  OAI211_X1 U19053 ( .C1(n20055), .C2(n15928), .A(n15927), .B(n15926), .ZN(
        P1_U3026) );
  OAI22_X1 U19054 ( .A1(n20574), .A2(n15931), .B1(n15930), .B2(n15929), .ZN(
        n20686) );
  OAI21_X1 U19055 ( .B1(n15933), .B2(n20686), .A(n15932), .ZN(n15934) );
  OAI221_X1 U19056 ( .B1(n15935), .B2(n20493), .C1(n15935), .C2(n20697), .A(
        n15934), .ZN(n15936) );
  AOI221_X1 U19057 ( .B1(n15938), .B2(n15937), .C1(n20098), .C2(n15937), .A(
        n15936), .ZN(P1_U3162) );
  NOR2_X1 U19058 ( .A1(n15938), .A2(n20098), .ZN(n15940) );
  OAI22_X1 U19059 ( .A1(n20493), .A2(n15940), .B1(n15939), .B2(n20098), .ZN(
        P1_U3466) );
  INV_X1 U19060 ( .A(n16020), .ZN(n15946) );
  INV_X1 U19061 ( .A(n15941), .ZN(n15944) );
  OAI22_X1 U19062 ( .A1(n18960), .A2(n16019), .B1(n10037), .B2(n18987), .ZN(
        n15942) );
  AOI21_X1 U19063 ( .B1(P2_REIP_REG_31__SCAN_IN), .B2(n18989), .A(n15942), 
        .ZN(n15943) );
  OAI21_X1 U19064 ( .B1(n15944), .B2(n18994), .A(n15943), .ZN(n15945) );
  AOI21_X1 U19065 ( .B1(n15946), .B2(n18997), .A(n15945), .ZN(n15950) );
  NAND4_X1 U19066 ( .A1(n18999), .A2(n15948), .A3(n18873), .A4(n15947), .ZN(
        n15949) );
  OAI211_X1 U19067 ( .C1(n15951), .C2(n18982), .A(n15950), .B(n15949), .ZN(
        P2_U2824) );
  AOI22_X1 U19068 ( .A1(n15952), .A2(n18950), .B1(P2_EBX_REG_29__SCAN_IN), 
        .B2(n18990), .ZN(n15961) );
  AOI22_X1 U19069 ( .A1(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n19002), .B1(
        P2_REIP_REG_29__SCAN_IN), .B2(n18989), .ZN(n15960) );
  AOI22_X1 U19070 ( .A1(n15954), .A2(n18997), .B1(n15953), .B2(n18991), .ZN(
        n15959) );
  OAI211_X1 U19071 ( .C1(n15957), .C2(n15956), .A(n18999), .B(n15955), .ZN(
        n15958) );
  NAND4_X1 U19072 ( .A1(n15961), .A2(n15960), .A3(n15959), .A4(n15958), .ZN(
        P2_U2826) );
  INV_X1 U19073 ( .A(P2_EBX_REG_27__SCAN_IN), .ZN(n15963) );
  OAI22_X1 U19074 ( .A1(n18960), .A2(n15963), .B1(n15962), .B2(n18987), .ZN(
        n15964) );
  AOI21_X1 U19075 ( .B1(P2_REIP_REG_27__SCAN_IN), .B2(n18989), .A(n15964), 
        .ZN(n15965) );
  OAI21_X1 U19076 ( .B1(n15966), .B2(n18994), .A(n15965), .ZN(n15967) );
  AOI21_X1 U19077 ( .B1(n15968), .B2(n18997), .A(n15967), .ZN(n15973) );
  OAI211_X1 U19078 ( .C1(n15971), .C2(n15970), .A(n18999), .B(n15969), .ZN(
        n15972) );
  OAI211_X1 U19079 ( .C1(n18982), .C2(n15974), .A(n15973), .B(n15972), .ZN(
        P2_U2828) );
  AOI22_X1 U19080 ( .A1(n15975), .A2(n18950), .B1(P2_REIP_REG_26__SCAN_IN), 
        .B2(n18989), .ZN(n15985) );
  AOI22_X1 U19081 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(n18990), .B1(
        P2_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n18964), .ZN(n15984) );
  OAI22_X1 U19082 ( .A1(n15977), .A2(n18981), .B1(n15976), .B2(n18982), .ZN(
        n15978) );
  INV_X1 U19083 ( .A(n15978), .ZN(n15983) );
  OAI211_X1 U19084 ( .C1(n15981), .C2(n15980), .A(n18999), .B(n15979), .ZN(
        n15982) );
  NAND4_X1 U19085 ( .A1(n15985), .A2(n15984), .A3(n15983), .A4(n15982), .ZN(
        P2_U2829) );
  AOI22_X1 U19086 ( .A1(n15986), .A2(n18950), .B1(P2_REIP_REG_25__SCAN_IN), 
        .B2(n18989), .ZN(n15996) );
  AOI22_X1 U19087 ( .A1(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n18964), .B1(
        P2_EBX_REG_25__SCAN_IN), .B2(n18990), .ZN(n15995) );
  OAI22_X1 U19088 ( .A1(n15988), .A2(n18981), .B1(n15987), .B2(n18982), .ZN(
        n15989) );
  INV_X1 U19089 ( .A(n15989), .ZN(n15994) );
  OAI211_X1 U19090 ( .C1(n15992), .C2(n15991), .A(n18999), .B(n15990), .ZN(
        n15993) );
  NAND4_X1 U19091 ( .A1(n15996), .A2(n15995), .A3(n15994), .A4(n15993), .ZN(
        P2_U2830) );
  AOI22_X1 U19092 ( .A1(n15997), .A2(n18950), .B1(P2_EBX_REG_24__SCAN_IN), 
        .B2(n18990), .ZN(n16006) );
  AOI22_X1 U19093 ( .A1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n19002), .B1(
        P2_REIP_REG_24__SCAN_IN), .B2(n18989), .ZN(n16005) );
  AOI22_X1 U19094 ( .A1(n15999), .A2(n18997), .B1(n18991), .B2(n15998), .ZN(
        n16004) );
  OAI211_X1 U19095 ( .C1(n16002), .C2(n16001), .A(n18999), .B(n16000), .ZN(
        n16003) );
  NAND4_X1 U19096 ( .A1(n16006), .A2(n16005), .A3(n16004), .A4(n16003), .ZN(
        P2_U2831) );
  NOR2_X1 U19097 ( .A1(n18960), .A2(n12132), .ZN(n16008) );
  OAI22_X1 U19098 ( .A1(n12091), .A2(n18987), .B1(n19756), .B2(n18973), .ZN(
        n16007) );
  NOR2_X1 U19099 ( .A1(n16008), .A2(n16007), .ZN(n16009) );
  OAI21_X1 U19100 ( .B1(n16010), .B2(n18981), .A(n16009), .ZN(n16011) );
  AOI21_X1 U19101 ( .B1(n16012), .B2(n18950), .A(n16011), .ZN(n16017) );
  OAI211_X1 U19102 ( .C1(n16015), .C2(n16014), .A(n18999), .B(n16013), .ZN(
        n16016) );
  OAI211_X1 U19103 ( .C1(n18982), .C2(n16018), .A(n16017), .B(n16016), .ZN(
        P2_U2832) );
  AOI22_X1 U19104 ( .A1(n19020), .A2(n16020), .B1(n16019), .B2(n19037), .ZN(
        P2_U2856) );
  INV_X1 U19105 ( .A(n16021), .ZN(n16023) );
  AOI21_X1 U19106 ( .B1(n16023), .B2(n9878), .A(n16022), .ZN(n16035) );
  AOI22_X1 U19107 ( .A1(n16035), .A2(n19038), .B1(P2_EBX_REG_22__SCAN_IN), 
        .B2(n19037), .ZN(n16024) );
  OAI21_X1 U19108 ( .B1(n19037), .B2(n16054), .A(n16024), .ZN(P2_U2865) );
  AND2_X1 U19109 ( .A1(n16026), .A2(n16025), .ZN(n16027) );
  OR2_X1 U19110 ( .A1(n16027), .A2(n14729), .ZN(n16041) );
  OAI22_X1 U19111 ( .A1(n16041), .A2(n19031), .B1(n19037), .B2(n18825), .ZN(
        n16028) );
  INV_X1 U19112 ( .A(n16028), .ZN(n16029) );
  OAI21_X1 U19113 ( .B1(n19020), .B2(n10112), .A(n16029), .ZN(P2_U2867) );
  AOI21_X1 U19114 ( .B1(n16031), .B2(n14734), .A(n16030), .ZN(n16050) );
  AOI22_X1 U19115 ( .A1(n16050), .A2(n19038), .B1(P2_EBX_REG_18__SCAN_IN), 
        .B2(n19037), .ZN(n16032) );
  OAI21_X1 U19116 ( .B1(n19037), .B2(n18851), .A(n16032), .ZN(P2_U2869) );
  AOI22_X1 U19117 ( .A1(n16047), .A2(n16033), .B1(P2_EAX_REG_22__SCAN_IN), 
        .B2(n19083), .ZN(n16038) );
  AOI22_X1 U19118 ( .A1(n16049), .A2(BUF1_REG_22__SCAN_IN), .B1(n16048), .B2(
        BUF2_REG_22__SCAN_IN), .ZN(n16037) );
  AOI22_X1 U19119 ( .A1(n16035), .A2(n19086), .B1(n19084), .B2(n16034), .ZN(
        n16036) );
  NAND3_X1 U19120 ( .A1(n16038), .A2(n16037), .A3(n16036), .ZN(P2_U2897) );
  AOI22_X1 U19121 ( .A1(n16047), .A2(n19062), .B1(P2_EAX_REG_20__SCAN_IN), 
        .B2(n19083), .ZN(n16045) );
  AOI22_X1 U19122 ( .A1(n16049), .A2(BUF1_REG_20__SCAN_IN), .B1(n16048), .B2(
        BUF2_REG_20__SCAN_IN), .ZN(n16044) );
  INV_X1 U19123 ( .A(n16039), .ZN(n18824) );
  OAI22_X1 U19124 ( .A1(n16041), .A2(n19079), .B1(n16040), .B2(n18824), .ZN(
        n16042) );
  INV_X1 U19125 ( .A(n16042), .ZN(n16043) );
  NAND3_X1 U19126 ( .A1(n16045), .A2(n16044), .A3(n16043), .ZN(P2_U2899) );
  AOI22_X1 U19127 ( .A1(n16047), .A2(n16046), .B1(P2_EAX_REG_18__SCAN_IN), 
        .B2(n19083), .ZN(n16053) );
  AOI22_X1 U19128 ( .A1(n16049), .A2(BUF1_REG_18__SCAN_IN), .B1(n16048), .B2(
        BUF2_REG_18__SCAN_IN), .ZN(n16052) );
  AOI22_X1 U19129 ( .A1(n16050), .A2(n19086), .B1(n19084), .B2(n18849), .ZN(
        n16051) );
  NAND3_X1 U19130 ( .A1(n16053), .A2(n16052), .A3(n16051), .ZN(P2_U2901) );
  AOI22_X1 U19131 ( .A1(n16062), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n18976), .ZN(n16060) );
  OAI22_X1 U19132 ( .A1(n16056), .A2(n16055), .B1(n16088), .B2(n16054), .ZN(
        n16057) );
  AOI21_X1 U19133 ( .B1(n16118), .B2(n16058), .A(n16057), .ZN(n16059) );
  OAI211_X1 U19134 ( .C1(n16068), .C2(n16061), .A(n16060), .B(n16059), .ZN(
        P2_U2992) );
  AOI22_X1 U19135 ( .A1(n16062), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B1(
        P2_REIP_REG_18__SCAN_IN), .B2(n18976), .ZN(n16067) );
  INV_X1 U19136 ( .A(n18851), .ZN(n16064) );
  AOI222_X1 U19137 ( .A1(n16065), .A2(n16118), .B1(n16117), .B2(n16064), .C1(
        n16120), .C2(n16063), .ZN(n16066) );
  OAI211_X1 U19138 ( .C1(n16068), .C2(n18855), .A(n16067), .B(n16066), .ZN(
        P2_U2996) );
  AOI22_X1 U19139 ( .A1(P2_REIP_REG_14__SCAN_IN), .A2(n18976), .B1(n16114), 
        .B2(n16069), .ZN(n16077) );
  AOI21_X1 U19140 ( .B1(n11105), .B2(n16071), .A(n16070), .ZN(n16142) );
  NAND2_X1 U19141 ( .A1(n16073), .A2(n16072), .ZN(n16074) );
  XNOR2_X1 U19142 ( .A(n16075), .B(n16074), .ZN(n16141) );
  INV_X1 U19143 ( .A(n19014), .ZN(n16140) );
  AOI222_X1 U19144 ( .A1(n16142), .A2(n16120), .B1(n16118), .B2(n16141), .C1(
        n16117), .C2(n16140), .ZN(n16076) );
  OAI211_X1 U19145 ( .C1(n16125), .C2(n16078), .A(n16077), .B(n16076), .ZN(
        P2_U3000) );
  AOI22_X1 U19146 ( .A1(P2_REIP_REG_12__SCAN_IN), .A2(n18976), .B1(n16114), 
        .B2(n16079), .ZN(n16091) );
  AOI21_X1 U19147 ( .B1(n16161), .B2(n16081), .A(n16080), .ZN(n16166) );
  NAND2_X1 U19148 ( .A1(n10103), .A2(n16083), .ZN(n16087) );
  NAND2_X1 U19149 ( .A1(n16085), .A2(n16084), .ZN(n16086) );
  XOR2_X1 U19150 ( .A(n16087), .B(n16086), .Z(n16169) );
  OAI22_X1 U19151 ( .A1(n16169), .A2(n15067), .B1(n16088), .B2(n19023), .ZN(
        n16089) );
  AOI21_X1 U19152 ( .B1(n16166), .B2(n16120), .A(n16089), .ZN(n16090) );
  OAI211_X1 U19153 ( .C1(n16125), .C2(n16092), .A(n16091), .B(n16090), .ZN(
        P2_U3002) );
  AOI22_X1 U19154 ( .A1(P2_REIP_REG_10__SCAN_IN), .A2(n18976), .B1(n16114), 
        .B2(n18924), .ZN(n16097) );
  AOI222_X1 U19155 ( .A1(n16095), .A2(n16118), .B1(n16117), .B2(n16094), .C1(
        n16120), .C2(n16093), .ZN(n16096) );
  OAI211_X1 U19156 ( .C1(n16125), .C2(n16098), .A(n16097), .B(n16096), .ZN(
        P2_U3004) );
  AOI22_X1 U19157 ( .A1(P2_REIP_REG_8__SCAN_IN), .A2(n18976), .B1(n16114), 
        .B2(n16099), .ZN(n16112) );
  AOI21_X1 U19158 ( .B1(n15101), .B2(n16101), .A(n16100), .ZN(n16106) );
  INV_X1 U19159 ( .A(n16102), .ZN(n16103) );
  NOR2_X1 U19160 ( .A1(n16104), .A2(n16103), .ZN(n16105) );
  XNOR2_X1 U19161 ( .A(n16106), .B(n16105), .ZN(n16185) );
  OAI21_X1 U19162 ( .B1(n16109), .B2(n16108), .A(n9797), .ZN(n16110) );
  INV_X1 U19163 ( .A(n16110), .ZN(n16183) );
  AOI222_X1 U19164 ( .A1(n16185), .A2(n16118), .B1(n16117), .B2(n16184), .C1(
        n16120), .C2(n16183), .ZN(n16111) );
  OAI211_X1 U19165 ( .C1(n16125), .C2(n16113), .A(n16112), .B(n16111), .ZN(
        P2_U3006) );
  AOI22_X1 U19166 ( .A1(P2_REIP_REG_6__SCAN_IN), .A2(n18976), .B1(n16114), 
        .B2(n18967), .ZN(n16123) );
  INV_X1 U19167 ( .A(n16115), .ZN(n16121) );
  INV_X1 U19168 ( .A(n16116), .ZN(n18968) );
  AOI222_X1 U19169 ( .A1(n16121), .A2(n16120), .B1(n16119), .B2(n16118), .C1(
        n16117), .C2(n18968), .ZN(n16122) );
  OAI211_X1 U19170 ( .C1(n16125), .C2(n16124), .A(n16123), .B(n16122), .ZN(
        P2_U3008) );
  INV_X1 U19171 ( .A(n18838), .ZN(n16126) );
  OAI22_X1 U19172 ( .A1(n21133), .A2(n16126), .B1(n21044), .B2(n9889), .ZN(
        n16127) );
  AOI221_X1 U19173 ( .B1(n16130), .B2(n16129), .C1(n16128), .C2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(n16127), .ZN(n16134) );
  INV_X1 U19174 ( .A(n16131), .ZN(n18839) );
  AOI22_X1 U19175 ( .A1(n16132), .A2(n21137), .B1(n21130), .B2(n18839), .ZN(
        n16133) );
  OAI211_X1 U19176 ( .C1(n21140), .C2(n16135), .A(n16134), .B(n16133), .ZN(
        P2_U3027) );
  INV_X1 U19177 ( .A(n16136), .ZN(n16137) );
  AOI21_X1 U19178 ( .B1(n16139), .B2(n16138), .A(n16137), .ZN(n16162) );
  OAI21_X1 U19179 ( .B1(n16149), .B2(n16143), .A(n16162), .ZN(n16152) );
  AOI22_X1 U19180 ( .A1(n16181), .A2(n19042), .B1(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n16152), .ZN(n16147) );
  AOI222_X1 U19181 ( .A1(n16142), .A2(n21137), .B1(n11126), .B2(n16141), .C1(
        n21130), .C2(n16140), .ZN(n16146) );
  NAND2_X1 U19182 ( .A1(P2_REIP_REG_14__SCAN_IN), .A2(n18976), .ZN(n16145) );
  NAND3_X1 U19183 ( .A1(n16143), .A2(n16158), .A3(n11105), .ZN(n16144) );
  NAND4_X1 U19184 ( .A1(n16147), .A2(n16146), .A3(n16145), .A4(n16144), .ZN(
        P2_U3032) );
  OAI21_X1 U19185 ( .B1(n16161), .B2(n16149), .A(n16148), .ZN(n16151) );
  OAI22_X1 U19186 ( .A1(n21133), .A2(n18906), .B1(n10995), .B2(n9889), .ZN(
        n16150) );
  AOI21_X1 U19187 ( .B1(n16152), .B2(n16151), .A(n16150), .ZN(n16155) );
  AOI22_X1 U19188 ( .A1(n16153), .A2(n11126), .B1(n21130), .B2(n18903), .ZN(
        n16154) );
  OAI211_X1 U19189 ( .C1(n16157), .C2(n16156), .A(n16155), .B(n16154), .ZN(
        P2_U3033) );
  NAND2_X1 U19190 ( .A1(n16158), .A2(n16161), .ZN(n16160) );
  NAND2_X1 U19191 ( .A1(P2_REIP_REG_12__SCAN_IN), .A2(n18976), .ZN(n16159) );
  OAI211_X1 U19192 ( .C1(n16162), .C2(n16161), .A(n16160), .B(n16159), .ZN(
        n16163) );
  AOI21_X1 U19193 ( .B1(n16164), .B2(n16181), .A(n16163), .ZN(n16168) );
  INV_X1 U19194 ( .A(n19023), .ZN(n16165) );
  AOI22_X1 U19195 ( .A1(n16166), .A2(n21137), .B1(n21130), .B2(n16165), .ZN(
        n16167) );
  OAI211_X1 U19196 ( .C1(n16169), .C2(n21140), .A(n16168), .B(n16167), .ZN(
        P2_U3034) );
  OAI21_X1 U19197 ( .B1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(n16170), .ZN(n16171) );
  OAI22_X1 U19198 ( .A1(n18914), .A2(n21133), .B1(n16172), .B2(n16171), .ZN(
        n16173) );
  AOI211_X1 U19199 ( .C1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n16175), .A(
        n16174), .B(n16173), .ZN(n16178) );
  AOI22_X1 U19200 ( .A1(n16176), .A2(n21137), .B1(n21130), .B2(n18907), .ZN(
        n16177) );
  OAI211_X1 U19201 ( .C1(n16179), .C2(n21140), .A(n16178), .B(n16177), .ZN(
        P2_U3035) );
  AOI22_X1 U19202 ( .A1(n16182), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B1(
        n16181), .B2(n16180), .ZN(n16192) );
  AOI222_X1 U19203 ( .A1(n16185), .A2(n11126), .B1(n21130), .B2(n16184), .C1(
        n21137), .C2(n16183), .ZN(n16191) );
  NAND2_X1 U19204 ( .A1(P2_REIP_REG_8__SCAN_IN), .A2(n16186), .ZN(n16190) );
  OAI211_X1 U19205 ( .C1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n16188), .B(n16187), .ZN(n16189) );
  NAND4_X1 U19206 ( .A1(n16192), .A2(n16191), .A3(n16190), .A4(n16189), .ZN(
        P2_U3038) );
  NAND2_X1 U19207 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19149), .ZN(n19702) );
  INV_X1 U19208 ( .A(n16232), .ZN(n16200) );
  NAND2_X1 U19209 ( .A1(n16193), .A2(n16200), .ZN(n16196) );
  NAND2_X1 U19210 ( .A1(n16232), .A2(n16194), .ZN(n16195) );
  NAND2_X1 U19211 ( .A1(n16196), .A2(n16195), .ZN(n16234) );
  INV_X1 U19212 ( .A(n16234), .ZN(n16209) );
  INV_X1 U19213 ( .A(n16197), .ZN(n16199) );
  AOI22_X1 U19214 ( .A1(n16199), .A2(n19353), .B1(n19813), .B2(n19821), .ZN(
        n16206) );
  OAI21_X1 U19215 ( .B1(n16199), .B2(n19813), .A(n16198), .ZN(n16205) );
  MUX2_X1 U19216 ( .A(n10330), .B(n16201), .S(n16200), .Z(n16235) );
  INV_X1 U19217 ( .A(n16235), .ZN(n16203) );
  AOI21_X1 U19218 ( .B1(n16234), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n16202) );
  AOI21_X1 U19219 ( .B1(n16203), .B2(n19804), .A(n16202), .ZN(n16204) );
  AOI211_X1 U19220 ( .C1(n16206), .C2(n16205), .A(n16232), .B(n16204), .ZN(
        n16207) );
  AOI21_X1 U19221 ( .B1(n16209), .B2(n16208), .A(n16207), .ZN(n16210) );
  AOI221_X1 U19222 ( .B1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n16210), 
        .C1(n16235), .C2(n16210), .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(
        n16237) );
  INV_X1 U19223 ( .A(n16211), .ZN(n16216) );
  INV_X1 U19224 ( .A(n16212), .ZN(n16221) );
  NAND2_X1 U19225 ( .A1(n16223), .A2(n16221), .ZN(n16215) );
  NAND2_X1 U19226 ( .A1(n16217), .A2(n16213), .ZN(n16214) );
  OAI211_X1 U19227 ( .C1(n16217), .C2(n16216), .A(n16215), .B(n16214), .ZN(
        n19830) );
  INV_X1 U19228 ( .A(n19830), .ZN(n16230) );
  NAND2_X1 U19229 ( .A1(n16219), .A2(n16218), .ZN(n16229) );
  OR2_X1 U19230 ( .A1(n10495), .A2(n16220), .ZN(n19843) );
  AOI21_X1 U19231 ( .B1(n19835), .B2(n19843), .A(n16221), .ZN(n16222) );
  AND2_X1 U19232 ( .A1(n16223), .A2(n16222), .ZN(n18789) );
  OAI21_X1 U19233 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(P2_MORE_REG_SCAN_IN), .A(
        n18789), .ZN(n16228) );
  INV_X1 U19234 ( .A(n16224), .ZN(n16225) );
  NAND3_X1 U19235 ( .A1(n16226), .A2(n9776), .A3(n16225), .ZN(n16227) );
  NAND4_X1 U19236 ( .A1(n16230), .A2(n16229), .A3(n16228), .A4(n16227), .ZN(
        n16231) );
  AOI21_X1 U19237 ( .B1(n16232), .B2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n16231), .ZN(n16233) );
  OAI21_X1 U19238 ( .B1(n16235), .B2(n16234), .A(n16233), .ZN(n16236) );
  OR2_X1 U19239 ( .A1(n16237), .A2(n16236), .ZN(n16241) );
  NAND2_X1 U19240 ( .A1(n9776), .A2(n16238), .ZN(n16239) );
  OR2_X1 U19241 ( .A1(n10953), .A2(n16239), .ZN(n16242) );
  OAI21_X1 U19242 ( .B1(n16241), .B2(n16242), .A(n19840), .ZN(n16240) );
  INV_X1 U19243 ( .A(n16240), .ZN(n16247) );
  OAI21_X1 U19244 ( .B1(n16241), .B2(n18788), .A(n19123), .ZN(n16243) );
  AOI21_X1 U19245 ( .B1(n19836), .B2(n16244), .A(n19849), .ZN(n16245) );
  AOI21_X1 U19246 ( .B1(n19707), .B2(n19844), .A(n16245), .ZN(n16246) );
  AOI211_X1 U19247 ( .C1(n16249), .C2(n16248), .A(n16247), .B(n16246), .ZN(
        n16251) );
  OAI211_X1 U19248 ( .C1(n19835), .C2(n19702), .A(n16251), .B(n16250), .ZN(
        P2_U3176) );
  INV_X1 U19249 ( .A(n19707), .ZN(n16253) );
  OAI221_X1 U19250 ( .B1(n19796), .B2(P2_STATE2_REG_0__SCAN_IN), .C1(n19796), 
        .C2(n16253), .A(n16252), .ZN(P2_U3593) );
  INV_X1 U19251 ( .A(n16254), .ZN(n16285) );
  NAND2_X1 U19252 ( .A1(n16285), .A2(n17587), .ZN(n17436) );
  INV_X1 U19253 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16457) );
  XNOR2_X1 U19254 ( .A(n16457), .B(n16277), .ZN(n16456) );
  OAI221_X1 U19255 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n16257), .C1(
        n16457), .C2(n16256), .A(n16255), .ZN(n16258) );
  AOI21_X1 U19256 ( .B1(n17638), .B2(n16456), .A(n16258), .ZN(n16264) );
  INV_X1 U19257 ( .A(n17696), .ZN(n17616) );
  NAND2_X1 U19258 ( .A1(n17773), .A2(n16259), .ZN(n16271) );
  OAI21_X1 U19259 ( .B1(n16260), .B2(n17616), .A(n16271), .ZN(n16262) );
  AOI22_X1 U19260 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16262), .B1(
        n17695), .B2(n16261), .ZN(n16263) );
  OAI211_X1 U19261 ( .C1(n16265), .C2(n17436), .A(n16264), .B(n16263), .ZN(
        P3_U2800) );
  OAI21_X1 U19262 ( .B1(n18428), .B2(n16266), .A(n16278), .ZN(n16268) );
  AOI21_X1 U19263 ( .B1(n16269), .B2(n16268), .A(n16267), .ZN(n16283) );
  NAND2_X1 U19264 ( .A1(n17791), .A2(n16270), .ZN(n16300) );
  AOI21_X1 U19265 ( .B1(n16272), .B2(n16300), .A(n16271), .ZN(n16273) );
  AOI21_X1 U19266 ( .B1(n16274), .B2(n17695), .A(n16273), .ZN(n16282) );
  NOR2_X1 U19267 ( .A1(n16275), .A2(n17793), .ZN(n16301) );
  OAI211_X1 U19268 ( .C1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n16301), .A(
        n17696), .B(n16276), .ZN(n16281) );
  AOI21_X1 U19269 ( .B1(n16278), .B2(n16439), .A(n16277), .ZN(n16467) );
  OAI21_X1 U19270 ( .B1(n16279), .B2(n17638), .A(n16467), .ZN(n16280) );
  NAND4_X1 U19271 ( .A1(n16283), .A2(n16282), .A3(n16281), .A4(n16280), .ZN(
        P3_U2801) );
  NOR3_X1 U19272 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n20896), .A3(
        n16284), .ZN(n16286) );
  NAND3_X1 U19273 ( .A1(n16286), .A2(n16285), .A3(n17813), .ZN(n16288) );
  OAI22_X1 U19274 ( .A1(n18084), .A2(n16288), .B1(n16287), .B2(n18728), .ZN(
        n16289) );
  AOI211_X1 U19275 ( .C1(n16292), .C2(n16291), .A(n16290), .B(n16289), .ZN(
        n16296) );
  AOI22_X1 U19276 ( .A1(n16294), .A2(n18017), .B1(n16293), .B2(n18015), .ZN(
        n16295) );
  OAI211_X1 U19277 ( .C1(n16297), .C2(n18097), .A(n16296), .B(n16295), .ZN(
        P3_U2831) );
  NAND2_X1 U19278 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n16298), .ZN(
        n17430) );
  AOI22_X1 U19279 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17628), .B1(
        n17694), .B2(n16298), .ZN(n17419) );
  AOI21_X1 U19280 ( .B1(n17694), .B2(n17433), .A(n16309), .ZN(n17418) );
  NOR2_X1 U19281 ( .A1(n17419), .A2(n17418), .ZN(n17417) );
  NOR4_X1 U19282 ( .A1(n16299), .A2(n17274), .A3(n17417), .A4(n18557), .ZN(
        n16307) );
  INV_X1 U19283 ( .A(n16300), .ZN(n16305) );
  OR2_X1 U19284 ( .A1(n16301), .A2(n17954), .ZN(n16303) );
  AND2_X1 U19285 ( .A1(n16303), .A2(n15563), .ZN(n16304) );
  OAI21_X1 U19286 ( .B1(n16305), .B2(n18072), .A(n16304), .ZN(n16306) );
  OR2_X1 U19287 ( .A1(n16307), .A2(n16306), .ZN(n16308) );
  AND2_X1 U19288 ( .A1(n16308), .A2(n18091), .ZN(n16313) );
  AND3_X1 U19289 ( .A1(n16309), .A2(n18015), .A3(n17419), .ZN(n16312) );
  NOR3_X1 U19290 ( .A1(n17433), .A2(n18095), .A3(n16310), .ZN(n16311) );
  AOI211_X1 U19291 ( .C1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .C2(n16313), .A(
        n16312), .B(n16311), .ZN(n16314) );
  NAND2_X1 U19292 ( .A1(n18093), .A2(P3_REIP_REG_28__SCAN_IN), .ZN(n17423) );
  OAI211_X1 U19293 ( .C1(n17794), .C2(n17430), .A(n16314), .B(n17423), .ZN(
        P3_U2834) );
  NOR3_X1 U19294 ( .A1(P3_W_R_N_REG_SCAN_IN), .A2(P3_BE_N_REG_0__SCAN_IN), 
        .A3(P3_BE_N_REG_1__SCAN_IN), .ZN(n16316) );
  NOR4_X1 U19295 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n16315) );
  NAND4_X1 U19296 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n16316), .A3(n16315), .A4(
        U215), .ZN(U213) );
  INV_X2 U19297 ( .A(U214), .ZN(n16370) );
  NOR2_X1 U19298 ( .A1(n16370), .A2(n16317), .ZN(n16322) );
  INV_X1 U19299 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n19093) );
  OAI222_X1 U19300 ( .A1(U214), .A2(n16406), .B1(n16373), .B2(n16318), .C1(
        U212), .C2(n19093), .ZN(U216) );
  INV_X1 U19301 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n16319) );
  INV_X1 U19302 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n20870) );
  INV_X1 U19303 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n19096) );
  OAI222_X1 U19304 ( .A1(U214), .A2(n16319), .B1(n16373), .B2(n20870), .C1(
        U212), .C2(n19096), .ZN(U217) );
  INV_X1 U19305 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n16321) );
  INV_X2 U19306 ( .A(U212), .ZN(n16371) );
  AOI22_X1 U19307 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(n16371), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n16370), .ZN(n16320) );
  OAI21_X1 U19308 ( .B1(n16321), .B2(n16373), .A(n16320), .ZN(U218) );
  AOI222_X1 U19309 ( .A1(n16370), .A2(P1_DATAO_REG_28__SCAN_IN), .B1(n16322), 
        .B2(BUF1_REG_28__SCAN_IN), .C1(n16371), .C2(P2_DATAO_REG_28__SCAN_IN), 
        .ZN(n16323) );
  INV_X1 U19310 ( .A(n16323), .ZN(U219) );
  AOI22_X1 U19311 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(n16371), .B1(
        P1_DATAO_REG_27__SCAN_IN), .B2(n16370), .ZN(n16324) );
  OAI21_X1 U19312 ( .B1(n16325), .B2(n16373), .A(n16324), .ZN(U220) );
  INV_X1 U19313 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n20863) );
  AOI22_X1 U19314 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(n16371), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n16370), .ZN(n16326) );
  OAI21_X1 U19315 ( .B1(n20863), .B2(n16373), .A(n16326), .ZN(U221) );
  INV_X1 U19316 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n16328) );
  AOI22_X1 U19317 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(n16371), .B1(
        P1_DATAO_REG_25__SCAN_IN), .B2(n16370), .ZN(n16327) );
  OAI21_X1 U19318 ( .B1(n16328), .B2(n16373), .A(n16327), .ZN(U222) );
  INV_X1 U19319 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n16330) );
  AOI22_X1 U19320 ( .A1(P2_DATAO_REG_24__SCAN_IN), .A2(n16371), .B1(
        P1_DATAO_REG_24__SCAN_IN), .B2(n16370), .ZN(n16329) );
  OAI21_X1 U19321 ( .B1(n16330), .B2(n16373), .A(n16329), .ZN(U223) );
  AOI22_X1 U19322 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(n16371), .B1(
        P1_DATAO_REG_23__SCAN_IN), .B2(n16370), .ZN(n16331) );
  OAI21_X1 U19323 ( .B1(n16332), .B2(n16373), .A(n16331), .ZN(U224) );
  INV_X1 U19324 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n16334) );
  AOI22_X1 U19325 ( .A1(P2_DATAO_REG_22__SCAN_IN), .A2(n16371), .B1(
        P1_DATAO_REG_22__SCAN_IN), .B2(n16370), .ZN(n16333) );
  OAI21_X1 U19326 ( .B1(n16334), .B2(n16373), .A(n16333), .ZN(U225) );
  AOI22_X1 U19327 ( .A1(P2_DATAO_REG_21__SCAN_IN), .A2(n16371), .B1(
        P1_DATAO_REG_21__SCAN_IN), .B2(n16370), .ZN(n16335) );
  OAI21_X1 U19328 ( .B1(n16336), .B2(n16373), .A(n16335), .ZN(U226) );
  INV_X1 U19329 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n16338) );
  AOI22_X1 U19330 ( .A1(P2_DATAO_REG_20__SCAN_IN), .A2(n16371), .B1(
        P1_DATAO_REG_20__SCAN_IN), .B2(n16370), .ZN(n16337) );
  OAI21_X1 U19331 ( .B1(n16338), .B2(n16373), .A(n16337), .ZN(U227) );
  INV_X1 U19332 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n16340) );
  AOI22_X1 U19333 ( .A1(P2_DATAO_REG_19__SCAN_IN), .A2(n16371), .B1(
        P1_DATAO_REG_19__SCAN_IN), .B2(n16370), .ZN(n16339) );
  OAI21_X1 U19334 ( .B1(n16340), .B2(n16373), .A(n16339), .ZN(U228) );
  INV_X1 U19335 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n16342) );
  AOI22_X1 U19336 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(n16371), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n16370), .ZN(n16341) );
  OAI21_X1 U19337 ( .B1(n16342), .B2(n16373), .A(n16341), .ZN(U229) );
  INV_X1 U19338 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n16344) );
  AOI22_X1 U19339 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(n16371), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n16370), .ZN(n16343) );
  OAI21_X1 U19340 ( .B1(n16344), .B2(n16373), .A(n16343), .ZN(U230) );
  INV_X1 U19341 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n16346) );
  AOI22_X1 U19342 ( .A1(P2_DATAO_REG_16__SCAN_IN), .A2(n16371), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n16370), .ZN(n16345) );
  OAI21_X1 U19343 ( .B1(n16346), .B2(n16373), .A(n16345), .ZN(U231) );
  AOI22_X1 U19344 ( .A1(P2_DATAO_REG_15__SCAN_IN), .A2(n16371), .B1(
        P1_DATAO_REG_15__SCAN_IN), .B2(n16370), .ZN(n16347) );
  OAI21_X1 U19345 ( .B1(n13530), .B2(n16373), .A(n16347), .ZN(U232) );
  AOI22_X1 U19346 ( .A1(P2_DATAO_REG_14__SCAN_IN), .A2(n16371), .B1(
        P1_DATAO_REG_14__SCAN_IN), .B2(n16370), .ZN(n16348) );
  OAI21_X1 U19347 ( .B1(n14223), .B2(n16373), .A(n16348), .ZN(U233) );
  AOI22_X1 U19348 ( .A1(P2_DATAO_REG_13__SCAN_IN), .A2(n16371), .B1(
        P1_DATAO_REG_13__SCAN_IN), .B2(n16370), .ZN(n16349) );
  OAI21_X1 U19349 ( .B1(n14229), .B2(n16373), .A(n16349), .ZN(U234) );
  AOI22_X1 U19350 ( .A1(P2_DATAO_REG_12__SCAN_IN), .A2(n16371), .B1(
        P1_DATAO_REG_12__SCAN_IN), .B2(n16370), .ZN(n16350) );
  OAI21_X1 U19351 ( .B1(n21043), .B2(n16373), .A(n16350), .ZN(U235) );
  AOI22_X1 U19352 ( .A1(P2_DATAO_REG_11__SCAN_IN), .A2(n16371), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n16370), .ZN(n16351) );
  OAI21_X1 U19353 ( .B1(n13295), .B2(n16373), .A(n16351), .ZN(U236) );
  AOI22_X1 U19354 ( .A1(P2_DATAO_REG_10__SCAN_IN), .A2(n16371), .B1(
        P1_DATAO_REG_10__SCAN_IN), .B2(n16370), .ZN(n16352) );
  OAI21_X1 U19355 ( .B1(n16353), .B2(n16373), .A(n16352), .ZN(U237) );
  AOI22_X1 U19356 ( .A1(P2_DATAO_REG_9__SCAN_IN), .A2(n16371), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n16370), .ZN(n16354) );
  OAI21_X1 U19357 ( .B1(n13920), .B2(n16373), .A(n16354), .ZN(U238) );
  AOI22_X1 U19358 ( .A1(P2_DATAO_REG_8__SCAN_IN), .A2(n16371), .B1(
        P1_DATAO_REG_8__SCAN_IN), .B2(n16370), .ZN(n16355) );
  OAI21_X1 U19359 ( .B1(n13906), .B2(n16373), .A(n16355), .ZN(U239) );
  INV_X1 U19360 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n16357) );
  AOI22_X1 U19361 ( .A1(P2_DATAO_REG_7__SCAN_IN), .A2(n16371), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(n16370), .ZN(n16356) );
  OAI21_X1 U19362 ( .B1(n16357), .B2(n16373), .A(n16356), .ZN(U240) );
  AOI22_X1 U19363 ( .A1(P2_DATAO_REG_6__SCAN_IN), .A2(n16371), .B1(
        P1_DATAO_REG_6__SCAN_IN), .B2(n16370), .ZN(n16358) );
  OAI21_X1 U19364 ( .B1(n16359), .B2(n16373), .A(n16358), .ZN(U241) );
  INV_X1 U19365 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n16361) );
  AOI22_X1 U19366 ( .A1(P2_DATAO_REG_5__SCAN_IN), .A2(n16371), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(n16370), .ZN(n16360) );
  OAI21_X1 U19367 ( .B1(n16361), .B2(n16373), .A(n16360), .ZN(U242) );
  AOI22_X1 U19368 ( .A1(P2_DATAO_REG_4__SCAN_IN), .A2(n16371), .B1(
        P1_DATAO_REG_4__SCAN_IN), .B2(n16370), .ZN(n16362) );
  OAI21_X1 U19369 ( .B1(n16363), .B2(n16373), .A(n16362), .ZN(U243) );
  INV_X1 U19370 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n16365) );
  AOI22_X1 U19371 ( .A1(P2_DATAO_REG_3__SCAN_IN), .A2(n16371), .B1(
        P1_DATAO_REG_3__SCAN_IN), .B2(n16370), .ZN(n16364) );
  OAI21_X1 U19372 ( .B1(n16365), .B2(n16373), .A(n16364), .ZN(U244) );
  INV_X1 U19373 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n16367) );
  AOI22_X1 U19374 ( .A1(P2_DATAO_REG_2__SCAN_IN), .A2(n16371), .B1(
        P1_DATAO_REG_2__SCAN_IN), .B2(n16370), .ZN(n16366) );
  OAI21_X1 U19375 ( .B1(n16367), .B2(n16373), .A(n16366), .ZN(U245) );
  INV_X1 U19376 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n16369) );
  AOI22_X1 U19377 ( .A1(P2_DATAO_REG_1__SCAN_IN), .A2(n16371), .B1(
        P1_DATAO_REG_1__SCAN_IN), .B2(n16370), .ZN(n16368) );
  OAI21_X1 U19378 ( .B1(n16369), .B2(n16373), .A(n16368), .ZN(U246) );
  INV_X1 U19379 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n20865) );
  AOI22_X1 U19380 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(n16371), .B1(
        P1_DATAO_REG_0__SCAN_IN), .B2(n16370), .ZN(n16372) );
  OAI21_X1 U19381 ( .B1(n20865), .B2(n16373), .A(n16372), .ZN(U247) );
  OAI22_X1 U19382 ( .A1(U215), .A2(P2_DATAO_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n16405), .ZN(n16374) );
  INV_X1 U19383 ( .A(n16374), .ZN(U251) );
  OAI22_X1 U19384 ( .A1(U215), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n16405), .ZN(n16375) );
  INV_X1 U19385 ( .A(n16375), .ZN(U252) );
  OAI22_X1 U19386 ( .A1(U215), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n16405), .ZN(n16376) );
  INV_X1 U19387 ( .A(n16376), .ZN(U253) );
  OAI22_X1 U19388 ( .A1(U215), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n16405), .ZN(n16377) );
  INV_X1 U19389 ( .A(n16377), .ZN(U254) );
  OAI22_X1 U19390 ( .A1(U215), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n16405), .ZN(n16378) );
  INV_X1 U19391 ( .A(n16378), .ZN(U255) );
  OAI22_X1 U19392 ( .A1(U215), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n16405), .ZN(n16379) );
  INV_X1 U19393 ( .A(n16379), .ZN(U256) );
  OAI22_X1 U19394 ( .A1(U215), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n16405), .ZN(n16380) );
  INV_X1 U19395 ( .A(n16380), .ZN(U257) );
  OAI22_X1 U19396 ( .A1(U215), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n16405), .ZN(n16381) );
  INV_X1 U19397 ( .A(n16381), .ZN(U258) );
  OAI22_X1 U19398 ( .A1(U215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n16405), .ZN(n16382) );
  INV_X1 U19399 ( .A(n16382), .ZN(U259) );
  OAI22_X1 U19400 ( .A1(U215), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(
        BUF2_REG_9__SCAN_IN), .B2(n16397), .ZN(n16383) );
  INV_X1 U19401 ( .A(n16383), .ZN(U260) );
  OAI22_X1 U19402 ( .A1(U215), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n16397), .ZN(n16384) );
  INV_X1 U19403 ( .A(n16384), .ZN(U261) );
  OAI22_X1 U19404 ( .A1(U215), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n16405), .ZN(n16385) );
  INV_X1 U19405 ( .A(n16385), .ZN(U262) );
  OAI22_X1 U19406 ( .A1(U215), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n16397), .ZN(n16386) );
  INV_X1 U19407 ( .A(n16386), .ZN(U263) );
  OAI22_X1 U19408 ( .A1(U215), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n16405), .ZN(n16387) );
  INV_X1 U19409 ( .A(n16387), .ZN(U264) );
  OAI22_X1 U19410 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n16405), .ZN(n16388) );
  INV_X1 U19411 ( .A(n16388), .ZN(U265) );
  OAI22_X1 U19412 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n16397), .ZN(n16389) );
  INV_X1 U19413 ( .A(n16389), .ZN(U266) );
  OAI22_X1 U19414 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n16397), .ZN(n16390) );
  INV_X1 U19415 ( .A(n16390), .ZN(U267) );
  OAI22_X1 U19416 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n16397), .ZN(n16391) );
  INV_X1 U19417 ( .A(n16391), .ZN(U268) );
  OAI22_X1 U19418 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n16397), .ZN(n16392) );
  INV_X1 U19419 ( .A(n16392), .ZN(U269) );
  OAI22_X1 U19420 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n16397), .ZN(n16393) );
  INV_X1 U19421 ( .A(n16393), .ZN(U270) );
  OAI22_X1 U19422 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n16397), .ZN(n16394) );
  INV_X1 U19423 ( .A(n16394), .ZN(U271) );
  OAI22_X1 U19424 ( .A1(U215), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n16405), .ZN(n16395) );
  INV_X1 U19425 ( .A(n16395), .ZN(U272) );
  OAI22_X1 U19426 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n16405), .ZN(n16396) );
  INV_X1 U19427 ( .A(n16396), .ZN(U273) );
  OAI22_X1 U19428 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n16397), .ZN(n16398) );
  INV_X1 U19429 ( .A(n16398), .ZN(U274) );
  OAI22_X1 U19430 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n16405), .ZN(n16399) );
  INV_X1 U19431 ( .A(n16399), .ZN(U275) );
  OAI22_X1 U19432 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n16405), .ZN(n16400) );
  INV_X1 U19433 ( .A(n16400), .ZN(U276) );
  OAI22_X1 U19434 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n16405), .ZN(n16401) );
  INV_X1 U19435 ( .A(n16401), .ZN(U277) );
  OAI22_X1 U19436 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n16405), .ZN(n16402) );
  INV_X1 U19437 ( .A(n16402), .ZN(U278) );
  INV_X1 U19438 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n19100) );
  INV_X1 U19439 ( .A(BUF2_REG_28__SCAN_IN), .ZN(n18128) );
  AOI22_X1 U19440 ( .A1(n16405), .A2(n19100), .B1(n18128), .B2(U215), .ZN(U279) );
  OAI22_X1 U19441 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n16405), .ZN(n16403) );
  INV_X1 U19442 ( .A(n16403), .ZN(U280) );
  INV_X1 U19443 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n18138) );
  AOI22_X1 U19444 ( .A1(n16405), .A2(n19096), .B1(n18138), .B2(U215), .ZN(U281) );
  INV_X1 U19445 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n16404) );
  AOI22_X1 U19446 ( .A1(n16405), .A2(n19093), .B1(n16404), .B2(U215), .ZN(U282) );
  INV_X1 U19447 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n16407) );
  AOI222_X1 U19448 ( .A1(n16407), .A2(P3_DATAO_REG_30__SCAN_IN), .B1(n16406), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .C1(n19093), .C2(
        P2_DATAO_REG_30__SCAN_IN), .ZN(n16408) );
  INV_X2 U19449 ( .A(n16410), .ZN(n16409) );
  INV_X1 U19450 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n18664) );
  INV_X1 U19451 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n19738) );
  AOI22_X1 U19452 ( .A1(n16409), .A2(n18664), .B1(n19738), .B2(n16410), .ZN(
        U347) );
  INV_X1 U19453 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n18662) );
  INV_X1 U19454 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n19737) );
  AOI22_X1 U19455 ( .A1(n16409), .A2(n18662), .B1(n19737), .B2(n16410), .ZN(
        U348) );
  INV_X1 U19456 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n18659) );
  INV_X1 U19457 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n19735) );
  AOI22_X1 U19458 ( .A1(n16409), .A2(n18659), .B1(n19735), .B2(n16410), .ZN(
        U349) );
  INV_X1 U19459 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n18658) );
  INV_X1 U19460 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n19734) );
  AOI22_X1 U19461 ( .A1(n16409), .A2(n18658), .B1(n19734), .B2(n16410), .ZN(
        U350) );
  INV_X1 U19462 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n18656) );
  INV_X1 U19463 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n21025) );
  AOI22_X1 U19464 ( .A1(n16409), .A2(n18656), .B1(n21025), .B2(n16410), .ZN(
        U351) );
  INV_X1 U19465 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n18654) );
  INV_X1 U19466 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n19731) );
  AOI22_X1 U19467 ( .A1(n16409), .A2(n18654), .B1(n19731), .B2(n16410), .ZN(
        U352) );
  INV_X1 U19468 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n18652) );
  AOI22_X1 U19469 ( .A1(n16409), .A2(n18652), .B1(n19730), .B2(n16410), .ZN(
        U353) );
  INV_X1 U19470 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n18650) );
  INV_X1 U19471 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n20933) );
  AOI22_X1 U19472 ( .A1(n16409), .A2(n18650), .B1(n20933), .B2(n16410), .ZN(
        U354) );
  INV_X1 U19473 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n18705) );
  INV_X1 U19474 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n19774) );
  AOI22_X1 U19475 ( .A1(n16409), .A2(n18705), .B1(n19774), .B2(n16410), .ZN(
        U355) );
  INV_X1 U19476 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n18702) );
  INV_X1 U19477 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n19769) );
  AOI22_X1 U19478 ( .A1(n16409), .A2(n18702), .B1(n19769), .B2(n16410), .ZN(
        U356) );
  INV_X1 U19479 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n18699) );
  INV_X1 U19480 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n19767) );
  AOI22_X1 U19481 ( .A1(n16409), .A2(n18699), .B1(n19767), .B2(n16410), .ZN(
        U357) );
  INV_X1 U19482 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n18698) );
  INV_X1 U19483 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n19764) );
  AOI22_X1 U19484 ( .A1(n16409), .A2(n18698), .B1(n19764), .B2(n16410), .ZN(
        U358) );
  INV_X1 U19485 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n18696) );
  INV_X1 U19486 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n19763) );
  AOI22_X1 U19487 ( .A1(n16409), .A2(n18696), .B1(n19763), .B2(n16410), .ZN(
        U359) );
  INV_X1 U19488 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n18694) );
  INV_X1 U19489 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n19761) );
  AOI22_X1 U19490 ( .A1(n16409), .A2(n18694), .B1(n19761), .B2(n16410), .ZN(
        U360) );
  INV_X1 U19491 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n18692) );
  INV_X1 U19492 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n19759) );
  AOI22_X1 U19493 ( .A1(n16409), .A2(n18692), .B1(n19759), .B2(n16410), .ZN(
        U361) );
  INV_X1 U19494 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n18689) );
  INV_X1 U19495 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n19757) );
  AOI22_X1 U19496 ( .A1(n16409), .A2(n18689), .B1(n19757), .B2(n16410), .ZN(
        U362) );
  INV_X1 U19497 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n18688) );
  INV_X1 U19498 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n19755) );
  AOI22_X1 U19499 ( .A1(n16409), .A2(n18688), .B1(n19755), .B2(n16410), .ZN(
        U363) );
  INV_X1 U19500 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n18685) );
  INV_X1 U19501 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n19754) );
  AOI22_X1 U19502 ( .A1(n16409), .A2(n18685), .B1(n19754), .B2(n16410), .ZN(
        U364) );
  INV_X1 U19503 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n18648) );
  INV_X1 U19504 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n19727) );
  AOI22_X1 U19505 ( .A1(n16409), .A2(n18648), .B1(n19727), .B2(n16410), .ZN(
        U365) );
  INV_X1 U19506 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n18684) );
  INV_X1 U19507 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n19752) );
  AOI22_X1 U19508 ( .A1(n16409), .A2(n18684), .B1(n19752), .B2(n16410), .ZN(
        U366) );
  INV_X1 U19509 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n18682) );
  INV_X1 U19510 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n19751) );
  AOI22_X1 U19511 ( .A1(n16409), .A2(n18682), .B1(n19751), .B2(n16410), .ZN(
        U367) );
  INV_X1 U19512 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n18680) );
  INV_X1 U19513 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n19750) );
  AOI22_X1 U19514 ( .A1(n16409), .A2(n18680), .B1(n19750), .B2(n16410), .ZN(
        U368) );
  INV_X1 U19515 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n18677) );
  INV_X1 U19516 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n19749) );
  AOI22_X1 U19517 ( .A1(n16409), .A2(n18677), .B1(n19749), .B2(n16410), .ZN(
        U369) );
  INV_X1 U19518 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n18676) );
  INV_X1 U19519 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n19747) );
  AOI22_X1 U19520 ( .A1(n16409), .A2(n18676), .B1(n19747), .B2(n16410), .ZN(
        U370) );
  INV_X1 U19521 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n18674) );
  INV_X1 U19522 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n19745) );
  AOI22_X1 U19523 ( .A1(n16409), .A2(n18674), .B1(n19745), .B2(n16410), .ZN(
        U371) );
  INV_X1 U19524 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n18671) );
  INV_X1 U19525 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n19743) );
  AOI22_X1 U19526 ( .A1(n16409), .A2(n18671), .B1(n19743), .B2(n16410), .ZN(
        U372) );
  INV_X1 U19527 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n18670) );
  INV_X1 U19528 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n19741) );
  AOI22_X1 U19529 ( .A1(n16409), .A2(n18670), .B1(n19741), .B2(n16410), .ZN(
        U373) );
  INV_X1 U19530 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n18668) );
  INV_X1 U19531 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n20990) );
  AOI22_X1 U19532 ( .A1(n16409), .A2(n18668), .B1(n20990), .B2(n16410), .ZN(
        U374) );
  INV_X1 U19533 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n18666) );
  INV_X1 U19534 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n19739) );
  AOI22_X1 U19535 ( .A1(n16409), .A2(n18666), .B1(n19739), .B2(n16410), .ZN(
        U375) );
  INV_X1 U19536 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n18646) );
  INV_X1 U19537 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n19726) );
  AOI22_X1 U19538 ( .A1(n16409), .A2(n18646), .B1(n19726), .B2(n16410), .ZN(
        U376) );
  INV_X1 U19539 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n18645) );
  NAND2_X1 U19540 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n18645), .ZN(n18637) );
  OR2_X1 U19541 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(P3_STATE_REG_1__SCAN_IN), 
        .ZN(n18630) );
  OAI21_X1 U19542 ( .B1(n18642), .B2(n18637), .A(n18630), .ZN(n18713) );
  AOI21_X1 U19543 ( .B1(P3_STATE_REG_0__SCAN_IN), .B2(P3_ADS_N_REG_SCAN_IN), 
        .A(n18713), .ZN(n16411) );
  INV_X1 U19544 ( .A(n16411), .ZN(P3_U2633) );
  NAND2_X1 U19545 ( .A1(n18776), .A2(n18775), .ZN(n18781) );
  INV_X1 U19546 ( .A(n16416), .ZN(n16412) );
  OAI21_X1 U19547 ( .B1(n16412), .B2(n17345), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n16413) );
  OAI21_X1 U19548 ( .B1(n18781), .B2(n18764), .A(n16413), .ZN(P3_U2634) );
  AOI21_X1 U19549 ( .B1(n18642), .B2(n18645), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n16414) );
  AOI22_X1 U19550 ( .A1(n18772), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n16414), 
        .B2(n18773), .ZN(P3_U2635) );
  NOR2_X1 U19551 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n18628) );
  OAI21_X1 U19552 ( .B1(n18628), .B2(BS16), .A(n18713), .ZN(n18711) );
  OAI21_X1 U19553 ( .B1(n18713), .B2(n18621), .A(n18711), .ZN(P3_U2636) );
  AND3_X1 U19554 ( .A1(n16416), .A2(n18555), .A3(n16415), .ZN(n18558) );
  NOR2_X1 U19555 ( .A1(n18558), .A2(n18619), .ZN(n18756) );
  OAI21_X1 U19556 ( .B1(n18756), .B2(n18101), .A(n16417), .ZN(P3_U2637) );
  NOR4_X1 U19557 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_20__SCAN_IN), .A3(P3_DATAWIDTH_REG_21__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_22__SCAN_IN), .ZN(n16421) );
  NOR4_X1 U19558 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_15__SCAN_IN), .A3(P3_DATAWIDTH_REG_16__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_17__SCAN_IN), .ZN(n16420) );
  NOR4_X1 U19559 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_29__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n16419) );
  NOR4_X1 U19560 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_24__SCAN_IN), .A3(P3_DATAWIDTH_REG_25__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_26__SCAN_IN), .ZN(n16418) );
  NAND4_X1 U19561 ( .A1(n16421), .A2(n16420), .A3(n16419), .A4(n16418), .ZN(
        n16427) );
  NOR4_X1 U19562 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_3__SCAN_IN), .A3(P3_DATAWIDTH_REG_4__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_5__SCAN_IN), .ZN(n16425) );
  AOI211_X1 U19563 ( .C1(P3_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_27__SCAN_IN), .B(
        P3_DATAWIDTH_REG_18__SCAN_IN), .ZN(n16424) );
  NOR4_X1 U19564 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_11__SCAN_IN), .A3(P3_DATAWIDTH_REG_12__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_13__SCAN_IN), .ZN(n16423) );
  NOR4_X1 U19565 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_7__SCAN_IN), .A3(P3_DATAWIDTH_REG_8__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_9__SCAN_IN), .ZN(n16422) );
  NAND4_X1 U19566 ( .A1(n16425), .A2(n16424), .A3(n16423), .A4(n16422), .ZN(
        n16426) );
  NOR2_X1 U19567 ( .A1(n16427), .A2(n16426), .ZN(n18752) );
  INV_X1 U19568 ( .A(n18752), .ZN(n16430) );
  INV_X1 U19569 ( .A(P3_REIP_REG_0__SCAN_IN), .ZN(n20968) );
  NAND2_X1 U19570 ( .A1(n18752), .A2(n20968), .ZN(n18748) );
  NOR3_X1 U19571 ( .A1(P3_DATAWIDTH_REG_1__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A3(n18748), .ZN(n16429) );
  AOI221_X1 U19572 ( .B1(n16430), .B2(P3_BYTEENABLE_REG_1__SCAN_IN), .C1(
        n18752), .C2(P3_REIP_REG_1__SCAN_IN), .A(n16429), .ZN(n16428) );
  INV_X1 U19573 ( .A(n16428), .ZN(P3_U2638) );
  INV_X1 U19574 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n18749) );
  NAND2_X1 U19575 ( .A1(n18752), .A2(n18749), .ZN(n18753) );
  AOI21_X1 U19576 ( .B1(P3_BYTEENABLE_REG_3__SCAN_IN), .B2(n16430), .A(n16429), 
        .ZN(n16431) );
  OAI21_X1 U19577 ( .B1(P3_DATAWIDTH_REG_1__SCAN_IN), .B2(n18753), .A(n16431), 
        .ZN(P3_U2639) );
  NAND3_X1 U19578 ( .A1(n18764), .A2(n18775), .A3(n18621), .ZN(n16434) );
  NOR2_X2 U19579 ( .A1(n18726), .A2(n16434), .ZN(n16776) );
  NAND2_X1 U19580 ( .A1(n18775), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18491) );
  INV_X1 U19581 ( .A(n18491), .ZN(n18623) );
  NAND3_X1 U19582 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18623), .A3(n18726), 
        .ZN(n18617) );
  INV_X1 U19583 ( .A(n18768), .ZN(n18761) );
  AOI211_X1 U19584 ( .C1(n18117), .C2(n18758), .A(n18761), .B(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n16435) );
  AOI211_X4 U19585 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n18760), .A(n16435), .B(
        n18780), .ZN(n16783) );
  INV_X1 U19586 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n18706) );
  INV_X1 U19587 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n18700) );
  INV_X1 U19588 ( .A(n16435), .ZN(n18612) );
  INV_X1 U19589 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n18693) );
  INV_X1 U19590 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n18667) );
  INV_X1 U19591 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n18660) );
  INV_X1 U19592 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n18657) );
  INV_X1 U19593 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n18655) );
  INV_X1 U19594 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n18651) );
  NAND3_X1 U19595 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_3__SCAN_IN), 
        .A3(P3_REIP_REG_2__SCAN_IN), .ZN(n16751) );
  NOR2_X1 U19596 ( .A1(n18651), .A2(n16751), .ZN(n16735) );
  NAND2_X1 U19597 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(n16735), .ZN(n16733) );
  NOR4_X1 U19598 ( .A1(n18660), .A2(n18657), .A3(n18655), .A4(n16733), .ZN(
        n16678) );
  NAND4_X1 U19599 ( .A1(P3_REIP_REG_11__SCAN_IN), .A2(n16678), .A3(
        P3_REIP_REG_10__SCAN_IN), .A4(P3_REIP_REG_9__SCAN_IN), .ZN(n16661) );
  NOR2_X1 U19600 ( .A1(n18667), .A2(n16661), .ZN(n16643) );
  NAND3_X1 U19601 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(P3_REIP_REG_13__SCAN_IN), 
        .A3(n16643), .ZN(n16609) );
  NAND3_X1 U19602 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(P3_REIP_REG_16__SCAN_IN), 
        .A3(P3_REIP_REG_15__SCAN_IN), .ZN(n16545) );
  INV_X1 U19603 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n18686) );
  INV_X1 U19604 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n18683) );
  INV_X1 U19605 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n18681) );
  INV_X1 U19606 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n18679) );
  NOR3_X1 U19607 ( .A1(n18683), .A2(n18681), .A3(n18679), .ZN(n16546) );
  INV_X1 U19608 ( .A(n16546), .ZN(n16547) );
  NOR2_X1 U19609 ( .A1(n18686), .A2(n16547), .ZN(n16536) );
  NAND3_X1 U19610 ( .A1(P3_REIP_REG_23__SCAN_IN), .A2(n16536), .A3(
        P3_REIP_REG_22__SCAN_IN), .ZN(n16436) );
  NOR3_X1 U19611 ( .A1(n16609), .A2(n16545), .A3(n16436), .ZN(n16519) );
  NAND2_X1 U19612 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n16519), .ZN(n16510) );
  NOR2_X1 U19613 ( .A1(n18693), .A2(n16510), .ZN(n16496) );
  NAND2_X1 U19614 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(n16496), .ZN(n16447) );
  NOR2_X1 U19615 ( .A1(n16794), .A2(n16447), .ZN(n16478) );
  NAND2_X1 U19616 ( .A1(P3_REIP_REG_27__SCAN_IN), .A2(n16478), .ZN(n16487) );
  NOR2_X1 U19617 ( .A1(n18700), .A2(n16487), .ZN(n16472) );
  NAND2_X1 U19618 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n16472), .ZN(n16450) );
  NOR3_X1 U19619 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n18706), .A3(n16450), 
        .ZN(n16437) );
  AOI21_X1 U19620 ( .B1(n16783), .B2(P3_EBX_REG_31__SCAN_IN), .A(n16437), .ZN(
        n16453) );
  NAND2_X1 U19621 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n18760), .ZN(n16438) );
  AOI211_X4 U19622 ( .C1(n18621), .C2(n18768), .A(n18780), .B(n16438), .ZN(
        n16767) );
  NOR3_X1 U19623 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n16774) );
  INV_X1 U19624 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n17132) );
  NAND2_X1 U19625 ( .A1(n16774), .A2(n17132), .ZN(n16766) );
  NOR2_X1 U19626 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n16766), .ZN(n16746) );
  INV_X1 U19627 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n17123) );
  NAND2_X1 U19628 ( .A1(n16746), .A2(n17123), .ZN(n16741) );
  INV_X1 U19629 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n17119) );
  NAND2_X1 U19630 ( .A1(n16722), .A2(n17119), .ZN(n16715) );
  INV_X1 U19631 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n17066) );
  NAND2_X1 U19632 ( .A1(n16702), .A2(n17066), .ZN(n16693) );
  INV_X1 U19633 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n16673) );
  NAND2_X1 U19634 ( .A1(n16685), .A2(n16673), .ZN(n16672) );
  NAND2_X1 U19635 ( .A1(n16656), .A2(n16648), .ZN(n16647) );
  INV_X1 U19636 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n16998) );
  NAND2_X1 U19637 ( .A1(n16637), .A2(n16998), .ZN(n16626) );
  NAND2_X1 U19638 ( .A1(n16607), .A2(n16603), .ZN(n16602) );
  INV_X1 U19639 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n16577) );
  NAND2_X1 U19640 ( .A1(n16587), .A2(n16577), .ZN(n16575) );
  NAND2_X1 U19641 ( .A1(n16560), .A2(n16556), .ZN(n16555) );
  NAND2_X1 U19642 ( .A1(n16540), .A2(n16813), .ZN(n16532) );
  INV_X1 U19643 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n16514) );
  NAND2_X1 U19644 ( .A1(n16520), .A2(n16514), .ZN(n16513) );
  NOR2_X1 U19645 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16513), .ZN(n16497) );
  INV_X1 U19646 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n16493) );
  NAND2_X1 U19647 ( .A1(n16497), .A2(n16493), .ZN(n16492) );
  NOR2_X1 U19648 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16492), .ZN(n16476) );
  INV_X1 U19649 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n16847) );
  NAND2_X1 U19650 ( .A1(n16476), .A2(n16847), .ZN(n16455) );
  NOR2_X1 U19651 ( .A1(n16801), .A2(n16455), .ZN(n16461) );
  INV_X1 U19652 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n16818) );
  INV_X1 U19653 ( .A(n9891), .ZN(n16441) );
  NOR2_X1 U19654 ( .A1(n10010), .A2(n16441), .ZN(n16440) );
  OAI21_X1 U19655 ( .B1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n16440), .A(
        n16439), .ZN(n17424) );
  INV_X1 U19656 ( .A(n17424), .ZN(n16481) );
  AOI21_X1 U19657 ( .B1(n10010), .B2(n16441), .A(n16440), .ZN(n17431) );
  AOI21_X1 U19658 ( .B1(n17447), .B2(n17416), .A(n9891), .ZN(n17449) );
  NOR2_X1 U19659 ( .A1(n17473), .A2(n16443), .ZN(n16442) );
  OAI21_X1 U19660 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n16442), .A(
        n17416), .ZN(n17461) );
  INV_X1 U19661 ( .A(n17461), .ZN(n16508) );
  AOI21_X1 U19662 ( .B1(n17473), .B2(n16443), .A(n16442), .ZN(n17480) );
  INV_X1 U19663 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n16528) );
  NAND2_X1 U19664 ( .A1(n17492), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17458) );
  AOI21_X1 U19665 ( .B1(n16528), .B2(n17458), .A(n16444), .ZN(n17493) );
  NAND2_X1 U19666 ( .A1(n17528), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n16571) );
  INV_X1 U19667 ( .A(n16571), .ZN(n17498) );
  NAND2_X1 U19668 ( .A1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n17498), .ZN(
        n16446) );
  XNOR2_X1 U19669 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B(n16446), .ZN(
        n17514) );
  OAI21_X1 U19670 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17498), .A(
        n16446), .ZN(n17533) );
  INV_X1 U19671 ( .A(n17533), .ZN(n16564) );
  INV_X1 U19672 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n17774) );
  NOR2_X1 U19673 ( .A1(n17579), .A2(n17774), .ZN(n17578) );
  NAND2_X1 U19674 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17578), .ZN(
        n16620) );
  NOR2_X1 U19675 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n16620), .ZN(
        n16594) );
  INV_X1 U19676 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n20951) );
  INV_X1 U19677 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n16541) );
  INV_X1 U19678 ( .A(n17458), .ZN(n16445) );
  AOI221_X1 U19679 ( .B1(n20951), .B2(n16541), .C1(n16446), .C2(n16541), .A(
        n16445), .ZN(n17501) );
  NOR2_X1 U19680 ( .A1(n16521), .A2(n16713), .ZN(n16507) );
  NOR2_X1 U19681 ( .A1(n16508), .A2(n16507), .ZN(n16506) );
  NOR2_X1 U19682 ( .A1(n16488), .A2(n16713), .ZN(n16480) );
  NOR2_X1 U19683 ( .A1(n16481), .A2(n16480), .ZN(n16479) );
  NOR2_X1 U19684 ( .A1(n16479), .A2(n16713), .ZN(n16466) );
  NAND3_X1 U19685 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .ZN(n16449) );
  NAND2_X1 U19686 ( .A1(n16772), .A2(n16447), .ZN(n16448) );
  NAND2_X1 U19687 ( .A1(n16677), .A2(n16448), .ZN(n16477) );
  AOI21_X1 U19688 ( .B1(n16772), .B2(n16449), .A(n16477), .ZN(n16475) );
  NOR2_X1 U19689 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n16450), .ZN(n16459) );
  INV_X1 U19690 ( .A(n16459), .ZN(n16451) );
  AOI21_X1 U19691 ( .B1(n16475), .B2(n16451), .A(n18704), .ZN(n16452) );
  OAI211_X1 U19692 ( .C1(n16454), .C2(n16791), .A(n16453), .B(n9867), .ZN(
        P3_U2640) );
  NAND2_X1 U19693 ( .A1(n16767), .A2(n16455), .ZN(n16468) );
  XOR2_X1 U19694 ( .A(n16456), .B(n9882), .Z(n16460) );
  OAI22_X1 U19695 ( .A1(n16475), .A2(n18706), .B1(n16457), .B2(n16791), .ZN(
        n16458) );
  AOI211_X1 U19696 ( .C1(n16460), .C2(n16776), .A(n16459), .B(n16458), .ZN(
        n16463) );
  OAI21_X1 U19697 ( .B1(n16783), .B2(n16461), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n16462) );
  OAI211_X1 U19698 ( .C1(P3_EBX_REG_30__SCAN_IN), .C2(n16468), .A(n16463), .B(
        n16462), .ZN(P3_U2641) );
  AOI22_X1 U19699 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n16773), .B1(
        n16783), .B2(P3_EBX_REG_29__SCAN_IN), .ZN(n16474) );
  INV_X1 U19700 ( .A(n16464), .ZN(n16465) );
  AOI211_X1 U19701 ( .C1(n16467), .C2(n16466), .A(n16465), .B(n16793), .ZN(
        n16471) );
  INV_X1 U19702 ( .A(n16476), .ZN(n16469) );
  AOI21_X1 U19703 ( .B1(P3_EBX_REG_29__SCAN_IN), .B2(n16469), .A(n16468), .ZN(
        n16470) );
  AOI211_X1 U19704 ( .C1(n16472), .C2(n18701), .A(n16471), .B(n16470), .ZN(
        n16473) );
  OAI211_X1 U19705 ( .C1(n16475), .C2(n18701), .A(n16474), .B(n16473), .ZN(
        P3_U2642) );
  AOI22_X1 U19706 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n16773), .B1(
        n16783), .B2(P3_EBX_REG_28__SCAN_IN), .ZN(n16486) );
  AOI211_X1 U19707 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n16492), .A(n16476), .B(
        n16801), .ZN(n16484) );
  INV_X1 U19708 ( .A(n16477), .ZN(n16505) );
  INV_X1 U19709 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n18697) );
  NAND2_X1 U19710 ( .A1(n16478), .A2(n18697), .ZN(n16489) );
  AOI21_X1 U19711 ( .B1(n16505), .B2(n16489), .A(n18700), .ZN(n16483) );
  AOI211_X1 U19712 ( .C1(n16481), .C2(n16480), .A(n16479), .B(n16793), .ZN(
        n16482) );
  NOR3_X1 U19713 ( .A1(n16484), .A2(n16483), .A3(n16482), .ZN(n16485) );
  OAI211_X1 U19714 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n16487), .A(n16486), 
        .B(n16485), .ZN(P3_U2643) );
  AOI211_X1 U19715 ( .C1(n17431), .C2(n9843), .A(n16488), .B(n16793), .ZN(
        n16491) );
  OAI21_X1 U19716 ( .B1(n16791), .B2(n10010), .A(n16489), .ZN(n16490) );
  AOI211_X1 U19717 ( .C1(P3_EBX_REG_27__SCAN_IN), .C2(n16783), .A(n16491), .B(
        n16490), .ZN(n16495) );
  OAI211_X1 U19718 ( .C1(n16497), .C2(n16493), .A(n16767), .B(n16492), .ZN(
        n16494) );
  OAI211_X1 U19719 ( .C1(n16505), .C2(n18697), .A(n16495), .B(n16494), .ZN(
        P3_U2644) );
  AOI21_X1 U19720 ( .B1(n16772), .B2(n16496), .A(P3_REIP_REG_26__SCAN_IN), 
        .ZN(n16504) );
  AOI22_X1 U19721 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n16773), .B1(
        n16783), .B2(P3_EBX_REG_26__SCAN_IN), .ZN(n16503) );
  AOI211_X1 U19722 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n16513), .A(n16497), .B(
        n16801), .ZN(n16501) );
  AOI211_X1 U19723 ( .C1(n17449), .C2(n16499), .A(n16498), .B(n16793), .ZN(
        n16500) );
  NOR2_X1 U19724 ( .A1(n16501), .A2(n16500), .ZN(n16502) );
  OAI211_X1 U19725 ( .C1(n16505), .C2(n16504), .A(n16503), .B(n16502), .ZN(
        P3_U2645) );
  INV_X1 U19726 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n18691) );
  OAI21_X1 U19727 ( .B1(n16519), .B2(n16794), .A(n16677), .ZN(n16531) );
  AOI21_X1 U19728 ( .B1(n16772), .B2(n18691), .A(n16531), .ZN(n16517) );
  AOI211_X1 U19729 ( .C1(n16508), .C2(n16507), .A(n16506), .B(n16793), .ZN(
        n16512) );
  NAND2_X1 U19730 ( .A1(n16772), .A2(n18693), .ZN(n16509) );
  OAI22_X1 U19731 ( .A1(n17462), .A2(n16791), .B1(n16510), .B2(n16509), .ZN(
        n16511) );
  AOI211_X1 U19732 ( .C1(P3_EBX_REG_25__SCAN_IN), .C2(n16783), .A(n16512), .B(
        n16511), .ZN(n16516) );
  OAI211_X1 U19733 ( .C1(n16520), .C2(n16514), .A(n16767), .B(n16513), .ZN(
        n16515) );
  OAI211_X1 U19734 ( .C1(n16517), .C2(n18693), .A(n16516), .B(n16515), .ZN(
        P3_U2646) );
  NOR2_X1 U19735 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n16794), .ZN(n16518) );
  AOI22_X1 U19736 ( .A1(n16783), .A2(P3_EBX_REG_24__SCAN_IN), .B1(n16519), 
        .B2(n16518), .ZN(n16526) );
  AOI211_X1 U19737 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n16532), .A(n16520), .B(
        n16801), .ZN(n16524) );
  AOI211_X1 U19738 ( .C1(n17480), .C2(n16522), .A(n16521), .B(n16793), .ZN(
        n16523) );
  AOI211_X1 U19739 ( .C1(P3_REIP_REG_24__SCAN_IN), .C2(n16531), .A(n16524), 
        .B(n16523), .ZN(n16525) );
  OAI211_X1 U19740 ( .C1(n17473), .C2(n16791), .A(n16526), .B(n16525), .ZN(
        P3_U2647) );
  NAND4_X1 U19741 ( .A1(n16772), .A2(P3_REIP_REG_14__SCAN_IN), .A3(
        P3_REIP_REG_13__SCAN_IN), .A4(n16643), .ZN(n16619) );
  NAND3_X1 U19742 ( .A1(n16536), .A2(P3_REIP_REG_22__SCAN_IN), .A3(n16581), 
        .ZN(n16535) );
  AOI211_X1 U19743 ( .C1(n17493), .C2(n16527), .A(n9897), .B(n16793), .ZN(
        n16530) );
  OAI22_X1 U19744 ( .A1(n16528), .A2(n16791), .B1(n16802), .B2(n16813), .ZN(
        n16529) );
  AOI211_X1 U19745 ( .C1(P3_REIP_REG_23__SCAN_IN), .C2(n16531), .A(n16530), 
        .B(n16529), .ZN(n16534) );
  OAI211_X1 U19746 ( .C1(n16540), .C2(n16813), .A(n16767), .B(n16532), .ZN(
        n16533) );
  OAI211_X1 U19747 ( .C1(P3_REIP_REG_23__SCAN_IN), .C2(n16535), .A(n16534), 
        .B(n16533), .ZN(P3_U2648) );
  NAND2_X1 U19748 ( .A1(n16536), .A2(n16581), .ZN(n16550) );
  INV_X1 U19749 ( .A(n16537), .ZN(n16538) );
  AOI211_X1 U19750 ( .C1(n17501), .C2(n16539), .A(n16538), .B(n16793), .ZN(
        n16544) );
  AOI211_X1 U19751 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n16555), .A(n16540), .B(
        n16801), .ZN(n16543) );
  OAI22_X1 U19752 ( .A1(n16541), .A2(n16791), .B1(n16802), .B2(n16812), .ZN(
        n16542) );
  NOR3_X1 U19753 ( .A1(n16544), .A2(n16543), .A3(n16542), .ZN(n16549) );
  NOR3_X1 U19754 ( .A1(n16804), .A2(n16545), .A3(n16609), .ZN(n16570) );
  NOR2_X1 U19755 ( .A1(n16772), .A2(n16804), .ZN(n16809) );
  AOI21_X1 U19756 ( .B1(n16546), .B2(n16570), .A(n16809), .ZN(n16567) );
  INV_X1 U19757 ( .A(n16581), .ZN(n16592) );
  NOR3_X1 U19758 ( .A1(P3_REIP_REG_21__SCAN_IN), .A2(n16547), .A3(n16592), 
        .ZN(n16554) );
  OAI21_X1 U19759 ( .B1(n16567), .B2(n16554), .A(P3_REIP_REG_22__SCAN_IN), 
        .ZN(n16548) );
  OAI211_X1 U19760 ( .C1(P3_REIP_REG_22__SCAN_IN), .C2(n16550), .A(n16549), 
        .B(n16548), .ZN(P3_U2649) );
  AOI22_X1 U19761 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n16773), .B1(
        n16783), .B2(P3_EBX_REG_21__SCAN_IN), .ZN(n16559) );
  AOI211_X1 U19762 ( .C1(n17514), .C2(n16552), .A(n16551), .B(n16793), .ZN(
        n16553) );
  AOI211_X1 U19763 ( .C1(n16567), .C2(P3_REIP_REG_21__SCAN_IN), .A(n16554), 
        .B(n16553), .ZN(n16558) );
  OAI211_X1 U19764 ( .C1(n16560), .C2(n16556), .A(n16767), .B(n16555), .ZN(
        n16557) );
  NAND3_X1 U19765 ( .A1(n16559), .A2(n16558), .A3(n16557), .ZN(P3_U2650) );
  INV_X1 U19766 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n17530) );
  AOI211_X1 U19767 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n16575), .A(n16560), .B(
        n16801), .ZN(n16561) );
  AOI21_X1 U19768 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n16783), .A(n16561), .ZN(
        n16569) );
  NAND2_X1 U19769 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(P3_REIP_REG_18__SCAN_IN), 
        .ZN(n16580) );
  NOR2_X1 U19770 ( .A1(n16580), .A2(n16592), .ZN(n16566) );
  AOI211_X1 U19771 ( .C1(n16564), .C2(n16563), .A(n16562), .B(n16793), .ZN(
        n16565) );
  AOI221_X1 U19772 ( .B1(n16567), .B2(P3_REIP_REG_20__SCAN_IN), .C1(n16566), 
        .C2(n18683), .A(n16565), .ZN(n16568) );
  OAI211_X1 U19773 ( .C1(n17530), .C2(n16791), .A(n16569), .B(n16568), .ZN(
        P3_U2651) );
  OR2_X1 U19774 ( .A1(n16809), .A2(n16570), .ZN(n16597) );
  NAND3_X1 U19775 ( .A1(n17566), .A2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n16593) );
  INV_X1 U19776 ( .A(n16593), .ZN(n17544) );
  NAND2_X1 U19777 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n17544), .ZN(
        n16584) );
  INV_X1 U19778 ( .A(n16584), .ZN(n16572) );
  OAI21_X1 U19779 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n16572), .A(
        n16571), .ZN(n17549) );
  INV_X1 U19780 ( .A(n16594), .ZN(n16611) );
  OAI21_X1 U19781 ( .B1(n16584), .B2(n16611), .A(n16790), .ZN(n16574) );
  OAI21_X1 U19782 ( .B1(n17549), .B2(n16574), .A(n16776), .ZN(n16573) );
  AOI21_X1 U19783 ( .B1(n17549), .B2(n16574), .A(n16573), .ZN(n16579) );
  OAI211_X1 U19784 ( .C1(n16587), .C2(n16577), .A(n16767), .B(n16575), .ZN(
        n16576) );
  OAI211_X1 U19785 ( .C1(n16802), .C2(n16577), .A(n18091), .B(n16576), .ZN(
        n16578) );
  AOI211_X1 U19786 ( .C1(n16773), .C2(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n16579), .B(n16578), .ZN(n16583) );
  OAI211_X1 U19787 ( .C1(P3_REIP_REG_19__SCAN_IN), .C2(P3_REIP_REG_18__SCAN_IN), .A(n16581), .B(n16580), .ZN(n16582) );
  OAI211_X1 U19788 ( .C1(n16597), .C2(n18681), .A(n16583), .B(n16582), .ZN(
        P3_U2652) );
  OAI21_X1 U19789 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n17544), .A(
        n16584), .ZN(n17556) );
  OAI21_X1 U19790 ( .B1(n16593), .B2(n16611), .A(n16790), .ZN(n16586) );
  OAI21_X1 U19791 ( .B1(n17556), .B2(n16586), .A(n16776), .ZN(n16585) );
  AOI21_X1 U19792 ( .B1(n17556), .B2(n16586), .A(n16585), .ZN(n16590) );
  AOI211_X1 U19793 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n16602), .A(n16587), .B(
        n16801), .ZN(n16589) );
  INV_X1 U19794 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n17559) );
  OAI22_X1 U19795 ( .A1(n17559), .A2(n16791), .B1(n16802), .B2(n16945), .ZN(
        n16588) );
  NOR4_X1 U19796 ( .A1(n18093), .A2(n16590), .A3(n16589), .A4(n16588), .ZN(
        n16591) );
  OAI221_X1 U19797 ( .B1(P3_REIP_REG_18__SCAN_IN), .B2(n16592), .C1(n18679), 
        .C2(n16597), .A(n16591), .ZN(P3_U2653) );
  AOI22_X1 U19798 ( .A1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n16773), .B1(
        n16783), .B2(P3_EBX_REG_17__SCAN_IN), .ZN(n16606) );
  AND2_X1 U19799 ( .A1(n17566), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n16610) );
  OAI21_X1 U19800 ( .B1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n16610), .A(
        n16593), .ZN(n17571) );
  AOI21_X1 U19801 ( .B1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n16594), .A(
        n16713), .ZN(n16595) );
  XNOR2_X1 U19802 ( .A(n17571), .B(n16595), .ZN(n16601) );
  NAND2_X1 U19803 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(P3_REIP_REG_15__SCAN_IN), 
        .ZN(n16596) );
  NOR2_X1 U19804 ( .A1(n16596), .A2(n16619), .ZN(n16599) );
  INV_X1 U19805 ( .A(n16597), .ZN(n16598) );
  MUX2_X1 U19806 ( .A(n16599), .B(n16598), .S(P3_REIP_REG_17__SCAN_IN), .Z(
        n16600) );
  AOI21_X1 U19807 ( .B1(n16601), .B2(n16776), .A(n16600), .ZN(n16605) );
  OAI211_X1 U19808 ( .C1(n16607), .C2(n16603), .A(n16767), .B(n16602), .ZN(
        n16604) );
  NAND4_X1 U19809 ( .A1(n16606), .A2(n16605), .A3(n18091), .A4(n16604), .ZN(
        P3_U2654) );
  INV_X1 U19810 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n16618) );
  AOI211_X1 U19811 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n16626), .A(n16607), .B(
        n16801), .ZN(n16608) );
  AOI211_X1 U19812 ( .C1(n16783), .C2(P3_EBX_REG_16__SCAN_IN), .A(n18093), .B(
        n16608), .ZN(n16617) );
  NOR2_X1 U19813 ( .A1(n16804), .A2(n16609), .ZN(n16635) );
  AOI21_X1 U19814 ( .B1(P3_REIP_REG_15__SCAN_IN), .B2(n16635), .A(n16809), 
        .ZN(n16625) );
  AOI21_X1 U19815 ( .B1(n16618), .B2(n16620), .A(n16610), .ZN(n16613) );
  NAND2_X1 U19816 ( .A1(n16611), .A2(n16790), .ZN(n16612) );
  INV_X1 U19817 ( .A(n16612), .ZN(n16627) );
  INV_X1 U19818 ( .A(n16613), .ZN(n17584) );
  AOI221_X1 U19819 ( .B1(n16613), .B2(n16627), .C1(n17584), .C2(n16612), .A(
        n16793), .ZN(n16615) );
  INV_X1 U19820 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n18673) );
  NOR3_X1 U19821 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(n18673), .A3(n16619), 
        .ZN(n16614) );
  AOI211_X1 U19822 ( .C1(P3_REIP_REG_16__SCAN_IN), .C2(n16625), .A(n16615), 
        .B(n16614), .ZN(n16616) );
  OAI211_X1 U19823 ( .C1(n16618), .C2(n16791), .A(n16617), .B(n16616), .ZN(
        P3_U2655) );
  NAND2_X1 U19824 ( .A1(n18673), .A2(n16619), .ZN(n16624) );
  OAI21_X1 U19825 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n17578), .A(
        n16620), .ZN(n17590) );
  AOI21_X1 U19826 ( .B1(n16790), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n16793), .ZN(n16797) );
  INV_X1 U19827 ( .A(n16797), .ZN(n16621) );
  AOI211_X1 U19828 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(n16790), .A(
        n17590), .B(n16621), .ZN(n16623) );
  INV_X1 U19829 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17594) );
  OAI22_X1 U19830 ( .A1(n17594), .A2(n16791), .B1(n16802), .B2(n16998), .ZN(
        n16622) );
  AOI211_X1 U19831 ( .C1(n16625), .C2(n16624), .A(n16623), .B(n16622), .ZN(
        n16630) );
  OAI211_X1 U19832 ( .C1(n16637), .C2(n16998), .A(n16767), .B(n16626), .ZN(
        n16629) );
  NAND3_X1 U19833 ( .A1(n16776), .A2(n16627), .A3(n17590), .ZN(n16628) );
  NAND4_X1 U19834 ( .A1(n16630), .A2(n18091), .A3(n16629), .A4(n16628), .ZN(
        P3_U2656) );
  INV_X1 U19835 ( .A(n16631), .ZN(n17602) );
  NOR2_X1 U19836 ( .A1(n17774), .A2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n16777) );
  INV_X1 U19837 ( .A(n16777), .ZN(n16760) );
  NOR3_X1 U19838 ( .A1(n17602), .A2(n16632), .A3(n16760), .ZN(n16646) );
  NOR2_X1 U19839 ( .A1(n16646), .A2(n16713), .ZN(n16634) );
  NAND2_X1 U19840 ( .A1(n16631), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17619) );
  NOR2_X1 U19841 ( .A1(n16632), .A2(n17619), .ZN(n16644) );
  INV_X1 U19842 ( .A(n17578), .ZN(n16633) );
  OAI21_X1 U19843 ( .B1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n16644), .A(
        n16633), .ZN(n17605) );
  XOR2_X1 U19844 ( .A(n16634), .B(n17605), .Z(n16642) );
  AOI21_X1 U19845 ( .B1(n16783), .B2(P3_EBX_REG_14__SCAN_IN), .A(n18093), .ZN(
        n16641) );
  INV_X1 U19846 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n18672) );
  NAND3_X1 U19847 ( .A1(n16772), .A2(P3_REIP_REG_13__SCAN_IN), .A3(n16643), 
        .ZN(n16636) );
  AOI211_X1 U19848 ( .C1(n18672), .C2(n16636), .A(n16635), .B(n16809), .ZN(
        n16639) );
  AOI211_X1 U19849 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n16647), .A(n16637), .B(
        n16801), .ZN(n16638) );
  AOI211_X1 U19850 ( .C1(n16773), .C2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n16639), .B(n16638), .ZN(n16640) );
  OAI211_X1 U19851 ( .C1(n16793), .C2(n16642), .A(n16641), .B(n16640), .ZN(
        P3_U2657) );
  INV_X1 U19852 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n18669) );
  AOI21_X1 U19853 ( .B1(n16772), .B2(n16661), .A(n16804), .ZN(n16670) );
  NAND2_X1 U19854 ( .A1(n16772), .A2(n18667), .ZN(n16660) );
  AND2_X1 U19855 ( .A1(n16772), .A2(n16643), .ZN(n16654) );
  INV_X1 U19856 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17620) );
  INV_X1 U19857 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n17634) );
  NOR2_X1 U19858 ( .A1(n17634), .A2(n17619), .ZN(n16658) );
  INV_X1 U19859 ( .A(n16658), .ZN(n16645) );
  AOI21_X1 U19860 ( .B1(n17620), .B2(n16645), .A(n16644), .ZN(n17625) );
  NOR4_X1 U19861 ( .A1(n17625), .A2(n16646), .A3(n16793), .A4(n16713), .ZN(
        n16653) );
  AOI22_X1 U19862 ( .A1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n16773), .B1(
        n16783), .B2(P3_EBX_REG_13__SCAN_IN), .ZN(n16651) );
  OAI211_X1 U19863 ( .C1(n16658), .C2(n16713), .A(n17625), .B(n16797), .ZN(
        n16650) );
  OAI211_X1 U19864 ( .C1(n16656), .C2(n16648), .A(n16767), .B(n16647), .ZN(
        n16649) );
  NAND4_X1 U19865 ( .A1(n16651), .A2(n18091), .A3(n16650), .A4(n16649), .ZN(
        n16652) );
  AOI211_X1 U19866 ( .C1(n16654), .C2(n18669), .A(n16653), .B(n16652), .ZN(
        n16655) );
  OAI221_X1 U19867 ( .B1(n18669), .B2(n16670), .C1(n18669), .C2(n16660), .A(
        n16655), .ZN(P3_U2658) );
  AOI211_X1 U19868 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n16672), .A(n16656), .B(
        n16801), .ZN(n16657) );
  AOI21_X1 U19869 ( .B1(P3_EBX_REG_12__SCAN_IN), .B2(n16783), .A(n16657), .ZN(
        n16665) );
  AOI21_X1 U19870 ( .B1(n17634), .B2(n17619), .A(n16658), .ZN(n17637) );
  OAI21_X1 U19871 ( .B1(n17602), .B2(n16760), .A(n16790), .ZN(n16659) );
  XNOR2_X1 U19872 ( .A(n17637), .B(n16659), .ZN(n16663) );
  OAI22_X1 U19873 ( .A1(n17634), .A2(n16791), .B1(n16661), .B2(n16660), .ZN(
        n16662) );
  AOI211_X1 U19874 ( .C1(n16776), .C2(n16663), .A(n18093), .B(n16662), .ZN(
        n16664) );
  OAI211_X1 U19875 ( .C1(n16670), .C2(n18667), .A(n16665), .B(n16664), .ZN(
        P3_U2659) );
  INV_X1 U19876 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n18663) );
  INV_X1 U19877 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n18661) );
  NOR2_X1 U19878 ( .A1(n18663), .A2(n18661), .ZN(n16684) );
  NAND2_X1 U19879 ( .A1(n16772), .A2(n16678), .ZN(n16695) );
  INV_X1 U19880 ( .A(n16695), .ZN(n16666) );
  AOI21_X1 U19881 ( .B1(n16684), .B2(n16666), .A(P3_REIP_REG_11__SCAN_IN), 
        .ZN(n16669) );
  NOR2_X1 U19882 ( .A1(n17711), .A2(n17774), .ZN(n16736) );
  NAND2_X1 U19883 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n16736), .ZN(
        n16724) );
  NOR2_X1 U19884 ( .A1(n16667), .A2(n16724), .ZN(n16679) );
  OAI21_X1 U19885 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n16679), .A(
        n17619), .ZN(n17647) );
  OAI21_X1 U19886 ( .B1(n17646), .B2(n16760), .A(n16790), .ZN(n16682) );
  XNOR2_X1 U19887 ( .A(n17647), .B(n16682), .ZN(n16668) );
  OAI22_X1 U19888 ( .A1(n16670), .A2(n16669), .B1(n16793), .B2(n16668), .ZN(
        n16671) );
  AOI211_X1 U19889 ( .C1(n16783), .C2(P3_EBX_REG_11__SCAN_IN), .A(n18093), .B(
        n16671), .ZN(n16675) );
  OAI211_X1 U19890 ( .C1(n16685), .C2(n16673), .A(n16767), .B(n16672), .ZN(
        n16674) );
  OAI211_X1 U19891 ( .C1(n16791), .C2(n16676), .A(n16675), .B(n16674), .ZN(
        P3_U2660) );
  OAI21_X1 U19892 ( .B1(n16794), .B2(n16678), .A(n16677), .ZN(n16706) );
  INV_X1 U19893 ( .A(n16706), .ZN(n16691) );
  AOI22_X1 U19894 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n16773), .B1(
        n16783), .B2(P3_EBX_REG_10__SCAN_IN), .ZN(n16690) );
  AND3_X1 U19895 ( .A1(n17684), .A2(n17685), .A3(n16777), .ZN(n16699) );
  AOI21_X1 U19896 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n16699), .A(
        n16713), .ZN(n16698) );
  INV_X1 U19897 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n17673) );
  NAND2_X1 U19898 ( .A1(n17684), .A2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17686) );
  NOR2_X1 U19899 ( .A1(n17774), .A2(n17686), .ZN(n16712) );
  NAND2_X1 U19900 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n16712), .ZN(
        n16704) );
  NOR2_X1 U19901 ( .A1(n17673), .A2(n16704), .ZN(n16681) );
  INV_X1 U19902 ( .A(n16679), .ZN(n16680) );
  OAI21_X1 U19903 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n16681), .A(
        n16680), .ZN(n17660) );
  INV_X1 U19904 ( .A(n17660), .ZN(n16683) );
  AOI221_X1 U19905 ( .B1(n16698), .B2(n16683), .C1(n16682), .C2(n17660), .A(
        n16793), .ZN(n16688) );
  AOI211_X1 U19906 ( .C1(n18663), .C2(n18661), .A(n16684), .B(n16695), .ZN(
        n16687) );
  AOI211_X1 U19907 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n16693), .A(n16685), .B(
        n16801), .ZN(n16686) );
  NOR4_X1 U19908 ( .A1(n18093), .A2(n16688), .A3(n16687), .A4(n16686), .ZN(
        n16689) );
  OAI211_X1 U19909 ( .C1(n16691), .C2(n18663), .A(n16690), .B(n16689), .ZN(
        P3_U2661) );
  NAND2_X1 U19910 ( .A1(n16713), .A2(n16776), .ZN(n16780) );
  INV_X1 U19911 ( .A(n16704), .ZN(n16692) );
  AOI22_X1 U19912 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n16704), .B1(
        n16692), .B2(n17673), .ZN(n17675) );
  OAI22_X1 U19913 ( .A1(n17673), .A2(n16791), .B1(n16802), .B2(n17066), .ZN(
        n16697) );
  OAI211_X1 U19914 ( .C1(n16702), .C2(n17066), .A(n16767), .B(n16693), .ZN(
        n16694) );
  OAI211_X1 U19915 ( .C1(P3_REIP_REG_9__SCAN_IN), .C2(n16695), .A(n18091), .B(
        n16694), .ZN(n16696) );
  AOI211_X1 U19916 ( .C1(P3_REIP_REG_9__SCAN_IN), .C2(n16706), .A(n16697), .B(
        n16696), .ZN(n16701) );
  OAI211_X1 U19917 ( .C1(n16699), .C2(n17675), .A(n16776), .B(n16698), .ZN(
        n16700) );
  OAI211_X1 U19918 ( .C1(n16780), .C2(n17675), .A(n16701), .B(n16700), .ZN(
        P3_U2662) );
  AOI211_X1 U19919 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n16715), .A(n16702), .B(
        n16801), .ZN(n16703) );
  AOI211_X1 U19920 ( .C1(n16783), .C2(P3_EBX_REG_8__SCAN_IN), .A(n18093), .B(
        n16703), .ZN(n16711) );
  OAI21_X1 U19921 ( .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n16712), .A(
        n16704), .ZN(n17688) );
  INV_X1 U19922 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n16803) );
  AOI21_X1 U19923 ( .B1(n16712), .B2(n16803), .A(n16713), .ZN(n16705) );
  XNOR2_X1 U19924 ( .A(n17688), .B(n16705), .ZN(n16709) );
  NOR2_X1 U19925 ( .A1(n16794), .A2(n16733), .ZN(n16730) );
  NAND2_X1 U19926 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n16730), .ZN(n16721) );
  NOR2_X1 U19927 ( .A1(n18657), .A2(n16721), .ZN(n16707) );
  MUX2_X1 U19928 ( .A(n16707), .B(n16706), .S(P3_REIP_REG_8__SCAN_IN), .Z(
        n16708) );
  AOI21_X1 U19929 ( .B1(n16709), .B2(n16776), .A(n16708), .ZN(n16710) );
  OAI211_X1 U19930 ( .C1(n17687), .C2(n16791), .A(n16711), .B(n16710), .ZN(
        P3_U2663) );
  AOI221_X1 U19931 ( .B1(n18655), .B2(n16772), .C1(n16733), .C2(n16772), .A(
        n16804), .ZN(n16720) );
  AOI21_X1 U19932 ( .B1(n17702), .B2(n16724), .A(n16712), .ZN(n17708) );
  AOI21_X1 U19933 ( .B1(n17684), .B2(n16777), .A(n16713), .ZN(n16725) );
  OAI21_X1 U19934 ( .B1(n17708), .B2(n16725), .A(n16776), .ZN(n16714) );
  AOI21_X1 U19935 ( .B1(n17708), .B2(n16725), .A(n16714), .ZN(n16718) );
  OAI211_X1 U19936 ( .C1(n16722), .C2(n17119), .A(n16767), .B(n16715), .ZN(
        n16716) );
  OAI211_X1 U19937 ( .C1(n16802), .C2(n17119), .A(n18091), .B(n16716), .ZN(
        n16717) );
  AOI211_X1 U19938 ( .C1(n16773), .C2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n16718), .B(n16717), .ZN(n16719) );
  OAI221_X1 U19939 ( .B1(P3_REIP_REG_7__SCAN_IN), .B2(n16721), .C1(n18657), 
        .C2(n16720), .A(n16719), .ZN(P3_U2664) );
  AOI211_X1 U19940 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n16741), .A(n16722), .B(
        n16801), .ZN(n16723) );
  AOI211_X1 U19941 ( .C1(n16783), .C2(P3_EBX_REG_6__SCAN_IN), .A(n18093), .B(
        n16723), .ZN(n16732) );
  OAI21_X1 U19942 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n16736), .A(
        n16724), .ZN(n17717) );
  AND3_X1 U19943 ( .A1(n16776), .A2(n16725), .A3(n17717), .ZN(n16729) );
  AOI21_X1 U19944 ( .B1(n16772), .B2(n16733), .A(n16804), .ZN(n16738) );
  INV_X1 U19945 ( .A(n16780), .ZN(n16726) );
  OAI21_X1 U19946 ( .B1(n16736), .B2(n16726), .A(n16797), .ZN(n16727) );
  OAI22_X1 U19947 ( .A1(n16738), .A2(n18655), .B1(n17717), .B2(n16727), .ZN(
        n16728) );
  AOI211_X1 U19948 ( .C1(n16730), .C2(n18655), .A(n16729), .B(n16728), .ZN(
        n16731) );
  OAI211_X1 U19949 ( .C1(n17722), .C2(n16791), .A(n16732), .B(n16731), .ZN(
        P3_U2665) );
  AOI22_X1 U19950 ( .A1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n16773), .B1(
        n16783), .B2(P3_EBX_REG_5__SCAN_IN), .ZN(n16745) );
  AND2_X1 U19951 ( .A1(n16733), .A2(n16772), .ZN(n16734) );
  AOI21_X1 U19952 ( .B1(n16735), .B2(n16734), .A(n18093), .ZN(n16744) );
  INV_X1 U19953 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n16737) );
  NAND2_X1 U19954 ( .A1(n17726), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n16747) );
  AOI21_X1 U19955 ( .B1(n16737), .B2(n16747), .A(n16736), .ZN(n17732) );
  OAI21_X1 U19956 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16747), .A(
        n16790), .ZN(n16748) );
  XNOR2_X1 U19957 ( .A(n17732), .B(n16748), .ZN(n16740) );
  INV_X1 U19958 ( .A(n16738), .ZN(n16739) );
  AOI22_X1 U19959 ( .A1(n16776), .A2(n16740), .B1(P3_REIP_REG_5__SCAN_IN), 
        .B2(n16739), .ZN(n16743) );
  OAI211_X1 U19960 ( .C1(n16746), .C2(n17123), .A(n16767), .B(n16741), .ZN(
        n16742) );
  NAND4_X1 U19961 ( .A1(n16745), .A2(n16744), .A3(n16743), .A4(n16742), .ZN(
        P3_U2666) );
  AOI21_X1 U19962 ( .B1(n16772), .B2(n16751), .A(n16804), .ZN(n16761) );
  AOI211_X1 U19963 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n16766), .A(n16746), .B(
        n16801), .ZN(n16757) );
  NOR2_X1 U19964 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n17734), .ZN(
        n17746) );
  NOR2_X1 U19965 ( .A1(n17734), .A2(n17774), .ZN(n16759) );
  OAI21_X1 U19966 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n16759), .A(
        n16747), .ZN(n17743) );
  INV_X1 U19967 ( .A(n17743), .ZN(n16749) );
  AOI22_X1 U19968 ( .A1(n16749), .A2(n16790), .B1(n16748), .B2(n17743), .ZN(
        n16750) );
  AOI21_X1 U19969 ( .B1(n17746), .B2(n16777), .A(n16750), .ZN(n16755) );
  NOR2_X1 U19970 ( .A1(n17308), .A2(n18777), .ZN(n16807) );
  INV_X1 U19971 ( .A(n16807), .ZN(n16762) );
  AOI21_X1 U19972 ( .B1(n10222), .B2(n18561), .A(n16762), .ZN(n16753) );
  NOR3_X1 U19973 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n16794), .A3(n16751), .ZN(
        n16752) );
  AOI211_X1 U19974 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n16783), .A(n16753), .B(
        n16752), .ZN(n16754) );
  OAI211_X1 U19975 ( .C1(n16755), .C2(n16793), .A(n16754), .B(n18091), .ZN(
        n16756) );
  AOI211_X1 U19976 ( .C1(n16773), .C2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n16757), .B(n16756), .ZN(n16758) );
  OAI21_X1 U19977 ( .B1(n18651), .B2(n16761), .A(n16758), .ZN(P3_U2667) );
  INV_X1 U19978 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n16770) );
  NAND2_X1 U19979 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n16775) );
  AOI21_X1 U19980 ( .B1(n16770), .B2(n16775), .A(n16759), .ZN(n17756) );
  INV_X1 U19981 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17767) );
  OAI21_X1 U19982 ( .B1(n17767), .B2(n16760), .A(n16790), .ZN(n16779) );
  XNOR2_X1 U19983 ( .A(n17756), .B(n16779), .ZN(n16765) );
  INV_X1 U19984 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n18649) );
  NAND2_X1 U19985 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_2__SCAN_IN), 
        .ZN(n16771) );
  AOI221_X1 U19986 ( .B1(n16794), .B2(n18649), .C1(n16771), .C2(n18649), .A(
        n16761), .ZN(n16764) );
  NOR2_X1 U19987 ( .A1(n18739), .A2(n18732), .ZN(n18573) );
  AND2_X1 U19988 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18573), .ZN(
        n18572) );
  OAI21_X1 U19989 ( .B1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n18572), .A(
        n10222), .ZN(n18717) );
  OAI22_X1 U19990 ( .A1(n16802), .A2(n17132), .B1(n18717), .B2(n16762), .ZN(
        n16763) );
  AOI211_X1 U19991 ( .C1(n16776), .C2(n16765), .A(n16764), .B(n16763), .ZN(
        n16769) );
  OAI211_X1 U19992 ( .C1(n16774), .C2(n17132), .A(n16767), .B(n16766), .ZN(
        n16768) );
  OAI211_X1 U19993 ( .C1(n16791), .C2(n16770), .A(n16769), .B(n16768), .ZN(
        P3_U2668) );
  NOR2_X1 U19994 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_2__SCAN_IN), 
        .ZN(n16787) );
  AOI22_X1 U19995 ( .A1(n16772), .A2(n16771), .B1(P3_REIP_REG_2__SCAN_IN), 
        .B2(n16804), .ZN(n16786) );
  AOI21_X1 U19996 ( .B1(n18576), .B2(n18732), .A(n18572), .ZN(n18729) );
  AOI22_X1 U19997 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n16773), .B1(
        n18729), .B2(n16807), .ZN(n16785) );
  INV_X1 U19998 ( .A(P3_EBX_REG_0__SCAN_IN), .ZN(n16800) );
  INV_X1 U19999 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n17147) );
  NAND2_X1 U20000 ( .A1(n16800), .A2(n17147), .ZN(n16788) );
  AOI211_X1 U20001 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n16788), .A(n16774), .B(
        n16801), .ZN(n16782) );
  OAI21_X1 U20002 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A(n16775), .ZN(n17764) );
  OAI21_X1 U20003 ( .B1(n16777), .B2(n17764), .A(n16776), .ZN(n16778) );
  OAI22_X1 U20004 ( .A1(n17764), .A2(n16780), .B1(n16779), .B2(n16778), .ZN(
        n16781) );
  AOI211_X1 U20005 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n16783), .A(n16782), .B(
        n16781), .ZN(n16784) );
  OAI211_X1 U20006 ( .C1(n16787), .C2(n16786), .A(n16785), .B(n16784), .ZN(
        P3_U2669) );
  NAND2_X1 U20007 ( .A1(n16788), .A2(n17131), .ZN(n17148) );
  NAND2_X1 U20008 ( .A1(n18576), .A2(n16789), .ZN(n18591) );
  INV_X1 U20009 ( .A(n18591), .ZN(n18736) );
  AOI22_X1 U20010 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n16804), .B1(n18736), 
        .B2(n16807), .ZN(n16799) );
  NAND2_X1 U20011 ( .A1(n16790), .A2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n16792) );
  OAI21_X1 U20012 ( .B1(n16793), .B2(n16792), .A(n16791), .ZN(n16796) );
  OAI22_X1 U20013 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n16794), .B1(n17147), 
        .B2(n16802), .ZN(n16795) );
  AOI221_X1 U20014 ( .B1(n16797), .B2(n17774), .C1(n16796), .C2(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A(n16795), .ZN(n16798) );
  OAI211_X1 U20015 ( .C1(n16801), .C2(n17148), .A(n16799), .B(n16798), .ZN(
        P3_U2670) );
  AOI21_X1 U20016 ( .B1(n16802), .B2(n16801), .A(n16800), .ZN(n16806) );
  NOR3_X1 U20017 ( .A1(n18776), .A2(n16804), .A3(n16803), .ZN(n16805) );
  AOI211_X1 U20018 ( .C1(n16807), .C2(n18745), .A(n16806), .B(n16805), .ZN(
        n16808) );
  OAI21_X1 U20019 ( .B1(n16809), .B2(n20968), .A(n16808), .ZN(P3_U2671) );
  INV_X1 U20020 ( .A(P3_EBX_REG_20__SCAN_IN), .ZN(n16810) );
  NOR2_X1 U20021 ( .A1(n16810), .A2(n16929), .ZN(n16888) );
  NAND4_X1 U20022 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .A3(P3_EBX_REG_24__SCAN_IN), .A4(P3_EBX_REG_21__SCAN_IN), .ZN(n16811)
         );
  NOR4_X1 U20023 ( .A1(n16847), .A2(n16813), .A3(n16812), .A4(n16811), .ZN(
        n16814) );
  NAND4_X1 U20024 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(P3_EBX_REG_25__SCAN_IN), 
        .A3(n16888), .A4(n16814), .ZN(n16817) );
  NOR2_X1 U20025 ( .A1(n16818), .A2(n16817), .ZN(n16843) );
  NAND2_X1 U20026 ( .A1(n16963), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n16816) );
  NAND2_X1 U20027 ( .A1(n16843), .A2(n18145), .ZN(n16815) );
  OAI22_X1 U20028 ( .A1(n16843), .A2(n16816), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n16815), .ZN(P3_U2672) );
  NAND2_X1 U20029 ( .A1(n16818), .A2(n16817), .ZN(n16819) );
  NAND2_X1 U20030 ( .A1(n16819), .A2(n17141), .ZN(n16842) );
  AOI22_X1 U20031 ( .A1(n17103), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n16830) );
  INV_X1 U20032 ( .A(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n16822) );
  AOI22_X1 U20033 ( .A1(n17095), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17083), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n16821) );
  AOI22_X1 U20034 ( .A1(n17002), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17100), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n16820) );
  OAI211_X1 U20035 ( .C1(n16933), .C2(n16822), .A(n16821), .B(n16820), .ZN(
        n16828) );
  AOI22_X1 U20036 ( .A1(n17089), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17093), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n16826) );
  AOI22_X1 U20037 ( .A1(n17101), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17049), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n16825) );
  AOI22_X1 U20038 ( .A1(n17070), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17074), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n16824) );
  NAND2_X1 U20039 ( .A1(n17110), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n16823) );
  NAND4_X1 U20040 ( .A1(n16826), .A2(n16825), .A3(n16824), .A4(n16823), .ZN(
        n16827) );
  AOI211_X1 U20041 ( .C1(n16967), .C2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A(
        n16828), .B(n16827), .ZN(n16829) );
  OAI211_X1 U20042 ( .C1(n17027), .C2(n17013), .A(n16830), .B(n16829), .ZN(
        n16845) );
  NAND2_X1 U20043 ( .A1(n16846), .A2(n16845), .ZN(n16844) );
  AOI22_X1 U20044 ( .A1(n17092), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17049), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n16840) );
  AOI22_X1 U20045 ( .A1(n17002), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17095), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n16832) );
  AOI22_X1 U20046 ( .A1(n17089), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17101), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n16831) );
  OAI211_X1 U20047 ( .C1(n16933), .C2(n21058), .A(n16832), .B(n16831), .ZN(
        n16838) );
  AOI22_X1 U20048 ( .A1(n17070), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n16836) );
  AOI22_X1 U20049 ( .A1(n17103), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17093), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n16835) );
  AOI22_X1 U20050 ( .A1(n17074), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17100), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n16834) );
  NAND2_X1 U20051 ( .A1(n17110), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n16833) );
  NAND4_X1 U20052 ( .A1(n16836), .A2(n16835), .A3(n16834), .A4(n16833), .ZN(
        n16837) );
  AOI211_X1 U20053 ( .C1(n16967), .C2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A(
        n16838), .B(n16837), .ZN(n16839) );
  OAI211_X1 U20054 ( .C1(n9847), .C2(n20943), .A(n16840), .B(n16839), .ZN(
        n16841) );
  XOR2_X1 U20055 ( .A(n16844), .B(n16841), .Z(n17163) );
  OAI22_X1 U20056 ( .A1(n16843), .A2(n16842), .B1(n17163), .B2(n17141), .ZN(
        P3_U2673) );
  OAI21_X1 U20057 ( .B1(n16846), .B2(n16845), .A(n16844), .ZN(n17167) );
  AOI22_X1 U20058 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n16849), .B1(n16848), 
        .B2(n16847), .ZN(n16850) );
  OAI21_X1 U20059 ( .B1(n17167), .B2(n17141), .A(n16850), .ZN(P3_U2674) );
  OAI21_X1 U20060 ( .B1(n16855), .B2(n16852), .A(n16851), .ZN(n17176) );
  NAND3_X1 U20061 ( .A1(n16854), .A2(P3_EBX_REG_27__SCAN_IN), .A3(n16963), 
        .ZN(n16853) );
  OAI221_X1 U20062 ( .B1(n16854), .B2(P3_EBX_REG_27__SCAN_IN), .C1(n16963), 
        .C2(n17176), .A(n16853), .ZN(P3_U2676) );
  AOI21_X1 U20063 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n16963), .A(n16863), .ZN(
        n16858) );
  AOI21_X1 U20064 ( .B1(n16856), .B2(n16860), .A(n16855), .ZN(n17177) );
  INV_X1 U20065 ( .A(n17177), .ZN(n16857) );
  OAI22_X1 U20066 ( .A1(n16859), .A2(n16858), .B1(n16963), .B2(n16857), .ZN(
        P3_U2677) );
  AOI21_X1 U20067 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n16963), .A(n16868), .ZN(
        n16862) );
  OAI21_X1 U20068 ( .B1(n16864), .B2(n16861), .A(n16860), .ZN(n17186) );
  OAI22_X1 U20069 ( .A1(n16863), .A2(n16862), .B1(n16963), .B2(n17186), .ZN(
        P3_U2678) );
  AOI21_X1 U20070 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17141), .A(n16874), .ZN(
        n16867) );
  AOI21_X1 U20071 ( .B1(n16865), .B2(n16870), .A(n16864), .ZN(n17187) );
  INV_X1 U20072 ( .A(n17187), .ZN(n16866) );
  OAI22_X1 U20073 ( .A1(n16868), .A2(n16867), .B1(n16963), .B2(n16866), .ZN(
        P3_U2679) );
  AOI22_X1 U20074 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(n17141), .B1(
        P3_EBX_REG_22__SCAN_IN), .B2(n16869), .ZN(n16873) );
  OAI21_X1 U20075 ( .B1(n16872), .B2(n16871), .A(n16870), .ZN(n17197) );
  OAI22_X1 U20076 ( .A1(n16874), .A2(n16873), .B1(n16963), .B2(n17197), .ZN(
        P3_U2680) );
  AOI22_X1 U20077 ( .A1(n17095), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17049), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n16884) );
  AOI22_X1 U20078 ( .A1(n17101), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17100), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n16883) );
  AOI22_X1 U20079 ( .A1(n17077), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17110), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n16882) );
  OAI22_X1 U20080 ( .A1(n17027), .A2(n17126), .B1(n11811), .B2(n17013), .ZN(
        n16880) );
  AOI22_X1 U20081 ( .A1(n17089), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17083), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n16878) );
  AOI22_X1 U20082 ( .A1(n17070), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17103), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n16877) );
  AOI22_X1 U20083 ( .A1(n17002), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n16876) );
  NAND2_X1 U20084 ( .A1(n17074), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n16875) );
  NAND4_X1 U20085 ( .A1(n16878), .A2(n16877), .A3(n16876), .A4(n16875), .ZN(
        n16879) );
  AOI211_X1 U20086 ( .C1(n17076), .C2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A(
        n16880), .B(n16879), .ZN(n16881) );
  NAND4_X1 U20087 ( .A1(n16884), .A2(n16883), .A3(n16882), .A4(n16881), .ZN(
        n17198) );
  INV_X1 U20088 ( .A(n17198), .ZN(n16886) );
  NAND3_X1 U20089 ( .A1(n16887), .A2(P3_EBX_REG_22__SCAN_IN), .A3(n16963), 
        .ZN(n16885) );
  OAI221_X1 U20090 ( .B1(n16887), .B2(P3_EBX_REG_22__SCAN_IN), .C1(n16963), 
        .C2(n16886), .A(n16885), .ZN(P3_U2681) );
  NOR2_X1 U20091 ( .A1(n17150), .A2(n16888), .ZN(n16914) );
  AOI22_X1 U20092 ( .A1(n17094), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17093), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n16889) );
  OAI21_X1 U20093 ( .B1(n11820), .B2(n21003), .A(n16889), .ZN(n16900) );
  AOI22_X1 U20094 ( .A1(n17095), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17049), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n16898) );
  INV_X1 U20095 ( .A(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n16891) );
  AOI22_X1 U20096 ( .A1(n17101), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17074), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n16890) );
  OAI21_X1 U20097 ( .B1(n16933), .B2(n16891), .A(n16890), .ZN(n16896) );
  AOI22_X1 U20098 ( .A1(n17103), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n15497), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n16893) );
  AOI22_X1 U20099 ( .A1(n17089), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n16892) );
  OAI211_X1 U20100 ( .C1(n16987), .C2(n16894), .A(n16893), .B(n16892), .ZN(
        n16895) );
  AOI211_X1 U20101 ( .C1(n16967), .C2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A(
        n16896), .B(n16895), .ZN(n16897) );
  OAI211_X1 U20102 ( .C1(n17027), .C2(n17128), .A(n16898), .B(n16897), .ZN(
        n16899) );
  AOI211_X1 U20103 ( .C1(n17065), .C2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A(
        n16900), .B(n16899), .ZN(n17206) );
  INV_X1 U20104 ( .A(n17206), .ZN(n16901) );
  AOI22_X1 U20105 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n16914), .B1(n17150), 
        .B2(n16901), .ZN(n16902) );
  OAI21_X1 U20106 ( .B1(P3_EBX_REG_21__SCAN_IN), .B2(n16903), .A(n16902), .ZN(
        P3_U2682) );
  AOI22_X1 U20107 ( .A1(n17103), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17110), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n16913) );
  AOI22_X1 U20108 ( .A1(n17095), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17083), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n16905) );
  AOI22_X1 U20109 ( .A1(n17089), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n16904) );
  OAI211_X1 U20110 ( .C1(n11811), .C2(n17018), .A(n16905), .B(n16904), .ZN(
        n16911) );
  AOI22_X1 U20111 ( .A1(n17101), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17093), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n16909) );
  AOI22_X1 U20112 ( .A1(n17002), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17049), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n16908) );
  AOI22_X1 U20113 ( .A1(n17070), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n15497), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n16907) );
  NAND2_X1 U20114 ( .A1(n17074), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n16906) );
  NAND4_X1 U20115 ( .A1(n16909), .A2(n16908), .A3(n16907), .A4(n16906), .ZN(
        n16910) );
  AOI211_X1 U20116 ( .C1(n17077), .C2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A(
        n16911), .B(n16910), .ZN(n16912) );
  OAI211_X1 U20117 ( .C1(n17027), .C2(n17133), .A(n16913), .B(n16912), .ZN(
        n17210) );
  INV_X1 U20118 ( .A(n17210), .ZN(n16917) );
  OAI21_X1 U20119 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n16915), .A(n16914), .ZN(
        n16916) );
  OAI21_X1 U20120 ( .B1(n16917), .B2(n17141), .A(n16916), .ZN(P3_U2683) );
  AOI22_X1 U20121 ( .A1(n17076), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n15497), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n16918) );
  OAI21_X1 U20122 ( .B1(n17114), .B2(n18443), .A(n16918), .ZN(n16928) );
  AOI22_X1 U20123 ( .A1(n17092), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11832), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n16926) );
  AOI22_X1 U20124 ( .A1(n17110), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17049), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n16919) );
  OAI21_X1 U20125 ( .B1(n11799), .B2(n17034), .A(n16919), .ZN(n16924) );
  AOI22_X1 U20126 ( .A1(n17101), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17103), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n16921) );
  AOI22_X1 U20127 ( .A1(n17095), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17083), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n16920) );
  OAI211_X1 U20128 ( .C1(n16933), .C2(n16922), .A(n16921), .B(n16920), .ZN(
        n16923) );
  AOI211_X1 U20129 ( .C1(n16967), .C2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A(
        n16924), .B(n16923), .ZN(n16925) );
  OAI211_X1 U20130 ( .C1(n16970), .C2(n17033), .A(n16926), .B(n16925), .ZN(
        n16927) );
  AOI211_X1 U20131 ( .C1(n17036), .C2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A(
        n16928), .B(n16927), .ZN(n17219) );
  OAI21_X1 U20132 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n16930), .A(n16929), .ZN(
        n16931) );
  AOI22_X1 U20133 ( .A1(n17150), .A2(n17219), .B1(n16931), .B2(n16963), .ZN(
        P3_U2684) );
  NAND2_X1 U20134 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n16932), .ZN(n16948) );
  INV_X1 U20135 ( .A(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n21100) );
  OAI22_X1 U20136 ( .A1(n11799), .A2(n16934), .B1(n16933), .B2(n21100), .ZN(
        n16944) );
  AOI22_X1 U20137 ( .A1(n17049), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n15497), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n16942) );
  AOI22_X1 U20138 ( .A1(n17094), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n16941) );
  AOI22_X1 U20139 ( .A1(n17092), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17103), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n16935) );
  OAI21_X1 U20140 ( .B1(n16970), .B2(n17052), .A(n16935), .ZN(n16939) );
  AOI22_X1 U20141 ( .A1(n17070), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17054), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n16937) );
  AOI22_X1 U20142 ( .A1(n17095), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17076), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n16936) );
  OAI211_X1 U20143 ( .C1(n11811), .C2(n17062), .A(n16937), .B(n16936), .ZN(
        n16938) );
  AOI211_X1 U20144 ( .C1(n17110), .C2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A(
        n16939), .B(n16938), .ZN(n16940) );
  NAND3_X1 U20145 ( .A1(n16942), .A2(n16941), .A3(n16940), .ZN(n16943) );
  AOI211_X1 U20146 ( .C1(n17065), .C2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A(
        n16944), .B(n16943), .ZN(n17223) );
  INV_X1 U20147 ( .A(n17115), .ZN(n17069) );
  NAND2_X1 U20148 ( .A1(P3_EBX_REG_11__SCAN_IN), .A2(n17068), .ZN(n17046) );
  NOR2_X1 U20149 ( .A1(n17291), .A2(n17046), .ZN(n17031) );
  NAND2_X1 U20150 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17031), .ZN(n16949) );
  INV_X1 U20151 ( .A(n16949), .ZN(n17000) );
  NAND3_X1 U20152 ( .A1(n16946), .A2(n17000), .A3(n16945), .ZN(n16947) );
  OAI221_X1 U20153 ( .B1(n17150), .B2(n16948), .C1(n17141), .C2(n17223), .A(
        n16947), .ZN(P3_U2685) );
  INV_X1 U20154 ( .A(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n20927) );
  AOI22_X1 U20155 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n17054), .B1(
        P3_INSTQUEUE_REG_14__1__SCAN_IN), .B2(n15497), .ZN(n16951) );
  OAI21_X1 U20156 ( .B1(n17114), .B2(n20927), .A(n16951), .ZN(n16961) );
  AOI22_X1 U20157 ( .A1(n17089), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n17103), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n16959) );
  AOI22_X1 U20158 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n17110), .B1(
        n17074), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n16952) );
  OAI21_X1 U20159 ( .B1(n11820), .B2(n17075), .A(n16952), .ZN(n16957) );
  AOI22_X1 U20160 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n17049), .B1(
        P3_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n17102), .ZN(n16954) );
  AOI22_X1 U20161 ( .A1(n17094), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n17076), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n16953) );
  OAI211_X1 U20162 ( .C1(n11811), .C2(n16955), .A(n16954), .B(n16953), .ZN(
        n16956) );
  AOI211_X1 U20163 ( .C1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .C2(n17077), .A(
        n16957), .B(n16956), .ZN(n16958) );
  OAI211_X1 U20164 ( .C1(n17027), .C2(n17145), .A(n16959), .B(n16958), .ZN(
        n16960) );
  AOI211_X1 U20165 ( .C1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .C2(n17095), .A(
        n16961), .B(n16960), .ZN(n17229) );
  NAND3_X1 U20166 ( .A1(n16980), .A2(P3_EBX_REG_17__SCAN_IN), .A3(n16963), 
        .ZN(n16962) );
  OAI221_X1 U20167 ( .B1(n16980), .B2(P3_EBX_REG_17__SCAN_IN), .C1(n16963), 
        .C2(n17229), .A(n16962), .ZN(P3_U2686) );
  AOI22_X1 U20168 ( .A1(n17076), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n15497), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n16964) );
  OAI21_X1 U20169 ( .B1(n16966), .B2(n16965), .A(n16964), .ZN(n16979) );
  AOI22_X1 U20170 ( .A1(n17092), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n16967), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n16977) );
  OAI22_X1 U20171 ( .A1(n16970), .A2(n16969), .B1(n16983), .B2(n16968), .ZN(
        n16975) );
  AOI22_X1 U20172 ( .A1(n17095), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17049), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n16973) );
  AOI22_X1 U20173 ( .A1(n17094), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n15498), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n16972) );
  AOI22_X1 U20174 ( .A1(n17077), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17110), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n16971) );
  NAND3_X1 U20175 ( .A1(n16973), .A2(n16972), .A3(n16971), .ZN(n16974) );
  AOI211_X1 U20176 ( .C1(n17074), .C2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A(
        n16975), .B(n16974), .ZN(n16976) );
  OAI211_X1 U20177 ( .C1(n17114), .C2(n21054), .A(n16977), .B(n16976), .ZN(
        n16978) );
  AOI211_X1 U20178 ( .C1(n17103), .C2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A(
        n16979), .B(n16978), .ZN(n17236) );
  NAND3_X1 U20179 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(P3_EBX_REG_13__SCAN_IN), 
        .A3(n17001), .ZN(n16997) );
  NOR2_X1 U20180 ( .A1(n16998), .A2(n16997), .ZN(n16996) );
  OAI211_X1 U20181 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n16996), .A(n16980), .B(
        n16963), .ZN(n16981) );
  OAI21_X1 U20182 ( .B1(n17236), .B2(n17141), .A(n16981), .ZN(P3_U2687) );
  AOI22_X1 U20183 ( .A1(n17095), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17074), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n16995) );
  AOI22_X1 U20184 ( .A1(n17070), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n15497), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n16982) );
  OAI21_X1 U20185 ( .B1(n16983), .B2(n21058), .A(n16982), .ZN(n16993) );
  AOI22_X1 U20186 ( .A1(n17094), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17092), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n16990) );
  AOI22_X1 U20187 ( .A1(n17036), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17049), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n16985) );
  AOI22_X1 U20188 ( .A1(n17089), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17103), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n16984) );
  OAI211_X1 U20189 ( .C1(n16987), .C2(n16986), .A(n16985), .B(n16984), .ZN(
        n16988) );
  AOI21_X1 U20190 ( .B1(n17077), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A(
        n16988), .ZN(n16989) );
  OAI211_X1 U20191 ( .C1(n11811), .C2(n16991), .A(n16990), .B(n16989), .ZN(
        n16992) );
  AOI211_X1 U20192 ( .C1(n17065), .C2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A(
        n16993), .B(n16992), .ZN(n16994) );
  OAI211_X1 U20193 ( .C1(n9848), .C2(n20943), .A(n16995), .B(n16994), .ZN(
        n17240) );
  AOI21_X1 U20194 ( .B1(n16998), .B2(n16997), .A(n16996), .ZN(n16999) );
  MUX2_X1 U20195 ( .A(n17240), .B(n16999), .S(n17141), .Z(P3_U2688) );
  NAND2_X1 U20196 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n17000), .ZN(n17016) );
  NAND2_X1 U20197 ( .A1(n18145), .A2(n17146), .ZN(n17152) );
  OAI22_X1 U20198 ( .A1(n17150), .A2(n17001), .B1(P3_EBX_REG_13__SCAN_IN), 
        .B2(n17152), .ZN(n17014) );
  AOI22_X1 U20199 ( .A1(n17074), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17077), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17012) );
  AOI22_X1 U20200 ( .A1(n17070), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17054), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n17004) );
  AOI22_X1 U20201 ( .A1(n17002), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17076), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17003) );
  OAI211_X1 U20202 ( .C1(n11811), .C2(n17126), .A(n17004), .B(n17003), .ZN(
        n17010) );
  AOI22_X1 U20203 ( .A1(n17095), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n15497), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17008) );
  AOI22_X1 U20204 ( .A1(n17094), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17007) );
  AOI22_X1 U20205 ( .A1(n17089), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17049), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17006) );
  NAND2_X1 U20206 ( .A1(n17092), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n17005) );
  NAND4_X1 U20207 ( .A1(n17008), .A2(n17007), .A3(n17006), .A4(n17005), .ZN(
        n17009) );
  AOI211_X1 U20208 ( .C1(n17110), .C2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A(
        n17010), .B(n17009), .ZN(n17011) );
  OAI211_X1 U20209 ( .C1(n10222), .C2(n17013), .A(n17012), .B(n17011), .ZN(
        n17245) );
  AOI22_X1 U20210 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n17014), .B1(n17150), 
        .B2(n17245), .ZN(n17015) );
  OAI21_X1 U20211 ( .B1(P3_EBX_REG_14__SCAN_IN), .B2(n17016), .A(n17015), .ZN(
        P3_U2689) );
  AOI22_X1 U20212 ( .A1(n17002), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17095), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n17017) );
  OAI21_X1 U20213 ( .B1(n10222), .B2(n17018), .A(n17017), .ZN(n17029) );
  INV_X1 U20214 ( .A(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17026) );
  AOI22_X1 U20215 ( .A1(n17036), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17049), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17025) );
  AOI22_X1 U20216 ( .A1(n17074), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17110), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17019) );
  OAI21_X1 U20217 ( .B1(n17051), .B2(n20935), .A(n17019), .ZN(n17023) );
  AOI22_X1 U20218 ( .A1(n17101), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17076), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17021) );
  AOI22_X1 U20219 ( .A1(n17094), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17070), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n17020) );
  OAI211_X1 U20220 ( .C1(n11811), .C2(n17133), .A(n17021), .B(n17020), .ZN(
        n17022) );
  AOI211_X1 U20221 ( .C1(n17077), .C2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A(
        n17023), .B(n17022), .ZN(n17024) );
  OAI211_X1 U20222 ( .C1(n17027), .C2(n17026), .A(n17025), .B(n17024), .ZN(
        n17028) );
  AOI211_X1 U20223 ( .C1(n17089), .C2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A(
        n17029), .B(n17028), .ZN(n17254) );
  OAI21_X1 U20224 ( .B1(P3_EBX_REG_12__SCAN_IN), .B2(n17031), .A(n17030), .ZN(
        n17032) );
  OAI21_X1 U20225 ( .B1(n17254), .B2(n17141), .A(n17032), .ZN(P3_U2691) );
  AOI22_X1 U20226 ( .A1(n17089), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17095), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17045) );
  AOI22_X1 U20227 ( .A1(n17101), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17049), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17044) );
  OAI22_X1 U20228 ( .A1(n9847), .A2(n17034), .B1(n9848), .B2(n17033), .ZN(
        n17042) );
  OAI22_X1 U20229 ( .A1(n11811), .A2(n17137), .B1(n17051), .B2(n18443), .ZN(
        n17035) );
  AOI21_X1 U20230 ( .B1(n17092), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A(
        n17035), .ZN(n17040) );
  AOI22_X1 U20231 ( .A1(n17070), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n17039) );
  AOI22_X1 U20232 ( .A1(n17002), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17103), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17038) );
  AOI22_X1 U20233 ( .A1(n17077), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17110), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17037) );
  NAND4_X1 U20234 ( .A1(n17040), .A2(n17039), .A3(n17038), .A4(n17037), .ZN(
        n17041) );
  AOI211_X1 U20235 ( .C1(n17074), .C2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A(
        n17042), .B(n17041), .ZN(n17043) );
  NAND3_X1 U20236 ( .A1(n17045), .A2(n17044), .A3(n17043), .ZN(n17258) );
  INV_X1 U20237 ( .A(n17258), .ZN(n17048) );
  OAI21_X1 U20238 ( .B1(P3_EBX_REG_11__SCAN_IN), .B2(n17068), .A(n17046), .ZN(
        n17047) );
  AOI22_X1 U20239 ( .A1(n17150), .A2(n17048), .B1(n17047), .B2(n16963), .ZN(
        P3_U2692) );
  AOI22_X1 U20240 ( .A1(n17102), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17049), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17050) );
  OAI21_X1 U20241 ( .B1(n17051), .B2(n18439), .A(n17050), .ZN(n17064) );
  AOI22_X1 U20242 ( .A1(n17092), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17110), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n17061) );
  OAI22_X1 U20243 ( .A1(n11799), .A2(n21070), .B1(n9848), .B2(n17052), .ZN(
        n17059) );
  AOI22_X1 U20244 ( .A1(n17089), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17095), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17057) );
  AOI22_X1 U20245 ( .A1(n17070), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17054), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17056) );
  AOI22_X1 U20246 ( .A1(n16967), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17077), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17055) );
  NAND3_X1 U20247 ( .A1(n17057), .A2(n17056), .A3(n17055), .ZN(n17058) );
  AOI211_X1 U20248 ( .C1(n17083), .C2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A(
        n17059), .B(n17058), .ZN(n17060) );
  OAI211_X1 U20249 ( .C1(n10222), .C2(n17062), .A(n17061), .B(n17060), .ZN(
        n17063) );
  AOI211_X1 U20250 ( .C1(n17065), .C2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A(
        n17064), .B(n17063), .ZN(n17261) );
  NOR2_X1 U20251 ( .A1(n17066), .A2(n17115), .ZN(n17091) );
  OAI21_X1 U20252 ( .B1(P3_EBX_REG_10__SCAN_IN), .B2(n17091), .A(n17141), .ZN(
        n17067) );
  OAI22_X1 U20253 ( .A1(n17261), .A2(n17141), .B1(n17068), .B2(n17067), .ZN(
        P3_U2693) );
  OAI21_X1 U20254 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n17069), .A(n17141), .ZN(
        n17090) );
  AOI22_X1 U20255 ( .A1(n17070), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n17103), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n17071) );
  OAI21_X1 U20256 ( .B1(n17073), .B2(n17072), .A(n17071), .ZN(n17088) );
  AOI22_X1 U20257 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n17074), .B1(
        P3_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n17102), .ZN(n17085) );
  OAI22_X1 U20258 ( .A1(n17027), .A2(n17075), .B1(n11811), .B2(n17145), .ZN(
        n17082) );
  AOI22_X1 U20259 ( .A1(n17002), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_13__1__SCAN_IN), .B2(n15497), .ZN(n17080) );
  AOI22_X1 U20260 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n17076), .B1(
        n17095), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n17079) );
  AOI22_X1 U20261 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n17077), .B1(
        n17110), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n17078) );
  NAND3_X1 U20262 ( .A1(n17080), .A2(n17079), .A3(n17078), .ZN(n17081) );
  AOI211_X1 U20263 ( .C1(n17083), .C2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A(
        n17082), .B(n17081), .ZN(n17084) );
  OAI211_X1 U20264 ( .C1(n16983), .C2(n17086), .A(n17085), .B(n17084), .ZN(
        n17087) );
  AOI211_X1 U20265 ( .C1(n17089), .C2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A(
        n17088), .B(n17087), .ZN(n17264) );
  OAI22_X1 U20266 ( .A1(n17091), .A2(n17090), .B1(n17264), .B2(n17141), .ZN(
        P3_U2694) );
  INV_X1 U20267 ( .A(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17113) );
  AOI22_X1 U20268 ( .A1(n17092), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11832), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n17112) );
  INV_X1 U20269 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17099) );
  AOI22_X1 U20270 ( .A1(n17094), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17093), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17098) );
  AOI22_X1 U20271 ( .A1(n17089), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17095), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17097) );
  OAI211_X1 U20272 ( .C1(n11811), .C2(n17099), .A(n17098), .B(n17097), .ZN(
        n17109) );
  AOI22_X1 U20273 ( .A1(n17101), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17100), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n17107) );
  AOI22_X1 U20274 ( .A1(n17103), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17102), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17106) );
  AOI22_X1 U20275 ( .A1(n17074), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17049), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17105) );
  NAND2_X1 U20276 ( .A1(n17077), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n17104) );
  NAND4_X1 U20277 ( .A1(n17107), .A2(n17106), .A3(n17105), .A4(n17104), .ZN(
        n17108) );
  AOI211_X1 U20278 ( .C1(n17110), .C2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A(
        n17109), .B(n17108), .ZN(n17111) );
  OAI211_X1 U20279 ( .C1(n17114), .C2(n17113), .A(n17112), .B(n17111), .ZN(
        n17268) );
  INV_X1 U20280 ( .A(n17268), .ZN(n17117) );
  OAI21_X1 U20281 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(n17118), .A(n17115), .ZN(
        n17116) );
  AOI22_X1 U20282 ( .A1(n17150), .A2(n17117), .B1(n17116), .B2(n16963), .ZN(
        P3_U2695) );
  NOR2_X1 U20283 ( .A1(n17291), .A2(n17122), .ZN(n17134) );
  NAND3_X1 U20284 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(P3_EBX_REG_5__SCAN_IN), 
        .A3(n17134), .ZN(n17124) );
  OAI21_X1 U20285 ( .B1(n17119), .B2(n17118), .A(n17141), .ZN(n17120) );
  OAI21_X1 U20286 ( .B1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B2(n17141), .A(
        n17120), .ZN(n17121) );
  OAI21_X1 U20287 ( .B1(P3_EBX_REG_7__SCAN_IN), .B2(n17124), .A(n17121), .ZN(
        P3_U2696) );
  NOR2_X1 U20288 ( .A1(n17123), .A2(n17122), .ZN(n17130) );
  OAI21_X1 U20289 ( .B1(P3_EBX_REG_6__SCAN_IN), .B2(n17130), .A(n17124), .ZN(
        n17125) );
  AOI22_X1 U20290 ( .A1(n17150), .A2(n17126), .B1(n17125), .B2(n17141), .ZN(
        P3_U2697) );
  OAI21_X1 U20291 ( .B1(P3_EBX_REG_5__SCAN_IN), .B2(n17127), .A(n17141), .ZN(
        n17129) );
  OAI22_X1 U20292 ( .A1(n17130), .A2(n17129), .B1(n17128), .B2(n17141), .ZN(
        P3_U2698) );
  NOR2_X1 U20293 ( .A1(n17131), .A2(n17152), .ZN(n17140) );
  NAND2_X1 U20294 ( .A1(P3_EBX_REG_2__SCAN_IN), .A2(n17140), .ZN(n17136) );
  NOR2_X1 U20295 ( .A1(n17132), .A2(n17136), .ZN(n17139) );
  AOI21_X1 U20296 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n16963), .A(n17139), .ZN(
        n17135) );
  OAI22_X1 U20297 ( .A1(n17135), .A2(n17134), .B1(n17133), .B2(n17141), .ZN(
        P3_U2699) );
  INV_X1 U20298 ( .A(n17136), .ZN(n17144) );
  AOI21_X1 U20299 ( .B1(P3_EBX_REG_3__SCAN_IN), .B2(n16963), .A(n17144), .ZN(
        n17138) );
  OAI22_X1 U20300 ( .A1(n17139), .A2(n17138), .B1(n17137), .B2(n17141), .ZN(
        P3_U2700) );
  AOI21_X1 U20301 ( .B1(P3_EBX_REG_2__SCAN_IN), .B2(n16963), .A(n17140), .ZN(
        n17143) );
  INV_X1 U20302 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17142) );
  OAI22_X1 U20303 ( .A1(n17144), .A2(n17143), .B1(n17142), .B2(n17141), .ZN(
        P3_U2701) );
  OAI222_X1 U20304 ( .A1(n17148), .A2(n17152), .B1(n17147), .B2(n17146), .C1(
        n17145), .C2(n16963), .ZN(P3_U2702) );
  AOI22_X1 U20305 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n17150), .B1(
        P3_EBX_REG_0__SCAN_IN), .B2(n17149), .ZN(n17151) );
  OAI21_X1 U20306 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(n17152), .A(n17151), .ZN(
        P3_U2703) );
  INV_X1 U20307 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n17373) );
  INV_X1 U20308 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n17369) );
  INV_X1 U20309 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n17361) );
  INV_X1 U20310 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n17351) );
  INV_X1 U20311 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n17413) );
  INV_X1 U20312 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n17393) );
  INV_X1 U20313 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n17391) );
  INV_X1 U20314 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n17389) );
  INV_X1 U20315 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n17387) );
  NOR4_X1 U20316 ( .A1(n17393), .A2(n17391), .A3(n17389), .A4(n17387), .ZN(
        n17153) );
  NAND3_X1 U20317 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(P3_EAX_REG_2__SCAN_IN), 
        .A3(n17153), .ZN(n17237) );
  NOR2_X2 U20318 ( .A1(n17302), .A2(n17237), .ZN(n17269) );
  INV_X1 U20319 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n17399) );
  NAND2_X1 U20320 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(P3_EAX_REG_8__SCAN_IN), 
        .ZN(n17243) );
  NAND4_X1 U20321 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(P3_EAX_REG_11__SCAN_IN), 
        .A3(P3_EAX_REG_14__SCAN_IN), .A4(P3_EAX_REG_13__SCAN_IN), .ZN(n17154)
         );
  NOR3_X1 U20322 ( .A1(n17399), .A2(n17243), .A3(n17154), .ZN(n17238) );
  NAND2_X1 U20323 ( .A1(n17269), .A2(n17238), .ZN(n17239) );
  NAND4_X1 U20324 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(P3_EAX_REG_21__SCAN_IN), 
        .A3(P3_EAX_REG_20__SCAN_IN), .A4(P3_EAX_REG_18__SCAN_IN), .ZN(n17204)
         );
  NAND2_X1 U20325 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n17194), .ZN(n17193) );
  NAND2_X1 U20326 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n17188), .ZN(n17189) );
  NAND2_X1 U20327 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n17169), .ZN(n17164) );
  NAND2_X1 U20328 ( .A1(n17160), .A2(P3_EAX_REG_30__SCAN_IN), .ZN(n17159) );
  NAND2_X1 U20329 ( .A1(n17156), .A2(n17270), .ZN(n17205) );
  OAI22_X1 U20330 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(n17199), .B1(n17270), 
        .B2(n17160), .ZN(n17157) );
  AOI22_X1 U20331 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n17230), .B1(
        P3_EAX_REG_31__SCAN_IN), .B2(n17157), .ZN(n17158) );
  OAI21_X1 U20332 ( .B1(P3_EAX_REG_31__SCAN_IN), .B2(n17159), .A(n17158), .ZN(
        P3_U2704) );
  NAND2_X1 U20333 ( .A1(n18135), .A2(n17270), .ZN(n17214) );
  AOI22_X1 U20334 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17231), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n17230), .ZN(n17162) );
  OAI211_X1 U20335 ( .C1(n17160), .C2(P3_EAX_REG_30__SCAN_IN), .A(n17303), .B(
        n17159), .ZN(n17161) );
  OAI211_X1 U20336 ( .C1(n17163), .C2(n17295), .A(n17162), .B(n17161), .ZN(
        P3_U2705) );
  AOI22_X1 U20337 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17231), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n17230), .ZN(n17166) );
  OAI211_X1 U20338 ( .C1(n17169), .C2(P3_EAX_REG_29__SCAN_IN), .A(n17303), .B(
        n17164), .ZN(n17165) );
  OAI211_X1 U20339 ( .C1(n17167), .C2(n17295), .A(n17166), .B(n17165), .ZN(
        P3_U2706) );
  AOI22_X1 U20340 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17231), .B1(n17300), .B2(
        n17168), .ZN(n17172) );
  AOI211_X1 U20341 ( .C1(n17373), .C2(n17173), .A(n17169), .B(n17270), .ZN(
        n17170) );
  INV_X1 U20342 ( .A(n17170), .ZN(n17171) );
  OAI211_X1 U20343 ( .C1(n17205), .C2(n18128), .A(n17172), .B(n17171), .ZN(
        P3_U2707) );
  AOI22_X1 U20344 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17231), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n17230), .ZN(n17175) );
  OAI211_X1 U20345 ( .C1(n17178), .C2(P3_EAX_REG_27__SCAN_IN), .A(n17303), .B(
        n17173), .ZN(n17174) );
  OAI211_X1 U20346 ( .C1(n17176), .C2(n17295), .A(n17175), .B(n17174), .ZN(
        P3_U2708) );
  INV_X1 U20347 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n20866) );
  AOI22_X1 U20348 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n17230), .B1(n17300), .B2(
        n17177), .ZN(n17181) );
  AOI211_X1 U20349 ( .C1(n17369), .C2(n17182), .A(n17178), .B(n17270), .ZN(
        n17179) );
  INV_X1 U20350 ( .A(n17179), .ZN(n17180) );
  OAI211_X1 U20351 ( .C1(n17214), .C2(n20866), .A(n17181), .B(n17180), .ZN(
        P3_U2709) );
  AOI22_X1 U20352 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17231), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n17230), .ZN(n17185) );
  OAI211_X1 U20353 ( .C1(n17183), .C2(P3_EAX_REG_25__SCAN_IN), .A(n17303), .B(
        n17182), .ZN(n17184) );
  OAI211_X1 U20354 ( .C1(n17186), .C2(n17295), .A(n17185), .B(n17184), .ZN(
        P3_U2710) );
  INV_X1 U20355 ( .A(BUF2_REG_24__SCAN_IN), .ZN(n17192) );
  AOI22_X1 U20356 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17231), .B1(n17300), .B2(
        n17187), .ZN(n17191) );
  OAI211_X1 U20357 ( .C1(n17188), .C2(P3_EAX_REG_24__SCAN_IN), .A(n17303), .B(
        n17189), .ZN(n17190) );
  OAI211_X1 U20358 ( .C1(n17205), .C2(n17192), .A(n17191), .B(n17190), .ZN(
        P3_U2711) );
  AOI22_X1 U20359 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17231), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n17230), .ZN(n17196) );
  OAI211_X1 U20360 ( .C1(P3_EAX_REG_23__SCAN_IN), .C2(n17194), .A(n17303), .B(
        n17193), .ZN(n17195) );
  OAI211_X1 U20361 ( .C1(n17197), .C2(n17295), .A(n17196), .B(n17195), .ZN(
        P3_U2712) );
  NAND2_X1 U20362 ( .A1(n17224), .A2(n17361), .ZN(n17203) );
  AOI22_X1 U20363 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n17230), .B1(n17300), .B2(
        n17198), .ZN(n17202) );
  INV_X1 U20364 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n17355) );
  NAND2_X1 U20365 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17224), .ZN(n17220) );
  NAND2_X1 U20366 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17215), .ZN(n17211) );
  NAND2_X1 U20367 ( .A1(n17303), .A2(n17211), .ZN(n17209) );
  OAI21_X1 U20368 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17199), .A(n17209), .ZN(
        n17200) );
  AOI22_X1 U20369 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17231), .B1(
        P3_EAX_REG_22__SCAN_IN), .B2(n17200), .ZN(n17201) );
  OAI211_X1 U20370 ( .C1(n17204), .C2(n17203), .A(n17202), .B(n17201), .ZN(
        P3_U2713) );
  INV_X1 U20371 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n17359) );
  INV_X1 U20372 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n18133) );
  OAI22_X1 U20373 ( .A1(n17206), .A2(n17295), .B1(n18133), .B2(n17205), .ZN(
        n17207) );
  AOI21_X1 U20374 ( .B1(BUF2_REG_5__SCAN_IN), .B2(n17231), .A(n17207), .ZN(
        n17208) );
  OAI221_X1 U20375 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17211), .C1(n17359), 
        .C2(n17209), .A(n17208), .ZN(P3_U2714) );
  AOI22_X1 U20376 ( .A1(BUF2_REG_20__SCAN_IN), .A2(n17230), .B1(n17300), .B2(
        n17210), .ZN(n17213) );
  OAI211_X1 U20377 ( .C1(n17215), .C2(P3_EAX_REG_20__SCAN_IN), .A(n17303), .B(
        n17211), .ZN(n17212) );
  OAI211_X1 U20378 ( .C1(n17214), .C2(n18129), .A(n17213), .B(n17212), .ZN(
        P3_U2715) );
  AOI22_X1 U20379 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17231), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n17230), .ZN(n17218) );
  AOI211_X1 U20380 ( .C1(n17355), .C2(n17220), .A(n17215), .B(n17270), .ZN(
        n17216) );
  INV_X1 U20381 ( .A(n17216), .ZN(n17217) );
  OAI211_X1 U20382 ( .C1(n17219), .C2(n17295), .A(n17218), .B(n17217), .ZN(
        P3_U2716) );
  AOI22_X1 U20383 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17231), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n17230), .ZN(n17222) );
  OAI211_X1 U20384 ( .C1(n17224), .C2(P3_EAX_REG_18__SCAN_IN), .A(n17303), .B(
        n17220), .ZN(n17221) );
  OAI211_X1 U20385 ( .C1(n17223), .C2(n17295), .A(n17222), .B(n17221), .ZN(
        P3_U2717) );
  AOI22_X1 U20386 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17231), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n17230), .ZN(n17228) );
  INV_X1 U20387 ( .A(n17232), .ZN(n17226) );
  INV_X1 U20388 ( .A(n17224), .ZN(n17225) );
  OAI211_X1 U20389 ( .C1(n17226), .C2(P3_EAX_REG_17__SCAN_IN), .A(n17303), .B(
        n17225), .ZN(n17227) );
  OAI211_X1 U20390 ( .C1(n17229), .C2(n17295), .A(n17228), .B(n17227), .ZN(
        P3_U2718) );
  AOI22_X1 U20391 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17231), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n17230), .ZN(n17235) );
  OAI211_X1 U20392 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n17233), .A(n17232), .B(
        n17303), .ZN(n17234) );
  OAI211_X1 U20393 ( .C1(n17236), .C2(n17295), .A(n17235), .B(n17234), .ZN(
        P3_U2719) );
  NAND2_X1 U20394 ( .A1(n17238), .A2(n17276), .ZN(n17242) );
  NAND2_X1 U20395 ( .A1(n17303), .A2(n17239), .ZN(n17247) );
  AOI22_X1 U20396 ( .A1(n17300), .A2(n17240), .B1(BUF2_REG_15__SCAN_IN), .B2(
        n17301), .ZN(n17241) );
  OAI221_X1 U20397 ( .B1(P3_EAX_REG_15__SCAN_IN), .B2(n17242), .C1(n17413), 
        .C2(n17247), .A(n17241), .ZN(P3_U2720) );
  NAND2_X1 U20398 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(P3_EAX_REG_11__SCAN_IN), 
        .ZN(n17244) );
  INV_X1 U20399 ( .A(n17276), .ZN(n17273) );
  NAND2_X1 U20400 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17266), .ZN(n17260) );
  NOR2_X1 U20401 ( .A1(n17244), .A2(n17260), .ZN(n17256) );
  NAND2_X1 U20402 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n17256), .ZN(n17248) );
  INV_X1 U20403 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n17408) );
  AOI22_X1 U20404 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17301), .B1(n17300), .B2(
        n17245), .ZN(n17246) );
  OAI221_X1 U20405 ( .B1(P3_EAX_REG_14__SCAN_IN), .B2(n17248), .C1(n17408), 
        .C2(n17247), .A(n17246), .ZN(P3_U2721) );
  INV_X1 U20406 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n17252) );
  INV_X1 U20407 ( .A(n17248), .ZN(n17251) );
  AOI21_X1 U20408 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(n17303), .A(n17256), .ZN(
        n17250) );
  OAI222_X1 U20409 ( .A1(n17298), .A2(n17252), .B1(n17251), .B2(n17250), .C1(
        n17295), .C2(n17249), .ZN(P3_U2722) );
  INV_X1 U20410 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n17257) );
  INV_X1 U20411 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n17401) );
  INV_X1 U20412 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n17404) );
  OAI22_X1 U20413 ( .A1(n17260), .A2(n17401), .B1(n17404), .B2(n17270), .ZN(
        n17253) );
  INV_X1 U20414 ( .A(n17253), .ZN(n17255) );
  OAI222_X1 U20415 ( .A1(n17298), .A2(n17257), .B1(n17256), .B2(n17255), .C1(
        n17295), .C2(n17254), .ZN(P3_U2723) );
  NAND2_X1 U20416 ( .A1(n17303), .A2(n17260), .ZN(n17263) );
  AOI22_X1 U20417 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17301), .B1(n17300), .B2(
        n17258), .ZN(n17259) );
  OAI221_X1 U20418 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n17260), .C1(n17401), 
        .C2(n17263), .A(n17259), .ZN(P3_U2724) );
  NOR2_X1 U20419 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17266), .ZN(n17262) );
  OAI222_X1 U20420 ( .A1(n17298), .A2(n20866), .B1(n17263), .B2(n17262), .C1(
        n17295), .C2(n17261), .ZN(P3_U2725) );
  INV_X1 U20421 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n17267) );
  AOI22_X1 U20422 ( .A1(n17276), .A2(P3_EAX_REG_8__SCAN_IN), .B1(
        P3_EAX_REG_9__SCAN_IN), .B2(n17303), .ZN(n17265) );
  OAI222_X1 U20423 ( .A1(n17298), .A2(n17267), .B1(n17266), .B2(n17265), .C1(
        n17295), .C2(n17264), .ZN(P3_U2726) );
  AOI22_X1 U20424 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17301), .B1(n17300), .B2(
        n17268), .ZN(n17272) );
  INV_X1 U20425 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n17395) );
  OR3_X1 U20426 ( .A1(n17395), .A2(n17270), .A3(n17269), .ZN(n17271) );
  OAI211_X1 U20427 ( .C1(P3_EAX_REG_8__SCAN_IN), .C2(n17273), .A(n17272), .B(
        n17271), .ZN(P3_U2727) );
  INV_X1 U20428 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n21002) );
  INV_X1 U20429 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n17383) );
  NOR3_X1 U20430 ( .A1(n17291), .A2(n17302), .A3(n17383), .ZN(n17297) );
  NAND2_X1 U20431 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n17297), .ZN(n17284) );
  NOR2_X1 U20432 ( .A1(n17387), .A2(n17284), .ZN(n17287) );
  NAND2_X1 U20433 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n17287), .ZN(n17277) );
  NOR2_X1 U20434 ( .A1(n17391), .A2(n17277), .ZN(n17280) );
  AOI21_X1 U20435 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n17303), .A(n17280), .ZN(
        n17275) );
  OAI222_X1 U20436 ( .A1(n17298), .A2(n21002), .B1(n17276), .B2(n17275), .C1(
        n17295), .C2(n17274), .ZN(P3_U2728) );
  INV_X1 U20437 ( .A(n17277), .ZN(n17283) );
  AOI21_X1 U20438 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n17303), .A(n17283), .ZN(
        n17279) );
  OAI222_X1 U20439 ( .A1(n18139), .A2(n17298), .B1(n17280), .B2(n17279), .C1(
        n17295), .C2(n17278), .ZN(P3_U2729) );
  INV_X1 U20440 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n18134) );
  AOI21_X1 U20441 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n17303), .A(n17287), .ZN(
        n17282) );
  OAI222_X1 U20442 ( .A1(n18134), .A2(n17298), .B1(n17283), .B2(n17282), .C1(
        n17295), .C2(n17281), .ZN(P3_U2730) );
  INV_X1 U20443 ( .A(n17284), .ZN(n17290) );
  AOI21_X1 U20444 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n17303), .A(n17290), .ZN(
        n17286) );
  OAI222_X1 U20445 ( .A1(n18129), .A2(n17298), .B1(n17287), .B2(n17286), .C1(
        n17295), .C2(n17285), .ZN(P3_U2731) );
  INV_X1 U20446 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n18124) );
  AOI21_X1 U20447 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n17303), .A(n17297), .ZN(
        n17289) );
  OAI222_X1 U20448 ( .A1(n18124), .A2(n17298), .B1(n17290), .B2(n17289), .C1(
        n17295), .C2(n17288), .ZN(P3_U2732) );
  INV_X1 U20449 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n18120) );
  NOR2_X1 U20450 ( .A1(n17291), .A2(n17302), .ZN(n17292) );
  AOI21_X1 U20451 ( .B1(P3_EAX_REG_2__SCAN_IN), .B2(n17303), .A(n17292), .ZN(
        n17296) );
  INV_X1 U20452 ( .A(n17293), .ZN(n17294) );
  OAI222_X1 U20453 ( .A1(n18120), .A2(n17298), .B1(n17297), .B2(n17296), .C1(
        n17295), .C2(n17294), .ZN(P3_U2733) );
  AOI22_X1 U20454 ( .A1(n17301), .A2(BUF2_REG_1__SCAN_IN), .B1(n17300), .B2(
        n17299), .ZN(n17306) );
  OAI211_X1 U20455 ( .C1(P3_EAX_REG_1__SCAN_IN), .C2(n17304), .A(n17303), .B(
        n17302), .ZN(n17305) );
  NAND2_X1 U20456 ( .A1(n17306), .A2(n17305), .ZN(P3_U2734) );
  NOR2_X2 U20457 ( .A1(n18726), .A2(n17781), .ZN(n18769) );
  NOR2_X4 U20458 ( .A1(n18769), .A2(n17325), .ZN(n17339) );
  AND2_X1 U20459 ( .A1(n17339), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  INV_X1 U20460 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n17377) );
  AOI22_X1 U20461 ( .A1(n18769), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n17339), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n17309) );
  OAI21_X1 U20462 ( .B1(n17377), .B2(n17324), .A(n17309), .ZN(P3_U2737) );
  INV_X1 U20463 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n17375) );
  AOI22_X1 U20464 ( .A1(P3_DATAO_REG_29__SCAN_IN), .A2(n17339), .B1(n18769), 
        .B2(P3_UWORD_REG_13__SCAN_IN), .ZN(n17310) );
  OAI21_X1 U20465 ( .B1(n17375), .B2(n17324), .A(n17310), .ZN(P3_U2738) );
  CLKBUF_X1 U20466 ( .A(n18769), .Z(n17342) );
  AOI22_X1 U20467 ( .A1(n17342), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n17339), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n17311) );
  OAI21_X1 U20468 ( .B1(n17373), .B2(n17324), .A(n17311), .ZN(P3_U2739) );
  INV_X1 U20469 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n17371) );
  AOI22_X1 U20470 ( .A1(P3_DATAO_REG_27__SCAN_IN), .A2(n17339), .B1(n18769), 
        .B2(P3_UWORD_REG_11__SCAN_IN), .ZN(n17312) );
  OAI21_X1 U20471 ( .B1(n17371), .B2(n17324), .A(n17312), .ZN(P3_U2740) );
  AOI22_X1 U20472 ( .A1(n17342), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n17339), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n17313) );
  OAI21_X1 U20473 ( .B1(n17369), .B2(n17324), .A(n17313), .ZN(P3_U2741) );
  INV_X1 U20474 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n17367) );
  AOI22_X1 U20475 ( .A1(P3_DATAO_REG_25__SCAN_IN), .A2(n17339), .B1(n18769), 
        .B2(P3_UWORD_REG_9__SCAN_IN), .ZN(n17314) );
  OAI21_X1 U20476 ( .B1(n17367), .B2(n17324), .A(n17314), .ZN(P3_U2742) );
  INV_X1 U20477 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n17365) );
  AOI22_X1 U20478 ( .A1(n17342), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n17339), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n17315) );
  OAI21_X1 U20479 ( .B1(n17365), .B2(n17324), .A(n17315), .ZN(P3_U2743) );
  INV_X1 U20480 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n17363) );
  AOI22_X1 U20481 ( .A1(n17342), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n17339), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n17316) );
  OAI21_X1 U20482 ( .B1(n17363), .B2(n17324), .A(n17316), .ZN(P3_U2744) );
  AOI22_X1 U20483 ( .A1(P3_DATAO_REG_22__SCAN_IN), .A2(n17339), .B1(n18769), 
        .B2(P3_UWORD_REG_6__SCAN_IN), .ZN(n17317) );
  OAI21_X1 U20484 ( .B1(n17361), .B2(n17324), .A(n17317), .ZN(P3_U2745) );
  AOI22_X1 U20485 ( .A1(n17342), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n17339), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n17318) );
  OAI21_X1 U20486 ( .B1(n17359), .B2(n17324), .A(n17318), .ZN(P3_U2746) );
  INV_X1 U20487 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n17357) );
  AOI22_X1 U20488 ( .A1(n17342), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n17339), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n17319) );
  OAI21_X1 U20489 ( .B1(n17357), .B2(n17324), .A(n17319), .ZN(P3_U2747) );
  AOI22_X1 U20490 ( .A1(n17342), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n17339), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n17320) );
  OAI21_X1 U20491 ( .B1(n17355), .B2(n17324), .A(n17320), .ZN(P3_U2748) );
  INV_X1 U20492 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n17353) );
  AOI22_X1 U20493 ( .A1(n17342), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n17339), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n17321) );
  OAI21_X1 U20494 ( .B1(n17353), .B2(n17324), .A(n17321), .ZN(P3_U2749) );
  AOI22_X1 U20495 ( .A1(n17342), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n17339), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n17322) );
  OAI21_X1 U20496 ( .B1(n17351), .B2(n17324), .A(n17322), .ZN(P3_U2750) );
  INV_X1 U20497 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n17349) );
  AOI22_X1 U20498 ( .A1(P3_UWORD_REG_0__SCAN_IN), .A2(n18769), .B1(n17339), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n17323) );
  OAI21_X1 U20499 ( .B1(n17349), .B2(n17324), .A(n17323), .ZN(P3_U2751) );
  AOI22_X1 U20500 ( .A1(n17342), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n17339), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n17326) );
  OAI21_X1 U20501 ( .B1(n17413), .B2(n17344), .A(n17326), .ZN(P3_U2752) );
  AOI22_X1 U20502 ( .A1(n17342), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n17339), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n17327) );
  OAI21_X1 U20503 ( .B1(n17408), .B2(n17344), .A(n17327), .ZN(P3_U2753) );
  INV_X1 U20504 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n17406) );
  AOI22_X1 U20505 ( .A1(n17342), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n17339), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n17328) );
  OAI21_X1 U20506 ( .B1(n17406), .B2(n17344), .A(n17328), .ZN(P3_U2754) );
  AOI22_X1 U20507 ( .A1(n17342), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n17339), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n17329) );
  OAI21_X1 U20508 ( .B1(n17404), .B2(n17344), .A(n17329), .ZN(P3_U2755) );
  AOI22_X1 U20509 ( .A1(n17342), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n17339), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n17330) );
  OAI21_X1 U20510 ( .B1(n17401), .B2(n17344), .A(n17330), .ZN(P3_U2756) );
  AOI22_X1 U20511 ( .A1(n17342), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n17339), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n17331) );
  OAI21_X1 U20512 ( .B1(n17399), .B2(n17344), .A(n17331), .ZN(P3_U2757) );
  INV_X1 U20513 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n17397) );
  AOI22_X1 U20514 ( .A1(n17342), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n17339), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n17332) );
  OAI21_X1 U20515 ( .B1(n17397), .B2(n17344), .A(n17332), .ZN(P3_U2758) );
  AOI22_X1 U20516 ( .A1(n17342), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n17339), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n17333) );
  OAI21_X1 U20517 ( .B1(n17395), .B2(n17344), .A(n17333), .ZN(P3_U2759) );
  AOI22_X1 U20518 ( .A1(P3_DATAO_REG_7__SCAN_IN), .A2(n17339), .B1(n18769), 
        .B2(P3_LWORD_REG_7__SCAN_IN), .ZN(n17334) );
  OAI21_X1 U20519 ( .B1(n17393), .B2(n17344), .A(n17334), .ZN(P3_U2760) );
  AOI22_X1 U20520 ( .A1(n17342), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n17339), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n17335) );
  OAI21_X1 U20521 ( .B1(n17391), .B2(n17344), .A(n17335), .ZN(P3_U2761) );
  AOI22_X1 U20522 ( .A1(n17342), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n17339), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n17336) );
  OAI21_X1 U20523 ( .B1(n17389), .B2(n17344), .A(n17336), .ZN(P3_U2762) );
  AOI22_X1 U20524 ( .A1(n17342), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n17339), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n17337) );
  OAI21_X1 U20525 ( .B1(n17387), .B2(n17344), .A(n17337), .ZN(P3_U2763) );
  INV_X1 U20526 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n17385) );
  AOI22_X1 U20527 ( .A1(n17342), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n17339), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n17338) );
  OAI21_X1 U20528 ( .B1(n17385), .B2(n17344), .A(n17338), .ZN(P3_U2764) );
  AOI22_X1 U20529 ( .A1(n17342), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n17339), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n17340) );
  OAI21_X1 U20530 ( .B1(n17383), .B2(n17344), .A(n17340), .ZN(P3_U2765) );
  INV_X1 U20531 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n17381) );
  AOI22_X1 U20532 ( .A1(n17342), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n17339), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n17341) );
  OAI21_X1 U20533 ( .B1(n17381), .B2(n17344), .A(n17341), .ZN(P3_U2766) );
  AOI22_X1 U20534 ( .A1(n17342), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n17339), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n17343) );
  OAI21_X1 U20535 ( .B1(n17379), .B2(n17344), .A(n17343), .ZN(P3_U2767) );
  AOI211_X1 U20536 ( .C1(n18760), .C2(n18761), .A(n17346), .B(n17345), .ZN(
        n17347) );
  INV_X2 U20537 ( .A(n17347), .ZN(n17409) );
  AOI22_X1 U20538 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17410), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n17409), .ZN(n17348) );
  OAI21_X1 U20539 ( .B1(n17349), .B2(n17412), .A(n17348), .ZN(P3_U2768) );
  AOI22_X1 U20540 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17410), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n17409), .ZN(n17350) );
  OAI21_X1 U20541 ( .B1(n17351), .B2(n17412), .A(n17350), .ZN(P3_U2769) );
  AOI22_X1 U20542 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17410), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n17409), .ZN(n17352) );
  OAI21_X1 U20543 ( .B1(n17353), .B2(n17412), .A(n17352), .ZN(P3_U2770) );
  AOI22_X1 U20544 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17402), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n17409), .ZN(n17354) );
  OAI21_X1 U20545 ( .B1(n17355), .B2(n17412), .A(n17354), .ZN(P3_U2771) );
  AOI22_X1 U20546 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17402), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n17409), .ZN(n17356) );
  OAI21_X1 U20547 ( .B1(n17357), .B2(n17412), .A(n17356), .ZN(P3_U2772) );
  AOI22_X1 U20548 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17402), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n17409), .ZN(n17358) );
  OAI21_X1 U20549 ( .B1(n17359), .B2(n17412), .A(n17358), .ZN(P3_U2773) );
  AOI22_X1 U20550 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17402), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n17409), .ZN(n17360) );
  OAI21_X1 U20551 ( .B1(n17361), .B2(n17412), .A(n17360), .ZN(P3_U2774) );
  AOI22_X1 U20552 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17402), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n17409), .ZN(n17362) );
  OAI21_X1 U20553 ( .B1(n17363), .B2(n17412), .A(n17362), .ZN(P3_U2775) );
  AOI22_X1 U20554 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17402), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n17409), .ZN(n17364) );
  OAI21_X1 U20555 ( .B1(n17365), .B2(n17412), .A(n17364), .ZN(P3_U2776) );
  AOI22_X1 U20556 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17402), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n17409), .ZN(n17366) );
  OAI21_X1 U20557 ( .B1(n17367), .B2(n17412), .A(n17366), .ZN(P3_U2777) );
  AOI22_X1 U20558 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17402), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n17409), .ZN(n17368) );
  OAI21_X1 U20559 ( .B1(n17369), .B2(n17412), .A(n17368), .ZN(P3_U2778) );
  AOI22_X1 U20560 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17402), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n17409), .ZN(n17370) );
  OAI21_X1 U20561 ( .B1(n17371), .B2(n17412), .A(n17370), .ZN(P3_U2779) );
  AOI22_X1 U20562 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17410), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n17409), .ZN(n17372) );
  OAI21_X1 U20563 ( .B1(n17373), .B2(n17412), .A(n17372), .ZN(P3_U2780) );
  AOI22_X1 U20564 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17410), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n17409), .ZN(n17374) );
  OAI21_X1 U20565 ( .B1(n17375), .B2(n17412), .A(n17374), .ZN(P3_U2781) );
  AOI22_X1 U20566 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17410), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n17409), .ZN(n17376) );
  OAI21_X1 U20567 ( .B1(n17377), .B2(n17412), .A(n17376), .ZN(P3_U2782) );
  AOI22_X1 U20568 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17410), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n17409), .ZN(n17378) );
  OAI21_X1 U20569 ( .B1(n17379), .B2(n17412), .A(n17378), .ZN(P3_U2783) );
  AOI22_X1 U20570 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17410), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n17409), .ZN(n17380) );
  OAI21_X1 U20571 ( .B1(n17381), .B2(n17412), .A(n17380), .ZN(P3_U2784) );
  AOI22_X1 U20572 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17410), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n17409), .ZN(n17382) );
  OAI21_X1 U20573 ( .B1(n17383), .B2(n17412), .A(n17382), .ZN(P3_U2785) );
  AOI22_X1 U20574 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17410), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n17409), .ZN(n17384) );
  OAI21_X1 U20575 ( .B1(n17385), .B2(n17412), .A(n17384), .ZN(P3_U2786) );
  AOI22_X1 U20576 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17410), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n17409), .ZN(n17386) );
  OAI21_X1 U20577 ( .B1(n17387), .B2(n17412), .A(n17386), .ZN(P3_U2787) );
  AOI22_X1 U20578 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17410), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n17409), .ZN(n17388) );
  OAI21_X1 U20579 ( .B1(n17389), .B2(n17412), .A(n17388), .ZN(P3_U2788) );
  AOI22_X1 U20580 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17410), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n17409), .ZN(n17390) );
  OAI21_X1 U20581 ( .B1(n17391), .B2(n17412), .A(n17390), .ZN(P3_U2789) );
  AOI22_X1 U20582 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17410), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n17409), .ZN(n17392) );
  OAI21_X1 U20583 ( .B1(n17393), .B2(n17412), .A(n17392), .ZN(P3_U2790) );
  AOI22_X1 U20584 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17410), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n17409), .ZN(n17394) );
  OAI21_X1 U20585 ( .B1(n17395), .B2(n17412), .A(n17394), .ZN(P3_U2791) );
  AOI22_X1 U20586 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17410), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n17409), .ZN(n17396) );
  OAI21_X1 U20587 ( .B1(n17397), .B2(n17412), .A(n17396), .ZN(P3_U2792) );
  AOI22_X1 U20588 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17402), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n17409), .ZN(n17398) );
  OAI21_X1 U20589 ( .B1(n17399), .B2(n17412), .A(n17398), .ZN(P3_U2793) );
  AOI22_X1 U20590 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17410), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n17409), .ZN(n17400) );
  OAI21_X1 U20591 ( .B1(n17401), .B2(n17412), .A(n17400), .ZN(P3_U2794) );
  AOI22_X1 U20592 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17402), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n17409), .ZN(n17403) );
  OAI21_X1 U20593 ( .B1(n17404), .B2(n17412), .A(n17403), .ZN(P3_U2795) );
  AOI22_X1 U20594 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17410), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n17409), .ZN(n17405) );
  OAI21_X1 U20595 ( .B1(n17406), .B2(n17412), .A(n17405), .ZN(P3_U2796) );
  AOI22_X1 U20596 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17410), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n17409), .ZN(n17407) );
  OAI21_X1 U20597 ( .B1(n17408), .B2(n17412), .A(n17407), .ZN(P3_U2797) );
  AOI22_X1 U20598 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17410), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n17409), .ZN(n17411) );
  OAI21_X1 U20599 ( .B1(n17413), .B2(n17412), .A(n17411), .ZN(P3_U2798) );
  INV_X1 U20600 ( .A(n17781), .ZN(n17459) );
  INV_X1 U20601 ( .A(n17735), .ZN(n17683) );
  OAI21_X1 U20602 ( .B1(n17414), .B2(n17683), .A(n17780), .ZN(n17415) );
  AOI21_X1 U20603 ( .B1(n17459), .B2(n17416), .A(n17415), .ZN(n17445) );
  OAI21_X1 U20604 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17500), .A(
        n17445), .ZN(n17432) );
  AOI211_X1 U20605 ( .C1(n17419), .C2(n17418), .A(n17417), .B(n17659), .ZN(
        n17426) );
  NAND2_X1 U20606 ( .A1(n17444), .A2(n17632), .ZN(n17474) );
  NOR2_X1 U20607 ( .A1(n17420), .A2(n17474), .ZN(n17435) );
  NAND2_X1 U20608 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17421) );
  OAI211_X1 U20609 ( .C1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A(n17435), .B(n17421), .ZN(n17422) );
  OAI211_X1 U20610 ( .C1(n17591), .C2(n17424), .A(n17423), .B(n17422), .ZN(
        n17425) );
  AOI211_X1 U20611 ( .C1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .C2(n17432), .A(
        n17426), .B(n17425), .ZN(n17429) );
  NOR2_X1 U20612 ( .A1(n17773), .A2(n17696), .ZN(n17626) );
  INV_X1 U20613 ( .A(n17626), .ZN(n17527) );
  OAI22_X1 U20614 ( .A1(n17785), .A2(n17791), .B1(n17616), .B2(n17427), .ZN(
        n17450) );
  OR2_X1 U20615 ( .A1(n17800), .A2(n17450), .ZN(n17437) );
  NAND3_X1 U20616 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17527), .A3(
        n17437), .ZN(n17428) );
  OAI211_X1 U20617 ( .C1(n17430), .C2(n17436), .A(n17429), .B(n17428), .ZN(
        P3_U2802) );
  AOI22_X1 U20618 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n17432), .B1(
        n17638), .B2(n17431), .ZN(n17441) );
  XOR2_X1 U20619 ( .A(n17694), .B(n17434), .Z(n17797) );
  AOI22_X1 U20620 ( .A1(n17695), .A2(n17797), .B1(n17435), .B2(n10010), .ZN(
        n17440) );
  INV_X1 U20621 ( .A(n17436), .ZN(n17438) );
  OAI21_X1 U20622 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n17438), .A(
        n17437), .ZN(n17439) );
  NAND2_X1 U20623 ( .A1(n18093), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n17798) );
  NAND4_X1 U20624 ( .A1(n17441), .A2(n17440), .A3(n17439), .A4(n17798), .ZN(
        P3_U2803) );
  AOI21_X1 U20625 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17443), .A(
        n17442), .ZN(n17807) );
  INV_X1 U20626 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n18695) );
  NOR2_X1 U20627 ( .A1(n18091), .A2(n18695), .ZN(n17804) );
  NAND3_X1 U20628 ( .A1(n18497), .A2(n17444), .A3(n17456), .ZN(n17446) );
  AOI21_X1 U20629 ( .B1(n17447), .B2(n17446), .A(n17445), .ZN(n17448) );
  AOI211_X1 U20630 ( .C1(n17449), .C2(n17775), .A(n17804), .B(n17448), .ZN(
        n17452) );
  NOR3_X1 U20631 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n17810), .A3(
        n17811), .ZN(n17805) );
  NAND2_X1 U20632 ( .A1(n17863), .A2(n17587), .ZN(n17554) );
  INV_X1 U20633 ( .A(n17554), .ZN(n17538) );
  AOI22_X1 U20634 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n17450), .B1(
        n17805), .B2(n17538), .ZN(n17451) );
  OAI211_X1 U20635 ( .C1(n17807), .C2(n17659), .A(n17452), .B(n17451), .ZN(
        P3_U2804) );
  OAI21_X1 U20636 ( .B1(n17628), .B2(n17454), .A(n17453), .ZN(n17455) );
  XOR2_X1 U20637 ( .A(n17455), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n17823) );
  AOI211_X1 U20638 ( .C1(n17473), .C2(n17462), .A(n17456), .B(n17474), .ZN(
        n17464) );
  NOR2_X1 U20639 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n17500), .ZN(
        n17494) );
  AOI22_X1 U20640 ( .A1(n17459), .A2(n17458), .B1(n18497), .B2(n17457), .ZN(
        n17460) );
  NAND2_X1 U20641 ( .A1(n17460), .A2(n17780), .ZN(n17491) );
  NOR2_X1 U20642 ( .A1(n17494), .A2(n17491), .ZN(n17472) );
  OAI22_X1 U20643 ( .A1(n17472), .A2(n17462), .B1(n17591), .B2(n17461), .ZN(
        n17463) );
  AOI211_X1 U20644 ( .C1(P3_REIP_REG_25__SCAN_IN), .C2(n18093), .A(n17464), 
        .B(n17463), .ZN(n17470) );
  NOR3_X1 U20645 ( .A1(n17811), .A2(n17812), .A3(n17465), .ZN(n17466) );
  XOR2_X1 U20646 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B(n17466), .Z(
        n17819) );
  NOR3_X1 U20647 ( .A1(n17467), .A2(n17811), .A3(n17812), .ZN(n17468) );
  XOR2_X1 U20648 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B(n17468), .Z(
        n17820) );
  AOI22_X1 U20649 ( .A1(n17773), .A2(n17819), .B1(n17696), .B2(n17820), .ZN(
        n17469) );
  OAI211_X1 U20650 ( .C1(n17659), .C2(n17823), .A(n17470), .B(n17469), .ZN(
        P3_U2805) );
  NAND2_X1 U20651 ( .A1(n17471), .A2(n17477), .ZN(n17824) );
  NAND2_X1 U20652 ( .A1(n18093), .A2(P3_REIP_REG_24__SCAN_IN), .ZN(n17837) );
  OAI221_X1 U20653 ( .B1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n17474), .C1(
        n17473), .C2(n17472), .A(n17837), .ZN(n17479) );
  AOI21_X1 U20654 ( .B1(n17919), .B2(n17827), .A(n17616), .ZN(n17486) );
  AOI21_X1 U20655 ( .B1(n17918), .B2(n17827), .A(n17785), .ZN(n17487) );
  NOR2_X1 U20656 ( .A1(n17486), .A2(n17487), .ZN(n17489) );
  AOI21_X1 U20657 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n17476), .A(
        n17475), .ZN(n17825) );
  OAI22_X1 U20658 ( .A1(n17489), .A2(n17477), .B1(n17825), .B2(n17659), .ZN(
        n17478) );
  AOI211_X1 U20659 ( .C1(n17638), .C2(n17480), .A(n17479), .B(n17478), .ZN(
        n17481) );
  OAI21_X1 U20660 ( .B1(n17554), .B2(n17824), .A(n17481), .ZN(P3_U2806) );
  INV_X1 U20661 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n17862) );
  OAI21_X1 U20662 ( .B1(n17483), .B2(n17482), .A(n17502), .ZN(n17484) );
  OAI211_X1 U20663 ( .C1(n17694), .C2(n17862), .A(n17536), .B(n17484), .ZN(
        n17485) );
  XOR2_X1 U20664 ( .A(n17832), .B(n17485), .Z(n17839) );
  AOI22_X1 U20665 ( .A1(n17918), .A2(n17487), .B1(n17919), .B2(n17486), .ZN(
        n17488) );
  OAI22_X1 U20666 ( .A1(n17489), .A2(n17832), .B1(n17488), .B2(n17854), .ZN(
        n17490) );
  AOI21_X1 U20667 ( .B1(n17695), .B2(n17839), .A(n17490), .ZN(n17497) );
  NAND2_X1 U20668 ( .A1(n18093), .A2(P3_REIP_REG_23__SCAN_IN), .ZN(n17843) );
  OAI221_X1 U20669 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17492), .C1(
        P3_PHYADDRPOINTER_REG_23__SCAN_IN), .C2(n18497), .A(n17491), .ZN(
        n17496) );
  OAI21_X1 U20670 ( .B1(n17638), .B2(n17494), .A(n17493), .ZN(n17495) );
  NAND4_X1 U20671 ( .A1(n17497), .A2(n17843), .A3(n17496), .A4(n17495), .ZN(
        P3_U2807) );
  OAI21_X1 U20672 ( .B1(n17498), .B2(n17781), .A(n17780), .ZN(n17499) );
  AOI21_X1 U20673 ( .B1(n17735), .B2(n17509), .A(n17499), .ZN(n17529) );
  OAI21_X1 U20674 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17500), .A(
        n17529), .ZN(n17517) );
  AOI22_X1 U20675 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n17517), .B1(
        n17638), .B2(n17501), .ZN(n17513) );
  INV_X1 U20676 ( .A(n17502), .ZN(n17503) );
  OAI221_X1 U20677 ( .B1(n17503), .B2(n17851), .C1(n17503), .C2(n17576), .A(
        n17536), .ZN(n17504) );
  XOR2_X1 U20678 ( .A(n17862), .B(n17504), .Z(n17859) );
  NOR2_X1 U20679 ( .A1(n17505), .A2(n17554), .ZN(n17507) );
  OAI22_X1 U20680 ( .A1(n17918), .A2(n17785), .B1(n17919), .B2(n17616), .ZN(
        n17586) );
  AOI21_X1 U20681 ( .B1(n17845), .B2(n17527), .A(n17586), .ZN(n17526) );
  INV_X1 U20682 ( .A(n17526), .ZN(n17506) );
  MUX2_X1 U20683 ( .A(n17507), .B(n17506), .S(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .Z(n17508) );
  AOI21_X1 U20684 ( .B1(n17695), .B2(n17859), .A(n17508), .ZN(n17512) );
  NAND2_X1 U20685 ( .A1(n18093), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n17860) );
  NOR2_X1 U20686 ( .A1(n17580), .A2(n17509), .ZN(n17518) );
  OAI211_X1 U20687 ( .C1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A(n17518), .B(n17510), .ZN(n17511) );
  NAND4_X1 U20688 ( .A1(n17513), .A2(n17512), .A3(n17860), .A4(n17511), .ZN(
        P3_U2808) );
  INV_X1 U20689 ( .A(n17514), .ZN(n17515) );
  OAI22_X1 U20690 ( .A1(n18091), .A2(n18686), .B1(n17591), .B2(n17515), .ZN(
        n17516) );
  AOI221_X1 U20691 ( .B1(n17518), .B2(n20951), .C1(n17517), .C2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(n17516), .ZN(n17524) );
  NOR3_X1 U20692 ( .A1(n10019), .A2(n17628), .A3(n17519), .ZN(n17542) );
  INV_X1 U20693 ( .A(n17520), .ZN(n17562) );
  AOI22_X1 U20694 ( .A1(n17865), .A2(n17542), .B1(n17562), .B2(n17521), .ZN(
        n17522) );
  XOR2_X1 U20695 ( .A(n17525), .B(n17522), .Z(n17868) );
  AND2_X1 U20696 ( .A1(n17525), .A2(n17865), .ZN(n17867) );
  AOI22_X1 U20697 ( .A1(n17695), .A2(n17868), .B1(n17538), .B2(n17867), .ZN(
        n17523) );
  OAI211_X1 U20698 ( .C1(n17526), .C2(n17525), .A(n17524), .B(n17523), .ZN(
        P3_U2809) );
  NAND2_X1 U20699 ( .A1(n17863), .A2(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n17877) );
  AOI21_X1 U20700 ( .B1(n17527), .B2(n17877), .A(n17586), .ZN(n17552) );
  INV_X1 U20701 ( .A(n17528), .ZN(n17531) );
  AOI221_X1 U20702 ( .B1(n17531), .B2(n17530), .C1(n18428), .C2(n17530), .A(
        n17529), .ZN(n17535) );
  AOI21_X1 U20703 ( .B1(n17591), .B2(n17500), .A(n17533), .ZN(n17534) );
  AOI211_X1 U20704 ( .C1(P3_REIP_REG_20__SCAN_IN), .C2(n18093), .A(n17535), 
        .B(n17534), .ZN(n17540) );
  OAI221_X1 U20705 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17561), 
        .C1(n17553), .C2(n17542), .A(n17536), .ZN(n17537) );
  XOR2_X1 U20706 ( .A(n17541), .B(n17537), .Z(n17873) );
  NOR2_X1 U20707 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17553), .ZN(
        n17871) );
  AOI22_X1 U20708 ( .A1(n17695), .A2(n17873), .B1(n17538), .B2(n17871), .ZN(
        n17539) );
  OAI211_X1 U20709 ( .C1(n17552), .C2(n17541), .A(n17540), .B(n17539), .ZN(
        P3_U2810) );
  AOI21_X1 U20710 ( .B1(n17561), .B2(n17562), .A(n17542), .ZN(n17543) );
  XOR2_X1 U20711 ( .A(n17553), .B(n17543), .Z(n17882) );
  AOI21_X1 U20712 ( .B1(n17735), .B2(n17545), .A(n17768), .ZN(n17574) );
  OAI21_X1 U20713 ( .B1(n17544), .B2(n17781), .A(n17574), .ZN(n17558) );
  AOI22_X1 U20714 ( .A1(n18093), .A2(P3_REIP_REG_19__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n17558), .ZN(n17548) );
  NOR2_X1 U20715 ( .A1(n17580), .A2(n17545), .ZN(n17560) );
  OAI211_X1 U20716 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n17560), .B(n17546), .ZN(n17547) );
  OAI211_X1 U20717 ( .C1(n17591), .C2(n17549), .A(n17548), .B(n17547), .ZN(
        n17550) );
  AOI21_X1 U20718 ( .B1(n17695), .B2(n17882), .A(n17550), .ZN(n17551) );
  OAI221_X1 U20719 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17554), 
        .C1(n17553), .C2(n17552), .A(n17551), .ZN(P3_U2811) );
  INV_X1 U20720 ( .A(n17555), .ZN(n17888) );
  AOI21_X1 U20721 ( .B1(n17587), .B2(n17888), .A(n17586), .ZN(n17570) );
  OAI22_X1 U20722 ( .A1(n18091), .A2(n18679), .B1(n17591), .B2(n17556), .ZN(
        n17557) );
  AOI221_X1 U20723 ( .B1(n17560), .B2(n17559), .C1(n17558), .C2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(n17557), .ZN(n17565) );
  AOI21_X1 U20724 ( .B1(n17694), .B2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n17561), .ZN(n17563) );
  XOR2_X1 U20725 ( .A(n17563), .B(n17562), .Z(n17897) );
  NOR2_X1 U20726 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17888), .ZN(
        n17896) );
  AOI22_X1 U20727 ( .A1(n17695), .A2(n17897), .B1(n17587), .B2(n17896), .ZN(
        n17564) );
  OAI211_X1 U20728 ( .C1(n17570), .C2(n10019), .A(n17565), .B(n17564), .ZN(
        P3_U2812) );
  AOI21_X1 U20729 ( .B1(n17566), .B2(n18497), .A(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17575) );
  OAI21_X1 U20730 ( .B1(n17568), .B2(n17893), .A(n17567), .ZN(n17901) );
  AOI21_X1 U20731 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17587), .A(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17569) );
  OAI22_X1 U20732 ( .A1(n17765), .A2(n17571), .B1(n17570), .B2(n17569), .ZN(
        n17572) );
  AOI21_X1 U20733 ( .B1(n17695), .B2(n17901), .A(n17572), .ZN(n17573) );
  NAND2_X1 U20734 ( .A1(n18093), .A2(P3_REIP_REG_17__SCAN_IN), .ZN(n17904) );
  OAI211_X1 U20735 ( .C1(n17575), .C2(n17574), .A(n17573), .B(n17904), .ZN(
        P3_U2813) );
  NOR2_X1 U20736 ( .A1(n17628), .A2(n17692), .ZN(n17669) );
  INV_X1 U20737 ( .A(n17669), .ZN(n17657) );
  OAI22_X1 U20738 ( .A1(n17694), .A2(n17576), .B1(n17895), .B2(n17657), .ZN(
        n17577) );
  XOR2_X1 U20739 ( .A(n17912), .B(n17577), .Z(n17917) );
  AOI21_X1 U20740 ( .B1(n17735), .B2(n17579), .A(n17768), .ZN(n17604) );
  OAI21_X1 U20741 ( .B1(n17578), .B2(n17781), .A(n17604), .ZN(n17593) );
  AOI22_X1 U20742 ( .A1(n18093), .A2(P3_REIP_REG_16__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n17593), .ZN(n17583) );
  NOR2_X1 U20743 ( .A1(n17580), .A2(n17579), .ZN(n17595) );
  OAI211_X1 U20744 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n17595), .B(n17581), .ZN(n17582) );
  OAI211_X1 U20745 ( .C1(n17591), .C2(n17584), .A(n17583), .B(n17582), .ZN(
        n17585) );
  AOI221_X1 U20746 ( .B1(n17587), .B2(n17912), .C1(n17586), .C2(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A(n17585), .ZN(n17588) );
  OAI21_X1 U20747 ( .B1(n17917), .B2(n17659), .A(n17588), .ZN(P3_U2814) );
  NOR2_X1 U20748 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17639), .ZN(
        n17611) );
  NOR2_X1 U20749 ( .A1(n17607), .A2(n17657), .ZN(n17612) );
  NOR2_X1 U20750 ( .A1(n17962), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n17617) );
  INV_X1 U20751 ( .A(n17617), .ZN(n17610) );
  OAI221_X1 U20752 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n17611), 
        .C1(n20946), .C2(n17612), .A(n17610), .ZN(n17589) );
  XOR2_X1 U20753 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n17589), .Z(
        n17925) );
  OAI22_X1 U20754 ( .A1(n18091), .A2(n18673), .B1(n17591), .B2(n17590), .ZN(
        n17592) );
  AOI221_X1 U20755 ( .B1(n17595), .B2(n17594), .C1(n17593), .C2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(n17592), .ZN(n17599) );
  NOR2_X1 U20756 ( .A1(n17918), .A2(n17785), .ZN(n17597) );
  OAI21_X1 U20757 ( .B1(n17974), .B2(n17910), .A(n17932), .ZN(n17928) );
  NOR2_X1 U20758 ( .A1(n17919), .A2(n17616), .ZN(n17596) );
  NAND3_X1 U20759 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n17934), .A3(
        n17951), .ZN(n17600) );
  NAND2_X1 U20760 ( .A1(n17932), .A2(n17600), .ZN(n17923) );
  AOI22_X1 U20761 ( .A1(n17597), .A2(n17928), .B1(n17596), .B2(n17923), .ZN(
        n17598) );
  OAI211_X1 U20762 ( .C1(n17659), .C2(n17925), .A(n17599), .B(n17598), .ZN(
        P3_U2815) );
  AND2_X1 U20763 ( .A1(n17934), .A2(n17951), .ZN(n17601) );
  OAI21_X1 U20764 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n17601), .A(
        n17600), .ZN(n17947) );
  NOR2_X1 U20765 ( .A1(n18428), .A2(n17602), .ZN(n17649) );
  AOI21_X1 U20766 ( .B1(n17622), .B2(n17649), .A(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17603) );
  OAI22_X1 U20767 ( .A1(n17765), .A2(n17605), .B1(n17604), .B2(n17603), .ZN(
        n17606) );
  AOI21_X1 U20768 ( .B1(n18093), .B2(P3_REIP_REG_14__SCAN_IN), .A(n17606), 
        .ZN(n17615) );
  INV_X1 U20769 ( .A(n17607), .ZN(n17955) );
  NAND2_X1 U20770 ( .A1(n17955), .A2(n17608), .ZN(n17952) );
  NOR2_X1 U20771 ( .A1(n17974), .A2(n17910), .ZN(n17609) );
  AOI221_X1 U20772 ( .B1(n17938), .B2(n20946), .C1(n17952), .C2(n20946), .A(
        n17609), .ZN(n17944) );
  OAI21_X1 U20773 ( .B1(n17612), .B2(n17611), .A(n17610), .ZN(n17613) );
  XOR2_X1 U20774 ( .A(n17613), .B(n20946), .Z(n17943) );
  AOI22_X1 U20775 ( .A1(n17773), .A2(n17944), .B1(n17695), .B2(n17943), .ZN(
        n17614) );
  OAI211_X1 U20776 ( .C1(n17616), .C2(n17947), .A(n17615), .B(n17614), .ZN(
        P3_U2816) );
  NAND2_X1 U20777 ( .A1(n17966), .A2(n17617), .ZN(n17961) );
  NOR2_X1 U20778 ( .A1(n18091), .A2(n18669), .ZN(n17624) );
  OAI211_X1 U20779 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(n16631), .B(n17632), .ZN(n17621) );
  OAI21_X1 U20780 ( .B1(n16631), .B2(n17683), .A(n17781), .ZN(n17618) );
  AOI21_X1 U20781 ( .B1(n17619), .B2(n17618), .A(n17768), .ZN(n17633) );
  OAI22_X1 U20782 ( .A1(n17622), .A2(n17621), .B1(n17633), .B2(n17620), .ZN(
        n17623) );
  AOI211_X1 U20783 ( .C1(n17638), .C2(n17625), .A(n17624), .B(n17623), .ZN(
        n17631) );
  AOI22_X1 U20784 ( .A1(n17773), .A2(n17974), .B1(n17696), .B2(n17692), .ZN(
        n17679) );
  OAI21_X1 U20785 ( .B1(n17955), .B2(n17626), .A(n17679), .ZN(n17641) );
  AOI22_X1 U20786 ( .A1(n17951), .A2(n17955), .B1(n17962), .B2(n17628), .ZN(
        n17627) );
  AOI21_X1 U20787 ( .B1(n17639), .B2(n17628), .A(n17627), .ZN(n17629) );
  XOR2_X1 U20788 ( .A(n17629), .B(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .Z(
        n17949) );
  AOI22_X1 U20789 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17641), .B1(
        n17695), .B2(n17949), .ZN(n17630) );
  OAI211_X1 U20790 ( .C1(n17680), .C2(n17961), .A(n17631), .B(n17630), .ZN(
        P3_U2817) );
  NAND2_X1 U20791 ( .A1(n17966), .A2(n17962), .ZN(n17644) );
  NAND2_X1 U20792 ( .A1(n16631), .A2(n17632), .ZN(n17635) );
  NAND2_X1 U20793 ( .A1(n18093), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n17968) );
  OAI221_X1 U20794 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n17635), .C1(
        n17634), .C2(n17633), .A(n17968), .ZN(n17636) );
  AOI21_X1 U20795 ( .B1(n17638), .B2(n17637), .A(n17636), .ZN(n17643) );
  NAND2_X1 U20796 ( .A1(n17651), .A2(n17669), .ZN(n17652) );
  OAI21_X1 U20797 ( .B1(n17645), .B2(n17652), .A(n17639), .ZN(n17640) );
  XOR2_X1 U20798 ( .A(n17640), .B(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .Z(
        n17967) );
  AOI22_X1 U20799 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17641), .B1(
        n17695), .B2(n17967), .ZN(n17642) );
  OAI211_X1 U20800 ( .C1(n17680), .C2(n17644), .A(n17643), .B(n17642), .ZN(
        P3_U2818) );
  NAND2_X1 U20801 ( .A1(n17651), .A2(n17645), .ZN(n17983) );
  INV_X1 U20802 ( .A(n17672), .ZN(n17776) );
  NOR2_X1 U20803 ( .A1(n18428), .A2(n17646), .ZN(n17667) );
  AOI21_X1 U20804 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n17776), .A(
        n17667), .ZN(n17648) );
  OAI22_X1 U20805 ( .A1(n17649), .A2(n17648), .B1(n17765), .B2(n17647), .ZN(
        n17650) );
  AOI21_X1 U20806 ( .B1(n18093), .B2(P3_REIP_REG_11__SCAN_IN), .A(n17650), 
        .ZN(n17655) );
  OAI21_X1 U20807 ( .B1(n17651), .B2(n17680), .A(n17679), .ZN(n17663) );
  OAI21_X1 U20808 ( .B1(n17656), .B2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n17652), .ZN(n17653) );
  XOR2_X1 U20809 ( .A(n17653), .B(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .Z(
        n17972) );
  AOI22_X1 U20810 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n17663), .B1(
        n17695), .B2(n17972), .ZN(n17654) );
  OAI211_X1 U20811 ( .C1(n17680), .C2(n17983), .A(n17655), .B(n17654), .ZN(
        P3_U2819) );
  NOR3_X1 U20812 ( .A1(n18428), .A2(n17711), .A3(n17722), .ZN(n17703) );
  NAND2_X1 U20813 ( .A1(n17685), .A2(n17703), .ZN(n17674) );
  NOR2_X1 U20814 ( .A1(n17673), .A2(n17674), .ZN(n17671) );
  AOI21_X1 U20815 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n17776), .A(
        n17671), .ZN(n17666) );
  OAI21_X1 U20816 ( .B1(n17680), .B2(n18001), .A(n17986), .ZN(n17662) );
  OAI21_X1 U20817 ( .B1(n18001), .B2(n17657), .A(n17656), .ZN(n17658) );
  XOR2_X1 U20818 ( .A(n17658), .B(n17986), .Z(n17993) );
  OAI22_X1 U20819 ( .A1(n17765), .A2(n17660), .B1(n17993), .B2(n17659), .ZN(
        n17661) );
  AOI21_X1 U20820 ( .B1(n17663), .B2(n17662), .A(n17661), .ZN(n17665) );
  NAND2_X1 U20821 ( .A1(n18093), .A2(P3_REIP_REG_10__SCAN_IN), .ZN(n17664) );
  OAI211_X1 U20822 ( .C1(n17667), .C2(n17666), .A(n17665), .B(n17664), .ZN(
        P3_U2820) );
  NOR2_X1 U20823 ( .A1(n17669), .A2(n17668), .ZN(n17670) );
  XOR2_X1 U20824 ( .A(n17670), .B(n18001), .Z(n17998) );
  AOI211_X1 U20825 ( .C1(n17674), .C2(n17673), .A(n17672), .B(n17671), .ZN(
        n17677) );
  OAI22_X1 U20826 ( .A1(n17765), .A2(n17675), .B1(n18091), .B2(n18661), .ZN(
        n17676) );
  AOI211_X1 U20827 ( .C1(n17695), .C2(n17998), .A(n17677), .B(n17676), .ZN(
        n17678) );
  OAI221_X1 U20828 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17680), .C1(
        n18001), .C2(n17679), .A(n17678), .ZN(P3_U2821) );
  OAI21_X1 U20829 ( .B1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n17682), .A(
        n17681), .ZN(n18020) );
  OAI21_X1 U20830 ( .B1(n17684), .B2(n17683), .A(n17780), .ZN(n17701) );
  AOI211_X1 U20831 ( .C1(n17687), .C2(n17686), .A(n17685), .B(n18428), .ZN(
        n17690) );
  OAI22_X1 U20832 ( .A1(n17765), .A2(n17688), .B1(n18091), .B2(n18660), .ZN(
        n17689) );
  AOI211_X1 U20833 ( .C1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(n17701), .A(
        n17690), .B(n17689), .ZN(n17698) );
  NAND2_X1 U20834 ( .A1(n17692), .A2(n17691), .ZN(n17693) );
  INV_X1 U20835 ( .A(n17693), .ZN(n18016) );
  XOR2_X1 U20836 ( .A(n17694), .B(n17693), .Z(n18014) );
  AOI22_X1 U20837 ( .A1(n17696), .A2(n18016), .B1(n17695), .B2(n18014), .ZN(
        n17697) );
  OAI211_X1 U20838 ( .C1(n17785), .C2(n18020), .A(n17698), .B(n17697), .ZN(
        P3_U2822) );
  OAI21_X1 U20839 ( .B1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n17700), .A(
        n17699), .ZN(n18030) );
  NOR2_X1 U20840 ( .A1(n18091), .A2(n18657), .ZN(n18021) );
  AOI221_X1 U20841 ( .B1(n17703), .B2(n17702), .C1(n17701), .C2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A(n18021), .ZN(n17710) );
  AOI21_X1 U20842 ( .B1(n17706), .B2(n17705), .A(n17704), .ZN(n17707) );
  XOR2_X1 U20843 ( .A(n17707), .B(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .Z(
        n18027) );
  AOI22_X1 U20844 ( .A1(n17773), .A2(n18027), .B1(n17708), .B2(n17775), .ZN(
        n17709) );
  OAI211_X1 U20845 ( .C1(n17784), .C2(n18030), .A(n17710), .B(n17709), .ZN(
        P3_U2823) );
  OAI21_X1 U20846 ( .B1(n17711), .B2(n18428), .A(n17776), .ZN(n17729) );
  NOR2_X1 U20847 ( .A1(n18428), .A2(n17711), .ZN(n17720) );
  OAI21_X1 U20848 ( .B1(n17714), .B2(n17713), .A(n17712), .ZN(n18034) );
  OAI22_X1 U20849 ( .A1(n17784), .A2(n18034), .B1(n18091), .B2(n18655), .ZN(
        n17719) );
  OAI21_X1 U20850 ( .B1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n17716), .A(
        n17715), .ZN(n18033) );
  OAI22_X1 U20851 ( .A1(n17765), .A2(n17717), .B1(n17785), .B2(n18033), .ZN(
        n17718) );
  AOI211_X1 U20852 ( .C1(n17720), .C2(n17722), .A(n17719), .B(n17718), .ZN(
        n17721) );
  OAI21_X1 U20853 ( .B1(n17722), .B2(n17729), .A(n17721), .ZN(P3_U2824) );
  OAI21_X1 U20854 ( .B1(n17725), .B2(n17724), .A(n17723), .ZN(n18040) );
  AOI21_X1 U20855 ( .B1(n17726), .B2(n17780), .A(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17730) );
  OAI21_X1 U20856 ( .B1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n17728), .A(
        n17727), .ZN(n18045) );
  OAI22_X1 U20857 ( .A1(n17730), .A2(n17729), .B1(n17784), .B2(n18045), .ZN(
        n17731) );
  AOI21_X1 U20858 ( .B1(n17732), .B2(n17775), .A(n17731), .ZN(n17733) );
  NAND2_X1 U20859 ( .A1(n18093), .A2(P3_REIP_REG_5__SCAN_IN), .ZN(n18039) );
  OAI211_X1 U20860 ( .C1(n17785), .C2(n18040), .A(n17733), .B(n18039), .ZN(
        P3_U2825) );
  AOI21_X1 U20861 ( .B1(n17735), .B2(n17734), .A(n17768), .ZN(n17754) );
  OAI21_X1 U20862 ( .B1(n17738), .B2(n17737), .A(n17736), .ZN(n17739) );
  XOR2_X1 U20863 ( .A(n17739), .B(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .Z(
        n18053) );
  OAI22_X1 U20864 ( .A1(n17785), .A2(n18053), .B1(n18091), .B2(n18651), .ZN(
        n17745) );
  OAI21_X1 U20865 ( .B1(n17742), .B2(n17741), .A(n17740), .ZN(n18047) );
  OAI22_X1 U20866 ( .A1(n17765), .A2(n17743), .B1(n17784), .B2(n18047), .ZN(
        n17744) );
  AOI211_X1 U20867 ( .C1(n18497), .C2(n17746), .A(n17745), .B(n17744), .ZN(
        n17747) );
  OAI21_X1 U20868 ( .B1(n17754), .B2(n20959), .A(n17747), .ZN(P3_U2826) );
  OAI21_X1 U20869 ( .B1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n17749), .A(
        n17748), .ZN(n18058) );
  AOI21_X1 U20870 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n17780), .A(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17753) );
  OAI21_X1 U20871 ( .B1(n17752), .B2(n17751), .A(n17750), .ZN(n18062) );
  OAI22_X1 U20872 ( .A1(n17754), .A2(n17753), .B1(n17785), .B2(n18062), .ZN(
        n17755) );
  AOI21_X1 U20873 ( .B1(n17756), .B2(n17775), .A(n17755), .ZN(n17757) );
  NAND2_X1 U20874 ( .A1(n18093), .A2(P3_REIP_REG_3__SCAN_IN), .ZN(n18057) );
  OAI211_X1 U20875 ( .C1(n17784), .C2(n18058), .A(n17757), .B(n18057), .ZN(
        P3_U2827) );
  OAI21_X1 U20876 ( .B1(n17760), .B2(n17759), .A(n17758), .ZN(n18073) );
  OAI21_X1 U20877 ( .B1(n17763), .B2(n17762), .A(n17761), .ZN(n18077) );
  OAI22_X1 U20878 ( .A1(n17765), .A2(n17764), .B1(n17784), .B2(n18077), .ZN(
        n17766) );
  AOI221_X1 U20879 ( .B1(n17768), .B2(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .C1(
        n18497), .C2(n17767), .A(n17766), .ZN(n17769) );
  NAND2_X1 U20880 ( .A1(n18093), .A2(P3_REIP_REG_2__SCAN_IN), .ZN(n18075) );
  OAI211_X1 U20881 ( .C1(n17785), .C2(n18073), .A(n17769), .B(n18075), .ZN(
        P3_U2828) );
  OAI21_X1 U20882 ( .B1(n17771), .B2(n17779), .A(n17770), .ZN(n18088) );
  NAND2_X1 U20883 ( .A1(n18742), .A2(n10241), .ZN(n17772) );
  XNOR2_X1 U20884 ( .A(n17772), .B(n17771), .ZN(n18081) );
  AOI22_X1 U20885 ( .A1(n17773), .A2(n18081), .B1(n18093), .B2(
        P3_REIP_REG_1__SCAN_IN), .ZN(n17778) );
  AOI22_X1 U20886 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17776), .B1(
        n17775), .B2(n17774), .ZN(n17777) );
  OAI211_X1 U20887 ( .C1(n17784), .C2(n18088), .A(n17778), .B(n17777), .ZN(
        P3_U2829) );
  AOI21_X1 U20888 ( .B1(n10241), .B2(n18742), .A(n17779), .ZN(n18098) );
  INV_X1 U20889 ( .A(n18098), .ZN(n18096) );
  NAND3_X1 U20890 ( .A1(n18726), .A2(n17781), .A3(n17780), .ZN(n17782) );
  AOI22_X1 U20891 ( .A1(n18093), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17782), .ZN(n17783) );
  OAI221_X1 U20892 ( .B1(n18098), .B2(n17785), .C1(n18096), .C2(n17784), .A(
        n17783), .ZN(P3_U2830) );
  NAND2_X1 U20893 ( .A1(n18089), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17795) );
  NOR2_X1 U20894 ( .A1(n18742), .A2(n17887), .ZN(n17907) );
  OAI211_X1 U20895 ( .C1(n18563), .C2(n17907), .A(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n17851), .ZN(n17786) );
  OAI21_X1 U20896 ( .B1(n17887), .B2(n17786), .A(n18068), .ZN(n17830) );
  OAI21_X1 U20897 ( .B1(n17892), .B2(n17787), .A(n17830), .ZN(n17808) );
  NAND2_X1 U20898 ( .A1(n17788), .A2(n18068), .ZN(n17789) );
  OAI211_X1 U20899 ( .C1(n17791), .C2(n18072), .A(n17790), .B(n17789), .ZN(
        n17792) );
  AOI211_X1 U20900 ( .C1(n17850), .C2(n17793), .A(n17808), .B(n17792), .ZN(
        n17802) );
  AOI22_X1 U20901 ( .A1(n17795), .A2(n17794), .B1(n17802), .B2(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n17796) );
  AOI21_X1 U20902 ( .B1(n18015), .B2(n17797), .A(n17796), .ZN(n17799) );
  OAI211_X1 U20903 ( .C1(n18046), .C2(n17800), .A(n17799), .B(n17798), .ZN(
        P3_U2835) );
  INV_X1 U20904 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17801) );
  AOI211_X1 U20905 ( .C1(n17802), .C2(n18089), .A(n18093), .B(n17801), .ZN(
        n17803) );
  AOI211_X1 U20906 ( .C1(n17805), .C2(n17872), .A(n17804), .B(n17803), .ZN(
        n17806) );
  OAI21_X1 U20907 ( .B1(n17807), .B2(n17992), .A(n17806), .ZN(P3_U2836) );
  NOR2_X1 U20908 ( .A1(n18091), .A2(n18693), .ZN(n17818) );
  NOR3_X1 U20909 ( .A1(n17810), .A2(n17809), .A3(n17808), .ZN(n17816) );
  NOR2_X1 U20910 ( .A1(n17812), .A2(n17811), .ZN(n17814) );
  AOI21_X1 U20911 ( .B1(n17814), .B2(n17813), .A(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17815) );
  NOR3_X1 U20912 ( .A1(n18084), .A2(n17816), .A3(n17815), .ZN(n17817) );
  AOI211_X1 U20913 ( .C1(n18085), .C2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n17818), .B(n17817), .ZN(n17822) );
  AOI22_X1 U20914 ( .A1(n18017), .A2(n17820), .B1(n18082), .B2(n17819), .ZN(
        n17821) );
  OAI211_X1 U20915 ( .C1(n17992), .C2(n17823), .A(n17822), .B(n17821), .ZN(
        P3_U2837) );
  INV_X1 U20916 ( .A(n17872), .ZN(n17886) );
  OAI22_X1 U20917 ( .A1(n17825), .A2(n17992), .B1(n17886), .B2(n17824), .ZN(
        n17826) );
  INV_X1 U20918 ( .A(n17826), .ZN(n17838) );
  NAND2_X1 U20919 ( .A1(n17918), .A2(n17827), .ZN(n17829) );
  NAND2_X1 U20920 ( .A1(n17919), .A2(n17827), .ZN(n17828) );
  AOI22_X1 U20921 ( .A1(n18551), .A2(n17829), .B1(n17850), .B2(n17828), .ZN(
        n17831) );
  NAND3_X1 U20922 ( .A1(n17831), .A2(n18046), .A3(n17830), .ZN(n17835) );
  NOR2_X1 U20923 ( .A1(n17832), .A2(n17835), .ZN(n17834) );
  AOI21_X1 U20924 ( .B1(n17834), .B2(n17833), .A(n18093), .ZN(n17840) );
  OAI211_X1 U20925 ( .C1(n18010), .C2(n17835), .A(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n17840), .ZN(n17836) );
  NAND3_X1 U20926 ( .A1(n17838), .A2(n17837), .A3(n17836), .ZN(P3_U2838) );
  INV_X1 U20927 ( .A(n17839), .ZN(n17844) );
  NOR3_X1 U20928 ( .A1(n18085), .A2(n17846), .A3(n17854), .ZN(n17841) );
  OAI21_X1 U20929 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n17841), .A(
        n17840), .ZN(n17842) );
  OAI211_X1 U20930 ( .C1(n17844), .C2(n17992), .A(n17843), .B(n17842), .ZN(
        P3_U2839) );
  AOI221_X1 U20931 ( .B1(n17846), .B2(n17862), .C1(n17845), .C2(n17862), .A(
        n18084), .ZN(n17858) );
  INV_X1 U20932 ( .A(n17984), .ZN(n17957) );
  OAI22_X1 U20933 ( .A1(n17918), .A2(n18072), .B1(n17919), .B2(n17954), .ZN(
        n17906) );
  AOI221_X1 U20934 ( .B1(n17887), .B2(n17847), .C1(n17877), .C2(n17847), .A(
        n17906), .ZN(n17849) );
  OAI21_X1 U20935 ( .B1(n17888), .B2(n17848), .A(n18567), .ZN(n17889) );
  OAI211_X1 U20936 ( .C1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .C2(n18582), .A(
        n17849), .B(n17889), .ZN(n17875) );
  NOR2_X1 U20937 ( .A1(n18551), .A2(n17850), .ZN(n17874) );
  OAI22_X1 U20938 ( .A1(n18589), .A2(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        n17851), .B2(n17874), .ZN(n17852) );
  NOR2_X1 U20939 ( .A1(n17875), .A2(n17852), .ZN(n17864) );
  INV_X1 U20940 ( .A(n17907), .ZN(n17853) );
  OAI22_X1 U20941 ( .A1(n18587), .A2(n17862), .B1(n17854), .B2(n17853), .ZN(
        n17855) );
  OAI211_X1 U20942 ( .C1(n17957), .C2(n17856), .A(n17864), .B(n17855), .ZN(
        n17857) );
  AOI22_X1 U20943 ( .A1(n18015), .A2(n17859), .B1(n17858), .B2(n17857), .ZN(
        n17861) );
  OAI211_X1 U20944 ( .C1(n18046), .C2(n17862), .A(n17861), .B(n17860), .ZN(
        P3_U2840) );
  OAI221_X1 U20945 ( .B1(n18563), .B2(n17863), .C1(n18563), .C2(n17907), .A(
        n18089), .ZN(n17876) );
  NAND2_X1 U20946 ( .A1(n18582), .A2(n18563), .ZN(n17937) );
  INV_X1 U20947 ( .A(n17937), .ZN(n18083) );
  OAI21_X1 U20948 ( .B1(n17865), .B2(n18083), .A(n17864), .ZN(n17866) );
  OAI21_X1 U20949 ( .B1(n17876), .B2(n17866), .A(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n17870) );
  AOI22_X1 U20950 ( .A1(n18015), .A2(n17868), .B1(n17872), .B2(n17867), .ZN(
        n17869) );
  OAI221_X1 U20951 ( .B1(n18093), .B2(n17870), .C1(n18091), .C2(n18686), .A(
        n17869), .ZN(P3_U2841) );
  AOI22_X1 U20952 ( .A1(n18015), .A2(n17873), .B1(n17872), .B2(n17871), .ZN(
        n17881) );
  INV_X1 U20953 ( .A(n17874), .ZN(n17977) );
  AOI211_X1 U20954 ( .C1(n17877), .C2(n17977), .A(n17876), .B(n17875), .ZN(
        n17878) );
  NOR2_X1 U20955 ( .A1(n18093), .A2(n17878), .ZN(n17883) );
  NOR3_X1 U20956 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18083), .A3(
        n18775), .ZN(n17879) );
  OAI21_X1 U20957 ( .B1(n17883), .B2(n17879), .A(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17880) );
  OAI211_X1 U20958 ( .C1(n18683), .C2(n18091), .A(n17881), .B(n17880), .ZN(
        P3_U2842) );
  AOI22_X1 U20959 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17883), .B1(
        n18015), .B2(n17882), .ZN(n17885) );
  NAND2_X1 U20960 ( .A1(n18093), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n17884) );
  OAI211_X1 U20961 ( .C1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n17886), .A(
        n17885), .B(n17884), .ZN(P3_U2843) );
  NOR2_X1 U20962 ( .A1(n18563), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n18069) );
  NOR3_X1 U20963 ( .A1(n18069), .A2(n17887), .A3(n17912), .ZN(n17891) );
  AOI211_X1 U20964 ( .C1(n17888), .C2(n17977), .A(n18084), .B(n17906), .ZN(
        n17890) );
  OAI211_X1 U20965 ( .C1(n17892), .C2(n17891), .A(n17890), .B(n17889), .ZN(
        n17902) );
  OAI221_X1 U20966 ( .B1(n17902), .B2(n17893), .C1(n17902), .C2(n18068), .A(
        P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17899) );
  OAI22_X1 U20967 ( .A1(n18005), .A2(n18582), .B1(n18064), .B2(n18006), .ZN(
        n18003) );
  INV_X1 U20968 ( .A(n18003), .ZN(n18055) );
  NOR2_X1 U20969 ( .A1(n18055), .A2(n17933), .ZN(n17920) );
  OAI21_X1 U20970 ( .B1(n17920), .B2(n17894), .A(n18089), .ZN(n18002) );
  NOR2_X1 U20971 ( .A1(n17895), .A2(n18002), .ZN(n17913) );
  AOI22_X1 U20972 ( .A1(n18015), .A2(n17897), .B1(n17896), .B2(n17913), .ZN(
        n17898) );
  OAI221_X1 U20973 ( .B1(n18093), .B2(n17899), .C1(n18091), .C2(n18679), .A(
        n17898), .ZN(P3_U2844) );
  NOR2_X1 U20974 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n17912), .ZN(
        n17900) );
  AOI22_X1 U20975 ( .A1(n18015), .A2(n17901), .B1(n17913), .B2(n17900), .ZN(
        n17905) );
  NAND3_X1 U20976 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n18091), .A3(
        n17902), .ZN(n17903) );
  NAND3_X1 U20977 ( .A1(n17905), .A2(n17904), .A3(n17903), .ZN(P3_U2845) );
  NOR2_X1 U20978 ( .A1(n18084), .A2(n17906), .ZN(n17911) );
  AOI21_X1 U20979 ( .B1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n18563), .A(
        n17907), .ZN(n17909) );
  NOR2_X1 U20980 ( .A1(n18589), .A2(n17908), .ZN(n17985) );
  INV_X1 U20981 ( .A(n17985), .ZN(n17994) );
  OAI21_X1 U20982 ( .B1(n17950), .B2(n18582), .A(n17994), .ZN(n17936) );
  AOI211_X1 U20983 ( .C1(n17984), .C2(n17910), .A(n17909), .B(n17936), .ZN(
        n17921) );
  AOI221_X1 U20984 ( .B1(n18008), .B2(n17911), .C1(n17921), .C2(n17911), .A(
        n18093), .ZN(n17914) );
  AOI22_X1 U20985 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n17914), .B1(
        n17913), .B2(n17912), .ZN(n17916) );
  NAND2_X1 U20986 ( .A1(n18093), .A2(P3_REIP_REG_16__SCAN_IN), .ZN(n17915) );
  OAI211_X1 U20987 ( .C1(n17917), .C2(n17992), .A(n17916), .B(n17915), .ZN(
        P3_U2846) );
  NOR2_X1 U20988 ( .A1(n17918), .A2(n18097), .ZN(n17929) );
  NOR2_X1 U20989 ( .A1(n17919), .A2(n17954), .ZN(n17924) );
  NAND2_X1 U20990 ( .A1(n17934), .A2(n17920), .ZN(n17940) );
  AOI221_X1 U20991 ( .B1(n20946), .B2(n17932), .C1(n17940), .C2(n17932), .A(
        n17921), .ZN(n17922) );
  AOI21_X1 U20992 ( .B1(n17924), .B2(n17923), .A(n17922), .ZN(n17926) );
  OAI22_X1 U20993 ( .A1(n18084), .A2(n17926), .B1(n17925), .B2(n17992), .ZN(
        n17927) );
  AOI21_X1 U20994 ( .B1(n17929), .B2(n17928), .A(n17927), .ZN(n17931) );
  NAND2_X1 U20995 ( .A1(n18093), .A2(P3_REIP_REG_15__SCAN_IN), .ZN(n17930) );
  OAI211_X1 U20996 ( .C1(n18046), .C2(n17932), .A(n17931), .B(n17930), .ZN(
        P3_U2847) );
  INV_X1 U20997 ( .A(n18017), .ZN(n17948) );
  NOR2_X1 U20998 ( .A1(n18091), .A2(n18672), .ZN(n17942) );
  NAND3_X1 U20999 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18063) );
  NOR2_X1 U21000 ( .A1(n17933), .A2(n18063), .ZN(n17995) );
  NAND2_X1 U21001 ( .A1(n17955), .A2(n17995), .ZN(n17964) );
  NAND2_X1 U21002 ( .A1(n18587), .A2(n17964), .ZN(n17956) );
  OAI211_X1 U21003 ( .C1(n17957), .C2(n17934), .A(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B(n17956), .ZN(n17935) );
  AOI211_X1 U21004 ( .C1(n17938), .C2(n17937), .A(n17936), .B(n17935), .ZN(
        n17939) );
  AOI211_X1 U21005 ( .C1(n20946), .C2(n17940), .A(n17939), .B(n18084), .ZN(
        n17941) );
  AOI211_X1 U21006 ( .C1(n18085), .C2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n17942), .B(n17941), .ZN(n17946) );
  AOI22_X1 U21007 ( .A1(n18082), .A2(n17944), .B1(n18015), .B2(n17943), .ZN(
        n17945) );
  OAI211_X1 U21008 ( .C1(n17948), .C2(n17947), .A(n17946), .B(n17945), .ZN(
        P3_U2848) );
  AOI22_X1 U21009 ( .A1(n18093), .A2(P3_REIP_REG_13__SCAN_IN), .B1(n18015), 
        .B2(n17949), .ZN(n17960) );
  OAI22_X1 U21010 ( .A1(n17951), .A2(n17954), .B1(n17950), .B2(n18582), .ZN(
        n17973) );
  OAI21_X1 U21011 ( .B1(n17957), .B2(n17966), .A(n17994), .ZN(n17980) );
  AOI211_X1 U21012 ( .C1(n18551), .C2(n17952), .A(n17973), .B(n17980), .ZN(
        n17953) );
  OAI21_X1 U21013 ( .B1(n17955), .B2(n17954), .A(n17953), .ZN(n17963) );
  OAI211_X1 U21014 ( .C1(n17957), .C2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n17956), .B(n18089), .ZN(n17958) );
  OAI211_X1 U21015 ( .C1(n17963), .C2(n17958), .A(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n18091), .ZN(n17959) );
  OAI211_X1 U21016 ( .C1(n17961), .C2(n18002), .A(n17960), .B(n17959), .ZN(
        P3_U2849) );
  AOI211_X1 U21017 ( .C1(n17964), .C2(n18587), .A(n17963), .B(n17962), .ZN(
        n17971) );
  INV_X1 U21018 ( .A(n18002), .ZN(n17965) );
  AOI22_X1 U21019 ( .A1(n17966), .A2(n17965), .B1(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n18089), .ZN(n17970) );
  AOI22_X1 U21020 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18085), .B1(
        n18015), .B2(n17967), .ZN(n17969) );
  OAI211_X1 U21021 ( .C1(n17971), .C2(n17970), .A(n17969), .B(n17968), .ZN(
        P3_U2850) );
  AOI22_X1 U21022 ( .A1(n18093), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n18015), 
        .B2(n17972), .ZN(n17982) );
  AOI21_X1 U21023 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17995), .A(
        n18563), .ZN(n17976) );
  AOI211_X1 U21024 ( .C1(n17974), .C2(n18551), .A(n17973), .B(n18084), .ZN(
        n17975) );
  INV_X1 U21025 ( .A(n17975), .ZN(n17997) );
  AOI211_X1 U21026 ( .C1(n17978), .C2(n17977), .A(n17976), .B(n17997), .ZN(
        n17988) );
  OAI21_X1 U21027 ( .B1(n18563), .B2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n17988), .ZN(n17979) );
  OAI211_X1 U21028 ( .C1(n17980), .C2(n17979), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n18091), .ZN(n17981) );
  OAI211_X1 U21029 ( .C1(n17983), .C2(n18002), .A(n17982), .B(n17981), .ZN(
        P3_U2851) );
  OAI21_X1 U21030 ( .B1(n17985), .B2(n18001), .A(n17984), .ZN(n17987) );
  AOI21_X1 U21031 ( .B1(n17988), .B2(n17987), .A(n17986), .ZN(n17990) );
  NOR3_X1 U21032 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n18001), .A3(
        n18002), .ZN(n17989) );
  AOI221_X1 U21033 ( .B1(P3_REIP_REG_10__SCAN_IN), .B2(n18093), .C1(n17990), 
        .C2(n18091), .A(n17989), .ZN(n17991) );
  OAI21_X1 U21034 ( .B1(n17993), .B2(n17992), .A(n17991), .ZN(P3_U2852) );
  OAI21_X1 U21035 ( .B1(n18563), .B2(n17995), .A(n17994), .ZN(n17996) );
  OAI21_X1 U21036 ( .B1(n17997), .B2(n17996), .A(n18091), .ZN(n18000) );
  AOI22_X1 U21037 ( .A1(n18093), .A2(P3_REIP_REG_9__SCAN_IN), .B1(n18015), 
        .B2(n17998), .ZN(n17999) );
  OAI221_X1 U21038 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18002), .C1(
        n18001), .C2(n18000), .A(n17999), .ZN(P3_U2853) );
  NAND2_X1 U21039 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n18009) );
  NAND3_X1 U21040 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n18089), .A3(
        n18003), .ZN(n18048) );
  NOR2_X1 U21041 ( .A1(n18004), .A2(n18048), .ZN(n18043) );
  NAND2_X1 U21042 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n18043), .ZN(
        n18038) );
  NOR2_X1 U21043 ( .A1(n18009), .A2(n18038), .ZN(n18013) );
  AND2_X1 U21044 ( .A1(n18567), .A2(n18005), .ZN(n18066) );
  AOI211_X1 U21045 ( .C1(n18068), .C2(n18006), .A(n18066), .B(n18069), .ZN(
        n18056) );
  OAI21_X1 U21046 ( .B1(n18008), .B2(n18007), .A(n18056), .ZN(n18031) );
  AOI21_X1 U21047 ( .B1(n18010), .B2(n18009), .A(n18031), .ZN(n18022) );
  OAI21_X1 U21048 ( .B1(n18022), .B2(n18078), .A(n18046), .ZN(n18012) );
  NOR2_X1 U21049 ( .A1(n18091), .A2(n18660), .ZN(n18011) );
  AOI221_X1 U21050 ( .B1(n18013), .B2(n20862), .C1(n18012), .C2(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A(n18011), .ZN(n18019) );
  AOI22_X1 U21051 ( .A1(n18017), .A2(n18016), .B1(n18015), .B2(n18014), .ZN(
        n18018) );
  OAI211_X1 U21052 ( .C1(n18097), .C2(n18020), .A(n18019), .B(n18018), .ZN(
        P3_U2854) );
  AOI21_X1 U21053 ( .B1(n18085), .B2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n18021), .ZN(n18029) );
  INV_X1 U21054 ( .A(n18022), .ZN(n18026) );
  INV_X1 U21055 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n18023) );
  OAI22_X1 U21056 ( .A1(n18084), .A2(n18024), .B1(n18023), .B2(n18038), .ZN(
        n18025) );
  AOI22_X1 U21057 ( .A1(n18082), .A2(n18027), .B1(n18026), .B2(n18025), .ZN(
        n18028) );
  OAI211_X1 U21058 ( .C1(n18095), .C2(n18030), .A(n18029), .B(n18028), .ZN(
        P3_U2855) );
  AOI21_X1 U21059 ( .B1(n18089), .B2(n18031), .A(n18085), .ZN(n18032) );
  INV_X1 U21060 ( .A(n18032), .ZN(n18042) );
  NOR2_X1 U21061 ( .A1(n18091), .A2(n18655), .ZN(n18036) );
  OAI22_X1 U21062 ( .A1(n18095), .A2(n18034), .B1(n18097), .B2(n18033), .ZN(
        n18035) );
  AOI211_X1 U21063 ( .C1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n18042), .A(
        n18036), .B(n18035), .ZN(n18037) );
  OAI21_X1 U21064 ( .B1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n18038), .A(
        n18037), .ZN(P3_U2856) );
  OAI21_X1 U21065 ( .B1(n18097), .B2(n18040), .A(n18039), .ZN(n18041) );
  AOI221_X1 U21066 ( .B1(n18043), .B2(n10013), .C1(n18042), .C2(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A(n18041), .ZN(n18044) );
  OAI21_X1 U21067 ( .B1(n18095), .B2(n18045), .A(n18044), .ZN(P3_U2857) );
  OAI221_X1 U21068 ( .B1(n18078), .B2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .C1(
        n18078), .C2(n18056), .A(n18046), .ZN(n18050) );
  OAI22_X1 U21069 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n18048), .B1(
        n18047), .B2(n18095), .ZN(n18049) );
  AOI21_X1 U21070 ( .B1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n18050), .A(
        n18049), .ZN(n18052) );
  NAND2_X1 U21071 ( .A1(n18093), .A2(P3_REIP_REG_4__SCAN_IN), .ZN(n18051) );
  OAI211_X1 U21072 ( .C1(n18097), .C2(n18053), .A(n18052), .B(n18051), .ZN(
        P3_U2858) );
  AOI221_X1 U21073 ( .B1(n18056), .B2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .C1(
        n18055), .C2(n18054), .A(n18084), .ZN(n18060) );
  OAI21_X1 U21074 ( .B1(n18095), .B2(n18058), .A(n18057), .ZN(n18059) );
  AOI211_X1 U21075 ( .C1(n18085), .C2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n18060), .B(n18059), .ZN(n18061) );
  OAI21_X1 U21076 ( .B1(n18097), .B2(n18062), .A(n18061), .ZN(P3_U2859) );
  INV_X1 U21077 ( .A(n18063), .ZN(n18067) );
  NOR3_X1 U21078 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n18727), .A3(
        n18064), .ZN(n18065) );
  AOI211_X1 U21079 ( .C1(n18067), .C2(n18567), .A(n18066), .B(n18065), .ZN(
        n18071) );
  OAI211_X1 U21080 ( .C1(n18069), .C2(n18727), .A(n18068), .B(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18070) );
  OAI211_X1 U21081 ( .C1(n18073), .C2(n18072), .A(n18071), .B(n18070), .ZN(
        n18074) );
  AOI22_X1 U21082 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n18085), .B1(
        n18089), .B2(n18074), .ZN(n18076) );
  OAI211_X1 U21083 ( .C1(n18077), .C2(n18095), .A(n18076), .B(n18075), .ZN(
        P3_U2860) );
  NOR2_X1 U21084 ( .A1(n18091), .A2(n18749), .ZN(n18080) );
  AOI211_X1 U21085 ( .C1(n18589), .C2(n18742), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B(n18078), .ZN(n18079) );
  AOI211_X1 U21086 ( .C1(n18082), .C2(n18081), .A(n18080), .B(n18079), .ZN(
        n18087) );
  NOR3_X1 U21087 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n18084), .A3(
        n18083), .ZN(n18090) );
  OAI21_X1 U21088 ( .B1(n18085), .B2(n18090), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18086) );
  OAI211_X1 U21089 ( .C1(n18088), .C2(n18095), .A(n18087), .B(n18086), .ZN(
        P3_U2861) );
  AOI21_X1 U21090 ( .B1(n18589), .B2(n18089), .A(n18742), .ZN(n18092) );
  AOI221_X1 U21091 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(n18093), .C1(n18092), 
        .C2(n18091), .A(n18090), .ZN(n18094) );
  OAI221_X1 U21092 ( .B1(n18098), .B2(n18097), .C1(n18096), .C2(n18095), .A(
        n18094), .ZN(P3_U2862) );
  AOI21_X1 U21093 ( .B1(n18101), .B2(n18100), .A(n18099), .ZN(n18614) );
  OAI21_X1 U21094 ( .B1(n18614), .B2(n18149), .A(n18110), .ZN(n18102) );
  OAI221_X1 U21095 ( .B1(n18169), .B2(n18766), .C1(n18169), .C2(n18110), .A(
        n18102), .ZN(P3_U2863) );
  NAND2_X1 U21096 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18326) );
  AOI221_X1 U21097 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18326), .C1(n18104), 
        .C2(n18326), .A(n18103), .ZN(n18109) );
  NOR2_X1 U21098 ( .A1(n18105), .A2(n18594), .ZN(n18106) );
  OAI21_X1 U21099 ( .B1(n18106), .B2(n18191), .A(n18110), .ZN(n18107) );
  AOI22_X1 U21100 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18109), .B1(
        n18107), .B2(n18599), .ZN(P3_U2865) );
  INV_X1 U21101 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18602) );
  NAND2_X1 U21102 ( .A1(n18599), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n18378) );
  INV_X1 U21103 ( .A(n18378), .ZN(n18377) );
  NAND2_X1 U21104 ( .A1(n18602), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n18282) );
  INV_X1 U21105 ( .A(n18282), .ZN(n18281) );
  NOR2_X1 U21106 ( .A1(n18377), .A2(n18281), .ZN(n18108) );
  OAI22_X1 U21107 ( .A1(n18109), .A2(n18602), .B1(n18108), .B2(n18107), .ZN(
        P3_U2866) );
  NOR2_X1 U21108 ( .A1(n20878), .A2(n18110), .ZN(P3_U2867) );
  NOR2_X1 U21109 ( .A1(n18602), .A2(n18326), .ZN(n18495) );
  NAND2_X1 U21110 ( .A1(n18495), .A2(n18169), .ZN(n18156) );
  NAND2_X1 U21111 ( .A1(n18497), .A2(BUF2_REG_16__SCAN_IN), .ZN(n18501) );
  NAND2_X1 U21112 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18430) );
  NAND2_X1 U21113 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18594), .ZN(
        n18330) );
  NOR2_X2 U21114 ( .A1(n18430), .A2(n18330), .ZN(n18543) );
  NAND2_X1 U21115 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n18497), .ZN(n18381) );
  INV_X1 U21116 ( .A(n18381), .ZN(n18493) );
  INV_X1 U21117 ( .A(n18401), .ZN(n18458) );
  AND2_X1 U21118 ( .A1(n18458), .A2(BUF2_REG_0__SCAN_IN), .ZN(n18492) );
  NAND2_X1 U21119 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18593) );
  NOR2_X2 U21120 ( .A1(n18593), .A2(n18430), .ZN(n18545) );
  NAND2_X1 U21121 ( .A1(n18594), .A2(n18169), .ZN(n18595) );
  NOR2_X1 U21122 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18193) );
  INV_X1 U21123 ( .A(n18193), .ZN(n18194) );
  NOR2_X2 U21124 ( .A1(n18595), .A2(n18194), .ZN(n18211) );
  NOR2_X1 U21125 ( .A1(n18545), .A2(n18211), .ZN(n18170) );
  NOR2_X1 U21126 ( .A1(n18623), .A2(n18170), .ZN(n18143) );
  AOI22_X1 U21127 ( .A1(n18543), .A2(n18493), .B1(n18492), .B2(n18143), .ZN(
        n18116) );
  NAND2_X1 U21128 ( .A1(n18539), .A2(n18156), .ZN(n18455) );
  AOI211_X1 U21129 ( .C1(P3_STATE2_REG_3__SCAN_IN), .C2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n18170), .B(n18401), .ZN(
        n18111) );
  AOI21_X1 U21130 ( .B1(n18497), .B2(n18455), .A(n18111), .ZN(n18146) );
  NAND2_X1 U21131 ( .A1(n18113), .A2(n18112), .ZN(n18144) );
  NOR2_X2 U21132 ( .A1(n18114), .A2(n18144), .ZN(n18498) );
  AOI22_X1 U21133 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18146), .B1(
        n18211), .B2(n18498), .ZN(n18115) );
  OAI211_X1 U21134 ( .C1(n18156), .C2(n18501), .A(n18116), .B(n18115), .ZN(
        P3_U2868) );
  NAND2_X1 U21135 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n18497), .ZN(n18507) );
  NAND2_X1 U21136 ( .A1(n18497), .A2(BUF2_REG_17__SCAN_IN), .ZN(n18465) );
  INV_X1 U21137 ( .A(n18465), .ZN(n18503) );
  AND2_X1 U21138 ( .A1(n18458), .A2(BUF2_REG_1__SCAN_IN), .ZN(n18502) );
  AOI22_X1 U21139 ( .A1(n18486), .A2(n18503), .B1(n18143), .B2(n18502), .ZN(
        n18119) );
  NOR2_X2 U21140 ( .A1(n18117), .A2(n18144), .ZN(n18504) );
  AOI22_X1 U21141 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n18146), .B1(
        n18211), .B2(n18504), .ZN(n18118) );
  OAI211_X1 U21142 ( .C1(n18539), .C2(n18507), .A(n18119), .B(n18118), .ZN(
        P3_U2869) );
  NAND2_X1 U21143 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n18497), .ZN(n18513) );
  NAND2_X1 U21144 ( .A1(n18497), .A2(BUF2_REG_18__SCAN_IN), .ZN(n18386) );
  INV_X1 U21145 ( .A(n18386), .ZN(n18509) );
  NOR2_X2 U21146 ( .A1(n18401), .A2(n18120), .ZN(n18508) );
  AOI22_X1 U21147 ( .A1(n18486), .A2(n18509), .B1(n18143), .B2(n18508), .ZN(
        n18123) );
  NOR2_X2 U21148 ( .A1(n18121), .A2(n18144), .ZN(n18510) );
  AOI22_X1 U21149 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n18146), .B1(
        n18211), .B2(n18510), .ZN(n18122) );
  OAI211_X1 U21150 ( .C1(n18539), .C2(n18513), .A(n18123), .B(n18122), .ZN(
        P3_U2870) );
  NAND2_X1 U21151 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n18497), .ZN(n18519) );
  NAND2_X1 U21152 ( .A1(n18497), .A2(BUF2_REG_19__SCAN_IN), .ZN(n18313) );
  INV_X1 U21153 ( .A(n18313), .ZN(n18515) );
  NOR2_X2 U21154 ( .A1(n18401), .A2(n18124), .ZN(n18514) );
  AOI22_X1 U21155 ( .A1(n18486), .A2(n18515), .B1(n18143), .B2(n18514), .ZN(
        n18127) );
  NOR2_X2 U21156 ( .A1(n9817), .A2(n18144), .ZN(n18516) );
  AOI22_X1 U21157 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n18146), .B1(
        n18211), .B2(n18516), .ZN(n18126) );
  OAI211_X1 U21158 ( .C1(n18539), .C2(n18519), .A(n18127), .B(n18126), .ZN(
        P3_U2871) );
  NOR2_X1 U21159 ( .A1(n18128), .A2(n18428), .ZN(n18521) );
  INV_X1 U21160 ( .A(n18521), .ZN(n18473) );
  NAND2_X1 U21161 ( .A1(n18497), .A2(BUF2_REG_20__SCAN_IN), .ZN(n18525) );
  INV_X1 U21162 ( .A(n18525), .ZN(n18470) );
  NOR2_X2 U21163 ( .A1(n18401), .A2(n18129), .ZN(n18520) );
  AOI22_X1 U21164 ( .A1(n18486), .A2(n18470), .B1(n18143), .B2(n18520), .ZN(
        n18132) );
  NOR2_X2 U21165 ( .A1(n18130), .A2(n18144), .ZN(n18522) );
  AOI22_X1 U21166 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n18146), .B1(
        n18211), .B2(n18522), .ZN(n18131) );
  OAI211_X1 U21167 ( .C1(n18539), .C2(n18473), .A(n18132), .B(n18131), .ZN(
        P3_U2872) );
  NOR2_X1 U21168 ( .A1(n18428), .A2(n18133), .ZN(n18527) );
  NAND2_X1 U21169 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n18497), .ZN(n18531) );
  INV_X1 U21170 ( .A(n18531), .ZN(n18474) );
  NOR2_X2 U21171 ( .A1(n18401), .A2(n18134), .ZN(n18526) );
  AOI22_X1 U21172 ( .A1(n18543), .A2(n18474), .B1(n18143), .B2(n18526), .ZN(
        n18137) );
  NOR2_X2 U21173 ( .A1(n18135), .A2(n18144), .ZN(n18528) );
  AOI22_X1 U21174 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n18146), .B1(
        n18211), .B2(n18528), .ZN(n18136) );
  OAI211_X1 U21175 ( .C1(n18156), .C2(n18477), .A(n18137), .B(n18136), .ZN(
        P3_U2873) );
  NAND2_X1 U21176 ( .A1(n18497), .A2(BUF2_REG_22__SCAN_IN), .ZN(n18538) );
  NOR2_X1 U21177 ( .A1(n18138), .A2(n18428), .ZN(n18534) );
  NOR2_X2 U21178 ( .A1(n18401), .A2(n18139), .ZN(n18532) );
  AOI22_X1 U21179 ( .A1(n18543), .A2(n18534), .B1(n18143), .B2(n18532), .ZN(
        n18142) );
  NOR2_X2 U21180 ( .A1(n18140), .A2(n18144), .ZN(n18535) );
  AOI22_X1 U21181 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n18146), .B1(
        n18211), .B2(n18535), .ZN(n18141) );
  OAI211_X1 U21182 ( .C1(n18156), .C2(n18538), .A(n18142), .B(n18141), .ZN(
        P3_U2874) );
  NAND2_X1 U21183 ( .A1(n18497), .A2(BUF2_REG_31__SCAN_IN), .ZN(n18550) );
  NAND2_X1 U21184 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n18497), .ZN(n18490) );
  INV_X1 U21185 ( .A(n18490), .ZN(n18542) );
  NOR2_X2 U21186 ( .A1(n21002), .A2(n18401), .ZN(n18541) );
  AOI22_X1 U21187 ( .A1(n18486), .A2(n18542), .B1(n18143), .B2(n18541), .ZN(
        n18148) );
  NOR2_X2 U21188 ( .A1(n18145), .A2(n18144), .ZN(n18544) );
  AOI22_X1 U21189 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n18146), .B1(
        n18211), .B2(n18544), .ZN(n18147) );
  OAI211_X1 U21190 ( .C1(n18539), .C2(n18550), .A(n18148), .B(n18147), .ZN(
        P3_U2875) );
  INV_X1 U21191 ( .A(n18501), .ZN(n18431) );
  NAND2_X1 U21192 ( .A1(n18594), .A2(n18491), .ZN(n18429) );
  NOR2_X1 U21193 ( .A1(n18194), .A2(n18429), .ZN(n18165) );
  AOI22_X1 U21194 ( .A1(n18545), .A2(n18431), .B1(n18492), .B2(n18165), .ZN(
        n18151) );
  NOR2_X1 U21195 ( .A1(n18401), .A2(n18149), .ZN(n18494) );
  INV_X1 U21196 ( .A(n18494), .ZN(n18328) );
  NOR2_X1 U21197 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18328), .ZN(
        n18425) );
  AOI22_X1 U21198 ( .A1(n18497), .A2(n18495), .B1(n18193), .B2(n18425), .ZN(
        n18166) );
  NOR2_X2 U21199 ( .A1(n18330), .A2(n18194), .ZN(n18227) );
  AOI22_X1 U21200 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n18166), .B1(
        n18498), .B2(n18227), .ZN(n18150) );
  OAI211_X1 U21201 ( .C1(n18156), .C2(n18381), .A(n18151), .B(n18150), .ZN(
        P3_U2876) );
  INV_X1 U21202 ( .A(n18545), .ZN(n18190) );
  INV_X1 U21203 ( .A(n18507), .ZN(n18462) );
  AOI22_X1 U21204 ( .A1(n18486), .A2(n18462), .B1(n18502), .B2(n18165), .ZN(
        n18153) );
  AOI22_X1 U21205 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18166), .B1(
        n18504), .B2(n18227), .ZN(n18152) );
  OAI211_X1 U21206 ( .C1(n18190), .C2(n18465), .A(n18153), .B(n18152), .ZN(
        P3_U2877) );
  AOI22_X1 U21207 ( .A1(n18545), .A2(n18509), .B1(n18508), .B2(n18165), .ZN(
        n18155) );
  AOI22_X1 U21208 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n18166), .B1(
        n18510), .B2(n18227), .ZN(n18154) );
  OAI211_X1 U21209 ( .C1(n18156), .C2(n18513), .A(n18155), .B(n18154), .ZN(
        P3_U2878) );
  INV_X1 U21210 ( .A(n18519), .ZN(n18440) );
  AOI22_X1 U21211 ( .A1(n18486), .A2(n18440), .B1(n18514), .B2(n18165), .ZN(
        n18158) );
  AOI22_X1 U21212 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n18166), .B1(
        n18516), .B2(n18227), .ZN(n18157) );
  OAI211_X1 U21213 ( .C1(n18190), .C2(n18313), .A(n18158), .B(n18157), .ZN(
        P3_U2879) );
  AOI22_X1 U21214 ( .A1(n18486), .A2(n18521), .B1(n18520), .B2(n18165), .ZN(
        n18160) );
  AOI22_X1 U21215 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18166), .B1(
        n18522), .B2(n18227), .ZN(n18159) );
  OAI211_X1 U21216 ( .C1(n18190), .C2(n18525), .A(n18160), .B(n18159), .ZN(
        P3_U2880) );
  AOI22_X1 U21217 ( .A1(n18486), .A2(n18474), .B1(n18526), .B2(n18165), .ZN(
        n18162) );
  AOI22_X1 U21218 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18166), .B1(
        n18528), .B2(n18227), .ZN(n18161) );
  OAI211_X1 U21219 ( .C1(n18190), .C2(n18477), .A(n18162), .B(n18161), .ZN(
        P3_U2881) );
  AOI22_X1 U21220 ( .A1(n18486), .A2(n18534), .B1(n18532), .B2(n18165), .ZN(
        n18164) );
  AOI22_X1 U21221 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n18166), .B1(
        n18535), .B2(n18227), .ZN(n18163) );
  OAI211_X1 U21222 ( .C1(n18190), .C2(n18538), .A(n18164), .B(n18163), .ZN(
        P3_U2882) );
  INV_X1 U21223 ( .A(n18550), .ZN(n18485) );
  AOI22_X1 U21224 ( .A1(n18486), .A2(n18485), .B1(n18541), .B2(n18165), .ZN(
        n18168) );
  AOI22_X1 U21225 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n18166), .B1(
        n18544), .B2(n18227), .ZN(n18167) );
  OAI211_X1 U21226 ( .C1(n18190), .C2(n18490), .A(n18168), .B(n18167), .ZN(
        P3_U2883) );
  INV_X1 U21227 ( .A(n18211), .ZN(n18209) );
  INV_X1 U21228 ( .A(n18227), .ZN(n18236) );
  NOR2_X1 U21229 ( .A1(n18594), .A2(n18194), .ZN(n18237) );
  NAND2_X1 U21230 ( .A1(n18237), .A2(n18169), .ZN(n18248) );
  AOI21_X1 U21231 ( .B1(n18236), .B2(n18248), .A(n18623), .ZN(n18186) );
  AOI22_X1 U21232 ( .A1(n18545), .A2(n18493), .B1(n18492), .B2(n18186), .ZN(
        n18173) );
  OAI21_X1 U21233 ( .B1(n18227), .B2(n18254), .A(n18458), .ZN(n18215) );
  OAI21_X1 U21234 ( .B1(n18170), .B2(n18428), .A(n18215), .ZN(n18171) );
  OAI21_X1 U21235 ( .B1(n18254), .B2(n18716), .A(n18171), .ZN(n18187) );
  AOI22_X1 U21236 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n18187), .B1(
        n18498), .B2(n18254), .ZN(n18172) );
  OAI211_X1 U21237 ( .C1(n18209), .C2(n18501), .A(n18173), .B(n18172), .ZN(
        P3_U2884) );
  AOI22_X1 U21238 ( .A1(n18211), .A2(n18503), .B1(n18502), .B2(n18186), .ZN(
        n18175) );
  AOI22_X1 U21239 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18187), .B1(
        n18504), .B2(n18254), .ZN(n18174) );
  OAI211_X1 U21240 ( .C1(n18190), .C2(n18507), .A(n18175), .B(n18174), .ZN(
        P3_U2885) );
  INV_X1 U21241 ( .A(n18513), .ZN(n18436) );
  AOI22_X1 U21242 ( .A1(n18545), .A2(n18436), .B1(n18508), .B2(n18186), .ZN(
        n18177) );
  AOI22_X1 U21243 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18187), .B1(
        n18510), .B2(n18254), .ZN(n18176) );
  OAI211_X1 U21244 ( .C1(n18209), .C2(n18386), .A(n18177), .B(n18176), .ZN(
        P3_U2886) );
  AOI22_X1 U21245 ( .A1(n18545), .A2(n18440), .B1(n18514), .B2(n18186), .ZN(
        n18179) );
  AOI22_X1 U21246 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18187), .B1(
        n18516), .B2(n18254), .ZN(n18178) );
  OAI211_X1 U21247 ( .C1(n18209), .C2(n18313), .A(n18179), .B(n18178), .ZN(
        P3_U2887) );
  AOI22_X1 U21248 ( .A1(n18545), .A2(n18521), .B1(n18520), .B2(n18186), .ZN(
        n18181) );
  AOI22_X1 U21249 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18187), .B1(
        n18522), .B2(n18254), .ZN(n18180) );
  OAI211_X1 U21250 ( .C1(n18209), .C2(n18525), .A(n18181), .B(n18180), .ZN(
        P3_U2888) );
  AOI22_X1 U21251 ( .A1(n18211), .A2(n18527), .B1(n18526), .B2(n18186), .ZN(
        n18183) );
  AOI22_X1 U21252 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18187), .B1(
        n18528), .B2(n18254), .ZN(n18182) );
  OAI211_X1 U21253 ( .C1(n18190), .C2(n18531), .A(n18183), .B(n18182), .ZN(
        P3_U2889) );
  AOI22_X1 U21254 ( .A1(n18545), .A2(n18534), .B1(n18532), .B2(n18186), .ZN(
        n18185) );
  AOI22_X1 U21255 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18187), .B1(
        n18535), .B2(n18254), .ZN(n18184) );
  OAI211_X1 U21256 ( .C1(n18209), .C2(n18538), .A(n18185), .B(n18184), .ZN(
        P3_U2890) );
  AOI22_X1 U21257 ( .A1(n18211), .A2(n18542), .B1(n18541), .B2(n18186), .ZN(
        n18189) );
  AOI22_X1 U21258 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18187), .B1(
        n18544), .B2(n18254), .ZN(n18188) );
  OAI211_X1 U21259 ( .C1(n18190), .C2(n18550), .A(n18189), .B(n18188), .ZN(
        P3_U2891) );
  OAI21_X1 U21260 ( .B1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n18191), .A(
        n18458), .ZN(n18192) );
  AOI21_X1 U21261 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18593), .A(n18192), 
        .ZN(n18280) );
  NAND2_X1 U21262 ( .A1(n18193), .A2(n18280), .ZN(n18212) );
  AND2_X1 U21263 ( .A1(n18491), .A2(n18237), .ZN(n18210) );
  AOI22_X1 U21264 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n18212), .B1(
        n18492), .B2(n18210), .ZN(n18196) );
  NOR2_X2 U21265 ( .A1(n18593), .A2(n18194), .ZN(n18270) );
  AOI22_X1 U21266 ( .A1(n18211), .A2(n18493), .B1(n18498), .B2(n18270), .ZN(
        n18195) );
  OAI211_X1 U21267 ( .C1(n18501), .C2(n18236), .A(n18196), .B(n18195), .ZN(
        P3_U2892) );
  AOI22_X1 U21268 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n18212), .B1(
        n18502), .B2(n18210), .ZN(n18198) );
  AOI22_X1 U21269 ( .A1(n18211), .A2(n18462), .B1(n18504), .B2(n18270), .ZN(
        n18197) );
  OAI211_X1 U21270 ( .C1(n18465), .C2(n18236), .A(n18198), .B(n18197), .ZN(
        P3_U2893) );
  AOI22_X1 U21271 ( .A1(n18509), .A2(n18227), .B1(n18508), .B2(n18210), .ZN(
        n18200) );
  AOI22_X1 U21272 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n18212), .B1(
        n18510), .B2(n18270), .ZN(n18199) );
  OAI211_X1 U21273 ( .C1(n18209), .C2(n18513), .A(n18200), .B(n18199), .ZN(
        P3_U2894) );
  AOI22_X1 U21274 ( .A1(n18515), .A2(n18227), .B1(n18514), .B2(n18210), .ZN(
        n18202) );
  AOI22_X1 U21275 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n18212), .B1(
        n18516), .B2(n18270), .ZN(n18201) );
  OAI211_X1 U21276 ( .C1(n18209), .C2(n18519), .A(n18202), .B(n18201), .ZN(
        P3_U2895) );
  AOI22_X1 U21277 ( .A1(n18470), .A2(n18227), .B1(n18520), .B2(n18210), .ZN(
        n18204) );
  AOI22_X1 U21278 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n18212), .B1(
        n18522), .B2(n18270), .ZN(n18203) );
  OAI211_X1 U21279 ( .C1(n18209), .C2(n18473), .A(n18204), .B(n18203), .ZN(
        P3_U2896) );
  AOI22_X1 U21280 ( .A1(n18527), .A2(n18227), .B1(n18526), .B2(n18210), .ZN(
        n18206) );
  AOI22_X1 U21281 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n18212), .B1(
        n18528), .B2(n18270), .ZN(n18205) );
  OAI211_X1 U21282 ( .C1(n18209), .C2(n18531), .A(n18206), .B(n18205), .ZN(
        P3_U2897) );
  INV_X1 U21283 ( .A(n18534), .ZN(n18482) );
  INV_X1 U21284 ( .A(n18538), .ZN(n18478) );
  AOI22_X1 U21285 ( .A1(n18478), .A2(n18227), .B1(n18532), .B2(n18210), .ZN(
        n18208) );
  AOI22_X1 U21286 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n18212), .B1(
        n18535), .B2(n18270), .ZN(n18207) );
  OAI211_X1 U21287 ( .C1(n18209), .C2(n18482), .A(n18208), .B(n18207), .ZN(
        P3_U2898) );
  AOI22_X1 U21288 ( .A1(n18211), .A2(n18485), .B1(n18541), .B2(n18210), .ZN(
        n18214) );
  AOI22_X1 U21289 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n18212), .B1(
        n18544), .B2(n18270), .ZN(n18213) );
  OAI211_X1 U21290 ( .C1(n18490), .C2(n18236), .A(n18214), .B(n18213), .ZN(
        P3_U2899) );
  NOR2_X2 U21291 ( .A1(n18595), .A2(n18282), .ZN(n18295) );
  NOR2_X1 U21292 ( .A1(n18270), .A2(n18295), .ZN(n18258) );
  NOR2_X1 U21293 ( .A1(n18623), .A2(n18258), .ZN(n18232) );
  AOI22_X1 U21294 ( .A1(n18431), .A2(n18254), .B1(n18492), .B2(n18232), .ZN(
        n18218) );
  OAI22_X1 U21295 ( .A1(n18258), .A2(n18401), .B1(n18456), .B2(n18215), .ZN(
        n18216) );
  OAI21_X1 U21296 ( .B1(n18295), .B2(n18716), .A(n18216), .ZN(n18233) );
  AOI22_X1 U21297 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n18233), .B1(
        n18498), .B2(n18295), .ZN(n18217) );
  OAI211_X1 U21298 ( .C1(n18381), .C2(n18236), .A(n18218), .B(n18217), .ZN(
        P3_U2900) );
  AOI22_X1 U21299 ( .A1(n18502), .A2(n18232), .B1(n18503), .B2(n18254), .ZN(
        n18220) );
  AOI22_X1 U21300 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18233), .B1(
        n18504), .B2(n18295), .ZN(n18219) );
  OAI211_X1 U21301 ( .C1(n18507), .C2(n18236), .A(n18220), .B(n18219), .ZN(
        P3_U2901) );
  AOI22_X1 U21302 ( .A1(n18509), .A2(n18254), .B1(n18508), .B2(n18232), .ZN(
        n18222) );
  AOI22_X1 U21303 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n18233), .B1(
        n18510), .B2(n18295), .ZN(n18221) );
  OAI211_X1 U21304 ( .C1(n18513), .C2(n18236), .A(n18222), .B(n18221), .ZN(
        P3_U2902) );
  AOI22_X1 U21305 ( .A1(n18515), .A2(n18254), .B1(n18514), .B2(n18232), .ZN(
        n18224) );
  AOI22_X1 U21306 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n18233), .B1(
        n18516), .B2(n18295), .ZN(n18223) );
  OAI211_X1 U21307 ( .C1(n18519), .C2(n18236), .A(n18224), .B(n18223), .ZN(
        P3_U2903) );
  AOI22_X1 U21308 ( .A1(n18521), .A2(n18227), .B1(n18520), .B2(n18232), .ZN(
        n18226) );
  AOI22_X1 U21309 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n18233), .B1(
        n18522), .B2(n18295), .ZN(n18225) );
  OAI211_X1 U21310 ( .C1(n18525), .C2(n18248), .A(n18226), .B(n18225), .ZN(
        P3_U2904) );
  AOI22_X1 U21311 ( .A1(n18526), .A2(n18232), .B1(n18474), .B2(n18227), .ZN(
        n18229) );
  AOI22_X1 U21312 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n18233), .B1(
        n18528), .B2(n18295), .ZN(n18228) );
  OAI211_X1 U21313 ( .C1(n18477), .C2(n18248), .A(n18229), .B(n18228), .ZN(
        P3_U2905) );
  AOI22_X1 U21314 ( .A1(n18478), .A2(n18254), .B1(n18532), .B2(n18232), .ZN(
        n18231) );
  AOI22_X1 U21315 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n18233), .B1(
        n18535), .B2(n18295), .ZN(n18230) );
  OAI211_X1 U21316 ( .C1(n18482), .C2(n18236), .A(n18231), .B(n18230), .ZN(
        P3_U2906) );
  AOI22_X1 U21317 ( .A1(n18542), .A2(n18254), .B1(n18541), .B2(n18232), .ZN(
        n18235) );
  AOI22_X1 U21318 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18233), .B1(
        n18544), .B2(n18295), .ZN(n18234) );
  OAI211_X1 U21319 ( .C1(n18550), .C2(n18236), .A(n18235), .B(n18234), .ZN(
        P3_U2907) );
  NOR2_X1 U21320 ( .A1(n18282), .A2(n18429), .ZN(n18253) );
  AOI22_X1 U21321 ( .A1(n18431), .A2(n18270), .B1(n18492), .B2(n18253), .ZN(
        n18239) );
  AOI22_X1 U21322 ( .A1(n18497), .A2(n18237), .B1(n18281), .B2(n18425), .ZN(
        n18255) );
  NOR2_X2 U21323 ( .A1(n18282), .A2(n18330), .ZN(n18322) );
  AOI22_X1 U21324 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n18255), .B1(
        n18498), .B2(n18322), .ZN(n18238) );
  OAI211_X1 U21325 ( .C1(n18381), .C2(n18248), .A(n18239), .B(n18238), .ZN(
        P3_U2908) );
  AOI22_X1 U21326 ( .A1(n18502), .A2(n18253), .B1(n18503), .B2(n18270), .ZN(
        n18241) );
  AOI22_X1 U21327 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18255), .B1(
        n18504), .B2(n18322), .ZN(n18240) );
  OAI211_X1 U21328 ( .C1(n18507), .C2(n18248), .A(n18241), .B(n18240), .ZN(
        P3_U2909) );
  AOI22_X1 U21329 ( .A1(n18509), .A2(n18270), .B1(n18508), .B2(n18253), .ZN(
        n18243) );
  AOI22_X1 U21330 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n18255), .B1(
        n18510), .B2(n18322), .ZN(n18242) );
  OAI211_X1 U21331 ( .C1(n18513), .C2(n18248), .A(n18243), .B(n18242), .ZN(
        P3_U2910) );
  INV_X1 U21332 ( .A(n18270), .ZN(n18279) );
  AOI22_X1 U21333 ( .A1(n18440), .A2(n18254), .B1(n18514), .B2(n18253), .ZN(
        n18245) );
  AOI22_X1 U21334 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n18255), .B1(
        n18516), .B2(n18322), .ZN(n18244) );
  OAI211_X1 U21335 ( .C1(n18313), .C2(n18279), .A(n18245), .B(n18244), .ZN(
        P3_U2911) );
  AOI22_X1 U21336 ( .A1(n18470), .A2(n18270), .B1(n18520), .B2(n18253), .ZN(
        n18247) );
  AOI22_X1 U21337 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n18255), .B1(
        n18522), .B2(n18322), .ZN(n18246) );
  OAI211_X1 U21338 ( .C1(n18473), .C2(n18248), .A(n18247), .B(n18246), .ZN(
        P3_U2912) );
  AOI22_X1 U21339 ( .A1(n18526), .A2(n18253), .B1(n18474), .B2(n18254), .ZN(
        n18250) );
  AOI22_X1 U21340 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n18255), .B1(
        n18528), .B2(n18322), .ZN(n18249) );
  OAI211_X1 U21341 ( .C1(n18477), .C2(n18279), .A(n18250), .B(n18249), .ZN(
        P3_U2913) );
  AOI22_X1 U21342 ( .A1(n18534), .A2(n18254), .B1(n18532), .B2(n18253), .ZN(
        n18252) );
  AOI22_X1 U21343 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n18255), .B1(
        n18535), .B2(n18322), .ZN(n18251) );
  OAI211_X1 U21344 ( .C1(n18538), .C2(n18279), .A(n18252), .B(n18251), .ZN(
        P3_U2914) );
  AOI22_X1 U21345 ( .A1(n18485), .A2(n18254), .B1(n18541), .B2(n18253), .ZN(
        n18257) );
  AOI22_X1 U21346 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n18255), .B1(
        n18544), .B2(n18322), .ZN(n18256) );
  OAI211_X1 U21347 ( .C1(n18490), .C2(n18279), .A(n18257), .B(n18256), .ZN(
        P3_U2915) );
  INV_X1 U21348 ( .A(n18295), .ZN(n18302) );
  NOR2_X1 U21349 ( .A1(n18322), .A2(n18351), .ZN(n18303) );
  NOR2_X1 U21350 ( .A1(n18623), .A2(n18303), .ZN(n18275) );
  AOI22_X1 U21351 ( .A1(n18493), .A2(n18270), .B1(n18492), .B2(n18275), .ZN(
        n18261) );
  OAI21_X1 U21352 ( .B1(n18258), .B2(n18456), .A(n18303), .ZN(n18259) );
  OAI211_X1 U21353 ( .C1(n18351), .C2(n18716), .A(n18458), .B(n18259), .ZN(
        n18276) );
  AOI22_X1 U21354 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n18276), .B1(
        n18498), .B2(n18351), .ZN(n18260) );
  OAI211_X1 U21355 ( .C1(n18501), .C2(n18302), .A(n18261), .B(n18260), .ZN(
        P3_U2916) );
  AOI22_X1 U21356 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18276), .B1(
        n18502), .B2(n18275), .ZN(n18263) );
  AOI22_X1 U21357 ( .A1(n18504), .A2(n18351), .B1(n18503), .B2(n18295), .ZN(
        n18262) );
  OAI211_X1 U21358 ( .C1(n18507), .C2(n18279), .A(n18263), .B(n18262), .ZN(
        P3_U2917) );
  AOI22_X1 U21359 ( .A1(n18436), .A2(n18270), .B1(n18508), .B2(n18275), .ZN(
        n18265) );
  AOI22_X1 U21360 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n18276), .B1(
        n18510), .B2(n18351), .ZN(n18264) );
  OAI211_X1 U21361 ( .C1(n18386), .C2(n18302), .A(n18265), .B(n18264), .ZN(
        P3_U2918) );
  AOI22_X1 U21362 ( .A1(n18515), .A2(n18295), .B1(n18514), .B2(n18275), .ZN(
        n18267) );
  AOI22_X1 U21363 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n18276), .B1(
        n18516), .B2(n18351), .ZN(n18266) );
  OAI211_X1 U21364 ( .C1(n18519), .C2(n18279), .A(n18267), .B(n18266), .ZN(
        P3_U2919) );
  AOI22_X1 U21365 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n18276), .B1(
        n18520), .B2(n18275), .ZN(n18269) );
  AOI22_X1 U21366 ( .A1(n18522), .A2(n18351), .B1(n18470), .B2(n18295), .ZN(
        n18268) );
  OAI211_X1 U21367 ( .C1(n18473), .C2(n18279), .A(n18269), .B(n18268), .ZN(
        P3_U2920) );
  AOI22_X1 U21368 ( .A1(n18526), .A2(n18275), .B1(n18474), .B2(n18270), .ZN(
        n18272) );
  AOI22_X1 U21369 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n18276), .B1(
        n18528), .B2(n18351), .ZN(n18271) );
  OAI211_X1 U21370 ( .C1(n18477), .C2(n18302), .A(n18272), .B(n18271), .ZN(
        P3_U2921) );
  AOI22_X1 U21371 ( .A1(n18478), .A2(n18295), .B1(n18532), .B2(n18275), .ZN(
        n18274) );
  AOI22_X1 U21372 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n18276), .B1(
        n18535), .B2(n18351), .ZN(n18273) );
  OAI211_X1 U21373 ( .C1(n18482), .C2(n18279), .A(n18274), .B(n18273), .ZN(
        P3_U2922) );
  AOI22_X1 U21374 ( .A1(n18542), .A2(n18295), .B1(n18541), .B2(n18275), .ZN(
        n18278) );
  AOI22_X1 U21375 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18276), .B1(
        n18544), .B2(n18351), .ZN(n18277) );
  OAI211_X1 U21376 ( .C1(n18550), .C2(n18279), .A(n18278), .B(n18277), .ZN(
        P3_U2923) );
  NAND2_X1 U21377 ( .A1(n18281), .A2(n18280), .ZN(n18299) );
  AOI22_X1 U21378 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n18299), .B1(
        n18492), .B2(n18298), .ZN(n18284) );
  NOR2_X2 U21379 ( .A1(n18593), .A2(n18282), .ZN(n18373) );
  AOI22_X1 U21380 ( .A1(n18431), .A2(n18322), .B1(n18498), .B2(n18373), .ZN(
        n18283) );
  OAI211_X1 U21381 ( .C1(n18381), .C2(n18302), .A(n18284), .B(n18283), .ZN(
        P3_U2924) );
  AOI22_X1 U21382 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18299), .B1(
        n18502), .B2(n18298), .ZN(n18286) );
  AOI22_X1 U21383 ( .A1(n18504), .A2(n18373), .B1(n18503), .B2(n18322), .ZN(
        n18285) );
  OAI211_X1 U21384 ( .C1(n18507), .C2(n18302), .A(n18286), .B(n18285), .ZN(
        P3_U2925) );
  INV_X1 U21385 ( .A(n18322), .ZN(n18320) );
  AOI22_X1 U21386 ( .A1(n18436), .A2(n18295), .B1(n18508), .B2(n18298), .ZN(
        n18288) );
  AOI22_X1 U21387 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n18299), .B1(
        n18510), .B2(n18373), .ZN(n18287) );
  OAI211_X1 U21388 ( .C1(n18386), .C2(n18320), .A(n18288), .B(n18287), .ZN(
        P3_U2926) );
  AOI22_X1 U21389 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n18299), .B1(
        n18514), .B2(n18298), .ZN(n18290) );
  AOI22_X1 U21390 ( .A1(n18516), .A2(n18373), .B1(n18515), .B2(n18322), .ZN(
        n18289) );
  OAI211_X1 U21391 ( .C1(n18519), .C2(n18302), .A(n18290), .B(n18289), .ZN(
        P3_U2927) );
  AOI22_X1 U21392 ( .A1(n18521), .A2(n18295), .B1(n18520), .B2(n18298), .ZN(
        n18292) );
  AOI22_X1 U21393 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n18299), .B1(
        n18522), .B2(n18373), .ZN(n18291) );
  OAI211_X1 U21394 ( .C1(n18525), .C2(n18320), .A(n18292), .B(n18291), .ZN(
        P3_U2928) );
  AOI22_X1 U21395 ( .A1(n18526), .A2(n18298), .B1(n18474), .B2(n18295), .ZN(
        n18294) );
  AOI22_X1 U21396 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n18299), .B1(
        n18528), .B2(n18373), .ZN(n18293) );
  OAI211_X1 U21397 ( .C1(n18477), .C2(n18320), .A(n18294), .B(n18293), .ZN(
        P3_U2929) );
  AOI22_X1 U21398 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n18299), .B1(
        n18532), .B2(n18298), .ZN(n18297) );
  AOI22_X1 U21399 ( .A1(n18535), .A2(n18373), .B1(n18534), .B2(n18295), .ZN(
        n18296) );
  OAI211_X1 U21400 ( .C1(n18538), .C2(n18320), .A(n18297), .B(n18296), .ZN(
        P3_U2930) );
  AOI22_X1 U21401 ( .A1(n18542), .A2(n18322), .B1(n18541), .B2(n18298), .ZN(
        n18301) );
  AOI22_X1 U21402 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n18299), .B1(
        n18544), .B2(n18373), .ZN(n18300) );
  OAI211_X1 U21403 ( .C1(n18550), .C2(n18302), .A(n18301), .B(n18300), .ZN(
        P3_U2931) );
  INV_X1 U21404 ( .A(n18351), .ZN(n18349) );
  NOR2_X2 U21405 ( .A1(n18595), .A2(n18378), .ZN(n18393) );
  NOR2_X1 U21406 ( .A1(n18373), .A2(n18393), .ZN(n18355) );
  NOR2_X1 U21407 ( .A1(n18623), .A2(n18355), .ZN(n18321) );
  AOI22_X1 U21408 ( .A1(n18493), .A2(n18322), .B1(n18492), .B2(n18321), .ZN(
        n18306) );
  OAI21_X1 U21409 ( .B1(n18303), .B2(n18456), .A(n18355), .ZN(n18304) );
  OAI211_X1 U21410 ( .C1(n18393), .C2(n18716), .A(n18458), .B(n18304), .ZN(
        n18323) );
  AOI22_X1 U21411 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n18323), .B1(
        n18498), .B2(n18393), .ZN(n18305) );
  OAI211_X1 U21412 ( .C1(n18501), .C2(n18349), .A(n18306), .B(n18305), .ZN(
        P3_U2932) );
  AOI22_X1 U21413 ( .A1(n18462), .A2(n18322), .B1(n18502), .B2(n18321), .ZN(
        n18308) );
  AOI22_X1 U21414 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18323), .B1(
        n18504), .B2(n18393), .ZN(n18307) );
  OAI211_X1 U21415 ( .C1(n18465), .C2(n18349), .A(n18308), .B(n18307), .ZN(
        P3_U2933) );
  AOI22_X1 U21416 ( .A1(n18436), .A2(n18322), .B1(n18508), .B2(n18321), .ZN(
        n18310) );
  AOI22_X1 U21417 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n18323), .B1(
        n18510), .B2(n18393), .ZN(n18309) );
  OAI211_X1 U21418 ( .C1(n18386), .C2(n18349), .A(n18310), .B(n18309), .ZN(
        P3_U2934) );
  AOI22_X1 U21419 ( .A1(n18440), .A2(n18322), .B1(n18514), .B2(n18321), .ZN(
        n18312) );
  AOI22_X1 U21420 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n18323), .B1(
        n18516), .B2(n18393), .ZN(n18311) );
  OAI211_X1 U21421 ( .C1(n18313), .C2(n18349), .A(n18312), .B(n18311), .ZN(
        P3_U2935) );
  AOI22_X1 U21422 ( .A1(n18521), .A2(n18322), .B1(n18520), .B2(n18321), .ZN(
        n18315) );
  AOI22_X1 U21423 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n18323), .B1(
        n18522), .B2(n18393), .ZN(n18314) );
  OAI211_X1 U21424 ( .C1(n18525), .C2(n18349), .A(n18315), .B(n18314), .ZN(
        P3_U2936) );
  AOI22_X1 U21425 ( .A1(n18527), .A2(n18351), .B1(n18526), .B2(n18321), .ZN(
        n18317) );
  AOI22_X1 U21426 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n18323), .B1(
        n18528), .B2(n18393), .ZN(n18316) );
  OAI211_X1 U21427 ( .C1(n18531), .C2(n18320), .A(n18317), .B(n18316), .ZN(
        P3_U2937) );
  AOI22_X1 U21428 ( .A1(n18478), .A2(n18351), .B1(n18532), .B2(n18321), .ZN(
        n18319) );
  AOI22_X1 U21429 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n18323), .B1(
        n18535), .B2(n18393), .ZN(n18318) );
  OAI211_X1 U21430 ( .C1(n18482), .C2(n18320), .A(n18319), .B(n18318), .ZN(
        P3_U2938) );
  AOI22_X1 U21431 ( .A1(n18485), .A2(n18322), .B1(n18541), .B2(n18321), .ZN(
        n18325) );
  AOI22_X1 U21432 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18323), .B1(
        n18544), .B2(n18393), .ZN(n18324) );
  OAI211_X1 U21433 ( .C1(n18490), .C2(n18349), .A(n18325), .B(n18324), .ZN(
        P3_U2939) );
  OR2_X1 U21434 ( .A1(n18326), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n18329) );
  NAND2_X1 U21435 ( .A1(n18377), .A2(n18594), .ZN(n18327) );
  OAI22_X1 U21436 ( .A1(n18428), .A2(n18329), .B1(n18328), .B2(n18327), .ZN(
        n18341) );
  NOR2_X1 U21437 ( .A1(n18378), .A2(n18429), .ZN(n18350) );
  AOI22_X1 U21438 ( .A1(n18431), .A2(n18373), .B1(n18492), .B2(n18350), .ZN(
        n18332) );
  NOR2_X2 U21439 ( .A1(n18378), .A2(n18330), .ZN(n18416) );
  AOI22_X1 U21440 ( .A1(n18498), .A2(n18416), .B1(n18493), .B2(n18351), .ZN(
        n18331) );
  OAI211_X1 U21441 ( .C1(n18333), .C2(n18341), .A(n18332), .B(n18331), .ZN(
        P3_U2940) );
  AOI22_X1 U21442 ( .A1(n18502), .A2(n18350), .B1(n18503), .B2(n18373), .ZN(
        n18335) );
  AOI22_X1 U21443 ( .A1(n18462), .A2(n18351), .B1(n18504), .B2(n18416), .ZN(
        n18334) );
  OAI211_X1 U21444 ( .C1(n18336), .C2(n18341), .A(n18335), .B(n18334), .ZN(
        P3_U2941) );
  AOI22_X1 U21445 ( .A1(n18509), .A2(n18373), .B1(n18508), .B2(n18350), .ZN(
        n18338) );
  INV_X1 U21446 ( .A(n18341), .ZN(n18352) );
  AOI22_X1 U21447 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n18352), .B1(
        n18510), .B2(n18416), .ZN(n18337) );
  OAI211_X1 U21448 ( .C1(n18513), .C2(n18349), .A(n18338), .B(n18337), .ZN(
        P3_U2942) );
  AOI22_X1 U21449 ( .A1(n18515), .A2(n18373), .B1(n18514), .B2(n18350), .ZN(
        n18340) );
  AOI22_X1 U21450 ( .A1(n18440), .A2(n18351), .B1(n18516), .B2(n18416), .ZN(
        n18339) );
  OAI211_X1 U21451 ( .C1(n18342), .C2(n18341), .A(n18340), .B(n18339), .ZN(
        P3_U2943) );
  AOI22_X1 U21452 ( .A1(n18470), .A2(n18373), .B1(n18520), .B2(n18350), .ZN(
        n18344) );
  AOI22_X1 U21453 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n18352), .B1(
        n18522), .B2(n18416), .ZN(n18343) );
  OAI211_X1 U21454 ( .C1(n18473), .C2(n18349), .A(n18344), .B(n18343), .ZN(
        P3_U2944) );
  AOI22_X1 U21455 ( .A1(n18527), .A2(n18373), .B1(n18526), .B2(n18350), .ZN(
        n18346) );
  AOI22_X1 U21456 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n18352), .B1(
        n18528), .B2(n18416), .ZN(n18345) );
  OAI211_X1 U21457 ( .C1(n18531), .C2(n18349), .A(n18346), .B(n18345), .ZN(
        P3_U2945) );
  AOI22_X1 U21458 ( .A1(n18478), .A2(n18373), .B1(n18532), .B2(n18350), .ZN(
        n18348) );
  AOI22_X1 U21459 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n18352), .B1(
        n18535), .B2(n18416), .ZN(n18347) );
  OAI211_X1 U21460 ( .C1(n18482), .C2(n18349), .A(n18348), .B(n18347), .ZN(
        P3_U2946) );
  INV_X1 U21461 ( .A(n18373), .ZN(n18371) );
  AOI22_X1 U21462 ( .A1(n18485), .A2(n18351), .B1(n18541), .B2(n18350), .ZN(
        n18354) );
  AOI22_X1 U21463 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n18352), .B1(
        n18544), .B2(n18416), .ZN(n18353) );
  OAI211_X1 U21464 ( .C1(n18490), .C2(n18371), .A(n18354), .B(n18353), .ZN(
        P3_U2947) );
  NAND2_X1 U21465 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18377), .ZN(
        n18427) );
  NOR2_X1 U21466 ( .A1(n18416), .A2(n9770), .ZN(n18402) );
  OAI21_X1 U21467 ( .B1(n18355), .B2(n18456), .A(n18402), .ZN(n18356) );
  OAI211_X1 U21468 ( .C1(n9770), .C2(n18716), .A(n18458), .B(n18356), .ZN(
        n18374) );
  NOR2_X1 U21469 ( .A1(n18623), .A2(n18402), .ZN(n18372) );
  AOI22_X1 U21470 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n18374), .B1(
        n18492), .B2(n18372), .ZN(n18358) );
  AOI22_X1 U21471 ( .A1(n18431), .A2(n18393), .B1(n18498), .B2(n9770), .ZN(
        n18357) );
  OAI211_X1 U21472 ( .C1(n18381), .C2(n18371), .A(n18358), .B(n18357), .ZN(
        P3_U2948) );
  INV_X1 U21473 ( .A(n18393), .ZN(n18400) );
  AOI22_X1 U21474 ( .A1(n18462), .A2(n18373), .B1(n18502), .B2(n18372), .ZN(
        n18360) );
  AOI22_X1 U21475 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n18374), .B1(
        n18504), .B2(n9770), .ZN(n18359) );
  OAI211_X1 U21476 ( .C1(n18465), .C2(n18400), .A(n18360), .B(n18359), .ZN(
        P3_U2949) );
  AOI22_X1 U21477 ( .A1(n18509), .A2(n18393), .B1(n18508), .B2(n18372), .ZN(
        n18362) );
  AOI22_X1 U21478 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n18374), .B1(
        n18510), .B2(n9770), .ZN(n18361) );
  OAI211_X1 U21479 ( .C1(n18513), .C2(n18371), .A(n18362), .B(n18361), .ZN(
        P3_U2950) );
  AOI22_X1 U21480 ( .A1(n18515), .A2(n18393), .B1(n18514), .B2(n18372), .ZN(
        n18364) );
  AOI22_X1 U21481 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n18374), .B1(
        n18516), .B2(n9770), .ZN(n18363) );
  OAI211_X1 U21482 ( .C1(n18519), .C2(n18371), .A(n18364), .B(n18363), .ZN(
        P3_U2951) );
  AOI22_X1 U21483 ( .A1(n18521), .A2(n18373), .B1(n18520), .B2(n18372), .ZN(
        n18366) );
  AOI22_X1 U21484 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n18374), .B1(
        n18522), .B2(n9770), .ZN(n18365) );
  OAI211_X1 U21485 ( .C1(n18525), .C2(n18400), .A(n18366), .B(n18365), .ZN(
        P3_U2952) );
  AOI22_X1 U21486 ( .A1(n18527), .A2(n18393), .B1(n18526), .B2(n18372), .ZN(
        n18368) );
  AOI22_X1 U21487 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n18374), .B1(
        n18528), .B2(n9770), .ZN(n18367) );
  OAI211_X1 U21488 ( .C1(n18531), .C2(n18371), .A(n18368), .B(n18367), .ZN(
        P3_U2953) );
  AOI22_X1 U21489 ( .A1(n18478), .A2(n18393), .B1(n18532), .B2(n18372), .ZN(
        n18370) );
  AOI22_X1 U21490 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n18374), .B1(
        n18535), .B2(n9770), .ZN(n18369) );
  OAI211_X1 U21491 ( .C1(n18482), .C2(n18371), .A(n18370), .B(n18369), .ZN(
        P3_U2954) );
  AOI22_X1 U21492 ( .A1(n18485), .A2(n18373), .B1(n18541), .B2(n18372), .ZN(
        n18376) );
  AOI22_X1 U21493 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n18374), .B1(
        n18544), .B2(n9770), .ZN(n18375) );
  OAI211_X1 U21494 ( .C1(n18490), .C2(n18400), .A(n18376), .B(n18375), .ZN(
        P3_U2955) );
  NOR2_X1 U21495 ( .A1(n18623), .A2(n18427), .ZN(n18396) );
  AOI22_X1 U21496 ( .A1(n18431), .A2(n18416), .B1(n18492), .B2(n18396), .ZN(
        n18380) );
  OAI211_X1 U21497 ( .C1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(n18497), .A(
        n18494), .B(n18377), .ZN(n18397) );
  NOR2_X2 U21498 ( .A1(n18593), .A2(n18378), .ZN(n18484) );
  AOI22_X1 U21499 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n18397), .B1(
        n18498), .B2(n18484), .ZN(n18379) );
  OAI211_X1 U21500 ( .C1(n18381), .C2(n18400), .A(n18380), .B(n18379), .ZN(
        P3_U2956) );
  INV_X1 U21501 ( .A(n18416), .ZN(n18424) );
  AOI22_X1 U21502 ( .A1(n18462), .A2(n18393), .B1(n18502), .B2(n18396), .ZN(
        n18383) );
  AOI22_X1 U21503 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n18397), .B1(
        n18504), .B2(n18484), .ZN(n18382) );
  OAI211_X1 U21504 ( .C1(n18465), .C2(n18424), .A(n18383), .B(n18382), .ZN(
        P3_U2957) );
  AOI22_X1 U21505 ( .A1(n18436), .A2(n18393), .B1(n18508), .B2(n18396), .ZN(
        n18385) );
  AOI22_X1 U21506 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n18397), .B1(
        n18510), .B2(n18484), .ZN(n18384) );
  OAI211_X1 U21507 ( .C1(n18386), .C2(n18424), .A(n18385), .B(n18384), .ZN(
        P3_U2958) );
  AOI22_X1 U21508 ( .A1(n18515), .A2(n18416), .B1(n18514), .B2(n18396), .ZN(
        n18388) );
  AOI22_X1 U21509 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n18397), .B1(
        n18516), .B2(n18484), .ZN(n18387) );
  OAI211_X1 U21510 ( .C1(n18519), .C2(n18400), .A(n18388), .B(n18387), .ZN(
        P3_U2959) );
  AOI22_X1 U21511 ( .A1(n18470), .A2(n18416), .B1(n18520), .B2(n18396), .ZN(
        n18390) );
  AOI22_X1 U21512 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n18397), .B1(
        n18522), .B2(n18484), .ZN(n18389) );
  OAI211_X1 U21513 ( .C1(n18473), .C2(n18400), .A(n18390), .B(n18389), .ZN(
        P3_U2960) );
  AOI22_X1 U21514 ( .A1(n18526), .A2(n18396), .B1(n18474), .B2(n18393), .ZN(
        n18392) );
  AOI22_X1 U21515 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n18397), .B1(
        n18528), .B2(n18484), .ZN(n18391) );
  OAI211_X1 U21516 ( .C1(n18477), .C2(n18424), .A(n18392), .B(n18391), .ZN(
        P3_U2961) );
  AOI22_X1 U21517 ( .A1(n18534), .A2(n18393), .B1(n18532), .B2(n18396), .ZN(
        n18395) );
  AOI22_X1 U21518 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n18397), .B1(
        n18535), .B2(n18484), .ZN(n18394) );
  OAI211_X1 U21519 ( .C1(n18538), .C2(n18424), .A(n18395), .B(n18394), .ZN(
        P3_U2962) );
  AOI22_X1 U21520 ( .A1(n18542), .A2(n18416), .B1(n18541), .B2(n18396), .ZN(
        n18399) );
  AOI22_X1 U21521 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n18397), .B1(
        n18544), .B2(n18484), .ZN(n18398) );
  OAI211_X1 U21522 ( .C1(n18550), .C2(n18400), .A(n18399), .B(n18398), .ZN(
        P3_U2963) );
  INV_X1 U21523 ( .A(n9770), .ZN(n18419) );
  NOR2_X2 U21524 ( .A1(n18595), .A2(n18430), .ZN(n18533) );
  NOR2_X1 U21525 ( .A1(n18484), .A2(n18533), .ZN(n18457) );
  NOR2_X1 U21526 ( .A1(n18623), .A2(n18457), .ZN(n18420) );
  AOI22_X1 U21527 ( .A1(n18493), .A2(n18416), .B1(n18492), .B2(n18420), .ZN(
        n18405) );
  OAI22_X1 U21528 ( .A1(n18402), .A2(n18428), .B1(n18457), .B2(n18401), .ZN(
        n18403) );
  OAI21_X1 U21529 ( .B1(n18533), .B2(n18716), .A(n18403), .ZN(n18421) );
  AOI22_X1 U21530 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n18421), .B1(
        n18498), .B2(n18533), .ZN(n18404) );
  OAI211_X1 U21531 ( .C1(n18501), .C2(n18419), .A(n18405), .B(n18404), .ZN(
        P3_U2964) );
  AOI22_X1 U21532 ( .A1(n18462), .A2(n18416), .B1(n18502), .B2(n18420), .ZN(
        n18407) );
  AOI22_X1 U21533 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18421), .B1(
        n18504), .B2(n18533), .ZN(n18406) );
  OAI211_X1 U21534 ( .C1(n18465), .C2(n18419), .A(n18407), .B(n18406), .ZN(
        P3_U2965) );
  AOI22_X1 U21535 ( .A1(n18509), .A2(n9770), .B1(n18508), .B2(n18420), .ZN(
        n18409) );
  AOI22_X1 U21536 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n18421), .B1(
        n18510), .B2(n18533), .ZN(n18408) );
  OAI211_X1 U21537 ( .C1(n18513), .C2(n18424), .A(n18409), .B(n18408), .ZN(
        P3_U2966) );
  AOI22_X1 U21538 ( .A1(n18515), .A2(n9770), .B1(n18514), .B2(n18420), .ZN(
        n18411) );
  AOI22_X1 U21539 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n18421), .B1(
        n18516), .B2(n18533), .ZN(n18410) );
  OAI211_X1 U21540 ( .C1(n18519), .C2(n18424), .A(n18411), .B(n18410), .ZN(
        P3_U2967) );
  AOI22_X1 U21541 ( .A1(n18521), .A2(n18416), .B1(n18520), .B2(n18420), .ZN(
        n18413) );
  AOI22_X1 U21542 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n18421), .B1(
        n18522), .B2(n18533), .ZN(n18412) );
  OAI211_X1 U21543 ( .C1(n18525), .C2(n18419), .A(n18413), .B(n18412), .ZN(
        P3_U2968) );
  AOI22_X1 U21544 ( .A1(n18526), .A2(n18420), .B1(n18474), .B2(n18416), .ZN(
        n18415) );
  AOI22_X1 U21545 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n18421), .B1(
        n18528), .B2(n18533), .ZN(n18414) );
  OAI211_X1 U21546 ( .C1(n18477), .C2(n18419), .A(n18415), .B(n18414), .ZN(
        P3_U2969) );
  AOI22_X1 U21547 ( .A1(n18534), .A2(n18416), .B1(n18532), .B2(n18420), .ZN(
        n18418) );
  AOI22_X1 U21548 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18421), .B1(
        n18535), .B2(n18533), .ZN(n18417) );
  OAI211_X1 U21549 ( .C1(n18538), .C2(n18419), .A(n18418), .B(n18417), .ZN(
        P3_U2970) );
  AOI22_X1 U21550 ( .A1(n18542), .A2(n9770), .B1(n18541), .B2(n18420), .ZN(
        n18423) );
  AOI22_X1 U21551 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n18421), .B1(
        n18544), .B2(n18533), .ZN(n18422) );
  OAI211_X1 U21552 ( .C1(n18550), .C2(n18424), .A(n18423), .B(n18422), .ZN(
        P3_U2971) );
  INV_X1 U21553 ( .A(n18425), .ZN(n18426) );
  OAI22_X1 U21554 ( .A1(n18428), .A2(n18427), .B1(n18430), .B2(n18426), .ZN(
        n18446) );
  NOR2_X1 U21555 ( .A1(n18430), .A2(n18429), .ZN(n18496) );
  AOI22_X1 U21556 ( .A1(n18493), .A2(n9770), .B1(n18492), .B2(n18496), .ZN(
        n18433) );
  AOI22_X1 U21557 ( .A1(n18543), .A2(n18498), .B1(n18431), .B2(n18484), .ZN(
        n18432) );
  OAI211_X1 U21558 ( .C1(n21054), .C2(n18446), .A(n18433), .B(n18432), .ZN(
        P3_U2972) );
  AOI22_X1 U21559 ( .A1(n18462), .A2(n9770), .B1(n18502), .B2(n18496), .ZN(
        n18435) );
  AOI22_X1 U21560 ( .A1(n18543), .A2(n18504), .B1(n18503), .B2(n18484), .ZN(
        n18434) );
  OAI211_X1 U21561 ( .C1(n20927), .C2(n18446), .A(n18435), .B(n18434), .ZN(
        P3_U2973) );
  AOI22_X1 U21562 ( .A1(n18436), .A2(n9770), .B1(n18508), .B2(n18496), .ZN(
        n18438) );
  AOI22_X1 U21563 ( .A1(n18543), .A2(n18510), .B1(n18509), .B2(n18484), .ZN(
        n18437) );
  OAI211_X1 U21564 ( .C1(n18439), .C2(n18446), .A(n18438), .B(n18437), .ZN(
        P3_U2974) );
  AOI22_X1 U21565 ( .A1(n18440), .A2(n9770), .B1(n18514), .B2(n18496), .ZN(
        n18442) );
  AOI22_X1 U21566 ( .A1(n18543), .A2(n18516), .B1(n18515), .B2(n18484), .ZN(
        n18441) );
  OAI211_X1 U21567 ( .C1(n18443), .C2(n18446), .A(n18442), .B(n18441), .ZN(
        P3_U2975) );
  AOI22_X1 U21568 ( .A1(n18470), .A2(n18484), .B1(n18520), .B2(n18496), .ZN(
        n18445) );
  AOI22_X1 U21569 ( .A1(n18543), .A2(n18522), .B1(n18521), .B2(n9770), .ZN(
        n18444) );
  OAI211_X1 U21570 ( .C1(n20935), .C2(n18446), .A(n18445), .B(n18444), .ZN(
        P3_U2976) );
  INV_X1 U21571 ( .A(n18484), .ZN(n18481) );
  AOI22_X1 U21572 ( .A1(n18526), .A2(n18496), .B1(n18474), .B2(n9770), .ZN(
        n18448) );
  INV_X1 U21573 ( .A(n18446), .ZN(n18452) );
  AOI22_X1 U21574 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n18452), .B1(
        n18543), .B2(n18528), .ZN(n18447) );
  OAI211_X1 U21575 ( .C1(n18477), .C2(n18481), .A(n18448), .B(n18447), .ZN(
        P3_U2977) );
  AOI22_X1 U21576 ( .A1(n18534), .A2(n9770), .B1(n18532), .B2(n18496), .ZN(
        n18451) );
  AOI22_X1 U21577 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n18452), .B1(
        n18543), .B2(n18535), .ZN(n18450) );
  OAI211_X1 U21578 ( .C1(n18538), .C2(n18481), .A(n18451), .B(n18450), .ZN(
        P3_U2978) );
  AOI22_X1 U21579 ( .A1(n18485), .A2(n9770), .B1(n18541), .B2(n18496), .ZN(
        n18454) );
  AOI22_X1 U21580 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n18452), .B1(
        n18543), .B2(n18544), .ZN(n18453) );
  OAI211_X1 U21581 ( .C1(n18490), .C2(n18481), .A(n18454), .B(n18453), .ZN(
        P3_U2979) );
  INV_X1 U21582 ( .A(n18533), .ZN(n18549) );
  AND2_X1 U21583 ( .A1(n18491), .A2(n18455), .ZN(n18483) );
  AOI22_X1 U21584 ( .A1(n18493), .A2(n18484), .B1(n18492), .B2(n18483), .ZN(
        n18461) );
  AOI221_X1 U21585 ( .B1(n18457), .B2(n18539), .C1(n18456), .C2(n18539), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18459) );
  OAI21_X1 U21586 ( .B1(n18486), .B2(n18459), .A(n18458), .ZN(n18487) );
  AOI22_X1 U21587 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n18487), .B1(
        n18486), .B2(n18498), .ZN(n18460) );
  OAI211_X1 U21588 ( .C1(n18501), .C2(n18549), .A(n18461), .B(n18460), .ZN(
        P3_U2980) );
  AOI22_X1 U21589 ( .A1(n18462), .A2(n18484), .B1(n18502), .B2(n18483), .ZN(
        n18464) );
  AOI22_X1 U21590 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18487), .B1(
        n18486), .B2(n18504), .ZN(n18463) );
  OAI211_X1 U21591 ( .C1(n18465), .C2(n18549), .A(n18464), .B(n18463), .ZN(
        P3_U2981) );
  AOI22_X1 U21592 ( .A1(n18509), .A2(n18533), .B1(n18508), .B2(n18483), .ZN(
        n18467) );
  AOI22_X1 U21593 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n18487), .B1(
        n18486), .B2(n18510), .ZN(n18466) );
  OAI211_X1 U21594 ( .C1(n18513), .C2(n18481), .A(n18467), .B(n18466), .ZN(
        P3_U2982) );
  AOI22_X1 U21595 ( .A1(n18515), .A2(n18533), .B1(n18514), .B2(n18483), .ZN(
        n18469) );
  AOI22_X1 U21596 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n18487), .B1(
        n18486), .B2(n18516), .ZN(n18468) );
  OAI211_X1 U21597 ( .C1(n18519), .C2(n18481), .A(n18469), .B(n18468), .ZN(
        P3_U2983) );
  AOI22_X1 U21598 ( .A1(n18470), .A2(n18533), .B1(n18520), .B2(n18483), .ZN(
        n18472) );
  AOI22_X1 U21599 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n18487), .B1(
        n18486), .B2(n18522), .ZN(n18471) );
  OAI211_X1 U21600 ( .C1(n18473), .C2(n18481), .A(n18472), .B(n18471), .ZN(
        P3_U2984) );
  AOI22_X1 U21601 ( .A1(n18526), .A2(n18483), .B1(n18474), .B2(n18484), .ZN(
        n18476) );
  AOI22_X1 U21602 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n18487), .B1(
        n18486), .B2(n18528), .ZN(n18475) );
  OAI211_X1 U21603 ( .C1(n18477), .C2(n18549), .A(n18476), .B(n18475), .ZN(
        P3_U2985) );
  AOI22_X1 U21604 ( .A1(n18478), .A2(n18533), .B1(n18532), .B2(n18483), .ZN(
        n18480) );
  AOI22_X1 U21605 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n18487), .B1(
        n18486), .B2(n18535), .ZN(n18479) );
  OAI211_X1 U21606 ( .C1(n18482), .C2(n18481), .A(n18480), .B(n18479), .ZN(
        P3_U2986) );
  AOI22_X1 U21607 ( .A1(n18485), .A2(n18484), .B1(n18541), .B2(n18483), .ZN(
        n18489) );
  AOI22_X1 U21608 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n18487), .B1(
        n18486), .B2(n18544), .ZN(n18488) );
  OAI211_X1 U21609 ( .C1(n18490), .C2(n18549), .A(n18489), .B(n18488), .ZN(
        P3_U2987) );
  AND2_X1 U21610 ( .A1(n18491), .A2(n18495), .ZN(n18540) );
  AOI22_X1 U21611 ( .A1(n18493), .A2(n18533), .B1(n18492), .B2(n18540), .ZN(
        n18500) );
  AOI22_X1 U21612 ( .A1(n18497), .A2(n18496), .B1(n18495), .B2(n18494), .ZN(
        n18546) );
  AOI22_X1 U21613 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n18546), .B1(
        n18545), .B2(n18498), .ZN(n18499) );
  OAI211_X1 U21614 ( .C1(n18539), .C2(n18501), .A(n18500), .B(n18499), .ZN(
        P3_U2988) );
  AOI22_X1 U21615 ( .A1(n18543), .A2(n18503), .B1(n18502), .B2(n18540), .ZN(
        n18506) );
  AOI22_X1 U21616 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n18546), .B1(
        n18545), .B2(n18504), .ZN(n18505) );
  OAI211_X1 U21617 ( .C1(n18507), .C2(n18549), .A(n18506), .B(n18505), .ZN(
        P3_U2989) );
  AOI22_X1 U21618 ( .A1(n18543), .A2(n18509), .B1(n18508), .B2(n18540), .ZN(
        n18512) );
  AOI22_X1 U21619 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n18546), .B1(
        n18545), .B2(n18510), .ZN(n18511) );
  OAI211_X1 U21620 ( .C1(n18513), .C2(n18549), .A(n18512), .B(n18511), .ZN(
        P3_U2990) );
  AOI22_X1 U21621 ( .A1(n18543), .A2(n18515), .B1(n18514), .B2(n18540), .ZN(
        n18518) );
  AOI22_X1 U21622 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n18546), .B1(
        n18545), .B2(n18516), .ZN(n18517) );
  OAI211_X1 U21623 ( .C1(n18519), .C2(n18549), .A(n18518), .B(n18517), .ZN(
        P3_U2991) );
  AOI22_X1 U21624 ( .A1(n18521), .A2(n18533), .B1(n18520), .B2(n18540), .ZN(
        n18524) );
  AOI22_X1 U21625 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n18546), .B1(
        n18545), .B2(n18522), .ZN(n18523) );
  OAI211_X1 U21626 ( .C1(n18539), .C2(n18525), .A(n18524), .B(n18523), .ZN(
        P3_U2992) );
  AOI22_X1 U21627 ( .A1(n18543), .A2(n18527), .B1(n18526), .B2(n18540), .ZN(
        n18530) );
  AOI22_X1 U21628 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n18546), .B1(
        n18545), .B2(n18528), .ZN(n18529) );
  OAI211_X1 U21629 ( .C1(n18531), .C2(n18549), .A(n18530), .B(n18529), .ZN(
        P3_U2993) );
  AOI22_X1 U21630 ( .A1(n18534), .A2(n18533), .B1(n18532), .B2(n18540), .ZN(
        n18537) );
  AOI22_X1 U21631 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n18546), .B1(
        n18545), .B2(n18535), .ZN(n18536) );
  OAI211_X1 U21632 ( .C1(n18539), .C2(n18538), .A(n18537), .B(n18536), .ZN(
        P3_U2994) );
  AOI22_X1 U21633 ( .A1(n18543), .A2(n18542), .B1(n18541), .B2(n18540), .ZN(
        n18548) );
  AOI22_X1 U21634 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n18546), .B1(
        n18545), .B2(n18544), .ZN(n18547) );
  OAI211_X1 U21635 ( .C1(n18550), .C2(n18549), .A(n18548), .B(n18547), .ZN(
        P3_U2995) );
  NOR2_X1 U21636 ( .A1(n18567), .A2(n18551), .ZN(n18553) );
  OAI222_X1 U21637 ( .A1(n18557), .A2(n18556), .B1(n18555), .B2(n18554), .C1(
        n18553), .C2(n18552), .ZN(n18757) );
  OAI21_X1 U21638 ( .B1(P3_MORE_REG_SCAN_IN), .B2(P3_FLUSH_REG_SCAN_IN), .A(
        n18558), .ZN(n18559) );
  OAI211_X1 U21639 ( .C1(n18561), .C2(n18586), .A(n18560), .B(n18559), .ZN(
        n18607) );
  NAND2_X1 U21640 ( .A1(n18576), .A2(n18732), .ZN(n18566) );
  OAI21_X1 U21641 ( .B1(n18745), .B2(n18563), .A(n18562), .ZN(n18579) );
  NOR2_X1 U21642 ( .A1(n18579), .A2(n18564), .ZN(n18590) );
  INV_X1 U21643 ( .A(n18590), .ZN(n18565) );
  AOI22_X1 U21644 ( .A1(n18567), .A2(n18566), .B1(n18573), .B2(n18565), .ZN(
        n18568) );
  NOR2_X1 U21645 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18568), .ZN(
        n18719) );
  AOI21_X1 U21646 ( .B1(n18571), .B2(n18570), .A(n18569), .ZN(n18577) );
  OAI22_X1 U21647 ( .A1(n18589), .A2(n18573), .B1(n18572), .B2(n18577), .ZN(
        n18574) );
  AOI21_X1 U21648 ( .B1(n18576), .B2(n18732), .A(n18574), .ZN(n18720) );
  NAND2_X1 U21649 ( .A1(n18586), .A2(n18720), .ZN(n18575) );
  AOI22_X1 U21650 ( .A1(n18586), .A2(n18719), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n18575), .ZN(n18605) );
  INV_X1 U21651 ( .A(n18586), .ZN(n18597) );
  AND2_X1 U21652 ( .A1(n18576), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n18585) );
  INV_X1 U21653 ( .A(n18577), .ZN(n18584) );
  NAND2_X1 U21654 ( .A1(n18739), .A2(n18732), .ZN(n18578) );
  OAI221_X1 U21655 ( .B1(n18739), .B2(n18732), .C1(n18580), .C2(n18579), .A(
        n18578), .ZN(n18581) );
  OAI21_X1 U21656 ( .B1(n18729), .B2(n18582), .A(n18581), .ZN(n18583) );
  AOI21_X1 U21657 ( .B1(n18585), .B2(n18584), .A(n18583), .ZN(n18725) );
  AOI22_X1 U21658 ( .A1(n18597), .A2(n18732), .B1(n18725), .B2(n18586), .ZN(
        n18601) );
  NOR2_X1 U21659 ( .A1(n18588), .A2(n18587), .ZN(n18592) );
  AOI22_X1 U21660 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18589), .B1(
        n18592), .B2(n18745), .ZN(n18741) );
  OAI22_X1 U21661 ( .A1(n18592), .A2(n18591), .B1(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18590), .ZN(n18737) );
  AOI222_X1 U21662 ( .A1(n18741), .A2(n18737), .B1(n18741), .B2(n18594), .C1(
        n18737), .C2(n18593), .ZN(n18596) );
  OAI21_X1 U21663 ( .B1(n18597), .B2(n18596), .A(n18595), .ZN(n18600) );
  AND2_X1 U21664 ( .A1(n18601), .A2(n18600), .ZN(n18598) );
  OAI221_X1 U21665 ( .B1(n18601), .B2(n18600), .C1(n18599), .C2(n18598), .A(
        n20878), .ZN(n18604) );
  AOI21_X1 U21666 ( .B1(n20878), .B2(n18602), .A(n18601), .ZN(n18603) );
  AOI222_X1 U21667 ( .A1(n18605), .A2(n18604), .B1(n18605), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C1(n18604), .C2(n18603), .ZN(
        n18606) );
  NOR4_X1 U21668 ( .A1(n18608), .A2(n18757), .A3(n18607), .A4(n18606), .ZN(
        n18620) );
  AOI22_X1 U21669 ( .A1(n18740), .A2(n18609), .B1(n18761), .B2(n18769), .ZN(
        n18610) );
  INV_X1 U21670 ( .A(n18610), .ZN(n18616) );
  OAI211_X1 U21671 ( .C1(n18613), .C2(n18612), .A(n18611), .B(n18620), .ZN(
        n18715) );
  OAI21_X1 U21672 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(n18768), .A(n18715), 
        .ZN(n18622) );
  NOR2_X1 U21673 ( .A1(n18614), .A2(n18622), .ZN(n18615) );
  MUX2_X1 U21674 ( .A(n18616), .B(n18615), .S(P3_STATE2_REG_0__SCAN_IN), .Z(
        n18618) );
  OAI211_X1 U21675 ( .C1(n18620), .C2(n18619), .A(n18618), .B(n18617), .ZN(
        P3_U2996) );
  OAI221_X1 U21676 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n18621), .C1(n18764), 
        .C2(n18761), .A(n18775), .ZN(n18626) );
  NAND2_X1 U21677 ( .A1(n18761), .A2(n18769), .ZN(n18624) );
  OAI211_X1 U21678 ( .C1(n18626), .C2(n18726), .A(n18625), .B(n18624), .ZN(
        P3_U2997) );
  AND3_X1 U21679 ( .A1(n18626), .A2(n18763), .A3(n18714), .ZN(P3_U2998) );
  AND2_X1 U21680 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n18627), .ZN(
        P3_U2999) );
  AND2_X1 U21681 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n18627), .ZN(
        P3_U3000) );
  AND2_X1 U21682 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n18627), .ZN(
        P3_U3001) );
  AND2_X1 U21683 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n18627), .ZN(
        P3_U3002) );
  AND2_X1 U21684 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n18627), .ZN(
        P3_U3003) );
  AND2_X1 U21685 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n18627), .ZN(
        P3_U3004) );
  AND2_X1 U21686 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n18627), .ZN(
        P3_U3005) );
  AND2_X1 U21687 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n18627), .ZN(
        P3_U3006) );
  AND2_X1 U21688 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n18627), .ZN(
        P3_U3007) );
  AND2_X1 U21689 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n18627), .ZN(
        P3_U3008) );
  AND2_X1 U21690 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n18627), .ZN(
        P3_U3009) );
  AND2_X1 U21691 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n18627), .ZN(
        P3_U3010) );
  AND2_X1 U21692 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n18627), .ZN(
        P3_U3011) );
  AND2_X1 U21693 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n18627), .ZN(
        P3_U3012) );
  AND2_X1 U21694 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n18627), .ZN(
        P3_U3013) );
  AND2_X1 U21695 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n18627), .ZN(
        P3_U3014) );
  AND2_X1 U21696 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n18627), .ZN(
        P3_U3015) );
  AND2_X1 U21697 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n18627), .ZN(
        P3_U3016) );
  AND2_X1 U21698 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n18627), .ZN(
        P3_U3017) );
  AND2_X1 U21699 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n18627), .ZN(
        P3_U3018) );
  AND2_X1 U21700 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n18627), .ZN(
        P3_U3019) );
  AND2_X1 U21701 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n18627), .ZN(
        P3_U3020) );
  AND2_X1 U21702 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n18627), .ZN(P3_U3021) );
  AND2_X1 U21703 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n18627), .ZN(P3_U3022) );
  AND2_X1 U21704 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n18627), .ZN(P3_U3023) );
  AND2_X1 U21705 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n18627), .ZN(P3_U3024) );
  AND2_X1 U21706 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n18627), .ZN(P3_U3025) );
  AND2_X1 U21707 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n18627), .ZN(P3_U3026) );
  AND2_X1 U21708 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n18627), .ZN(P3_U3027) );
  AND2_X1 U21709 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n18627), .ZN(P3_U3028) );
  OAI21_X1 U21710 ( .B1(n20703), .B2(n18628), .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18629) );
  INV_X1 U21711 ( .A(n18629), .ZN(n18632) );
  NAND2_X1 U21712 ( .A1(n18761), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n18638) );
  INV_X1 U21713 ( .A(n18638), .ZN(n18634) );
  NOR2_X1 U21714 ( .A1(n18634), .A2(n18642), .ZN(n18644) );
  INV_X1 U21715 ( .A(NA), .ZN(n20690) );
  OAI21_X1 U21716 ( .B1(n20690), .B2(n18630), .A(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n18643) );
  INV_X1 U21717 ( .A(n18643), .ZN(n18631) );
  OAI22_X1 U21718 ( .A1(n18772), .A2(n18632), .B1(n18644), .B2(n18631), .ZN(
        P3_U3029) );
  NOR2_X1 U21719 ( .A1(n18645), .A2(n20703), .ZN(n18640) );
  INV_X1 U21720 ( .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18633) );
  NOR3_X1 U21721 ( .A1(n18640), .A2(n18633), .A3(n18642), .ZN(n18635) );
  NOR2_X1 U21722 ( .A1(n18635), .A2(n18634), .ZN(n18636) );
  OAI211_X1 U21723 ( .C1(n20703), .C2(n18637), .A(n18636), .B(n18758), .ZN(
        P3_U3030) );
  OAI22_X1 U21724 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(NA), .B2(n18638), .ZN(n18639) );
  OAI22_X1 U21725 ( .A1(n18640), .A2(n18639), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n18641) );
  OAI22_X1 U21726 ( .A1(n18644), .A2(n18643), .B1(n18642), .B2(n18641), .ZN(
        P3_U3031) );
  INV_X1 U21727 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n18647) );
  OAI222_X1 U21728 ( .A1(n18749), .A2(n18707), .B1(n18646), .B2(n18772), .C1(
        n18647), .C2(n18703), .ZN(P3_U3032) );
  OAI222_X1 U21729 ( .A1(n18703), .A2(n18649), .B1(n18648), .B2(n18772), .C1(
        n18647), .C2(n18707), .ZN(P3_U3033) );
  OAI222_X1 U21730 ( .A1(n18703), .A2(n18651), .B1(n18650), .B2(n18772), .C1(
        n18649), .C2(n18707), .ZN(P3_U3034) );
  INV_X1 U21731 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n18653) );
  OAI222_X1 U21732 ( .A1(n18703), .A2(n18653), .B1(n18652), .B2(n18772), .C1(
        n18651), .C2(n18707), .ZN(P3_U3035) );
  OAI222_X1 U21733 ( .A1(n18703), .A2(n18655), .B1(n18654), .B2(n18772), .C1(
        n18653), .C2(n18707), .ZN(P3_U3036) );
  OAI222_X1 U21734 ( .A1(n18703), .A2(n18657), .B1(n18656), .B2(n18772), .C1(
        n18655), .C2(n18707), .ZN(P3_U3037) );
  OAI222_X1 U21735 ( .A1(n18703), .A2(n18660), .B1(n18658), .B2(n18772), .C1(
        n18657), .C2(n18707), .ZN(P3_U3038) );
  OAI222_X1 U21736 ( .A1(n18660), .A2(n18707), .B1(n18659), .B2(n18772), .C1(
        n18661), .C2(n18703), .ZN(P3_U3039) );
  OAI222_X1 U21737 ( .A1(n18703), .A2(n18663), .B1(n18662), .B2(n18772), .C1(
        n18661), .C2(n18707), .ZN(P3_U3040) );
  INV_X1 U21738 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n18665) );
  OAI222_X1 U21739 ( .A1(n18703), .A2(n18665), .B1(n18664), .B2(n18772), .C1(
        n18663), .C2(n18707), .ZN(P3_U3041) );
  OAI222_X1 U21740 ( .A1(n18703), .A2(n18667), .B1(n18666), .B2(n18772), .C1(
        n18665), .C2(n18707), .ZN(P3_U3042) );
  OAI222_X1 U21741 ( .A1(n18703), .A2(n18669), .B1(n18668), .B2(n18772), .C1(
        n18667), .C2(n18707), .ZN(P3_U3043) );
  OAI222_X1 U21742 ( .A1(n18703), .A2(n18672), .B1(n18670), .B2(n18772), .C1(
        n18669), .C2(n18707), .ZN(P3_U3044) );
  OAI222_X1 U21743 ( .A1(n18672), .A2(n18707), .B1(n18671), .B2(n18772), .C1(
        n18673), .C2(n18703), .ZN(P3_U3045) );
  INV_X1 U21744 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n18675) );
  OAI222_X1 U21745 ( .A1(n18703), .A2(n18675), .B1(n18674), .B2(n18772), .C1(
        n18673), .C2(n18707), .ZN(P3_U3046) );
  INV_X1 U21746 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n18678) );
  OAI222_X1 U21747 ( .A1(n18703), .A2(n18678), .B1(n18676), .B2(n18772), .C1(
        n18675), .C2(n18707), .ZN(P3_U3047) );
  OAI222_X1 U21748 ( .A1(n18678), .A2(n18707), .B1(n18677), .B2(n18772), .C1(
        n18679), .C2(n18703), .ZN(P3_U3048) );
  OAI222_X1 U21749 ( .A1(n18703), .A2(n18681), .B1(n18680), .B2(n18772), .C1(
        n18679), .C2(n18707), .ZN(P3_U3049) );
  OAI222_X1 U21750 ( .A1(n18703), .A2(n18683), .B1(n18682), .B2(n18772), .C1(
        n18681), .C2(n18707), .ZN(P3_U3050) );
  OAI222_X1 U21751 ( .A1(n18703), .A2(n18686), .B1(n18684), .B2(n18772), .C1(
        n18683), .C2(n18707), .ZN(P3_U3051) );
  INV_X1 U21752 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n18687) );
  OAI222_X1 U21753 ( .A1(n18686), .A2(n18707), .B1(n18685), .B2(n18772), .C1(
        n18687), .C2(n18703), .ZN(P3_U3052) );
  INV_X1 U21754 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n18690) );
  OAI222_X1 U21755 ( .A1(n18703), .A2(n18690), .B1(n18688), .B2(n18772), .C1(
        n18687), .C2(n18707), .ZN(P3_U3053) );
  OAI222_X1 U21756 ( .A1(n18690), .A2(n18707), .B1(n18689), .B2(n18772), .C1(
        n18691), .C2(n18703), .ZN(P3_U3054) );
  OAI222_X1 U21757 ( .A1(n18703), .A2(n18693), .B1(n18692), .B2(n18772), .C1(
        n18691), .C2(n18707), .ZN(P3_U3055) );
  OAI222_X1 U21758 ( .A1(n18703), .A2(n18695), .B1(n18694), .B2(n18772), .C1(
        n18693), .C2(n18707), .ZN(P3_U3056) );
  OAI222_X1 U21759 ( .A1(n18703), .A2(n18697), .B1(n18696), .B2(n18772), .C1(
        n18695), .C2(n18707), .ZN(P3_U3057) );
  OAI222_X1 U21760 ( .A1(n18703), .A2(n18700), .B1(n18698), .B2(n18772), .C1(
        n18697), .C2(n18707), .ZN(P3_U3058) );
  OAI222_X1 U21761 ( .A1(n18700), .A2(n18707), .B1(n18699), .B2(n18772), .C1(
        n18701), .C2(n18703), .ZN(P3_U3059) );
  OAI222_X1 U21762 ( .A1(n18703), .A2(n18706), .B1(n18702), .B2(n18772), .C1(
        n18701), .C2(n18707), .ZN(P3_U3060) );
  OAI222_X1 U21763 ( .A1(n18707), .A2(n18706), .B1(n18705), .B2(n18772), .C1(
        n18704), .C2(n18703), .ZN(P3_U3061) );
  MUX2_X1 U21764 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .B(P3_BE_N_REG_3__SCAN_IN), .S(n18773), .Z(P3_U3274) );
  MUX2_X1 U21765 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .B(P3_BE_N_REG_2__SCAN_IN), .S(n18773), .Z(P3_U3275) );
  OAI22_X1 U21766 ( .A1(n18773), .A2(P3_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P3_BE_N_REG_1__SCAN_IN), .B2(n18772), .ZN(n18708) );
  INV_X1 U21767 ( .A(n18708), .ZN(P3_U3276) );
  OAI22_X1 U21768 ( .A1(n18773), .A2(P3_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P3_BE_N_REG_0__SCAN_IN), .B2(n18772), .ZN(n18709) );
  INV_X1 U21769 ( .A(n18709), .ZN(P3_U3277) );
  OAI21_X1 U21770 ( .B1(n18713), .B2(P3_DATAWIDTH_REG_0__SCAN_IN), .A(n18711), 
        .ZN(n18710) );
  INV_X1 U21771 ( .A(n18710), .ZN(P3_U3280) );
  INV_X1 U21772 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n18712) );
  OAI21_X1 U21773 ( .B1(n18713), .B2(n18712), .A(n18711), .ZN(P3_U3281) );
  OAI221_X1 U21774 ( .B1(n18716), .B2(P3_STATE2_REG_0__SCAN_IN), .C1(n18716), 
        .C2(n18715), .A(n18714), .ZN(P3_U3282) );
  INV_X1 U21775 ( .A(n18717), .ZN(n18718) );
  AOI22_X1 U21776 ( .A1(n18776), .A2(n18719), .B1(n18740), .B2(n18718), .ZN(
        n18724) );
  INV_X1 U21777 ( .A(n18720), .ZN(n18721) );
  AOI21_X1 U21778 ( .B1(n18776), .B2(n18721), .A(n18746), .ZN(n18723) );
  OAI22_X1 U21779 ( .A1(n18746), .A2(n18724), .B1(n18723), .B2(n18722), .ZN(
        P3_U3285) );
  INV_X1 U21780 ( .A(n18725), .ZN(n18730) );
  NOR2_X1 U21781 ( .A1(n18726), .A2(n18742), .ZN(n18734) );
  OAI22_X1 U21782 ( .A1(n18728), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n18727), .B2(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18733) );
  AOI222_X1 U21783 ( .A1(n18730), .A2(n18776), .B1(n18734), .B2(n18733), .C1(
        n18740), .C2(n18729), .ZN(n18731) );
  AOI22_X1 U21784 ( .A1(n18746), .A2(n18732), .B1(n18731), .B2(n18743), .ZN(
        P3_U3288) );
  INV_X1 U21785 ( .A(n18733), .ZN(n18735) );
  AOI222_X1 U21786 ( .A1(n18737), .A2(n18776), .B1(n18740), .B2(n18736), .C1(
        n18735), .C2(n18734), .ZN(n18738) );
  AOI22_X1 U21787 ( .A1(n18746), .A2(n18739), .B1(n18738), .B2(n18743), .ZN(
        P3_U3289) );
  AOI222_X1 U21788 ( .A1(n18742), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n18776), 
        .B2(n18741), .C1(n18745), .C2(n18740), .ZN(n18744) );
  AOI22_X1 U21789 ( .A1(n18746), .A2(n18745), .B1(n18744), .B2(n18743), .ZN(
        P3_U3290) );
  NOR2_X1 U21790 ( .A1(P3_DATAWIDTH_REG_1__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18747) );
  AOI211_X1 U21791 ( .C1(P3_DATAWIDTH_REG_0__SCAN_IN), .C2(n20968), .A(n18747), 
        .B(n18753), .ZN(n18751) );
  OAI22_X1 U21792 ( .A1(n18752), .A2(P3_BYTEENABLE_REG_2__SCAN_IN), .B1(n18749), .B2(n18748), .ZN(n18750) );
  NOR2_X1 U21793 ( .A1(n18751), .A2(n18750), .ZN(P3_U3292) );
  OAI22_X1 U21794 ( .A1(n18753), .A2(P3_REIP_REG_0__SCAN_IN), .B1(n18752), 
        .B2(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18754) );
  INV_X1 U21795 ( .A(n18754), .ZN(P3_U3293) );
  INV_X1 U21796 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n18755) );
  AOI22_X1 U21797 ( .A1(n18772), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n18755), 
        .B2(n18773), .ZN(P3_U3294) );
  MUX2_X1 U21798 ( .A(P3_MORE_REG_SCAN_IN), .B(n18757), .S(n18756), .Z(
        P3_U3295) );
  INV_X1 U21799 ( .A(n18758), .ZN(n18759) );
  OAI21_X1 U21800 ( .B1(P3_STATEBS16_REG_SCAN_IN), .B2(n18760), .A(n18759), 
        .ZN(n18762) );
  AOI211_X1 U21801 ( .C1(n18779), .C2(n18762), .A(n18761), .B(n18775), .ZN(
        n18765) );
  OAI21_X1 U21802 ( .B1(n18765), .B2(n18764), .A(n18763), .ZN(n18771) );
  AOI21_X1 U21803 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(
        P3_STATE2_REG_2__SCAN_IN), .A(n18766), .ZN(n18767) );
  AOI211_X1 U21804 ( .C1(n18769), .C2(n18768), .A(n18767), .B(n18783), .ZN(
        n18770) );
  MUX2_X1 U21805 ( .A(n18771), .B(P3_REQUESTPENDING_REG_SCAN_IN), .S(n18770), 
        .Z(P3_U3296) );
  OAI22_X1 U21806 ( .A1(n18773), .A2(P3_MEMORYFETCH_REG_SCAN_IN), .B1(
        P3_M_IO_N_REG_SCAN_IN), .B2(n18772), .ZN(n18774) );
  INV_X1 U21807 ( .A(n18774), .ZN(P3_U3297) );
  AOI21_X1 U21808 ( .B1(n18776), .B2(n18775), .A(P3_READREQUEST_REG_SCAN_IN), 
        .ZN(n18778) );
  AOI22_X1 U21809 ( .A1(n18783), .A2(n18779), .B1(n18778), .B2(n18777), .ZN(
        P3_U3298) );
  INV_X1 U21810 ( .A(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n18782) );
  OAI211_X1 U21811 ( .C1(n18783), .C2(n18782), .A(n18781), .B(n18780), .ZN(
        P3_U3299) );
  INV_X1 U21812 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n19725) );
  NAND2_X1 U21813 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19725), .ZN(n19715) );
  INV_X1 U21814 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n19709) );
  AOI22_X1 U21815 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n19715), .B1(
        P2_STATE_REG_1__SCAN_IN), .B2(n19709), .ZN(n19783) );
  AOI21_X1 U21816 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(P2_ADS_N_REG_SCAN_IN), 
        .A(n19783), .ZN(n18784) );
  INV_X1 U21817 ( .A(n18784), .ZN(P2_U2815) );
  AOI22_X1 U21818 ( .A1(n19838), .A2(P2_CODEFETCH_REG_SCAN_IN), .B1(n18785), 
        .B2(n19786), .ZN(n18786) );
  INV_X1 U21819 ( .A(n18786), .ZN(P2_U2816) );
  INV_X1 U21820 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n19718) );
  AOI22_X1 U21821 ( .A1(P2_D_C_N_REG_SCAN_IN), .A2(n19856), .B1(n19717), .B2(
        n19709), .ZN(n18787) );
  OAI21_X1 U21822 ( .B1(P2_CODEFETCH_REG_SCAN_IN), .B2(n19856), .A(n18787), 
        .ZN(P2_U2817) );
  OAI21_X1 U21823 ( .B1(n19717), .B2(BS16), .A(n19783), .ZN(n19781) );
  OAI21_X1 U21824 ( .B1(n19783), .B2(n19846), .A(n19781), .ZN(P2_U2818) );
  NOR2_X1 U21825 ( .A1(n18789), .A2(n18788), .ZN(n19824) );
  OAI21_X1 U21826 ( .B1(n19824), .B2(n21000), .A(n18790), .ZN(P2_U2819) );
  NOR4_X1 U21827 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_21__SCAN_IN), .A3(P2_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_23__SCAN_IN), .ZN(n18794) );
  NOR4_X1 U21828 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_17__SCAN_IN), .A3(P2_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_19__SCAN_IN), .ZN(n18793) );
  NOR4_X1 U21829 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n18792) );
  NOR4_X1 U21830 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_25__SCAN_IN), .A3(P2_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n18791) );
  NAND4_X1 U21831 ( .A1(n18794), .A2(n18793), .A3(n18792), .A4(n18791), .ZN(
        n18800) );
  NOR4_X1 U21832 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_2__SCAN_IN), .A3(P2_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_5__SCAN_IN), .ZN(n18798) );
  AOI211_X1 U21833 ( .C1(P2_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_0__SCAN_IN), .A(P2_DATAWIDTH_REG_4__SCAN_IN), .B(
        P2_DATAWIDTH_REG_16__SCAN_IN), .ZN(n18797) );
  NOR4_X1 U21834 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_11__SCAN_IN), .A3(P2_DATAWIDTH_REG_12__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_13__SCAN_IN), .ZN(n18796) );
  NOR4_X1 U21835 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_7__SCAN_IN), .A3(P2_DATAWIDTH_REG_8__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_9__SCAN_IN), .ZN(n18795) );
  NAND4_X1 U21836 ( .A1(n18798), .A2(n18797), .A3(n18796), .A4(n18795), .ZN(
        n18799) );
  NOR2_X1 U21837 ( .A1(n18800), .A2(n18799), .ZN(n18810) );
  INV_X1 U21838 ( .A(n18810), .ZN(n18808) );
  NOR2_X1 U21839 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n18808), .ZN(n18803) );
  INV_X1 U21840 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18801) );
  AOI22_X1 U21841 ( .A1(n18803), .A2(n10122), .B1(n18808), .B2(n18801), .ZN(
        P2_U2820) );
  OR3_X1 U21842 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18807) );
  INV_X1 U21843 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n18802) );
  AOI22_X1 U21844 ( .A1(n18803), .A2(n18807), .B1(n18808), .B2(n18802), .ZN(
        P2_U2821) );
  INV_X1 U21845 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19782) );
  NAND2_X1 U21846 ( .A1(n18803), .A2(n19782), .ZN(n18806) );
  OAI21_X1 U21847 ( .B1(n10122), .B2(n10543), .A(n18810), .ZN(n18804) );
  OAI21_X1 U21848 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n18810), .A(n18804), 
        .ZN(n18805) );
  OAI221_X1 U21849 ( .B1(n18806), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n18806), .C2(P2_REIP_REG_0__SCAN_IN), .A(n18805), .ZN(P2_U2822) );
  INV_X1 U21850 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n18809) );
  OAI221_X1 U21851 ( .B1(n18810), .B2(n18809), .C1(n18808), .C2(n18807), .A(
        n18806), .ZN(P2_U2823) );
  OAI22_X1 U21852 ( .A1(n18811), .A2(n18994), .B1(n19753), .B2(n18973), .ZN(
        n18812) );
  INV_X1 U21853 ( .A(n18812), .ZN(n18822) );
  AOI22_X1 U21854 ( .A1(P2_EBX_REG_21__SCAN_IN), .A2(n18990), .B1(
        P2_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n18964), .ZN(n18821) );
  OAI22_X1 U21855 ( .A1(n18814), .A2(n18981), .B1(n18813), .B2(n18982), .ZN(
        n18815) );
  INV_X1 U21856 ( .A(n18815), .ZN(n18820) );
  OAI211_X1 U21857 ( .C1(n18818), .C2(n18817), .A(n18999), .B(n18816), .ZN(
        n18819) );
  NAND4_X1 U21858 ( .A1(n18822), .A2(n18821), .A3(n18820), .A4(n18819), .ZN(
        P2_U2834) );
  AOI22_X1 U21859 ( .A1(n18823), .A2(n18950), .B1(P2_EBX_REG_20__SCAN_IN), 
        .B2(n18990), .ZN(n18833) );
  AOI22_X1 U21860 ( .A1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n19002), .B1(
        P2_REIP_REG_20__SCAN_IN), .B2(n18989), .ZN(n18832) );
  OAI22_X1 U21861 ( .A1(n18825), .A2(n18981), .B1(n18824), .B2(n18982), .ZN(
        n18826) );
  INV_X1 U21862 ( .A(n18826), .ZN(n18831) );
  OAI211_X1 U21863 ( .C1(n18829), .C2(n18828), .A(n18999), .B(n18827), .ZN(
        n18830) );
  NAND4_X1 U21864 ( .A1(n18833), .A2(n18832), .A3(n18831), .A4(n18830), .ZN(
        P2_U2835) );
  OAI21_X1 U21865 ( .B1(n21044), .B2(n18973), .A(n9889), .ZN(n18837) );
  OAI22_X1 U21866 ( .A1(n18835), .A2(n18994), .B1(n18834), .B2(n18987), .ZN(
        n18836) );
  AOI211_X1 U21867 ( .C1(P2_EBX_REG_19__SCAN_IN), .C2(n18990), .A(n18837), .B(
        n18836), .ZN(n18845) );
  AOI22_X1 U21868 ( .A1(n18839), .A2(n18997), .B1(n18991), .B2(n18838), .ZN(
        n18844) );
  OAI211_X1 U21869 ( .C1(n18842), .C2(n18841), .A(n18999), .B(n18840), .ZN(
        n18843) );
  NAND3_X1 U21870 ( .A1(n18845), .A2(n18844), .A3(n18843), .ZN(P2_U2836) );
  AOI22_X1 U21871 ( .A1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n18964), .B1(
        P2_REIP_REG_18__SCAN_IN), .B2(n18989), .ZN(n18846) );
  OAI21_X1 U21872 ( .B1(n18847), .B2(n18994), .A(n18846), .ZN(n18848) );
  AOI211_X1 U21873 ( .C1(P2_EBX_REG_18__SCAN_IN), .C2(n18990), .A(n18976), .B(
        n18848), .ZN(n18858) );
  INV_X1 U21874 ( .A(n18849), .ZN(n18850) );
  OAI22_X1 U21875 ( .A1(n18851), .A2(n18981), .B1(n18982), .B2(n18850), .ZN(
        n18852) );
  INV_X1 U21876 ( .A(n18852), .ZN(n18857) );
  OAI211_X1 U21877 ( .C1(n18855), .C2(n18854), .A(n18999), .B(n18853), .ZN(
        n18856) );
  NAND3_X1 U21878 ( .A1(n18858), .A2(n18857), .A3(n18856), .ZN(P2_U2837) );
  AOI22_X1 U21879 ( .A1(n18859), .A2(n18950), .B1(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n18964), .ZN(n18860) );
  OAI211_X1 U21880 ( .C1(n19748), .C2(n18973), .A(n18860), .B(n9889), .ZN(
        n18861) );
  AOI21_X1 U21881 ( .B1(P2_EBX_REG_17__SCAN_IN), .B2(n18990), .A(n18861), .ZN(
        n18869) );
  AOI22_X1 U21882 ( .A1(n18863), .A2(n18997), .B1(n18991), .B2(n18862), .ZN(
        n18868) );
  OAI211_X1 U21883 ( .C1(n18866), .C2(n18865), .A(n18999), .B(n18864), .ZN(
        n18867) );
  NAND3_X1 U21884 ( .A1(n18869), .A2(n18868), .A3(n18867), .ZN(P2_U2838) );
  INV_X1 U21885 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n19746) );
  OAI22_X1 U21886 ( .A1(n18870), .A2(n18994), .B1(n19746), .B2(n18973), .ZN(
        n18871) );
  AOI211_X1 U21887 ( .C1(P2_EBX_REG_16__SCAN_IN), .C2(n18990), .A(n18976), .B(
        n18871), .ZN(n18881) );
  NAND2_X1 U21888 ( .A1(n18873), .A2(n18872), .ZN(n18874) );
  XNOR2_X1 U21889 ( .A(n18875), .B(n18874), .ZN(n18879) );
  INV_X1 U21890 ( .A(n18876), .ZN(n18877) );
  OAI22_X1 U21891 ( .A1(n19010), .A2(n18981), .B1(n18982), .B2(n18877), .ZN(
        n18878) );
  AOI21_X1 U21892 ( .B1(n18999), .B2(n18879), .A(n18878), .ZN(n18880) );
  OAI211_X1 U21893 ( .C1(n18882), .C2(n18987), .A(n18881), .B(n18880), .ZN(
        P2_U2839) );
  INV_X1 U21894 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n18894) );
  OAI22_X1 U21895 ( .A1(n18883), .A2(n18994), .B1(n19744), .B2(n18973), .ZN(
        n18884) );
  AOI211_X1 U21896 ( .C1(P2_EBX_REG_15__SCAN_IN), .C2(n18990), .A(n18976), .B(
        n18884), .ZN(n18893) );
  NOR2_X1 U21897 ( .A1(n14665), .A2(n18885), .ZN(n18886) );
  XNOR2_X1 U21898 ( .A(n18887), .B(n18886), .ZN(n18891) );
  OAI22_X1 U21899 ( .A1(n18889), .A2(n18981), .B1(n18888), .B2(n18982), .ZN(
        n18890) );
  AOI21_X1 U21900 ( .B1(n18891), .B2(n18999), .A(n18890), .ZN(n18892) );
  OAI211_X1 U21901 ( .C1(n18894), .C2(n18987), .A(n18893), .B(n18892), .ZN(
        P2_U2840) );
  OAI211_X1 U21902 ( .C1(n18897), .C2(n18896), .A(n18999), .B(n18895), .ZN(
        n18899) );
  AOI22_X1 U21903 ( .A1(n18990), .A2(P2_EBX_REG_13__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n18964), .ZN(n18898) );
  OAI211_X1 U21904 ( .C1(n18900), .C2(n18994), .A(n18899), .B(n18898), .ZN(
        n18901) );
  AOI211_X1 U21905 ( .C1(P2_REIP_REG_13__SCAN_IN), .C2(n18989), .A(n18976), 
        .B(n18901), .ZN(n18905) );
  INV_X1 U21906 ( .A(n18922), .ZN(n19001) );
  AOI22_X1 U21907 ( .A1(n18903), .A2(n18997), .B1(n18902), .B2(n19001), .ZN(
        n18904) );
  OAI211_X1 U21908 ( .C1(n18982), .C2(n18906), .A(n18905), .B(n18904), .ZN(
        P2_U2842) );
  NAND2_X1 U21909 ( .A1(n18907), .A2(n18997), .ZN(n18910) );
  AOI22_X1 U21910 ( .A1(P2_EBX_REG_11__SCAN_IN), .A2(n18990), .B1(
        P2_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n18964), .ZN(n18909) );
  NAND2_X1 U21911 ( .A1(n18989), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n18908) );
  NAND4_X1 U21912 ( .A1(n18910), .A2(n18909), .A3(n9889), .A4(n18908), .ZN(
        n18911) );
  AOI21_X1 U21913 ( .B1(n18912), .B2(n18950), .A(n18911), .ZN(n18913) );
  OAI21_X1 U21914 ( .B1(n18914), .B2(n18982), .A(n18913), .ZN(n18915) );
  INV_X1 U21915 ( .A(n18915), .ZN(n18920) );
  NOR2_X1 U21916 ( .A1(n14665), .A2(n19705), .ZN(n18917) );
  OAI211_X1 U21917 ( .C1(n18918), .C2(n18921), .A(n18917), .B(n18916), .ZN(
        n18919) );
  OAI211_X1 U21918 ( .C1(n18922), .C2(n18921), .A(n18920), .B(n18919), .ZN(
        P2_U2844) );
  NAND2_X1 U21919 ( .A1(n12116), .A2(n18923), .ZN(n18925) );
  XOR2_X1 U21920 ( .A(n18925), .B(n18924), .Z(n18934) );
  OAI22_X1 U21921 ( .A1(n18927), .A2(n18994), .B1(n18926), .B2(n18973), .ZN(
        n18928) );
  INV_X1 U21922 ( .A(n18928), .ZN(n18929) );
  OAI211_X1 U21923 ( .C1(n18930), .C2(n18960), .A(n18929), .B(n9889), .ZN(
        n18932) );
  OAI22_X1 U21924 ( .A1(n19027), .A2(n18981), .B1(n18982), .B2(n19053), .ZN(
        n18931) );
  AOI211_X1 U21925 ( .C1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .C2(n18964), .A(
        n18932), .B(n18931), .ZN(n18933) );
  OAI21_X1 U21926 ( .B1(n18934), .B2(n19705), .A(n18933), .ZN(P2_U2845) );
  INV_X1 U21927 ( .A(n18935), .ZN(n18936) );
  OAI22_X1 U21928 ( .A1(n18936), .A2(n18994), .B1(n11075), .B2(n18960), .ZN(
        n18937) );
  AOI211_X1 U21929 ( .C1(P2_REIP_REG_9__SCAN_IN), .C2(n18989), .A(n18976), .B(
        n18937), .ZN(n18946) );
  NOR2_X1 U21930 ( .A1(n14665), .A2(n18938), .ZN(n18939) );
  XNOR2_X1 U21931 ( .A(n18940), .B(n18939), .ZN(n18944) );
  OAI22_X1 U21932 ( .A1(n18942), .A2(n18981), .B1(n18982), .B2(n18941), .ZN(
        n18943) );
  AOI21_X1 U21933 ( .B1(n18944), .B2(n18999), .A(n18943), .ZN(n18945) );
  OAI211_X1 U21934 ( .C1(n10049), .C2(n18987), .A(n18946), .B(n18945), .ZN(
        P2_U2846) );
  NOR2_X1 U21935 ( .A1(n14665), .A2(n18947), .ZN(n18948) );
  XOR2_X1 U21936 ( .A(n18949), .B(n18948), .Z(n18958) );
  AOI22_X1 U21937 ( .A1(n18951), .A2(n18950), .B1(n18989), .B2(
        P2_REIP_REG_7__SCAN_IN), .ZN(n18952) );
  OAI211_X1 U21938 ( .C1(n11061), .C2(n18960), .A(n18952), .B(n9889), .ZN(
        n18956) );
  OAI22_X1 U21939 ( .A1(n18954), .A2(n18982), .B1(n18981), .B2(n18953), .ZN(
        n18955) );
  AOI211_X1 U21940 ( .C1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .C2(n19002), .A(
        n18956), .B(n18955), .ZN(n18957) );
  OAI21_X1 U21941 ( .B1(n19705), .B2(n18958), .A(n18957), .ZN(P2_U2848) );
  OAI21_X1 U21942 ( .B1(n19732), .B2(n18973), .A(n9889), .ZN(n18963) );
  INV_X1 U21943 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n18959) );
  OAI22_X1 U21944 ( .A1(n18961), .A2(n18994), .B1(n18960), .B2(n18959), .ZN(
        n18962) );
  AOI211_X1 U21945 ( .C1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n18964), .A(
        n18963), .B(n18962), .ZN(n18971) );
  NAND2_X1 U21946 ( .A1(n12116), .A2(n18965), .ZN(n18966) );
  XNOR2_X1 U21947 ( .A(n18967), .B(n18966), .ZN(n18969) );
  AOI22_X1 U21948 ( .A1(n18969), .A2(n18999), .B1(n18997), .B2(n18968), .ZN(
        n18970) );
  OAI211_X1 U21949 ( .C1(n18982), .C2(n18972), .A(n18971), .B(n18970), .ZN(
        P2_U2849) );
  OAI22_X1 U21950 ( .A1(n18974), .A2(n18994), .B1(n13900), .B2(n18973), .ZN(
        n18975) );
  AOI211_X1 U21951 ( .C1(P2_EBX_REG_5__SCAN_IN), .C2(n18990), .A(n18976), .B(
        n18975), .ZN(n18986) );
  NOR2_X1 U21952 ( .A1(n14665), .A2(n18977), .ZN(n18978) );
  XNOR2_X1 U21953 ( .A(n18979), .B(n18978), .ZN(n18984) );
  OAI22_X1 U21954 ( .A1(n19060), .A2(n18982), .B1(n18981), .B2(n18980), .ZN(
        n18983) );
  AOI21_X1 U21955 ( .B1(n18984), .B2(n18999), .A(n18983), .ZN(n18985) );
  OAI211_X1 U21956 ( .C1(n18988), .C2(n18987), .A(n18986), .B(n18985), .ZN(
        P2_U2850) );
  AOI22_X1 U21957 ( .A1(n18990), .A2(P2_EBX_REG_0__SCAN_IN), .B1(n18989), .B2(
        P2_REIP_REG_0__SCAN_IN), .ZN(n18993) );
  NAND2_X1 U21958 ( .A1(n19088), .A2(n18991), .ZN(n18992) );
  OAI211_X1 U21959 ( .C1(n18995), .C2(n18994), .A(n18993), .B(n18992), .ZN(
        n18996) );
  AOI21_X1 U21960 ( .B1(n12319), .B2(n18997), .A(n18996), .ZN(n19005) );
  AOI22_X1 U21961 ( .A1(n19000), .A2(n18999), .B1(n19381), .B2(n18998), .ZN(
        n19004) );
  OAI21_X1 U21962 ( .B1(n19002), .B2(n19001), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n19003) );
  NAND3_X1 U21963 ( .A1(n19005), .A2(n19004), .A3(n19003), .ZN(P2_U2855) );
  OAI22_X1 U21964 ( .A1(n19007), .A2(n19031), .B1(n19020), .B2(n19006), .ZN(
        n19008) );
  INV_X1 U21965 ( .A(n19008), .ZN(n19009) );
  OAI21_X1 U21966 ( .B1(n19037), .B2(n19010), .A(n19009), .ZN(P2_U2871) );
  AOI21_X1 U21967 ( .B1(n13761), .B2(n19011), .A(n19031), .ZN(n19012) );
  AOI22_X1 U21968 ( .A1(n19012), .A2(n14745), .B1(P2_EBX_REG_14__SCAN_IN), 
        .B2(n19037), .ZN(n19013) );
  OAI21_X1 U21969 ( .B1(n19014), .B2(n19037), .A(n19013), .ZN(P2_U2873) );
  AOI21_X1 U21970 ( .B1(n13716), .B2(n19016), .A(n19015), .ZN(n19017) );
  OR3_X1 U21971 ( .A1(n13760), .A2(n19017), .A3(n19031), .ZN(n19018) );
  OAI21_X1 U21972 ( .B1(n19020), .B2(n19019), .A(n19018), .ZN(n19021) );
  INV_X1 U21973 ( .A(n19021), .ZN(n19022) );
  OAI21_X1 U21974 ( .B1(n19023), .B2(n19037), .A(n19022), .ZN(P2_U2875) );
  AOI211_X1 U21975 ( .C1(n19024), .C2(n13679), .A(n19031), .B(n13716), .ZN(
        n19025) );
  AOI21_X1 U21976 ( .B1(P2_EBX_REG_10__SCAN_IN), .B2(n19037), .A(n19025), .ZN(
        n19026) );
  OAI21_X1 U21977 ( .B1(n19027), .B2(n19037), .A(n19026), .ZN(P2_U2877) );
  INV_X1 U21978 ( .A(n19028), .ZN(n19033) );
  INV_X1 U21979 ( .A(n19029), .ZN(n19032) );
  AOI211_X1 U21980 ( .C1(n19033), .C2(n19032), .A(n19031), .B(n19030), .ZN(
        n19034) );
  AOI21_X1 U21981 ( .B1(P2_EBX_REG_8__SCAN_IN), .B2(n19037), .A(n19034), .ZN(
        n19035) );
  OAI21_X1 U21982 ( .B1(n19036), .B2(n19037), .A(n19035), .ZN(P2_U2879) );
  INV_X1 U21983 ( .A(n19065), .ZN(n19039) );
  AOI22_X1 U21984 ( .A1(n19039), .A2(n19038), .B1(P2_EBX_REG_4__SCAN_IN), .B2(
        n19037), .ZN(n19040) );
  OAI21_X1 U21985 ( .B1(n19037), .B2(n19041), .A(n19040), .ZN(P2_U2883) );
  INV_X1 U21986 ( .A(n19042), .ZN(n19047) );
  INV_X1 U21987 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n19043) );
  OAI22_X1 U21988 ( .A1(n19091), .A2(n19137), .B1(n19044), .B2(n19043), .ZN(
        n19045) );
  INV_X1 U21989 ( .A(n19045), .ZN(n19046) );
  OAI21_X1 U21990 ( .B1(n19061), .B2(n19047), .A(n19046), .ZN(P2_U2905) );
  INV_X1 U21991 ( .A(n19048), .ZN(n19134) );
  AOI22_X1 U21992 ( .A1(n19055), .A2(n19134), .B1(P2_EAX_REG_12__SCAN_IN), 
        .B2(n19083), .ZN(n19049) );
  OAI21_X1 U21993 ( .B1(n19061), .B2(n19050), .A(n19049), .ZN(P2_U2907) );
  AOI22_X1 U21994 ( .A1(n19055), .A2(n19051), .B1(P2_EAX_REG_10__SCAN_IN), 
        .B2(n19083), .ZN(n19052) );
  OAI21_X1 U21995 ( .B1(n19061), .B2(n19053), .A(n19052), .ZN(P2_U2909) );
  AOI22_X1 U21996 ( .A1(n19055), .A2(n19054), .B1(P2_EAX_REG_5__SCAN_IN), .B2(
        n19083), .ZN(n19059) );
  AOI21_X1 U21997 ( .B1(n19797), .B2(n19147), .A(n19056), .ZN(n19071) );
  XNOR2_X1 U21998 ( .A(n19788), .B(n21134), .ZN(n19072) );
  NOR2_X1 U21999 ( .A1(n19071), .A2(n19072), .ZN(n19070) );
  AOI21_X1 U22000 ( .B1(n19788), .B2(n21134), .A(n19070), .ZN(n19057) );
  NOR2_X1 U22001 ( .A1(n19057), .A2(n19063), .ZN(n19064) );
  OR3_X1 U22002 ( .A1(n19064), .A2(n19065), .A3(n19079), .ZN(n19058) );
  OAI211_X1 U22003 ( .C1(n19061), .C2(n19060), .A(n19059), .B(n19058), .ZN(
        P2_U2914) );
  INV_X1 U22004 ( .A(n19062), .ZN(n19168) );
  AOI22_X1 U22005 ( .A1(n19084), .A2(n19063), .B1(P2_EAX_REG_4__SCAN_IN), .B2(
        n19083), .ZN(n19068) );
  XOR2_X1 U22006 ( .A(n19065), .B(n19064), .Z(n19066) );
  NAND2_X1 U22007 ( .A1(n19066), .A2(n19086), .ZN(n19067) );
  OAI211_X1 U22008 ( .C1(n19168), .C2(n19091), .A(n19068), .B(n19067), .ZN(
        P2_U2915) );
  INV_X1 U22009 ( .A(n21134), .ZN(n19069) );
  AOI22_X1 U22010 ( .A1(n19069), .A2(n19084), .B1(P2_EAX_REG_3__SCAN_IN), .B2(
        n19083), .ZN(n19075) );
  AOI21_X1 U22011 ( .B1(n19072), .B2(n19071), .A(n19070), .ZN(n19073) );
  OR2_X1 U22012 ( .A1(n19073), .A2(n19079), .ZN(n19074) );
  OAI211_X1 U22013 ( .C1(n19076), .C2(n19091), .A(n19075), .B(n19074), .ZN(
        P2_U2916) );
  AOI22_X1 U22014 ( .A1(n19084), .A2(n19811), .B1(P2_EAX_REG_1__SCAN_IN), .B2(
        n19083), .ZN(n19082) );
  AOI21_X1 U22015 ( .B1(n19085), .B2(n19078), .A(n19077), .ZN(n19080) );
  OR2_X1 U22016 ( .A1(n19080), .A2(n19079), .ZN(n19081) );
  OAI211_X1 U22017 ( .C1(n19158), .C2(n19091), .A(n19082), .B(n19081), .ZN(
        P2_U2918) );
  AOI22_X1 U22018 ( .A1(n19084), .A2(n19088), .B1(P2_EAX_REG_0__SCAN_IN), .B2(
        n19083), .ZN(n19090) );
  INV_X1 U22019 ( .A(n19085), .ZN(n19087) );
  OAI211_X1 U22020 ( .C1(n19381), .C2(n19088), .A(n19087), .B(n19086), .ZN(
        n19089) );
  OAI211_X1 U22021 ( .C1(n19092), .C2(n19091), .A(n19090), .B(n19089), .ZN(
        P2_U2919) );
  NOR2_X1 U22022 ( .A1(n19093), .A2(n19099), .ZN(P2_U2920) );
  INV_X1 U22023 ( .A(n19094), .ZN(n19097) );
  AOI22_X1 U22024 ( .A1(n19097), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n19131), 
        .B2(P2_UWORD_REG_14__SCAN_IN), .ZN(n19095) );
  OAI21_X1 U22025 ( .B1(n19099), .B2(n19096), .A(n19095), .ZN(P2_U2921) );
  AOI22_X1 U22026 ( .A1(n19097), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n19131), 
        .B2(P2_UWORD_REG_12__SCAN_IN), .ZN(n19098) );
  OAI21_X1 U22027 ( .B1(n19100), .B2(n19099), .A(n19098), .ZN(P2_U2923) );
  AOI22_X1 U22028 ( .A1(n19131), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n19128), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n19101) );
  OAI21_X1 U22029 ( .B1(n19133), .B2(n13271), .A(n19101), .ZN(P2_U2936) );
  AOI22_X1 U22030 ( .A1(n19131), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n19128), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n19102) );
  OAI21_X1 U22031 ( .B1(n19133), .B2(n19043), .A(n19102), .ZN(P2_U2937) );
  AOI22_X1 U22032 ( .A1(n19131), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n19128), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n19103) );
  OAI21_X1 U22033 ( .B1(n19133), .B2(n19104), .A(n19103), .ZN(P2_U2938) );
  INV_X1 U22034 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n19106) );
  AOI22_X1 U22035 ( .A1(n19131), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n19128), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n19105) );
  OAI21_X1 U22036 ( .B1(n19133), .B2(n19106), .A(n19105), .ZN(P2_U2939) );
  AOI22_X1 U22037 ( .A1(n19131), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n19128), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n19107) );
  OAI21_X1 U22038 ( .B1(n19133), .B2(n19108), .A(n19107), .ZN(P2_U2940) );
  AOI22_X1 U22039 ( .A1(n19131), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n19128), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n19109) );
  OAI21_X1 U22040 ( .B1(n19133), .B2(n19110), .A(n19109), .ZN(P2_U2941) );
  AOI22_X1 U22041 ( .A1(n19131), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n19128), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n19111) );
  OAI21_X1 U22042 ( .B1(n19133), .B2(n19112), .A(n19111), .ZN(P2_U2942) );
  AOI22_X1 U22043 ( .A1(n19131), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n19128), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n19113) );
  OAI21_X1 U22044 ( .B1(n19133), .B2(n19114), .A(n19113), .ZN(P2_U2943) );
  AOI22_X1 U22045 ( .A1(n19131), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19128), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n19115) );
  OAI21_X1 U22046 ( .B1(n19133), .B2(n19116), .A(n19115), .ZN(P2_U2944) );
  AOI22_X1 U22047 ( .A1(n19131), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19128), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n19117) );
  OAI21_X1 U22048 ( .B1(n19133), .B2(n19118), .A(n19117), .ZN(P2_U2945) );
  INV_X1 U22049 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n19120) );
  AOI22_X1 U22050 ( .A1(n19131), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19128), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n19119) );
  OAI21_X1 U22051 ( .B1(n19133), .B2(n19120), .A(n19119), .ZN(P2_U2946) );
  INV_X1 U22052 ( .A(P2_LWORD_REG_4__SCAN_IN), .ZN(n20971) );
  AOI22_X1 U22053 ( .A1(P2_EAX_REG_4__SCAN_IN), .A2(n19121), .B1(n19128), .B2(
        P2_DATAO_REG_4__SCAN_IN), .ZN(n19122) );
  OAI21_X1 U22054 ( .B1(n20971), .B2(n19123), .A(n19122), .ZN(P2_U2947) );
  INV_X1 U22055 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n19125) );
  AOI22_X1 U22056 ( .A1(n19131), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n19128), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n19124) );
  OAI21_X1 U22057 ( .B1(n19133), .B2(n19125), .A(n19124), .ZN(P2_U2948) );
  INV_X1 U22058 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n19127) );
  AOI22_X1 U22059 ( .A1(n19131), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n19128), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n19126) );
  OAI21_X1 U22060 ( .B1(n19133), .B2(n19127), .A(n19126), .ZN(P2_U2949) );
  INV_X1 U22061 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n19130) );
  AOI22_X1 U22062 ( .A1(n19131), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19128), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n19129) );
  OAI21_X1 U22063 ( .B1(n19133), .B2(n19130), .A(n19129), .ZN(P2_U2950) );
  AOI22_X1 U22064 ( .A1(P2_LWORD_REG_0__SCAN_IN), .A2(n19131), .B1(n19128), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n19132) );
  OAI21_X1 U22065 ( .B1(n19133), .B2(n10817), .A(n19132), .ZN(P2_U2951) );
  AOI22_X1 U22066 ( .A1(n13338), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(
        P2_EAX_REG_28__SCAN_IN), .B2(n19143), .ZN(n19135) );
  NAND2_X1 U22067 ( .A1(n19139), .A2(n19134), .ZN(n19141) );
  NAND2_X1 U22068 ( .A1(n19135), .A2(n19141), .ZN(P2_U2964) );
  AOI22_X1 U22069 ( .A1(n13338), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(
        P2_EAX_REG_30__SCAN_IN), .B2(n19136), .ZN(n19140) );
  INV_X1 U22070 ( .A(n19137), .ZN(n19138) );
  NAND2_X1 U22071 ( .A1(n19139), .A2(n19138), .ZN(n19144) );
  NAND2_X1 U22072 ( .A1(n19140), .A2(n19144), .ZN(P2_U2966) );
  AOI22_X1 U22073 ( .A1(n13338), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(
        P2_EAX_REG_12__SCAN_IN), .B2(n19143), .ZN(n19142) );
  NAND2_X1 U22074 ( .A1(n19142), .A2(n19141), .ZN(P2_U2979) );
  AOI22_X1 U22075 ( .A1(n13338), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(
        P2_EAX_REG_14__SCAN_IN), .B2(n19143), .ZN(n19145) );
  NAND2_X1 U22076 ( .A1(n19145), .A2(n19144), .ZN(P2_U2981) );
  NOR2_X1 U22077 ( .A1(n19382), .A2(n19215), .ZN(n19180) );
  AOI22_X1 U22078 ( .A1(n19551), .A2(n19685), .B1(n19640), .B2(n19180), .ZN(
        n19157) );
  AOI21_X1 U22079 ( .B1(n19699), .B2(n19213), .A(n19846), .ZN(n19148) );
  INV_X1 U22080 ( .A(n19786), .ZN(n19789) );
  NOR2_X1 U22081 ( .A1(n19148), .A2(n19789), .ZN(n19152) );
  OAI21_X1 U22082 ( .B1(n19153), .B2(n19149), .A(n19796), .ZN(n19150) );
  AOI21_X1 U22083 ( .B1(n19152), .B2(n19644), .A(n19150), .ZN(n19151) );
  OAI21_X1 U22084 ( .B1(n19151), .B2(n19180), .A(n19647), .ZN(n19183) );
  INV_X1 U22085 ( .A(n19644), .ZN(n19691) );
  OAI21_X1 U22086 ( .B1(n19691), .B2(n19180), .A(n19152), .ZN(n19155) );
  OAI21_X1 U22087 ( .B1(n19153), .B2(n19180), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19154) );
  NAND2_X1 U22088 ( .A1(n19155), .A2(n19154), .ZN(n19182) );
  AOI22_X1 U22089 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n19183), .B1(
        n13777), .B2(n19182), .ZN(n19156) );
  OAI211_X1 U22090 ( .C1(n19554), .C2(n19213), .A(n19157), .B(n19156), .ZN(
        P2_U3048) );
  AOI22_X1 U22091 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n19178), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n19177), .ZN(n19658) );
  AOI22_X1 U22092 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n19178), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n19177), .ZN(n19614) );
  AOI22_X1 U22093 ( .A1(n19655), .A2(n19685), .B1(n19653), .B2(n19180), .ZN(
        n19160) );
  NOR2_X2 U22094 ( .A1(n19158), .A2(n19268), .ZN(n19654) );
  AOI22_X1 U22095 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n19183), .B1(
        n19654), .B2(n19182), .ZN(n19159) );
  OAI211_X1 U22096 ( .C1(n19658), .C2(n19213), .A(n19160), .B(n19159), .ZN(
        P2_U3049) );
  AOI22_X1 U22097 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n19178), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19177), .ZN(n19663) );
  AOI22_X1 U22098 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n19177), .B1(
        BUF1_REG_26__SCAN_IN), .B2(n19178), .ZN(n19489) );
  NOR2_X2 U22099 ( .A1(n10511), .A2(n19167), .ZN(n19659) );
  AOI22_X1 U22100 ( .A1(n19660), .A2(n19685), .B1(n19659), .B2(n19180), .ZN(
        n19164) );
  AOI22_X1 U22101 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n19183), .B1(
        n19162), .B2(n19182), .ZN(n19163) );
  OAI211_X1 U22102 ( .C1(n19663), .C2(n19213), .A(n19164), .B(n19163), .ZN(
        P2_U3050) );
  AOI22_X1 U22103 ( .A1(n19568), .A2(n19685), .B1(n19664), .B2(n19180), .ZN(
        n19166) );
  AOI22_X1 U22104 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19183), .B1(
        n19665), .B2(n19182), .ZN(n19165) );
  OAI211_X1 U22105 ( .C1(n19571), .C2(n19213), .A(n19166), .B(n19165), .ZN(
        P2_U3051) );
  AOI22_X1 U22106 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n19178), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n19177), .ZN(n19623) );
  AOI22_X1 U22107 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n19178), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n19177), .ZN(n19675) );
  NOR2_X2 U22108 ( .A1(n10371), .A2(n19167), .ZN(n19670) );
  AOI22_X1 U22109 ( .A1(n19620), .A2(n19685), .B1(n19670), .B2(n19180), .ZN(
        n19170) );
  NOR2_X2 U22110 ( .A1(n19168), .A2(n19268), .ZN(n19671) );
  AOI22_X1 U22111 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n19183), .B1(
        n19671), .B2(n19182), .ZN(n19169) );
  OAI211_X1 U22112 ( .C1(n19623), .C2(n19213), .A(n19170), .B(n19169), .ZN(
        P2_U3052) );
  AOI22_X1 U22113 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n19178), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n19177), .ZN(n19681) );
  AOI22_X1 U22114 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n19177), .B1(
        BUF1_REG_29__SCAN_IN), .B2(n19178), .ZN(n19627) );
  AOI22_X1 U22115 ( .A1(n19678), .A2(n19685), .B1(n19676), .B2(n19180), .ZN(
        n19173) );
  NOR2_X2 U22116 ( .A1(n19171), .A2(n19268), .ZN(n19677) );
  AOI22_X1 U22117 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19183), .B1(
        n19677), .B2(n19182), .ZN(n19172) );
  OAI211_X1 U22118 ( .C1(n19681), .C2(n19213), .A(n19173), .B(n19172), .ZN(
        P2_U3053) );
  AOI22_X1 U22119 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n19178), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n19177), .ZN(n19588) );
  AOI22_X1 U22120 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n19178), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n19177), .ZN(n19689) );
  AND2_X1 U22121 ( .A1(n12305), .A2(n19179), .ZN(n19682) );
  AOI22_X1 U22122 ( .A1(n19585), .A2(n19685), .B1(n19682), .B2(n19180), .ZN(
        n19176) );
  NOR2_X2 U22123 ( .A1(n19174), .A2(n19268), .ZN(n19683) );
  AOI22_X1 U22124 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19183), .B1(
        n19683), .B2(n19182), .ZN(n19175) );
  OAI211_X1 U22125 ( .C1(n19588), .C2(n19213), .A(n19176), .B(n19175), .ZN(
        P2_U3054) );
  AOI22_X1 U22126 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n19178), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n19177), .ZN(n19700) );
  AOI22_X1 U22127 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n19178), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n19177), .ZN(n19637) );
  AOI22_X1 U22128 ( .A1(n19694), .A2(n19685), .B1(n19690), .B2(n19180), .ZN(
        n19185) );
  NOR2_X2 U22129 ( .A1(n19181), .A2(n19268), .ZN(n19692) );
  AOI22_X1 U22130 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19183), .B1(
        n19692), .B2(n19182), .ZN(n19184) );
  OAI211_X1 U22131 ( .C1(n19700), .C2(n19213), .A(n19185), .B(n19184), .ZN(
        P2_U3055) );
  NOR2_X1 U22132 ( .A1(n19215), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19193) );
  INV_X1 U22133 ( .A(n19193), .ZN(n19186) );
  OR2_X1 U22134 ( .A1(n19186), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19188) );
  NAND2_X1 U22135 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19193), .ZN(
        n19190) );
  INV_X1 U22136 ( .A(n19190), .ZN(n19208) );
  NOR3_X1 U22137 ( .A1(n19187), .A2(n19208), .A3(n19149), .ZN(n19189) );
  AOI21_X1 U22138 ( .B1(n19149), .B2(n19188), .A(n19189), .ZN(n19209) );
  AOI22_X1 U22139 ( .A1(n19209), .A2(n13777), .B1(n19640), .B2(n19208), .ZN(
        n19195) );
  AOI211_X1 U22140 ( .C1(P2_STATE2_REG_3__SCAN_IN), .C2(n19190), .A(n19268), 
        .B(n19189), .ZN(n19191) );
  OAI221_X1 U22141 ( .B1(n19193), .B2(n19192), .C1(n19193), .C2(n19357), .A(
        n19191), .ZN(n19210) );
  AOI22_X1 U22142 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19210), .B1(
        n19237), .B2(n19649), .ZN(n19194) );
  OAI211_X1 U22143 ( .C1(n19652), .C2(n19213), .A(n19195), .B(n19194), .ZN(
        P2_U3056) );
  AOI22_X1 U22144 ( .A1(n19209), .A2(n19654), .B1(n19653), .B2(n19208), .ZN(
        n19197) );
  INV_X1 U22145 ( .A(n19658), .ZN(n19611) );
  AOI22_X1 U22146 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19210), .B1(
        n19237), .B2(n19611), .ZN(n19196) );
  OAI211_X1 U22147 ( .C1(n19614), .C2(n19213), .A(n19197), .B(n19196), .ZN(
        P2_U3057) );
  AOI22_X1 U22148 ( .A1(n19209), .A2(n19162), .B1(n19659), .B2(n19208), .ZN(
        n19199) );
  INV_X1 U22149 ( .A(n19663), .ZN(n19517) );
  AOI22_X1 U22150 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19210), .B1(
        n19237), .B2(n19517), .ZN(n19198) );
  OAI211_X1 U22151 ( .C1(n19489), .C2(n19213), .A(n19199), .B(n19198), .ZN(
        P2_U3058) );
  AOI22_X1 U22152 ( .A1(n19209), .A2(n19665), .B1(n19664), .B2(n19208), .ZN(
        n19201) );
  AOI22_X1 U22153 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19210), .B1(
        n19237), .B2(n19666), .ZN(n19200) );
  OAI211_X1 U22154 ( .C1(n19669), .C2(n19213), .A(n19201), .B(n19200), .ZN(
        P2_U3059) );
  AOI22_X1 U22155 ( .A1(n19209), .A2(n19671), .B1(n19670), .B2(n19208), .ZN(
        n19203) );
  INV_X1 U22156 ( .A(n19623), .ZN(n19672) );
  AOI22_X1 U22157 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19210), .B1(
        n19237), .B2(n19672), .ZN(n19202) );
  OAI211_X1 U22158 ( .C1(n19675), .C2(n19213), .A(n19203), .B(n19202), .ZN(
        P2_U3060) );
  AOI22_X1 U22159 ( .A1(n19209), .A2(n19677), .B1(n19676), .B2(n19208), .ZN(
        n19205) );
  INV_X1 U22160 ( .A(n19681), .ZN(n19624) );
  AOI22_X1 U22161 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19210), .B1(
        n19237), .B2(n19624), .ZN(n19204) );
  OAI211_X1 U22162 ( .C1(n19627), .C2(n19213), .A(n19205), .B(n19204), .ZN(
        P2_U3061) );
  AOI22_X1 U22163 ( .A1(n19209), .A2(n19683), .B1(n19682), .B2(n19208), .ZN(
        n19207) );
  INV_X1 U22164 ( .A(n19588), .ZN(n19684) );
  AOI22_X1 U22165 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19210), .B1(
        n19237), .B2(n19684), .ZN(n19206) );
  OAI211_X1 U22166 ( .C1(n19689), .C2(n19213), .A(n19207), .B(n19206), .ZN(
        P2_U3062) );
  AOI22_X1 U22167 ( .A1(n19209), .A2(n19692), .B1(n19690), .B2(n19208), .ZN(
        n19212) );
  INV_X1 U22168 ( .A(n19700), .ZN(n19631) );
  AOI22_X1 U22169 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19210), .B1(
        n19237), .B2(n19631), .ZN(n19211) );
  OAI211_X1 U22170 ( .C1(n19637), .C2(n19213), .A(n19212), .B(n19211), .ZN(
        P2_U3063) );
  NOR2_X1 U22171 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19214), .ZN(
        n19235) );
  OAI21_X1 U22172 ( .B1(n10732), .B2(n19235), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19216) );
  OR2_X1 U22173 ( .A1(n19445), .A2(n19215), .ZN(n19217) );
  NAND2_X1 U22174 ( .A1(n19216), .A2(n19217), .ZN(n19236) );
  AOI22_X1 U22175 ( .A1(n19236), .A2(n13777), .B1(n19640), .B2(n19235), .ZN(
        n19222) );
  AOI21_X1 U22176 ( .B1(n10686), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19220) );
  OAI21_X1 U22177 ( .B1(n19237), .B2(n19256), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19218) );
  NAND3_X1 U22178 ( .A1(n19218), .A2(n19786), .A3(n19217), .ZN(n19219) );
  OAI211_X1 U22179 ( .C1(n19235), .C2(n19220), .A(n19219), .B(n19647), .ZN(
        n19238) );
  AOI22_X1 U22180 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19238), .B1(
        n19237), .B2(n19551), .ZN(n19221) );
  OAI211_X1 U22181 ( .C1(n19554), .C2(n19246), .A(n19222), .B(n19221), .ZN(
        P2_U3064) );
  AOI22_X1 U22182 ( .A1(n19236), .A2(n19654), .B1(n19653), .B2(n19235), .ZN(
        n19224) );
  AOI22_X1 U22183 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19238), .B1(
        n19237), .B2(n19655), .ZN(n19223) );
  OAI211_X1 U22184 ( .C1(n19658), .C2(n19246), .A(n19224), .B(n19223), .ZN(
        P2_U3065) );
  AOI22_X1 U22185 ( .A1(n19236), .A2(n19162), .B1(n19659), .B2(n19235), .ZN(
        n19226) );
  AOI22_X1 U22186 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19238), .B1(
        n19237), .B2(n19660), .ZN(n19225) );
  OAI211_X1 U22187 ( .C1(n19663), .C2(n19246), .A(n19226), .B(n19225), .ZN(
        P2_U3066) );
  AOI22_X1 U22188 ( .A1(n19236), .A2(n19665), .B1(n19664), .B2(n19235), .ZN(
        n19228) );
  AOI22_X1 U22189 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19238), .B1(
        n19237), .B2(n19568), .ZN(n19227) );
  OAI211_X1 U22190 ( .C1(n19571), .C2(n19246), .A(n19228), .B(n19227), .ZN(
        P2_U3067) );
  AOI22_X1 U22191 ( .A1(n19236), .A2(n19671), .B1(n19670), .B2(n19235), .ZN(
        n19230) );
  AOI22_X1 U22192 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19238), .B1(
        n19237), .B2(n19620), .ZN(n19229) );
  OAI211_X1 U22193 ( .C1(n19623), .C2(n19246), .A(n19230), .B(n19229), .ZN(
        P2_U3068) );
  AOI22_X1 U22194 ( .A1(n19236), .A2(n19677), .B1(n19676), .B2(n19235), .ZN(
        n19232) );
  AOI22_X1 U22195 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19238), .B1(
        n19237), .B2(n19678), .ZN(n19231) );
  OAI211_X1 U22196 ( .C1(n19681), .C2(n19246), .A(n19232), .B(n19231), .ZN(
        P2_U3069) );
  AOI22_X1 U22197 ( .A1(n19236), .A2(n19683), .B1(n19682), .B2(n19235), .ZN(
        n19234) );
  AOI22_X1 U22198 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19238), .B1(
        n19237), .B2(n19585), .ZN(n19233) );
  OAI211_X1 U22199 ( .C1(n19588), .C2(n19246), .A(n19234), .B(n19233), .ZN(
        P2_U3070) );
  AOI22_X1 U22200 ( .A1(n19236), .A2(n19692), .B1(n19690), .B2(n19235), .ZN(
        n19240) );
  AOI22_X1 U22201 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19238), .B1(
        n19237), .B2(n19694), .ZN(n19239) );
  OAI211_X1 U22202 ( .C1(n19700), .C2(n19246), .A(n19240), .B(n19239), .ZN(
        P2_U3071) );
  AOI22_X1 U22203 ( .A1(n19655), .A2(n19256), .B1(n19255), .B2(n19653), .ZN(
        n19242) );
  AOI22_X1 U22204 ( .A1(n19654), .A2(n19257), .B1(n19289), .B2(n19611), .ZN(
        n19241) );
  OAI211_X1 U22205 ( .C1(n19243), .C2(n12465), .A(n19242), .B(n19241), .ZN(
        P2_U3073) );
  AOI22_X1 U22206 ( .A1(n19517), .A2(n19289), .B1(n19255), .B2(n19659), .ZN(
        n19245) );
  AOI22_X1 U22207 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19258), .B1(
        n19162), .B2(n19257), .ZN(n19244) );
  OAI211_X1 U22208 ( .C1(n19489), .C2(n19246), .A(n19245), .B(n19244), .ZN(
        P2_U3074) );
  AOI22_X1 U22209 ( .A1(n19568), .A2(n19256), .B1(n19255), .B2(n19664), .ZN(
        n19248) );
  AOI22_X1 U22210 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19258), .B1(
        n19665), .B2(n19257), .ZN(n19247) );
  OAI211_X1 U22211 ( .C1(n19571), .C2(n19261), .A(n19248), .B(n19247), .ZN(
        P2_U3075) );
  AOI22_X1 U22212 ( .A1(n19620), .A2(n19256), .B1(n19255), .B2(n19670), .ZN(
        n19250) );
  AOI22_X1 U22213 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19258), .B1(
        n19671), .B2(n19257), .ZN(n19249) );
  OAI211_X1 U22214 ( .C1(n19623), .C2(n19261), .A(n19250), .B(n19249), .ZN(
        P2_U3076) );
  AOI22_X1 U22215 ( .A1(n19678), .A2(n19256), .B1(n19255), .B2(n19676), .ZN(
        n19252) );
  AOI22_X1 U22216 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19258), .B1(
        n19677), .B2(n19257), .ZN(n19251) );
  OAI211_X1 U22217 ( .C1(n19681), .C2(n19261), .A(n19252), .B(n19251), .ZN(
        P2_U3077) );
  AOI22_X1 U22218 ( .A1(n19585), .A2(n19256), .B1(n19255), .B2(n19682), .ZN(
        n19254) );
  AOI22_X1 U22219 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19258), .B1(
        n19683), .B2(n19257), .ZN(n19253) );
  OAI211_X1 U22220 ( .C1(n19588), .C2(n19261), .A(n19254), .B(n19253), .ZN(
        P2_U3078) );
  AOI22_X1 U22221 ( .A1(n19694), .A2(n19256), .B1(n19255), .B2(n19690), .ZN(
        n19260) );
  AOI22_X1 U22222 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19258), .B1(
        n19692), .B2(n19257), .ZN(n19259) );
  OAI211_X1 U22223 ( .C1(n19700), .C2(n19261), .A(n19260), .B(n19259), .ZN(
        P2_U3079) );
  INV_X1 U22224 ( .A(n19262), .ZN(n19263) );
  NOR2_X1 U22225 ( .A1(n19263), .A2(n19321), .ZN(n19504) );
  NAND2_X1 U22226 ( .A1(n19504), .A2(n19794), .ZN(n19269) );
  NOR2_X1 U22227 ( .A1(n19382), .A2(n19264), .ZN(n19287) );
  OAI21_X1 U22228 ( .B1(n19265), .B2(n19287), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19266) );
  OAI21_X1 U22229 ( .B1(n19789), .B2(n19269), .A(n19266), .ZN(n19288) );
  AOI22_X1 U22230 ( .A1(n19288), .A2(n13777), .B1(n19640), .B2(n19287), .ZN(
        n19274) );
  AOI21_X1 U22231 ( .B1(n19267), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19272) );
  OAI21_X1 U22232 ( .B1(n19289), .B2(n19302), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19270) );
  AOI21_X1 U22233 ( .B1(n19270), .B2(n19269), .A(n19268), .ZN(n19271) );
  AOI22_X1 U22234 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19290), .B1(
        n19289), .B2(n19551), .ZN(n19273) );
  OAI211_X1 U22235 ( .C1(n19554), .C2(n19313), .A(n19274), .B(n19273), .ZN(
        P2_U3080) );
  AOI22_X1 U22236 ( .A1(n19288), .A2(n19654), .B1(n19653), .B2(n19287), .ZN(
        n19276) );
  AOI22_X1 U22237 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19290), .B1(
        n19289), .B2(n19655), .ZN(n19275) );
  OAI211_X1 U22238 ( .C1(n19658), .C2(n19313), .A(n19276), .B(n19275), .ZN(
        P2_U3081) );
  AOI22_X1 U22239 ( .A1(n19288), .A2(n19162), .B1(n19659), .B2(n19287), .ZN(
        n19278) );
  AOI22_X1 U22240 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19290), .B1(
        n19289), .B2(n19660), .ZN(n19277) );
  OAI211_X1 U22241 ( .C1(n19663), .C2(n19313), .A(n19278), .B(n19277), .ZN(
        P2_U3082) );
  AOI22_X1 U22242 ( .A1(n19288), .A2(n19665), .B1(n19664), .B2(n19287), .ZN(
        n19280) );
  AOI22_X1 U22243 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19290), .B1(
        n19289), .B2(n19568), .ZN(n19279) );
  OAI211_X1 U22244 ( .C1(n19571), .C2(n19313), .A(n19280), .B(n19279), .ZN(
        P2_U3083) );
  AOI22_X1 U22245 ( .A1(n19288), .A2(n19671), .B1(n19670), .B2(n19287), .ZN(
        n19282) );
  AOI22_X1 U22246 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19290), .B1(
        n19289), .B2(n19620), .ZN(n19281) );
  OAI211_X1 U22247 ( .C1(n19623), .C2(n19313), .A(n19282), .B(n19281), .ZN(
        P2_U3084) );
  AOI22_X1 U22248 ( .A1(n19288), .A2(n19677), .B1(n19676), .B2(n19287), .ZN(
        n19284) );
  AOI22_X1 U22249 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19290), .B1(
        n19289), .B2(n19678), .ZN(n19283) );
  OAI211_X1 U22250 ( .C1(n19681), .C2(n19313), .A(n19284), .B(n19283), .ZN(
        P2_U3085) );
  AOI22_X1 U22251 ( .A1(n19288), .A2(n19683), .B1(n19682), .B2(n19287), .ZN(
        n19286) );
  AOI22_X1 U22252 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19290), .B1(
        n19289), .B2(n19585), .ZN(n19285) );
  OAI211_X1 U22253 ( .C1(n19588), .C2(n19313), .A(n19286), .B(n19285), .ZN(
        P2_U3086) );
  AOI22_X1 U22254 ( .A1(n19288), .A2(n19692), .B1(n19690), .B2(n19287), .ZN(
        n19292) );
  AOI22_X1 U22255 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19290), .B1(
        n19289), .B2(n19694), .ZN(n19291) );
  OAI211_X1 U22256 ( .C1(n19700), .C2(n19313), .A(n19292), .B(n19291), .ZN(
        P2_U3087) );
  INV_X1 U22257 ( .A(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n19295) );
  AOI22_X1 U22258 ( .A1(n19655), .A2(n19302), .B1(n19308), .B2(n19653), .ZN(
        n19294) );
  AOI22_X1 U22259 ( .A1(n19654), .A2(n19309), .B1(n19347), .B2(n19611), .ZN(
        n19293) );
  OAI211_X1 U22260 ( .C1(n19305), .C2(n19295), .A(n19294), .B(n19293), .ZN(
        P2_U3089) );
  INV_X1 U22261 ( .A(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n19298) );
  AOI22_X1 U22262 ( .A1(n19660), .A2(n19302), .B1(n19308), .B2(n19659), .ZN(
        n19297) );
  AOI22_X1 U22263 ( .A1(n19162), .A2(n19309), .B1(n19347), .B2(n19517), .ZN(
        n19296) );
  OAI211_X1 U22264 ( .C1(n19305), .C2(n19298), .A(n19297), .B(n19296), .ZN(
        P2_U3090) );
  INV_X1 U22265 ( .A(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n19301) );
  AOI22_X1 U22266 ( .A1(n19620), .A2(n19302), .B1(n19308), .B2(n19670), .ZN(
        n19300) );
  AOI22_X1 U22267 ( .A1(n19671), .A2(n19309), .B1(n19347), .B2(n19672), .ZN(
        n19299) );
  OAI211_X1 U22268 ( .C1(n19305), .C2(n19301), .A(n19300), .B(n19299), .ZN(
        P2_U3092) );
  AOI22_X1 U22269 ( .A1(n19678), .A2(n19302), .B1(n19308), .B2(n19676), .ZN(
        n19304) );
  AOI22_X1 U22270 ( .A1(n19677), .A2(n19309), .B1(n19347), .B2(n19624), .ZN(
        n19303) );
  OAI211_X1 U22271 ( .C1(n19305), .C2(n10689), .A(n19304), .B(n19303), .ZN(
        P2_U3093) );
  AOI22_X1 U22272 ( .A1(n19684), .A2(n19347), .B1(n19308), .B2(n19682), .ZN(
        n19307) );
  AOI22_X1 U22273 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19310), .B1(
        n19683), .B2(n19309), .ZN(n19306) );
  OAI211_X1 U22274 ( .C1(n19689), .C2(n19313), .A(n19307), .B(n19306), .ZN(
        P2_U3094) );
  AOI22_X1 U22275 ( .A1(n19631), .A2(n19347), .B1(n19308), .B2(n19690), .ZN(
        n19312) );
  AOI22_X1 U22276 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19310), .B1(
        n19692), .B2(n19309), .ZN(n19311) );
  OAI211_X1 U22277 ( .C1(n19637), .C2(n19313), .A(n19312), .B(n19311), .ZN(
        P2_U3095) );
  NOR2_X2 U22278 ( .A1(n19642), .A2(n19314), .ZN(n19377) );
  OAI21_X1 U22279 ( .B1(n19347), .B2(n19377), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19320) );
  NAND2_X1 U22280 ( .A1(n19321), .A2(n19354), .ZN(n19319) );
  NAND2_X1 U22281 ( .A1(n19599), .A2(n19794), .ZN(n19359) );
  NOR2_X1 U22282 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19359), .ZN(
        n19345) );
  INV_X1 U22283 ( .A(n19345), .ZN(n19315) );
  NAND2_X1 U22284 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19315), .ZN(n19316) );
  NOR2_X1 U22285 ( .A1(n19317), .A2(n19316), .ZN(n19322) );
  OAI21_X1 U22286 ( .B1(n19345), .B2(n19796), .A(n19647), .ZN(n19318) );
  NAND3_X1 U22287 ( .A1(n19321), .A2(n19354), .A3(n19796), .ZN(n19323) );
  AOI21_X1 U22288 ( .B1(n19149), .B2(n19323), .A(n19322), .ZN(n19346) );
  AOI22_X1 U22289 ( .A1(n19346), .A2(n13777), .B1(n19640), .B2(n19345), .ZN(
        n19325) );
  AOI22_X1 U22290 ( .A1(n19347), .A2(n19551), .B1(n19377), .B2(n19649), .ZN(
        n19324) );
  OAI211_X1 U22291 ( .C1(n19351), .C2(n19326), .A(n19325), .B(n19324), .ZN(
        P2_U3096) );
  INV_X1 U22292 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n19329) );
  AOI22_X1 U22293 ( .A1(n19346), .A2(n19654), .B1(n19653), .B2(n19345), .ZN(
        n19328) );
  AOI22_X1 U22294 ( .A1(n19347), .A2(n19655), .B1(n19377), .B2(n19611), .ZN(
        n19327) );
  OAI211_X1 U22295 ( .C1(n19351), .C2(n19329), .A(n19328), .B(n19327), .ZN(
        P2_U3097) );
  INV_X1 U22296 ( .A(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n19332) );
  AOI22_X1 U22297 ( .A1(n19346), .A2(n19162), .B1(n19659), .B2(n19345), .ZN(
        n19331) );
  AOI22_X1 U22298 ( .A1(n19377), .A2(n19517), .B1(n19347), .B2(n19660), .ZN(
        n19330) );
  OAI211_X1 U22299 ( .C1(n19351), .C2(n19332), .A(n19331), .B(n19330), .ZN(
        P2_U3098) );
  INV_X1 U22300 ( .A(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n19335) );
  AOI22_X1 U22301 ( .A1(n19346), .A2(n19665), .B1(n19664), .B2(n19345), .ZN(
        n19334) );
  AOI22_X1 U22302 ( .A1(n19347), .A2(n19568), .B1(n19377), .B2(n19666), .ZN(
        n19333) );
  OAI211_X1 U22303 ( .C1(n19351), .C2(n19335), .A(n19334), .B(n19333), .ZN(
        P2_U3099) );
  INV_X1 U22304 ( .A(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n19338) );
  AOI22_X1 U22305 ( .A1(n19346), .A2(n19671), .B1(n19670), .B2(n19345), .ZN(
        n19337) );
  AOI22_X1 U22306 ( .A1(n19347), .A2(n19620), .B1(n19377), .B2(n19672), .ZN(
        n19336) );
  OAI211_X1 U22307 ( .C1(n19351), .C2(n19338), .A(n19337), .B(n19336), .ZN(
        P2_U3100) );
  INV_X1 U22308 ( .A(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n19341) );
  AOI22_X1 U22309 ( .A1(n19346), .A2(n19677), .B1(n19676), .B2(n19345), .ZN(
        n19340) );
  AOI22_X1 U22310 ( .A1(n19377), .A2(n19624), .B1(n19347), .B2(n19678), .ZN(
        n19339) );
  OAI211_X1 U22311 ( .C1(n19351), .C2(n19341), .A(n19340), .B(n19339), .ZN(
        P2_U3101) );
  INV_X1 U22312 ( .A(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n19344) );
  AOI22_X1 U22313 ( .A1(n19346), .A2(n19683), .B1(n19682), .B2(n19345), .ZN(
        n19343) );
  AOI22_X1 U22314 ( .A1(n19377), .A2(n19684), .B1(n19347), .B2(n19585), .ZN(
        n19342) );
  OAI211_X1 U22315 ( .C1(n19351), .C2(n19344), .A(n19343), .B(n19342), .ZN(
        P2_U3102) );
  INV_X1 U22316 ( .A(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n19350) );
  AOI22_X1 U22317 ( .A1(n19346), .A2(n19692), .B1(n19690), .B2(n19345), .ZN(
        n19349) );
  AOI22_X1 U22318 ( .A1(n19377), .A2(n19631), .B1(n19347), .B2(n19694), .ZN(
        n19348) );
  OAI211_X1 U22319 ( .C1(n19351), .C2(n19350), .A(n19349), .B(n19348), .ZN(
        P2_U3103) );
  INV_X1 U22320 ( .A(n19353), .ZN(n19472) );
  NAND2_X1 U22321 ( .A1(n19472), .A2(n19354), .ZN(n19385) );
  INV_X1 U22322 ( .A(n19385), .ZN(n19388) );
  OAI21_X1 U22323 ( .B1(n19355), .B2(n19388), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19356) );
  OAI21_X1 U22324 ( .B1(n19359), .B2(n19789), .A(n19356), .ZN(n19376) );
  AOI22_X1 U22325 ( .A1(n19376), .A2(n13777), .B1(n19640), .B2(n19388), .ZN(
        n19363) );
  NAND3_X1 U22326 ( .A1(n10695), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(n19385), 
        .ZN(n19361) );
  NAND2_X1 U22327 ( .A1(n19358), .A2(n19357), .ZN(n19790) );
  AOI22_X1 U22328 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19385), .B1(n19359), 
        .B2(n19790), .ZN(n19360) );
  NAND3_X1 U22329 ( .A1(n19361), .A2(n19360), .A3(n19647), .ZN(n19378) );
  AOI22_X1 U22330 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19378), .B1(
        n19377), .B2(n19551), .ZN(n19362) );
  OAI211_X1 U22331 ( .C1(n19554), .C2(n19412), .A(n19363), .B(n19362), .ZN(
        P2_U3104) );
  AOI22_X1 U22332 ( .A1(n19376), .A2(n19654), .B1(n19388), .B2(n19653), .ZN(
        n19365) );
  AOI22_X1 U22333 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19378), .B1(
        n19377), .B2(n19655), .ZN(n19364) );
  OAI211_X1 U22334 ( .C1(n19658), .C2(n19412), .A(n19365), .B(n19364), .ZN(
        P2_U3105) );
  AOI22_X1 U22335 ( .A1(n19376), .A2(n19162), .B1(n19388), .B2(n19659), .ZN(
        n19367) );
  AOI22_X1 U22336 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19378), .B1(
        n19377), .B2(n19660), .ZN(n19366) );
  OAI211_X1 U22337 ( .C1(n19663), .C2(n19412), .A(n19367), .B(n19366), .ZN(
        P2_U3106) );
  AOI22_X1 U22338 ( .A1(n19376), .A2(n19665), .B1(n19664), .B2(n19388), .ZN(
        n19369) );
  AOI22_X1 U22339 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19378), .B1(
        n19377), .B2(n19568), .ZN(n19368) );
  OAI211_X1 U22340 ( .C1(n19571), .C2(n19412), .A(n19369), .B(n19368), .ZN(
        P2_U3107) );
  AOI22_X1 U22341 ( .A1(n19376), .A2(n19671), .B1(n19388), .B2(n19670), .ZN(
        n19371) );
  AOI22_X1 U22342 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19378), .B1(
        n19377), .B2(n19620), .ZN(n19370) );
  OAI211_X1 U22343 ( .C1(n19623), .C2(n19412), .A(n19371), .B(n19370), .ZN(
        P2_U3108) );
  AOI22_X1 U22344 ( .A1(n19376), .A2(n19677), .B1(n19388), .B2(n19676), .ZN(
        n19373) );
  AOI22_X1 U22345 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19378), .B1(
        n19377), .B2(n19678), .ZN(n19372) );
  OAI211_X1 U22346 ( .C1(n19681), .C2(n19412), .A(n19373), .B(n19372), .ZN(
        P2_U3109) );
  AOI22_X1 U22347 ( .A1(n19376), .A2(n19683), .B1(n19388), .B2(n19682), .ZN(
        n19375) );
  AOI22_X1 U22348 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19378), .B1(
        n19377), .B2(n19585), .ZN(n19374) );
  OAI211_X1 U22349 ( .C1(n19588), .C2(n19412), .A(n19375), .B(n19374), .ZN(
        P2_U3110) );
  AOI22_X1 U22350 ( .A1(n19376), .A2(n19692), .B1(n19388), .B2(n19690), .ZN(
        n19380) );
  AOI22_X1 U22351 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19378), .B1(
        n19377), .B2(n19694), .ZN(n19379) );
  OAI211_X1 U22352 ( .C1(n19700), .C2(n19412), .A(n19380), .B(n19379), .ZN(
        P2_U3111) );
  INV_X1 U22353 ( .A(n19412), .ZN(n19400) );
  NOR2_X1 U22354 ( .A1(n19794), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n19474) );
  INV_X1 U22355 ( .A(n19474), .ZN(n19478) );
  NOR2_X1 U22356 ( .A1(n19382), .A2(n19478), .ZN(n19407) );
  AOI22_X1 U22357 ( .A1(n19551), .A2(n19400), .B1(n19640), .B2(n19407), .ZN(
        n19393) );
  AOI21_X1 U22358 ( .B1(n19432), .B2(n19412), .A(n19846), .ZN(n19383) );
  NOR2_X1 U22359 ( .A1(n19383), .A2(n19789), .ZN(n19387) );
  OAI21_X1 U22360 ( .B1(n19389), .B2(n19149), .A(n19796), .ZN(n19384) );
  AOI21_X1 U22361 ( .B1(n19387), .B2(n19385), .A(n19384), .ZN(n19386) );
  OAI21_X1 U22362 ( .B1(n19407), .B2(n19386), .A(n19647), .ZN(n19409) );
  OAI21_X1 U22363 ( .B1(n19388), .B2(n19407), .A(n19387), .ZN(n19391) );
  OAI21_X1 U22364 ( .B1(n19389), .B2(n19407), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19390) );
  NAND2_X1 U22365 ( .A1(n19391), .A2(n19390), .ZN(n19408) );
  AOI22_X1 U22366 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19409), .B1(
        n13777), .B2(n19408), .ZN(n19392) );
  OAI211_X1 U22367 ( .C1(n19554), .C2(n19432), .A(n19393), .B(n19392), .ZN(
        P2_U3112) );
  AOI22_X1 U22368 ( .A1(n19655), .A2(n19400), .B1(n19407), .B2(n19653), .ZN(
        n19395) );
  AOI22_X1 U22369 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19409), .B1(
        n19408), .B2(n19654), .ZN(n19394) );
  OAI211_X1 U22370 ( .C1(n19658), .C2(n19432), .A(n19395), .B(n19394), .ZN(
        P2_U3113) );
  AOI22_X1 U22371 ( .A1(n19517), .A2(n19438), .B1(n19659), .B2(n19407), .ZN(
        n19397) );
  AOI22_X1 U22372 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19409), .B1(
        n19408), .B2(n19162), .ZN(n19396) );
  OAI211_X1 U22373 ( .C1(n19489), .C2(n19412), .A(n19397), .B(n19396), .ZN(
        P2_U3114) );
  AOI22_X1 U22374 ( .A1(n19568), .A2(n19400), .B1(n19664), .B2(n19407), .ZN(
        n19399) );
  AOI22_X1 U22375 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19409), .B1(
        n19408), .B2(n19665), .ZN(n19398) );
  OAI211_X1 U22376 ( .C1(n19571), .C2(n19432), .A(n19399), .B(n19398), .ZN(
        P2_U3115) );
  AOI22_X1 U22377 ( .A1(n19620), .A2(n19400), .B1(n19670), .B2(n19407), .ZN(
        n19402) );
  AOI22_X1 U22378 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19409), .B1(
        n19408), .B2(n19671), .ZN(n19401) );
  OAI211_X1 U22379 ( .C1(n19623), .C2(n19432), .A(n19402), .B(n19401), .ZN(
        P2_U3116) );
  AOI22_X1 U22380 ( .A1(n19624), .A2(n19438), .B1(n19407), .B2(n19676), .ZN(
        n19404) );
  AOI22_X1 U22381 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19409), .B1(
        n19408), .B2(n19677), .ZN(n19403) );
  OAI211_X1 U22382 ( .C1(n19627), .C2(n19412), .A(n19404), .B(n19403), .ZN(
        P2_U3117) );
  AOI22_X1 U22383 ( .A1(n19684), .A2(n19438), .B1(n19407), .B2(n19682), .ZN(
        n19406) );
  AOI22_X1 U22384 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19409), .B1(
        n19408), .B2(n19683), .ZN(n19405) );
  OAI211_X1 U22385 ( .C1(n19689), .C2(n19412), .A(n19406), .B(n19405), .ZN(
        P2_U3118) );
  AOI22_X1 U22386 ( .A1(n19631), .A2(n19438), .B1(n19407), .B2(n19690), .ZN(
        n19411) );
  AOI22_X1 U22387 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19409), .B1(
        n19408), .B2(n19692), .ZN(n19410) );
  OAI211_X1 U22388 ( .C1(n19637), .C2(n19412), .A(n19411), .B(n19410), .ZN(
        P2_U3119) );
  NOR2_X1 U22389 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19478), .ZN(
        n19417) );
  NAND2_X1 U22390 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19417), .ZN(
        n19448) );
  INV_X1 U22391 ( .A(n19448), .ZN(n19437) );
  AOI22_X1 U22392 ( .A1(n19551), .A2(n19438), .B1(n19640), .B2(n19437), .ZN(
        n19423) );
  INV_X1 U22393 ( .A(n19788), .ZN(n19413) );
  NAND2_X1 U22394 ( .A1(n19413), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19643) );
  OAI21_X1 U22395 ( .B1(n19643), .B2(n19414), .A(n19786), .ZN(n19421) );
  OAI211_X1 U22396 ( .C1(n19415), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19448), 
        .B(n19789), .ZN(n19416) );
  OAI211_X1 U22397 ( .C1(n19421), .C2(n19417), .A(n19647), .B(n19416), .ZN(
        n19440) );
  INV_X1 U22398 ( .A(n19417), .ZN(n19420) );
  OAI21_X1 U22399 ( .B1(n19418), .B2(n19437), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19419) );
  OAI21_X1 U22400 ( .B1(n19421), .B2(n19420), .A(n19419), .ZN(n19439) );
  AOI22_X1 U22401 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19440), .B1(
        n13777), .B2(n19439), .ZN(n19422) );
  OAI211_X1 U22402 ( .C1(n19554), .C2(n19449), .A(n19423), .B(n19422), .ZN(
        P2_U3120) );
  AOI22_X1 U22403 ( .A1(n19655), .A2(n19438), .B1(n19437), .B2(n19653), .ZN(
        n19425) );
  AOI22_X1 U22404 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19440), .B1(
        n19654), .B2(n19439), .ZN(n19424) );
  OAI211_X1 U22405 ( .C1(n19658), .C2(n19449), .A(n19425), .B(n19424), .ZN(
        P2_U3121) );
  AOI22_X1 U22406 ( .A1(n19660), .A2(n19438), .B1(n19437), .B2(n19659), .ZN(
        n19427) );
  AOI22_X1 U22407 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19440), .B1(
        n19162), .B2(n19439), .ZN(n19426) );
  OAI211_X1 U22408 ( .C1(n19663), .C2(n19449), .A(n19427), .B(n19426), .ZN(
        P2_U3122) );
  AOI22_X1 U22409 ( .A1(n19568), .A2(n19438), .B1(n19664), .B2(n19437), .ZN(
        n19429) );
  AOI22_X1 U22410 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19440), .B1(
        n19665), .B2(n19439), .ZN(n19428) );
  OAI211_X1 U22411 ( .C1(n19571), .C2(n19449), .A(n19429), .B(n19428), .ZN(
        P2_U3123) );
  AOI22_X1 U22412 ( .A1(n19672), .A2(n19468), .B1(n19670), .B2(n19437), .ZN(
        n19431) );
  AOI22_X1 U22413 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19440), .B1(
        n19671), .B2(n19439), .ZN(n19430) );
  OAI211_X1 U22414 ( .C1(n19675), .C2(n19432), .A(n19431), .B(n19430), .ZN(
        P2_U3124) );
  AOI22_X1 U22415 ( .A1(n19678), .A2(n19438), .B1(n19437), .B2(n19676), .ZN(
        n19434) );
  AOI22_X1 U22416 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19440), .B1(
        n19677), .B2(n19439), .ZN(n19433) );
  OAI211_X1 U22417 ( .C1(n19681), .C2(n19449), .A(n19434), .B(n19433), .ZN(
        P2_U3125) );
  AOI22_X1 U22418 ( .A1(n19585), .A2(n19438), .B1(n19437), .B2(n19682), .ZN(
        n19436) );
  AOI22_X1 U22419 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19440), .B1(
        n19683), .B2(n19439), .ZN(n19435) );
  OAI211_X1 U22420 ( .C1(n19588), .C2(n19449), .A(n19436), .B(n19435), .ZN(
        P2_U3126) );
  AOI22_X1 U22421 ( .A1(n19694), .A2(n19438), .B1(n19437), .B2(n19690), .ZN(
        n19442) );
  AOI22_X1 U22422 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19440), .B1(
        n19692), .B2(n19439), .ZN(n19441) );
  OAI211_X1 U22423 ( .C1(n19700), .C2(n19449), .A(n19442), .B(n19441), .ZN(
        P2_U3127) );
  INV_X1 U22424 ( .A(n19598), .ZN(n19443) );
  NAND3_X1 U22425 ( .A1(n19821), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(
        n19474), .ZN(n19446) );
  INV_X1 U22426 ( .A(n19446), .ZN(n19466) );
  OAI21_X1 U22427 ( .B1(n10639), .B2(n19466), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19444) );
  OAI21_X1 U22428 ( .B1(n19478), .B2(n19445), .A(n19444), .ZN(n19467) );
  AOI22_X1 U22429 ( .A1(n19467), .A2(n13777), .B1(n19640), .B2(n19466), .ZN(
        n19453) );
  NAND3_X1 U22430 ( .A1(n10639), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(n19796), 
        .ZN(n19447) );
  NAND2_X1 U22431 ( .A1(n19447), .A2(n19446), .ZN(n19451) );
  OAI221_X1 U22432 ( .B1(n19846), .B2(n19503), .C1(n19846), .C2(n19449), .A(
        n19448), .ZN(n19450) );
  OAI221_X1 U22433 ( .B1(n19451), .B2(n19786), .C1(n19451), .C2(n19450), .A(
        n19647), .ZN(n19469) );
  AOI22_X1 U22434 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19469), .B1(
        n19468), .B2(n19551), .ZN(n19452) );
  OAI211_X1 U22435 ( .C1(n19554), .C2(n19503), .A(n19453), .B(n19452), .ZN(
        P2_U3128) );
  AOI22_X1 U22436 ( .A1(n19467), .A2(n19654), .B1(n19653), .B2(n19466), .ZN(
        n19455) );
  AOI22_X1 U22437 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19469), .B1(
        n19468), .B2(n19655), .ZN(n19454) );
  OAI211_X1 U22438 ( .C1(n19658), .C2(n19503), .A(n19455), .B(n19454), .ZN(
        P2_U3129) );
  AOI22_X1 U22439 ( .A1(n19467), .A2(n19162), .B1(n19659), .B2(n19466), .ZN(
        n19457) );
  AOI22_X1 U22440 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19469), .B1(
        n19468), .B2(n19660), .ZN(n19456) );
  OAI211_X1 U22441 ( .C1(n19663), .C2(n19503), .A(n19457), .B(n19456), .ZN(
        P2_U3130) );
  AOI22_X1 U22442 ( .A1(n19467), .A2(n19665), .B1(n19664), .B2(n19466), .ZN(
        n19459) );
  AOI22_X1 U22443 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19469), .B1(
        n19468), .B2(n19568), .ZN(n19458) );
  OAI211_X1 U22444 ( .C1(n19571), .C2(n19503), .A(n19459), .B(n19458), .ZN(
        P2_U3131) );
  AOI22_X1 U22445 ( .A1(n19467), .A2(n19671), .B1(n19670), .B2(n19466), .ZN(
        n19461) );
  AOI22_X1 U22446 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19469), .B1(
        n19468), .B2(n19620), .ZN(n19460) );
  OAI211_X1 U22447 ( .C1(n19623), .C2(n19503), .A(n19461), .B(n19460), .ZN(
        P2_U3132) );
  AOI22_X1 U22448 ( .A1(n19467), .A2(n19677), .B1(n19676), .B2(n19466), .ZN(
        n19463) );
  AOI22_X1 U22449 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19469), .B1(
        n19468), .B2(n19678), .ZN(n19462) );
  OAI211_X1 U22450 ( .C1(n19681), .C2(n19503), .A(n19463), .B(n19462), .ZN(
        P2_U3133) );
  AOI22_X1 U22451 ( .A1(n19467), .A2(n19683), .B1(n19682), .B2(n19466), .ZN(
        n19465) );
  AOI22_X1 U22452 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19469), .B1(
        n19468), .B2(n19585), .ZN(n19464) );
  OAI211_X1 U22453 ( .C1(n19588), .C2(n19503), .A(n19465), .B(n19464), .ZN(
        P2_U3134) );
  AOI22_X1 U22454 ( .A1(n19467), .A2(n19692), .B1(n19690), .B2(n19466), .ZN(
        n19471) );
  AOI22_X1 U22455 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19469), .B1(
        n19468), .B2(n19694), .ZN(n19470) );
  OAI211_X1 U22456 ( .C1(n19700), .C2(n19503), .A(n19471), .B(n19470), .ZN(
        P2_U3135) );
  NAND2_X1 U22457 ( .A1(n19474), .A2(n19472), .ZN(n19477) );
  NAND3_X1 U22458 ( .A1(n19473), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(n19477), 
        .ZN(n19479) );
  NAND2_X1 U22459 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19474), .ZN(
        n19475) );
  OAI21_X1 U22460 ( .B1(n19475), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19149), 
        .ZN(n19476) );
  INV_X1 U22461 ( .A(n19477), .ZN(n19498) );
  AOI22_X1 U22462 ( .A1(n19499), .A2(n13777), .B1(n19640), .B2(n19498), .ZN(
        n19484) );
  NOR3_X1 U22463 ( .A1(n19643), .A2(P2_STATE2_REG_3__SCAN_IN), .A3(n19482), 
        .ZN(n19481) );
  NOR3_X1 U22464 ( .A1(n19818), .A2(n19813), .A3(n19478), .ZN(n19480) );
  OAI211_X1 U22465 ( .C1(n19481), .C2(n19480), .A(n19647), .B(n19479), .ZN(
        n19500) );
  AOI22_X1 U22466 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19500), .B1(
        n19531), .B2(n19649), .ZN(n19483) );
  OAI211_X1 U22467 ( .C1(n19652), .C2(n19503), .A(n19484), .B(n19483), .ZN(
        P2_U3136) );
  AOI22_X1 U22468 ( .A1(n19499), .A2(n19654), .B1(n19653), .B2(n19498), .ZN(
        n19486) );
  AOI22_X1 U22469 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19500), .B1(
        n19531), .B2(n19611), .ZN(n19485) );
  OAI211_X1 U22470 ( .C1(n19614), .C2(n19503), .A(n19486), .B(n19485), .ZN(
        P2_U3137) );
  AOI22_X1 U22471 ( .A1(n19499), .A2(n19162), .B1(n19659), .B2(n19498), .ZN(
        n19488) );
  AOI22_X1 U22472 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19500), .B1(
        n19531), .B2(n19517), .ZN(n19487) );
  OAI211_X1 U22473 ( .C1(n19489), .C2(n19503), .A(n19488), .B(n19487), .ZN(
        P2_U3138) );
  AOI22_X1 U22474 ( .A1(n19499), .A2(n19665), .B1(n19664), .B2(n19498), .ZN(
        n19491) );
  AOI22_X1 U22475 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19500), .B1(
        n19531), .B2(n19666), .ZN(n19490) );
  OAI211_X1 U22476 ( .C1(n19669), .C2(n19503), .A(n19491), .B(n19490), .ZN(
        P2_U3139) );
  AOI22_X1 U22477 ( .A1(n19499), .A2(n19671), .B1(n19670), .B2(n19498), .ZN(
        n19493) );
  AOI22_X1 U22478 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19500), .B1(
        n19531), .B2(n19672), .ZN(n19492) );
  OAI211_X1 U22479 ( .C1(n19675), .C2(n19503), .A(n19493), .B(n19492), .ZN(
        P2_U3140) );
  AOI22_X1 U22480 ( .A1(n19499), .A2(n19677), .B1(n19676), .B2(n19498), .ZN(
        n19495) );
  AOI22_X1 U22481 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19500), .B1(
        n19531), .B2(n19624), .ZN(n19494) );
  OAI211_X1 U22482 ( .C1(n19627), .C2(n19503), .A(n19495), .B(n19494), .ZN(
        P2_U3141) );
  AOI22_X1 U22483 ( .A1(n19499), .A2(n19683), .B1(n19682), .B2(n19498), .ZN(
        n19497) );
  AOI22_X1 U22484 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19500), .B1(
        n19531), .B2(n19684), .ZN(n19496) );
  OAI211_X1 U22485 ( .C1(n19689), .C2(n19503), .A(n19497), .B(n19496), .ZN(
        P2_U3142) );
  AOI22_X1 U22486 ( .A1(n19499), .A2(n19692), .B1(n19690), .B2(n19498), .ZN(
        n19502) );
  AOI22_X1 U22487 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19500), .B1(
        n19531), .B2(n19631), .ZN(n19501) );
  OAI211_X1 U22488 ( .C1(n19637), .C2(n19503), .A(n19502), .B(n19501), .ZN(
        P2_U3143) );
  NOR2_X2 U22489 ( .A1(n19598), .A2(n19536), .ZN(n19594) );
  OAI21_X1 U22490 ( .B1(n19594), .B2(n19531), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19508) );
  NAND2_X1 U22491 ( .A1(n19504), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19509) );
  NAND3_X1 U22492 ( .A1(n19813), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19548) );
  NOR2_X1 U22493 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19548), .ZN(
        n19529) );
  INV_X1 U22494 ( .A(n19529), .ZN(n19505) );
  AND2_X1 U22495 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19505), .ZN(n19506) );
  NAND2_X1 U22496 ( .A1(n10701), .A2(n19506), .ZN(n19511) );
  OAI211_X1 U22497 ( .C1(n19529), .C2(n19796), .A(n19511), .B(n19647), .ZN(
        n19507) );
  INV_X1 U22498 ( .A(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n19514) );
  OAI21_X1 U22499 ( .B1(n19509), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19149), 
        .ZN(n19510) );
  AND2_X1 U22500 ( .A1(n19511), .A2(n19510), .ZN(n19530) );
  AOI22_X1 U22501 ( .A1(n19530), .A2(n13777), .B1(n19640), .B2(n19529), .ZN(
        n19513) );
  AOI22_X1 U22502 ( .A1(n19531), .A2(n19551), .B1(n19594), .B2(n19649), .ZN(
        n19512) );
  OAI211_X1 U22503 ( .C1(n19535), .C2(n19514), .A(n19513), .B(n19512), .ZN(
        P2_U3144) );
  AOI22_X1 U22504 ( .A1(n19530), .A2(n19654), .B1(n19653), .B2(n19529), .ZN(
        n19516) );
  AOI22_X1 U22505 ( .A1(n19531), .A2(n19655), .B1(n19594), .B2(n19611), .ZN(
        n19515) );
  OAI211_X1 U22506 ( .C1(n19535), .C2(n12474), .A(n19516), .B(n19515), .ZN(
        P2_U3145) );
  AOI22_X1 U22507 ( .A1(n19530), .A2(n19162), .B1(n19659), .B2(n19529), .ZN(
        n19519) );
  AOI22_X1 U22508 ( .A1(n19594), .A2(n19517), .B1(n19531), .B2(n19660), .ZN(
        n19518) );
  OAI211_X1 U22509 ( .C1(n19535), .C2(n12499), .A(n19519), .B(n19518), .ZN(
        P2_U3146) );
  AOI22_X1 U22510 ( .A1(n19530), .A2(n19665), .B1(n19664), .B2(n19529), .ZN(
        n19521) );
  AOI22_X1 U22511 ( .A1(n19531), .A2(n19568), .B1(n19594), .B2(n19666), .ZN(
        n19520) );
  OAI211_X1 U22512 ( .C1(n19535), .C2(n12526), .A(n19521), .B(n19520), .ZN(
        P2_U3147) );
  AOI22_X1 U22513 ( .A1(n19530), .A2(n19671), .B1(n19670), .B2(n19529), .ZN(
        n19523) );
  AOI22_X1 U22514 ( .A1(n19531), .A2(n19620), .B1(n19594), .B2(n19672), .ZN(
        n19522) );
  OAI211_X1 U22515 ( .C1(n19535), .C2(n12549), .A(n19523), .B(n19522), .ZN(
        P2_U3148) );
  AOI22_X1 U22516 ( .A1(n19530), .A2(n19677), .B1(n19676), .B2(n19529), .ZN(
        n19525) );
  AOI22_X1 U22517 ( .A1(n19594), .A2(n19624), .B1(n19531), .B2(n19678), .ZN(
        n19524) );
  OAI211_X1 U22518 ( .C1(n19535), .C2(n12582), .A(n19525), .B(n19524), .ZN(
        P2_U3149) );
  INV_X1 U22519 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n19528) );
  AOI22_X1 U22520 ( .A1(n19530), .A2(n19683), .B1(n19682), .B2(n19529), .ZN(
        n19527) );
  AOI22_X1 U22521 ( .A1(n19594), .A2(n19684), .B1(n19531), .B2(n19585), .ZN(
        n19526) );
  OAI211_X1 U22522 ( .C1(n19535), .C2(n19528), .A(n19527), .B(n19526), .ZN(
        P2_U3150) );
  INV_X1 U22523 ( .A(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n19534) );
  AOI22_X1 U22524 ( .A1(n19530), .A2(n19692), .B1(n19690), .B2(n19529), .ZN(
        n19533) );
  AOI22_X1 U22525 ( .A1(n19594), .A2(n19631), .B1(n19531), .B2(n19694), .ZN(
        n19532) );
  OAI211_X1 U22526 ( .C1(n19535), .C2(n19534), .A(n19533), .B(n19532), .ZN(
        P2_U3151) );
  NOR2_X1 U22527 ( .A1(n19821), .A2(n19548), .ZN(n19601) );
  INV_X1 U22528 ( .A(n19601), .ZN(n19589) );
  NAND2_X1 U22529 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19589), .ZN(n19538) );
  NOR2_X1 U22530 ( .A1(n19539), .A2(n19538), .ZN(n19547) );
  INV_X1 U22531 ( .A(n19548), .ZN(n19540) );
  AOI21_X1 U22532 ( .B1(n19796), .B2(n19540), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19541) );
  INV_X1 U22533 ( .A(n13777), .ZN(n19543) );
  INV_X1 U22534 ( .A(n19640), .ZN(n19542) );
  OAI22_X1 U22535 ( .A1(n19592), .A2(n19543), .B1(n19542), .B2(n19589), .ZN(
        n19544) );
  INV_X1 U22536 ( .A(n19544), .ZN(n19553) );
  INV_X1 U22537 ( .A(n19643), .ZN(n19546) );
  NAND2_X1 U22538 ( .A1(n19546), .A2(n19545), .ZN(n19549) );
  AOI21_X1 U22539 ( .B1(n19549), .B2(n19548), .A(n19547), .ZN(n19550) );
  OAI211_X1 U22540 ( .C1(n19601), .C2(n19796), .A(n19550), .B(n19647), .ZN(
        n19595) );
  AOI22_X1 U22541 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19595), .B1(
        n19594), .B2(n19551), .ZN(n19552) );
  OAI211_X1 U22542 ( .C1(n19554), .C2(n19636), .A(n19553), .B(n19552), .ZN(
        P2_U3152) );
  INV_X1 U22543 ( .A(n19654), .ZN(n19556) );
  INV_X1 U22544 ( .A(n19653), .ZN(n19555) );
  OAI22_X1 U22545 ( .A1(n19592), .A2(n19556), .B1(n19555), .B2(n19589), .ZN(
        n19557) );
  INV_X1 U22546 ( .A(n19557), .ZN(n19559) );
  AOI22_X1 U22547 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19595), .B1(
        n19594), .B2(n19655), .ZN(n19558) );
  OAI211_X1 U22548 ( .C1(n19658), .C2(n19636), .A(n19559), .B(n19558), .ZN(
        P2_U3153) );
  INV_X1 U22549 ( .A(n19162), .ZN(n19561) );
  INV_X1 U22550 ( .A(n19659), .ZN(n19560) );
  OAI22_X1 U22551 ( .A1(n19592), .A2(n19561), .B1(n19560), .B2(n19589), .ZN(
        n19562) );
  INV_X1 U22552 ( .A(n19562), .ZN(n19564) );
  AOI22_X1 U22553 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19595), .B1(
        n19594), .B2(n19660), .ZN(n19563) );
  OAI211_X1 U22554 ( .C1(n19663), .C2(n19636), .A(n19564), .B(n19563), .ZN(
        P2_U3154) );
  INV_X1 U22555 ( .A(n19665), .ZN(n19566) );
  INV_X1 U22556 ( .A(n19664), .ZN(n19565) );
  OAI22_X1 U22557 ( .A1(n19592), .A2(n19566), .B1(n19565), .B2(n19589), .ZN(
        n19567) );
  INV_X1 U22558 ( .A(n19567), .ZN(n19570) );
  AOI22_X1 U22559 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19595), .B1(
        n19594), .B2(n19568), .ZN(n19569) );
  OAI211_X1 U22560 ( .C1(n19571), .C2(n19636), .A(n19570), .B(n19569), .ZN(
        P2_U3155) );
  INV_X1 U22561 ( .A(n19671), .ZN(n19573) );
  INV_X1 U22562 ( .A(n19670), .ZN(n19572) );
  OAI22_X1 U22563 ( .A1(n19592), .A2(n19573), .B1(n19572), .B2(n19589), .ZN(
        n19574) );
  INV_X1 U22564 ( .A(n19574), .ZN(n19576) );
  AOI22_X1 U22565 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19595), .B1(
        n19594), .B2(n19620), .ZN(n19575) );
  OAI211_X1 U22566 ( .C1(n19623), .C2(n19636), .A(n19576), .B(n19575), .ZN(
        P2_U3156) );
  INV_X1 U22567 ( .A(n19677), .ZN(n19578) );
  INV_X1 U22568 ( .A(n19676), .ZN(n19577) );
  OAI22_X1 U22569 ( .A1(n19592), .A2(n19578), .B1(n19577), .B2(n19589), .ZN(
        n19579) );
  INV_X1 U22570 ( .A(n19579), .ZN(n19581) );
  AOI22_X1 U22571 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19595), .B1(
        n19594), .B2(n19678), .ZN(n19580) );
  OAI211_X1 U22572 ( .C1(n19681), .C2(n19636), .A(n19581), .B(n19580), .ZN(
        P2_U3157) );
  INV_X1 U22573 ( .A(n19683), .ZN(n19583) );
  INV_X1 U22574 ( .A(n19682), .ZN(n19582) );
  OAI22_X1 U22575 ( .A1(n19592), .A2(n19583), .B1(n19582), .B2(n19589), .ZN(
        n19584) );
  INV_X1 U22576 ( .A(n19584), .ZN(n19587) );
  AOI22_X1 U22577 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19595), .B1(
        n19594), .B2(n19585), .ZN(n19586) );
  OAI211_X1 U22578 ( .C1(n19588), .C2(n19636), .A(n19587), .B(n19586), .ZN(
        P2_U3158) );
  INV_X1 U22579 ( .A(n19692), .ZN(n19591) );
  INV_X1 U22580 ( .A(n19690), .ZN(n19590) );
  OAI22_X1 U22581 ( .A1(n19592), .A2(n19591), .B1(n19590), .B2(n19589), .ZN(
        n19593) );
  INV_X1 U22582 ( .A(n19593), .ZN(n19597) );
  AOI22_X1 U22583 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19595), .B1(
        n19594), .B2(n19694), .ZN(n19596) );
  OAI211_X1 U22584 ( .C1(n19700), .C2(n19636), .A(n19597), .B(n19596), .ZN(
        P2_U3159) );
  NAND2_X1 U22585 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19599), .ZN(
        n19641) );
  NOR2_X1 U22586 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19641), .ZN(
        n19630) );
  AOI22_X1 U22587 ( .A1(n19649), .A2(n19695), .B1(n19640), .B2(n19630), .ZN(
        n19610) );
  OAI21_X1 U22588 ( .B1(n19695), .B2(n19619), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19600) );
  NAND2_X1 U22589 ( .A1(n19600), .A2(n19786), .ZN(n19608) );
  NOR2_X1 U22590 ( .A1(n19630), .A2(n19601), .ZN(n19607) );
  INV_X1 U22591 ( .A(n19607), .ZN(n19604) );
  INV_X1 U22592 ( .A(n19630), .ZN(n19602) );
  OAI211_X1 U22593 ( .C1(n10702), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19602), 
        .B(n19789), .ZN(n19603) );
  OAI211_X1 U22594 ( .C1(n19608), .C2(n19604), .A(n19647), .B(n19603), .ZN(
        n19633) );
  OAI21_X1 U22595 ( .B1(n19605), .B2(n19630), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19606) );
  AOI22_X1 U22596 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19633), .B1(
        n13777), .B2(n19632), .ZN(n19609) );
  OAI211_X1 U22597 ( .C1(n19652), .C2(n19636), .A(n19610), .B(n19609), .ZN(
        P2_U3160) );
  AOI22_X1 U22598 ( .A1(n19611), .A2(n19695), .B1(n19630), .B2(n19653), .ZN(
        n19613) );
  AOI22_X1 U22599 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19633), .B1(
        n19654), .B2(n19632), .ZN(n19612) );
  OAI211_X1 U22600 ( .C1(n19614), .C2(n19636), .A(n19613), .B(n19612), .ZN(
        P2_U3161) );
  AOI22_X1 U22601 ( .A1(n19660), .A2(n19619), .B1(n19659), .B2(n19630), .ZN(
        n19616) );
  AOI22_X1 U22602 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19633), .B1(
        n19162), .B2(n19632), .ZN(n19615) );
  OAI211_X1 U22603 ( .C1(n19663), .C2(n19688), .A(n19616), .B(n19615), .ZN(
        P2_U3162) );
  AOI22_X1 U22604 ( .A1(n19666), .A2(n19695), .B1(n19664), .B2(n19630), .ZN(
        n19618) );
  AOI22_X1 U22605 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19633), .B1(
        n19665), .B2(n19632), .ZN(n19617) );
  OAI211_X1 U22606 ( .C1(n19669), .C2(n19636), .A(n19618), .B(n19617), .ZN(
        P2_U3163) );
  AOI22_X1 U22607 ( .A1(n19620), .A2(n19619), .B1(n19670), .B2(n19630), .ZN(
        n19622) );
  AOI22_X1 U22608 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19633), .B1(
        n19671), .B2(n19632), .ZN(n19621) );
  OAI211_X1 U22609 ( .C1(n19623), .C2(n19688), .A(n19622), .B(n19621), .ZN(
        P2_U3164) );
  AOI22_X1 U22610 ( .A1(n19624), .A2(n19695), .B1(n19630), .B2(n19676), .ZN(
        n19626) );
  AOI22_X1 U22611 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19633), .B1(
        n19677), .B2(n19632), .ZN(n19625) );
  OAI211_X1 U22612 ( .C1(n19627), .C2(n19636), .A(n19626), .B(n19625), .ZN(
        P2_U3165) );
  AOI22_X1 U22613 ( .A1(n19684), .A2(n19695), .B1(n19630), .B2(n19682), .ZN(
        n19629) );
  AOI22_X1 U22614 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19633), .B1(
        n19683), .B2(n19632), .ZN(n19628) );
  OAI211_X1 U22615 ( .C1(n19689), .C2(n19636), .A(n19629), .B(n19628), .ZN(
        P2_U3166) );
  AOI22_X1 U22616 ( .A1(n19631), .A2(n19695), .B1(n19630), .B2(n19690), .ZN(
        n19635) );
  AOI22_X1 U22617 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19633), .B1(
        n19692), .B2(n19632), .ZN(n19634) );
  OAI211_X1 U22618 ( .C1(n19637), .C2(n19636), .A(n19635), .B(n19634), .ZN(
        P2_U3167) );
  OAI21_X1 U22619 ( .B1(n19638), .B2(n19691), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19639) );
  OAI21_X1 U22620 ( .B1(n19641), .B2(n19789), .A(n19639), .ZN(n19693) );
  AOI22_X1 U22621 ( .A1(n19693), .A2(n13777), .B1(n19691), .B2(n19640), .ZN(
        n19651) );
  OAI21_X1 U22622 ( .B1(n19643), .B2(n19642), .A(n19641), .ZN(n19648) );
  OAI211_X1 U22623 ( .C1(n19645), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19789), 
        .B(n19644), .ZN(n19646) );
  NAND3_X1 U22624 ( .A1(n19648), .A2(n19647), .A3(n19646), .ZN(n19696) );
  AOI22_X1 U22625 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19696), .B1(
        n19685), .B2(n19649), .ZN(n19650) );
  OAI211_X1 U22626 ( .C1(n19652), .C2(n19688), .A(n19651), .B(n19650), .ZN(
        P2_U3168) );
  AOI22_X1 U22627 ( .A1(n19693), .A2(n19654), .B1(n19691), .B2(n19653), .ZN(
        n19657) );
  AOI22_X1 U22628 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19696), .B1(
        n19695), .B2(n19655), .ZN(n19656) );
  OAI211_X1 U22629 ( .C1(n19658), .C2(n19699), .A(n19657), .B(n19656), .ZN(
        P2_U3169) );
  AOI22_X1 U22630 ( .A1(n19693), .A2(n19162), .B1(n19691), .B2(n19659), .ZN(
        n19662) );
  AOI22_X1 U22631 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19696), .B1(
        n19695), .B2(n19660), .ZN(n19661) );
  OAI211_X1 U22632 ( .C1(n19663), .C2(n19699), .A(n19662), .B(n19661), .ZN(
        P2_U3170) );
  AOI22_X1 U22633 ( .A1(n19693), .A2(n19665), .B1(n19691), .B2(n19664), .ZN(
        n19668) );
  AOI22_X1 U22634 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19696), .B1(
        n19685), .B2(n19666), .ZN(n19667) );
  OAI211_X1 U22635 ( .C1(n19669), .C2(n19688), .A(n19668), .B(n19667), .ZN(
        P2_U3171) );
  AOI22_X1 U22636 ( .A1(n19693), .A2(n19671), .B1(n19691), .B2(n19670), .ZN(
        n19674) );
  AOI22_X1 U22637 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19696), .B1(
        n19685), .B2(n19672), .ZN(n19673) );
  OAI211_X1 U22638 ( .C1(n19675), .C2(n19688), .A(n19674), .B(n19673), .ZN(
        P2_U3172) );
  AOI22_X1 U22639 ( .A1(n19693), .A2(n19677), .B1(n19691), .B2(n19676), .ZN(
        n19680) );
  AOI22_X1 U22640 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19696), .B1(
        n19695), .B2(n19678), .ZN(n19679) );
  OAI211_X1 U22641 ( .C1(n19681), .C2(n19699), .A(n19680), .B(n19679), .ZN(
        P2_U3173) );
  AOI22_X1 U22642 ( .A1(n19693), .A2(n19683), .B1(n19691), .B2(n19682), .ZN(
        n19687) );
  AOI22_X1 U22643 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19696), .B1(
        n19685), .B2(n19684), .ZN(n19686) );
  OAI211_X1 U22644 ( .C1(n19689), .C2(n19688), .A(n19687), .B(n19686), .ZN(
        P2_U3174) );
  AOI22_X1 U22645 ( .A1(n19693), .A2(n19692), .B1(n19691), .B2(n19690), .ZN(
        n19698) );
  AOI22_X1 U22646 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19696), .B1(
        n19695), .B2(n19694), .ZN(n19697) );
  OAI211_X1 U22647 ( .C1(n19700), .C2(n19699), .A(n19698), .B(n19697), .ZN(
        P2_U3175) );
  AOI21_X1 U22648 ( .B1(n19784), .B2(n19701), .A(n19840), .ZN(n19706) );
  INV_X1 U22649 ( .A(n19702), .ZN(n19703) );
  OAI211_X1 U22650 ( .C1(n19707), .C2(n19703), .A(n19844), .B(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n19704) );
  OAI211_X1 U22651 ( .C1(n19707), .C2(n19706), .A(n19705), .B(n19704), .ZN(
        P2_U3177) );
  AND2_X1 U22652 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n19708), .ZN(
        P2_U3179) );
  AND2_X1 U22653 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n19708), .ZN(
        P2_U3180) );
  AND2_X1 U22654 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n19708), .ZN(
        P2_U3181) );
  AND2_X1 U22655 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n19708), .ZN(
        P2_U3182) );
  AND2_X1 U22656 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n19708), .ZN(
        P2_U3183) );
  AND2_X1 U22657 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n19708), .ZN(
        P2_U3184) );
  AND2_X1 U22658 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n19708), .ZN(
        P2_U3185) );
  AND2_X1 U22659 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n19708), .ZN(
        P2_U3186) );
  AND2_X1 U22660 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n19708), .ZN(
        P2_U3187) );
  AND2_X1 U22661 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n19708), .ZN(
        P2_U3188) );
  AND2_X1 U22662 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n19708), .ZN(
        P2_U3189) );
  AND2_X1 U22663 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n19708), .ZN(
        P2_U3190) );
  AND2_X1 U22664 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n19708), .ZN(
        P2_U3191) );
  AND2_X1 U22665 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n19708), .ZN(
        P2_U3192) );
  AND2_X1 U22666 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n19708), .ZN(
        P2_U3193) );
  AND2_X1 U22667 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n19708), .ZN(
        P2_U3194) );
  AND2_X1 U22668 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n19708), .ZN(
        P2_U3195) );
  AND2_X1 U22669 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n19708), .ZN(
        P2_U3196) );
  AND2_X1 U22670 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n19708), .ZN(
        P2_U3197) );
  AND2_X1 U22671 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n19708), .ZN(
        P2_U3198) );
  AND2_X1 U22672 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n19708), .ZN(
        P2_U3199) );
  AND2_X1 U22673 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n19708), .ZN(
        P2_U3200) );
  AND2_X1 U22674 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n19708), .ZN(P2_U3201) );
  AND2_X1 U22675 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n19708), .ZN(P2_U3202) );
  AND2_X1 U22676 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n19708), .ZN(P2_U3203) );
  AND2_X1 U22677 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n19708), .ZN(P2_U3204) );
  AND2_X1 U22678 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n19708), .ZN(P2_U3205) );
  AND2_X1 U22679 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n19708), .ZN(P2_U3206) );
  AND2_X1 U22680 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n19708), .ZN(P2_U3207) );
  AND2_X1 U22681 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n19708), .ZN(P2_U3208) );
  NOR2_X1 U22682 ( .A1(n19718), .A2(n19835), .ZN(n19716) );
  INV_X1 U22683 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n19854) );
  OR3_X1 U22684 ( .A1(n19716), .A2(n19854), .A3(n19709), .ZN(n19711) );
  INV_X2 U22685 ( .A(n19856), .ZN(n19773) );
  AOI211_X1 U22686 ( .C1(n20703), .C2(P2_REQUESTPENDING_REG_SCAN_IN), .A(
        n19717), .B(n19773), .ZN(n19710) );
  NOR3_X1 U22687 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_0__SCAN_IN), 
        .A3(n20690), .ZN(n19722) );
  AOI211_X1 U22688 ( .C1(n19725), .C2(n19711), .A(n19710), .B(n19722), .ZN(
        n19712) );
  INV_X1 U22689 ( .A(n19712), .ZN(P2_U3209) );
  AOI21_X1 U22690 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n20703), .A(n19725), 
        .ZN(n19719) );
  NOR3_X1 U22691 ( .A1(n19719), .A2(n19854), .A3(n19709), .ZN(n19713) );
  NOR2_X1 U22692 ( .A1(n19713), .A2(n19716), .ZN(n19714) );
  OAI211_X1 U22693 ( .C1(n20703), .C2(n19715), .A(n19714), .B(n19847), .ZN(
        P2_U3210) );
  AOI22_X1 U22694 ( .A1(n19717), .A2(n19854), .B1(n19716), .B2(n20690), .ZN(
        n19724) );
  OAI21_X1 U22695 ( .B1(P2_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .ZN(n19723) );
  NOR2_X1 U22696 ( .A1(n19725), .A2(n19718), .ZN(n19720) );
  AOI21_X1 U22697 ( .B1(n19844), .B2(n19720), .A(n19719), .ZN(n19721) );
  OAI22_X1 U22698 ( .A1(n19724), .A2(n19723), .B1(n19722), .B2(n19721), .ZN(
        P2_U3211) );
  NAND2_X1 U22699 ( .A1(n19773), .A2(n19725), .ZN(n19776) );
  OAI222_X1 U22700 ( .A1(n19771), .A2(n10543), .B1(n19726), .B2(n19773), .C1(
        n10566), .C2(n19770), .ZN(P2_U3212) );
  OAI222_X1 U22701 ( .A1(n19771), .A2(n10566), .B1(n19727), .B2(n19773), .C1(
        n19728), .C2(n19770), .ZN(P2_U3213) );
  OAI222_X1 U22702 ( .A1(n19770), .A2(n19729), .B1(n20933), .B2(n19773), .C1(
        n19728), .C2(n19771), .ZN(P2_U3214) );
  OAI222_X1 U22703 ( .A1(n19776), .A2(n13900), .B1(n19730), .B2(n19773), .C1(
        n19729), .C2(n19771), .ZN(P2_U3215) );
  OAI222_X1 U22704 ( .A1(n19776), .A2(n19732), .B1(n19731), .B2(n19773), .C1(
        n13900), .C2(n19771), .ZN(P2_U3216) );
  OAI222_X1 U22705 ( .A1(n19776), .A2(n19733), .B1(n21025), .B2(n19773), .C1(
        n19732), .C2(n19771), .ZN(P2_U3217) );
  OAI222_X1 U22706 ( .A1(n19776), .A2(n14607), .B1(n19734), .B2(n19773), .C1(
        n19733), .C2(n19771), .ZN(P2_U3218) );
  OAI222_X1 U22707 ( .A1(n19776), .A2(n19736), .B1(n19735), .B2(n19773), .C1(
        n14607), .C2(n19771), .ZN(P2_U3219) );
  OAI222_X1 U22708 ( .A1(n19776), .A2(n18926), .B1(n19737), .B2(n19773), .C1(
        n19736), .C2(n19771), .ZN(P2_U3220) );
  OAI222_X1 U22709 ( .A1(n19770), .A2(n15087), .B1(n19738), .B2(n19773), .C1(
        n18926), .C2(n19771), .ZN(P2_U3221) );
  INV_X1 U22710 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n19740) );
  OAI222_X1 U22711 ( .A1(n19770), .A2(n19740), .B1(n19739), .B2(n19773), .C1(
        n15087), .C2(n19771), .ZN(P2_U3222) );
  OAI222_X1 U22712 ( .A1(n19770), .A2(n10995), .B1(n20990), .B2(n19773), .C1(
        n19740), .C2(n19771), .ZN(P2_U3223) );
  INV_X1 U22713 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n19742) );
  OAI222_X1 U22714 ( .A1(n19770), .A2(n19742), .B1(n19741), .B2(n19773), .C1(
        n10995), .C2(n19771), .ZN(P2_U3224) );
  OAI222_X1 U22715 ( .A1(n19770), .A2(n19744), .B1(n19743), .B2(n19773), .C1(
        n19742), .C2(n19771), .ZN(P2_U3225) );
  OAI222_X1 U22716 ( .A1(n19770), .A2(n19746), .B1(n19745), .B2(n19773), .C1(
        n19744), .C2(n19771), .ZN(P2_U3226) );
  OAI222_X1 U22717 ( .A1(n19770), .A2(n19748), .B1(n19747), .B2(n19773), .C1(
        n19746), .C2(n19771), .ZN(P2_U3227) );
  OAI222_X1 U22718 ( .A1(n19776), .A2(n12180), .B1(n19749), .B2(n19773), .C1(
        n19748), .C2(n19771), .ZN(P2_U3228) );
  OAI222_X1 U22719 ( .A1(n19776), .A2(n21044), .B1(n19750), .B2(n19773), .C1(
        n12180), .C2(n19771), .ZN(P2_U3229) );
  OAI222_X1 U22720 ( .A1(n19776), .A2(n15020), .B1(n19751), .B2(n19773), .C1(
        n21044), .C2(n19771), .ZN(P2_U3230) );
  OAI222_X1 U22721 ( .A1(n19776), .A2(n19753), .B1(n19752), .B2(n19773), .C1(
        n15020), .C2(n19771), .ZN(P2_U3231) );
  OAI222_X1 U22722 ( .A1(n19770), .A2(n12191), .B1(n19754), .B2(n19773), .C1(
        n19753), .C2(n19771), .ZN(P2_U3232) );
  OAI222_X1 U22723 ( .A1(n19770), .A2(n19756), .B1(n19755), .B2(n19773), .C1(
        n12191), .C2(n19771), .ZN(P2_U3233) );
  INV_X1 U22724 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n19758) );
  OAI222_X1 U22725 ( .A1(n19770), .A2(n19758), .B1(n19757), .B2(n19773), .C1(
        n19756), .C2(n19771), .ZN(P2_U3234) );
  OAI222_X1 U22726 ( .A1(n19770), .A2(n19760), .B1(n19759), .B2(n19773), .C1(
        n19758), .C2(n19771), .ZN(P2_U3235) );
  OAI222_X1 U22727 ( .A1(n19770), .A2(n19762), .B1(n19761), .B2(n19773), .C1(
        n19760), .C2(n19771), .ZN(P2_U3236) );
  OAI222_X1 U22728 ( .A1(n19770), .A2(n19765), .B1(n19763), .B2(n19773), .C1(
        n19762), .C2(n19771), .ZN(P2_U3237) );
  INV_X1 U22729 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n19766) );
  OAI222_X1 U22730 ( .A1(n19771), .A2(n19765), .B1(n19764), .B2(n19773), .C1(
        n19766), .C2(n19770), .ZN(P2_U3238) );
  OAI222_X1 U22731 ( .A1(n19770), .A2(n19768), .B1(n19767), .B2(n19773), .C1(
        n19766), .C2(n19771), .ZN(P2_U3239) );
  OAI222_X1 U22732 ( .A1(n19770), .A2(n19772), .B1(n19769), .B2(n19773), .C1(
        n19768), .C2(n19771), .ZN(P2_U3240) );
  OAI222_X1 U22733 ( .A1(n19776), .A2(n19775), .B1(n19774), .B2(n19773), .C1(
        n19772), .C2(n19771), .ZN(P2_U3241) );
  OAI22_X1 U22734 ( .A1(n19856), .A2(P2_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P2_BE_N_REG_3__SCAN_IN), .B2(n19773), .ZN(n19777) );
  INV_X1 U22735 ( .A(n19777), .ZN(P2_U3585) );
  MUX2_X1 U22736 ( .A(P2_BYTEENABLE_REG_2__SCAN_IN), .B(P2_BE_N_REG_2__SCAN_IN), .S(n19856), .Z(P2_U3586) );
  OAI22_X1 U22737 ( .A1(n19856), .A2(P2_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P2_BE_N_REG_1__SCAN_IN), .B2(n19773), .ZN(n19778) );
  INV_X1 U22738 ( .A(n19778), .ZN(P2_U3587) );
  OAI22_X1 U22739 ( .A1(n19856), .A2(P2_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P2_BE_N_REG_0__SCAN_IN), .B2(n19773), .ZN(n19779) );
  INV_X1 U22740 ( .A(n19779), .ZN(P2_U3588) );
  OAI21_X1 U22741 ( .B1(n19783), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n19781), 
        .ZN(n19780) );
  INV_X1 U22742 ( .A(n19780), .ZN(P2_U3591) );
  OAI21_X1 U22743 ( .B1(n19783), .B2(n19782), .A(n19781), .ZN(P2_U3592) );
  INV_X1 U22744 ( .A(n19822), .ZN(n19814) );
  NAND2_X1 U22745 ( .A1(n19807), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19785) );
  AOI21_X1 U22746 ( .B1(n19785), .B2(n19786), .A(n19784), .ZN(n19795) );
  AND2_X1 U22747 ( .A1(n19786), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19809) );
  NAND2_X1 U22748 ( .A1(n19787), .A2(n19809), .ZN(n19798) );
  AOI21_X1 U22749 ( .B1(n19795), .B2(n19798), .A(n19788), .ZN(n19792) );
  OAI22_X1 U22750 ( .A1(n21134), .A2(n19796), .B1(n19790), .B2(n19789), .ZN(
        n19791) );
  NOR2_X1 U22751 ( .A1(n19792), .A2(n19791), .ZN(n19793) );
  AOI22_X1 U22752 ( .A1(n19814), .A2(n19794), .B1(n19793), .B2(n19822), .ZN(
        P2_U3602) );
  INV_X1 U22753 ( .A(n19795), .ZN(n19801) );
  NOR2_X1 U22754 ( .A1(n19797), .A2(n19796), .ZN(n19800) );
  INV_X1 U22755 ( .A(n19798), .ZN(n19799) );
  AOI211_X1 U22756 ( .C1(n19802), .C2(n19801), .A(n19800), .B(n19799), .ZN(
        n19803) );
  AOI22_X1 U22757 ( .A1(n19814), .A2(n19804), .B1(n19803), .B2(n19822), .ZN(
        P2_U3603) );
  INV_X1 U22758 ( .A(n19805), .ZN(n19839) );
  NOR2_X1 U22759 ( .A1(n19839), .A2(n19806), .ZN(n19808) );
  MUX2_X1 U22760 ( .A(n19809), .B(n19808), .S(n19807), .Z(n19810) );
  AOI21_X1 U22761 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19811), .A(n19810), 
        .ZN(n19812) );
  AOI22_X1 U22762 ( .A1(n19814), .A2(n19813), .B1(n19812), .B2(n19822), .ZN(
        P2_U3604) );
  OAI22_X1 U22763 ( .A1(n19817), .A2(n19839), .B1(n19816), .B2(n19815), .ZN(
        n19819) );
  OAI21_X1 U22764 ( .B1(n19819), .B2(n19818), .A(n19822), .ZN(n19820) );
  OAI21_X1 U22765 ( .B1(n19822), .B2(n19821), .A(n19820), .ZN(P2_U3605) );
  INV_X1 U22766 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n19823) );
  AOI22_X1 U22767 ( .A1(n19773), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n19823), 
        .B2(n19856), .ZN(P2_U3608) );
  INV_X1 U22768 ( .A(P2_MORE_REG_SCAN_IN), .ZN(n19834) );
  INV_X1 U22769 ( .A(n19824), .ZN(n19833) );
  INV_X1 U22770 ( .A(n19825), .ZN(n19829) );
  AOI22_X1 U22771 ( .A1(n19829), .A2(n19828), .B1(n19827), .B2(n19826), .ZN(
        n19832) );
  NOR2_X1 U22772 ( .A1(n19833), .A2(n19830), .ZN(n19831) );
  AOI22_X1 U22773 ( .A1(n19834), .A2(n19833), .B1(n19832), .B2(n19831), .ZN(
        P2_U3609) );
  NAND4_X1 U22774 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_STATE2_REG_2__SCAN_IN), .A3(n19836), .A4(n19835), .ZN(n19837) );
  OAI211_X1 U22775 ( .C1(n19840), .C2(n19839), .A(n19838), .B(n19837), .ZN(
        n19855) );
  INV_X1 U22776 ( .A(n19841), .ZN(n19842) );
  NOR2_X1 U22777 ( .A1(n19843), .A2(n19842), .ZN(n19852) );
  NOR2_X1 U22778 ( .A1(n19844), .A2(n19149), .ZN(n19850) );
  OAI211_X1 U22779 ( .C1(n19847), .C2(n19846), .A(n19845), .B(n9776), .ZN(
        n19848) );
  OAI21_X1 U22780 ( .B1(n19850), .B2(n19849), .A(n19848), .ZN(n19851) );
  OAI21_X1 U22781 ( .B1(n19852), .B2(n19851), .A(n19855), .ZN(n19853) );
  OAI21_X1 U22782 ( .B1(n19855), .B2(n19854), .A(n19853), .ZN(P2_U3610) );
  OAI22_X1 U22783 ( .A1(n19856), .A2(P2_MEMORYFETCH_REG_SCAN_IN), .B1(
        P2_M_IO_N_REG_SCAN_IN), .B2(n19773), .ZN(n19857) );
  INV_X1 U22784 ( .A(n19857), .ZN(P2_U3611) );
  AOI21_X1 U22785 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n19858), .A(n20698), 
        .ZN(n20701) );
  INV_X1 U22786 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n19859) );
  NAND2_X1 U22787 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n20698), .ZN(n20740) );
  AOI21_X1 U22788 ( .B1(n20701), .B2(n19859), .A(n20796), .ZN(P1_U2802) );
  INV_X1 U22789 ( .A(n19860), .ZN(n19862) );
  OAI21_X1 U22790 ( .B1(n19862), .B2(n19861), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n19863) );
  OAI21_X1 U22791 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n19864), .A(n19863), 
        .ZN(P1_U2803) );
  INV_X1 U22792 ( .A(n20796), .ZN(n20783) );
  NOR2_X1 U22793 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n19866) );
  OAI21_X1 U22794 ( .B1(n19866), .B2(P1_D_C_N_REG_SCAN_IN), .A(n20740), .ZN(
        n19865) );
  OAI21_X1 U22795 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n20783), .A(n19865), 
        .ZN(P1_U2804) );
  NOR2_X1 U22796 ( .A1(n20796), .A2(n20701), .ZN(n20757) );
  OAI21_X1 U22797 ( .B1(BS16), .B2(n19866), .A(n20757), .ZN(n20755) );
  OAI21_X1 U22798 ( .B1(n20757), .B2(n20574), .A(n20755), .ZN(P1_U2805) );
  OAI21_X1 U22799 ( .B1(n19869), .B2(n19868), .A(n19867), .ZN(P1_U2806) );
  NOR4_X1 U22800 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_21__SCAN_IN), .A3(P1_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_23__SCAN_IN), .ZN(n19873) );
  NOR4_X1 U22801 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_16__SCAN_IN), .A3(P1_DATAWIDTH_REG_17__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_18__SCAN_IN), .ZN(n19872) );
  NOR4_X1 U22802 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A3(P1_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n19871) );
  NOR4_X1 U22803 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_25__SCAN_IN), .A3(P1_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_27__SCAN_IN), .ZN(n19870) );
  NAND4_X1 U22804 ( .A1(n19873), .A2(n19872), .A3(n19871), .A4(n19870), .ZN(
        n19879) );
  NOR4_X1 U22805 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_2__SCAN_IN), .A3(P1_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_4__SCAN_IN), .ZN(n19877) );
  AOI211_X1 U22806 ( .C1(P1_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_20__SCAN_IN), .B(
        P1_DATAWIDTH_REG_8__SCAN_IN), .ZN(n19876) );
  NOR4_X1 U22807 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_11__SCAN_IN), .A3(P1_DATAWIDTH_REG_12__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_14__SCAN_IN), .ZN(n19875) );
  NOR4_X1 U22808 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_6__SCAN_IN), .A3(P1_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_9__SCAN_IN), .ZN(n19874) );
  NAND4_X1 U22809 ( .A1(n19877), .A2(n19876), .A3(n19875), .A4(n19874), .ZN(
        n19878) );
  NOR2_X1 U22810 ( .A1(n19879), .A2(n19878), .ZN(n20778) );
  INV_X1 U22811 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19881) );
  NOR3_X1 U22812 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n19882) );
  OAI21_X1 U22813 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n19882), .A(n20778), .ZN(
        n19880) );
  OAI21_X1 U22814 ( .B1(n20778), .B2(n19881), .A(n19880), .ZN(P1_U2807) );
  INV_X1 U22815 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20756) );
  AOI21_X1 U22816 ( .B1(n13748), .B2(n20756), .A(n19882), .ZN(n19884) );
  INV_X1 U22817 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n19883) );
  INV_X1 U22818 ( .A(n20778), .ZN(n20781) );
  AOI22_X1 U22819 ( .A1(n20778), .A2(n19884), .B1(n19883), .B2(n20781), .ZN(
        P1_U2808) );
  NAND2_X1 U22820 ( .A1(n19950), .A2(n19885), .ZN(n19887) );
  AOI22_X1 U22821 ( .A1(n19948), .A2(n19958), .B1(n19937), .B2(
        P1_EBX_REG_9__SCAN_IN), .ZN(n19886) );
  OAI21_X1 U22822 ( .B1(P1_REIP_REG_9__SCAN_IN), .B2(n19887), .A(n19886), .ZN(
        n19888) );
  AOI211_X1 U22823 ( .C1(n19940), .C2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n19909), .B(n19888), .ZN(n19893) );
  INV_X1 U22824 ( .A(n19889), .ZN(n19959) );
  AOI22_X1 U22825 ( .A1(n19959), .A2(n19912), .B1(n19891), .B2(n19890), .ZN(
        n19892) );
  OAI211_X1 U22826 ( .C1(n19894), .C2(n13939), .A(n19893), .B(n19892), .ZN(
        P1_U2831) );
  NAND2_X1 U22827 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .ZN(n19896) );
  AOI221_X1 U22828 ( .B1(n19923), .B2(n19950), .C1(n19896), .C2(n19950), .A(
        n19895), .ZN(n19911) );
  INV_X1 U22829 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n19908) );
  NAND4_X1 U22830 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .A3(n19922), .A4(n19908), .ZN(n19903) );
  OAI22_X1 U22831 ( .A1(n19900), .A2(n19899), .B1(n19898), .B2(n19897), .ZN(
        n19901) );
  AOI211_X1 U22832 ( .C1(n19940), .C2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n19909), .B(n19901), .ZN(n19902) );
  OAI211_X1 U22833 ( .C1(n19904), .C2(n19957), .A(n19903), .B(n19902), .ZN(
        n19905) );
  AOI21_X1 U22834 ( .B1(n19906), .B2(n19912), .A(n19905), .ZN(n19907) );
  OAI21_X1 U22835 ( .B1(n19911), .B2(n19908), .A(n19907), .ZN(P1_U2833) );
  AOI21_X1 U22836 ( .B1(n19940), .B2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n19909), .ZN(n19921) );
  AOI22_X1 U22837 ( .A1(n19948), .A2(n19910), .B1(n19937), .B2(
        P1_EBX_REG_6__SCAN_IN), .ZN(n19920) );
  INV_X1 U22838 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n20886) );
  OR2_X1 U22839 ( .A1(n19911), .A2(n20886), .ZN(n19915) );
  NAND2_X1 U22840 ( .A1(n19913), .A2(n19912), .ZN(n19914) );
  OAI211_X1 U22841 ( .C1(n19916), .C2(n19957), .A(n19915), .B(n19914), .ZN(
        n19917) );
  INV_X1 U22842 ( .A(n19917), .ZN(n19919) );
  NAND3_X1 U22843 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(n19922), .A3(n20886), 
        .ZN(n19918) );
  NAND4_X1 U22844 ( .A1(n19921), .A2(n19920), .A3(n19919), .A4(n19918), .ZN(
        P1_U2834) );
  INV_X1 U22845 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n20712) );
  AOI22_X1 U22846 ( .A1(n19922), .A2(n20712), .B1(n19937), .B2(
        P1_EBX_REG_5__SCAN_IN), .ZN(n19935) );
  INV_X1 U22847 ( .A(n19923), .ZN(n19925) );
  OAI21_X1 U22848 ( .B1(n19926), .B2(n19925), .A(n19924), .ZN(n19945) );
  NAND2_X1 U22849 ( .A1(n19948), .A2(n19961), .ZN(n19928) );
  NAND2_X1 U22850 ( .A1(n19940), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n19927) );
  NAND3_X1 U22851 ( .A1(n19928), .A2(n19942), .A3(n19927), .ZN(n19929) );
  AOI21_X1 U22852 ( .B1(P1_REIP_REG_5__SCAN_IN), .B2(n19945), .A(n19929), .ZN(
        n19930) );
  OAI21_X1 U22853 ( .B1(n19932), .B2(n19931), .A(n19930), .ZN(n19933) );
  INV_X1 U22854 ( .A(n19933), .ZN(n19934) );
  OAI211_X1 U22855 ( .C1(n19936), .C2(n19957), .A(n19935), .B(n19934), .ZN(
        P1_U2835) );
  NAND2_X1 U22856 ( .A1(n19937), .A2(P1_EBX_REG_4__SCAN_IN), .ZN(n19944) );
  NAND2_X1 U22857 ( .A1(n19939), .A2(n19938), .ZN(n19943) );
  NAND2_X1 U22858 ( .A1(n19940), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n19941) );
  AND4_X1 U22859 ( .A1(n19944), .A2(n19943), .A3(n19942), .A4(n19941), .ZN(
        n19956) );
  NAND2_X1 U22860 ( .A1(n19945), .A2(P1_REIP_REG_4__SCAN_IN), .ZN(n19952) );
  NAND3_X1 U22861 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(P1_REIP_REG_1__SCAN_IN), 
        .A3(P1_REIP_REG_2__SCAN_IN), .ZN(n19946) );
  NOR2_X1 U22862 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(n19946), .ZN(n19949) );
  INV_X1 U22863 ( .A(n20056), .ZN(n19947) );
  AOI22_X1 U22864 ( .A1(n19950), .A2(n19949), .B1(n19948), .B2(n19947), .ZN(
        n19951) );
  NAND2_X1 U22865 ( .A1(n19952), .A2(n19951), .ZN(n19953) );
  AOI21_X1 U22866 ( .B1(n20037), .B2(n19954), .A(n19953), .ZN(n19955) );
  OAI211_X1 U22867 ( .C1(n20042), .C2(n19957), .A(n19956), .B(n19955), .ZN(
        P1_U2836) );
  INV_X1 U22868 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n21074) );
  AOI22_X1 U22869 ( .A1(n19959), .A2(n13156), .B1(n19962), .B2(n19958), .ZN(
        n19960) );
  OAI21_X1 U22870 ( .B1(n19966), .B2(n21074), .A(n19960), .ZN(P1_U2863) );
  INV_X1 U22871 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n19965) );
  AOI22_X1 U22872 ( .A1(n19963), .A2(n13156), .B1(n19962), .B2(n19961), .ZN(
        n19964) );
  OAI21_X1 U22873 ( .B1(n19966), .B2(n19965), .A(n19964), .ZN(P1_U2867) );
  INV_X1 U22874 ( .A(n19967), .ZN(n19968) );
  AOI22_X1 U22875 ( .A1(n19968), .A2(P1_EAX_REG_27__SCAN_IN), .B1(n19993), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n19969) );
  OAI21_X1 U22876 ( .B1(n20997), .B2(n19970), .A(n19969), .ZN(P1_U2909) );
  AOI22_X1 U22877 ( .A1(P1_LWORD_REG_15__SCAN_IN), .A2(n19994), .B1(n19993), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n19971) );
  OAI21_X1 U22878 ( .B1(n13534), .B2(n19996), .A(n19971), .ZN(P1_U2921) );
  AOI22_X1 U22879 ( .A1(P1_LWORD_REG_14__SCAN_IN), .A2(n19994), .B1(n19993), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n19972) );
  OAI21_X1 U22880 ( .B1(n14291), .B2(n19996), .A(n19972), .ZN(P1_U2922) );
  AOI22_X1 U22881 ( .A1(P1_LWORD_REG_13__SCAN_IN), .A2(n19994), .B1(n19993), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n19973) );
  OAI21_X1 U22882 ( .B1(n14293), .B2(n19996), .A(n19973), .ZN(P1_U2923) );
  AOI22_X1 U22883 ( .A1(P1_LWORD_REG_12__SCAN_IN), .A2(n19994), .B1(n19993), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n19974) );
  OAI21_X1 U22884 ( .B1(n14295), .B2(n19996), .A(n19974), .ZN(P1_U2924) );
  INV_X1 U22885 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n19976) );
  AOI22_X1 U22886 ( .A1(P1_LWORD_REG_11__SCAN_IN), .A2(n19994), .B1(n19993), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n19975) );
  OAI21_X1 U22887 ( .B1(n19976), .B2(n19996), .A(n19975), .ZN(P1_U2925) );
  AOI22_X1 U22888 ( .A1(P1_LWORD_REG_10__SCAN_IN), .A2(n19994), .B1(n19993), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n19977) );
  OAI21_X1 U22889 ( .B1(n13934), .B2(n19996), .A(n19977), .ZN(P1_U2926) );
  AOI22_X1 U22890 ( .A1(P1_LWORD_REG_9__SCAN_IN), .A2(n19994), .B1(n19993), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n19978) );
  OAI21_X1 U22891 ( .B1(n13922), .B2(n19996), .A(n19978), .ZN(P1_U2927) );
  AOI22_X1 U22892 ( .A1(P1_LWORD_REG_8__SCAN_IN), .A2(n19994), .B1(n19993), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n19979) );
  OAI21_X1 U22893 ( .B1(n13908), .B2(n19996), .A(n19979), .ZN(P1_U2928) );
  AOI22_X1 U22894 ( .A1(P1_LWORD_REG_7__SCAN_IN), .A2(n19994), .B1(n19993), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n19980) );
  OAI21_X1 U22895 ( .B1(n19981), .B2(n19996), .A(n19980), .ZN(P1_U2929) );
  AOI22_X1 U22896 ( .A1(P1_LWORD_REG_6__SCAN_IN), .A2(n19994), .B1(n19993), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n19982) );
  OAI21_X1 U22897 ( .B1(n19983), .B2(n19996), .A(n19982), .ZN(P1_U2930) );
  AOI22_X1 U22898 ( .A1(P1_LWORD_REG_5__SCAN_IN), .A2(n19994), .B1(n19993), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n19984) );
  OAI21_X1 U22899 ( .B1(n13759), .B2(n19996), .A(n19984), .ZN(P1_U2931) );
  AOI22_X1 U22900 ( .A1(P1_LWORD_REG_4__SCAN_IN), .A2(n19994), .B1(n19993), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n19985) );
  OAI21_X1 U22901 ( .B1(n19986), .B2(n19996), .A(n19985), .ZN(P1_U2932) );
  AOI22_X1 U22902 ( .A1(P1_LWORD_REG_3__SCAN_IN), .A2(n19994), .B1(n19993), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n19987) );
  OAI21_X1 U22903 ( .B1(n19988), .B2(n19996), .A(n19987), .ZN(P1_U2933) );
  AOI22_X1 U22904 ( .A1(P1_LWORD_REG_2__SCAN_IN), .A2(n19994), .B1(n19993), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n19989) );
  OAI21_X1 U22905 ( .B1(n19990), .B2(n19996), .A(n19989), .ZN(P1_U2934) );
  AOI22_X1 U22906 ( .A1(P1_LWORD_REG_1__SCAN_IN), .A2(n19994), .B1(n19993), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n19991) );
  OAI21_X1 U22907 ( .B1(n19992), .B2(n19996), .A(n19991), .ZN(P1_U2935) );
  AOI22_X1 U22908 ( .A1(P1_LWORD_REG_0__SCAN_IN), .A2(n19994), .B1(n19993), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n19995) );
  OAI21_X1 U22909 ( .B1(n19997), .B2(n19996), .A(n19995), .ZN(P1_U2936) );
  AOI22_X1 U22910 ( .A1(n9778), .A2(P1_EAX_REG_24__SCAN_IN), .B1(
        P1_UWORD_REG_8__SCAN_IN), .B2(n20030), .ZN(n20000) );
  INV_X1 U22911 ( .A(n19998), .ZN(n19999) );
  NAND2_X1 U22912 ( .A1(n20015), .A2(n19999), .ZN(n20017) );
  NAND2_X1 U22913 ( .A1(n20000), .A2(n20017), .ZN(P1_U2945) );
  AOI22_X1 U22914 ( .A1(n9778), .A2(P1_EAX_REG_25__SCAN_IN), .B1(
        P1_UWORD_REG_9__SCAN_IN), .B2(n20030), .ZN(n20003) );
  INV_X1 U22915 ( .A(n20001), .ZN(n20002) );
  NAND2_X1 U22916 ( .A1(n20015), .A2(n20002), .ZN(n20019) );
  NAND2_X1 U22917 ( .A1(n20003), .A2(n20019), .ZN(P1_U2946) );
  AOI22_X1 U22918 ( .A1(n9778), .A2(P1_EAX_REG_26__SCAN_IN), .B1(
        P1_UWORD_REG_10__SCAN_IN), .B2(n20025), .ZN(n20006) );
  INV_X1 U22919 ( .A(n20004), .ZN(n20005) );
  NAND2_X1 U22920 ( .A1(n20015), .A2(n20005), .ZN(n20021) );
  NAND2_X1 U22921 ( .A1(n20006), .A2(n20021), .ZN(P1_U2947) );
  AOI22_X1 U22922 ( .A1(n9778), .A2(P1_EAX_REG_28__SCAN_IN), .B1(
        P1_UWORD_REG_12__SCAN_IN), .B2(n20025), .ZN(n20009) );
  INV_X1 U22923 ( .A(n20007), .ZN(n20008) );
  NAND2_X1 U22924 ( .A1(n20015), .A2(n20008), .ZN(n20026) );
  NAND2_X1 U22925 ( .A1(n20009), .A2(n20026), .ZN(P1_U2949) );
  AOI22_X1 U22926 ( .A1(n9778), .A2(P1_EAX_REG_29__SCAN_IN), .B1(
        P1_UWORD_REG_13__SCAN_IN), .B2(n20030), .ZN(n20012) );
  INV_X1 U22927 ( .A(n20010), .ZN(n20011) );
  NAND2_X1 U22928 ( .A1(n20015), .A2(n20011), .ZN(n20028) );
  NAND2_X1 U22929 ( .A1(n20012), .A2(n20028), .ZN(P1_U2950) );
  AOI22_X1 U22930 ( .A1(n9778), .A2(P1_EAX_REG_30__SCAN_IN), .B1(
        P1_UWORD_REG_14__SCAN_IN), .B2(n20030), .ZN(n20016) );
  INV_X1 U22931 ( .A(n20013), .ZN(n20014) );
  NAND2_X1 U22932 ( .A1(n20015), .A2(n20014), .ZN(n20031) );
  NAND2_X1 U22933 ( .A1(n20016), .A2(n20031), .ZN(P1_U2951) );
  AOI22_X1 U22934 ( .A1(n9778), .A2(P1_EAX_REG_8__SCAN_IN), .B1(
        P1_LWORD_REG_8__SCAN_IN), .B2(n20025), .ZN(n20018) );
  NAND2_X1 U22935 ( .A1(n20018), .A2(n20017), .ZN(P1_U2960) );
  AOI22_X1 U22936 ( .A1(n9778), .A2(P1_EAX_REG_9__SCAN_IN), .B1(
        P1_LWORD_REG_9__SCAN_IN), .B2(n20030), .ZN(n20020) );
  NAND2_X1 U22937 ( .A1(n20020), .A2(n20019), .ZN(P1_U2961) );
  AOI22_X1 U22938 ( .A1(n9778), .A2(P1_EAX_REG_10__SCAN_IN), .B1(
        P1_LWORD_REG_10__SCAN_IN), .B2(n20025), .ZN(n20022) );
  NAND2_X1 U22939 ( .A1(n20022), .A2(n20021), .ZN(P1_U2962) );
  AOI22_X1 U22940 ( .A1(n9778), .A2(P1_EAX_REG_11__SCAN_IN), .B1(
        P1_LWORD_REG_11__SCAN_IN), .B2(n20030), .ZN(n20024) );
  NAND2_X1 U22941 ( .A1(n20024), .A2(n20023), .ZN(P1_U2963) );
  AOI22_X1 U22942 ( .A1(n9778), .A2(P1_EAX_REG_12__SCAN_IN), .B1(
        P1_LWORD_REG_12__SCAN_IN), .B2(n20025), .ZN(n20027) );
  NAND2_X1 U22943 ( .A1(n20027), .A2(n20026), .ZN(P1_U2964) );
  AOI22_X1 U22944 ( .A1(n9778), .A2(P1_EAX_REG_13__SCAN_IN), .B1(
        P1_LWORD_REG_13__SCAN_IN), .B2(n20030), .ZN(n20029) );
  NAND2_X1 U22945 ( .A1(n20029), .A2(n20028), .ZN(P1_U2965) );
  AOI22_X1 U22946 ( .A1(n9778), .A2(P1_EAX_REG_14__SCAN_IN), .B1(
        P1_LWORD_REG_14__SCAN_IN), .B2(n20030), .ZN(n20032) );
  NAND2_X1 U22947 ( .A1(n20032), .A2(n20031), .ZN(P1_U2966) );
  AOI22_X1 U22948 ( .A1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n20043), .B1(
        n11744), .B2(P1_REIP_REG_4__SCAN_IN), .ZN(n20040) );
  OAI21_X1 U22949 ( .B1(n20035), .B2(n20034), .A(n20033), .ZN(n20036) );
  INV_X1 U22950 ( .A(n20036), .ZN(n20059) );
  AOI22_X1 U22951 ( .A1(n20059), .A2(n20046), .B1(n20038), .B2(n20037), .ZN(
        n20039) );
  OAI211_X1 U22952 ( .C1(n20042), .C2(n20041), .A(n20040), .B(n20039), .ZN(
        P1_U2995) );
  AOI22_X1 U22953 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n20043), .B1(
        n11744), .B2(P1_REIP_REG_1__SCAN_IN), .ZN(n20049) );
  AOI22_X1 U22954 ( .A1(n20047), .A2(n20046), .B1(n20045), .B2(n20044), .ZN(
        n20048) );
  OAI211_X1 U22955 ( .C1(n20094), .C2(n20050), .A(n20049), .B(n20048), .ZN(
        P1_U2998) );
  INV_X1 U22956 ( .A(n20051), .ZN(n20077) );
  AOI21_X1 U22957 ( .B1(n20053), .B2(n20077), .A(n20052), .ZN(n20070) );
  AOI211_X1 U22958 ( .C1(n20061), .C2(n20069), .A(n20055), .B(n20054), .ZN(
        n20058) );
  INV_X1 U22959 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n20710) );
  OAI22_X1 U22960 ( .A1(n20083), .A2(n20056), .B1(n20710), .B2(n20081), .ZN(
        n20057) );
  AOI211_X1 U22961 ( .C1(n20059), .C2(n20086), .A(n20058), .B(n20057), .ZN(
        n20060) );
  OAI21_X1 U22962 ( .B1(n20070), .B2(n20061), .A(n20060), .ZN(P1_U3027) );
  AOI22_X1 U22963 ( .A1(n11744), .A2(P1_REIP_REG_3__SCAN_IN), .B1(n20063), 
        .B2(n20062), .ZN(n20068) );
  INV_X1 U22964 ( .A(n20064), .ZN(n20066) );
  AOI22_X1 U22965 ( .A1(n20066), .A2(n20086), .B1(n20069), .B2(n20065), .ZN(
        n20067) );
  OAI211_X1 U22966 ( .C1(n20070), .C2(n20069), .A(n20068), .B(n20067), .ZN(
        P1_U3028) );
  NAND2_X1 U22967 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n20071), .ZN(
        n20091) );
  AOI21_X1 U22968 ( .B1(n20075), .B2(n20073), .A(n20072), .ZN(n20089) );
  INV_X1 U22969 ( .A(n20074), .ZN(n20087) );
  NOR2_X1 U22970 ( .A1(n20076), .A2(n20075), .ZN(n20078) );
  AOI21_X1 U22971 ( .B1(n20078), .B2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n20077), .ZN(n20079) );
  NOR2_X1 U22972 ( .A1(n20080), .A2(n20079), .ZN(n20085) );
  INV_X1 U22973 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n20708) );
  OAI22_X1 U22974 ( .A1(n20083), .A2(n20082), .B1(n20708), .B2(n20081), .ZN(
        n20084) );
  AOI211_X1 U22975 ( .C1(n20087), .C2(n20086), .A(n20085), .B(n20084), .ZN(
        n20088) );
  OAI221_X1 U22976 ( .B1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n20091), .C1(
        n20090), .C2(n20089), .A(n20088), .ZN(P1_U3029) );
  NOR2_X1 U22977 ( .A1(n20869), .A2(n20771), .ZN(P1_U3032) );
  NOR2_X2 U22978 ( .A1(n20092), .A2(n20094), .ZN(n20142) );
  NOR2_X2 U22979 ( .A1(n20094), .A2(n20093), .ZN(n20141) );
  AOI22_X1 U22980 ( .A1(DATAI_16_), .A2(n20142), .B1(BUF1_REG_16__SCAN_IN), 
        .B2(n20141), .ZN(n20585) );
  INV_X1 U22981 ( .A(n20179), .ZN(n20095) );
  NAND2_X1 U22982 ( .A1(n14544), .A2(n20252), .ZN(n20629) );
  INV_X1 U22983 ( .A(n20450), .ZN(n20096) );
  AOI22_X1 U22984 ( .A1(DATAI_24_), .A2(n20142), .B1(BUF1_REG_24__SCAN_IN), 
        .B2(n20141), .ZN(n20638) );
  NAND2_X1 U22985 ( .A1(n20143), .A2(n9822), .ZN(n20486) );
  NAND2_X1 U22986 ( .A1(n20367), .A2(n20773), .ZN(n20180) );
  OR2_X1 U22987 ( .A1(n20485), .A2(n20180), .ZN(n20144) );
  OAI22_X1 U22988 ( .A1(n20634), .A2(n20638), .B1(n20486), .B2(n20144), .ZN(
        n20099) );
  INV_X1 U22989 ( .A(n20099), .ZN(n20112) );
  INV_X1 U22990 ( .A(n20144), .ZN(n20105) );
  INV_X1 U22991 ( .A(n20108), .ZN(n20100) );
  NOR2_X1 U22992 ( .A1(n20100), .A2(n20623), .ZN(n20484) );
  NAND3_X1 U22993 ( .A1(n20172), .A2(n20765), .A3(n20634), .ZN(n20101) );
  NAND2_X1 U22994 ( .A1(n20574), .A2(n20765), .ZN(n20480) );
  NAND2_X1 U22995 ( .A1(n20101), .A2(n20480), .ZN(n20107) );
  NAND2_X1 U22996 ( .A1(n9890), .A2(n13609), .ZN(n20109) );
  INV_X1 U22997 ( .A(n20103), .ZN(n20369) );
  NAND2_X1 U22998 ( .A1(n20369), .A2(n20421), .ZN(n20256) );
  AOI22_X1 U22999 ( .A1(n20107), .A2(n20109), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20256), .ZN(n20104) );
  NOR2_X2 U23000 ( .A1(n20106), .A2(n20259), .ZN(n20625) );
  INV_X1 U23001 ( .A(n20107), .ZN(n20110) );
  OR2_X1 U23002 ( .A1(n20108), .A2(n20623), .ZN(n20370) );
  AOI22_X1 U23003 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n20148), .B1(
        n20625), .B2(n20147), .ZN(n20111) );
  OAI211_X1 U23004 ( .C1(n20585), .C2(n20172), .A(n20112), .B(n20111), .ZN(
        P1_U3033) );
  AOI22_X1 U23005 ( .A1(DATAI_17_), .A2(n20142), .B1(BUF1_REG_17__SCAN_IN), 
        .B2(n20141), .ZN(n20589) );
  AOI22_X1 U23006 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n20141), .B1(DATAI_25_), 
        .B2(n20142), .ZN(n20644) );
  NAND2_X1 U23007 ( .A1(n20143), .A2(n20113), .ZN(n20499) );
  OAI22_X1 U23008 ( .A1(n20634), .A2(n20644), .B1(n20499), .B2(n20144), .ZN(
        n20114) );
  INV_X1 U23009 ( .A(n20114), .ZN(n20117) );
  NOR2_X2 U23010 ( .A1(n20115), .A2(n20259), .ZN(n20639) );
  AOI22_X1 U23011 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20148), .B1(
        n20639), .B2(n20147), .ZN(n20116) );
  OAI211_X1 U23012 ( .C1(n20589), .C2(n20172), .A(n20117), .B(n20116), .ZN(
        P1_U3034) );
  AOI22_X1 U23013 ( .A1(DATAI_18_), .A2(n20142), .B1(BUF1_REG_18__SCAN_IN), 
        .B2(n20141), .ZN(n20593) );
  AOI22_X1 U23014 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n20141), .B1(DATAI_26_), 
        .B2(n20142), .ZN(n20650) );
  NAND2_X1 U23015 ( .A1(n20143), .A2(n11267), .ZN(n20504) );
  OAI22_X1 U23016 ( .A1(n20634), .A2(n20650), .B1(n20504), .B2(n20144), .ZN(
        n20118) );
  INV_X1 U23017 ( .A(n20118), .ZN(n20121) );
  NOR2_X2 U23018 ( .A1(n20119), .A2(n20259), .ZN(n20645) );
  AOI22_X1 U23019 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20148), .B1(
        n20645), .B2(n20147), .ZN(n20120) );
  OAI211_X1 U23020 ( .C1(n20593), .C2(n20172), .A(n20121), .B(n20120), .ZN(
        P1_U3035) );
  AOI22_X1 U23021 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n20141), .B1(DATAI_19_), 
        .B2(n20142), .ZN(n20597) );
  AOI22_X1 U23022 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n20141), .B1(DATAI_27_), 
        .B2(n20142), .ZN(n20656) );
  NAND2_X1 U23023 ( .A1(n20143), .A2(n20122), .ZN(n20509) );
  OAI22_X1 U23024 ( .A1(n20634), .A2(n20656), .B1(n20509), .B2(n20144), .ZN(
        n20123) );
  INV_X1 U23025 ( .A(n20123), .ZN(n20126) );
  NOR2_X2 U23026 ( .A1(n20124), .A2(n20259), .ZN(n20651) );
  AOI22_X1 U23027 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20148), .B1(
        n20651), .B2(n20147), .ZN(n20125) );
  OAI211_X1 U23028 ( .C1(n20597), .C2(n20172), .A(n20126), .B(n20125), .ZN(
        P1_U3036) );
  AOI22_X1 U23029 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n20141), .B1(DATAI_20_), 
        .B2(n20142), .ZN(n20601) );
  AOI22_X1 U23030 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n20141), .B1(DATAI_28_), 
        .B2(n20142), .ZN(n20662) );
  NAND2_X1 U23031 ( .A1(n20143), .A2(n20127), .ZN(n20514) );
  OAI22_X1 U23032 ( .A1(n20634), .A2(n20662), .B1(n20514), .B2(n20144), .ZN(
        n20128) );
  INV_X1 U23033 ( .A(n20128), .ZN(n20131) );
  NOR2_X2 U23034 ( .A1(n20129), .A2(n20259), .ZN(n20657) );
  AOI22_X1 U23035 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20148), .B1(
        n20657), .B2(n20147), .ZN(n20130) );
  OAI211_X1 U23036 ( .C1(n20601), .C2(n20172), .A(n20131), .B(n20130), .ZN(
        P1_U3037) );
  AOI22_X1 U23037 ( .A1(DATAI_21_), .A2(n20142), .B1(BUF1_REG_21__SCAN_IN), 
        .B2(n20141), .ZN(n20605) );
  AOI22_X1 U23038 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n20141), .B1(DATAI_29_), 
        .B2(n20142), .ZN(n20668) );
  NAND2_X1 U23039 ( .A1(n20143), .A2(n11251), .ZN(n20519) );
  OAI22_X1 U23040 ( .A1(n20634), .A2(n20668), .B1(n20519), .B2(n20144), .ZN(
        n20132) );
  INV_X1 U23041 ( .A(n20132), .ZN(n20135) );
  NOR2_X2 U23042 ( .A1(n20133), .A2(n20259), .ZN(n20663) );
  AOI22_X1 U23043 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20148), .B1(
        n20663), .B2(n20147), .ZN(n20134) );
  OAI211_X1 U23044 ( .C1(n20605), .C2(n20172), .A(n20135), .B(n20134), .ZN(
        P1_U3038) );
  AOI22_X1 U23045 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n20141), .B1(DATAI_22_), 
        .B2(n20142), .ZN(n20609) );
  AOI22_X1 U23046 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n20141), .B1(DATAI_30_), 
        .B2(n20142), .ZN(n20674) );
  NAND2_X1 U23047 ( .A1(n20143), .A2(n20136), .ZN(n20524) );
  OAI22_X1 U23048 ( .A1(n20634), .A2(n20674), .B1(n20524), .B2(n20144), .ZN(
        n20137) );
  INV_X1 U23049 ( .A(n20137), .ZN(n20140) );
  NOR2_X2 U23050 ( .A1(n20138), .A2(n20259), .ZN(n20669) );
  AOI22_X1 U23051 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20148), .B1(
        n20669), .B2(n20147), .ZN(n20139) );
  OAI211_X1 U23052 ( .C1(n20609), .C2(n20172), .A(n20140), .B(n20139), .ZN(
        P1_U3039) );
  AOI22_X1 U23053 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n20141), .B1(DATAI_23_), 
        .B2(n20142), .ZN(n20617) );
  AOI22_X1 U23054 ( .A1(DATAI_31_), .A2(n20142), .B1(BUF1_REG_31__SCAN_IN), 
        .B2(n20141), .ZN(n20685) );
  NAND2_X1 U23055 ( .A1(n20143), .A2(n9790), .ZN(n20530) );
  OAI22_X1 U23056 ( .A1(n20634), .A2(n20685), .B1(n20530), .B2(n20144), .ZN(
        n20145) );
  INV_X1 U23057 ( .A(n20145), .ZN(n20150) );
  NOR2_X2 U23058 ( .A1(n20146), .A2(n20259), .ZN(n20676) );
  AOI22_X1 U23059 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20148), .B1(
        n20676), .B2(n20147), .ZN(n20149) );
  OAI211_X1 U23060 ( .C1(n20617), .C2(n20172), .A(n20150), .B(n20149), .ZN(
        P1_U3040) );
  NOR2_X1 U23061 ( .A1(n20180), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20156) );
  INV_X1 U23062 ( .A(n20156), .ZN(n20152) );
  NOR2_X1 U23063 ( .A1(n20538), .A2(n20152), .ZN(n20174) );
  INV_X1 U23064 ( .A(n20151), .ZN(n20540) );
  AOI21_X1 U23065 ( .B1(n9890), .B2(n20540), .A(n20174), .ZN(n20153) );
  OAI22_X1 U23066 ( .A1(n20153), .A2(n20632), .B1(n20152), .B2(n20623), .ZN(
        n20173) );
  AOI22_X1 U23067 ( .A1(n20626), .A2(n20174), .B1(n20173), .B2(n20625), .ZN(
        n20158) );
  INV_X1 U23068 ( .A(n20219), .ZN(n20154) );
  OAI211_X1 U23069 ( .C1(n20154), .C2(n20574), .A(n20458), .B(n20153), .ZN(
        n20155) );
  OAI211_X1 U23070 ( .C1(n20765), .C2(n20156), .A(n20630), .B(n20155), .ZN(
        n20176) );
  INV_X1 U23071 ( .A(n20638), .ZN(n20582) );
  AOI22_X1 U23072 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20176), .B1(
        n20175), .B2(n20582), .ZN(n20157) );
  OAI211_X1 U23073 ( .C1(n20585), .C2(n20213), .A(n20158), .B(n20157), .ZN(
        P1_U3041) );
  AOI22_X1 U23074 ( .A1(n20640), .A2(n20174), .B1(n20173), .B2(n20639), .ZN(
        n20160) );
  INV_X1 U23075 ( .A(n20644), .ZN(n20586) );
  AOI22_X1 U23076 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20176), .B1(
        n20175), .B2(n20586), .ZN(n20159) );
  OAI211_X1 U23077 ( .C1(n20589), .C2(n20213), .A(n20160), .B(n20159), .ZN(
        P1_U3042) );
  AOI22_X1 U23078 ( .A1(n20646), .A2(n20174), .B1(n20173), .B2(n20645), .ZN(
        n20162) );
  INV_X1 U23079 ( .A(n20650), .ZN(n20590) );
  AOI22_X1 U23080 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20176), .B1(
        n20175), .B2(n20590), .ZN(n20161) );
  OAI211_X1 U23081 ( .C1(n20593), .C2(n20213), .A(n20162), .B(n20161), .ZN(
        P1_U3043) );
  AOI22_X1 U23082 ( .A1(n20652), .A2(n20174), .B1(n20173), .B2(n20651), .ZN(
        n20164) );
  INV_X1 U23083 ( .A(n20656), .ZN(n20594) );
  AOI22_X1 U23084 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20176), .B1(
        n20175), .B2(n20594), .ZN(n20163) );
  OAI211_X1 U23085 ( .C1(n20597), .C2(n20213), .A(n20164), .B(n20163), .ZN(
        P1_U3044) );
  AOI22_X1 U23086 ( .A1(n20658), .A2(n20174), .B1(n20173), .B2(n20657), .ZN(
        n20166) );
  INV_X1 U23087 ( .A(n20662), .ZN(n20598) );
  AOI22_X1 U23088 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20176), .B1(
        n20175), .B2(n20598), .ZN(n20165) );
  OAI211_X1 U23089 ( .C1(n20601), .C2(n20213), .A(n20166), .B(n20165), .ZN(
        P1_U3045) );
  AOI22_X1 U23090 ( .A1(n20664), .A2(n20174), .B1(n20173), .B2(n20663), .ZN(
        n20168) );
  INV_X1 U23091 ( .A(n20668), .ZN(n20602) );
  AOI22_X1 U23092 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20176), .B1(
        n20175), .B2(n20602), .ZN(n20167) );
  OAI211_X1 U23093 ( .C1(n20605), .C2(n20213), .A(n20168), .B(n20167), .ZN(
        P1_U3046) );
  AOI22_X1 U23094 ( .A1(n20670), .A2(n20174), .B1(n20173), .B2(n20669), .ZN(
        n20171) );
  INV_X1 U23095 ( .A(n20213), .ZN(n20169) );
  INV_X1 U23096 ( .A(n20609), .ZN(n20671) );
  AOI22_X1 U23097 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20176), .B1(
        n20169), .B2(n20671), .ZN(n20170) );
  OAI211_X1 U23098 ( .C1(n20674), .C2(n20172), .A(n20171), .B(n20170), .ZN(
        P1_U3047) );
  AOI22_X1 U23099 ( .A1(n20678), .A2(n20174), .B1(n20173), .B2(n20676), .ZN(
        n20178) );
  INV_X1 U23100 ( .A(n20685), .ZN(n20612) );
  AOI22_X1 U23101 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20176), .B1(
        n20175), .B2(n20612), .ZN(n20177) );
  OAI211_X1 U23102 ( .C1(n20617), .C2(n20213), .A(n20178), .B(n20177), .ZN(
        P1_U3048) );
  INV_X1 U23103 ( .A(n20180), .ZN(n20214) );
  NAND2_X1 U23104 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20214), .ZN(
        n20222) );
  OR2_X1 U23105 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20222), .ZN(
        n20207) );
  OAI22_X1 U23106 ( .A1(n20213), .A2(n20638), .B1(n20486), .B2(n20207), .ZN(
        n20181) );
  INV_X1 U23107 ( .A(n20181), .ZN(n20188) );
  NAND2_X1 U23108 ( .A1(n20251), .A2(n20213), .ZN(n20182) );
  AOI21_X1 U23109 ( .B1(n20182), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n20632), 
        .ZN(n20184) );
  NAND2_X1 U23110 ( .A1(n9890), .A2(n20577), .ZN(n20185) );
  AOI22_X1 U23111 ( .A1(n20184), .A2(n20185), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20207), .ZN(n20183) );
  OAI21_X1 U23112 ( .B1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n20421), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n20316) );
  NAND3_X1 U23113 ( .A1(n20429), .A2(n20183), .A3(n20316), .ZN(n20210) );
  INV_X1 U23114 ( .A(n20184), .ZN(n20186) );
  INV_X1 U23115 ( .A(n20421), .ZN(n20368) );
  NAND2_X1 U23116 ( .A1(n20368), .A2(n20773), .ZN(n20309) );
  AOI22_X1 U23117 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20210), .B1(
        n20625), .B2(n20209), .ZN(n20187) );
  OAI211_X1 U23118 ( .C1(n20585), .C2(n20251), .A(n20188), .B(n20187), .ZN(
        P1_U3049) );
  OAI22_X1 U23119 ( .A1(n20213), .A2(n20644), .B1(n20499), .B2(n20207), .ZN(
        n20189) );
  INV_X1 U23120 ( .A(n20189), .ZN(n20191) );
  AOI22_X1 U23121 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20210), .B1(
        n20639), .B2(n20209), .ZN(n20190) );
  OAI211_X1 U23122 ( .C1(n20589), .C2(n20251), .A(n20191), .B(n20190), .ZN(
        P1_U3050) );
  OAI22_X1 U23123 ( .A1(n20213), .A2(n20650), .B1(n20504), .B2(n20207), .ZN(
        n20192) );
  INV_X1 U23124 ( .A(n20192), .ZN(n20194) );
  AOI22_X1 U23125 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20210), .B1(
        n20645), .B2(n20209), .ZN(n20193) );
  OAI211_X1 U23126 ( .C1(n20593), .C2(n20251), .A(n20194), .B(n20193), .ZN(
        P1_U3051) );
  OAI22_X1 U23127 ( .A1(n20251), .A2(n20597), .B1(n20509), .B2(n20207), .ZN(
        n20195) );
  INV_X1 U23128 ( .A(n20195), .ZN(n20197) );
  AOI22_X1 U23129 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20210), .B1(
        n20651), .B2(n20209), .ZN(n20196) );
  OAI211_X1 U23130 ( .C1(n20656), .C2(n20213), .A(n20197), .B(n20196), .ZN(
        P1_U3052) );
  OAI22_X1 U23131 ( .A1(n20213), .A2(n20662), .B1(n20514), .B2(n20207), .ZN(
        n20198) );
  INV_X1 U23132 ( .A(n20198), .ZN(n20200) );
  AOI22_X1 U23133 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20210), .B1(
        n20657), .B2(n20209), .ZN(n20199) );
  OAI211_X1 U23134 ( .C1(n20601), .C2(n20251), .A(n20200), .B(n20199), .ZN(
        P1_U3053) );
  OAI22_X1 U23135 ( .A1(n20251), .A2(n20605), .B1(n20519), .B2(n20207), .ZN(
        n20201) );
  INV_X1 U23136 ( .A(n20201), .ZN(n20203) );
  AOI22_X1 U23137 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20210), .B1(
        n20663), .B2(n20209), .ZN(n20202) );
  OAI211_X1 U23138 ( .C1(n20668), .C2(n20213), .A(n20203), .B(n20202), .ZN(
        P1_U3054) );
  OAI22_X1 U23139 ( .A1(n20251), .A2(n20609), .B1(n20524), .B2(n20207), .ZN(
        n20204) );
  INV_X1 U23140 ( .A(n20204), .ZN(n20206) );
  AOI22_X1 U23141 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20210), .B1(
        n20669), .B2(n20209), .ZN(n20205) );
  OAI211_X1 U23142 ( .C1(n20674), .C2(n20213), .A(n20206), .B(n20205), .ZN(
        P1_U3055) );
  OAI22_X1 U23143 ( .A1(n20251), .A2(n20617), .B1(n20530), .B2(n20207), .ZN(
        n20208) );
  INV_X1 U23144 ( .A(n20208), .ZN(n20212) );
  AOI22_X1 U23145 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20210), .B1(
        n20676), .B2(n20209), .ZN(n20211) );
  OAI211_X1 U23146 ( .C1(n20685), .C2(n20213), .A(n20212), .B(n20211), .ZN(
        P1_U3056) );
  NAND2_X1 U23147 ( .A1(n20215), .A2(n20214), .ZN(n20245) );
  OAI22_X1 U23148 ( .A1(n20251), .A2(n20638), .B1(n20486), .B2(n20245), .ZN(
        n20216) );
  INV_X1 U23149 ( .A(n20216), .ZN(n20226) );
  NOR2_X1 U23150 ( .A1(n20217), .A2(n9801), .ZN(n20619) );
  INV_X1 U23151 ( .A(n20245), .ZN(n20218) );
  AOI21_X1 U23152 ( .B1(n9890), .B2(n20619), .A(n20218), .ZN(n20223) );
  INV_X1 U23153 ( .A(n20628), .ZN(n20764) );
  AOI21_X1 U23154 ( .B1(n20219), .B2(n20764), .A(n20632), .ZN(n20221) );
  AOI22_X1 U23155 ( .A1(n20223), .A2(n20221), .B1(n20632), .B2(n20222), .ZN(
        n20220) );
  NAND2_X1 U23156 ( .A1(n20630), .A2(n20220), .ZN(n20248) );
  INV_X1 U23157 ( .A(n20221), .ZN(n20224) );
  OAI22_X1 U23158 ( .A1(n20224), .A2(n20223), .B1(n20623), .B2(n20222), .ZN(
        n20247) );
  AOI22_X1 U23159 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20248), .B1(
        n20625), .B2(n20247), .ZN(n20225) );
  OAI211_X1 U23160 ( .C1(n20585), .C2(n20281), .A(n20226), .B(n20225), .ZN(
        P1_U3057) );
  OAI22_X1 U23161 ( .A1(n20281), .A2(n20589), .B1(n20499), .B2(n20245), .ZN(
        n20227) );
  INV_X1 U23162 ( .A(n20227), .ZN(n20229) );
  AOI22_X1 U23163 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20248), .B1(
        n20639), .B2(n20247), .ZN(n20228) );
  OAI211_X1 U23164 ( .C1(n20644), .C2(n20251), .A(n20229), .B(n20228), .ZN(
        P1_U3058) );
  OAI22_X1 U23165 ( .A1(n20251), .A2(n20650), .B1(n20504), .B2(n20245), .ZN(
        n20230) );
  INV_X1 U23166 ( .A(n20230), .ZN(n20232) );
  AOI22_X1 U23167 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20248), .B1(
        n20645), .B2(n20247), .ZN(n20231) );
  OAI211_X1 U23168 ( .C1(n20593), .C2(n20281), .A(n20232), .B(n20231), .ZN(
        P1_U3059) );
  OAI22_X1 U23169 ( .A1(n20281), .A2(n20597), .B1(n20509), .B2(n20245), .ZN(
        n20233) );
  INV_X1 U23170 ( .A(n20233), .ZN(n20235) );
  AOI22_X1 U23171 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20248), .B1(
        n20651), .B2(n20247), .ZN(n20234) );
  OAI211_X1 U23172 ( .C1(n20656), .C2(n20251), .A(n20235), .B(n20234), .ZN(
        P1_U3060) );
  OAI22_X1 U23173 ( .A1(n20281), .A2(n20601), .B1(n20514), .B2(n20245), .ZN(
        n20236) );
  INV_X1 U23174 ( .A(n20236), .ZN(n20238) );
  AOI22_X1 U23175 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20248), .B1(
        n20657), .B2(n20247), .ZN(n20237) );
  OAI211_X1 U23176 ( .C1(n20662), .C2(n20251), .A(n20238), .B(n20237), .ZN(
        P1_U3061) );
  OAI22_X1 U23177 ( .A1(n20281), .A2(n20605), .B1(n20519), .B2(n20245), .ZN(
        n20239) );
  INV_X1 U23178 ( .A(n20239), .ZN(n20241) );
  AOI22_X1 U23179 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20248), .B1(
        n20663), .B2(n20247), .ZN(n20240) );
  OAI211_X1 U23180 ( .C1(n20668), .C2(n20251), .A(n20241), .B(n20240), .ZN(
        P1_U3062) );
  OAI22_X1 U23181 ( .A1(n20251), .A2(n20674), .B1(n20524), .B2(n20245), .ZN(
        n20242) );
  INV_X1 U23182 ( .A(n20242), .ZN(n20244) );
  AOI22_X1 U23183 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20248), .B1(
        n20669), .B2(n20247), .ZN(n20243) );
  OAI211_X1 U23184 ( .C1(n20609), .C2(n20281), .A(n20244), .B(n20243), .ZN(
        P1_U3063) );
  OAI22_X1 U23185 ( .A1(n20281), .A2(n20617), .B1(n20530), .B2(n20245), .ZN(
        n20246) );
  INV_X1 U23186 ( .A(n20246), .ZN(n20250) );
  AOI22_X1 U23187 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20248), .B1(
        n20676), .B2(n20247), .ZN(n20249) );
  OAI211_X1 U23188 ( .C1(n20685), .C2(n20251), .A(n20250), .B(n20249), .ZN(
        P1_U3064) );
  INV_X1 U23189 ( .A(n20252), .ZN(n20253) );
  INV_X1 U23190 ( .A(n20484), .ZN(n20573) );
  OR2_X1 U23191 ( .A1(n13438), .A2(n20254), .ZN(n20308) );
  NAND3_X1 U23192 ( .A1(n20339), .A2(n20765), .A3(n13609), .ZN(n20255) );
  OAI21_X1 U23193 ( .B1(n20256), .B2(n20573), .A(n20255), .ZN(n20276) );
  AOI22_X1 U23194 ( .A1(n20626), .A2(n10242), .B1(n20625), .B2(n20276), .ZN(
        n20262) );
  AOI21_X1 U23195 ( .B1(n20281), .B2(n20305), .A(n20574), .ZN(n20257) );
  AOI21_X1 U23196 ( .B1(n20339), .B2(n13609), .A(n20257), .ZN(n20258) );
  NOR2_X1 U23197 ( .A1(n20258), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20260) );
  INV_X1 U23198 ( .A(n20370), .ZN(n20422) );
  INV_X1 U23199 ( .A(n20281), .ZN(n20269) );
  AOI22_X1 U23200 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20278), .B1(
        n20269), .B2(n20582), .ZN(n20261) );
  OAI211_X1 U23201 ( .C1(n20585), .C2(n20305), .A(n20262), .B(n20261), .ZN(
        P1_U3065) );
  AOI22_X1 U23202 ( .A1(n20640), .A2(n10242), .B1(n20639), .B2(n20276), .ZN(
        n20264) );
  AOI22_X1 U23203 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20278), .B1(
        n20269), .B2(n20586), .ZN(n20263) );
  OAI211_X1 U23204 ( .C1(n20589), .C2(n20305), .A(n20264), .B(n20263), .ZN(
        P1_U3066) );
  AOI22_X1 U23205 ( .A1(n20646), .A2(n10242), .B1(n20645), .B2(n20276), .ZN(
        n20266) );
  AOI22_X1 U23206 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20278), .B1(
        n20269), .B2(n20590), .ZN(n20265) );
  OAI211_X1 U23207 ( .C1(n20593), .C2(n20305), .A(n20266), .B(n20265), .ZN(
        P1_U3067) );
  AOI22_X1 U23208 ( .A1(n20652), .A2(n10242), .B1(n20651), .B2(n20276), .ZN(
        n20268) );
  INV_X1 U23209 ( .A(n20305), .ZN(n20277) );
  INV_X1 U23210 ( .A(n20597), .ZN(n20653) );
  AOI22_X1 U23211 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20278), .B1(
        n20277), .B2(n20653), .ZN(n20267) );
  OAI211_X1 U23212 ( .C1(n20656), .C2(n20281), .A(n20268), .B(n20267), .ZN(
        P1_U3068) );
  AOI22_X1 U23213 ( .A1(n20658), .A2(n10242), .B1(n20657), .B2(n20276), .ZN(
        n20271) );
  AOI22_X1 U23214 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20278), .B1(
        n20269), .B2(n20598), .ZN(n20270) );
  OAI211_X1 U23215 ( .C1(n20601), .C2(n20305), .A(n20271), .B(n20270), .ZN(
        P1_U3069) );
  AOI22_X1 U23216 ( .A1(n20664), .A2(n10242), .B1(n20663), .B2(n20276), .ZN(
        n20273) );
  INV_X1 U23217 ( .A(n20605), .ZN(n20665) );
  AOI22_X1 U23218 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20278), .B1(
        n20277), .B2(n20665), .ZN(n20272) );
  OAI211_X1 U23219 ( .C1(n20668), .C2(n20281), .A(n20273), .B(n20272), .ZN(
        P1_U3070) );
  AOI22_X1 U23220 ( .A1(n20670), .A2(n10242), .B1(n20669), .B2(n20276), .ZN(
        n20275) );
  AOI22_X1 U23221 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20278), .B1(
        n20277), .B2(n20671), .ZN(n20274) );
  OAI211_X1 U23222 ( .C1(n20674), .C2(n20281), .A(n20275), .B(n20274), .ZN(
        P1_U3071) );
  AOI22_X1 U23223 ( .A1(n20678), .A2(n10242), .B1(n20676), .B2(n20276), .ZN(
        n20280) );
  INV_X1 U23224 ( .A(n20617), .ZN(n20679) );
  AOI22_X1 U23225 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20278), .B1(
        n20277), .B2(n20679), .ZN(n20279) );
  OAI211_X1 U23226 ( .C1(n20685), .C2(n20281), .A(n20280), .B(n20279), .ZN(
        P1_U3072) );
  NOR2_X1 U23227 ( .A1(n20311), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20285) );
  INV_X1 U23228 ( .A(n20285), .ZN(n20282) );
  NOR2_X1 U23229 ( .A1(n20538), .A2(n20282), .ZN(n20301) );
  AOI21_X1 U23230 ( .B1(n20339), .B2(n20540), .A(n20301), .ZN(n20283) );
  OAI22_X1 U23231 ( .A1(n20283), .A2(n20632), .B1(n20282), .B2(n20623), .ZN(
        n20300) );
  AOI22_X1 U23232 ( .A1(n20626), .A2(n20301), .B1(n20625), .B2(n20300), .ZN(
        n20287) );
  INV_X1 U23233 ( .A(n20766), .ZN(n20342) );
  OAI211_X1 U23234 ( .C1(n20342), .C2(n20574), .A(n20458), .B(n20283), .ZN(
        n20284) );
  OAI211_X1 U23235 ( .C1(n20458), .C2(n20285), .A(n20630), .B(n20284), .ZN(
        n20302) );
  INV_X1 U23236 ( .A(n20585), .ZN(n20635) );
  AOI22_X1 U23237 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20302), .B1(
        n20333), .B2(n20635), .ZN(n20286) );
  OAI211_X1 U23238 ( .C1(n20638), .C2(n20305), .A(n20287), .B(n20286), .ZN(
        P1_U3073) );
  AOI22_X1 U23239 ( .A1(n20640), .A2(n20301), .B1(n20639), .B2(n20300), .ZN(
        n20289) );
  INV_X1 U23240 ( .A(n20589), .ZN(n20641) );
  AOI22_X1 U23241 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20302), .B1(
        n20333), .B2(n20641), .ZN(n20288) );
  OAI211_X1 U23242 ( .C1(n20644), .C2(n20305), .A(n20289), .B(n20288), .ZN(
        P1_U3074) );
  AOI22_X1 U23243 ( .A1(n20646), .A2(n20301), .B1(n20645), .B2(n20300), .ZN(
        n20291) );
  INV_X1 U23244 ( .A(n20593), .ZN(n20647) );
  AOI22_X1 U23245 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20302), .B1(
        n20333), .B2(n20647), .ZN(n20290) );
  OAI211_X1 U23246 ( .C1(n20650), .C2(n20305), .A(n20291), .B(n20290), .ZN(
        P1_U3075) );
  AOI22_X1 U23247 ( .A1(n20652), .A2(n20301), .B1(n20651), .B2(n20300), .ZN(
        n20293) );
  AOI22_X1 U23248 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20302), .B1(
        n20333), .B2(n20653), .ZN(n20292) );
  OAI211_X1 U23249 ( .C1(n20656), .C2(n20305), .A(n20293), .B(n20292), .ZN(
        P1_U3076) );
  AOI22_X1 U23250 ( .A1(n20658), .A2(n20301), .B1(n20657), .B2(n20300), .ZN(
        n20295) );
  INV_X1 U23251 ( .A(n20601), .ZN(n20659) );
  AOI22_X1 U23252 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20302), .B1(
        n20333), .B2(n20659), .ZN(n20294) );
  OAI211_X1 U23253 ( .C1(n20662), .C2(n20305), .A(n20295), .B(n20294), .ZN(
        P1_U3077) );
  AOI22_X1 U23254 ( .A1(n20664), .A2(n20301), .B1(n20663), .B2(n20300), .ZN(
        n20297) );
  AOI22_X1 U23255 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20302), .B1(
        n20333), .B2(n20665), .ZN(n20296) );
  OAI211_X1 U23256 ( .C1(n20668), .C2(n20305), .A(n20297), .B(n20296), .ZN(
        P1_U3078) );
  AOI22_X1 U23257 ( .A1(n20670), .A2(n20301), .B1(n20669), .B2(n20300), .ZN(
        n20299) );
  AOI22_X1 U23258 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20302), .B1(
        n20333), .B2(n20671), .ZN(n20298) );
  OAI211_X1 U23259 ( .C1(n20674), .C2(n20305), .A(n20299), .B(n20298), .ZN(
        P1_U3079) );
  AOI22_X1 U23260 ( .A1(n20678), .A2(n20301), .B1(n20676), .B2(n20300), .ZN(
        n20304) );
  AOI22_X1 U23261 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20302), .B1(
        n20333), .B2(n20679), .ZN(n20303) );
  OAI211_X1 U23262 ( .C1(n20685), .C2(n20305), .A(n20304), .B(n20303), .ZN(
        P1_U3080) );
  INV_X1 U23263 ( .A(n20333), .ZN(n20306) );
  NAND2_X1 U23264 ( .A1(n20306), .A2(n20765), .ZN(n20307) );
  OAI21_X1 U23265 ( .B1(n20307), .B2(n20361), .A(n20480), .ZN(n20315) );
  NOR2_X1 U23266 ( .A1(n20308), .A2(n13609), .ZN(n20312) );
  INV_X1 U23267 ( .A(n20309), .ZN(n20310) );
  INV_X1 U23268 ( .A(n20625), .ZN(n20498) );
  NOR2_X1 U23269 ( .A1(n20622), .A2(n20311), .ZN(n20344) );
  NAND2_X1 U23270 ( .A1(n20538), .A2(n20344), .ZN(n20313) );
  INV_X1 U23271 ( .A(n20313), .ZN(n20332) );
  AOI22_X1 U23272 ( .A1(n20361), .A2(n20635), .B1(n20626), .B2(n20332), .ZN(
        n20319) );
  INV_X1 U23273 ( .A(n20312), .ZN(n20314) );
  AOI22_X1 U23274 ( .A1(n20315), .A2(n20314), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20313), .ZN(n20317) );
  NAND3_X1 U23275 ( .A1(n20580), .A2(n20317), .A3(n20316), .ZN(n20334) );
  AOI22_X1 U23276 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20334), .B1(
        n20333), .B2(n20582), .ZN(n20318) );
  OAI211_X1 U23277 ( .C1(n20337), .C2(n20498), .A(n20319), .B(n20318), .ZN(
        P1_U3081) );
  INV_X1 U23278 ( .A(n20639), .ZN(n20503) );
  AOI22_X1 U23279 ( .A1(n20361), .A2(n20641), .B1(n20640), .B2(n20332), .ZN(
        n20321) );
  AOI22_X1 U23280 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20334), .B1(
        n20333), .B2(n20586), .ZN(n20320) );
  OAI211_X1 U23281 ( .C1(n20337), .C2(n20503), .A(n20321), .B(n20320), .ZN(
        P1_U3082) );
  INV_X1 U23282 ( .A(n20645), .ZN(n20508) );
  AOI22_X1 U23283 ( .A1(n20333), .A2(n20590), .B1(n20646), .B2(n20332), .ZN(
        n20323) );
  AOI22_X1 U23284 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20334), .B1(
        n20361), .B2(n20647), .ZN(n20322) );
  OAI211_X1 U23285 ( .C1(n20337), .C2(n20508), .A(n20323), .B(n20322), .ZN(
        P1_U3083) );
  INV_X1 U23286 ( .A(n20651), .ZN(n20513) );
  AOI22_X1 U23287 ( .A1(n20333), .A2(n20594), .B1(n20652), .B2(n20332), .ZN(
        n20325) );
  AOI22_X1 U23288 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20334), .B1(
        n20361), .B2(n20653), .ZN(n20324) );
  OAI211_X1 U23289 ( .C1(n20337), .C2(n20513), .A(n20325), .B(n20324), .ZN(
        P1_U3084) );
  INV_X1 U23290 ( .A(n20657), .ZN(n20518) );
  AOI22_X1 U23291 ( .A1(n20333), .A2(n20598), .B1(n20658), .B2(n20332), .ZN(
        n20327) );
  AOI22_X1 U23292 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20334), .B1(
        n20361), .B2(n20659), .ZN(n20326) );
  OAI211_X1 U23293 ( .C1(n20337), .C2(n20518), .A(n20327), .B(n20326), .ZN(
        P1_U3085) );
  INV_X1 U23294 ( .A(n20663), .ZN(n20523) );
  AOI22_X1 U23295 ( .A1(n20333), .A2(n20602), .B1(n20664), .B2(n20332), .ZN(
        n20329) );
  AOI22_X1 U23296 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20334), .B1(
        n20361), .B2(n20665), .ZN(n20328) );
  OAI211_X1 U23297 ( .C1(n20337), .C2(n20523), .A(n20329), .B(n20328), .ZN(
        P1_U3086) );
  INV_X1 U23298 ( .A(n20669), .ZN(n20528) );
  INV_X1 U23299 ( .A(n20674), .ZN(n20606) );
  AOI22_X1 U23300 ( .A1(n20333), .A2(n20606), .B1(n20670), .B2(n20332), .ZN(
        n20331) );
  AOI22_X1 U23301 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20334), .B1(
        n20361), .B2(n20671), .ZN(n20330) );
  OAI211_X1 U23302 ( .C1(n20337), .C2(n20528), .A(n20331), .B(n20330), .ZN(
        P1_U3087) );
  INV_X1 U23303 ( .A(n20676), .ZN(n20536) );
  AOI22_X1 U23304 ( .A1(n20361), .A2(n20679), .B1(n20678), .B2(n20332), .ZN(
        n20336) );
  AOI22_X1 U23305 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20334), .B1(
        n20333), .B2(n20612), .ZN(n20335) );
  OAI211_X1 U23306 ( .C1(n20337), .C2(n20536), .A(n20336), .B(n20335), .ZN(
        P1_U3088) );
  INV_X1 U23307 ( .A(n20338), .ZN(n20360) );
  AOI21_X1 U23308 ( .B1(n20339), .B2(n20619), .A(n20360), .ZN(n20341) );
  INV_X1 U23309 ( .A(n20344), .ZN(n20340) );
  OAI22_X1 U23310 ( .A1(n20341), .A2(n20632), .B1(n20340), .B2(n20623), .ZN(
        n20359) );
  AOI22_X1 U23311 ( .A1(n20626), .A2(n20360), .B1(n20625), .B2(n20359), .ZN(
        n20346) );
  OAI211_X1 U23312 ( .C1(n20342), .C2(n20628), .A(n20765), .B(n20341), .ZN(
        n20343) );
  OAI211_X1 U23313 ( .C1(n20458), .C2(n20344), .A(n20630), .B(n20343), .ZN(
        n20362) );
  AOI22_X1 U23314 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20362), .B1(
        n20361), .B2(n20582), .ZN(n20345) );
  OAI211_X1 U23315 ( .C1(n20585), .C2(n20371), .A(n20346), .B(n20345), .ZN(
        P1_U3089) );
  AOI22_X1 U23316 ( .A1(n20640), .A2(n20360), .B1(n20639), .B2(n20359), .ZN(
        n20348) );
  AOI22_X1 U23317 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20362), .B1(
        n20361), .B2(n20586), .ZN(n20347) );
  OAI211_X1 U23318 ( .C1(n20589), .C2(n20371), .A(n20348), .B(n20347), .ZN(
        P1_U3090) );
  AOI22_X1 U23319 ( .A1(n20646), .A2(n20360), .B1(n20645), .B2(n20359), .ZN(
        n20350) );
  AOI22_X1 U23320 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20362), .B1(
        n20361), .B2(n20590), .ZN(n20349) );
  OAI211_X1 U23321 ( .C1(n20593), .C2(n20371), .A(n20350), .B(n20349), .ZN(
        P1_U3091) );
  AOI22_X1 U23322 ( .A1(n20652), .A2(n20360), .B1(n20651), .B2(n20359), .ZN(
        n20352) );
  AOI22_X1 U23323 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20362), .B1(
        n20361), .B2(n20594), .ZN(n20351) );
  OAI211_X1 U23324 ( .C1(n20597), .C2(n20371), .A(n20352), .B(n20351), .ZN(
        P1_U3092) );
  AOI22_X1 U23325 ( .A1(n20658), .A2(n20360), .B1(n20657), .B2(n20359), .ZN(
        n20354) );
  AOI22_X1 U23326 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20362), .B1(
        n20361), .B2(n20598), .ZN(n20353) );
  OAI211_X1 U23327 ( .C1(n20601), .C2(n20371), .A(n20354), .B(n20353), .ZN(
        P1_U3093) );
  AOI22_X1 U23328 ( .A1(n20664), .A2(n20360), .B1(n20663), .B2(n20359), .ZN(
        n20356) );
  AOI22_X1 U23329 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20362), .B1(
        n20361), .B2(n20602), .ZN(n20355) );
  OAI211_X1 U23330 ( .C1(n20605), .C2(n20371), .A(n20356), .B(n20355), .ZN(
        P1_U3094) );
  AOI22_X1 U23331 ( .A1(n20670), .A2(n20360), .B1(n20669), .B2(n20359), .ZN(
        n20358) );
  AOI22_X1 U23332 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20362), .B1(
        n20361), .B2(n20606), .ZN(n20357) );
  OAI211_X1 U23333 ( .C1(n20609), .C2(n20371), .A(n20358), .B(n20357), .ZN(
        P1_U3095) );
  AOI22_X1 U23334 ( .A1(n20678), .A2(n20360), .B1(n20676), .B2(n20359), .ZN(
        n20364) );
  AOI22_X1 U23335 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20362), .B1(
        n20361), .B2(n20612), .ZN(n20363) );
  OAI211_X1 U23336 ( .C1(n20617), .C2(n20371), .A(n20364), .B(n20363), .ZN(
        P1_U3096) );
  NAND2_X1 U23337 ( .A1(n20367), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20451) );
  AND2_X1 U23338 ( .A1(n20760), .A2(n13438), .ZN(n20452) );
  AOI21_X1 U23339 ( .B1(n20452), .B2(n13609), .A(n10240), .ZN(n20373) );
  NOR2_X1 U23340 ( .A1(n20369), .A2(n20368), .ZN(n20483) );
  INV_X1 U23341 ( .A(n20483), .ZN(n20489) );
  OAI22_X1 U23342 ( .A1(n20373), .A2(n20632), .B1(n20370), .B2(n20489), .ZN(
        n20390) );
  AOI22_X1 U23343 ( .A1(n20626), .A2(n10240), .B1(n20625), .B2(n20390), .ZN(
        n20377) );
  INV_X1 U23344 ( .A(n20418), .ZN(n20372) );
  OAI21_X1 U23345 ( .B1(n20372), .B2(n20391), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20374) );
  NAND2_X1 U23346 ( .A1(n20374), .A2(n20373), .ZN(n20375) );
  AOI22_X1 U23347 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20392), .B1(
        n20391), .B2(n20582), .ZN(n20376) );
  OAI211_X1 U23348 ( .C1(n20585), .C2(n20418), .A(n20377), .B(n20376), .ZN(
        P1_U3097) );
  AOI22_X1 U23349 ( .A1(n20640), .A2(n10240), .B1(n20639), .B2(n20390), .ZN(
        n20379) );
  AOI22_X1 U23350 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20392), .B1(
        n20391), .B2(n20586), .ZN(n20378) );
  OAI211_X1 U23351 ( .C1(n20589), .C2(n20418), .A(n20379), .B(n20378), .ZN(
        P1_U3098) );
  AOI22_X1 U23352 ( .A1(n20646), .A2(n10240), .B1(n20645), .B2(n20390), .ZN(
        n20381) );
  AOI22_X1 U23353 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20392), .B1(
        n20391), .B2(n20590), .ZN(n20380) );
  OAI211_X1 U23354 ( .C1(n20593), .C2(n20418), .A(n20381), .B(n20380), .ZN(
        P1_U3099) );
  AOI22_X1 U23355 ( .A1(n20652), .A2(n10240), .B1(n20651), .B2(n20390), .ZN(
        n20383) );
  AOI22_X1 U23356 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20392), .B1(
        n20391), .B2(n20594), .ZN(n20382) );
  OAI211_X1 U23357 ( .C1(n20597), .C2(n20418), .A(n20383), .B(n20382), .ZN(
        P1_U3100) );
  AOI22_X1 U23358 ( .A1(n20658), .A2(n10240), .B1(n20657), .B2(n20390), .ZN(
        n20385) );
  AOI22_X1 U23359 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20392), .B1(
        n20391), .B2(n20598), .ZN(n20384) );
  OAI211_X1 U23360 ( .C1(n20601), .C2(n20418), .A(n20385), .B(n20384), .ZN(
        P1_U3101) );
  AOI22_X1 U23361 ( .A1(n20664), .A2(n10240), .B1(n20663), .B2(n20390), .ZN(
        n20387) );
  AOI22_X1 U23362 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20392), .B1(
        n20391), .B2(n20602), .ZN(n20386) );
  OAI211_X1 U23363 ( .C1(n20605), .C2(n20418), .A(n20387), .B(n20386), .ZN(
        P1_U3102) );
  AOI22_X1 U23364 ( .A1(n20670), .A2(n10240), .B1(n20669), .B2(n20390), .ZN(
        n20389) );
  AOI22_X1 U23365 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20392), .B1(
        n20391), .B2(n20606), .ZN(n20388) );
  OAI211_X1 U23366 ( .C1(n20609), .C2(n20418), .A(n20389), .B(n20388), .ZN(
        P1_U3103) );
  AOI22_X1 U23367 ( .A1(n20678), .A2(n10240), .B1(n20676), .B2(n20390), .ZN(
        n20394) );
  AOI22_X1 U23368 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20392), .B1(
        n20391), .B2(n20612), .ZN(n20393) );
  OAI211_X1 U23369 ( .C1(n20617), .C2(n20418), .A(n20394), .B(n20393), .ZN(
        P1_U3104) );
  NOR2_X1 U23370 ( .A1(n20451), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20398) );
  INV_X1 U23371 ( .A(n20398), .ZN(n20395) );
  NOR2_X1 U23372 ( .A1(n20538), .A2(n20395), .ZN(n20414) );
  AOI21_X1 U23373 ( .B1(n20452), .B2(n20540), .A(n20414), .ZN(n20396) );
  OAI22_X1 U23374 ( .A1(n20396), .A2(n20632), .B1(n20395), .B2(n20623), .ZN(
        n20413) );
  AOI22_X1 U23375 ( .A1(n20626), .A2(n20414), .B1(n20625), .B2(n20413), .ZN(
        n20400) );
  INV_X1 U23376 ( .A(n20759), .ZN(n20455) );
  OAI211_X1 U23377 ( .C1(n20455), .C2(n20574), .A(n20765), .B(n20396), .ZN(
        n20397) );
  OAI211_X1 U23378 ( .C1(n20458), .C2(n20398), .A(n20630), .B(n20397), .ZN(
        n20415) );
  AOI22_X1 U23379 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20415), .B1(
        n20445), .B2(n20635), .ZN(n20399) );
  OAI211_X1 U23380 ( .C1(n20638), .C2(n20418), .A(n20400), .B(n20399), .ZN(
        P1_U3105) );
  AOI22_X1 U23381 ( .A1(n20640), .A2(n20414), .B1(n20639), .B2(n20413), .ZN(
        n20402) );
  AOI22_X1 U23382 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20415), .B1(
        n20445), .B2(n20641), .ZN(n20401) );
  OAI211_X1 U23383 ( .C1(n20644), .C2(n20418), .A(n20402), .B(n20401), .ZN(
        P1_U3106) );
  AOI22_X1 U23384 ( .A1(n20646), .A2(n20414), .B1(n20645), .B2(n20413), .ZN(
        n20404) );
  AOI22_X1 U23385 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20415), .B1(
        n20445), .B2(n20647), .ZN(n20403) );
  OAI211_X1 U23386 ( .C1(n20650), .C2(n20418), .A(n20404), .B(n20403), .ZN(
        P1_U3107) );
  AOI22_X1 U23387 ( .A1(n20652), .A2(n20414), .B1(n20651), .B2(n20413), .ZN(
        n20406) );
  AOI22_X1 U23388 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20415), .B1(
        n20445), .B2(n20653), .ZN(n20405) );
  OAI211_X1 U23389 ( .C1(n20656), .C2(n20418), .A(n20406), .B(n20405), .ZN(
        P1_U3108) );
  AOI22_X1 U23390 ( .A1(n20658), .A2(n20414), .B1(n20657), .B2(n20413), .ZN(
        n20408) );
  AOI22_X1 U23391 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20415), .B1(
        n20445), .B2(n20659), .ZN(n20407) );
  OAI211_X1 U23392 ( .C1(n20662), .C2(n20418), .A(n20408), .B(n20407), .ZN(
        P1_U3109) );
  AOI22_X1 U23393 ( .A1(n20664), .A2(n20414), .B1(n20663), .B2(n20413), .ZN(
        n20410) );
  AOI22_X1 U23394 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20415), .B1(
        n20445), .B2(n20665), .ZN(n20409) );
  OAI211_X1 U23395 ( .C1(n20668), .C2(n20418), .A(n20410), .B(n20409), .ZN(
        P1_U3110) );
  AOI22_X1 U23396 ( .A1(n20670), .A2(n20414), .B1(n20669), .B2(n20413), .ZN(
        n20412) );
  AOI22_X1 U23397 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20415), .B1(
        n20445), .B2(n20671), .ZN(n20411) );
  OAI211_X1 U23398 ( .C1(n20674), .C2(n20418), .A(n20412), .B(n20411), .ZN(
        P1_U3111) );
  AOI22_X1 U23399 ( .A1(n20678), .A2(n20414), .B1(n20676), .B2(n20413), .ZN(
        n20417) );
  AOI22_X1 U23400 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20415), .B1(
        n20445), .B2(n20679), .ZN(n20416) );
  OAI211_X1 U23401 ( .C1(n20685), .C2(n20418), .A(n20417), .B(n20416), .ZN(
        P1_U3112) );
  INV_X1 U23402 ( .A(n20445), .ZN(n20419) );
  NAND2_X1 U23403 ( .A1(n20419), .A2(n20765), .ZN(n20420) );
  OAI21_X1 U23404 ( .B1(n20420), .B2(n20475), .A(n20480), .ZN(n20427) );
  AND2_X1 U23405 ( .A1(n20452), .A2(n20577), .ZN(n20424) );
  OR2_X1 U23406 ( .A1(n20421), .A2(n20773), .ZN(n20572) );
  INV_X1 U23407 ( .A(n20572), .ZN(n20423) );
  NOR2_X1 U23408 ( .A1(n20622), .A2(n20451), .ZN(n20457) );
  NAND2_X1 U23409 ( .A1(n20538), .A2(n20457), .ZN(n20425) );
  INV_X1 U23410 ( .A(n20425), .ZN(n20444) );
  AOI22_X1 U23411 ( .A1(n20475), .A2(n20635), .B1(n20626), .B2(n20444), .ZN(
        n20431) );
  INV_X1 U23412 ( .A(n20424), .ZN(n20426) );
  AOI22_X1 U23413 ( .A1(n20427), .A2(n20426), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20425), .ZN(n20428) );
  NAND2_X1 U23414 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20572), .ZN(n20579) );
  NAND3_X1 U23415 ( .A1(n20429), .A2(n20428), .A3(n20579), .ZN(n20446) );
  AOI22_X1 U23416 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20446), .B1(
        n20445), .B2(n20582), .ZN(n20430) );
  OAI211_X1 U23417 ( .C1(n20449), .C2(n20498), .A(n20431), .B(n20430), .ZN(
        P1_U3113) );
  AOI22_X1 U23418 ( .A1(n20445), .A2(n20586), .B1(n20444), .B2(n20640), .ZN(
        n20433) );
  AOI22_X1 U23419 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20446), .B1(
        n20475), .B2(n20641), .ZN(n20432) );
  OAI211_X1 U23420 ( .C1(n20449), .C2(n20503), .A(n20433), .B(n20432), .ZN(
        P1_U3114) );
  AOI22_X1 U23421 ( .A1(n20445), .A2(n20590), .B1(n20444), .B2(n20646), .ZN(
        n20435) );
  AOI22_X1 U23422 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20446), .B1(
        n20475), .B2(n20647), .ZN(n20434) );
  OAI211_X1 U23423 ( .C1(n20449), .C2(n20508), .A(n20435), .B(n20434), .ZN(
        P1_U3115) );
  AOI22_X1 U23424 ( .A1(n20475), .A2(n20653), .B1(n20444), .B2(n20652), .ZN(
        n20437) );
  AOI22_X1 U23425 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20446), .B1(
        n20445), .B2(n20594), .ZN(n20436) );
  OAI211_X1 U23426 ( .C1(n20449), .C2(n20513), .A(n20437), .B(n20436), .ZN(
        P1_U3116) );
  AOI22_X1 U23427 ( .A1(n20445), .A2(n20598), .B1(n20444), .B2(n20658), .ZN(
        n20439) );
  AOI22_X1 U23428 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20446), .B1(
        n20475), .B2(n20659), .ZN(n20438) );
  OAI211_X1 U23429 ( .C1(n20449), .C2(n20518), .A(n20439), .B(n20438), .ZN(
        P1_U3117) );
  AOI22_X1 U23430 ( .A1(n20445), .A2(n20602), .B1(n20444), .B2(n20664), .ZN(
        n20441) );
  AOI22_X1 U23431 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20446), .B1(
        n20475), .B2(n20665), .ZN(n20440) );
  OAI211_X1 U23432 ( .C1(n20449), .C2(n20523), .A(n20441), .B(n20440), .ZN(
        P1_U3118) );
  AOI22_X1 U23433 ( .A1(n20475), .A2(n20671), .B1(n20444), .B2(n20670), .ZN(
        n20443) );
  AOI22_X1 U23434 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20446), .B1(
        n20445), .B2(n20606), .ZN(n20442) );
  OAI211_X1 U23435 ( .C1(n20449), .C2(n20528), .A(n20443), .B(n20442), .ZN(
        P1_U3119) );
  AOI22_X1 U23436 ( .A1(n20445), .A2(n20612), .B1(n20444), .B2(n20678), .ZN(
        n20448) );
  AOI22_X1 U23437 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20446), .B1(
        n20475), .B2(n20679), .ZN(n20447) );
  OAI211_X1 U23438 ( .C1(n20449), .C2(n20536), .A(n20448), .B(n20447), .ZN(
        P1_U3120) );
  NOR2_X1 U23439 ( .A1(n20618), .A2(n20451), .ZN(n20474) );
  AOI21_X1 U23440 ( .B1(n20452), .B2(n20619), .A(n20474), .ZN(n20454) );
  INV_X1 U23441 ( .A(n20457), .ZN(n20453) );
  OAI22_X1 U23442 ( .A1(n20454), .A2(n20632), .B1(n20453), .B2(n20623), .ZN(
        n20473) );
  AOI22_X1 U23443 ( .A1(n20626), .A2(n20474), .B1(n20625), .B2(n20473), .ZN(
        n20460) );
  OAI211_X1 U23444 ( .C1(n20455), .C2(n20628), .A(n20765), .B(n20454), .ZN(
        n20456) );
  OAI211_X1 U23445 ( .C1(n20458), .C2(n20457), .A(n20630), .B(n20456), .ZN(
        n20476) );
  AOI22_X1 U23446 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20476), .B1(
        n20475), .B2(n20582), .ZN(n20459) );
  OAI211_X1 U23447 ( .C1(n20585), .C2(n20495), .A(n20460), .B(n20459), .ZN(
        P1_U3121) );
  AOI22_X1 U23448 ( .A1(n20640), .A2(n20474), .B1(n20639), .B2(n20473), .ZN(
        n20462) );
  AOI22_X1 U23449 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20476), .B1(
        n20475), .B2(n20586), .ZN(n20461) );
  OAI211_X1 U23450 ( .C1(n20589), .C2(n20495), .A(n20462), .B(n20461), .ZN(
        P1_U3122) );
  AOI22_X1 U23451 ( .A1(n20646), .A2(n20474), .B1(n20645), .B2(n20473), .ZN(
        n20464) );
  AOI22_X1 U23452 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20476), .B1(
        n20475), .B2(n20590), .ZN(n20463) );
  OAI211_X1 U23453 ( .C1(n20593), .C2(n20495), .A(n20464), .B(n20463), .ZN(
        P1_U3123) );
  AOI22_X1 U23454 ( .A1(n20652), .A2(n20474), .B1(n20651), .B2(n20473), .ZN(
        n20466) );
  AOI22_X1 U23455 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20476), .B1(
        n20475), .B2(n20594), .ZN(n20465) );
  OAI211_X1 U23456 ( .C1(n20597), .C2(n20495), .A(n20466), .B(n20465), .ZN(
        P1_U3124) );
  AOI22_X1 U23457 ( .A1(n20658), .A2(n20474), .B1(n20657), .B2(n20473), .ZN(
        n20468) );
  AOI22_X1 U23458 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20476), .B1(
        n20475), .B2(n20598), .ZN(n20467) );
  OAI211_X1 U23459 ( .C1(n20601), .C2(n20495), .A(n20468), .B(n20467), .ZN(
        P1_U3125) );
  AOI22_X1 U23460 ( .A1(n20664), .A2(n20474), .B1(n20663), .B2(n20473), .ZN(
        n20470) );
  AOI22_X1 U23461 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20476), .B1(
        n20475), .B2(n20602), .ZN(n20469) );
  OAI211_X1 U23462 ( .C1(n20605), .C2(n20495), .A(n20470), .B(n20469), .ZN(
        P1_U3126) );
  AOI22_X1 U23463 ( .A1(n20670), .A2(n20474), .B1(n20669), .B2(n20473), .ZN(
        n20472) );
  AOI22_X1 U23464 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20476), .B1(
        n20475), .B2(n20606), .ZN(n20471) );
  OAI211_X1 U23465 ( .C1(n20609), .C2(n20495), .A(n20472), .B(n20471), .ZN(
        P1_U3127) );
  AOI22_X1 U23466 ( .A1(n20678), .A2(n20474), .B1(n20676), .B2(n20473), .ZN(
        n20478) );
  AOI22_X1 U23467 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20476), .B1(
        n20475), .B2(n20612), .ZN(n20477) );
  OAI211_X1 U23468 ( .C1(n20617), .C2(n20495), .A(n20478), .B(n20477), .ZN(
        P1_U3128) );
  NAND3_X1 U23469 ( .A1(n20495), .A2(n20765), .A3(n20568), .ZN(n20481) );
  NAND2_X1 U23470 ( .A1(n20481), .A2(n20480), .ZN(n20491) );
  OR2_X1 U23471 ( .A1(n13438), .A2(n20482), .ZN(n20539) );
  NOR2_X1 U23472 ( .A1(n20539), .A2(n20577), .ZN(n20488) );
  NAND2_X1 U23473 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20621) );
  OR2_X1 U23474 ( .A1(n20485), .A2(n20621), .ZN(n20529) );
  OAI22_X1 U23475 ( .A1(n20568), .A2(n20585), .B1(n20486), .B2(n20529), .ZN(
        n20487) );
  INV_X1 U23476 ( .A(n20487), .ZN(n20497) );
  INV_X1 U23477 ( .A(n20529), .ZN(n20494) );
  INV_X1 U23478 ( .A(n20488), .ZN(n20490) );
  AOI22_X1 U23479 ( .A1(n20491), .A2(n20490), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20489), .ZN(n20492) );
  AOI22_X1 U23480 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20533), .B1(
        n20532), .B2(n20582), .ZN(n20496) );
  OAI211_X1 U23481 ( .C1(n20537), .C2(n20498), .A(n20497), .B(n20496), .ZN(
        P1_U3129) );
  OAI22_X1 U23482 ( .A1(n20568), .A2(n20589), .B1(n20499), .B2(n20529), .ZN(
        n20500) );
  INV_X1 U23483 ( .A(n20500), .ZN(n20502) );
  AOI22_X1 U23484 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20533), .B1(
        n20532), .B2(n20586), .ZN(n20501) );
  OAI211_X1 U23485 ( .C1(n20537), .C2(n20503), .A(n20502), .B(n20501), .ZN(
        P1_U3130) );
  OAI22_X1 U23486 ( .A1(n20568), .A2(n20593), .B1(n20504), .B2(n20529), .ZN(
        n20505) );
  INV_X1 U23487 ( .A(n20505), .ZN(n20507) );
  AOI22_X1 U23488 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20533), .B1(
        n20532), .B2(n20590), .ZN(n20506) );
  OAI211_X1 U23489 ( .C1(n20537), .C2(n20508), .A(n20507), .B(n20506), .ZN(
        P1_U3131) );
  OAI22_X1 U23490 ( .A1(n20568), .A2(n20597), .B1(n20509), .B2(n20529), .ZN(
        n20510) );
  INV_X1 U23491 ( .A(n20510), .ZN(n20512) );
  AOI22_X1 U23492 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20533), .B1(
        n20532), .B2(n20594), .ZN(n20511) );
  OAI211_X1 U23493 ( .C1(n20537), .C2(n20513), .A(n20512), .B(n20511), .ZN(
        P1_U3132) );
  OAI22_X1 U23494 ( .A1(n20568), .A2(n20601), .B1(n20514), .B2(n20529), .ZN(
        n20515) );
  INV_X1 U23495 ( .A(n20515), .ZN(n20517) );
  AOI22_X1 U23496 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20533), .B1(
        n20532), .B2(n20598), .ZN(n20516) );
  OAI211_X1 U23497 ( .C1(n20537), .C2(n20518), .A(n20517), .B(n20516), .ZN(
        P1_U3133) );
  OAI22_X1 U23498 ( .A1(n20568), .A2(n20605), .B1(n20519), .B2(n20529), .ZN(
        n20520) );
  INV_X1 U23499 ( .A(n20520), .ZN(n20522) );
  AOI22_X1 U23500 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20533), .B1(
        n20532), .B2(n20602), .ZN(n20521) );
  OAI211_X1 U23501 ( .C1(n20537), .C2(n20523), .A(n20522), .B(n20521), .ZN(
        P1_U3134) );
  OAI22_X1 U23502 ( .A1(n20568), .A2(n20609), .B1(n20524), .B2(n20529), .ZN(
        n20525) );
  INV_X1 U23503 ( .A(n20525), .ZN(n20527) );
  AOI22_X1 U23504 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20533), .B1(
        n20532), .B2(n20606), .ZN(n20526) );
  OAI211_X1 U23505 ( .C1(n20537), .C2(n20528), .A(n20527), .B(n20526), .ZN(
        P1_U3135) );
  OAI22_X1 U23506 ( .A1(n20568), .A2(n20617), .B1(n20530), .B2(n20529), .ZN(
        n20531) );
  INV_X1 U23507 ( .A(n20531), .ZN(n20535) );
  AOI22_X1 U23508 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20533), .B1(
        n20532), .B2(n20612), .ZN(n20534) );
  OAI211_X1 U23509 ( .C1(n20537), .C2(n20536), .A(n20535), .B(n20534), .ZN(
        P1_U3136) );
  NOR3_X2 U23510 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20538), .A3(
        n20621), .ZN(n20564) );
  AOI21_X1 U23511 ( .B1(n20620), .B2(n20540), .A(n20564), .ZN(n20542) );
  NOR2_X1 U23512 ( .A1(n20621), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20545) );
  INV_X1 U23513 ( .A(n20545), .ZN(n20541) );
  OAI22_X1 U23514 ( .A1(n20542), .A2(n20632), .B1(n20541), .B2(n20623), .ZN(
        n20563) );
  AOI22_X1 U23515 ( .A1(n20626), .A2(n20564), .B1(n20625), .B2(n20563), .ZN(
        n20550) );
  OR3_X1 U23516 ( .A1(n20629), .A2(n20544), .A3(n20543), .ZN(n20768) );
  INV_X1 U23517 ( .A(n20768), .ZN(n20546) );
  INV_X1 U23518 ( .A(n20547), .ZN(n20548) );
  AOI22_X1 U23519 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20565), .B1(
        n20613), .B2(n20635), .ZN(n20549) );
  OAI211_X1 U23520 ( .C1(n20638), .C2(n20568), .A(n20550), .B(n20549), .ZN(
        P1_U3137) );
  AOI22_X1 U23521 ( .A1(n20640), .A2(n20564), .B1(n20639), .B2(n20563), .ZN(
        n20552) );
  AOI22_X1 U23522 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20565), .B1(
        n20613), .B2(n20641), .ZN(n20551) );
  OAI211_X1 U23523 ( .C1(n20644), .C2(n20568), .A(n20552), .B(n20551), .ZN(
        P1_U3138) );
  AOI22_X1 U23524 ( .A1(n20646), .A2(n20564), .B1(n20645), .B2(n20563), .ZN(
        n20554) );
  AOI22_X1 U23525 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20565), .B1(
        n20613), .B2(n20647), .ZN(n20553) );
  OAI211_X1 U23526 ( .C1(n20650), .C2(n20568), .A(n20554), .B(n20553), .ZN(
        P1_U3139) );
  AOI22_X1 U23527 ( .A1(n20652), .A2(n20564), .B1(n20651), .B2(n20563), .ZN(
        n20556) );
  AOI22_X1 U23528 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20565), .B1(
        n20613), .B2(n20653), .ZN(n20555) );
  OAI211_X1 U23529 ( .C1(n20656), .C2(n20568), .A(n20556), .B(n20555), .ZN(
        P1_U3140) );
  AOI22_X1 U23530 ( .A1(n20658), .A2(n20564), .B1(n20657), .B2(n20563), .ZN(
        n20558) );
  AOI22_X1 U23531 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20565), .B1(
        n20613), .B2(n20659), .ZN(n20557) );
  OAI211_X1 U23532 ( .C1(n20662), .C2(n20568), .A(n20558), .B(n20557), .ZN(
        P1_U3141) );
  AOI22_X1 U23533 ( .A1(n20664), .A2(n20564), .B1(n20663), .B2(n20563), .ZN(
        n20560) );
  AOI22_X1 U23534 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20565), .B1(
        n20613), .B2(n20665), .ZN(n20559) );
  OAI211_X1 U23535 ( .C1(n20668), .C2(n20568), .A(n20560), .B(n20559), .ZN(
        P1_U3142) );
  AOI22_X1 U23536 ( .A1(n20670), .A2(n20564), .B1(n20669), .B2(n20563), .ZN(
        n20562) );
  AOI22_X1 U23537 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20565), .B1(
        n20613), .B2(n20671), .ZN(n20561) );
  OAI211_X1 U23538 ( .C1(n20674), .C2(n20568), .A(n20562), .B(n20561), .ZN(
        P1_U3143) );
  AOI22_X1 U23539 ( .A1(n20678), .A2(n20564), .B1(n20676), .B2(n20563), .ZN(
        n20567) );
  AOI22_X1 U23540 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20565), .B1(
        n20613), .B2(n20679), .ZN(n20566) );
  OAI211_X1 U23541 ( .C1(n20685), .C2(n20568), .A(n20567), .B(n20566), .ZN(
        P1_U3144) );
  INV_X1 U23542 ( .A(n20629), .ZN(n20570) );
  NOR3_X2 U23543 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20622), .A3(
        n20621), .ZN(n20611) );
  NAND3_X1 U23544 ( .A1(n20620), .A2(n20577), .A3(n20765), .ZN(n20571) );
  OAI21_X1 U23545 ( .B1(n20573), .B2(n20572), .A(n20571), .ZN(n20610) );
  AOI22_X1 U23546 ( .A1(n20626), .A2(n20611), .B1(n20625), .B2(n20610), .ZN(
        n20584) );
  AOI21_X1 U23547 ( .B1(n20684), .B2(n20575), .A(n20574), .ZN(n20576) );
  AOI21_X1 U23548 ( .B1(n20620), .B2(n20577), .A(n20576), .ZN(n20578) );
  NOR2_X1 U23549 ( .A1(n20578), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20581) );
  AOI22_X1 U23550 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20614), .B1(
        n20613), .B2(n20582), .ZN(n20583) );
  OAI211_X1 U23551 ( .C1(n20585), .C2(n20684), .A(n20584), .B(n20583), .ZN(
        P1_U3145) );
  AOI22_X1 U23552 ( .A1(n20640), .A2(n20611), .B1(n20639), .B2(n20610), .ZN(
        n20588) );
  AOI22_X1 U23553 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20614), .B1(
        n20613), .B2(n20586), .ZN(n20587) );
  OAI211_X1 U23554 ( .C1(n20589), .C2(n20684), .A(n20588), .B(n20587), .ZN(
        P1_U3146) );
  AOI22_X1 U23555 ( .A1(n20646), .A2(n20611), .B1(n20645), .B2(n20610), .ZN(
        n20592) );
  AOI22_X1 U23556 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20614), .B1(
        n20613), .B2(n20590), .ZN(n20591) );
  OAI211_X1 U23557 ( .C1(n20593), .C2(n20684), .A(n20592), .B(n20591), .ZN(
        P1_U3147) );
  AOI22_X1 U23558 ( .A1(n20652), .A2(n20611), .B1(n20651), .B2(n20610), .ZN(
        n20596) );
  AOI22_X1 U23559 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20614), .B1(
        n20613), .B2(n20594), .ZN(n20595) );
  OAI211_X1 U23560 ( .C1(n20597), .C2(n20684), .A(n20596), .B(n20595), .ZN(
        P1_U3148) );
  AOI22_X1 U23561 ( .A1(n20658), .A2(n20611), .B1(n20657), .B2(n20610), .ZN(
        n20600) );
  AOI22_X1 U23562 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20614), .B1(
        n20613), .B2(n20598), .ZN(n20599) );
  OAI211_X1 U23563 ( .C1(n20601), .C2(n20684), .A(n20600), .B(n20599), .ZN(
        P1_U3149) );
  AOI22_X1 U23564 ( .A1(n20664), .A2(n20611), .B1(n20663), .B2(n20610), .ZN(
        n20604) );
  AOI22_X1 U23565 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20614), .B1(
        n20613), .B2(n20602), .ZN(n20603) );
  OAI211_X1 U23566 ( .C1(n20605), .C2(n20684), .A(n20604), .B(n20603), .ZN(
        P1_U3150) );
  AOI22_X1 U23567 ( .A1(n20670), .A2(n20611), .B1(n20669), .B2(n20610), .ZN(
        n20608) );
  AOI22_X1 U23568 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20614), .B1(
        n20613), .B2(n20606), .ZN(n20607) );
  OAI211_X1 U23569 ( .C1(n20609), .C2(n20684), .A(n20608), .B(n20607), .ZN(
        P1_U3151) );
  AOI22_X1 U23570 ( .A1(n20678), .A2(n20611), .B1(n20676), .B2(n20610), .ZN(
        n20616) );
  AOI22_X1 U23571 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20614), .B1(
        n20613), .B2(n20612), .ZN(n20615) );
  OAI211_X1 U23572 ( .C1(n20617), .C2(n20684), .A(n20616), .B(n20615), .ZN(
        P1_U3152) );
  NOR2_X1 U23573 ( .A1(n20618), .A2(n20621), .ZN(n20677) );
  AOI21_X1 U23574 ( .B1(n20620), .B2(n20619), .A(n20677), .ZN(n20627) );
  NOR2_X1 U23575 ( .A1(n20622), .A2(n20621), .ZN(n20633) );
  INV_X1 U23576 ( .A(n20633), .ZN(n20624) );
  OAI22_X1 U23577 ( .A1(n20627), .A2(n20632), .B1(n20624), .B2(n20623), .ZN(
        n20675) );
  AOI22_X1 U23578 ( .A1(n20626), .A2(n20677), .B1(n20625), .B2(n20675), .ZN(
        n20637) );
  OAI21_X1 U23579 ( .B1(n20629), .B2(n20628), .A(n20627), .ZN(n20631) );
  OAI221_X1 U23580 ( .B1(n20765), .B2(n20633), .C1(n20632), .C2(n20631), .A(
        n20630), .ZN(n20681) );
  AOI22_X1 U23581 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20681), .B1(
        n20680), .B2(n20635), .ZN(n20636) );
  OAI211_X1 U23582 ( .C1(n20638), .C2(n20684), .A(n20637), .B(n20636), .ZN(
        P1_U3153) );
  AOI22_X1 U23583 ( .A1(n20640), .A2(n20677), .B1(n20639), .B2(n20675), .ZN(
        n20643) );
  AOI22_X1 U23584 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20681), .B1(
        n20680), .B2(n20641), .ZN(n20642) );
  OAI211_X1 U23585 ( .C1(n20644), .C2(n20684), .A(n20643), .B(n20642), .ZN(
        P1_U3154) );
  AOI22_X1 U23586 ( .A1(n20646), .A2(n20677), .B1(n20645), .B2(n20675), .ZN(
        n20649) );
  AOI22_X1 U23587 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20681), .B1(
        n20680), .B2(n20647), .ZN(n20648) );
  OAI211_X1 U23588 ( .C1(n20650), .C2(n20684), .A(n20649), .B(n20648), .ZN(
        P1_U3155) );
  AOI22_X1 U23589 ( .A1(n20652), .A2(n20677), .B1(n20651), .B2(n20675), .ZN(
        n20655) );
  AOI22_X1 U23590 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20681), .B1(
        n20680), .B2(n20653), .ZN(n20654) );
  OAI211_X1 U23591 ( .C1(n20656), .C2(n20684), .A(n20655), .B(n20654), .ZN(
        P1_U3156) );
  AOI22_X1 U23592 ( .A1(n20658), .A2(n20677), .B1(n20657), .B2(n20675), .ZN(
        n20661) );
  AOI22_X1 U23593 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20681), .B1(
        n20680), .B2(n20659), .ZN(n20660) );
  OAI211_X1 U23594 ( .C1(n20662), .C2(n20684), .A(n20661), .B(n20660), .ZN(
        P1_U3157) );
  AOI22_X1 U23595 ( .A1(n20664), .A2(n20677), .B1(n20663), .B2(n20675), .ZN(
        n20667) );
  AOI22_X1 U23596 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20681), .B1(
        n20680), .B2(n20665), .ZN(n20666) );
  OAI211_X1 U23597 ( .C1(n20668), .C2(n20684), .A(n20667), .B(n20666), .ZN(
        P1_U3158) );
  AOI22_X1 U23598 ( .A1(n20670), .A2(n20677), .B1(n20669), .B2(n20675), .ZN(
        n20673) );
  AOI22_X1 U23599 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20681), .B1(
        n20680), .B2(n20671), .ZN(n20672) );
  OAI211_X1 U23600 ( .C1(n20674), .C2(n20684), .A(n20673), .B(n20672), .ZN(
        P1_U3159) );
  AOI22_X1 U23601 ( .A1(n20678), .A2(n20677), .B1(n20676), .B2(n20675), .ZN(
        n20683) );
  AOI22_X1 U23602 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20681), .B1(
        n20680), .B2(n20679), .ZN(n20682) );
  OAI211_X1 U23603 ( .C1(n20685), .C2(n20684), .A(n20683), .B(n20682), .ZN(
        P1_U3160) );
  OR3_X1 U23604 ( .A1(n20687), .A2(n20788), .A3(n20686), .ZN(P1_U3163) );
  AND2_X1 U23605 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n20688), .ZN(
        P1_U3164) );
  AND2_X1 U23606 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n20688), .ZN(
        P1_U3165) );
  AND2_X1 U23607 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n20688), .ZN(
        P1_U3166) );
  AND2_X1 U23608 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n20688), .ZN(
        P1_U3167) );
  AND2_X1 U23609 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n20688), .ZN(
        P1_U3168) );
  AND2_X1 U23610 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n20688), .ZN(
        P1_U3169) );
  AND2_X1 U23611 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n20688), .ZN(
        P1_U3170) );
  AND2_X1 U23612 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n20688), .ZN(
        P1_U3171) );
  AND2_X1 U23613 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n20688), .ZN(
        P1_U3172) );
  AND2_X1 U23614 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n20688), .ZN(
        P1_U3173) );
  AND2_X1 U23615 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n20688), .ZN(
        P1_U3174) );
  INV_X1 U23616 ( .A(P1_DATAWIDTH_REG_20__SCAN_IN), .ZN(n21022) );
  NOR2_X1 U23617 ( .A1(n20757), .A2(n21022), .ZN(P1_U3175) );
  AND2_X1 U23618 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n20688), .ZN(
        P1_U3176) );
  AND2_X1 U23619 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n20688), .ZN(
        P1_U3177) );
  AND2_X1 U23620 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n20688), .ZN(
        P1_U3178) );
  AND2_X1 U23621 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n20688), .ZN(
        P1_U3179) );
  AND2_X1 U23622 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n20688), .ZN(
        P1_U3180) );
  AND2_X1 U23623 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n20688), .ZN(
        P1_U3181) );
  INV_X1 U23624 ( .A(P1_DATAWIDTH_REG_13__SCAN_IN), .ZN(n20994) );
  NOR2_X1 U23625 ( .A1(n20757), .A2(n20994), .ZN(P1_U3182) );
  AND2_X1 U23626 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n20688), .ZN(
        P1_U3183) );
  AND2_X1 U23627 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n20688), .ZN(
        P1_U3184) );
  AND2_X1 U23628 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n20688), .ZN(
        P1_U3185) );
  AND2_X1 U23629 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n20688), .ZN(P1_U3186) );
  AND2_X1 U23630 ( .A1(n20688), .A2(P1_DATAWIDTH_REG_8__SCAN_IN), .ZN(P1_U3187) );
  AND2_X1 U23631 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n20688), .ZN(P1_U3188) );
  AND2_X1 U23632 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n20688), .ZN(P1_U3189) );
  AND2_X1 U23633 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n20688), .ZN(P1_U3190) );
  AND2_X1 U23634 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n20688), .ZN(P1_U3191) );
  AND2_X1 U23635 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n20688), .ZN(P1_U3192) );
  AND2_X1 U23636 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n20688), .ZN(P1_U3193) );
  NAND2_X1 U23637 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n20689) );
  OAI211_X1 U23638 ( .C1(P1_STATE_REG_0__SCAN_IN), .C2(n20690), .A(
        P1_REQUESTPENDING_REG_SCAN_IN), .B(n20689), .ZN(n20691) );
  OAI21_X1 U23639 ( .B1(n20692), .B2(n20691), .A(n20740), .ZN(n20693) );
  OAI221_X1 U23640 ( .B1(P1_STATE_REG_2__SCAN_IN), .B2(P1_STATE_REG_0__SCAN_IN), .C1(P1_STATE_REG_2__SCAN_IN), .C2(n20695), .A(n20693), .ZN(P1_U3194) );
  NOR2_X1 U23641 ( .A1(NA), .A2(n20698), .ZN(n20694) );
  AOI21_X1 U23642 ( .B1(P1_REQUESTPENDING_REG_SCAN_IN), .B2(n20694), .A(
        P1_STATE_REG_2__SCAN_IN), .ZN(n20705) );
  NAND2_X1 U23643 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20796), .ZN(n20744) );
  OAI211_X1 U23644 ( .C1(P1_STATE_REG_0__SCAN_IN), .C2(NA), .A(n20695), .B(
        n20744), .ZN(n20696) );
  INV_X1 U23645 ( .A(n20696), .ZN(n20704) );
  NOR3_X1 U23646 ( .A1(NA), .A2(n20698), .A3(n20697), .ZN(n20700) );
  INV_X1 U23647 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20699) );
  OAI22_X1 U23648 ( .A1(n20701), .A2(n20700), .B1(P1_STATE_REG_2__SCAN_IN), 
        .B2(n20699), .ZN(n20702) );
  OAI22_X1 U23649 ( .A1(n20705), .A2(n20704), .B1(n20703), .B2(n20702), .ZN(
        P1_U3196) );
  NOR2_X1 U23650 ( .A1(n20783), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n20739) );
  INV_X1 U23651 ( .A(n20739), .ZN(n20748) );
  INV_X1 U23652 ( .A(n20744), .ZN(n20746) );
  AOI22_X1 U23653 ( .A1(P1_ADDRESS_REG_0__SCAN_IN), .A2(n20740), .B1(
        P1_REIP_REG_1__SCAN_IN), .B2(n20746), .ZN(n20706) );
  OAI21_X1 U23654 ( .B1(n20708), .B2(n20748), .A(n20706), .ZN(P1_U3197) );
  AOI22_X1 U23655 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(n20740), .B1(
        P1_REIP_REG_3__SCAN_IN), .B2(n20742), .ZN(n20707) );
  OAI21_X1 U23656 ( .B1(n20708), .B2(n20744), .A(n20707), .ZN(P1_U3198) );
  AOI222_X1 U23657 ( .A1(n20746), .A2(P1_REIP_REG_3__SCAN_IN), .B1(
        P1_ADDRESS_REG_2__SCAN_IN), .B2(n20783), .C1(P1_REIP_REG_4__SCAN_IN), 
        .C2(n20739), .ZN(n20709) );
  INV_X1 U23658 ( .A(n20709), .ZN(P1_U3199) );
  OAI222_X1 U23659 ( .A1(n20748), .A2(n20712), .B1(n20711), .B2(n20796), .C1(
        n20710), .C2(n20744), .ZN(P1_U3200) );
  AOI222_X1 U23660 ( .A1(n20746), .A2(P1_REIP_REG_5__SCAN_IN), .B1(
        P1_ADDRESS_REG_4__SCAN_IN), .B2(n20740), .C1(P1_REIP_REG_6__SCAN_IN), 
        .C2(n20739), .ZN(n20713) );
  INV_X1 U23661 ( .A(n20713), .ZN(P1_U3201) );
  AOI222_X1 U23662 ( .A1(n20746), .A2(P1_REIP_REG_6__SCAN_IN), .B1(
        P1_ADDRESS_REG_5__SCAN_IN), .B2(n20740), .C1(P1_REIP_REG_7__SCAN_IN), 
        .C2(n20742), .ZN(n20714) );
  INV_X1 U23663 ( .A(n20714), .ZN(P1_U3202) );
  AOI222_X1 U23664 ( .A1(n20746), .A2(P1_REIP_REG_7__SCAN_IN), .B1(
        P1_ADDRESS_REG_6__SCAN_IN), .B2(n20740), .C1(P1_REIP_REG_8__SCAN_IN), 
        .C2(n20742), .ZN(n20715) );
  INV_X1 U23665 ( .A(n20715), .ZN(P1_U3203) );
  AOI222_X1 U23666 ( .A1(n20746), .A2(P1_REIP_REG_8__SCAN_IN), .B1(
        P1_ADDRESS_REG_7__SCAN_IN), .B2(n20783), .C1(P1_REIP_REG_9__SCAN_IN), 
        .C2(n20742), .ZN(n20716) );
  INV_X1 U23667 ( .A(n20716), .ZN(P1_U3204) );
  AOI222_X1 U23668 ( .A1(n20746), .A2(P1_REIP_REG_9__SCAN_IN), .B1(
        P1_ADDRESS_REG_8__SCAN_IN), .B2(n20740), .C1(P1_REIP_REG_10__SCAN_IN), 
        .C2(n20742), .ZN(n20717) );
  INV_X1 U23669 ( .A(n20717), .ZN(P1_U3205) );
  AOI222_X1 U23670 ( .A1(n20746), .A2(P1_REIP_REG_10__SCAN_IN), .B1(
        P1_ADDRESS_REG_9__SCAN_IN), .B2(n20783), .C1(P1_REIP_REG_11__SCAN_IN), 
        .C2(n20742), .ZN(n20718) );
  INV_X1 U23671 ( .A(n20718), .ZN(P1_U3206) );
  AOI222_X1 U23672 ( .A1(n20742), .A2(P1_REIP_REG_12__SCAN_IN), .B1(
        P1_ADDRESS_REG_10__SCAN_IN), .B2(n20783), .C1(P1_REIP_REG_11__SCAN_IN), 
        .C2(n20746), .ZN(n20719) );
  INV_X1 U23673 ( .A(n20719), .ZN(P1_U3207) );
  AOI222_X1 U23674 ( .A1(n20746), .A2(P1_REIP_REG_12__SCAN_IN), .B1(
        P1_ADDRESS_REG_11__SCAN_IN), .B2(n20783), .C1(P1_REIP_REG_13__SCAN_IN), 
        .C2(n20742), .ZN(n20720) );
  INV_X1 U23675 ( .A(n20720), .ZN(P1_U3208) );
  AOI22_X1 U23676 ( .A1(P1_ADDRESS_REG_12__SCAN_IN), .A2(n20740), .B1(
        P1_REIP_REG_14__SCAN_IN), .B2(n20739), .ZN(n20721) );
  OAI21_X1 U23677 ( .B1(n20722), .B2(n20744), .A(n20721), .ZN(P1_U3209) );
  AOI22_X1 U23678 ( .A1(P1_ADDRESS_REG_13__SCAN_IN), .A2(n20783), .B1(
        P1_REIP_REG_14__SCAN_IN), .B2(n20746), .ZN(n20723) );
  OAI21_X1 U23679 ( .B1(n20724), .B2(n20748), .A(n20723), .ZN(P1_U3210) );
  AOI222_X1 U23680 ( .A1(n20746), .A2(P1_REIP_REG_15__SCAN_IN), .B1(
        P1_ADDRESS_REG_14__SCAN_IN), .B2(n20783), .C1(P1_REIP_REG_16__SCAN_IN), 
        .C2(n20742), .ZN(n20725) );
  INV_X1 U23681 ( .A(n20725), .ZN(P1_U3211) );
  AOI222_X1 U23682 ( .A1(n20746), .A2(P1_REIP_REG_16__SCAN_IN), .B1(
        P1_ADDRESS_REG_15__SCAN_IN), .B2(n20783), .C1(P1_REIP_REG_17__SCAN_IN), 
        .C2(n20742), .ZN(n20726) );
  INV_X1 U23683 ( .A(n20726), .ZN(P1_U3212) );
  AOI22_X1 U23684 ( .A1(P1_ADDRESS_REG_16__SCAN_IN), .A2(n20740), .B1(
        P1_REIP_REG_18__SCAN_IN), .B2(n20739), .ZN(n20727) );
  OAI21_X1 U23685 ( .B1(n20728), .B2(n20744), .A(n20727), .ZN(P1_U3213) );
  AOI222_X1 U23686 ( .A1(n20746), .A2(P1_REIP_REG_18__SCAN_IN), .B1(
        P1_ADDRESS_REG_17__SCAN_IN), .B2(n20783), .C1(P1_REIP_REG_19__SCAN_IN), 
        .C2(n20742), .ZN(n20729) );
  INV_X1 U23687 ( .A(n20729), .ZN(P1_U3214) );
  AOI222_X1 U23688 ( .A1(n20742), .A2(P1_REIP_REG_20__SCAN_IN), .B1(
        P1_ADDRESS_REG_18__SCAN_IN), .B2(n20740), .C1(P1_REIP_REG_19__SCAN_IN), 
        .C2(n20746), .ZN(n20730) );
  INV_X1 U23689 ( .A(n20730), .ZN(P1_U3215) );
  AOI222_X1 U23690 ( .A1(n20746), .A2(P1_REIP_REG_20__SCAN_IN), .B1(
        P1_ADDRESS_REG_19__SCAN_IN), .B2(n20740), .C1(P1_REIP_REG_21__SCAN_IN), 
        .C2(n20742), .ZN(n20731) );
  INV_X1 U23691 ( .A(n20731), .ZN(P1_U3216) );
  INV_X1 U23692 ( .A(P1_ADDRESS_REG_20__SCAN_IN), .ZN(n20999) );
  OAI222_X1 U23693 ( .A1(n20748), .A2(n20732), .B1(n20999), .B2(n20796), .C1(
        n14372), .C2(n20744), .ZN(P1_U3217) );
  AOI222_X1 U23694 ( .A1(n20746), .A2(P1_REIP_REG_22__SCAN_IN), .B1(
        P1_ADDRESS_REG_21__SCAN_IN), .B2(n20740), .C1(P1_REIP_REG_23__SCAN_IN), 
        .C2(n20742), .ZN(n20733) );
  INV_X1 U23695 ( .A(n20733), .ZN(P1_U3218) );
  AOI222_X1 U23696 ( .A1(n20746), .A2(P1_REIP_REG_23__SCAN_IN), .B1(
        P1_ADDRESS_REG_22__SCAN_IN), .B2(n20740), .C1(P1_REIP_REG_24__SCAN_IN), 
        .C2(n20742), .ZN(n20734) );
  INV_X1 U23697 ( .A(n20734), .ZN(P1_U3219) );
  AOI222_X1 U23698 ( .A1(n20746), .A2(P1_REIP_REG_24__SCAN_IN), .B1(
        P1_ADDRESS_REG_23__SCAN_IN), .B2(n20740), .C1(P1_REIP_REG_25__SCAN_IN), 
        .C2(n20739), .ZN(n20735) );
  INV_X1 U23699 ( .A(n20735), .ZN(P1_U3220) );
  AOI222_X1 U23700 ( .A1(n20746), .A2(P1_REIP_REG_25__SCAN_IN), .B1(
        P1_ADDRESS_REG_24__SCAN_IN), .B2(n20740), .C1(P1_REIP_REG_26__SCAN_IN), 
        .C2(n20739), .ZN(n20736) );
  INV_X1 U23701 ( .A(n20736), .ZN(P1_U3221) );
  AOI222_X1 U23702 ( .A1(n20746), .A2(P1_REIP_REG_26__SCAN_IN), .B1(
        P1_ADDRESS_REG_25__SCAN_IN), .B2(n20740), .C1(P1_REIP_REG_27__SCAN_IN), 
        .C2(n20739), .ZN(n20737) );
  INV_X1 U23703 ( .A(n20737), .ZN(P1_U3222) );
  AOI222_X1 U23704 ( .A1(n20746), .A2(P1_REIP_REG_27__SCAN_IN), .B1(
        P1_ADDRESS_REG_26__SCAN_IN), .B2(n20740), .C1(P1_REIP_REG_28__SCAN_IN), 
        .C2(n20742), .ZN(n20738) );
  INV_X1 U23705 ( .A(n20738), .ZN(P1_U3223) );
  AOI222_X1 U23706 ( .A1(n20746), .A2(P1_REIP_REG_28__SCAN_IN), .B1(
        P1_ADDRESS_REG_27__SCAN_IN), .B2(n20740), .C1(P1_REIP_REG_29__SCAN_IN), 
        .C2(n20739), .ZN(n20741) );
  INV_X1 U23707 ( .A(n20741), .ZN(P1_U3224) );
  AOI22_X1 U23708 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(n20742), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n20783), .ZN(n20743) );
  OAI21_X1 U23709 ( .B1(n20745), .B2(n20744), .A(n20743), .ZN(P1_U3225) );
  AOI22_X1 U23710 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(n20746), .B1(
        P1_ADDRESS_REG_29__SCAN_IN), .B2(n20783), .ZN(n20747) );
  OAI21_X1 U23711 ( .B1(n20749), .B2(n20748), .A(n20747), .ZN(P1_U3226) );
  OAI22_X1 U23712 ( .A1(n20783), .A2(P1_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P1_BE_N_REG_3__SCAN_IN), .B2(n20796), .ZN(n20750) );
  INV_X1 U23713 ( .A(n20750), .ZN(P1_U3458) );
  OAI22_X1 U23714 ( .A1(n20740), .A2(P1_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P1_BE_N_REG_2__SCAN_IN), .B2(n20796), .ZN(n20751) );
  INV_X1 U23715 ( .A(n20751), .ZN(P1_U3459) );
  OAI22_X1 U23716 ( .A1(n20740), .A2(P1_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P1_BE_N_REG_1__SCAN_IN), .B2(n20796), .ZN(n20752) );
  INV_X1 U23717 ( .A(n20752), .ZN(P1_U3460) );
  OAI22_X1 U23718 ( .A1(n20740), .A2(P1_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P1_BE_N_REG_0__SCAN_IN), .B2(n20796), .ZN(n20753) );
  INV_X1 U23719 ( .A(n20753), .ZN(P1_U3461) );
  OAI21_X1 U23720 ( .B1(P1_DATAWIDTH_REG_0__SCAN_IN), .B2(n20757), .A(n20755), 
        .ZN(n20754) );
  INV_X1 U23721 ( .A(n20754), .ZN(P1_U3464) );
  OAI21_X1 U23722 ( .B1(n20757), .B2(n20756), .A(n20755), .ZN(P1_U3465) );
  INV_X1 U23723 ( .A(n20771), .ZN(n20774) );
  NAND2_X1 U23724 ( .A1(n20759), .A2(n20758), .ZN(n20770) );
  AOI22_X1 U23725 ( .A1(n20763), .A2(n20762), .B1(n20761), .B2(n20760), .ZN(
        n20769) );
  NAND3_X1 U23726 ( .A1(n20766), .A2(n20765), .A3(n20764), .ZN(n20767) );
  AND4_X1 U23727 ( .A1(n20770), .A2(n20769), .A3(n20768), .A4(n20767), .ZN(
        n20772) );
  AOI22_X1 U23728 ( .A1(n20774), .A2(n20773), .B1(n20772), .B2(n20771), .ZN(
        P1_U3475) );
  AOI21_X1 U23729 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n20775) );
  AOI22_X1 U23730 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .B1(n20775), .B2(n13748), .ZN(n20777) );
  INV_X1 U23731 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n20776) );
  AOI22_X1 U23732 ( .A1(n20778), .A2(n20777), .B1(n20776), .B2(n20781), .ZN(
        P1_U3481) );
  INV_X1 U23733 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20782) );
  NOR2_X1 U23734 ( .A1(n20781), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n20779) );
  AOI22_X1 U23735 ( .A1(n20782), .A2(n20781), .B1(n20780), .B2(n20779), .ZN(
        P1_U3482) );
  AOI22_X1 U23736 ( .A1(n20796), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n20784), 
        .B2(n20783), .ZN(P1_U3483) );
  AOI211_X1 U23737 ( .C1(n20788), .C2(n20787), .A(n20786), .B(n20785), .ZN(
        n20795) );
  INV_X1 U23738 ( .A(n20789), .ZN(n20790) );
  OAI211_X1 U23739 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n11280), .A(n20790), 
        .B(P1_STATE2_REG_2__SCAN_IN), .ZN(n20792) );
  AOI21_X1 U23740 ( .B1(n20792), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n20791), 
        .ZN(n20794) );
  NAND2_X1 U23741 ( .A1(n20795), .A2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n20793) );
  OAI21_X1 U23742 ( .B1(n20795), .B2(n20794), .A(n20793), .ZN(P1_U3485) );
  OAI22_X1 U23743 ( .A1(n20740), .A2(P1_MEMORYFETCH_REG_SCAN_IN), .B1(
        P1_M_IO_N_REG_SCAN_IN), .B2(n20796), .ZN(n20797) );
  INV_X1 U23744 ( .A(n20797), .ZN(P1_U3486) );
  OR4_X1 U23745 ( .A1(keyinput63), .A2(keyinput21), .A3(keyinput98), .A4(
        keyinput56), .ZN(n20804) );
  INV_X1 U23746 ( .A(keyinput32), .ZN(n20798) );
  NAND4_X1 U23747 ( .A1(keyinput90), .A2(keyinput87), .A3(keyinput11), .A4(
        n20798), .ZN(n20803) );
  NOR2_X1 U23748 ( .A1(keyinput72), .A2(keyinput44), .ZN(n20799) );
  NAND3_X1 U23749 ( .A1(keyinput86), .A2(keyinput22), .A3(n20799), .ZN(n20802)
         );
  NOR2_X1 U23750 ( .A1(keyinput114), .A2(keyinput25), .ZN(n20800) );
  NAND3_X1 U23751 ( .A1(keyinput117), .A2(keyinput78), .A3(n20800), .ZN(n20801) );
  NOR4_X1 U23752 ( .A1(n20804), .A2(n20803), .A3(n20802), .A4(n20801), .ZN(
        n20826) );
  NOR2_X1 U23753 ( .A1(keyinput54), .A2(keyinput48), .ZN(n20805) );
  NAND3_X1 U23754 ( .A1(keyinput29), .A2(keyinput112), .A3(n20805), .ZN(n20809) );
  NAND4_X1 U23755 ( .A1(keyinput0), .A2(keyinput115), .A3(keyinput42), .A4(
        keyinput67), .ZN(n20808) );
  NAND4_X1 U23756 ( .A1(keyinput36), .A2(keyinput125), .A3(keyinput70), .A4(
        keyinput74), .ZN(n20807) );
  INV_X1 U23757 ( .A(keyinput88), .ZN(n21046) );
  NAND4_X1 U23758 ( .A1(keyinput85), .A2(keyinput34), .A3(keyinput66), .A4(
        n21046), .ZN(n20806) );
  NOR4_X1 U23759 ( .A1(n20809), .A2(n20808), .A3(n20807), .A4(n20806), .ZN(
        n20825) );
  NOR2_X1 U23760 ( .A1(keyinput79), .A2(keyinput124), .ZN(n20810) );
  NAND3_X1 U23761 ( .A1(keyinput105), .A2(keyinput53), .A3(n20810), .ZN(n20816) );
  INV_X1 U23762 ( .A(keyinput12), .ZN(n20811) );
  NAND4_X1 U23763 ( .A1(keyinput19), .A2(keyinput92), .A3(keyinput120), .A4(
        n20811), .ZN(n20815) );
  NAND4_X1 U23764 ( .A1(keyinput75), .A2(keyinput55), .A3(keyinput38), .A4(
        keyinput94), .ZN(n20814) );
  NOR2_X1 U23765 ( .A1(keyinput51), .A2(keyinput20), .ZN(n20812) );
  NAND3_X1 U23766 ( .A1(keyinput59), .A2(keyinput50), .A3(n20812), .ZN(n20813)
         );
  NOR4_X1 U23767 ( .A1(n20816), .A2(n20815), .A3(n20814), .A4(n20813), .ZN(
        n20824) );
  NOR4_X1 U23768 ( .A1(keyinput84), .A2(keyinput111), .A3(keyinput60), .A4(
        keyinput91), .ZN(n20822) );
  NOR4_X1 U23769 ( .A1(keyinput104), .A2(keyinput65), .A3(keyinput9), .A4(
        keyinput26), .ZN(n20821) );
  NAND2_X1 U23770 ( .A1(keyinput58), .A2(keyinput46), .ZN(n20817) );
  NOR3_X1 U23771 ( .A1(keyinput96), .A2(keyinput101), .A3(n20817), .ZN(n20820)
         );
  NAND2_X1 U23772 ( .A1(keyinput95), .A2(keyinput16), .ZN(n20818) );
  NOR3_X1 U23773 ( .A1(keyinput57), .A2(keyinput123), .A3(n20818), .ZN(n20819)
         );
  AND4_X1 U23774 ( .A1(n20822), .A2(n20821), .A3(n20820), .A4(n20819), .ZN(
        n20823) );
  NAND4_X1 U23775 ( .A1(n20826), .A2(n20825), .A3(n20824), .A4(n20823), .ZN(
        n20860) );
  NAND2_X1 U23776 ( .A1(keyinput17), .A2(keyinput15), .ZN(n20827) );
  NOR3_X1 U23777 ( .A1(keyinput40), .A2(keyinput77), .A3(n20827), .ZN(n20829)
         );
  INV_X1 U23778 ( .A(keyinput102), .ZN(n20828) );
  NAND4_X1 U23779 ( .A1(keyinput39), .A2(keyinput7), .A3(n20829), .A4(n20828), 
        .ZN(n20842) );
  NAND4_X1 U23780 ( .A1(keyinput23), .A2(keyinput82), .A3(keyinput30), .A4(
        keyinput68), .ZN(n20841) );
  NOR3_X1 U23781 ( .A1(keyinput108), .A2(keyinput106), .A3(keyinput64), .ZN(
        n20830) );
  NAND2_X1 U23782 ( .A1(keyinput52), .A2(n20830), .ZN(n20840) );
  NAND3_X1 U23783 ( .A1(keyinput1), .A2(keyinput71), .A3(keyinput100), .ZN(
        n20831) );
  NOR2_X1 U23784 ( .A1(keyinput4), .A2(n20831), .ZN(n20838) );
  INV_X1 U23785 ( .A(keyinput61), .ZN(n20832) );
  NOR4_X1 U23786 ( .A1(keyinput33), .A2(keyinput121), .A3(keyinput69), .A4(
        n20832), .ZN(n20837) );
  NAND2_X1 U23787 ( .A1(keyinput14), .A2(keyinput113), .ZN(n20833) );
  NOR3_X1 U23788 ( .A1(keyinput27), .A2(keyinput107), .A3(n20833), .ZN(n20836)
         );
  NAND2_X1 U23789 ( .A1(keyinput45), .A2(keyinput49), .ZN(n20834) );
  NOR3_X1 U23790 ( .A1(keyinput80), .A2(keyinput99), .A3(n20834), .ZN(n20835)
         );
  NAND4_X1 U23791 ( .A1(n20838), .A2(n20837), .A3(n20836), .A4(n20835), .ZN(
        n20839) );
  NOR4_X1 U23792 ( .A1(n20842), .A2(n20841), .A3(n20840), .A4(n20839), .ZN(
        n20858) );
  NOR4_X1 U23793 ( .A1(keyinput62), .A2(keyinput81), .A3(keyinput110), .A4(
        keyinput31), .ZN(n20857) );
  NAND3_X1 U23794 ( .A1(keyinput83), .A2(keyinput47), .A3(keyinput6), .ZN(
        n20843) );
  NOR2_X1 U23795 ( .A1(keyinput109), .A2(n20843), .ZN(n20856) );
  NAND2_X1 U23796 ( .A1(keyinput122), .A2(keyinput73), .ZN(n20844) );
  NOR3_X1 U23797 ( .A1(keyinput3), .A2(keyinput18), .A3(n20844), .ZN(n20845)
         );
  NAND3_X1 U23798 ( .A1(keyinput41), .A2(keyinput8), .A3(n20845), .ZN(n20854)
         );
  NAND2_X1 U23799 ( .A1(keyinput76), .A2(keyinput37), .ZN(n20846) );
  NOR3_X1 U23800 ( .A1(keyinput43), .A2(keyinput116), .A3(n20846), .ZN(n20852)
         );
  NAND2_X1 U23801 ( .A1(keyinput118), .A2(keyinput5), .ZN(n20847) );
  NOR3_X1 U23802 ( .A1(keyinput126), .A2(keyinput127), .A3(n20847), .ZN(n20851) );
  NAND2_X1 U23803 ( .A1(keyinput93), .A2(keyinput35), .ZN(n20848) );
  NOR3_X1 U23804 ( .A1(keyinput13), .A2(keyinput2), .A3(n20848), .ZN(n20850)
         );
  NOR4_X1 U23805 ( .A1(keyinput119), .A2(keyinput10), .A3(keyinput97), .A4(
        keyinput89), .ZN(n20849) );
  NAND4_X1 U23806 ( .A1(n20852), .A2(n20851), .A3(n20850), .A4(n20849), .ZN(
        n20853) );
  NOR4_X1 U23807 ( .A1(keyinput24), .A2(keyinput28), .A3(n20854), .A4(n20853), 
        .ZN(n20855) );
  NAND4_X1 U23808 ( .A1(n20858), .A2(n20857), .A3(n20856), .A4(n20855), .ZN(
        n20859) );
  OAI21_X1 U23809 ( .B1(n20860), .B2(n20859), .A(keyinput103), .ZN(n21125) );
  AOI22_X1 U23810 ( .A1(n20863), .A2(keyinput111), .B1(keyinput60), .B2(n20862), .ZN(n20861) );
  OAI221_X1 U23811 ( .B1(n20863), .B2(keyinput111), .C1(n20862), .C2(
        keyinput60), .A(n20861), .ZN(n20876) );
  AOI22_X1 U23812 ( .A1(n20866), .A2(keyinput26), .B1(keyinput84), .B2(n20865), 
        .ZN(n20864) );
  OAI221_X1 U23813 ( .B1(n20866), .B2(keyinput26), .C1(n20865), .C2(keyinput84), .A(n20864), .ZN(n20875) );
  INV_X1 U23814 ( .A(keyinput65), .ZN(n20868) );
  AOI22_X1 U23815 ( .A1(n20869), .A2(keyinput9), .B1(READY22_REG_SCAN_IN), 
        .B2(n20868), .ZN(n20867) );
  OAI221_X1 U23816 ( .B1(n20869), .B2(keyinput9), .C1(n20868), .C2(
        READY22_REG_SCAN_IN), .A(n20867), .ZN(n20874) );
  XOR2_X1 U23817 ( .A(n20870), .B(keyinput92), .Z(n20872) );
  XNOR2_X1 U23818 ( .A(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B(keyinput91), .ZN(
        n20871) );
  NAND2_X1 U23819 ( .A1(n20872), .A2(n20871), .ZN(n20873) );
  NOR4_X1 U23820 ( .A1(n20876), .A2(n20875), .A3(n20874), .A4(n20873), .ZN(
        n20924) );
  INV_X1 U23821 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n20879) );
  AOI22_X1 U23822 ( .A1(n20879), .A2(keyinput12), .B1(keyinput79), .B2(n20878), 
        .ZN(n20877) );
  OAI221_X1 U23823 ( .B1(n20879), .B2(keyinput12), .C1(n20878), .C2(keyinput79), .A(n20877), .ZN(n20890) );
  INV_X1 U23824 ( .A(keyinput105), .ZN(n20881) );
  AOI22_X1 U23825 ( .A1(n14408), .A2(keyinput124), .B1(P3_UWORD_REG_0__SCAN_IN), .B2(n20881), .ZN(n20880) );
  OAI221_X1 U23826 ( .B1(n14408), .B2(keyinput124), .C1(n20881), .C2(
        P3_UWORD_REG_0__SCAN_IN), .A(n20880), .ZN(n20889) );
  INV_X1 U23827 ( .A(keyinput120), .ZN(n20882) );
  XOR2_X1 U23828 ( .A(P3_EAX_REG_27__SCAN_IN), .B(n20882), .Z(n20885) );
  XNOR2_X1 U23829 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B(keyinput19), .ZN(
        n20884) );
  XNOR2_X1 U23830 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(keyinput53), 
        .ZN(n20883) );
  NAND3_X1 U23831 ( .A1(n20885), .A2(n20884), .A3(n20883), .ZN(n20888) );
  XNOR2_X1 U23832 ( .A(n20886), .B(keyinput59), .ZN(n20887) );
  NOR4_X1 U23833 ( .A1(n20890), .A2(n20889), .A3(n20888), .A4(n20887), .ZN(
        n20923) );
  INV_X1 U23834 ( .A(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n20893) );
  INV_X1 U23835 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n20892) );
  AOI22_X1 U23836 ( .A1(n20893), .A2(keyinput55), .B1(keyinput50), .B2(n20892), 
        .ZN(n20891) );
  OAI221_X1 U23837 ( .B1(n20893), .B2(keyinput55), .C1(n20892), .C2(keyinput50), .A(n20891), .ZN(n20905) );
  INV_X1 U23838 ( .A(keyinput75), .ZN(n20895) );
  AOI22_X1 U23839 ( .A1(n20896), .A2(keyinput51), .B1(P1_ADS_N_REG_SCAN_IN), 
        .B2(n20895), .ZN(n20894) );
  OAI221_X1 U23840 ( .B1(n20896), .B2(keyinput51), .C1(n20895), .C2(
        P1_ADS_N_REG_SCAN_IN), .A(n20894), .ZN(n20904) );
  INV_X1 U23841 ( .A(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n20899) );
  INV_X1 U23842 ( .A(keyinput57), .ZN(n20898) );
  AOI22_X1 U23843 ( .A1(n20899), .A2(keyinput94), .B1(P3_DATAO_REG_22__SCAN_IN), .B2(n20898), .ZN(n20897) );
  OAI221_X1 U23844 ( .B1(n20899), .B2(keyinput94), .C1(n20898), .C2(
        P3_DATAO_REG_22__SCAN_IN), .A(n20897), .ZN(n20903) );
  XNOR2_X1 U23845 ( .A(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B(keyinput38), .ZN(
        n20901) );
  XNOR2_X1 U23846 ( .A(keyinput20), .B(P2_EBX_REG_1__SCAN_IN), .ZN(n20900) );
  NAND2_X1 U23847 ( .A1(n20901), .A2(n20900), .ZN(n20902) );
  NOR4_X1 U23848 ( .A1(n20905), .A2(n20904), .A3(n20903), .A4(n20902), .ZN(
        n20922) );
  INV_X1 U23849 ( .A(keyinput16), .ZN(n20908) );
  INV_X1 U23850 ( .A(keyinput95), .ZN(n20907) );
  AOI22_X1 U23851 ( .A1(n20908), .A2(P2_DATAWIDTH_REG_15__SCAN_IN), .B1(
        P2_REQUESTPENDING_REG_SCAN_IN), .B2(n20907), .ZN(n20906) );
  OAI221_X1 U23852 ( .B1(n20908), .B2(P2_DATAWIDTH_REG_15__SCAN_IN), .C1(
        n20907), .C2(P2_REQUESTPENDING_REG_SCAN_IN), .A(n20906), .ZN(n20920)
         );
  INV_X1 U23853 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n20911) );
  INV_X1 U23854 ( .A(keyinput96), .ZN(n20910) );
  AOI22_X1 U23855 ( .A1(n20911), .A2(keyinput123), .B1(P1_LWORD_REG_8__SCAN_IN), .B2(n20910), .ZN(n20909) );
  OAI221_X1 U23856 ( .B1(n20911), .B2(keyinput123), .C1(n20910), .C2(
        P1_LWORD_REG_8__SCAN_IN), .A(n20909), .ZN(n20919) );
  INV_X1 U23857 ( .A(keyinput46), .ZN(n20914) );
  INV_X1 U23858 ( .A(keyinput101), .ZN(n20913) );
  AOI22_X1 U23859 ( .A1(n20914), .A2(P3_DATAO_REG_25__SCAN_IN), .B1(
        P3_DATAO_REG_7__SCAN_IN), .B2(n20913), .ZN(n20912) );
  OAI221_X1 U23860 ( .B1(n20914), .B2(P3_DATAO_REG_25__SCAN_IN), .C1(n20913), 
        .C2(P3_DATAO_REG_7__SCAN_IN), .A(n20912), .ZN(n20918) );
  INV_X1 U23861 ( .A(DATAI_19_), .ZN(n20916) );
  AOI22_X1 U23862 ( .A1(n20916), .A2(keyinput39), .B1(n10122), .B2(keyinput58), 
        .ZN(n20915) );
  OAI221_X1 U23863 ( .B1(n20916), .B2(keyinput39), .C1(n10122), .C2(keyinput58), .A(n20915), .ZN(n20917) );
  NOR4_X1 U23864 ( .A1(n20920), .A2(n20919), .A3(n20918), .A4(n20917), .ZN(
        n20921) );
  NAND4_X1 U23865 ( .A1(n20924), .A2(n20923), .A3(n20922), .A4(n20921), .ZN(
        n21124) );
  INV_X1 U23866 ( .A(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n20926) );
  AOI22_X1 U23867 ( .A1(n20927), .A2(keyinput18), .B1(n20926), .B2(keyinput24), 
        .ZN(n20925) );
  OAI221_X1 U23868 ( .B1(n20927), .B2(keyinput18), .C1(n20926), .C2(keyinput24), .A(n20925), .ZN(n20940) );
  INV_X1 U23869 ( .A(DATAI_24_), .ZN(n20930) );
  INV_X1 U23870 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n20929) );
  AOI22_X1 U23871 ( .A1(n20930), .A2(keyinput28), .B1(n20929), .B2(keyinput3), 
        .ZN(n20928) );
  OAI221_X1 U23872 ( .B1(n20930), .B2(keyinput28), .C1(n20929), .C2(keyinput3), 
        .A(n20928), .ZN(n20939) );
  INV_X1 U23873 ( .A(keyinput41), .ZN(n20932) );
  AOI22_X1 U23874 ( .A1(n20933), .A2(keyinput122), .B1(
        P3_BYTEENABLE_REG_1__SCAN_IN), .B2(n20932), .ZN(n20931) );
  OAI221_X1 U23875 ( .B1(n20933), .B2(keyinput122), .C1(n20932), .C2(
        P3_BYTEENABLE_REG_1__SCAN_IN), .A(n20931), .ZN(n20938) );
  AOI22_X1 U23876 ( .A1(n20936), .A2(keyinput8), .B1(keyinput6), .B2(n20935), 
        .ZN(n20934) );
  OAI221_X1 U23877 ( .B1(n20936), .B2(keyinput8), .C1(n20935), .C2(keyinput6), 
        .A(n20934), .ZN(n20937) );
  NOR4_X1 U23878 ( .A1(n20940), .A2(n20939), .A3(n20938), .A4(n20937), .ZN(
        n21122) );
  INV_X1 U23879 ( .A(keyinput13), .ZN(n20942) );
  AOI22_X1 U23880 ( .A1(n20943), .A2(keyinput10), .B1(P3_DATAO_REG_29__SCAN_IN), .B2(n20942), .ZN(n20941) );
  OAI221_X1 U23881 ( .B1(n20943), .B2(keyinput10), .C1(n20942), .C2(
        P3_DATAO_REG_29__SCAN_IN), .A(n20941), .ZN(n20956) );
  INV_X1 U23882 ( .A(keyinput35), .ZN(n20945) );
  AOI22_X1 U23883 ( .A1(n20946), .A2(keyinput97), .B1(
        P3_ADDRESS_REG_6__SCAN_IN), .B2(n20945), .ZN(n20944) );
  OAI221_X1 U23884 ( .B1(n20946), .B2(keyinput97), .C1(n20945), .C2(
        P3_ADDRESS_REG_6__SCAN_IN), .A(n20944), .ZN(n20955) );
  INV_X1 U23885 ( .A(keyinput2), .ZN(n20948) );
  AOI22_X1 U23886 ( .A1(n20949), .A2(keyinput89), .B1(P2_DATAO_REG_28__SCAN_IN), .B2(n20948), .ZN(n20947) );
  OAI221_X1 U23887 ( .B1(n20949), .B2(keyinput89), .C1(n20948), .C2(
        P2_DATAO_REG_28__SCAN_IN), .A(n20947), .ZN(n20954) );
  AOI22_X1 U23888 ( .A1(n20952), .A2(keyinput93), .B1(keyinput104), .B2(n20951), .ZN(n20950) );
  OAI221_X1 U23889 ( .B1(n20952), .B2(keyinput93), .C1(n20951), .C2(
        keyinput104), .A(n20950), .ZN(n20953) );
  NOR4_X1 U23890 ( .A1(n20956), .A2(n20955), .A3(n20954), .A4(n20953), .ZN(
        n21121) );
  AOI22_X1 U23891 ( .A1(n20959), .A2(keyinput81), .B1(n20958), .B2(keyinput110), .ZN(n20957) );
  OAI221_X1 U23892 ( .B1(n20959), .B2(keyinput81), .C1(n20958), .C2(
        keyinput110), .A(n20957), .ZN(n20988) );
  INV_X1 U23893 ( .A(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n20962) );
  INV_X1 U23894 ( .A(keyinput31), .ZN(n20961) );
  AOI22_X1 U23895 ( .A1(n20962), .A2(keyinput47), .B1(P1_BE_N_REG_3__SCAN_IN), 
        .B2(n20961), .ZN(n20960) );
  OAI221_X1 U23896 ( .B1(n20962), .B2(keyinput47), .C1(n20961), .C2(
        P1_BE_N_REG_3__SCAN_IN), .A(n20960), .ZN(n20987) );
  XOR2_X1 U23897 ( .A(keyinput109), .B(P2_DATAWIDTH_REG_4__SCAN_IN), .Z(n20966) );
  INV_X1 U23898 ( .A(keyinput5), .ZN(n20964) );
  AOI22_X1 U23899 ( .A1(n12548), .A2(keyinput83), .B1(P2_DATAO_REG_31__SCAN_IN), .B2(n20964), .ZN(n20963) );
  OAI221_X1 U23900 ( .B1(n12548), .B2(keyinput83), .C1(n20964), .C2(
        P2_DATAO_REG_31__SCAN_IN), .A(n20963), .ZN(n20965) );
  AOI211_X1 U23901 ( .C1(n20968), .C2(keyinput62), .A(n20966), .B(n20965), 
        .ZN(n20967) );
  OAI21_X1 U23902 ( .B1(n20968), .B2(keyinput62), .A(n20967), .ZN(n20986) );
  INV_X1 U23903 ( .A(keyinput126), .ZN(n20970) );
  OAI22_X1 U23904 ( .A1(keyinput127), .A2(n20971), .B1(n20970), .B2(
        P3_DATAWIDTH_REG_27__SCAN_IN), .ZN(n20969) );
  AOI221_X1 U23905 ( .B1(n20971), .B2(keyinput127), .C1(n20970), .C2(
        P3_DATAWIDTH_REG_27__SCAN_IN), .A(n20969), .ZN(n20984) );
  OAI22_X1 U23906 ( .A1(n20974), .A2(keyinput118), .B1(n20973), .B2(keyinput43), .ZN(n20972) );
  AOI221_X1 U23907 ( .B1(n20974), .B2(keyinput118), .C1(keyinput43), .C2(
        n20973), .A(n20972), .ZN(n20983) );
  INV_X1 U23908 ( .A(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n20977) );
  OAI22_X1 U23909 ( .A1(n20977), .A2(keyinput37), .B1(n20976), .B2(keyinput116), .ZN(n20975) );
  AOI221_X1 U23910 ( .B1(n20977), .B2(keyinput37), .C1(keyinput116), .C2(
        n20976), .A(n20975), .ZN(n20982) );
  INV_X1 U23911 ( .A(DATAI_5_), .ZN(n20980) );
  INV_X1 U23912 ( .A(keyinput119), .ZN(n20979) );
  OAI22_X1 U23913 ( .A1(n20980), .A2(keyinput76), .B1(n20979), .B2(
        P3_DATAWIDTH_REG_18__SCAN_IN), .ZN(n20978) );
  AOI221_X1 U23914 ( .B1(n20980), .B2(keyinput76), .C1(
        P3_DATAWIDTH_REG_18__SCAN_IN), .C2(n20979), .A(n20978), .ZN(n20981) );
  NAND4_X1 U23915 ( .A1(n20984), .A2(n20983), .A3(n20982), .A4(n20981), .ZN(
        n20985) );
  NOR4_X1 U23916 ( .A1(n20988), .A2(n20987), .A3(n20986), .A4(n20985), .ZN(
        n21120) );
  XOR2_X1 U23917 ( .A(keyinput15), .B(P2_LWORD_REG_0__SCAN_IN), .Z(n20993) );
  AOI22_X1 U23918 ( .A1(n20991), .A2(keyinput102), .B1(keyinput7), .B2(n20990), 
        .ZN(n20989) );
  OAI221_X1 U23919 ( .B1(n20991), .B2(keyinput102), .C1(n20990), .C2(keyinput7), .A(n20989), .ZN(n20992) );
  AOI211_X1 U23920 ( .C1(keyinput103), .C2(n20994), .A(n20993), .B(n20992), 
        .ZN(n21019) );
  INV_X1 U23921 ( .A(keyinput1), .ZN(n20996) );
  OAI22_X1 U23922 ( .A1(keyinput4), .A2(n20997), .B1(n20996), .B2(
        P2_DATAO_REG_27__SCAN_IN), .ZN(n20995) );
  AOI221_X1 U23923 ( .B1(n20997), .B2(keyinput4), .C1(n20996), .C2(
        P2_DATAO_REG_27__SCAN_IN), .A(n20995), .ZN(n21018) );
  OAI22_X1 U23924 ( .A1(n21000), .A2(keyinput100), .B1(n20999), .B2(keyinput80), .ZN(n20998) );
  AOI221_X1 U23925 ( .B1(n21000), .B2(keyinput100), .C1(keyinput80), .C2(
        n20999), .A(n20998), .ZN(n21017) );
  AOI22_X1 U23926 ( .A1(n21003), .A2(keyinput17), .B1(n21002), .B2(keyinput33), 
        .ZN(n21001) );
  OAI221_X1 U23927 ( .B1(n21003), .B2(keyinput17), .C1(n21002), .C2(keyinput33), .A(n21001), .ZN(n21015) );
  INV_X1 U23928 ( .A(DATAI_21_), .ZN(n21005) );
  AOI22_X1 U23929 ( .A1(n21005), .A2(keyinput77), .B1(n12180), .B2(keyinput40), 
        .ZN(n21004) );
  OAI221_X1 U23930 ( .B1(n21005), .B2(keyinput77), .C1(n12180), .C2(keyinput40), .A(n21004), .ZN(n21014) );
  INV_X1 U23931 ( .A(DATAI_22_), .ZN(n21008) );
  INV_X1 U23932 ( .A(keyinput69), .ZN(n21007) );
  AOI22_X1 U23933 ( .A1(n21008), .A2(keyinput71), .B1(P3_EAX_REG_19__SCAN_IN), 
        .B2(n21007), .ZN(n21006) );
  OAI221_X1 U23934 ( .B1(n21008), .B2(keyinput71), .C1(n21007), .C2(
        P3_EAX_REG_19__SCAN_IN), .A(n21006), .ZN(n21013) );
  INV_X1 U23935 ( .A(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n21010) );
  AOI22_X1 U23936 ( .A1(n21011), .A2(keyinput121), .B1(n21010), .B2(keyinput61), .ZN(n21009) );
  OAI221_X1 U23937 ( .B1(n21011), .B2(keyinput121), .C1(n21010), .C2(
        keyinput61), .A(n21009), .ZN(n21012) );
  NOR4_X1 U23938 ( .A1(n21015), .A2(n21014), .A3(n21013), .A4(n21012), .ZN(
        n21016) );
  NAND4_X1 U23939 ( .A1(n21019), .A2(n21018), .A3(n21017), .A4(n21016), .ZN(
        n21118) );
  INV_X1 U23940 ( .A(keyinput36), .ZN(n21021) );
  OAI22_X1 U23941 ( .A1(keyinput66), .A2(n21022), .B1(n21021), .B2(
        P3_DATAO_REG_27__SCAN_IN), .ZN(n21020) );
  AOI221_X1 U23942 ( .B1(n21022), .B2(keyinput66), .C1(n21021), .C2(
        P3_DATAO_REG_27__SCAN_IN), .A(n21020), .ZN(n21035) );
  INV_X1 U23943 ( .A(keyinput34), .ZN(n21024) );
  OAI22_X1 U23944 ( .A1(n21025), .A2(keyinput85), .B1(n21024), .B2(
        P1_UWORD_REG_0__SCAN_IN), .ZN(n21023) );
  AOI221_X1 U23945 ( .B1(n21025), .B2(keyinput85), .C1(P1_UWORD_REG_0__SCAN_IN), .C2(n21024), .A(n21023), .ZN(n21034) );
  INV_X1 U23946 ( .A(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n21028) );
  INV_X1 U23947 ( .A(keyinput87), .ZN(n21027) );
  OAI22_X1 U23948 ( .A1(n21028), .A2(keyinput74), .B1(n21027), .B2(
        P1_BE_N_REG_1__SCAN_IN), .ZN(n21026) );
  AOI221_X1 U23949 ( .B1(n21028), .B2(keyinput74), .C1(P1_BE_N_REG_1__SCAN_IN), 
        .C2(n21027), .A(n21026), .ZN(n21033) );
  INV_X1 U23950 ( .A(keyinput125), .ZN(n21030) );
  OAI22_X1 U23951 ( .A1(n21031), .A2(keyinput70), .B1(n21030), .B2(
        P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n21029) );
  AOI221_X1 U23952 ( .B1(n21031), .B2(keyinput70), .C1(
        P3_INSTQUEUE_REG_15__7__SCAN_IN), .C2(n21030), .A(n21029), .ZN(n21032)
         );
  NAND4_X1 U23953 ( .A1(n21035), .A2(n21034), .A3(n21033), .A4(n21032), .ZN(
        n21117) );
  INV_X1 U23954 ( .A(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n21038) );
  INV_X1 U23955 ( .A(keyinput67), .ZN(n21037) );
  OAI22_X1 U23956 ( .A1(n21038), .A2(keyinput54), .B1(n21037), .B2(
        P1_UWORD_REG_9__SCAN_IN), .ZN(n21036) );
  AOI221_X1 U23957 ( .B1(n21038), .B2(keyinput54), .C1(P1_UWORD_REG_9__SCAN_IN), .C2(n21037), .A(n21036), .ZN(n21051) );
  INV_X1 U23958 ( .A(P1_ADDRESS_REG_17__SCAN_IN), .ZN(n21041) );
  INV_X1 U23959 ( .A(keyinput42), .ZN(n21040) );
  OAI22_X1 U23960 ( .A1(n21041), .A2(keyinput115), .B1(n21040), .B2(
        P3_ADDRESS_REG_16__SCAN_IN), .ZN(n21039) );
  AOI221_X1 U23961 ( .B1(n21041), .B2(keyinput115), .C1(
        P3_ADDRESS_REG_16__SCAN_IN), .C2(n21040), .A(n21039), .ZN(n21050) );
  OAI22_X1 U23962 ( .A1(n21044), .A2(keyinput112), .B1(n21043), .B2(keyinput48), .ZN(n21042) );
  AOI221_X1 U23963 ( .B1(n21044), .B2(keyinput112), .C1(keyinput48), .C2(
        n21043), .A(n21042), .ZN(n21049) );
  INV_X1 U23964 ( .A(P1_LWORD_REG_1__SCAN_IN), .ZN(n21047) );
  OAI22_X1 U23965 ( .A1(keyinput29), .A2(n21047), .B1(n21046), .B2(
        P3_REIP_REG_1__SCAN_IN), .ZN(n21045) );
  AOI221_X1 U23966 ( .B1(n21047), .B2(keyinput29), .C1(n21046), .C2(
        P3_REIP_REG_1__SCAN_IN), .A(n21045), .ZN(n21048) );
  NAND4_X1 U23967 ( .A1(n21051), .A2(n21050), .A3(n21049), .A4(n21048), .ZN(
        n21116) );
  INV_X1 U23968 ( .A(keyinput106), .ZN(n21053) );
  AOI22_X1 U23969 ( .A1(n21054), .A2(keyinput82), .B1(
        P2_DATAWIDTH_REG_16__SCAN_IN), .B2(n21053), .ZN(n21052) );
  OAI221_X1 U23970 ( .B1(n21054), .B2(keyinput82), .C1(n21053), .C2(
        P2_DATAWIDTH_REG_16__SCAN_IN), .A(n21052), .ZN(n21065) );
  AOI22_X1 U23971 ( .A1(n13934), .A2(keyinput64), .B1(n21056), .B2(keyinput23), 
        .ZN(n21055) );
  OAI221_X1 U23972 ( .B1(n13934), .B2(keyinput64), .C1(n21056), .C2(keyinput23), .A(n21055), .ZN(n21064) );
  AOI22_X1 U23973 ( .A1(n21058), .A2(keyinput68), .B1(n12571), .B2(keyinput0), 
        .ZN(n21057) );
  OAI221_X1 U23974 ( .B1(n21058), .B2(keyinput68), .C1(n12571), .C2(keyinput0), 
        .A(n21057), .ZN(n21063) );
  INV_X1 U23975 ( .A(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n21061) );
  AOI22_X1 U23976 ( .A1(n21061), .A2(keyinput52), .B1(n21060), .B2(keyinput30), 
        .ZN(n21059) );
  OAI221_X1 U23977 ( .B1(n21061), .B2(keyinput52), .C1(n21060), .C2(keyinput30), .A(n21059), .ZN(n21062) );
  NOR4_X1 U23978 ( .A1(n21065), .A2(n21064), .A3(n21063), .A4(n21062), .ZN(
        n21114) );
  INV_X1 U23979 ( .A(keyinput14), .ZN(n21067) );
  AOI22_X1 U23980 ( .A1(n21068), .A2(keyinput27), .B1(P3_EAX_REG_16__SCAN_IN), 
        .B2(n21067), .ZN(n21066) );
  OAI221_X1 U23981 ( .B1(n21068), .B2(keyinput27), .C1(n21067), .C2(
        P3_EAX_REG_16__SCAN_IN), .A(n21066), .ZN(n21080) );
  AOI22_X1 U23982 ( .A1(n14731), .A2(keyinput107), .B1(keyinput108), .B2(
        n21070), .ZN(n21069) );
  OAI221_X1 U23983 ( .B1(n14731), .B2(keyinput107), .C1(n21070), .C2(
        keyinput108), .A(n21069), .ZN(n21079) );
  INV_X1 U23984 ( .A(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n21073) );
  INV_X1 U23985 ( .A(keyinput49), .ZN(n21072) );
  AOI22_X1 U23986 ( .A1(n21073), .A2(keyinput99), .B1(P2_DATAO_REG_23__SCAN_IN), .B2(n21072), .ZN(n21071) );
  OAI221_X1 U23987 ( .B1(n21073), .B2(keyinput99), .C1(n21072), .C2(
        P2_DATAO_REG_23__SCAN_IN), .A(n21071), .ZN(n21078) );
  XOR2_X1 U23988 ( .A(n21074), .B(keyinput113), .Z(n21076) );
  XNOR2_X1 U23989 ( .A(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B(keyinput45), .ZN(
        n21075) );
  NAND2_X1 U23990 ( .A1(n21076), .A2(n21075), .ZN(n21077) );
  NOR4_X1 U23991 ( .A1(n21080), .A2(n21079), .A3(n21078), .A4(n21077), .ZN(
        n21113) );
  INV_X1 U23992 ( .A(keyinput22), .ZN(n21082) );
  AOI22_X1 U23993 ( .A1(n21083), .A2(keyinput73), .B1(P2_UWORD_REG_6__SCAN_IN), 
        .B2(n21082), .ZN(n21081) );
  OAI221_X1 U23994 ( .B1(n21083), .B2(keyinput73), .C1(n21082), .C2(
        P2_UWORD_REG_6__SCAN_IN), .A(n21081), .ZN(n21095) );
  INV_X1 U23995 ( .A(keyinput78), .ZN(n21085) );
  AOI22_X1 U23996 ( .A1(n11511), .A2(keyinput117), .B1(
        P1_DATAWIDTH_REG_8__SCAN_IN), .B2(n21085), .ZN(n21084) );
  OAI221_X1 U23997 ( .B1(n11511), .B2(keyinput117), .C1(n21085), .C2(
        P1_DATAWIDTH_REG_8__SCAN_IN), .A(n21084), .ZN(n21094) );
  INV_X1 U23998 ( .A(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n21088) );
  INV_X1 U23999 ( .A(keyinput25), .ZN(n21087) );
  AOI22_X1 U24000 ( .A1(n21088), .A2(keyinput86), .B1(P1_UWORD_REG_12__SCAN_IN), .B2(n21087), .ZN(n21086) );
  OAI221_X1 U24001 ( .B1(n21088), .B2(keyinput86), .C1(n21087), .C2(
        P1_UWORD_REG_12__SCAN_IN), .A(n21086), .ZN(n21093) );
  INV_X1 U24002 ( .A(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n21089) );
  XOR2_X1 U24003 ( .A(n21089), .B(keyinput44), .Z(n21091) );
  XNOR2_X1 U24004 ( .A(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B(keyinput72), .ZN(
        n21090) );
  NAND2_X1 U24005 ( .A1(n21091), .A2(n21090), .ZN(n21092) );
  NOR4_X1 U24006 ( .A1(n21095), .A2(n21094), .A3(n21093), .A4(n21092), .ZN(
        n21112) );
  INV_X1 U24007 ( .A(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n21097) );
  AOI22_X1 U24008 ( .A1(n21097), .A2(keyinput21), .B1(keyinput98), .B2(n14276), 
        .ZN(n21096) );
  OAI221_X1 U24009 ( .B1(n21097), .B2(keyinput21), .C1(n14276), .C2(keyinput98), .A(n21096), .ZN(n21110) );
  INV_X1 U24010 ( .A(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n21099) );
  AOI22_X1 U24011 ( .A1(n21100), .A2(keyinput90), .B1(n21099), .B2(keyinput63), 
        .ZN(n21098) );
  OAI221_X1 U24012 ( .B1(n21100), .B2(keyinput90), .C1(n21099), .C2(keyinput63), .A(n21098), .ZN(n21109) );
  INV_X1 U24013 ( .A(keyinput11), .ZN(n21102) );
  AOI22_X1 U24014 ( .A1(n21103), .A2(keyinput114), .B1(
        P3_ADDRESS_REG_12__SCAN_IN), .B2(n21102), .ZN(n21101) );
  OAI221_X1 U24015 ( .B1(n21103), .B2(keyinput114), .C1(n21102), .C2(
        P3_ADDRESS_REG_12__SCAN_IN), .A(n21101), .ZN(n21108) );
  INV_X1 U24016 ( .A(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n21106) );
  INV_X1 U24017 ( .A(keyinput56), .ZN(n21105) );
  AOI22_X1 U24018 ( .A1(n21106), .A2(keyinput32), .B1(P1_LWORD_REG_0__SCAN_IN), 
        .B2(n21105), .ZN(n21104) );
  OAI221_X1 U24019 ( .B1(n21106), .B2(keyinput32), .C1(n21105), .C2(
        P1_LWORD_REG_0__SCAN_IN), .A(n21104), .ZN(n21107) );
  NOR4_X1 U24020 ( .A1(n21110), .A2(n21109), .A3(n21108), .A4(n21107), .ZN(
        n21111) );
  NAND4_X1 U24021 ( .A1(n21114), .A2(n21113), .A3(n21112), .A4(n21111), .ZN(
        n21115) );
  NOR4_X1 U24022 ( .A1(n21118), .A2(n21117), .A3(n21116), .A4(n21115), .ZN(
        n21119) );
  NAND4_X1 U24023 ( .A1(n21122), .A2(n21121), .A3(n21120), .A4(n21119), .ZN(
        n21123) );
  AOI211_X1 U24024 ( .C1(P1_DATAWIDTH_REG_13__SCAN_IN), .C2(n21125), .A(n21124), .B(n21123), .ZN(n21143) );
  INV_X1 U24025 ( .A(n21126), .ZN(n21129) );
  MUX2_X1 U24026 ( .A(n21129), .B(n21128), .S(n21127), .Z(n21136) );
  NAND2_X1 U24027 ( .A1(n12304), .A2(n21130), .ZN(n21131) );
  OAI211_X1 U24028 ( .C1(n21134), .C2(n21133), .A(n21132), .B(n21131), .ZN(
        n21135) );
  AOI211_X1 U24029 ( .C1(n21138), .C2(n21137), .A(n21136), .B(n21135), .ZN(
        n21139) );
  OAI21_X1 U24030 ( .B1(n21141), .B2(n21140), .A(n21139), .ZN(n21142) );
  XOR2_X1 U24031 ( .A(n21143), .B(n21142), .Z(P2_U3043) );
  AND2_X2 U11300 ( .A1(n11141), .A2(n11140), .ZN(n11228) );
  INV_X1 U11235 ( .A(n10480), .ZN(n12636) );
  AND2_X1 U13364 ( .A1(n12622), .A2(n10330), .ZN(n10658) );
  NAND2_X1 U11286 ( .A1(n9919), .A2(n10574), .ZN(n9953) );
  INV_X2 U11319 ( .A(n14352), .ZN(n11524) );
  INV_X2 U11315 ( .A(n19912), .ZN(n15726) );
  NAND2_X2 U11664 ( .A1(n10325), .A2(n10324), .ZN(n10511) );
  NOR2_X1 U11236 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10269) );
  CLKBUF_X1 U11256 ( .A(n11263), .Z(n13151) );
  CLKBUF_X1 U11302 ( .A(n13529), .Z(n9787) );
  CLKBUF_X1 U11329 ( .A(n12670), .Z(n20179) );
  XNOR2_X1 U11344 ( .A(n12458), .B(n12459), .ZN(n14719) );
  CLKBUF_X1 U11349 ( .A(n10441), .Z(n16218) );
  CLKBUF_X1 U11368 ( .A(n11821), .Z(n17027) );
  CLKBUF_X1 U11498 ( .A(n18125), .Z(n9817) );
  XNOR2_X1 U11577 ( .A(n14957), .B(n14959), .ZN(n14970) );
  CLKBUF_X1 U11589 ( .A(n16397), .Z(n16405) );
  CLKBUF_X1 U11712 ( .A(n11228), .Z(n12901) );
  CLKBUF_X1 U11938 ( .A(n17402), .Z(n17410) );
endmodule

