

module b15_C_AntiSAT_k_256_9 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, 
        keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, 
        keyinput133, keyinput134, keyinput135, keyinput136, keyinput137, 
        keyinput138, keyinput139, keyinput140, keyinput141, keyinput142, 
        keyinput143, keyinput144, keyinput145, keyinput146, keyinput147, 
        keyinput148, keyinput149, keyinput150, keyinput151, keyinput152, 
        keyinput153, keyinput154, keyinput155, keyinput156, keyinput157, 
        keyinput158, keyinput159, keyinput160, keyinput161, keyinput162, 
        keyinput163, keyinput164, keyinput165, keyinput166, keyinput167, 
        keyinput168, keyinput169, keyinput170, keyinput171, keyinput172, 
        keyinput173, keyinput174, keyinput175, keyinput176, keyinput177, 
        keyinput178, keyinput179, keyinput180, keyinput181, keyinput182, 
        keyinput183, keyinput184, keyinput185, keyinput186, keyinput187, 
        keyinput188, keyinput189, keyinput190, keyinput191, keyinput192, 
        keyinput193, keyinput194, keyinput195, keyinput196, keyinput197, 
        keyinput198, keyinput199, keyinput200, keyinput201, keyinput202, 
        keyinput203, keyinput204, keyinput205, keyinput206, keyinput207, 
        keyinput208, keyinput209, keyinput210, keyinput211, keyinput212, 
        keyinput213, keyinput214, keyinput215, keyinput216, keyinput217, 
        keyinput218, keyinput219, keyinput220, keyinput221, keyinput222, 
        keyinput223, keyinput224, keyinput225, keyinput226, keyinput227, 
        keyinput228, keyinput229, keyinput230, keyinput231, keyinput232, 
        keyinput233, keyinput234, keyinput235, keyinput236, keyinput237, 
        keyinput238, keyinput239, keyinput240, keyinput241, keyinput242, 
        keyinput243, keyinput244, keyinput245, keyinput246, keyinput247, 
        keyinput248, keyinput249, keyinput250, keyinput251, keyinput252, 
        keyinput253, keyinput254, keyinput255, U3445, U3446, U3447, U3448, 
        U3213, U3212, U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, 
        U3203, U3202, U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, 
        U3193, U3192, U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, 
        U3183, U3182, U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, 
        U3175, U3174, U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, 
        U3165, U3164, U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, 
        U3155, U3154, U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, 
        U3146, U3145, U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, 
        U3136, U3135, U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, 
        U3126, U3125, U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, 
        U3116, U3115, U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, 
        U3106, U3105, U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, 
        U3096, U3095, U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, 
        U3086, U3085, U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, 
        U3076, U3075, U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, 
        U3066, U3065, U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, 
        U3056, U3055, U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, 
        U3046, U3045, U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, 
        U3036, U3035, U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, 
        U3026, U3025, U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, 
        U3460, U3461, U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, 
        U3015, U3014, U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, 
        U3005, U3004, U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, 
        U2995, U2994, U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, 
        U2985, U2984, U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, 
        U2975, U2974, U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, 
        U2965, U2964, U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, 
        U2955, U2954, U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, 
        U2945, U2944, U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, 
        U2935, U2934, U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, 
        U2925, U2924, U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, 
        U2915, U2914, U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, 
        U2905, U2904, U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, 
        U2895, U2894, U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, 
        U2885, U2884, U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, 
        U2875, U2874, U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, 
        U2865, U2864, U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, 
        U2855, U2854, U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, 
        U2845, U2844, U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, 
        U2835, U2834, U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, 
        U2825, U2824, U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, 
        U2815, U2814, U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, 
        U2805, U2804, U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, 
        U2795, U3468, U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, 
        U3473, U2790, U2789, U3474, U2788 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1,
         keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7,
         keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13,
         keyinput14, keyinput15, keyinput16, keyinput17, keyinput18,
         keyinput19, keyinput20, keyinput21, keyinput22, keyinput23,
         keyinput24, keyinput25, keyinput26, keyinput27, keyinput28,
         keyinput29, keyinput30, keyinput31, keyinput32, keyinput33,
         keyinput34, keyinput35, keyinput36, keyinput37, keyinput38,
         keyinput39, keyinput40, keyinput41, keyinput42, keyinput43,
         keyinput44, keyinput45, keyinput46, keyinput47, keyinput48,
         keyinput49, keyinput50, keyinput51, keyinput52, keyinput53,
         keyinput54, keyinput55, keyinput56, keyinput57, keyinput58,
         keyinput59, keyinput60, keyinput61, keyinput62, keyinput63,
         keyinput64, keyinput65, keyinput66, keyinput67, keyinput68,
         keyinput69, keyinput70, keyinput71, keyinput72, keyinput73,
         keyinput74, keyinput75, keyinput76, keyinput77, keyinput78,
         keyinput79, keyinput80, keyinput81, keyinput82, keyinput83,
         keyinput84, keyinput85, keyinput86, keyinput87, keyinput88,
         keyinput89, keyinput90, keyinput91, keyinput92, keyinput93,
         keyinput94, keyinput95, keyinput96, keyinput97, keyinput98,
         keyinput99, keyinput100, keyinput101, keyinput102, keyinput103,
         keyinput104, keyinput105, keyinput106, keyinput107, keyinput108,
         keyinput109, keyinput110, keyinput111, keyinput112, keyinput113,
         keyinput114, keyinput115, keyinput116, keyinput117, keyinput118,
         keyinput119, keyinput120, keyinput121, keyinput122, keyinput123,
         keyinput124, keyinput125, keyinput126, keyinput127, keyinput128,
         keyinput129, keyinput130, keyinput131, keyinput132, keyinput133,
         keyinput134, keyinput135, keyinput136, keyinput137, keyinput138,
         keyinput139, keyinput140, keyinput141, keyinput142, keyinput143,
         keyinput144, keyinput145, keyinput146, keyinput147, keyinput148,
         keyinput149, keyinput150, keyinput151, keyinput152, keyinput153,
         keyinput154, keyinput155, keyinput156, keyinput157, keyinput158,
         keyinput159, keyinput160, keyinput161, keyinput162, keyinput163,
         keyinput164, keyinput165, keyinput166, keyinput167, keyinput168,
         keyinput169, keyinput170, keyinput171, keyinput172, keyinput173,
         keyinput174, keyinput175, keyinput176, keyinput177, keyinput178,
         keyinput179, keyinput180, keyinput181, keyinput182, keyinput183,
         keyinput184, keyinput185, keyinput186, keyinput187, keyinput188,
         keyinput189, keyinput190, keyinput191, keyinput192, keyinput193,
         keyinput194, keyinput195, keyinput196, keyinput197, keyinput198,
         keyinput199, keyinput200, keyinput201, keyinput202, keyinput203,
         keyinput204, keyinput205, keyinput206, keyinput207, keyinput208,
         keyinput209, keyinput210, keyinput211, keyinput212, keyinput213,
         keyinput214, keyinput215, keyinput216, keyinput217, keyinput218,
         keyinput219, keyinput220, keyinput221, keyinput222, keyinput223,
         keyinput224, keyinput225, keyinput226, keyinput227, keyinput228,
         keyinput229, keyinput230, keyinput231, keyinput232, keyinput233,
         keyinput234, keyinput235, keyinput236, keyinput237, keyinput238,
         keyinput239, keyinput240, keyinput241, keyinput242, keyinput243,
         keyinput244, keyinput245, keyinput246, keyinput247, keyinput248,
         keyinput249, keyinput250, keyinput251, keyinput252, keyinput253,
         keyinput254, keyinput255;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n3193, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203,
         n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213,
         n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223,
         n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233,
         n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243,
         n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253,
         n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263,
         n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273,
         n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283,
         n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293,
         n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303,
         n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313,
         n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323,
         n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333,
         n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343,
         n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353,
         n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363,
         n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373,
         n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383,
         n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393,
         n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403,
         n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413,
         n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423,
         n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433,
         n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443,
         n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453,
         n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463,
         n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473,
         n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483,
         n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493,
         n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503,
         n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513,
         n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523,
         n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533,
         n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543,
         n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553,
         n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563,
         n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
         n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583,
         n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593,
         n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603,
         n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613,
         n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
         n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633,
         n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
         n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653,
         n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663,
         n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673,
         n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683,
         n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693,
         n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703,
         n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713,
         n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723,
         n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733,
         n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743,
         n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753,
         n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763,
         n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773,
         n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783,
         n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793,
         n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803,
         n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813,
         n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823,
         n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833,
         n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843,
         n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853,
         n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863,
         n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873,
         n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883,
         n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893,
         n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903,
         n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913,
         n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923,
         n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933,
         n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943,
         n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953,
         n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963,
         n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973,
         n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983,
         n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993,
         n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003,
         n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013,
         n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023,
         n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033,
         n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043,
         n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053,
         n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063,
         n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073,
         n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083,
         n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093,
         n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103,
         n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113,
         n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123,
         n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133,
         n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143,
         n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153,
         n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163,
         n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173,
         n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183,
         n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193,
         n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203,
         n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213,
         n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223,
         n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233,
         n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243,
         n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253,
         n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263,
         n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273,
         n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283,
         n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293,
         n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303,
         n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313,
         n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323,
         n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333,
         n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343,
         n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353,
         n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363,
         n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373,
         n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383,
         n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393,
         n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403,
         n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413,
         n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423,
         n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433,
         n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443,
         n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453,
         n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463,
         n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473,
         n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483,
         n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493,
         n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503,
         n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
         n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
         n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
         n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
         n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
         n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
         n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613,
         n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623,
         n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
         n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643,
         n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653,
         n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663,
         n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673,
         n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683,
         n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693,
         n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703,
         n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713,
         n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723,
         n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733,
         n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743,
         n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753,
         n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763,
         n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773,
         n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783,
         n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793,
         n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803,
         n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813,
         n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823,
         n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833,
         n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843,
         n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853,
         n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863,
         n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873,
         n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883,
         n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893,
         n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903,
         n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913,
         n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923,
         n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933,
         n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943,
         n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953,
         n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963,
         n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973,
         n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983,
         n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993,
         n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003,
         n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013,
         n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023,
         n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033,
         n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043,
         n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053,
         n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063,
         n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073,
         n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
         n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104,
         n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114,
         n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124,
         n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
         n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144,
         n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154,
         n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164,
         n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174,
         n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184,
         n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194,
         n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204,
         n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214,
         n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224,
         n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234,
         n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244,
         n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
         n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264,
         n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274,
         n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284,
         n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294,
         n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304,
         n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314,
         n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324,
         n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334,
         n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344,
         n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354,
         n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364,
         n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374,
         n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384,
         n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394,
         n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404,
         n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414,
         n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424,
         n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434,
         n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444,
         n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5453, n5454, n5455,
         n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5465, n5466,
         n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476,
         n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486,
         n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496,
         n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506,
         n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516,
         n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526,
         n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536,
         n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546,
         n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556,
         n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566,
         n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576,
         n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586,
         n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596,
         n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606,
         n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616,
         n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626,
         n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636,
         n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646,
         n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656,
         n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666,
         n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676,
         n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686,
         n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696,
         n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706,
         n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716,
         n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726,
         n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736,
         n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746,
         n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756,
         n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766,
         n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776,
         n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786,
         n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796,
         n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806,
         n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816,
         n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826,
         n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836,
         n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846,
         n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856,
         n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866,
         n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876,
         n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886,
         n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896,
         n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906,
         n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916,
         n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926,
         n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936,
         n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946,
         n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956,
         n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966,
         n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976,
         n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986,
         n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996,
         n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006,
         n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016,
         n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026,
         n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036,
         n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046,
         n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056,
         n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066,
         n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076,
         n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086,
         n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096,
         n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106,
         n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116,
         n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126,
         n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136,
         n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146,
         n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156,
         n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166,
         n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176,
         n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186,
         n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196,
         n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206,
         n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216,
         n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226,
         n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236,
         n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246,
         n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256,
         n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266,
         n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276,
         n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286,
         n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296,
         n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306,
         n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316,
         n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326,
         n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336,
         n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346,
         n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356,
         n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366,
         n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376,
         n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386,
         n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6396, n6397,
         n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407,
         n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417,
         n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427,
         n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437,
         n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447,
         n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457,
         n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467,
         n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477,
         n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487,
         n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497,
         n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507,
         n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517,
         n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527,
         n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537,
         n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547,
         n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557,
         n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567,
         n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577,
         n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587,
         n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597,
         n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607,
         n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617,
         n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627,
         n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637,
         n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647,
         n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657,
         n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667,
         n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677,
         n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687,
         n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697,
         n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707,
         n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717,
         n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727,
         n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737,
         n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747,
         n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757,
         n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767,
         n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777,
         n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787,
         n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797,
         n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807,
         n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817,
         n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827,
         n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837,
         n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847,
         n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857,
         n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867,
         n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877,
         n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887,
         n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897,
         n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907,
         n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917,
         n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927,
         n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937,
         n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947,
         n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957,
         n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967,
         n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975;

  INV_X1 U3640 ( .A(n6967), .ZN(n6005) );
  INV_X1 U3641 ( .A(n5604), .ZN(n5592) );
  NAND2_X1 U3642 ( .A1(n3361), .A2(n3494), .ZN(n4470) );
  OR2_X1 U3643 ( .A1(n3518), .A2(n3517), .ZN(n4733) );
  BUF_X2 U3644 ( .A(n3571), .Z(n4156) );
  CLKBUF_X2 U3645 ( .A(n3573), .Z(n4158) );
  BUF_X2 U3646 ( .A(n3666), .Z(n4150) );
  CLKBUF_X2 U3647 ( .A(n3597), .Z(n4131) );
  CLKBUF_X2 U3648 ( .A(n3467), .Z(n3988) );
  CLKBUF_X2 U3649 ( .A(n3572), .Z(n4735) );
  CLKBUF_X2 U3650 ( .A(n3550), .Z(n4157) );
  CLKBUF_X2 U3651 ( .A(n3667), .Z(n3197) );
  BUF_X2 U3652 ( .A(n3198), .Z(n4148) );
  CLKBUF_X2 U3653 ( .A(n4050), .Z(n3943) );
  CLKBUF_X2 U3654 ( .A(n3584), .Z(n3896) );
  AND4_X1 U3655 ( .A1(n3248), .A2(n3247), .A3(n3246), .A4(n3245), .ZN(n3264)
         );
  AND2_X2 U3656 ( .A1(n3237), .A2(n5332), .ZN(n4049) );
  AND2_X1 U3657 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4722) );
  INV_X1 U3659 ( .A(n6974), .ZN(n3193) );
  INV_X2 U3661 ( .A(n6975), .ZN(n3195) );
  CLKBUF_X2 U3662 ( .A(n3544), .Z(n4160) );
  CLKBUF_X2 U3663 ( .A(n3443), .Z(n4055) );
  INV_X1 U3664 ( .A(n4171), .ZN(n3701) );
  OR2_X1 U3665 ( .A1(n3244), .A2(n3243), .ZN(n4208) );
  NAND2_X1 U3666 ( .A1(n5093), .A2(n4497), .ZN(n4496) );
  OR2_X1 U3667 ( .A1(n4584), .A2(n3623), .ZN(n3624) );
  AOI211_X1 U3668 ( .C1(n5652), .C2(n6227), .A(n4368), .B(n4367), .ZN(n4390)
         );
  CLKBUF_X3 U3669 ( .A(n3287), .Z(n3196) );
  AOI21_X2 U3671 ( .B1(n4547), .B2(n4548), .A(n4228), .ZN(n6149) );
  OR2_X2 U3675 ( .A1(n4331), .A2(n3218), .ZN(n4500) );
  AOI21_X2 U3676 ( .B1(n3498), .B2(n3497), .A(n3496), .ZN(n3499) );
  INV_X2 U3677 ( .A(n3527), .ZN(n3528) );
  NAND2_X2 U3679 ( .A1(n4289), .A2(n6091), .ZN(n5205) );
  AND2_X4 U3680 ( .A1(n3237), .A2(n4750), .ZN(n3852) );
  AND2_X4 U3681 ( .A1(n3231), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3237)
         );
  AND4_X2 U3683 ( .A1(n3272), .A2(n3271), .A3(n3270), .A4(n3269), .ZN(n3273)
         );
  AND4_X2 U3684 ( .A1(n3268), .A2(n3267), .A3(n3266), .A4(n3265), .ZN(n3274)
         );
  NAND2_X1 U3685 ( .A1(n3392), .A2(n3391), .ZN(n3485) );
  AND4_X2 U3686 ( .A1(n3390), .A2(n3389), .A3(n3388), .A4(n3387), .ZN(n3391)
         );
  AND4_X2 U3687 ( .A1(n3457), .A2(n3456), .A3(n3455), .A4(n3454), .ZN(n3229)
         );
  INV_X2 U3688 ( .A(n4208), .ZN(n4605) );
  AND4_X2 U3689 ( .A1(n3461), .A2(n3460), .A3(n3459), .A4(n3458), .ZN(n3221)
         );
  AND2_X4 U3690 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n5332) );
  AND2_X4 U3691 ( .A1(n4504), .A2(n4738), .ZN(n3584) );
  NOR2_X2 U3692 ( .A1(n5489), .A2(n5314), .ZN(n5310) );
  NAND2_X2 U3693 ( .A1(n4427), .A2(n4428), .ZN(n5489) );
  AOI21_X2 U3694 ( .B1(n5532), .B2(n5343), .A(n5342), .ZN(n5344) );
  OAI211_X2 U3695 ( .C1(n5363), .C2(n3529), .A(n4347), .B(n4334), .ZN(n3532)
         );
  NAND2_X1 U3696 ( .A1(n3561), .A2(n3562), .ZN(n3613) );
  CLKBUF_X1 U3697 ( .A(n3525), .Z(n5275) );
  CLKBUF_X2 U3698 ( .A(n3482), .Z(n4346) );
  CLKBUF_X2 U3699 ( .A(n4049), .Z(n4149) );
  NOR2_X4 U3700 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4738) );
  INV_X1 U3701 ( .A(n5252), .ZN(n5511) );
  CLKBUF_X1 U3702 ( .A(n5429), .Z(n5434) );
  CLKBUF_X1 U3703 ( .A(n3845), .Z(n5221) );
  NAND2_X1 U3704 ( .A1(n5142), .A2(n5192), .ZN(n5191) );
  NAND2_X1 U3705 ( .A1(n3727), .A2(n3726), .ZN(n4715) );
  NAND2_X1 U3706 ( .A1(n3760), .A2(n3759), .ZN(n5119) );
  XNOR2_X1 U3707 ( .A(n4249), .B(n6202), .ZN(n6129) );
  AND2_X1 U3708 ( .A1(n4233), .A2(n4232), .ZN(n6141) );
  OR2_X1 U3709 ( .A1(n3749), .A2(n3748), .ZN(n4283) );
  XNOR2_X1 U3710 ( .A(n4241), .B(n6802), .ZN(n6139) );
  NAND2_X1 U3711 ( .A1(n4240), .A2(n4239), .ZN(n4241) );
  CLKBUF_X1 U3712 ( .A(n5274), .Z(n6006) );
  NOR2_X1 U3713 ( .A1(n6890), .A2(n4807), .ZN(n6396) );
  NOR2_X1 U3714 ( .A1(n6968), .A2(n4807), .ZN(n6408) );
  NOR2_X1 U3715 ( .A1(n6065), .A2(n4807), .ZN(n6414) );
  NOR2_X1 U3716 ( .A1(n6060), .A2(n4807), .ZN(n6402) );
  NOR2_X1 U3717 ( .A1(n6067), .A2(n4807), .ZN(n6423) );
  NAND2_X1 U3718 ( .A1(n3640), .A2(n3639), .ZN(n4218) );
  NAND2_X1 U3719 ( .A1(n3658), .A2(n3657), .ZN(n4464) );
  OAI22_X1 U3720 ( .A1(n4499), .A2(STATE2_REG_0__SCAN_IN), .B1(n3616), .B2(
        n3615), .ZN(n3625) );
  NAND2_X1 U3721 ( .A1(n3665), .A2(n3664), .ZN(n6268) );
  NAND4_X1 U3722 ( .A1(n4356), .A2(n3522), .A3(n3521), .A4(n3520), .ZN(n3562)
         );
  AND4_X1 U3723 ( .A1(n4353), .A2(n3519), .A3(n4733), .A4(n6464), .ZN(n3520)
         );
  NAND2_X1 U3724 ( .A1(n4593), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3610) );
  BUF_X2 U3725 ( .A(n3493), .Z(n4555) );
  INV_X1 U3726 ( .A(n3482), .ZN(n4601) );
  AND2_X2 U3727 ( .A1(n3473), .A2(n3472), .ZN(n3205) );
  INV_X2 U3728 ( .A(n3622), .ZN(n3641) );
  NAND2_X1 U3729 ( .A1(n3473), .A2(n3472), .ZN(n3483) );
  AND2_X1 U3730 ( .A1(n3622), .A2(n3516), .ZN(n3525) );
  AND4_X1 U3731 ( .A1(n3471), .A2(n3470), .A3(n3469), .A4(n3468), .ZN(n3472)
         );
  AND4_X1 U3732 ( .A1(n3384), .A2(n3383), .A3(n3382), .A4(n3381), .ZN(n3392)
         );
  AND4_X1 U3733 ( .A1(n3375), .A2(n3374), .A3(n3373), .A4(n3372), .ZN(n3380)
         );
  AND4_X1 U3734 ( .A1(n3447), .A2(n3446), .A3(n3445), .A4(n3444), .ZN(n3453)
         );
  AND2_X1 U3735 ( .A1(n3206), .A2(n3207), .ZN(n3468) );
  AND4_X1 U3736 ( .A1(n3466), .A2(n3465), .A3(n3464), .A4(n3463), .ZN(n3473)
         );
  AND4_X1 U3737 ( .A1(n3256), .A2(n3255), .A3(n3254), .A4(n3253), .ZN(n3262)
         );
  AND2_X1 U3738 ( .A1(n3571), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3386) );
  BUF_X2 U3739 ( .A(n3545), .Z(n4159) );
  AND2_X2 U3740 ( .A1(n4505), .A2(n4722), .ZN(n3597) );
  AND2_X2 U3741 ( .A1(n3393), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4505)
         );
  INV_X1 U3742 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3393) );
  BUF_X1 U3743 ( .A(n3566), .Z(n3198) );
  OR3_X1 U3744 ( .A1(n4438), .A2(n4440), .A3(n4439), .ZN(n3199) );
  OR2_X1 U3745 ( .A1(n4441), .A2(n3199), .ZN(U2992) );
  NAND2_X2 U3746 ( .A1(n3620), .A2(n3619), .ZN(n3200) );
  OAI21_X1 U3747 ( .B1(n5627), .B2(n4299), .A(n4298), .ZN(n3201) );
  OAI21_X1 U3749 ( .B1(n5627), .B2(n4299), .A(n4298), .ZN(n5286) );
  XNOR2_X1 U3750 ( .A(n3200), .B(n4586), .ZN(n4234) );
  NAND2_X1 U3751 ( .A1(n4303), .A2(n3223), .ZN(n5248) );
  NAND2_X1 U3752 ( .A1(n3392), .A2(n3391), .ZN(n3203) );
  NAND2_X1 U3753 ( .A1(n3392), .A2(n3391), .ZN(n3204) );
  NAND2_X1 U3754 ( .A1(n3667), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3206) );
  NAND2_X1 U3755 ( .A1(n3566), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3207)
         );
  AND2_X2 U3756 ( .A1(n3238), .A2(n5332), .ZN(n3667) );
  AND2_X2 U3757 ( .A1(n4722), .A2(n4504), .ZN(n3566) );
  NAND2_X1 U3758 ( .A1(n3505), .A2(n3504), .ZN(n3561) );
  INV_X1 U3759 ( .A(n3485), .ZN(n3208) );
  INV_X1 U3760 ( .A(n3485), .ZN(n4678) );
  NAND2_X1 U3761 ( .A1(n6108), .A2(n6107), .ZN(n6106) );
  OR2_X2 U3762 ( .A1(n5292), .A2(n5440), .ZN(n5442) );
  NOR2_X2 U3763 ( .A1(n4582), .A2(n3301), .ZN(n4640) );
  NOR2_X4 U3764 ( .A1(n5442), .A2(n5437), .ZN(n5436) );
  AOI211_X2 U3765 ( .C1(n4340), .C2(n4339), .A(n4341), .B(n4338), .ZN(n4344)
         );
  NAND2_X1 U3766 ( .A1(n6106), .A2(n4279), .ZN(n3209) );
  NAND2_X1 U3767 ( .A1(n6129), .A2(n6131), .ZN(n3210) );
  NAND3_X1 U3768 ( .A1(n3537), .A2(n3536), .A3(n3535), .ZN(n3211) );
  NOR2_X1 U3771 ( .A1(n5488), .A2(n5534), .ZN(n5342) );
  NOR4_X1 U3772 ( .A1(n5488), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_30__SCAN_IN), .A4(n5534), .ZN(n5309) );
  XNOR2_X1 U3773 ( .A(n3214), .B(n5311), .ZN(n3222) );
  INV_X1 U3774 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n3214) );
  NAND2_X1 U3775 ( .A1(n5590), .A2(n5249), .ZN(n3215) );
  NAND2_X1 U3776 ( .A1(n5590), .A2(n5249), .ZN(n5496) );
  NAND2_X1 U3777 ( .A1(n6141), .A2(n6139), .ZN(n3216) );
  NAND2_X1 U3778 ( .A1(n4601), .A2(n3204), .ZN(n4331) );
  AND2_X1 U3779 ( .A1(n3237), .A2(n5332), .ZN(n3217) );
  AND2_X2 U3780 ( .A1(n5429), .A2(n4023), .ZN(n5266) );
  NOR2_X2 U3781 ( .A1(n5433), .A2(n5435), .ZN(n5429) );
  NOR2_X1 U3782 ( .A1(n5770), .A2(n5771), .ZN(n5769) );
  NAND2_X2 U3783 ( .A1(n5248), .A2(n4305), .ZN(n5589) );
  NAND2_X1 U3784 ( .A1(n4208), .A2(n3205), .ZN(n4354) );
  OAI22_X2 U3785 ( .A1(n5498), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .B1(n5504), .B2(n5253), .ZN(n5254) );
  NAND2_X1 U3786 ( .A1(n4314), .A2(n3474), .ZN(n4323) );
  NAND2_X4 U3787 ( .A1(n3229), .A2(n3221), .ZN(n3516) );
  NOR2_X2 U3788 ( .A1(n5430), .A2(n5418), .ZN(n5417) );
  NAND2_X1 U3789 ( .A1(n4248), .A2(n4247), .ZN(n4249) );
  OAI21_X2 U3790 ( .B1(n5770), .B2(n5771), .A(n4311), .ZN(n4312) );
  NAND2_X2 U3791 ( .A1(n4310), .A2(n4309), .ZN(n5770) );
  OAI21_X2 U3792 ( .B1(n5228), .B2(n5231), .A(n5229), .ZN(n5798) );
  OAI21_X2 U3793 ( .B1(n6083), .B2(n4293), .A(n4292), .ZN(n5228) );
  NAND2_X1 U3794 ( .A1(n4208), .A2(n3401), .ZN(n3218) );
  NAND2_X1 U3795 ( .A1(n4208), .A2(n3401), .ZN(n3219) );
  INV_X1 U3796 ( .A(n3494), .ZN(n5419) );
  XNOR2_X2 U3798 ( .A(n3560), .B(n3559), .ZN(n3620) );
  NAND2_X1 U3799 ( .A1(n3688), .A2(n4586), .ZN(n3728) );
  NAND2_X1 U3800 ( .A1(n3700), .A2(n3699), .ZN(n3731) );
  AOI21_X1 U3801 ( .B1(n4589), .B2(n6567), .A(n3557), .ZN(n3560) );
  OR2_X1 U3802 ( .A1(n3506), .A2(n3524), .ZN(n4356) );
  NAND2_X1 U3803 ( .A1(n3592), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3615) );
  NAND2_X1 U3804 ( .A1(n3744), .A2(n4269), .ZN(n3431) );
  NOR2_X2 U3805 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n4176) );
  INV_X1 U3806 ( .A(n4176), .ZN(n4145) );
  INV_X1 U3807 ( .A(n3431), .ZN(n3438) );
  CLKBUF_X1 U3808 ( .A(n3527), .Z(n5354) );
  NAND2_X1 U3809 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n5953), .ZN(n5080) );
  OR2_X1 U3810 ( .A1(n5364), .A2(n6461), .ZN(n4551) );
  INV_X1 U3811 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6564) );
  NAND2_X1 U3812 ( .A1(n4537), .A2(n4208), .ZN(n3514) );
  CLKBUF_X1 U3813 ( .A(n3852), .Z(n4151) );
  NAND2_X1 U3814 ( .A1(n3733), .A2(n3732), .ZN(n3749) );
  AND2_X1 U3815 ( .A1(n3731), .A2(n3730), .ZN(n3732) );
  INV_X1 U3816 ( .A(n3728), .ZN(n3733) );
  OR2_X1 U3817 ( .A1(n3677), .A2(n3676), .ZN(n4244) );
  NAND2_X1 U3818 ( .A1(n4593), .A2(n3401), .ZN(n5081) );
  AND3_X1 U3819 ( .A1(n4503), .A2(n4360), .A3(n4501), .ZN(n4362) );
  NAND2_X1 U3820 ( .A1(n5451), .A2(n5450), .ZN(n5300) );
  NOR2_X2 U3821 ( .A1(n5191), .A2(n5222), .ZN(n3845) );
  NOR2_X1 U3822 ( .A1(n4715), .A2(n4716), .ZN(n4714) );
  INV_X1 U3823 ( .A(n4579), .ZN(n3709) );
  NOR2_X2 U3824 ( .A1(n3622), .A2(n5155), .ZN(n3873) );
  NOR2_X2 U3825 ( .A1(n5382), .A2(n5381), .ZN(n5371) );
  NAND2_X1 U3826 ( .A1(n4208), .A2(n3401), .ZN(n3494) );
  INV_X1 U3827 ( .A(n3636), .ZN(n3637) );
  NAND2_X1 U3828 ( .A1(n3532), .A2(n3531), .ZN(n3611) );
  AND2_X1 U3829 ( .A1(n3530), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3531) );
  NAND2_X1 U3830 ( .A1(n3528), .A2(n4702), .ZN(n4334) );
  INV_X1 U3831 ( .A(n4807), .ZN(n4845) );
  OAI21_X1 U3832 ( .B1(n6471), .B2(n4760), .A(n5327), .ZN(n4592) );
  INV_X1 U3833 ( .A(n5953), .ZN(n5103) );
  AND2_X1 U3834 ( .A1(n4362), .A2(n4361), .ZN(n5357) );
  NOR2_X2 U3835 ( .A1(n5375), .A2(n4406), .ZN(n4407) );
  AND2_X1 U3836 ( .A1(n5266), .A2(n5279), .ZN(n5378) );
  AND2_X1 U3837 ( .A1(n4102), .A2(n4101), .ZN(n5267) );
  AND2_X1 U3838 ( .A1(n3911), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n3975)
         );
  NOR2_X2 U3839 ( .A1(n5300), .A2(n5302), .ZN(n5301) );
  NAND2_X1 U3840 ( .A1(n3832), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3849)
         );
  NOR2_X1 U3841 ( .A1(n3801), .A2(n5935), .ZN(n3804) );
  NAND2_X1 U3842 ( .A1(n4714), .A2(n5119), .ZN(n5117) );
  NOR2_X2 U3843 ( .A1(n5137), .A2(n5126), .ZN(n5200) );
  AND2_X1 U3844 ( .A1(n4330), .A2(n4329), .ZN(n4370) );
  XNOR2_X1 U3845 ( .A(n3627), .B(n3626), .ZN(n3628) );
  OR2_X1 U3846 ( .A1(n5354), .A2(n4702), .ZN(n4731) );
  NAND2_X1 U3847 ( .A1(n3442), .A2(n3441), .ZN(n5364) );
  NAND2_X1 U3848 ( .A1(n3478), .A2(n3750), .ZN(n3441) );
  CLKBUF_X1 U3849 ( .A(n4334), .Z(n4719) );
  NOR2_X1 U3850 ( .A1(n4688), .A2(n4765), .ZN(n4697) );
  CLKBUF_X1 U3851 ( .A(n3202), .Z(n4857) );
  NAND2_X1 U3852 ( .A1(n6567), .A2(n4592), .ZN(n4807) );
  INV_X1 U3853 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6567) );
  NAND2_X1 U3854 ( .A1(REIP_REG_18__SCAN_IN), .A2(n5852), .ZN(n5736) );
  INV_X1 U3855 ( .A(n5967), .ZN(n5952) );
  OR2_X1 U3856 ( .A1(n3196), .A2(n3489), .ZN(n5969) );
  INV_X1 U3857 ( .A(n5983), .ZN(n5970) );
  INV_X1 U3858 ( .A(n5964), .ZN(n5990) );
  AND2_X1 U3859 ( .A1(n4420), .A2(n4419), .ZN(n5982) );
  INV_X1 U3860 ( .A(n5969), .ZN(n5981) );
  AND2_X1 U3861 ( .A1(n5320), .A2(n4414), .ZN(n5964) );
  NOR2_X2 U3862 ( .A1(n5103), .A2(n6547), .ZN(n5983) );
  INV_X1 U3863 ( .A(n5453), .ZN(n5462) );
  AND2_X1 U3864 ( .A1(n5453), .A2(n5468), .ZN(n5445) );
  AND2_X1 U3865 ( .A1(n5791), .A2(n4396), .ZN(n6134) );
  INV_X1 U3866 ( .A(n5831), .ZN(n6152) );
  OR2_X1 U3867 ( .A1(n4551), .A2(n6444), .ZN(n5831) );
  INV_X1 U3868 ( .A(n5815), .ZN(n6231) );
  INV_X1 U3869 ( .A(n4218), .ZN(n4866) );
  INV_X1 U3870 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6441) );
  NAND2_X1 U3871 ( .A1(n3506), .A2(n4702), .ZN(n3498) );
  NOR2_X1 U3872 ( .A1(n4331), .A2(n4555), .ZN(n3511) );
  AND2_X1 U3873 ( .A1(n3426), .A2(n3425), .ZN(n3428) );
  AOI22_X1 U3874 ( .A1(n4049), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3852), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3447) );
  AND2_X2 U3875 ( .A1(n3237), .A2(n4505), .ZN(n3666) );
  OR2_X1 U3876 ( .A1(n3743), .A2(n3742), .ZN(n4272) );
  OR2_X1 U3877 ( .A1(n3698), .A2(n3697), .ZN(n4261) );
  OR2_X1 U3878 ( .A1(n3515), .A2(n4345), .ZN(n3519) );
  AOI22_X1 U3879 ( .A1(n3666), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3550), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3465) );
  AOI22_X1 U3880 ( .A1(n4050), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3443), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3265) );
  AOI22_X1 U3881 ( .A1(n3573), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3584), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3268) );
  AND2_X1 U3882 ( .A1(n5407), .A2(n5412), .ZN(n5401) );
  NAND2_X1 U3883 ( .A1(n5301), .A2(n5444), .ZN(n5433) );
  INV_X1 U3884 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3848) );
  OR2_X1 U3885 ( .A1(n3590), .A2(n3589), .ZN(n4220) );
  NAND2_X1 U3886 ( .A1(n3679), .A2(n3678), .ZN(n4586) );
  NAND2_X1 U3887 ( .A1(n3621), .A2(n3200), .ZN(n4584) );
  AND2_X2 U3888 ( .A1(n4722), .A2(n5332), .ZN(n3572) );
  AND4_X1 U3889 ( .A1(n4358), .A2(n4357), .A3(n4356), .A4(n4355), .ZN(n4503)
         );
  NAND2_X1 U3890 ( .A1(n3615), .A2(n3610), .ZN(n3750) );
  AND2_X1 U3891 ( .A1(n3481), .A2(n3752), .ZN(n3433) );
  OR2_X1 U3892 ( .A1(n5084), .A2(n4767), .ZN(n4858) );
  INV_X1 U3893 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4859) );
  AND2_X1 U3894 ( .A1(n3540), .A2(n4950), .ZN(n4652) );
  XNOR2_X1 U3895 ( .A(n4464), .B(n6268), .ZN(n4588) );
  AND2_X1 U3896 ( .A1(n4316), .A2(n4317), .ZN(n4333) );
  INV_X1 U3897 ( .A(n4323), .ZN(n3475) );
  OR2_X1 U3898 ( .A1(n4512), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4392) );
  INV_X1 U3899 ( .A(n5976), .ZN(n5986) );
  INV_X1 U3900 ( .A(n4472), .ZN(n3281) );
  INV_X1 U3901 ( .A(n3283), .ZN(n3282) );
  OR2_X1 U3902 ( .A1(n6569), .A2(n3488), .ZN(n5953) );
  INV_X1 U3903 ( .A(n5371), .ZN(n5384) );
  AND2_X1 U3904 ( .A1(n3354), .A2(n3353), .ZN(n5256) );
  AND2_X1 U3905 ( .A1(n3331), .A2(n3330), .ZN(n5440) );
  AND2_X1 U3906 ( .A1(n3319), .A2(n3318), .ZN(n5225) );
  NAND2_X1 U3907 ( .A1(n4125), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4181)
         );
  NOR2_X1 U3908 ( .A1(n4092), .A2(n5265), .ZN(n4086) );
  NAND2_X1 U3909 ( .A1(PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n4086), .ZN(n4085)
         );
  NAND2_X1 U3910 ( .A1(n3976), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4092)
         );
  NOR2_X1 U3911 ( .A1(n3959), .A2(n5733), .ZN(n3911) );
  NOR2_X1 U3912 ( .A1(n4007), .A2(n3910), .ZN(n3960) );
  NOR2_X1 U3913 ( .A1(n3894), .A2(n5870), .ZN(n3895) );
  NAND2_X1 U3914 ( .A1(PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n3895), .ZN(n4007)
         );
  NAND2_X1 U3916 ( .A1(PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n3877), .ZN(n3894)
         );
  OR2_X1 U3917 ( .A1(n3849), .A2(n3848), .ZN(n3850) );
  INV_X1 U3918 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3851) );
  NOR2_X1 U3919 ( .A1(n3851), .A2(n3850), .ZN(n3877) );
  NAND2_X1 U3920 ( .A1(n5460), .A2(n3847), .ZN(n5451) );
  NAND2_X1 U3921 ( .A1(n5458), .A2(n5459), .ZN(n5460) );
  NOR2_X1 U3922 ( .A1(n3829), .A2(n3828), .ZN(n3832) );
  NAND2_X1 U3923 ( .A1(n3804), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3829)
         );
  CLKBUF_X1 U3924 ( .A(n5142), .Z(n5193) );
  INV_X1 U3925 ( .A(n3776), .ZN(n3777) );
  NOR2_X1 U3926 ( .A1(n3755), .A2(n3754), .ZN(n3756) );
  INV_X1 U3927 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3754) );
  INV_X1 U3928 ( .A(n4578), .ZN(n3727) );
  AOI21_X1 U3929 ( .B1(n4259), .B2(n3873), .A(n3747), .ZN(n4716) );
  CLKBUF_X1 U3930 ( .A(n4714), .Z(n5120) );
  NAND2_X1 U3931 ( .A1(n3723), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3755)
         );
  NOR2_X1 U3932 ( .A1(n6897), .A2(n3705), .ZN(n3723) );
  INV_X1 U3933 ( .A(n3680), .ZN(n3681) );
  NAND2_X1 U3934 ( .A1(PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n3680) );
  NAND2_X1 U3935 ( .A1(n4495), .A2(n3651), .ZN(n4542) );
  INV_X1 U3936 ( .A(n5372), .ZN(n3364) );
  OR2_X1 U3937 ( .A1(n5255), .A2(n5256), .ZN(n5392) );
  NOR2_X2 U3938 ( .A1(n5392), .A2(n5391), .ZN(n5390) );
  BUF_X1 U3940 ( .A(n5603), .Z(n5785) );
  AND2_X1 U3941 ( .A1(n3316), .A2(n3315), .ZN(n5196) );
  INV_X1 U3942 ( .A(n4632), .ZN(n5289) );
  AND2_X1 U3943 ( .A1(n3309), .A2(n3308), .ZN(n5136) );
  NAND2_X1 U3944 ( .A1(n3294), .A2(n3293), .ZN(n4582) );
  AND2_X1 U3945 ( .A1(n4575), .A2(n4574), .ZN(n3293) );
  OR2_X1 U3946 ( .A1(n4370), .A2(n4724), .ZN(n4382) );
  NAND2_X1 U3947 ( .A1(n3638), .A2(n3637), .ZN(n3639) );
  XNOR2_X1 U3948 ( .A(n3614), .B(n3613), .ZN(n4499) );
  INV_X1 U3949 ( .A(n4586), .ZN(n4689) );
  OR2_X1 U3951 ( .A1(n4537), .A2(n3889), .ZN(n5325) );
  OR2_X1 U3952 ( .A1(n4857), .A2(n4646), .ZN(n4955) );
  OAI21_X1 U3953 ( .B1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n6547), .A(n4845), 
        .ZN(n4958) );
  AND2_X1 U3954 ( .A1(n5084), .A2(n4767), .ZN(n4842) );
  CLKBUF_X1 U3955 ( .A(n4588), .Z(n6311) );
  NAND3_X1 U3956 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n6567), .A3(n4592), .ZN(
        n4703) );
  INV_X1 U3957 ( .A(n4958), .ZN(n6272) );
  INV_X1 U3958 ( .A(n4345), .ZN(n6565) );
  NAND2_X1 U3959 ( .A1(n4448), .A2(n4442), .ZN(n6569) );
  NOR2_X1 U3960 ( .A1(n4190), .A2(n5685), .ZN(n5669) );
  NOR2_X1 U3961 ( .A1(n4188), .A2(n5866), .ZN(n5852) );
  INV_X1 U3962 ( .A(n5982), .ZN(n5961) );
  INV_X1 U3963 ( .A(n5973), .ZN(n5958) );
  NOR2_X1 U3964 ( .A1(n5103), .A2(n5827), .ZN(n5973) );
  NAND2_X1 U3965 ( .A1(n4478), .A2(n4477), .ZN(n5453) );
  INV_X1 U3966 ( .A(n5445), .ZN(n5466) );
  AND2_X1 U3967 ( .A1(n5380), .A2(n5379), .ZN(n5748) );
  AND2_X1 U3968 ( .A1(n6967), .A2(n5275), .ZN(n5996) );
  AND2_X1 U3969 ( .A1(n6967), .A2(n4538), .ZN(n5997) );
  INV_X1 U3970 ( .A(n5479), .ZN(n6969) );
  INV_X1 U3971 ( .A(n5997), .ZN(n6970) );
  AND2_X1 U3972 ( .A1(n4554), .A2(n4553), .ZN(n6029) );
  OR2_X1 U3973 ( .A1(n4551), .A2(n4731), .ZN(n4552) );
  INV_X2 U3974 ( .A(n6035), .ZN(n6039) );
  INV_X1 U3975 ( .A(n6029), .ZN(n6042) );
  INV_X1 U3976 ( .A(n6045), .ZN(n6079) );
  OR3_X1 U3977 ( .A1(n4551), .A2(n4452), .A3(READY_N), .ZN(n6081) );
  OR2_X1 U3978 ( .A1(n4448), .A2(n3401), .ZN(n6045) );
  OAI21_X1 U3979 ( .B1(n4123), .B2(n3225), .A(n5375), .ZN(n5661) );
  INV_X1 U3980 ( .A(n5748), .ZN(n5495) );
  INV_X1 U3981 ( .A(n5281), .ZN(n5768) );
  AOI21_X1 U3982 ( .B1(n5389), .B2(n5388), .A(n5387), .ZN(n5773) );
  INV_X1 U3983 ( .A(n6134), .ZN(n6157) );
  INV_X1 U3984 ( .A(n5791), .ZN(n6147) );
  NOR2_X1 U3985 ( .A1(n5568), .A2(n4366), .ZN(n5802) );
  NOR2_X1 U3986 ( .A1(n5812), .A2(n4372), .ZN(n5560) );
  OAI21_X1 U3987 ( .B1(n5609), .B2(n5238), .A(n5629), .ZN(n6159) );
  OR2_X1 U3988 ( .A1(n4512), .A2(n6466), .ZN(n6175) );
  OR2_X1 U3989 ( .A1(n4370), .A2(n4336), .ZN(n5815) );
  OR2_X1 U3990 ( .A1(n4370), .A2(n4731), .ZN(n5633) );
  CLKBUF_X1 U3991 ( .A(n4585), .Z(n5642) );
  CLKBUF_X1 U3992 ( .A(n4499), .Z(n5644) );
  INV_X1 U3994 ( .A(n6313), .ZN(n6275) );
  INV_X1 U3995 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6237) );
  OAI21_X1 U3996 ( .B1(n4752), .B2(n6545), .A(n4807), .ZN(n6236) );
  INV_X1 U3997 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n6736) );
  INV_X1 U3998 ( .A(n6548), .ZN(n5327) );
  CLKBUF_X1 U3999 ( .A(n3393), .Z(n3394) );
  INV_X1 U4000 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n6876) );
  NOR2_X1 U4001 ( .A1(n5364), .A2(n6547), .ZN(n6548) );
  OAI21_X1 U4002 ( .B1(n6245), .B2(n6260), .A(n6244), .ZN(n6263) );
  INV_X1 U4003 ( .A(n6266), .ZN(n6241) );
  OR3_X1 U4004 ( .A1(n6321), .A2(n6320), .A3(n6319), .ZN(n6352) );
  NAND2_X1 U4005 ( .A1(n4697), .A2(n6276), .ZN(n5015) );
  OR3_X1 U4006 ( .A1(n4756), .A2(n6276), .A3(n4646), .ZN(n6427) );
  INV_X1 U4007 ( .A(n5062), .ZN(n6419) );
  OR2_X1 U4008 ( .A1(n4892), .A2(n4891), .ZN(n5055) );
  NOR2_X1 U4009 ( .A1(n4703), .A2(n5468), .ZN(n6369) );
  NOR2_X1 U4010 ( .A1(n6069), .A2(n4807), .ZN(n6373) );
  INV_X1 U4011 ( .A(n4851), .ZN(n4934) );
  NOR2_X1 U4012 ( .A1(n6861), .A2(n4807), .ZN(n6383) );
  INV_X1 U4013 ( .A(n6369), .ZN(n5010) );
  INV_X1 U4014 ( .A(n6463), .ZN(n6461) );
  INV_X1 U4015 ( .A(STATE_REG_0__SCAN_IN), .ZN(n6798) );
  NAND2_X1 U4016 ( .A1(n5367), .A2(n5981), .ZN(n4207) );
  OAI22_X1 U4017 ( .A1(n5718), .A2(n5967), .B1(n5717), .B2(n5969), .ZN(n5719)
         );
  NAND2_X1 U4018 ( .A1(n5741), .A2(n4403), .ZN(n4404) );
  NAND2_X1 U4019 ( .A1(n4400), .A2(n6231), .ZN(n4391) );
  OR2_X2 U4020 ( .A1(n5413), .A2(n3343), .ZN(n3220) );
  OAI21_X1 U4021 ( .B1(n4314), .B2(n4345), .A(n4500), .ZN(n3507) );
  BUF_X1 U4022 ( .A(n3508), .Z(n4316) );
  INV_X1 U4023 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3232) );
  INV_X1 U4024 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4734) );
  INV_X1 U4025 ( .A(n4544), .ZN(n3294) );
  NAND2_X1 U4026 ( .A1(n5604), .A2(n4302), .ZN(n3223) );
  AND2_X1 U4027 ( .A1(n4497), .A2(n5349), .ZN(n3224) );
  AND2_X1 U4028 ( .A1(n4122), .A2(n4121), .ZN(n3225) );
  XNOR2_X1 U4029 ( .A(n4180), .B(n4179), .ZN(n5319) );
  OR2_X1 U4030 ( .A1(n5430), .A2(n5394), .ZN(n3226) );
  INV_X1 U4031 ( .A(n5266), .ZN(n5268) );
  AOI21_X1 U4032 ( .B1(n4251), .B2(n3873), .A(n3725), .ZN(n4794) );
  INV_X1 U4033 ( .A(n4794), .ZN(n3726) );
  NOR2_X1 U4034 ( .A1(n5084), .A2(n5644), .ZN(n3227) );
  OR2_X1 U4035 ( .A1(n4408), .A2(n4407), .ZN(n5341) );
  AND4_X1 U4036 ( .A1(n3379), .A2(n3378), .A3(n3377), .A4(n3376), .ZN(n3228)
         );
  INV_X1 U4037 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3436) );
  INV_X1 U4038 ( .A(n6074), .ZN(n6044) );
  NAND2_X1 U4039 ( .A1(n3543), .A2(n3542), .ZN(n3657) );
  INV_X1 U4040 ( .A(n3356), .ZN(n3297) );
  NOR2_X1 U4041 ( .A1(n4423), .A2(n4422), .ZN(n3230) );
  INV_X1 U4042 ( .A(n3617), .ZN(n3619) );
  INV_X1 U4043 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n5155) );
  INV_X1 U4044 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n4463) );
  AND2_X1 U4045 ( .A1(n3744), .A2(n4537), .ZN(n3496) );
  OR2_X1 U4046 ( .A1(n3410), .A2(n3409), .ZN(n3412) );
  INV_X1 U4047 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3231) );
  AND2_X2 U4048 ( .A1(n4734), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3238)
         );
  OR2_X1 U4049 ( .A1(n3579), .A2(n3578), .ZN(n4274) );
  NOR2_X1 U4050 ( .A1(n3556), .A2(n3555), .ZN(n4235) );
  NAND2_X1 U4051 ( .A1(n3205), .A2(n5081), .ZN(n3512) );
  INV_X1 U4052 ( .A(n3744), .ZN(n3752) );
  INV_X1 U4053 ( .A(n4212), .ZN(n3616) );
  AOI22_X1 U4054 ( .A1(n3443), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3572), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3466) );
  AOI22_X1 U4055 ( .A1(n3443), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3572), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3458) );
  AND2_X2 U4056 ( .A1(n4750), .A2(n4738), .ZN(n3544) );
  OR2_X1 U4057 ( .A1(n5394), .A2(n5395), .ZN(n4022) );
  OR2_X1 U4058 ( .A1(n3607), .A2(n3606), .ZN(n4212) );
  INV_X1 U4059 ( .A(n4274), .ZN(n4284) );
  OR2_X1 U4060 ( .A1(n3721), .A2(n3720), .ZN(n4260) );
  NAND2_X1 U4061 ( .A1(n3513), .A2(n3512), .ZN(n4353) );
  AOI21_X1 U4062 ( .B1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n6441), .A(n3428), 
        .ZN(n3437) );
  BUF_X1 U4063 ( .A(n3533), .Z(n3659) );
  NAND2_X1 U4064 ( .A1(n5982), .A2(EBX_REG_29__SCAN_IN), .ZN(n4421) );
  NOR2_X1 U4065 ( .A1(n4085), .A2(n4024), .ZN(n4025) );
  OR2_X1 U4066 ( .A1(n3516), .A2(n4463), .ZN(n4171) );
  OR2_X1 U4067 ( .A1(n3615), .A2(n4284), .ZN(n4281) );
  NAND2_X1 U4068 ( .A1(n4497), .A2(n3494), .ZN(n3365) );
  AOI221_X1 U4069 ( .B1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n3437), .C1(
        n3436), .C2(n3437), .A(n3435), .ZN(n3478) );
  AND2_X1 U4070 ( .A1(n4124), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4125)
         );
  INV_X1 U4071 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3828) );
  NAND2_X1 U4072 ( .A1(n4702), .A2(n4593), .ZN(n3524) );
  NAND2_X1 U4073 ( .A1(n3286), .A2(n3196), .ZN(n3352) );
  AND2_X1 U4074 ( .A1(n3328), .A2(n3327), .ZN(n5290) );
  NAND2_X1 U4075 ( .A1(n3282), .A2(n3281), .ZN(n3285) );
  OR2_X1 U4076 ( .A1(n3974), .A2(n5418), .ZN(n5394) );
  AND2_X1 U4077 ( .A1(n5275), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3685) );
  AND4_X1 U4078 ( .A1(n3260), .A2(n3259), .A3(n3258), .A4(n3257), .ZN(n3261)
         );
  AND2_X1 U4079 ( .A1(n4025), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4124)
         );
  AND2_X1 U4080 ( .A1(n3975), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n3976)
         );
  INV_X1 U4081 ( .A(n3846), .ZN(n3833) );
  NOR2_X1 U4082 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n6564), .ZN(n4177) );
  XNOR2_X1 U4083 ( .A(n3728), .B(n3731), .ZN(n4243) );
  AND2_X1 U4084 ( .A1(n5604), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n4428)
         );
  NOR2_X1 U4085 ( .A1(n4281), .A2(n4280), .ZN(n4282) );
  AND2_X1 U4086 ( .A1(n3203), .A2(n3401), .ZN(n4269) );
  NOR2_X1 U4087 ( .A1(n4688), .A2(n5642), .ZN(n6277) );
  XNOR2_X1 U4088 ( .A(n3625), .B(n3628), .ZN(n4585) );
  NAND2_X1 U4089 ( .A1(n3380), .A2(n3228), .ZN(n3482) );
  OR2_X1 U4090 ( .A1(n5655), .A2(n6829), .ZN(n4203) );
  AND2_X1 U4091 ( .A1(n3350), .A2(n3349), .ZN(n5396) );
  INV_X1 U4092 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5870) );
  INV_X1 U4093 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n5935) );
  OR2_X1 U4094 ( .A1(n4181), .A2(n6707), .ZN(n4183) );
  NAND2_X1 U4095 ( .A1(n4325), .A2(n4187), .ZN(n5976) );
  AND2_X1 U4096 ( .A1(n3325), .A2(n3324), .ZN(n5447) );
  AND2_X1 U4097 ( .A1(n3942), .A2(n3941), .ZN(n5412) );
  INV_X1 U4098 ( .A(n4177), .ZN(n4096) );
  NAND2_X1 U4099 ( .A1(n5266), .A2(n4104), .ZN(n5380) );
  XNOR2_X1 U4100 ( .A(n3845), .B(n3833), .ZN(n5458) );
  NAND2_X1 U4101 ( .A1(n3777), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3801)
         );
  INV_X1 U4102 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n6897) );
  NAND2_X1 U4103 ( .A1(n5390), .A2(n4436), .ZN(n5382) );
  AND2_X1 U4104 ( .A1(n3305), .A2(n3304), .ZN(n5128) );
  AND2_X1 U4105 ( .A1(n5633), .A2(n5630), .ZN(n5609) );
  OR2_X1 U4106 ( .A1(n4551), .A2(n4328), .ZN(n4329) );
  INV_X1 U4108 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6436) );
  INV_X1 U4109 ( .A(n5642), .ZN(n4765) );
  AND2_X1 U4110 ( .A1(n6736), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3662) );
  NAND2_X1 U4111 ( .A1(n3475), .A2(n4555), .ZN(n5363) );
  NAND2_X1 U4112 ( .A1(n4204), .A2(n4203), .ZN(n4205) );
  NOR2_X1 U4113 ( .A1(n4189), .A2(n5736), .ZN(n5706) );
  AND2_X1 U4114 ( .A1(n4196), .A2(n5986), .ZN(n5906) );
  XNOR2_X1 U4115 ( .A(n4183), .B(n4182), .ZN(n5320) );
  AND2_X1 U4116 ( .A1(n5200), .A2(n5199), .ZN(n5202) );
  AND2_X1 U4118 ( .A1(n3958), .A2(n3957), .ZN(n5403) );
  AND2_X1 U4119 ( .A1(n6967), .A2(n4539), .ZN(n5479) );
  INV_X1 U4120 ( .A(n6044), .ZN(n6051) );
  INV_X1 U4121 ( .A(n6081), .ZN(n6075) );
  OR2_X1 U4122 ( .A1(n4323), .A2(n3196), .ZN(n4452) );
  NAND2_X1 U4123 ( .A1(n4123), .A2(n3225), .ZN(n5375) );
  NAND2_X1 U4124 ( .A1(n3960), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3959)
         );
  NAND2_X1 U4125 ( .A1(n5429), .A2(n5431), .ZN(n5430) );
  NAND2_X1 U4126 ( .A1(n3756), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3776)
         );
  NAND2_X1 U4127 ( .A1(PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n3681), .ZN(n3705)
         );
  AND2_X1 U4128 ( .A1(n4226), .A2(n4227), .ZN(n4548) );
  OR2_X1 U4129 ( .A1(n6224), .A2(n6223), .ZN(n4632) );
  CLKBUF_X1 U4130 ( .A(n4628), .Z(n4629) );
  INV_X1 U4131 ( .A(n4382), .ZN(n6212) );
  INV_X1 U4132 ( .A(n6177), .ZN(n6227) );
  OAI21_X1 U4133 ( .B1(n4987), .B2(n4985), .A(n4984), .ZN(n5063) );
  OR2_X1 U4134 ( .A1(n4857), .A2(n4856), .ZN(n4867) );
  OAI21_X1 U4135 ( .B1(n4961), .B2(n4960), .A(n4959), .ZN(n5051) );
  OAI21_X1 U4136 ( .B1(n4650), .B2(n4649), .A(n4648), .ZN(n5071) );
  INV_X1 U4137 ( .A(n6314), .ZN(n6350) );
  INV_X1 U4138 ( .A(n5015), .ZN(n6370) );
  INV_X1 U4139 ( .A(n5148), .ZN(n6389) );
  INV_X1 U4140 ( .A(n4866), .ZN(n6276) );
  NOR2_X1 U4141 ( .A1(n6063), .A2(n4807), .ZN(n6360) );
  AND2_X1 U4142 ( .A1(n3662), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6463) );
  NOR2_X1 U4143 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6573), .ZN(n6534) );
  OR2_X1 U4144 ( .A1(n4551), .A2(n5363), .ZN(n4448) );
  AOI21_X1 U4145 ( .B1(n5319), .B2(n5952), .A(n4205), .ZN(n4206) );
  OAI21_X1 U4146 ( .B1(n4424), .B2(REIP_REG_29__SCAN_IN), .A(n3230), .ZN(n4425) );
  AOI211_X1 U4147 ( .C1(EBX_REG_21__SCAN_IN), .C2(n5982), .A(n5720), .B(n5719), 
        .ZN(n5722) );
  INV_X1 U4148 ( .A(n5894), .ZN(n5865) );
  OR2_X1 U4149 ( .A1(n5320), .A2(n4413), .ZN(n5967) );
  OAI21_X1 U4150 ( .B1(n5266), .B2(n5269), .A(n5388), .ZN(n5692) );
  OAI21_X1 U4151 ( .B1(n5403), .B2(n5402), .A(n3226), .ZN(n5711) );
  OAI211_X2 U4152 ( .C1(n4551), .C2(n4723), .A(n4536), .B(n6081), .ZN(n6967)
         );
  OR2_X1 U4153 ( .A1(n6029), .A2(n6040), .ZN(n6035) );
  NAND2_X1 U4154 ( .A1(n5831), .A2(n4393), .ZN(n5791) );
  NAND2_X1 U4155 ( .A1(n4402), .A2(n6313), .ZN(n6138) );
  OR2_X1 U4156 ( .A1(n5312), .A2(n5313), .ZN(n4389) );
  AND2_X1 U4157 ( .A1(n5549), .A2(n4385), .ZN(n5808) );
  OR2_X1 U4158 ( .A1(n4370), .A2(n4349), .ZN(n6177) );
  AND2_X1 U4159 ( .A1(n4486), .A2(n4488), .ZN(n6235) );
  INV_X1 U4160 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6430) );
  OR2_X1 U4161 ( .A1(n4867), .A2(n6276), .ZN(n5070) );
  OR2_X1 U4162 ( .A1(n4955), .A2(n6276), .ZN(n6266) );
  OR2_X1 U4163 ( .A1(n4955), .A2(n4866), .ZN(n5078) );
  AOI21_X1 U4164 ( .B1(n6275), .B2(n6281), .A(n6274), .ZN(n6306) );
  NAND2_X1 U4165 ( .A1(n4697), .A2(n4866), .ZN(n6377) );
  NOR2_X1 U4166 ( .A1(n4809), .A2(n4808), .ZN(n5008) );
  OR2_X1 U4167 ( .A1(n4775), .A2(n4866), .ZN(n5148) );
  AOI21_X1 U4168 ( .B1(n5153), .B2(n5150), .A(n5147), .ZN(n5190) );
  INV_X1 U4169 ( .A(n6360), .ZN(n5179) );
  NAND2_X1 U4170 ( .A1(n4668), .A2(n6276), .ZN(n4851) );
  INV_X1 U4171 ( .A(n4914), .ZN(n4938) );
  INV_X1 U4172 ( .A(n4800), .ZN(n4709) );
  INV_X1 U4173 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6547) );
  INV_X1 U4174 ( .A(n6544), .ZN(n6540) );
  INV_X1 U4175 ( .A(n6534), .ZN(n6533) );
  NAND2_X1 U4176 ( .A1(n4207), .A2(n4206), .ZN(U2796) );
  NOR2_X4 U4177 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4750) );
  AOI22_X1 U4178 ( .A1(n4049), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3852), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3236) );
  AND2_X4 U4179 ( .A1(n3232), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4504)
         );
  AND2_X2 U4180 ( .A1(n4738), .A2(n5332), .ZN(n3545) );
  AOI22_X1 U4181 ( .A1(n3584), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3545), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3235) );
  AOI22_X1 U4182 ( .A1(n3667), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3566), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3234) );
  AND2_X2 U4184 ( .A1(n4505), .A2(n4738), .ZN(n3467) );
  AOI22_X1 U4185 ( .A1(n4050), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3467), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3233) );
  NAND4_X1 U4186 ( .A1(n3236), .A2(n3235), .A3(n3234), .A4(n3233), .ZN(n3244)
         );
  AND2_X4 U4187 ( .A1(n3237), .A2(n4504), .ZN(n3571) );
  AND2_X2 U4188 ( .A1(n3238), .A2(n4750), .ZN(n3550) );
  AOI22_X1 U4189 ( .A1(n3571), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3550), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3242) );
  AOI22_X1 U4190 ( .A1(n3666), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3597), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3241) );
  AND2_X2 U4191 ( .A1(n4750), .A2(n4722), .ZN(n3443) );
  AOI22_X1 U4192 ( .A1(n3443), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3572), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3240) );
  AND2_X4 U4193 ( .A1(n4504), .A2(n3238), .ZN(n3573) );
  AOI22_X1 U4194 ( .A1(n3573), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3544), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3239) );
  NAND4_X1 U4195 ( .A1(n3242), .A2(n3241), .A3(n3240), .A4(n3239), .ZN(n3243)
         );
  NAND2_X1 U4196 ( .A1(n3852), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3248) );
  NAND2_X1 U4197 ( .A1(n3571), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3247)
         );
  NAND2_X1 U4198 ( .A1(n3550), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3246) );
  NAND2_X1 U4199 ( .A1(n4049), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3245)
         );
  NAND2_X1 U4200 ( .A1(n3198), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3252)
         );
  NAND2_X1 U4201 ( .A1(n3597), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3251)
         );
  NAND2_X1 U4202 ( .A1(n3666), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3250) );
  NAND2_X1 U4203 ( .A1(n3667), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3249) );
  AND4_X2 U4204 ( .A1(n3252), .A2(n3251), .A3(n3250), .A4(n3249), .ZN(n3263)
         );
  NAND2_X1 U4205 ( .A1(n4050), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3256) );
  NAND2_X1 U4206 ( .A1(n3467), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3255) );
  NAND2_X1 U4207 ( .A1(n3443), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3254)
         );
  NAND2_X1 U4208 ( .A1(n3572), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3253)
         );
  NAND2_X1 U4209 ( .A1(n3573), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3260) );
  NAND2_X1 U4210 ( .A1(n3584), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3259) );
  NAND2_X1 U4211 ( .A1(n3544), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3258) );
  NAND2_X1 U4212 ( .A1(n3545), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3257) );
  NAND4_X4 U4213 ( .A1(n3264), .A2(n3263), .A3(n3262), .A4(n3261), .ZN(n3493)
         );
  NAND2_X2 U4214 ( .A1(n4605), .A2(n4555), .ZN(n3361) );
  AOI22_X1 U4215 ( .A1(n3597), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3566), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3267) );
  AOI22_X1 U4216 ( .A1(n4049), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3852), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3266) );
  AOI22_X1 U4217 ( .A1(n3467), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3572), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3272) );
  AOI22_X1 U4218 ( .A1(n3571), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3550), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3271) );
  AOI22_X1 U4219 ( .A1(n3544), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n3545), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3270) );
  AOI22_X1 U4220 ( .A1(n3666), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3667), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3269) );
  NAND2_X1 U4221 ( .A1(n3401), .A2(n4555), .ZN(n3287) );
  AOI22_X1 U4222 ( .A1(n4470), .A2(EBX_REG_30__SCAN_IN), .B1(
        INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n3196), .ZN(n4341) );
  NOR2_X2 U4223 ( .A1(n3219), .A2(n3287), .ZN(n3356) );
  INV_X1 U4224 ( .A(EBX_REG_1__SCAN_IN), .ZN(n3275) );
  NAND2_X1 U4225 ( .A1(n3356), .A2(n3275), .ZN(n3278) );
  INV_X1 U4226 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n6234) );
  NAND2_X1 U4227 ( .A1(n3361), .A2(n6234), .ZN(n3276) );
  OAI211_X1 U4228 ( .C1(n3287), .C2(EBX_REG_1__SCAN_IN), .A(n3276), .B(n3494), 
        .ZN(n3277) );
  NAND2_X1 U4229 ( .A1(n3278), .A2(n3277), .ZN(n3283) );
  NAND2_X1 U4230 ( .A1(n3361), .A2(EBX_REG_0__SCAN_IN), .ZN(n3280) );
  INV_X1 U4231 ( .A(EBX_REG_0__SCAN_IN), .ZN(n5109) );
  NAND2_X1 U4232 ( .A1(n3494), .A2(n5109), .ZN(n3279) );
  AND2_X1 U4233 ( .A1(n3280), .A2(n3279), .ZN(n4472) );
  NAND2_X1 U4234 ( .A1(n3283), .A2(n4472), .ZN(n3284) );
  AND2_X2 U4235 ( .A1(n3285), .A2(n3284), .ZN(n5093) );
  INV_X1 U4236 ( .A(n3287), .ZN(n4497) );
  NAND2_X1 U4237 ( .A1(n4496), .A2(n3285), .ZN(n4544) );
  MUX2_X1 U4238 ( .A(n3297), .B(n3361), .S(EBX_REG_2__SCAN_IN), .Z(n3290) );
  INV_X1 U4239 ( .A(n3361), .ZN(n3286) );
  NAND3_X1 U4240 ( .A1(n3219), .A2(n3196), .A3(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .ZN(n3288) );
  AND2_X1 U4241 ( .A1(n3352), .A2(n3288), .ZN(n3289) );
  NAND2_X1 U4242 ( .A1(n3290), .A2(n3289), .ZN(n4575) );
  OR2_X1 U4243 ( .A1(n4470), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3292)
         );
  MUX2_X1 U4244 ( .A(n3365), .B(n3219), .S(EBX_REG_3__SCAN_IN), .Z(n3291) );
  AND2_X1 U4245 ( .A1(n3292), .A2(n3291), .ZN(n4574) );
  OR2_X1 U4246 ( .A1(n4470), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3296)
         );
  MUX2_X1 U4247 ( .A(n3365), .B(n3494), .S(EBX_REG_5__SCAN_IN), .Z(n3295) );
  AND2_X1 U4248 ( .A1(n3296), .A2(n3295), .ZN(n4637) );
  OR2_X1 U4249 ( .A1(n3297), .A2(EBX_REG_4__SCAN_IN), .ZN(n3300) );
  INV_X1 U4250 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6202) );
  NAND2_X1 U4251 ( .A1(n3361), .A2(n6202), .ZN(n3298) );
  OAI211_X1 U4252 ( .C1(n3196), .C2(EBX_REG_4__SCAN_IN), .A(n3298), .B(n3219), 
        .ZN(n3299) );
  NAND2_X1 U4253 ( .A1(n3300), .A2(n3299), .ZN(n4638) );
  NAND2_X1 U4254 ( .A1(n4637), .A2(n4638), .ZN(n3301) );
  MUX2_X1 U4255 ( .A(n3365), .B(n3494), .S(EBX_REG_7__SCAN_IN), .Z(n3302) );
  OAI21_X1 U4256 ( .B1(INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n4470), .A(n3302), 
        .ZN(n5133) );
  OR2_X1 U4257 ( .A1(n3297), .A2(EBX_REG_6__SCAN_IN), .ZN(n3305) );
  INV_X1 U4258 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n6752) );
  NAND2_X1 U4259 ( .A1(n3361), .A2(n6752), .ZN(n3303) );
  OAI211_X1 U4260 ( .C1(n3196), .C2(EBX_REG_6__SCAN_IN), .A(n3303), .B(n3219), 
        .ZN(n3304) );
  NOR2_X1 U4261 ( .A1(n5133), .A2(n5128), .ZN(n3306) );
  NAND2_X1 U4262 ( .A1(n4640), .A2(n3306), .ZN(n5131) );
  INV_X1 U4263 ( .A(EBX_REG_8__SCAN_IN), .ZN(n5944) );
  NAND2_X1 U4264 ( .A1(n3356), .A2(n5944), .ZN(n3309) );
  INV_X1 U4265 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n6816) );
  NAND2_X1 U4266 ( .A1(n3361), .A2(n6816), .ZN(n3307) );
  OAI211_X1 U4267 ( .C1(n3196), .C2(EBX_REG_8__SCAN_IN), .A(n3307), .B(n3494), 
        .ZN(n3308) );
  OR2_X2 U4268 ( .A1(n5131), .A2(n5136), .ZN(n5137) );
  MUX2_X1 U4269 ( .A(n3365), .B(n3219), .S(EBX_REG_9__SCAN_IN), .Z(n3310) );
  OAI21_X1 U4270 ( .B1(INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n4470), .A(n3310), 
        .ZN(n5126) );
  MUX2_X1 U4271 ( .A(n3297), .B(n3361), .S(EBX_REG_10__SCAN_IN), .Z(n3313) );
  NAND2_X1 U4272 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n3196), .ZN(n3311) );
  AND2_X1 U4273 ( .A1(n3352), .A2(n3311), .ZN(n3312) );
  NAND2_X1 U4274 ( .A1(n3313), .A2(n3312), .ZN(n5199) );
  OR2_X1 U4275 ( .A1(n3365), .A2(EBX_REG_11__SCAN_IN), .ZN(n3316) );
  NAND2_X1 U4276 ( .A1(n3494), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n3314) );
  OAI211_X1 U4277 ( .C1(n3196), .C2(EBX_REG_11__SCAN_IN), .A(n3361), .B(n3314), 
        .ZN(n3315) );
  NAND2_X1 U4278 ( .A1(n5202), .A2(n5196), .ZN(n5195) );
  MUX2_X1 U4279 ( .A(n3297), .B(n3361), .S(EBX_REG_12__SCAN_IN), .Z(n3319) );
  NAND2_X1 U4280 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n3196), .ZN(n3317) );
  AND2_X1 U4281 ( .A1(n3352), .A2(n3317), .ZN(n3318) );
  OR2_X2 U4282 ( .A1(n5195), .A2(n5225), .ZN(n5456) );
  OR2_X1 U4283 ( .A1(n3365), .A2(EBX_REG_13__SCAN_IN), .ZN(n3322) );
  NAND2_X1 U4284 ( .A1(n3219), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n3320) );
  OAI211_X1 U4285 ( .C1(n3196), .C2(EBX_REG_13__SCAN_IN), .A(n3361), .B(n3320), 
        .ZN(n3321) );
  NAND2_X1 U4286 ( .A1(n3322), .A2(n3321), .ZN(n5457) );
  OR2_X2 U4287 ( .A1(n5456), .A2(n5457), .ZN(n5454) );
  MUX2_X1 U4288 ( .A(n3297), .B(n3361), .S(EBX_REG_14__SCAN_IN), .Z(n3325) );
  NAND2_X1 U4289 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n3196), .ZN(n3323) );
  AND2_X1 U4290 ( .A1(n3352), .A2(n3323), .ZN(n3324) );
  NOR2_X2 U4291 ( .A1(n5454), .A2(n5447), .ZN(n5291) );
  OR2_X1 U4292 ( .A1(n3365), .A2(EBX_REG_15__SCAN_IN), .ZN(n3328) );
  NAND2_X1 U4293 ( .A1(n3219), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n3326) );
  OAI211_X1 U4294 ( .C1(n3196), .C2(EBX_REG_15__SCAN_IN), .A(n3361), .B(n3326), 
        .ZN(n3327) );
  NAND2_X1 U4295 ( .A1(n5291), .A2(n5290), .ZN(n5292) );
  MUX2_X1 U4296 ( .A(n3297), .B(n3361), .S(EBX_REG_16__SCAN_IN), .Z(n3331) );
  NAND2_X1 U4297 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n3196), .ZN(n3329) );
  AND2_X1 U4298 ( .A1(n3352), .A2(n3329), .ZN(n3330) );
  OR2_X1 U4299 ( .A1(n3365), .A2(EBX_REG_17__SCAN_IN), .ZN(n3334) );
  NAND2_X1 U4300 ( .A1(n3494), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n3332) );
  OAI211_X1 U4301 ( .C1(n3196), .C2(EBX_REG_17__SCAN_IN), .A(n3361), .B(n3332), 
        .ZN(n3333) );
  NAND2_X1 U4302 ( .A1(n3334), .A2(n3333), .ZN(n5437) );
  MUX2_X1 U4303 ( .A(n3297), .B(n3361), .S(EBX_REG_19__SCAN_IN), .Z(n3337) );
  NAND2_X1 U4304 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n3196), .ZN(n3335) );
  AND2_X1 U4305 ( .A1(n3352), .A2(n3335), .ZN(n3336) );
  NAND2_X1 U4306 ( .A1(n3337), .A2(n3336), .ZN(n5423) );
  NAND2_X1 U4307 ( .A1(n5436), .A2(n5423), .ZN(n5413) );
  OR2_X1 U4308 ( .A1(n4470), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n3339)
         );
  INV_X1 U4309 ( .A(EBX_REG_20__SCAN_IN), .ZN(n5416) );
  NAND2_X1 U4310 ( .A1(n4497), .A2(n5416), .ZN(n3338) );
  AND2_X1 U4311 ( .A1(n3339), .A2(n3338), .ZN(n5414) );
  OR2_X1 U4312 ( .A1(n4470), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n3340)
         );
  OR2_X1 U4313 ( .A1(n3196), .A2(EBX_REG_18__SCAN_IN), .ZN(n5420) );
  NAND2_X1 U4314 ( .A1(n3340), .A2(n5420), .ZN(n5421) );
  NAND2_X1 U4315 ( .A1(n5419), .A2(EBX_REG_20__SCAN_IN), .ZN(n3342) );
  NAND2_X1 U4316 ( .A1(n5421), .A2(n3219), .ZN(n3341) );
  OAI211_X1 U4317 ( .C1(n5414), .C2(n5421), .A(n3342), .B(n3341), .ZN(n3343)
         );
  MUX2_X1 U4318 ( .A(n3365), .B(n3494), .S(EBX_REG_21__SCAN_IN), .Z(n3344) );
  OAI21_X1 U4319 ( .B1(INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n4470), .A(n3344), 
        .ZN(n5410) );
  NOR2_X2 U4320 ( .A1(n3220), .A2(n5410), .ZN(n5404) );
  MUX2_X1 U4321 ( .A(n3297), .B(n3361), .S(EBX_REG_22__SCAN_IN), .Z(n3347) );
  NAND2_X1 U4322 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n3196), .ZN(n3345) );
  AND2_X1 U4323 ( .A1(n3352), .A2(n3345), .ZN(n3346) );
  NAND2_X1 U4324 ( .A1(n3347), .A2(n3346), .ZN(n5405) );
  AND2_X2 U4325 ( .A1(n5404), .A2(n5405), .ZN(n5397) );
  OR2_X1 U4326 ( .A1(n3365), .A2(EBX_REG_23__SCAN_IN), .ZN(n3350) );
  NAND2_X1 U4327 ( .A1(n3494), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n3348) );
  OAI211_X1 U4328 ( .C1(n3196), .C2(EBX_REG_23__SCAN_IN), .A(n3361), .B(n3348), 
        .ZN(n3349) );
  NAND2_X1 U4329 ( .A1(n5397), .A2(n5396), .ZN(n5255) );
  MUX2_X1 U4330 ( .A(n3297), .B(n3361), .S(EBX_REG_24__SCAN_IN), .Z(n3354) );
  NAND2_X1 U4331 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n3196), .ZN(n3351) );
  AND2_X1 U4332 ( .A1(n3352), .A2(n3351), .ZN(n3353) );
  MUX2_X1 U4333 ( .A(n3365), .B(n3219), .S(EBX_REG_25__SCAN_IN), .Z(n3355) );
  OAI21_X1 U4334 ( .B1(INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n4470), .A(n3355), 
        .ZN(n5391) );
  INV_X1 U4335 ( .A(EBX_REG_26__SCAN_IN), .ZN(n5679) );
  NAND2_X1 U4336 ( .A1(n3356), .A2(n5679), .ZN(n3359) );
  INV_X1 U4337 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n4435) );
  NAND2_X1 U4338 ( .A1(n3361), .A2(n4435), .ZN(n3357) );
  OAI211_X1 U4339 ( .C1(n3196), .C2(EBX_REG_26__SCAN_IN), .A(n3357), .B(n3219), 
        .ZN(n3358) );
  NAND2_X1 U4340 ( .A1(n3359), .A2(n3358), .ZN(n4436) );
  MUX2_X1 U4341 ( .A(n3365), .B(n3494), .S(EBX_REG_27__SCAN_IN), .Z(n3360) );
  OAI21_X1 U4342 ( .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n4470), .A(n3360), 
        .ZN(n5381) );
  MUX2_X1 U4343 ( .A(n3297), .B(n3361), .S(EBX_REG_28__SCAN_IN), .Z(n3363) );
  NAND2_X1 U4344 ( .A1(INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n3196), .ZN(n3362) );
  AND2_X1 U4345 ( .A1(n3363), .A2(n3362), .ZN(n5372) );
  NAND2_X2 U4346 ( .A1(n5371), .A2(n3364), .ZN(n5374) );
  INV_X1 U4347 ( .A(n5374), .ZN(n4340) );
  NOR2_X1 U4348 ( .A1(n4470), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n3368)
         );
  MUX2_X1 U4349 ( .A(EBX_REG_29__SCAN_IN), .B(n3368), .S(n3219), .Z(n3367) );
  NOR2_X1 U4350 ( .A1(n3365), .A2(EBX_REG_29__SCAN_IN), .ZN(n3366) );
  NOR2_X1 U4351 ( .A1(n3367), .A2(n3366), .ZN(n4409) );
  NAND2_X1 U4352 ( .A1(n4340), .A2(n4409), .ZN(n4412) );
  INV_X1 U4353 ( .A(n4412), .ZN(n3369) );
  INV_X1 U4354 ( .A(EBX_REG_29__SCAN_IN), .ZN(n5349) );
  NOR3_X4 U4355 ( .A1(n5374), .A2(n3368), .A3(n3224), .ZN(n4337) );
  NOR2_X1 U4356 ( .A1(n4337), .A2(n5419), .ZN(n4338) );
  AOI21_X1 U4357 ( .B1(n4341), .B2(n3369), .A(n4338), .ZN(n3371) );
  OAI22_X1 U4358 ( .A1(n4470), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        EBX_REG_31__SCAN_IN), .B2(n3196), .ZN(n3370) );
  XNOR2_X1 U4359 ( .A(n3371), .B(n3370), .ZN(n5367) );
  NAND2_X1 U4360 ( .A1(n4324), .A2(n6564), .ZN(n4416) );
  INV_X1 U4361 ( .A(EBX_REG_31__SCAN_IN), .ZN(n4415) );
  AOI22_X1 U4362 ( .A1(n3571), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3852), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3375) );
  AOI22_X1 U4363 ( .A1(n4049), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3550), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3374) );
  AOI22_X1 U4364 ( .A1(n4050), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3443), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3373) );
  AOI22_X1 U4365 ( .A1(n3467), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3572), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3372) );
  AOI22_X1 U4366 ( .A1(n3597), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3566), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3379) );
  AOI22_X1 U4367 ( .A1(n3666), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3667), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3378) );
  AOI22_X1 U4368 ( .A1(n3573), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3584), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3377) );
  AOI22_X1 U4369 ( .A1(n3544), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n3545), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3376) );
  AND3_X4 U4370 ( .A1(n4346), .A2(STATE2_REG_0__SCAN_IN), .A3(n3493), .ZN(
        n3744) );
  AOI22_X1 U4371 ( .A1(n3467), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3443), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3384) );
  AOI22_X1 U4372 ( .A1(n3597), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3852), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3383) );
  AOI22_X1 U4373 ( .A1(n3584), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3545), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3382) );
  AOI22_X1 U4374 ( .A1(n3666), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3667), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3381) );
  AND2_X1 U4375 ( .A1(n3217), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3385) );
  NOR2_X1 U4376 ( .A1(n3386), .A2(n3385), .ZN(n3390) );
  AOI22_X1 U4377 ( .A1(n3550), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3566), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3389) );
  AOI22_X1 U4378 ( .A1(n4050), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3572), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3388) );
  AOI22_X1 U4379 ( .A1(n3573), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3544), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3387) );
  NAND2_X1 U4380 ( .A1(n6436), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3411) );
  NAND2_X1 U4381 ( .A1(n3394), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3395) );
  NAND2_X1 U4382 ( .A1(n3411), .A2(n3395), .ZN(n3410) );
  NAND2_X1 U4383 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n6430), .ZN(n3409) );
  INV_X1 U4384 ( .A(n3409), .ZN(n3396) );
  XNOR2_X1 U4385 ( .A(n3410), .B(n3396), .ZN(n3476) );
  INV_X1 U4386 ( .A(n4346), .ZN(n3592) );
  INV_X4 U4387 ( .A(n3493), .ZN(n4593) );
  NAND2_X1 U4388 ( .A1(n3750), .A2(n3401), .ZN(n3397) );
  NAND2_X1 U4389 ( .A1(n3397), .A2(n3203), .ZN(n3406) );
  OAI21_X1 U4390 ( .B1(n6430), .B2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(n3409), 
        .ZN(n3398) );
  INV_X1 U4391 ( .A(n3398), .ZN(n3400) );
  NAND2_X1 U4392 ( .A1(n3750), .A2(n3400), .ZN(n3399) );
  NAND2_X1 U4393 ( .A1(n3399), .A2(n3431), .ZN(n3405) );
  AOI21_X1 U4394 ( .B1(n4331), .B2(n3400), .A(n4593), .ZN(n3403) );
  INV_X4 U4395 ( .A(n3401), .ZN(n4702) );
  NAND2_X1 U4396 ( .A1(n4702), .A2(n3203), .ZN(n3402) );
  NAND2_X1 U4397 ( .A1(n3524), .A2(n3402), .ZN(n3414) );
  OR2_X1 U4398 ( .A1(n3403), .A2(n3414), .ZN(n3404) );
  OAI211_X1 U4399 ( .C1(n3406), .C2(n3476), .A(n3405), .B(n3404), .ZN(n3408)
         );
  NAND3_X1 U4400 ( .A1(n3406), .A2(STATE2_REG_0__SCAN_IN), .A3(n3476), .ZN(
        n3407) );
  OAI211_X1 U4401 ( .C1(n3431), .C2(n3476), .A(n3408), .B(n3407), .ZN(n3419)
         );
  NAND2_X1 U4402 ( .A1(n3412), .A2(n3411), .ZN(n3422) );
  NAND2_X1 U4403 ( .A1(n4859), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3423) );
  NAND2_X1 U4404 ( .A1(n6876), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3413) );
  NAND2_X1 U4405 ( .A1(n3423), .A2(n3413), .ZN(n3420) );
  XNOR2_X1 U4406 ( .A(n3422), .B(n3420), .ZN(n3477) );
  NAND2_X1 U4407 ( .A1(n3750), .A2(n3477), .ZN(n3416) );
  INV_X1 U4408 ( .A(n3414), .ZN(n3415) );
  OAI211_X1 U4409 ( .C1(n3477), .C2(n3752), .A(n3416), .B(n3415), .ZN(n3418)
         );
  NOR2_X1 U4410 ( .A1(n3416), .A2(n3415), .ZN(n3417) );
  AOI21_X1 U4411 ( .B1(n3419), .B2(n3418), .A(n3417), .ZN(n3434) );
  INV_X1 U4412 ( .A(n3420), .ZN(n3421) );
  NAND2_X1 U4413 ( .A1(n3422), .A2(n3421), .ZN(n3424) );
  NAND2_X1 U4414 ( .A1(n3424), .A2(n3423), .ZN(n3426) );
  XNOR2_X1 U4415 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3425) );
  NAND3_X1 U4416 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n3437), .A3(n3436), .ZN(n3430) );
  NOR2_X1 U4417 ( .A1(n3426), .A2(n3425), .ZN(n3427) );
  NOR2_X1 U4418 ( .A1(n3428), .A2(n3427), .ZN(n3429) );
  NAND2_X1 U4419 ( .A1(n3430), .A2(n3429), .ZN(n3481) );
  AOI22_X1 U4420 ( .A1(n3481), .A2(n3438), .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n6567), .ZN(n3432) );
  OAI21_X1 U4421 ( .B1(n3434), .B2(n3433), .A(n3432), .ZN(n3440) );
  NOR2_X1 U4422 ( .A1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n6237), .ZN(n3435)
         );
  NAND2_X1 U4423 ( .A1(n3478), .A2(n3438), .ZN(n3439) );
  NAND2_X1 U4424 ( .A1(n3440), .A2(n3439), .ZN(n3442) );
  AOI22_X1 U4425 ( .A1(n3667), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3566), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3446) );
  AOI22_X1 U4426 ( .A1(n3467), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3443), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3445) );
  AOI22_X1 U4427 ( .A1(n3544), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3545), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3444) );
  AOI22_X1 U4428 ( .A1(INSTQUEUE_REG_10__6__SCAN_IN), .A2(n3571), .B1(n3550), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3451) );
  AOI22_X1 U4429 ( .A1(n3666), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3597), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3450) );
  AOI22_X1 U4430 ( .A1(n3573), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3584), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3449) );
  AOI22_X1 U4431 ( .A1(n4050), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3572), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3448) );
  NAND2_X2 U4432 ( .A1(n3453), .A2(n3452), .ZN(n3622) );
  NAND2_X1 U4433 ( .A1(n4678), .A2(n3622), .ZN(n3462) );
  AOI22_X1 U4434 ( .A1(n4050), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3467), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3457) );
  AOI22_X1 U4435 ( .A1(n3566), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3852), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3456) );
  AOI22_X1 U4436 ( .A1(n3666), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3584), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3455) );
  AOI22_X1 U4437 ( .A1(n3544), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3545), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3454) );
  AOI22_X1 U4438 ( .A1(n3571), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4049), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3461) );
  AOI22_X1 U4439 ( .A1(n3597), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3550), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3460) );
  AOI22_X1 U4440 ( .A1(n3573), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3667), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3459) );
  NAND2_X1 U4441 ( .A1(n3462), .A2(n3516), .ZN(n3490) );
  NOR2_X2 U4442 ( .A1(n3490), .A2(n4346), .ZN(n4314) );
  AOI22_X1 U4443 ( .A1(n3571), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4049), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3464) );
  AOI22_X1 U4444 ( .A1(n3584), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3544), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3463) );
  AOI22_X1 U4445 ( .A1(n3597), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3852), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3471) );
  AOI22_X1 U4446 ( .A1(n4050), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3467), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3470) );
  AOI22_X1 U4447 ( .A1(n3573), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3545), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3469) );
  NOR2_X1 U4448 ( .A1(n4354), .A2(n3204), .ZN(n3474) );
  NAND2_X1 U4449 ( .A1(n3477), .A2(n3476), .ZN(n3480) );
  INV_X1 U4450 ( .A(n3478), .ZN(n3479) );
  OAI21_X1 U4451 ( .B1(n3481), .B2(n3480), .A(n3479), .ZN(n5355) );
  INV_X1 U4452 ( .A(n5355), .ZN(n5361) );
  NAND2_X1 U4453 ( .A1(n3641), .A2(n3205), .ZN(n3517) );
  NAND2_X1 U4454 ( .A1(n3516), .A2(n3482), .ZN(n3889) );
  OAI21_X1 U4455 ( .B1(n3208), .B2(n3483), .A(n3525), .ZN(n3484) );
  OAI21_X1 U4456 ( .B1(n3517), .B2(n3889), .A(n3484), .ZN(n3486) );
  NAND2_X2 U4457 ( .A1(n3203), .A2(n3641), .ZN(n4537) );
  AND2_X2 U4458 ( .A1(n3486), .A2(n3514), .ZN(n3506) );
  NAND2_X1 U4459 ( .A1(n3506), .A2(n3511), .ZN(n3527) );
  NOR2_X1 U4460 ( .A1(n5354), .A2(n6461), .ZN(n3487) );
  NAND2_X1 U4461 ( .A1(n5361), .A2(n3487), .ZN(n4442) );
  NOR2_X1 U4462 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6471) );
  NAND3_X1 U4463 ( .A1(STATE2_REG_0__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), 
        .A3(n6471), .ZN(n6459) );
  NAND2_X1 U4464 ( .A1(n6567), .A2(n5155), .ZN(n6466) );
  INV_X1 U4465 ( .A(n6466), .ZN(n6474) );
  NAND3_X1 U4466 ( .A1(n6474), .A2(STATE2_REG_1__SCAN_IN), .A3(n6564), .ZN(
        n6468) );
  NAND2_X1 U4467 ( .A1(n6736), .A2(n6547), .ZN(n4512) );
  NAND3_X1 U4468 ( .A1(n6459), .A2(n6468), .A3(n6175), .ZN(n3488) );
  NOR2_X1 U4469 ( .A1(n4415), .A2(n5080), .ZN(n4191) );
  NAND2_X1 U4470 ( .A1(n4416), .A2(n4191), .ZN(n3489) );
  INV_X1 U4471 ( .A(n4537), .ZN(n3491) );
  AOI21_X2 U4472 ( .B1(n3491), .B2(n3592), .A(n3490), .ZN(n3508) );
  XNOR2_X1 U4473 ( .A(STATE_REG_1__SCAN_IN), .B(STATE_REG_2__SCAN_IN), .ZN(
        n4184) );
  NAND2_X1 U4474 ( .A1(n4702), .A2(n4184), .ZN(n3523) );
  AOI21_X1 U4475 ( .B1(n3208), .B2(n3523), .A(n4354), .ZN(n3492) );
  NAND2_X1 U4476 ( .A1(n3508), .A2(n3492), .ZN(n3495) );
  NAND2_X2 U4477 ( .A1(n4702), .A2(n3493), .ZN(n4345) );
  OAI21_X1 U4478 ( .B1(n3495), .B2(n3507), .A(STATE2_REG_0__SCAN_IN), .ZN(
        n3500) );
  INV_X1 U4479 ( .A(n3610), .ZN(n3497) );
  NAND2_X1 U4480 ( .A1(n3500), .A2(n3499), .ZN(n3533) );
  NAND2_X1 U4481 ( .A1(n3533), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3505) );
  INV_X1 U4482 ( .A(n3662), .ZN(n3502) );
  INV_X1 U4483 ( .A(n4392), .ZN(n3501) );
  MUX2_X1 U4484 ( .A(n3502), .B(n3501), .S(n6430), .Z(n3503) );
  INV_X1 U4485 ( .A(n3503), .ZN(n3504) );
  INV_X1 U4486 ( .A(n3507), .ZN(n3522) );
  AOI21_X1 U4487 ( .B1(n4537), .B2(n4346), .A(n4605), .ZN(n3509) );
  NAND2_X1 U4488 ( .A1(n4316), .A2(n3509), .ZN(n3510) );
  NAND2_X1 U4489 ( .A1(n3510), .A2(n3401), .ZN(n3521) );
  INV_X1 U4490 ( .A(n3511), .ZN(n3513) );
  INV_X1 U4491 ( .A(n3514), .ZN(n3515) );
  NAND4_X1 U4492 ( .A1(n4605), .A2(n4593), .A3(n3516), .A4(n4346), .ZN(n3518)
         );
  NOR2_X1 U4493 ( .A1(n4512), .A2(n6567), .ZN(n6464) );
  INV_X1 U4494 ( .A(n3523), .ZN(n3529) );
  NAND3_X1 U4495 ( .A1(n4605), .A2(n3205), .A3(n3208), .ZN(n4474) );
  OR2_X2 U4496 ( .A1(n4474), .A2(n3524), .ZN(n4533) );
  INV_X1 U4497 ( .A(n4533), .ZN(n3526) );
  NAND2_X1 U4498 ( .A1(n3526), .A2(n5275), .ZN(n4347) );
  XNOR2_X1 U4499 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n5146) );
  OAI22_X1 U4500 ( .A1(n4392), .A2(n5146), .B1(n3662), .B2(n6436), .ZN(n3534)
         );
  OR2_X1 U4501 ( .A1(n3534), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3530)
         );
  NAND2_X1 U4502 ( .A1(n3613), .A2(n3611), .ZN(n3538) );
  NAND2_X1 U4503 ( .A1(n3532), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3537) );
  NAND2_X1 U4504 ( .A1(n3659), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3536) );
  INV_X1 U4505 ( .A(n3534), .ZN(n3535) );
  NAND3_X1 U4506 ( .A1(n3537), .A2(n3536), .A3(n3535), .ZN(n3612) );
  NAND2_X1 U4507 ( .A1(n3538), .A2(n3612), .ZN(n3656) );
  NAND2_X1 U4508 ( .A1(n3659), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3543) );
  NAND2_X1 U4509 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n3539) );
  NAND2_X1 U4510 ( .A1(n3539), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3540) );
  NOR2_X1 U4511 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n6436), .ZN(n4953)
         );
  NAND2_X1 U4512 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4953), .ZN(n4950) );
  OAI22_X1 U4513 ( .A1(n4392), .A2(n4652), .B1(n3662), .B2(n4859), .ZN(n3541)
         );
  INV_X1 U4514 ( .A(n3541), .ZN(n3542) );
  XNOR2_X1 U4515 ( .A(n3656), .B(n3657), .ZN(n4589) );
  AOI22_X1 U4516 ( .A1(n4131), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4148), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3549) );
  AOI22_X1 U4517 ( .A1(n4150), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3197), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3548) );
  AOI22_X1 U4518 ( .A1(n4158), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3896), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3547) );
  AOI22_X1 U4519 ( .A1(n4160), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4159), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3546) );
  NAND4_X1 U4520 ( .A1(n3549), .A2(n3548), .A3(n3547), .A4(n3546), .ZN(n3556)
         );
  AOI22_X1 U4521 ( .A1(n4156), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3852), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3554) );
  AOI22_X1 U4522 ( .A1(n4049), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4157), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3553) );
  AOI22_X1 U4523 ( .A1(n3943), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3552) );
  AOI22_X1 U4524 ( .A1(n3988), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n4735), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3551) );
  NAND4_X1 U4525 ( .A1(n3554), .A2(n3553), .A3(n3552), .A4(n3551), .ZN(n3555)
         );
  NOR2_X1 U4526 ( .A1(n3615), .A2(n4235), .ZN(n3557) );
  NAND2_X1 U4527 ( .A1(n3744), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3558) );
  OAI21_X1 U4528 ( .B1(n4235), .B2(n3610), .A(n3558), .ZN(n3559) );
  INV_X1 U4529 ( .A(n3620), .ZN(n3618) );
  INV_X1 U4530 ( .A(n3561), .ZN(n3564) );
  INV_X1 U4531 ( .A(n3562), .ZN(n3563) );
  NAND2_X1 U4532 ( .A1(n3564), .A2(n3563), .ZN(n3565) );
  NAND2_X1 U4533 ( .A1(n3613), .A2(n3565), .ZN(n3643) );
  INV_X1 U4534 ( .A(n3615), .ZN(n4473) );
  AOI22_X1 U4535 ( .A1(n4131), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4157), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3570) );
  AOI22_X1 U4536 ( .A1(INSTQUEUE_REG_15__7__SCAN_IN), .A2(n4148), .B1(n3197), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3569) );
  AOI22_X1 U4537 ( .A1(INSTQUEUE_REG_12__7__SCAN_IN), .A2(n4049), .B1(n4055), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3568) );
  AOI22_X1 U4538 ( .A1(n3896), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n4160), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3567) );
  NAND4_X1 U4539 ( .A1(n3570), .A2(n3569), .A3(n3568), .A4(n3567), .ZN(n3579)
         );
  AOI22_X1 U4540 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n4156), .B1(n3988), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3577) );
  AOI22_X1 U4541 ( .A1(INSTQUEUE_REG_10__7__SCAN_IN), .A2(n4150), .B1(n3852), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3576) );
  AOI22_X1 U4542 ( .A1(n3943), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4735), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3575) );
  AOI22_X1 U4543 ( .A1(n4158), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3545), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3574) );
  NAND4_X1 U4544 ( .A1(n3577), .A2(n3576), .A3(n3575), .A4(n3574), .ZN(n3578)
         );
  AOI22_X1 U4545 ( .A1(n4156), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3852), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3583) );
  AOI22_X1 U4546 ( .A1(n3197), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4148), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3582) );
  AOI22_X1 U4547 ( .A1(n3988), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n4735), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3581) );
  AOI22_X1 U4548 ( .A1(n4150), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3545), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3580) );
  NAND4_X1 U4549 ( .A1(n3583), .A2(n3582), .A3(n3581), .A4(n3580), .ZN(n3590)
         );
  AOI22_X1 U4550 ( .A1(n4049), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4157), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3588) );
  AOI22_X1 U4551 ( .A1(n4158), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4131), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3587) );
  AOI22_X1 U4552 ( .A1(n3943), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3586) );
  AOI22_X1 U4553 ( .A1(n3896), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n4160), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3585) );
  NAND4_X1 U4554 ( .A1(n3588), .A2(n3587), .A3(n3586), .A4(n3585), .ZN(n3589)
         );
  XNOR2_X1 U4555 ( .A(n4284), .B(n4220), .ZN(n3591) );
  NAND2_X1 U4556 ( .A1(n4473), .A2(n3591), .ZN(n3635) );
  OAI21_X2 U4557 ( .B1(n3643), .B2(STATE2_REG_0__SCAN_IN), .A(n3635), .ZN(
        n3633) );
  INV_X1 U4558 ( .A(n4220), .ZN(n3595) );
  NAND2_X1 U4559 ( .A1(n3744), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3594) );
  AOI21_X1 U4560 ( .B1(n3592), .B2(n4274), .A(n6567), .ZN(n3593) );
  OAI211_X1 U4561 ( .C1(n3595), .C2(n4555), .A(n3594), .B(n3593), .ZN(n3636)
         );
  NAND2_X1 U4562 ( .A1(n3633), .A2(n3636), .ZN(n3596) );
  NAND2_X1 U4563 ( .A1(n3596), .A2(n4281), .ZN(n3627) );
  AOI22_X1 U4564 ( .A1(n4156), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3852), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3601) );
  AOI22_X1 U4565 ( .A1(n4131), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4157), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3600) );
  AOI22_X1 U4566 ( .A1(n4150), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3197), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3599) );
  AOI22_X1 U4567 ( .A1(n3943), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3598) );
  NAND4_X1 U4568 ( .A1(n3601), .A2(n3600), .A3(n3599), .A4(n3598), .ZN(n3607)
         );
  AOI22_X1 U4569 ( .A1(n4049), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4148), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3605) );
  AOI22_X1 U4570 ( .A1(n4158), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3896), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3604) );
  AOI22_X1 U4571 ( .A1(n3988), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n4735), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3603) );
  AOI22_X1 U4572 ( .A1(n4160), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n4159), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3602) );
  NAND4_X1 U4573 ( .A1(n3605), .A2(n3604), .A3(n3603), .A4(n3602), .ZN(n3606)
         );
  OR2_X1 U4574 ( .A1(n3615), .A2(n4274), .ZN(n3609) );
  NAND2_X1 U4575 ( .A1(n3744), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3608) );
  OAI211_X1 U4576 ( .C1(n3610), .C2(n3616), .A(n3609), .B(n3608), .ZN(n3626)
         );
  NAND2_X1 U4577 ( .A1(n3211), .A2(n3611), .ZN(n3614) );
  OAI21_X1 U4578 ( .B1(n3627), .B2(n3626), .A(n3625), .ZN(n3617) );
  NAND2_X1 U4579 ( .A1(n3618), .A2(n3617), .ZN(n3621) );
  INV_X1 U4580 ( .A(n3873), .ZN(n3623) );
  NAND2_X1 U4581 ( .A1(n3624), .A2(n4096), .ZN(n4543) );
  NAND2_X1 U4582 ( .A1(n4585), .A2(n3873), .ZN(n3632) );
  INV_X1 U4583 ( .A(EAX_REG_1__SCAN_IN), .ZN(n3629) );
  INV_X1 U4584 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n5096) );
  OAI22_X1 U4585 ( .A1(n4171), .A2(n3629), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5096), .ZN(n3630) );
  AOI21_X1 U4586 ( .B1(n3685), .B2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(n3630), 
        .ZN(n3631) );
  NAND2_X1 U4587 ( .A1(n3632), .A2(n3631), .ZN(n4492) );
  INV_X1 U4588 ( .A(n3633), .ZN(n3634) );
  NAND2_X1 U4589 ( .A1(n3634), .A2(n3636), .ZN(n3640) );
  INV_X1 U4590 ( .A(n3635), .ZN(n3638) );
  NAND2_X1 U4591 ( .A1(n3641), .A2(n3516), .ZN(n3642) );
  OAI21_X1 U4592 ( .B1(n4218), .B2(n3642), .A(STATE2_REG_2__SCAN_IN), .ZN(
        n4479) );
  INV_X1 U4593 ( .A(n6267), .ZN(n4860) );
  INV_X1 U4594 ( .A(n3685), .ZN(n3704) );
  AOI22_X1 U4595 ( .A1(n3701), .A2(EAX_REG_0__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n5155), .ZN(n3644) );
  OAI21_X1 U4596 ( .B1(n3232), .B2(n3704), .A(n3644), .ZN(n3645) );
  AOI21_X1 U4597 ( .B1(n4860), .B2(n3873), .A(n3645), .ZN(n3646) );
  OR2_X1 U4598 ( .A1(n4479), .A2(n3646), .ZN(n4480) );
  INV_X1 U4599 ( .A(n3646), .ZN(n4481) );
  OR2_X1 U4600 ( .A1(n4481), .A2(n4145), .ZN(n3647) );
  NAND2_X1 U4601 ( .A1(n4480), .A2(n3647), .ZN(n4493) );
  NAND2_X1 U4602 ( .A1(n4492), .A2(n4493), .ZN(n4495) );
  INV_X1 U4603 ( .A(EAX_REG_2__SCAN_IN), .ZN(n3649) );
  OAI21_X1 U4604 ( .B1(PHYADDRPOINTER_REG_2__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_1__SCAN_IN), .A(n3680), .ZN(n6156) );
  AOI22_X1 U4605 ( .A1(n6156), .A2(n4176), .B1(n4177), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3648) );
  OAI21_X1 U4606 ( .B1(n4171), .B2(n3649), .A(n3648), .ZN(n3650) );
  AOI21_X1 U4607 ( .B1(n3685), .B2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n3650), 
        .ZN(n3651) );
  NAND2_X1 U4608 ( .A1(n4543), .A2(n4542), .ZN(n3655) );
  INV_X1 U4609 ( .A(n4495), .ZN(n3653) );
  INV_X1 U4610 ( .A(n3651), .ZN(n3652) );
  NAND2_X1 U4611 ( .A1(n3653), .A2(n3652), .ZN(n3654) );
  NAND2_X2 U4612 ( .A1(n3655), .A2(n3654), .ZN(n4540) );
  INV_X1 U4613 ( .A(n3656), .ZN(n3658) );
  NAND2_X1 U4614 ( .A1(n3659), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3665) );
  NAND3_X1 U4615 ( .A1(n6441), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6307) );
  INV_X1 U4616 ( .A(n6307), .ZN(n3660) );
  NAND2_X1 U4617 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n3660), .ZN(n4692) );
  NAND2_X1 U4618 ( .A1(n6441), .A2(n4692), .ZN(n3661) );
  NAND3_X1 U4619 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n4840) );
  INV_X1 U4620 ( .A(n4840), .ZN(n4595) );
  NAND2_X1 U4621 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4595), .ZN(n4798) );
  NAND2_X1 U4622 ( .A1(n3661), .A2(n4798), .ZN(n4647) );
  OAI22_X1 U4623 ( .A1(n4392), .A2(n4647), .B1(n3662), .B2(n6441), .ZN(n3663)
         );
  INV_X1 U4624 ( .A(n3663), .ZN(n3664) );
  NAND2_X1 U4625 ( .A1(n4588), .A2(n6567), .ZN(n3679) );
  AOI22_X1 U4626 ( .A1(n4131), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4148), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3671) );
  AOI22_X1 U4627 ( .A1(n4150), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3197), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3670) );
  AOI22_X1 U4628 ( .A1(n4158), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3896), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3669) );
  AOI22_X1 U4629 ( .A1(n4160), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n4159), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3668) );
  NAND4_X1 U4630 ( .A1(n3671), .A2(n3670), .A3(n3669), .A4(n3668), .ZN(n3677)
         );
  INV_X1 U4631 ( .A(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n6804) );
  AOI22_X1 U4632 ( .A1(n4156), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3852), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3675) );
  AOI22_X1 U4633 ( .A1(n4049), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4157), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3674) );
  AOI22_X1 U4634 ( .A1(n3943), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3673) );
  AOI22_X1 U4635 ( .A1(n3988), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n4735), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3672) );
  NAND4_X1 U4636 ( .A1(n3675), .A2(n3674), .A3(n3673), .A4(n3672), .ZN(n3676)
         );
  AOI22_X1 U4637 ( .A1(n3750), .A2(n4244), .B1(INSTQUEUE_REG_0__3__SCAN_IN), 
        .B2(n3744), .ZN(n3678) );
  NAND2_X1 U4638 ( .A1(n3202), .A2(n3873), .ZN(n3687) );
  INV_X1 U4639 ( .A(EAX_REG_3__SCAN_IN), .ZN(n3683) );
  OAI21_X1 U4640 ( .B1(PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n3681), .A(n3705), 
        .ZN(n6146) );
  AOI22_X1 U4641 ( .A1(PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n4177), .B1(n4176), 
        .B2(n6146), .ZN(n3682) );
  OAI21_X1 U4642 ( .B1(n4171), .B2(n3683), .A(n3682), .ZN(n3684) );
  AOI21_X1 U4643 ( .B1(n3685), .B2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(n3684), 
        .ZN(n3686) );
  NAND2_X1 U4644 ( .A1(n3687), .A2(n3686), .ZN(n4573) );
  NAND2_X1 U4645 ( .A1(n4540), .A2(n4573), .ZN(n4580) );
  INV_X1 U4646 ( .A(n4580), .ZN(n3710) );
  INV_X1 U4647 ( .A(n3200), .ZN(n3688) );
  AOI22_X1 U4648 ( .A1(n4131), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4148), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3692) );
  AOI22_X1 U4649 ( .A1(n4150), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3197), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3691) );
  AOI22_X1 U4650 ( .A1(n4158), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3896), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3690) );
  AOI22_X1 U4651 ( .A1(n4160), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n4159), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3689) );
  NAND4_X1 U4652 ( .A1(n3692), .A2(n3691), .A3(n3690), .A4(n3689), .ZN(n3698)
         );
  AOI22_X1 U4653 ( .A1(n4156), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4151), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3696) );
  AOI22_X1 U4654 ( .A1(n4149), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4157), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3695) );
  AOI22_X1 U4655 ( .A1(n3943), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3694) );
  AOI22_X1 U4656 ( .A1(n3988), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n4735), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3693) );
  NAND4_X1 U4657 ( .A1(n3696), .A2(n3695), .A3(n3694), .A4(n3693), .ZN(n3697)
         );
  NAND2_X1 U4658 ( .A1(n3750), .A2(n4261), .ZN(n3700) );
  NAND2_X1 U4659 ( .A1(n3744), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3699) );
  OAI21_X1 U4660 ( .B1(PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n6564), .A(n5155), 
        .ZN(n3703) );
  NAND2_X1 U4661 ( .A1(n3701), .A2(EAX_REG_4__SCAN_IN), .ZN(n3702) );
  OAI211_X1 U4662 ( .C1(n3704), .C2(n3436), .A(n3703), .B(n3702), .ZN(n3707)
         );
  AOI21_X1 U4663 ( .B1(n6897), .B2(n3705), .A(n3723), .ZN(n6133) );
  NAND2_X1 U4664 ( .A1(n6133), .A2(n4176), .ZN(n3706) );
  AND2_X1 U4665 ( .A1(n3707), .A2(n3706), .ZN(n3708) );
  AOI21_X1 U4666 ( .B1(n4243), .B2(n3873), .A(n3708), .ZN(n4579) );
  NAND2_X1 U4667 ( .A1(n3710), .A2(n3709), .ZN(n4578) );
  INV_X1 U4668 ( .A(n3731), .ZN(n3711) );
  NOR2_X1 U4669 ( .A1(n3728), .A2(n3711), .ZN(n3722) );
  AOI22_X1 U4670 ( .A1(n4131), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4148), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3715) );
  AOI22_X1 U4671 ( .A1(n4150), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3197), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3714) );
  AOI22_X1 U4672 ( .A1(n4158), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3896), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3713) );
  AOI22_X1 U4673 ( .A1(n4160), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n4159), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3712) );
  NAND4_X1 U4674 ( .A1(n3715), .A2(n3714), .A3(n3713), .A4(n3712), .ZN(n3721)
         );
  INV_X1 U4675 ( .A(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n6723) );
  AOI22_X1 U4676 ( .A1(n4156), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4151), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3719) );
  AOI22_X1 U4677 ( .A1(n4149), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4157), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3718) );
  AOI22_X1 U4678 ( .A1(n3943), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3717) );
  AOI22_X1 U4679 ( .A1(n3988), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n4735), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3716) );
  NAND4_X1 U4680 ( .A1(n3719), .A2(n3718), .A3(n3717), .A4(n3716), .ZN(n3720)
         );
  AOI22_X1 U4681 ( .A1(n3750), .A2(n4260), .B1(n3744), .B2(
        INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3729) );
  XNOR2_X1 U4682 ( .A(n3722), .B(n3729), .ZN(n4251) );
  INV_X1 U4683 ( .A(EAX_REG_5__SCAN_IN), .ZN(n4796) );
  OAI21_X1 U4684 ( .B1(n3723), .B2(PHYADDRPOINTER_REG_5__SCAN_IN), .A(n3755), 
        .ZN(n6128) );
  AOI22_X1 U4685 ( .A1(PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n4177), .B1(n4176), 
        .B2(n6128), .ZN(n3724) );
  OAI21_X1 U4686 ( .B1(n4171), .B2(n4796), .A(n3724), .ZN(n3725) );
  INV_X1 U4687 ( .A(n3729), .ZN(n3730) );
  AOI22_X1 U4688 ( .A1(n4131), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4148), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3737) );
  AOI22_X1 U4689 ( .A1(n4150), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3197), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3736) );
  AOI22_X1 U4690 ( .A1(n4158), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3896), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3735) );
  AOI22_X1 U4691 ( .A1(n4160), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n4159), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3734) );
  NAND4_X1 U4692 ( .A1(n3737), .A2(n3736), .A3(n3735), .A4(n3734), .ZN(n3743)
         );
  AOI22_X1 U4693 ( .A1(n4156), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4151), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3741) );
  AOI22_X1 U4694 ( .A1(n4149), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4157), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3740) );
  AOI22_X1 U4695 ( .A1(n3943), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3739) );
  AOI22_X1 U4696 ( .A1(n3988), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n4735), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3738) );
  NAND4_X1 U4697 ( .A1(n3741), .A2(n3740), .A3(n3739), .A4(n3738), .ZN(n3742)
         );
  AOI22_X1 U4698 ( .A1(n3750), .A2(n4272), .B1(n3744), .B2(
        INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3748) );
  NAND2_X1 U4699 ( .A1(n3749), .A2(n3748), .ZN(n4259) );
  OAI21_X1 U4700 ( .B1(PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n6564), .A(n5155), 
        .ZN(n3746) );
  NAND2_X1 U4701 ( .A1(n3701), .A2(EAX_REG_6__SCAN_IN), .ZN(n3745) );
  XNOR2_X1 U4702 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .B(n3755), .ZN(n6118) );
  AOI22_X1 U4703 ( .A1(n3746), .A2(n3745), .B1(n6118), .B2(n4176), .ZN(n3747)
         );
  INV_X1 U4704 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n6831) );
  NAND2_X1 U4705 ( .A1(n3750), .A2(n4274), .ZN(n3751) );
  OAI21_X1 U4706 ( .B1(n3752), .B2(n6831), .A(n3751), .ZN(n3753) );
  XNOR2_X1 U4707 ( .A(n4283), .B(n3753), .ZN(n4270) );
  NAND2_X1 U4708 ( .A1(n4270), .A2(n3873), .ZN(n3760) );
  OAI21_X1 U4709 ( .B1(n3756), .B2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n3776), 
        .ZN(n6113) );
  AOI22_X1 U4710 ( .A1(PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n4177), .B1(n4176), 
        .B2(n6113), .ZN(n3758) );
  NAND2_X1 U4711 ( .A1(n3701), .A2(EAX_REG_7__SCAN_IN), .ZN(n3757) );
  AND2_X1 U4712 ( .A1(n3758), .A2(n3757), .ZN(n3759) );
  XNOR2_X1 U4713 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .B(n3776), .ZN(n6102) );
  INV_X1 U4714 ( .A(n6102), .ZN(n3775) );
  AOI22_X1 U4715 ( .A1(n3988), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n4151), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3764) );
  AOI22_X1 U4716 ( .A1(n4158), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4150), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3763) );
  AOI22_X1 U4717 ( .A1(n4131), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4148), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3762) );
  AOI22_X1 U4718 ( .A1(n3943), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4735), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3761) );
  NAND4_X1 U4719 ( .A1(n3764), .A2(n3763), .A3(n3762), .A4(n3761), .ZN(n3770)
         );
  AOI22_X1 U4720 ( .A1(n4149), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4157), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3768) );
  AOI22_X1 U4721 ( .A1(n3197), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3896), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3767) );
  AOI22_X1 U4722 ( .A1(n4156), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3766) );
  AOI22_X1 U4723 ( .A1(n4160), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n4159), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3765) );
  NAND4_X1 U4724 ( .A1(n3768), .A2(n3767), .A3(n3766), .A4(n3765), .ZN(n3769)
         );
  OAI21_X1 U4725 ( .B1(n3770), .B2(n3769), .A(n3873), .ZN(n3773) );
  NAND2_X1 U4726 ( .A1(n3701), .A2(EAX_REG_8__SCAN_IN), .ZN(n3772) );
  NAND2_X1 U4727 ( .A1(PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n4177), .ZN(n3771)
         );
  NAND3_X1 U4728 ( .A1(n3773), .A2(n3772), .A3(n3771), .ZN(n3774) );
  AOI21_X1 U4729 ( .B1(n3775), .B2(n4176), .A(n3774), .ZN(n5116) );
  NOR2_X2 U4730 ( .A1(n5117), .A2(n5116), .ZN(n5124) );
  XNOR2_X1 U4731 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .B(n3801), .ZN(n6094) );
  AOI22_X1 U4732 ( .A1(n3701), .A2(EAX_REG_9__SCAN_IN), .B1(n4177), .B2(
        PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3789) );
  AOI22_X1 U4733 ( .A1(n4158), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4150), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3781) );
  AOI22_X1 U4734 ( .A1(n3943), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3780) );
  AOI22_X1 U4735 ( .A1(n4151), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4735), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3779) );
  AOI22_X1 U4736 ( .A1(n3896), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n4159), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3778) );
  NAND4_X1 U4737 ( .A1(n3781), .A2(n3780), .A3(n3779), .A4(n3778), .ZN(n3787)
         );
  AOI22_X1 U4738 ( .A1(n4156), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3988), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3785) );
  AOI22_X1 U4739 ( .A1(n4149), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4157), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3784) );
  AOI22_X1 U4740 ( .A1(n4131), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4148), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3783) );
  AOI22_X1 U4741 ( .A1(n3197), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4160), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3782) );
  NAND4_X1 U4742 ( .A1(n3785), .A2(n3784), .A3(n3783), .A4(n3782), .ZN(n3786)
         );
  OAI21_X1 U4743 ( .B1(n3787), .B2(n3786), .A(n3873), .ZN(n3788) );
  OAI211_X1 U4744 ( .C1(n6094), .C2(n4145), .A(n3789), .B(n3788), .ZN(n5123)
         );
  NAND2_X1 U4745 ( .A1(n5124), .A2(n5123), .ZN(n5122) );
  INV_X1 U4746 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n5216) );
  AOI22_X1 U4747 ( .A1(n4149), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4131), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3793) );
  AOI22_X1 U4748 ( .A1(n3197), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3896), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3792) );
  AOI22_X1 U4749 ( .A1(n3943), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3791) );
  AOI22_X1 U4750 ( .A1(n4151), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4735), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3790) );
  NAND4_X1 U4751 ( .A1(n3793), .A2(n3792), .A3(n3791), .A4(n3790), .ZN(n3799)
         );
  AOI22_X1 U4752 ( .A1(n4156), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3988), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3797) );
  AOI22_X1 U4753 ( .A1(n4158), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4150), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3796) );
  AOI22_X1 U4754 ( .A1(n4157), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4148), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3795) );
  AOI22_X1 U4755 ( .A1(n4160), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n4159), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3794) );
  NAND4_X1 U4756 ( .A1(n3797), .A2(n3796), .A3(n3795), .A4(n3794), .ZN(n3798)
         );
  OAI21_X1 U4757 ( .B1(n3799), .B2(n3798), .A(n3873), .ZN(n3800) );
  OAI21_X1 U4758 ( .B1(n5216), .B2(n4096), .A(n3800), .ZN(n3803) );
  XOR2_X1 U4759 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .B(n3804), .Z(n5926) );
  NOR2_X1 U4760 ( .A1(n5926), .A2(n4145), .ZN(n3802) );
  AOI211_X1 U4761 ( .C1(n3701), .C2(EAX_REG_10__SCAN_IN), .A(n3803), .B(n3802), 
        .ZN(n5143) );
  NOR2_X2 U4762 ( .A1(n5122), .A2(n5143), .ZN(n5142) );
  XNOR2_X1 U4763 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .B(n3829), .ZN(n6086)
         );
  AOI22_X1 U4764 ( .A1(n3701), .A2(EAX_REG_11__SCAN_IN), .B1(n4177), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3816) );
  AOI22_X1 U4765 ( .A1(n4150), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4151), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3808) );
  AOI22_X1 U4766 ( .A1(n3943), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3807) );
  AOI22_X1 U4767 ( .A1(n4158), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4159), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3806) );
  AOI22_X1 U4768 ( .A1(n3988), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n4735), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3805) );
  NAND4_X1 U4769 ( .A1(n3808), .A2(n3807), .A3(n3806), .A4(n3805), .ZN(n3814)
         );
  AOI22_X1 U4770 ( .A1(n4156), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4149), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3812) );
  AOI22_X1 U4771 ( .A1(n4131), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4157), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3811) );
  AOI22_X1 U4772 ( .A1(n3197), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4148), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3810) );
  AOI22_X1 U4773 ( .A1(n3896), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4160), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3809) );
  NAND4_X1 U4774 ( .A1(n3812), .A2(n3811), .A3(n3810), .A4(n3809), .ZN(n3813)
         );
  OAI21_X1 U4775 ( .B1(n3814), .B2(n3813), .A(n3873), .ZN(n3815) );
  OAI211_X1 U4776 ( .C1(n6086), .C2(n4145), .A(n3816), .B(n3815), .ZN(n5192)
         );
  INV_X1 U4777 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5234) );
  AOI22_X1 U4778 ( .A1(n4156), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4149), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3820) );
  AOI22_X1 U4779 ( .A1(n4157), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n4148), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3819) );
  AOI22_X1 U4780 ( .A1(n3943), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3818) );
  AOI22_X1 U4781 ( .A1(n4150), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4159), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3817) );
  NAND4_X1 U4782 ( .A1(n3820), .A2(n3819), .A3(n3818), .A4(n3817), .ZN(n3826)
         );
  AOI22_X1 U4783 ( .A1(n4131), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n4151), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3824) );
  AOI22_X1 U4784 ( .A1(n4158), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3197), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3823) );
  AOI22_X1 U4785 ( .A1(n3988), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n4735), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3822) );
  AOI22_X1 U4786 ( .A1(n3896), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n4160), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3821) );
  NAND4_X1 U4787 ( .A1(n3824), .A2(n3823), .A3(n3822), .A4(n3821), .ZN(n3825)
         );
  OAI21_X1 U4788 ( .B1(n3826), .B2(n3825), .A(n3873), .ZN(n3827) );
  OAI21_X1 U4789 ( .B1(n5234), .B2(n4096), .A(n3827), .ZN(n3831) );
  XOR2_X1 U4790 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .B(n3832), .Z(n5909) );
  NOR2_X1 U4791 ( .A1(n5909), .A2(n4145), .ZN(n3830) );
  AOI211_X1 U4792 ( .C1(n3701), .C2(EAX_REG_12__SCAN_IN), .A(n3831), .B(n3830), 
        .ZN(n5222) );
  XNOR2_X1 U4793 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .B(n3849), .ZN(n5901)
         );
  INV_X1 U4794 ( .A(EAX_REG_13__SCAN_IN), .ZN(n6019) );
  OAI222_X1 U4795 ( .A1(n4145), .A2(n5901), .B1(n4171), .B2(n6019), .C1(n3848), 
        .C2(n4096), .ZN(n3846) );
  AOI22_X1 U4796 ( .A1(n4131), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4148), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3837) );
  AOI22_X1 U4797 ( .A1(n4150), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3197), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3836) );
  AOI22_X1 U4798 ( .A1(n4158), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3896), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3835) );
  AOI22_X1 U4799 ( .A1(n4160), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n4159), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3834) );
  NAND4_X1 U4800 ( .A1(n3837), .A2(n3836), .A3(n3835), .A4(n3834), .ZN(n3843)
         );
  AOI22_X1 U4801 ( .A1(n4156), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4151), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3841) );
  AOI22_X1 U4802 ( .A1(n4149), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4157), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3840) );
  AOI22_X1 U4803 ( .A1(n3943), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3839) );
  AOI22_X1 U4804 ( .A1(n3988), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n4735), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3838) );
  NAND4_X1 U4805 ( .A1(n3841), .A2(n3840), .A3(n3839), .A4(n3838), .ZN(n3842)
         );
  OR2_X1 U4806 ( .A1(n3843), .A2(n3842), .ZN(n3844) );
  AND2_X1 U4807 ( .A1(n3873), .A2(n3844), .ZN(n5459) );
  NAND2_X1 U4808 ( .A1(n5221), .A2(n3846), .ZN(n3847) );
  AOI21_X1 U4809 ( .B1(n3851), .B2(n3850), .A(n3877), .ZN(n5888) );
  AOI22_X1 U4810 ( .A1(n3701), .A2(EAX_REG_14__SCAN_IN), .B1(n4177), .B2(
        PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3864) );
  AOI22_X1 U4811 ( .A1(n4156), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3988), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3856) );
  AOI22_X1 U4812 ( .A1(n4131), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3852), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3855) );
  AOI22_X1 U4813 ( .A1(n3943), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4735), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3854) );
  AOI22_X1 U4814 ( .A1(n3896), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4160), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3853) );
  NAND4_X1 U4815 ( .A1(n3856), .A2(n3855), .A3(n3854), .A4(n3853), .ZN(n3862)
         );
  AOI22_X1 U4816 ( .A1(n4157), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4148), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3860) );
  AOI22_X1 U4817 ( .A1(n4150), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3197), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3859) );
  AOI22_X1 U4818 ( .A1(n4149), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3858) );
  AOI22_X1 U4819 ( .A1(n4158), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4159), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3857) );
  NAND4_X1 U4820 ( .A1(n3860), .A2(n3859), .A3(n3858), .A4(n3857), .ZN(n3861)
         );
  OAI21_X1 U4821 ( .B1(n3862), .B2(n3861), .A(n3873), .ZN(n3863) );
  OAI211_X1 U4822 ( .C1(n5888), .C2(n4145), .A(n3864), .B(n3863), .ZN(n5450)
         );
  INV_X1 U4823 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n5305) );
  AOI22_X1 U4824 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n4150), .B1(n4158), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3868) );
  AOI22_X1 U4825 ( .A1(INSTQUEUE_REG_15__7__SCAN_IN), .A2(n4131), .B1(n3988), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3867) );
  AOI22_X1 U4826 ( .A1(n3943), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4735), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3866) );
  AOI22_X1 U4827 ( .A1(INSTQUEUE_REG_4__7__SCAN_IN), .A2(n3896), .B1(n4160), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3865) );
  NAND4_X1 U4828 ( .A1(n3868), .A2(n3867), .A3(n3866), .A4(n3865), .ZN(n3875)
         );
  AOI22_X1 U4829 ( .A1(n4149), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4151), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3872) );
  AOI22_X1 U4830 ( .A1(n4157), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4148), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3871) );
  AOI22_X1 U4831 ( .A1(n4156), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3870) );
  AOI22_X1 U4832 ( .A1(n3197), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4159), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3869) );
  NAND4_X1 U4833 ( .A1(n3872), .A2(n3871), .A3(n3870), .A4(n3869), .ZN(n3874)
         );
  OAI21_X1 U4834 ( .B1(n3875), .B2(n3874), .A(n3873), .ZN(n3876) );
  OAI21_X1 U4835 ( .B1(n5305), .B2(n4096), .A(n3876), .ZN(n3880) );
  OAI21_X1 U4836 ( .B1(PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n3877), .A(n3894), 
        .ZN(n3878) );
  INV_X1 U4837 ( .A(n3878), .ZN(n5882) );
  NOR2_X1 U4838 ( .A1(n5882), .A2(n4145), .ZN(n3879) );
  AOI211_X1 U4839 ( .C1(n3701), .C2(EAX_REG_15__SCAN_IN), .A(n3880), .B(n3879), 
        .ZN(n5302) );
  XNOR2_X1 U4840 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .B(n3894), .ZN(n5873)
         );
  AOI22_X1 U4841 ( .A1(n3701), .A2(EAX_REG_16__SCAN_IN), .B1(n4177), .B2(
        PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3893) );
  AOI22_X1 U4842 ( .A1(n3943), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3988), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3884) );
  AOI22_X1 U4843 ( .A1(n4149), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4157), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3883) );
  AOI22_X1 U4844 ( .A1(n4158), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3896), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3882) );
  AOI22_X1 U4845 ( .A1(n4160), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n4159), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3881) );
  NAND4_X1 U4846 ( .A1(n3884), .A2(n3883), .A3(n3882), .A4(n3881), .ZN(n3891)
         );
  AOI22_X1 U4847 ( .A1(n4156), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4151), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3888) );
  AOI22_X1 U4848 ( .A1(n4131), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n4148), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3887) );
  AOI22_X1 U4849 ( .A1(n4150), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3197), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3886) );
  AOI22_X1 U4850 ( .A1(n4055), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4735), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3885) );
  NAND4_X1 U4851 ( .A1(n3888), .A2(n3887), .A3(n3886), .A4(n3885), .ZN(n3890)
         );
  NOR2_X2 U4852 ( .A1(n5325), .A2(n6567), .ZN(n4173) );
  OAI21_X1 U4853 ( .B1(n3891), .B2(n3890), .A(n4173), .ZN(n3892) );
  OAI211_X1 U4854 ( .C1(n5873), .C2(n4145), .A(n3893), .B(n3892), .ZN(n5444)
         );
  OAI21_X1 U4855 ( .B1(PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n3895), .A(n4007), 
        .ZN(n5857) );
  AOI22_X1 U4856 ( .A1(n3701), .A2(EAX_REG_17__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n5155), .ZN(n3908) );
  AOI22_X1 U4857 ( .A1(n4157), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3988), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3900) );
  AOI22_X1 U4858 ( .A1(n4131), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n4148), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3899) );
  AOI22_X1 U4859 ( .A1(n4150), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3896), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3898) );
  AOI22_X1 U4860 ( .A1(n3943), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4735), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3897) );
  NAND4_X1 U4861 ( .A1(n3900), .A2(n3899), .A3(n3898), .A4(n3897), .ZN(n3906)
         );
  AOI22_X1 U4862 ( .A1(n4149), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4151), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3904) );
  AOI22_X1 U4863 ( .A1(n4158), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3197), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3903) );
  AOI22_X1 U4864 ( .A1(n4156), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3902) );
  AOI22_X1 U4865 ( .A1(n4160), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n4159), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3901) );
  NAND4_X1 U4866 ( .A1(n3904), .A2(n3903), .A3(n3902), .A4(n3901), .ZN(n3905)
         );
  OAI21_X1 U4867 ( .B1(n3906), .B2(n3905), .A(n4173), .ZN(n3907) );
  NAND3_X1 U4868 ( .A1(n4145), .A2(n3908), .A3(n3907), .ZN(n3909) );
  OAI21_X1 U4869 ( .B1(n4145), .B2(n5857), .A(n3909), .ZN(n5435) );
  INV_X1 U4870 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3910) );
  INV_X1 U4871 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5733) );
  NOR2_X1 U4872 ( .A1(n3911), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n3912)
         );
  OR2_X1 U4873 ( .A1(n3975), .A2(n3912), .ZN(n5723) );
  INV_X1 U4874 ( .A(n5723), .ZN(n3926) );
  INV_X1 U4875 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5715) );
  AOI22_X1 U4876 ( .A1(n4055), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4156), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3916) );
  AOI22_X1 U4877 ( .A1(n4157), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4151), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3915) );
  AOI22_X1 U4878 ( .A1(n4158), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4148), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3914) );
  AOI22_X1 U4879 ( .A1(n4160), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n4159), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3913) );
  NAND4_X1 U4880 ( .A1(n3916), .A2(n3915), .A3(n3914), .A4(n3913), .ZN(n3922)
         );
  AOI22_X1 U4881 ( .A1(n4735), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3943), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3920) );
  AOI22_X1 U4882 ( .A1(n4149), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3988), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3919) );
  AOI22_X1 U4883 ( .A1(n4131), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n3197), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3918) );
  AOI22_X1 U4884 ( .A1(n3896), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4150), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3917) );
  NAND4_X1 U4885 ( .A1(n3920), .A2(n3919), .A3(n3918), .A4(n3917), .ZN(n3921)
         );
  OAI21_X1 U4886 ( .B1(n3922), .B2(n3921), .A(n4173), .ZN(n3923) );
  OAI211_X1 U4887 ( .C1(n5715), .C2(STATE2_REG_2__SCAN_IN), .A(n3923), .B(
        n4145), .ZN(n3924) );
  AOI21_X1 U4888 ( .B1(n3701), .B2(EAX_REG_21__SCAN_IN), .A(n3924), .ZN(n3925)
         );
  AOI21_X1 U4889 ( .B1(n3926), .B2(n4176), .A(n3925), .ZN(n5407) );
  INV_X1 U4890 ( .A(EAX_REG_20__SCAN_IN), .ZN(n3940) );
  AOI22_X1 U4891 ( .A1(n4055), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3943), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3930) );
  AOI22_X1 U4892 ( .A1(n3988), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n4151), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3929) );
  AOI22_X1 U4893 ( .A1(n4149), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4150), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3928) );
  AOI22_X1 U4894 ( .A1(n3896), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n4159), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3927) );
  NAND4_X1 U4895 ( .A1(n3930), .A2(n3929), .A3(n3928), .A4(n3927), .ZN(n3936)
         );
  AOI22_X1 U4896 ( .A1(n4735), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n4156), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3934) );
  AOI22_X1 U4897 ( .A1(n4131), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n4157), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3933) );
  AOI22_X1 U4898 ( .A1(n3197), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4148), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3932) );
  AOI22_X1 U4899 ( .A1(n4158), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4160), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3931) );
  NAND4_X1 U4900 ( .A1(n3934), .A2(n3933), .A3(n3932), .A4(n3931), .ZN(n3935)
         );
  AOI221_X1 U4901 ( .B1(n3936), .B2(n4173), .C1(n3935), .C2(n4173), .A(n4176), 
        .ZN(n3937) );
  INV_X1 U4902 ( .A(n3937), .ZN(n3938) );
  AOI21_X1 U4903 ( .B1(n5155), .B2(PHYADDRPOINTER_REG_20__SCAN_IN), .A(n3938), 
        .ZN(n3939) );
  OAI21_X1 U4904 ( .B1(n4171), .B2(n3940), .A(n3939), .ZN(n3942) );
  XNOR2_X1 U4905 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .B(n3959), .ZN(n5724)
         );
  NAND2_X1 U4906 ( .A1(n4176), .A2(n5724), .ZN(n3941) );
  INV_X1 U4907 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5507) );
  XNOR2_X1 U4908 ( .A(n3975), .B(n5507), .ZN(n5707) );
  NAND2_X1 U4909 ( .A1(n5707), .A2(n4176), .ZN(n3958) );
  AOI22_X1 U4910 ( .A1(n4156), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4157), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3947) );
  AOI22_X1 U4911 ( .A1(n3943), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3946) );
  AOI22_X1 U4912 ( .A1(n4160), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n4159), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3945) );
  AOI22_X1 U4913 ( .A1(n3988), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4735), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3944) );
  NAND4_X1 U4914 ( .A1(n3947), .A2(n3946), .A3(n3945), .A4(n3944), .ZN(n3953)
         );
  AOI22_X1 U4915 ( .A1(n4149), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4151), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3951) );
  AOI22_X1 U4916 ( .A1(n4131), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n4148), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3950) );
  AOI22_X1 U4917 ( .A1(n4150), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3197), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3949) );
  AOI22_X1 U4918 ( .A1(n4158), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3896), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3948) );
  NAND4_X1 U4919 ( .A1(n3951), .A2(n3950), .A3(n3949), .A4(n3948), .ZN(n3952)
         );
  OAI21_X1 U4920 ( .B1(n3953), .B2(n3952), .A(n4173), .ZN(n3956) );
  AOI21_X1 U4921 ( .B1(n5155), .B2(PHYADDRPOINTER_REG_22__SCAN_IN), .A(n4176), 
        .ZN(n3955) );
  NAND2_X1 U4922 ( .A1(n3701), .A2(EAX_REG_22__SCAN_IN), .ZN(n3954) );
  NAND3_X1 U4923 ( .A1(n3956), .A2(n3955), .A3(n3954), .ZN(n3957) );
  NAND2_X1 U4924 ( .A1(n5401), .A2(n5403), .ZN(n3974) );
  OAI21_X1 U4925 ( .B1(n3960), .B2(PHYADDRPOINTER_REG_19__SCAN_IN), .A(n3959), 
        .ZN(n5781) );
  AOI22_X1 U4926 ( .A1(n3701), .A2(EAX_REG_19__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n5155), .ZN(n3972) );
  AOI22_X1 U4927 ( .A1(n3943), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3988), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3964) );
  AOI22_X1 U4928 ( .A1(n4149), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4151), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3963) );
  AOI22_X1 U4929 ( .A1(n4158), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3197), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3962) );
  AOI22_X1 U4930 ( .A1(n3896), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4159), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3961) );
  NAND4_X1 U4931 ( .A1(n3964), .A2(n3963), .A3(n3962), .A4(n3961), .ZN(n3970)
         );
  AOI22_X1 U4932 ( .A1(n4156), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4157), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3968) );
  AOI22_X1 U4933 ( .A1(n4131), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n4148), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3967) );
  AOI22_X1 U4934 ( .A1(n4055), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4735), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3966) );
  AOI22_X1 U4935 ( .A1(n4150), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4160), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3965) );
  NAND4_X1 U4936 ( .A1(n3968), .A2(n3967), .A3(n3966), .A4(n3965), .ZN(n3969)
         );
  OAI21_X1 U4937 ( .B1(n3970), .B2(n3969), .A(n4173), .ZN(n3971) );
  NAND3_X1 U4938 ( .A1(n4145), .A2(n3972), .A3(n3971), .ZN(n3973) );
  OAI21_X1 U4939 ( .B1(n4145), .B2(n5781), .A(n3973), .ZN(n5418) );
  OR2_X1 U4940 ( .A1(n3976), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n3977)
         );
  NAND2_X1 U4941 ( .A1(n4092), .A2(n3977), .ZN(n5697) );
  INV_X1 U4942 ( .A(n5697), .ZN(n4005) );
  AOI22_X1 U4943 ( .A1(n4157), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3988), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3981) );
  AOI22_X1 U4944 ( .A1(n4158), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3896), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3980) );
  AOI22_X1 U4945 ( .A1(n3943), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3979) );
  AOI22_X1 U4946 ( .A1(n4160), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n4159), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3978) );
  NAND4_X1 U4947 ( .A1(n3981), .A2(n3980), .A3(n3979), .A4(n3978), .ZN(n3987)
         );
  AOI22_X1 U4948 ( .A1(n4149), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3852), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3985) );
  AOI22_X1 U4949 ( .A1(n4131), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n4148), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3984) );
  AOI22_X1 U4950 ( .A1(INSTQUEUE_REG_12__7__SCAN_IN), .A2(n4150), .B1(n3197), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3983) );
  AOI22_X1 U4951 ( .A1(n4156), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4735), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3982) );
  NAND4_X1 U4952 ( .A1(n3985), .A2(n3984), .A3(n3983), .A4(n3982), .ZN(n3986)
         );
  NOR2_X1 U4953 ( .A1(n3987), .A2(n3986), .ZN(n4048) );
  AOI22_X1 U4954 ( .A1(n3988), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3852), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3992) );
  AOI22_X1 U4955 ( .A1(n4158), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4150), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3991) );
  AOI22_X1 U4956 ( .A1(n4149), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4157), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3990) );
  AOI22_X1 U4957 ( .A1(n3943), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3989) );
  NAND4_X1 U4958 ( .A1(n3992), .A2(n3991), .A3(n3990), .A4(n3989), .ZN(n3998)
         );
  AOI22_X1 U4959 ( .A1(n4131), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n4148), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3996) );
  AOI22_X1 U4960 ( .A1(n3197), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3896), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3995) );
  AOI22_X1 U4961 ( .A1(n4156), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4735), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3994) );
  AOI22_X1 U4962 ( .A1(n4160), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n4159), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3993) );
  NAND4_X1 U4963 ( .A1(n3996), .A2(n3995), .A3(n3994), .A4(n3993), .ZN(n3997)
         );
  NOR2_X1 U4964 ( .A1(n3998), .A2(n3997), .ZN(n4047) );
  XOR2_X1 U4965 ( .A(n4048), .B(n4047), .Z(n4003) );
  INV_X1 U4966 ( .A(EAX_REG_23__SCAN_IN), .ZN(n4561) );
  INV_X1 U4967 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n3999) );
  AOI21_X1 U4968 ( .B1(STATEBS16_REG_SCAN_IN), .B2(n3999), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4000) );
  INV_X1 U4969 ( .A(n4000), .ZN(n4001) );
  OAI21_X1 U4970 ( .B1(n4171), .B2(n4561), .A(n4001), .ZN(n4002) );
  AOI21_X1 U4971 ( .B1(n4173), .B2(n4003), .A(n4002), .ZN(n4004) );
  AOI21_X1 U4972 ( .B1(n4005), .B2(n4176), .A(n4004), .ZN(n4006) );
  INV_X1 U4973 ( .A(n4006), .ZN(n5395) );
  XNOR2_X1 U4974 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .B(n4007), .ZN(n5850)
         );
  AOI22_X1 U4975 ( .A1(n4156), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4151), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n4011) );
  AOI22_X1 U4976 ( .A1(n4149), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4157), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4010) );
  AOI22_X1 U4977 ( .A1(n3943), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4009) );
  AOI22_X1 U4978 ( .A1(n3988), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4735), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4008) );
  NAND4_X1 U4979 ( .A1(n4011), .A2(n4010), .A3(n4009), .A4(n4008), .ZN(n4017)
         );
  AOI22_X1 U4980 ( .A1(n4131), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4148), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4015) );
  AOI22_X1 U4981 ( .A1(n4150), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3197), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n4014) );
  AOI22_X1 U4982 ( .A1(n4158), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3896), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4013) );
  AOI22_X1 U4983 ( .A1(n4160), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n4159), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4012) );
  NAND4_X1 U4984 ( .A1(n4015), .A2(n4014), .A3(n4013), .A4(n4012), .ZN(n4016)
         );
  OR2_X1 U4985 ( .A1(n4017), .A2(n4016), .ZN(n4018) );
  AOI22_X1 U4986 ( .A1(n4173), .A2(n4018), .B1(n3701), .B2(EAX_REG_18__SCAN_IN), .ZN(n4020) );
  OAI21_X1 U4987 ( .B1(PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n6564), .A(n5155), 
        .ZN(n4019) );
  AOI22_X1 U4988 ( .A1(n4176), .A2(n5850), .B1(n4020), .B2(n4019), .ZN(n5431)
         );
  INV_X1 U4989 ( .A(n5431), .ZN(n4021) );
  NOR2_X1 U4990 ( .A1(n4022), .A2(n4021), .ZN(n4023) );
  INV_X1 U4991 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5265) );
  INV_X1 U4992 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4024) );
  NOR2_X1 U4993 ( .A1(n4025), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4026)
         );
  OR2_X1 U4994 ( .A1(n4124), .A2(n4026), .ZN(n5667) );
  AOI22_X1 U4995 ( .A1(n4158), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4150), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n4030) );
  AOI22_X1 U4996 ( .A1(n3197), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4151), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4029) );
  AOI22_X1 U4997 ( .A1(n3943), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4735), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4028) );
  AOI22_X1 U4998 ( .A1(n4160), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n4159), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4027) );
  NAND4_X1 U4999 ( .A1(n4030), .A2(n4029), .A3(n4028), .A4(n4027), .ZN(n4036)
         );
  AOI22_X1 U5000 ( .A1(n4156), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4149), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4034) );
  AOI22_X1 U5001 ( .A1(n4131), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n4157), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4033) );
  AOI22_X1 U5002 ( .A1(n4148), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3896), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4032) );
  AOI22_X1 U5003 ( .A1(n3988), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4031) );
  NAND4_X1 U5004 ( .A1(n4034), .A2(n4033), .A3(n4032), .A4(n4031), .ZN(n4035)
         );
  NOR2_X1 U5005 ( .A1(n4036), .A2(n4035), .ZN(n4116) );
  AOI22_X1 U5006 ( .A1(n4156), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4151), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4040) );
  AOI22_X1 U5007 ( .A1(n4149), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4157), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4039) );
  AOI22_X1 U5008 ( .A1(n3943), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4038) );
  AOI22_X1 U5009 ( .A1(n3988), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4735), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4037) );
  NAND4_X1 U5010 ( .A1(n4040), .A2(n4039), .A3(n4038), .A4(n4037), .ZN(n4046)
         );
  AOI22_X1 U5011 ( .A1(n4131), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4148), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4044) );
  AOI22_X1 U5012 ( .A1(n4150), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3197), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n4043) );
  AOI22_X1 U5013 ( .A1(n4158), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3896), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4042) );
  AOI22_X1 U5014 ( .A1(n4160), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4159), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4041) );
  NAND4_X1 U5015 ( .A1(n4044), .A2(n4043), .A3(n4042), .A4(n4041), .ZN(n4045)
         );
  NOR2_X1 U5016 ( .A1(n4046), .A2(n4045), .ZN(n4088) );
  OR2_X1 U5017 ( .A1(n4048), .A2(n4047), .ZN(n4095) );
  AOI22_X1 U5018 ( .A1(n4150), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3896), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4054) );
  AOI22_X1 U5019 ( .A1(n4149), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4148), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4053) );
  AOI22_X1 U5020 ( .A1(n4156), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3197), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n4052) );
  AOI22_X1 U5021 ( .A1(n3943), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4160), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4051) );
  NAND4_X1 U5022 ( .A1(n4054), .A2(n4053), .A3(n4052), .A4(n4051), .ZN(n4061)
         );
  AOI22_X1 U5023 ( .A1(n3988), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n4151), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n4059) );
  AOI22_X1 U5024 ( .A1(n4131), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n4157), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4058) );
  AOI22_X1 U5025 ( .A1(n4158), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4057) );
  AOI22_X1 U5026 ( .A1(n4159), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4735), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4056) );
  NAND4_X1 U5027 ( .A1(n4059), .A2(n4058), .A3(n4057), .A4(n4056), .ZN(n4060)
         );
  NOR2_X1 U5028 ( .A1(n4061), .A2(n4060), .ZN(n4094) );
  OR2_X1 U5029 ( .A1(n4095), .A2(n4094), .ZN(n4087) );
  NOR2_X1 U5030 ( .A1(n4088), .A2(n4087), .ZN(n4077) );
  AOI22_X1 U5031 ( .A1(n4156), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4151), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4065) );
  AOI22_X1 U5032 ( .A1(n4149), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4157), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4064) );
  AOI22_X1 U5033 ( .A1(n3943), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4063) );
  AOI22_X1 U5034 ( .A1(n3988), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4735), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4062) );
  NAND4_X1 U5035 ( .A1(n4065), .A2(n4064), .A3(n4063), .A4(n4062), .ZN(n4071)
         );
  AOI22_X1 U5036 ( .A1(n4131), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n4148), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4069) );
  AOI22_X1 U5037 ( .A1(n4150), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3197), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n4068) );
  AOI22_X1 U5038 ( .A1(n4158), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3896), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4067) );
  AOI22_X1 U5039 ( .A1(n4160), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4159), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4066) );
  NAND4_X1 U5040 ( .A1(n4069), .A2(n4068), .A3(n4067), .A4(n4066), .ZN(n4070)
         );
  OR2_X1 U5041 ( .A1(n4071), .A2(n4070), .ZN(n4078) );
  NAND2_X1 U5042 ( .A1(n4077), .A2(n4078), .ZN(n4115) );
  XNOR2_X1 U5043 ( .A(n4116), .B(n4115), .ZN(n4074) );
  INV_X1 U5044 ( .A(n4173), .ZN(n4142) );
  INV_X1 U5045 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5491) );
  OAI21_X1 U5046 ( .B1(n5491), .B2(STATE2_REG_2__SCAN_IN), .A(n4145), .ZN(
        n4072) );
  AOI21_X1 U5047 ( .B1(n3701), .B2(EAX_REG_27__SCAN_IN), .A(n4072), .ZN(n4073)
         );
  OAI21_X1 U5048 ( .B1(n4074), .B2(n4142), .A(n4073), .ZN(n4075) );
  OAI21_X1 U5049 ( .B1(n5667), .B2(n4145), .A(n4075), .ZN(n4076) );
  INV_X1 U5050 ( .A(n4076), .ZN(n5377) );
  XOR2_X1 U5051 ( .A(n4078), .B(n4077), .Z(n4079) );
  AOI21_X1 U5052 ( .B1(n4079), .B2(n4173), .A(n4176), .ZN(n4082) );
  NAND2_X1 U5053 ( .A1(n5155), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4081)
         );
  NAND2_X1 U5054 ( .A1(n3701), .A2(EAX_REG_26__SCAN_IN), .ZN(n4080) );
  NAND3_X1 U5055 ( .A1(n4082), .A2(n4081), .A3(n4080), .ZN(n4084) );
  XNOR2_X1 U5056 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .B(n4085), .ZN(n5764)
         );
  NAND2_X1 U5057 ( .A1(n4176), .A2(n5764), .ZN(n4083) );
  NAND2_X1 U5058 ( .A1(n4084), .A2(n4083), .ZN(n5280) );
  OAI21_X1 U5059 ( .B1(PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n4086), .A(n4085), 
        .ZN(n5776) );
  XNOR2_X1 U5060 ( .A(n4088), .B(n4087), .ZN(n4090) );
  AOI22_X1 U5061 ( .A1(n3701), .A2(EAX_REG_25__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n5155), .ZN(n4089) );
  OAI21_X1 U5062 ( .B1(n4142), .B2(n4090), .A(n4089), .ZN(n4091) );
  AOI22_X1 U5063 ( .A1(n4176), .A2(n5776), .B1(n4091), .B2(n4145), .ZN(n5389)
         );
  OR2_X1 U5064 ( .A1(n5280), .A2(n5389), .ZN(n4103) );
  XNOR2_X1 U5065 ( .A(n4092), .B(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5689)
         );
  OR2_X1 U5066 ( .A1(n5689), .A2(n4145), .ZN(n4102) );
  AOI21_X1 U5067 ( .B1(n4094), .B2(n4095), .A(n4142), .ZN(n4093) );
  OAI21_X1 U5068 ( .B1(n4095), .B2(n4094), .A(n4093), .ZN(n4100) );
  INV_X1 U5069 ( .A(EAX_REG_24__SCAN_IN), .ZN(n4097) );
  OAI22_X1 U5070 ( .A1(n4171), .A2(n4097), .B1(n4096), .B2(n5265), .ZN(n4098)
         );
  INV_X1 U5071 ( .A(n4098), .ZN(n4099) );
  AND2_X1 U5072 ( .A1(n4100), .A2(n4099), .ZN(n4101) );
  NOR2_X1 U5073 ( .A1(n4103), .A2(n5267), .ZN(n5279) );
  AND2_X1 U5074 ( .A1(n5377), .A2(n5279), .ZN(n4104) );
  INV_X1 U5075 ( .A(n5380), .ZN(n4123) );
  INV_X1 U5076 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5485) );
  XNOR2_X1 U5077 ( .A(n4124), .B(n5485), .ZN(n5656) );
  NAND2_X1 U5078 ( .A1(n5656), .A2(n4176), .ZN(n4122) );
  AOI22_X1 U5079 ( .A1(n4156), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4151), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4108) );
  AOI22_X1 U5080 ( .A1(n4149), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4157), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4107) );
  AOI22_X1 U5081 ( .A1(n3943), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4106) );
  AOI22_X1 U5082 ( .A1(n3988), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4735), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4105) );
  NAND4_X1 U5083 ( .A1(n4108), .A2(n4107), .A3(n4106), .A4(n4105), .ZN(n4114)
         );
  AOI22_X1 U5084 ( .A1(n4131), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n4148), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4112) );
  AOI22_X1 U5085 ( .A1(n4150), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3197), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n4111) );
  AOI22_X1 U5086 ( .A1(n4158), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3896), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4110) );
  AOI22_X1 U5087 ( .A1(n4160), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n4159), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4109) );
  NAND4_X1 U5088 ( .A1(n4112), .A2(n4111), .A3(n4110), .A4(n4109), .ZN(n4113)
         );
  OR2_X1 U5089 ( .A1(n4114), .A2(n4113), .ZN(n4138) );
  NOR2_X1 U5090 ( .A1(n4116), .A2(n4115), .ZN(n4139) );
  XOR2_X1 U5091 ( .A(n4138), .B(n4139), .Z(n4117) );
  NAND2_X1 U5092 ( .A1(n4117), .A2(n4173), .ZN(n4120) );
  OAI21_X1 U5093 ( .B1(n5485), .B2(STATE2_REG_2__SCAN_IN), .A(n4145), .ZN(
        n4118) );
  AOI21_X1 U5094 ( .B1(n3701), .B2(EAX_REG_28__SCAN_IN), .A(n4118), .ZN(n4119)
         );
  NAND2_X1 U5095 ( .A1(n4120), .A2(n4119), .ZN(n4121) );
  OR2_X1 U5096 ( .A1(n4125), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4126)
         );
  NAND2_X1 U5097 ( .A1(n4181), .A2(n4126), .ZN(n5346) );
  AOI22_X1 U5098 ( .A1(n4149), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4148), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4130) );
  AOI22_X1 U5099 ( .A1(n4150), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3584), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4129) );
  AOI22_X1 U5100 ( .A1(n3943), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4128) );
  AOI22_X1 U5101 ( .A1(n4156), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4735), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4127) );
  NAND4_X1 U5102 ( .A1(n4130), .A2(n4129), .A3(n4128), .A4(n4127), .ZN(n4137)
         );
  AOI22_X1 U5103 ( .A1(n3988), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4151), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4135) );
  AOI22_X1 U5104 ( .A1(n4131), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n4157), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4134) );
  AOI22_X1 U5105 ( .A1(n4158), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3197), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n4133) );
  AOI22_X1 U5106 ( .A1(n4160), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4159), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4132) );
  NAND4_X1 U5107 ( .A1(n4135), .A2(n4134), .A3(n4133), .A4(n4132), .ZN(n4136)
         );
  NOR2_X1 U5108 ( .A1(n4137), .A2(n4136), .ZN(n4147) );
  NAND2_X1 U5109 ( .A1(n4139), .A2(n4138), .ZN(n4146) );
  XNOR2_X1 U5110 ( .A(n4147), .B(n4146), .ZN(n4143) );
  INV_X1 U5111 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n6884) );
  AOI21_X1 U5112 ( .B1(STATEBS16_REG_SCAN_IN), .B2(n6884), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4140) );
  AOI21_X1 U5113 ( .B1(n3701), .B2(EAX_REG_29__SCAN_IN), .A(n4140), .ZN(n4141)
         );
  OAI21_X1 U5114 ( .B1(n4143), .B2(n4142), .A(n4141), .ZN(n4144) );
  OAI21_X1 U5115 ( .B1(n5346), .B2(n4145), .A(n4144), .ZN(n4406) );
  XNOR2_X1 U5116 ( .A(n4181), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5651)
         );
  NOR2_X1 U5117 ( .A1(n4147), .A2(n4146), .ZN(n4168) );
  AOI22_X1 U5118 ( .A1(INSTQUEUE_REG_15__7__SCAN_IN), .A2(n4149), .B1(n4148), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4155) );
  AOI22_X1 U5119 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n4150), .B1(n3584), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4154) );
  AOI22_X1 U5120 ( .A1(n3943), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4153) );
  AOI22_X1 U5121 ( .A1(n4151), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4735), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4152) );
  NAND4_X1 U5122 ( .A1(n4155), .A2(n4154), .A3(n4153), .A4(n4152), .ZN(n4166)
         );
  AOI22_X1 U5123 ( .A1(n4156), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3988), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4164) );
  AOI22_X1 U5124 ( .A1(n4131), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n4157), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4163) );
  AOI22_X1 U5125 ( .A1(INSTQUEUE_REG_10__7__SCAN_IN), .A2(n4158), .B1(n3197), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n4162) );
  AOI22_X1 U5126 ( .A1(INSTQUEUE_REG_4__7__SCAN_IN), .A2(n4160), .B1(n4159), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4161) );
  NAND4_X1 U5127 ( .A1(n4164), .A2(n4163), .A3(n4162), .A4(n4161), .ZN(n4165)
         );
  NOR2_X1 U5128 ( .A1(n4166), .A2(n4165), .ZN(n4167) );
  XNOR2_X1 U5129 ( .A(n4168), .B(n4167), .ZN(n4174) );
  INV_X1 U5130 ( .A(EAX_REG_30__SCAN_IN), .ZN(n4170) );
  OAI21_X1 U5131 ( .B1(PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n6564), .A(n5155), 
        .ZN(n4169) );
  OAI21_X1 U5132 ( .B1(n4171), .B2(n4170), .A(n4169), .ZN(n4172) );
  AOI21_X1 U5133 ( .B1(n4174), .B2(n4173), .A(n4172), .ZN(n4175) );
  AOI21_X1 U5134 ( .B1(n5651), .B2(n4176), .A(n4175), .ZN(n4401) );
  NAND2_X1 U5135 ( .A1(n4407), .A2(n4401), .ZN(n4180) );
  AOI22_X1 U5136 ( .A1(n3701), .A2(EAX_REG_31__SCAN_IN), .B1(n4177), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4178) );
  INV_X1 U5137 ( .A(n4178), .ZN(n4179) );
  INV_X1 U5138 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n6707) );
  INV_X1 U5139 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4182) );
  NAND2_X1 U5140 ( .A1(n5953), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4413) );
  INV_X1 U5141 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6530) );
  INV_X1 U5142 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6523) );
  INV_X1 U5143 ( .A(REIP_REG_26__SCAN_IN), .ZN(n6526) );
  INV_X1 U5144 ( .A(REIP_REG_25__SCAN_IN), .ZN(n6525) );
  NOR3_X1 U5145 ( .A1(n6523), .A2(n6526), .A3(n6525), .ZN(n4199) );
  INV_X1 U5146 ( .A(n4199), .ZN(n4190) );
  NAND2_X1 U5147 ( .A1(REIP_REG_20__SCAN_IN), .A2(REIP_REG_19__SCAN_IN), .ZN(
        n4189) );
  NAND3_X1 U5148 ( .A1(REIP_REG_15__SCAN_IN), .A2(REIP_REG_17__SCAN_IN), .A3(
        REIP_REG_16__SCAN_IN), .ZN(n4188) );
  INV_X1 U5149 ( .A(REIP_REG_11__SCAN_IN), .ZN(n6503) );
  INV_X1 U5150 ( .A(REIP_REG_8__SCAN_IN), .ZN(n6499) );
  INV_X1 U5151 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6719) );
  NAND3_X1 U5152 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_3__SCAN_IN), .A3(
        REIP_REG_2__SCAN_IN), .ZN(n5985) );
  NOR2_X1 U5153 ( .A1(n6719), .A2(n5985), .ZN(n5974) );
  AND2_X1 U5154 ( .A1(REIP_REG_5__SCAN_IN), .A2(n5974), .ZN(n5954) );
  NAND3_X1 U5155 ( .A1(REIP_REG_7__SCAN_IN), .A2(REIP_REG_6__SCAN_IN), .A3(
        n5954), .ZN(n5941) );
  OR2_X1 U5156 ( .A1(n6499), .A2(n5941), .ZN(n5928) );
  NAND2_X1 U5157 ( .A1(REIP_REG_9__SCAN_IN), .A2(REIP_REG_10__SCAN_IN), .ZN(
        n5914) );
  NOR3_X1 U5158 ( .A1(n6503), .A2(n5928), .A3(n5914), .ZN(n4196) );
  INV_X1 U5159 ( .A(n4184), .ZN(n4185) );
  NAND2_X1 U5160 ( .A1(n4185), .A2(n6798), .ZN(n6481) );
  NAND2_X1 U5161 ( .A1(n4702), .A2(n6481), .ZN(n4325) );
  NOR2_X1 U5162 ( .A1(n5080), .A2(n4416), .ZN(n4186) );
  AND2_X1 U5163 ( .A1(n4555), .A2(n4186), .ZN(n4187) );
  NAND4_X1 U5164 ( .A1(REIP_REG_14__SCAN_IN), .A2(REIP_REG_13__SCAN_IN), .A3(
        REIP_REG_12__SCAN_IN), .A4(n5906), .ZN(n5866) );
  NAND4_X1 U5165 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .A4(n5706), .ZN(n5685) );
  NAND3_X1 U5166 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .A3(
        n5669), .ZN(n4424) );
  NOR2_X1 U5167 ( .A1(n6530), .A2(n4424), .ZN(n5648) );
  NAND2_X1 U5168 ( .A1(REIP_REG_30__SCAN_IN), .A2(n5648), .ZN(n4194) );
  INV_X1 U5169 ( .A(n4191), .ZN(n4193) );
  INV_X1 U5170 ( .A(n6481), .ZN(n4553) );
  NAND3_X1 U5171 ( .A1(n4553), .A2(n4324), .A3(n6564), .ZN(n6451) );
  INV_X1 U5172 ( .A(n6451), .ZN(n4192) );
  OR2_X1 U5173 ( .A1(n4345), .A2(n4192), .ZN(n4418) );
  OAI22_X1 U5174 ( .A1(n4194), .A2(REIP_REG_31__SCAN_IN), .B1(n4193), .B2(
        n4418), .ZN(n4195) );
  AOI21_X1 U5175 ( .B1(PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n5983), .A(n4195), 
        .ZN(n4204) );
  INV_X1 U5176 ( .A(REIP_REG_30__SCAN_IN), .ZN(n6537) );
  INV_X1 U5177 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6513) );
  NAND2_X1 U5178 ( .A1(n4196), .A2(n5953), .ZN(n5893) );
  NAND3_X1 U5179 ( .A1(REIP_REG_14__SCAN_IN), .A2(REIP_REG_13__SCAN_IN), .A3(
        REIP_REG_12__SCAN_IN), .ZN(n4197) );
  NOR2_X1 U5180 ( .A1(n5893), .A2(n4197), .ZN(n5864) );
  NAND4_X1 U5181 ( .A1(n5864), .A2(REIP_REG_15__SCAN_IN), .A3(
        REIP_REG_17__SCAN_IN), .A4(REIP_REG_16__SCAN_IN), .ZN(n5856) );
  NOR2_X1 U5182 ( .A1(n6513), .A2(n5856), .ZN(n5734) );
  NAND3_X1 U5183 ( .A1(n5734), .A2(REIP_REG_20__SCAN_IN), .A3(
        REIP_REG_19__SCAN_IN), .ZN(n5705) );
  NAND3_X1 U5184 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .ZN(n4198) );
  NOR2_X1 U5185 ( .A1(n5705), .A2(n4198), .ZN(n5684) );
  NAND2_X1 U5186 ( .A1(n5953), .A2(n5976), .ZN(n5894) );
  AOI21_X1 U5187 ( .B1(n5684), .B2(n4199), .A(n5865), .ZN(n5676) );
  AND2_X1 U5188 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .ZN(
        n4200) );
  NOR2_X1 U5189 ( .A1(n5976), .A2(n4200), .ZN(n4201) );
  NOR2_X1 U5190 ( .A1(n5676), .A2(n4201), .ZN(n5659) );
  NAND2_X1 U5191 ( .A1(REIP_REG_29__SCAN_IN), .A2(n5659), .ZN(n4202) );
  OAI21_X1 U5192 ( .B1(n6537), .B2(n4202), .A(n5894), .ZN(n5655) );
  INV_X1 U5193 ( .A(REIP_REG_31__SCAN_IN), .ZN(n6829) );
  INV_X1 U5194 ( .A(n4269), .ZN(n4280) );
  NAND2_X1 U5195 ( .A1(n4212), .A2(n4220), .ZN(n4236) );
  XNOR2_X1 U5196 ( .A(n4236), .B(n4235), .ZN(n4210) );
  NAND2_X1 U5197 ( .A1(n4593), .A2(n4208), .ZN(n4219) );
  INV_X1 U5198 ( .A(n4219), .ZN(n4209) );
  AOI21_X1 U5199 ( .B1(n4210), .B2(n6565), .A(n4209), .ZN(n4211) );
  OAI21_X2 U5200 ( .B1(n4584), .B2(n4280), .A(n4211), .ZN(n6150) );
  NAND2_X1 U5201 ( .A1(n6150), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4229)
         );
  NAND2_X1 U5202 ( .A1(n4585), .A2(n4269), .ZN(n4217) );
  OAI21_X1 U5203 ( .B1(n4220), .B2(n4212), .A(n4236), .ZN(n4214) );
  INV_X1 U5204 ( .A(n4354), .ZN(n4213) );
  OAI211_X1 U5205 ( .C1(n4214), .C2(n4345), .A(n4213), .B(n3204), .ZN(n4215)
         );
  INV_X1 U5206 ( .A(n4215), .ZN(n4216) );
  NAND2_X1 U5207 ( .A1(n4217), .A2(n4216), .ZN(n4547) );
  NAND2_X1 U5208 ( .A1(n4218), .A2(n4269), .ZN(n4223) );
  OAI21_X1 U5209 ( .B1(n4345), .B2(n4220), .A(n4219), .ZN(n4221) );
  INV_X1 U5210 ( .A(n4221), .ZN(n4222) );
  NAND2_X1 U5211 ( .A1(n4223), .A2(n4222), .ZN(n4483) );
  NAND2_X1 U5212 ( .A1(n4483), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4224)
         );
  NAND2_X1 U5213 ( .A1(n4224), .A2(n6234), .ZN(n4226) );
  AND2_X1 U5214 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4225) );
  NAND2_X1 U5215 ( .A1(n4483), .A2(n4225), .ZN(n4227) );
  INV_X1 U5216 ( .A(n4227), .ZN(n4228) );
  NAND2_X1 U5217 ( .A1(n4229), .A2(n6149), .ZN(n4233) );
  INV_X1 U5218 ( .A(n6150), .ZN(n4231) );
  INV_X1 U5219 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4230) );
  NAND2_X1 U5220 ( .A1(n4231), .A2(n4230), .ZN(n4232) );
  NAND2_X1 U5221 ( .A1(n4234), .A2(n4269), .ZN(n4240) );
  NAND2_X1 U5222 ( .A1(n4236), .A2(n4235), .ZN(n4245) );
  INV_X1 U5223 ( .A(n4244), .ZN(n4237) );
  XNOR2_X1 U5224 ( .A(n4245), .B(n4237), .ZN(n4238) );
  NAND2_X1 U5225 ( .A1(n4238), .A2(n6565), .ZN(n4239) );
  INV_X1 U5226 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n6802) );
  NAND2_X1 U5227 ( .A1(n6141), .A2(n6139), .ZN(n6140) );
  NAND2_X1 U5228 ( .A1(n4241), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4242)
         );
  NAND2_X1 U5229 ( .A1(n6140), .A2(n4242), .ZN(n6131) );
  NAND2_X1 U5230 ( .A1(n4243), .A2(n4269), .ZN(n4248) );
  NAND2_X1 U5231 ( .A1(n4245), .A2(n4244), .ZN(n4263) );
  XNOR2_X1 U5232 ( .A(n4263), .B(n4261), .ZN(n4246) );
  NAND2_X1 U5233 ( .A1(n4246), .A2(n6565), .ZN(n4247) );
  NAND2_X1 U5234 ( .A1(n6131), .A2(n6129), .ZN(n6130) );
  NAND2_X1 U5235 ( .A1(n4249), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4250)
         );
  NAND2_X1 U5236 ( .A1(n6130), .A2(n4250), .ZN(n4627) );
  NAND2_X1 U5237 ( .A1(n4251), .A2(n4269), .ZN(n4256) );
  INV_X1 U5238 ( .A(n4261), .ZN(n4252) );
  OR2_X1 U5239 ( .A1(n4263), .A2(n4252), .ZN(n4253) );
  XNOR2_X1 U5240 ( .A(n4253), .B(n4260), .ZN(n4254) );
  NAND2_X1 U5241 ( .A1(n4254), .A2(n6565), .ZN(n4255) );
  NAND2_X1 U5242 ( .A1(n4256), .A2(n4255), .ZN(n4257) );
  INV_X1 U5243 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4635) );
  XNOR2_X1 U5244 ( .A(n4257), .B(n4635), .ZN(n4630) );
  NAND2_X1 U5245 ( .A1(n4627), .A2(n4630), .ZN(n4628) );
  NAND2_X1 U5246 ( .A1(n4257), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4258)
         );
  NAND2_X1 U5247 ( .A1(n4628), .A2(n4258), .ZN(n6116) );
  NAND3_X1 U5248 ( .A1(n4283), .A2(n4259), .A3(n4269), .ZN(n4266) );
  NAND2_X1 U5249 ( .A1(n4261), .A2(n4260), .ZN(n4262) );
  OR2_X1 U5250 ( .A1(n4263), .A2(n4262), .ZN(n4271) );
  XNOR2_X1 U5251 ( .A(n4271), .B(n4272), .ZN(n4264) );
  NAND2_X1 U5252 ( .A1(n4264), .A2(n6565), .ZN(n4265) );
  NAND2_X1 U5253 ( .A1(n4266), .A2(n4265), .ZN(n4267) );
  XNOR2_X1 U5254 ( .A(n4267), .B(n6752), .ZN(n6115) );
  NAND2_X1 U5255 ( .A1(n6116), .A2(n6115), .ZN(n6114) );
  NAND2_X1 U5256 ( .A1(n4267), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4268)
         );
  NAND2_X1 U5257 ( .A1(n6114), .A2(n4268), .ZN(n6108) );
  NAND2_X1 U5258 ( .A1(n4270), .A2(n4269), .ZN(n4277) );
  INV_X1 U5259 ( .A(n4271), .ZN(n4273) );
  NAND2_X1 U5260 ( .A1(n4273), .A2(n4272), .ZN(n4285) );
  XNOR2_X1 U5261 ( .A(n4285), .B(n4274), .ZN(n4275) );
  NAND2_X1 U5262 ( .A1(n4275), .A2(n6565), .ZN(n4276) );
  NAND2_X1 U5263 ( .A1(n4277), .A2(n4276), .ZN(n4278) );
  INV_X1 U5264 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6174) );
  XNOR2_X1 U5265 ( .A(n4278), .B(n6174), .ZN(n6107) );
  NAND2_X1 U5266 ( .A1(n4278), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4279)
         );
  NAND2_X1 U5267 ( .A1(n6106), .A2(n4279), .ZN(n6100) );
  NAND2_X4 U5268 ( .A1(n4283), .A2(n4282), .ZN(n5604) );
  OR3_X1 U5269 ( .A1(n4285), .A2(n4284), .A3(n4345), .ZN(n4286) );
  NAND2_X1 U5270 ( .A1(n5604), .A2(n4286), .ZN(n4287) );
  XNOR2_X1 U5271 ( .A(n4287), .B(n6816), .ZN(n6099) );
  NAND2_X1 U5272 ( .A1(n6100), .A2(n6099), .ZN(n6098) );
  NAND2_X1 U5273 ( .A1(n4287), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4288)
         );
  INV_X1 U5274 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n6171) );
  NAND2_X1 U5275 ( .A1(n5604), .A2(n6171), .ZN(n6090) );
  NAND2_X1 U5276 ( .A1(n6093), .A2(n6090), .ZN(n4289) );
  NAND2_X1 U5277 ( .A1(n5592), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n6091)
         );
  INV_X1 U5278 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n4290) );
  NAND2_X1 U5279 ( .A1(n5604), .A2(n4290), .ZN(n5204) );
  AND2_X1 U5280 ( .A1(n5604), .A2(n6163), .ZN(n4293) );
  OR2_X1 U5281 ( .A1(n5604), .A2(n4290), .ZN(n6082) );
  OAI21_X1 U5282 ( .B1(n6163), .B2(n5604), .A(n6082), .ZN(n4291) );
  INV_X1 U5283 ( .A(n4291), .ZN(n4292) );
  INV_X1 U5284 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5242) );
  NOR2_X1 U5285 ( .A1(n5604), .A2(n5242), .ZN(n5231) );
  NAND2_X1 U5286 ( .A1(n5604), .A2(n5242), .ZN(n5229) );
  XNOR2_X1 U5287 ( .A(n5604), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5799)
         );
  NAND2_X1 U5288 ( .A1(n5798), .A2(n5799), .ZN(n4296) );
  INV_X1 U5289 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n4294) );
  NAND2_X1 U5290 ( .A1(n5604), .A2(n4294), .ZN(n4295) );
  NAND2_X1 U5291 ( .A1(n4296), .A2(n4295), .ZN(n5627) );
  INV_X1 U5292 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n4297) );
  AND2_X1 U5293 ( .A1(n5604), .A2(n4297), .ZN(n4299) );
  NAND2_X1 U5294 ( .A1(n5592), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n4298) );
  INV_X1 U5295 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5618) );
  NOR2_X1 U5296 ( .A1(n5604), .A2(n5618), .ZN(n4301) );
  NAND2_X1 U5297 ( .A1(n5604), .A2(n5618), .ZN(n4300) );
  OAI21_X1 U5298 ( .B1(n5286), .B2(n4301), .A(n4300), .ZN(n5603) );
  INV_X1 U5299 ( .A(n5603), .ZN(n4303) );
  NAND2_X1 U5300 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5594) );
  INV_X1 U5301 ( .A(n5594), .ZN(n5579) );
  NAND2_X1 U5302 ( .A1(n5579), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n4302) );
  INV_X1 U5303 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5625) );
  INV_X1 U5304 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5608) );
  INV_X1 U5305 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5811) );
  NAND3_X1 U5306 ( .A1(n5625), .A2(n5608), .A3(n5811), .ZN(n4304) );
  NAND2_X1 U5307 ( .A1(n5592), .A2(n4304), .ZN(n4305) );
  NAND2_X1 U5308 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5582) );
  AND2_X1 U5309 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5497) );
  AND2_X1 U5310 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4306) );
  NAND2_X1 U5311 ( .A1(n5497), .A2(n4306), .ZN(n4366) );
  OAI21_X1 U5312 ( .B1(n5582), .B2(n4366), .A(n5604), .ZN(n4307) );
  NAND2_X1 U5313 ( .A1(n5589), .A2(n4307), .ZN(n4310) );
  NOR2_X1 U5314 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5580) );
  NOR2_X1 U5315 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5258) );
  NOR2_X1 U5316 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5557) );
  NAND3_X1 U5317 ( .A1(n5580), .A2(n5258), .A3(n5557), .ZN(n4308) );
  NAND2_X1 U5318 ( .A1(n5592), .A2(n4308), .ZN(n4309) );
  INV_X1 U5319 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5807) );
  XNOR2_X1 U5320 ( .A(n5604), .B(n5807), .ZN(n5771) );
  NAND2_X1 U5321 ( .A1(n5604), .A2(n5807), .ZN(n4311) );
  NOR2_X1 U5322 ( .A1(n5604), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n4429)
         );
  NAND2_X1 U5323 ( .A1(n4312), .A2(n4429), .ZN(n5488) );
  INV_X1 U5324 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n6749) );
  INV_X1 U5325 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5482) );
  NAND2_X1 U5326 ( .A1(n6749), .A2(n5482), .ZN(n5534) );
  INV_X1 U5327 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5523) );
  INV_X1 U5328 ( .A(n4312), .ZN(n4427) );
  AND2_X1 U5329 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5532) );
  NAND2_X1 U5330 ( .A1(n5532), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5314) );
  AOI21_X1 U5331 ( .B1(n5342), .B2(n5523), .A(n5310), .ZN(n4313) );
  XNOR2_X1 U5332 ( .A(n4313), .B(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4400)
         );
  NOR2_X1 U5333 ( .A1(n5325), .A2(n4702), .ZN(n4361) );
  NAND2_X1 U5334 ( .A1(n5364), .A2(n4361), .ZN(n4321) );
  OR2_X1 U5335 ( .A1(n4314), .A2(n4593), .ZN(n4315) );
  MUX2_X1 U5336 ( .A(n4315), .B(n4345), .S(n3491), .Z(n4501) );
  AOI21_X1 U5337 ( .B1(n5325), .B2(n4593), .A(n4354), .ZN(n4317) );
  NAND2_X1 U5338 ( .A1(n4501), .A2(n4333), .ZN(n4318) );
  NAND2_X1 U5339 ( .A1(n4318), .A2(n5354), .ZN(n4457) );
  NAND2_X1 U5340 ( .A1(n3401), .A2(n6481), .ZN(n4319) );
  NOR2_X1 U5341 ( .A1(READY_N), .A2(n5355), .ZN(n4531) );
  NAND3_X1 U5342 ( .A1(n4319), .A2(n4531), .A3(n3483), .ZN(n4320) );
  NAND3_X1 U5343 ( .A1(n4321), .A2(n4457), .A3(n4320), .ZN(n4322) );
  NAND2_X1 U5344 ( .A1(n4322), .A2(n6463), .ZN(n4330) );
  INV_X1 U5345 ( .A(READY_N), .ZN(n4324) );
  NAND2_X1 U5346 ( .A1(n4325), .A2(n4324), .ZN(n4326) );
  INV_X1 U5347 ( .A(n5275), .ZN(n4351) );
  OAI211_X1 U5348 ( .C1(n4323), .C2(n4326), .A(n4555), .B(n4351), .ZN(n4327)
         );
  NAND2_X1 U5349 ( .A1(n4327), .A2(n3205), .ZN(n4328) );
  INV_X1 U5350 ( .A(n3524), .ZN(n4445) );
  NAND2_X1 U5351 ( .A1(n4333), .A2(n4445), .ZN(n4723) );
  INV_X1 U5352 ( .A(n4331), .ZN(n4332) );
  NAND2_X1 U5353 ( .A1(n4333), .A2(n4332), .ZN(n6444) );
  NAND2_X1 U5354 ( .A1(n4723), .A2(n6444), .ZN(n5353) );
  OAI211_X1 U5355 ( .C1(n4601), .C2(n4347), .A(n4719), .B(n4452), .ZN(n4335)
         );
  NOR2_X1 U5356 ( .A1(n5353), .A2(n4335), .ZN(n4336) );
  INV_X1 U5357 ( .A(n4337), .ZN(n4339) );
  INV_X1 U5358 ( .A(n4341), .ZN(n4342) );
  AOI211_X1 U5359 ( .C1(n5419), .C2(n5374), .A(n4342), .B(n4337), .ZN(n4343)
         );
  NOR2_X1 U5360 ( .A1(n4344), .A2(n4343), .ZN(n5652) );
  OR2_X1 U5361 ( .A1(n4323), .A2(n4345), .ZN(n6452) );
  OAI21_X1 U5362 ( .B1(n4347), .B2(n4346), .A(n6452), .ZN(n4348) );
  INV_X1 U5363 ( .A(n4348), .ZN(n4349) );
  INV_X2 U5364 ( .A(n6175), .ZN(n6210) );
  NAND2_X1 U5365 ( .A1(n6210), .A2(REIP_REG_30__SCAN_IN), .ZN(n4397) );
  INV_X1 U5366 ( .A(n4397), .ZN(n4368) );
  NAND2_X1 U5367 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5631) );
  NOR2_X1 U5368 ( .A1(n4294), .A2(n5631), .ZN(n5635) );
  NAND2_X1 U5369 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n5635), .ZN(n5617) );
  NAND2_X1 U5370 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5621) );
  NOR2_X1 U5371 ( .A1(n5617), .A2(n5621), .ZN(n4377) );
  INV_X1 U5372 ( .A(n4316), .ZN(n4350) );
  NAND2_X1 U5373 ( .A1(n4350), .A2(n5419), .ZN(n4358) );
  NAND2_X1 U5374 ( .A1(n4351), .A2(n3483), .ZN(n4352) );
  AND2_X1 U5375 ( .A1(n4353), .A2(n4352), .ZN(n4357) );
  NOR2_X1 U5376 ( .A1(n5081), .A2(n3483), .ZN(n4456) );
  OAI21_X1 U5377 ( .B1(n4456), .B2(n4470), .A(n4354), .ZN(n4355) );
  OAI21_X1 U5378 ( .B1(n4500), .B2(n4555), .A(n4733), .ZN(n4359) );
  INV_X1 U5379 ( .A(n4359), .ZN(n4360) );
  NOR2_X1 U5380 ( .A1(n4370), .A2(n4362), .ZN(n4369) );
  NAND2_X1 U5381 ( .A1(n4369), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n5630)
         );
  NOR2_X1 U5382 ( .A1(n4230), .A2(n6234), .ZN(n6213) );
  NAND3_X1 U5383 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .A3(n6213), .ZN(n4636) );
  NAND2_X1 U5384 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4363) );
  NOR2_X1 U5385 ( .A1(n4636), .A2(n4363), .ZN(n5208) );
  NAND2_X1 U5386 ( .A1(INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n5210) );
  NAND2_X1 U5387 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5211) );
  NOR2_X1 U5388 ( .A1(n5210), .A2(n5211), .ZN(n4364) );
  NAND2_X1 U5389 ( .A1(n5208), .A2(n4364), .ZN(n5238) );
  INV_X1 U5390 ( .A(n5357), .ZN(n4724) );
  AOI21_X1 U5391 ( .B1(INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .A(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .ZN(n6214) );
  NAND2_X1 U5392 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6199) );
  NOR2_X1 U5393 ( .A1(n6214), .A2(n6199), .ZN(n4631) );
  NAND2_X1 U5394 ( .A1(n6212), .A2(n4631), .ZN(n4634) );
  NOR2_X1 U5395 ( .A1(n4363), .A2(n4634), .ZN(n5207) );
  NAND2_X1 U5396 ( .A1(n4364), .A2(n5207), .ZN(n5629) );
  NAND2_X1 U5397 ( .A1(n4377), .A2(n6159), .ZN(n5812) );
  INV_X1 U5398 ( .A(n5582), .ZN(n4365) );
  NAND2_X1 U5399 ( .A1(n5579), .A2(n4365), .ZN(n4372) );
  INV_X1 U5400 ( .A(n5560), .ZN(n5568) );
  AND2_X1 U5401 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n4434) );
  NAND2_X1 U5402 ( .A1(n5802), .A2(n4434), .ZN(n5522) );
  NOR3_X1 U5403 ( .A1(n5522), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(n5314), 
        .ZN(n4367) );
  INV_X1 U5404 ( .A(n4369), .ZN(n4371) );
  NAND2_X1 U5405 ( .A1(n4371), .A2(n4382), .ZN(n6224) );
  INV_X1 U5406 ( .A(n5633), .ZN(n6223) );
  INV_X1 U5407 ( .A(n4434), .ZN(n4387) );
  INV_X1 U5408 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4487) );
  NAND2_X1 U5409 ( .A1(n4487), .A2(n6224), .ZN(n4486) );
  NAND2_X1 U5410 ( .A1(n4370), .A2(n6175), .ZN(n4488) );
  NAND2_X1 U5411 ( .A1(n4382), .A2(n6235), .ZN(n5237) );
  NAND2_X1 U5412 ( .A1(n4371), .A2(n5633), .ZN(n5239) );
  OAI21_X1 U5413 ( .B1(n5237), .B2(n5239), .A(n4372), .ZN(n4376) );
  INV_X1 U5414 ( .A(n5238), .ZN(n4373) );
  NAND2_X1 U5415 ( .A1(n4377), .A2(n4373), .ZN(n4374) );
  AND2_X1 U5416 ( .A1(n5239), .A2(n4374), .ZN(n5575) );
  INV_X1 U5417 ( .A(n5575), .ZN(n4375) );
  AND2_X1 U5418 ( .A1(n4376), .A2(n4375), .ZN(n4380) );
  INV_X1 U5419 ( .A(n4377), .ZN(n4378) );
  NOR2_X1 U5420 ( .A1(n4378), .A2(n5629), .ZN(n5574) );
  INV_X1 U5421 ( .A(n5237), .ZN(n5573) );
  OR2_X1 U5422 ( .A1(n5574), .A2(n5573), .ZN(n4379) );
  NAND2_X1 U5423 ( .A1(n4380), .A2(n4379), .ZN(n5570) );
  INV_X1 U5424 ( .A(n5497), .ZN(n5559) );
  AND2_X1 U5425 ( .A1(n4632), .A2(n5559), .ZN(n4381) );
  NOR2_X1 U5426 ( .A1(n5570), .A2(n4381), .ZN(n5549) );
  NAND2_X1 U5427 ( .A1(n5609), .A2(n4382), .ZN(n4384) );
  NAND2_X1 U5428 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4383) );
  NAND2_X1 U5429 ( .A1(n4384), .A2(n4383), .ZN(n4385) );
  INV_X1 U5430 ( .A(n5808), .ZN(n4386) );
  AOI21_X1 U5431 ( .B1(n4632), .B2(n4387), .A(n4386), .ZN(n5548) );
  OAI21_X1 U5432 ( .B1(n5532), .B2(n5289), .A(n5548), .ZN(n5528) );
  AOI21_X1 U5433 ( .B1(INSTADDRPOINTER_REG_30__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_29__SCAN_IN), .A(n5289), .ZN(n4388) );
  NOR2_X1 U5434 ( .A1(n5528), .A2(n4388), .ZN(n5312) );
  INV_X1 U5435 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5313) );
  NAND3_X1 U5436 ( .A1(n4391), .A2(n4390), .A3(n4389), .ZN(U2988) );
  NOR2_X2 U5437 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .ZN(
        n6313) );
  NAND2_X1 U5438 ( .A1(n6275), .A2(n4392), .ZN(n6570) );
  NAND2_X1 U5439 ( .A1(n6570), .A2(n6567), .ZN(n4393) );
  NAND2_X1 U5440 ( .A1(n6567), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4395) );
  NAND2_X1 U5441 ( .A1(n6564), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4394) );
  AND2_X1 U5442 ( .A1(n4395), .A2(n4394), .ZN(n4525) );
  INV_X1 U5443 ( .A(n4525), .ZN(n4396) );
  NAND2_X1 U5444 ( .A1(n5651), .A2(n6134), .ZN(n4398) );
  OAI211_X1 U5445 ( .C1(n5791), .C2(n6707), .A(n4398), .B(n4397), .ZN(n4399)
         );
  AOI21_X1 U5446 ( .B1(n4400), .B2(n6152), .A(n4399), .ZN(n4405) );
  XOR2_X2 U5447 ( .A(n4401), .B(n4407), .Z(n5741) );
  NAND3_X1 U5448 ( .A1(n6567), .A2(STATEBS16_REG_SCAN_IN), .A3(
        STATE2_REG_1__SCAN_IN), .ZN(n6472) );
  INV_X1 U5449 ( .A(n6472), .ZN(n4402) );
  INV_X1 U5450 ( .A(n6138), .ZN(n4403) );
  NAND2_X1 U5451 ( .A1(n4405), .A2(n4404), .ZN(U2956) );
  AND2_X1 U5452 ( .A1(n5375), .A2(n4406), .ZN(n4408) );
  INV_X1 U5453 ( .A(n4409), .ZN(n4410) );
  NAND2_X1 U5454 ( .A1(n5374), .A2(n4410), .ZN(n4411) );
  NAND2_X1 U5455 ( .A1(n4412), .A2(n4411), .ZN(n5526) );
  OAI22_X1 U5456 ( .A1(n5341), .A2(n5967), .B1(n5526), .B2(n5969), .ZN(n4426)
         );
  INV_X1 U5457 ( .A(n4413), .ZN(n4414) );
  OAI22_X1 U5458 ( .A1(n6884), .A2(n5970), .B1(n5346), .B2(n5990), .ZN(n4423)
         );
  NAND3_X1 U5459 ( .A1(n4555), .A2(n4416), .A3(n4415), .ZN(n4417) );
  NAND2_X1 U5460 ( .A1(n4418), .A2(n4417), .ZN(n4420) );
  INV_X1 U5461 ( .A(n5080), .ZN(n4419) );
  OAI21_X1 U5462 ( .B1(n5659), .B2(n6530), .A(n4421), .ZN(n4422) );
  OR2_X1 U5463 ( .A1(n4426), .A2(n4425), .ZN(U2798) );
  INV_X1 U5464 ( .A(n4428), .ZN(n4432) );
  NOR2_X1 U5465 ( .A1(n4429), .A2(n4428), .ZN(n4430) );
  NAND2_X1 U5466 ( .A1(n3212), .A2(n4430), .ZN(n4431) );
  OAI211_X1 U5467 ( .C1(n3212), .C2(n4432), .A(n5488), .B(n4431), .ZN(n5765)
         );
  AND2_X1 U5468 ( .A1(n5765), .A2(n6231), .ZN(n4441) );
  INV_X1 U5469 ( .A(n5802), .ZN(n4433) );
  AOI211_X1 U5470 ( .C1(n4435), .C2(n5807), .A(n4434), .B(n4433), .ZN(n4440)
         );
  NOR2_X1 U5471 ( .A1(n5808), .A2(n4435), .ZN(n4439) );
  OR2_X1 U5472 ( .A1(n5390), .A2(n4436), .ZN(n4437) );
  NAND2_X1 U5473 ( .A1(n5382), .A2(n4437), .ZN(n5673) );
  OAI22_X1 U5474 ( .A1(n5673), .A2(n6177), .B1(n6175), .B2(n6526), .ZN(n4438)
         );
  INV_X1 U5475 ( .A(n4442), .ZN(n4443) );
  INV_X1 U5476 ( .A(MEMORYFETCH_REG_SCAN_IN), .ZN(n6574) );
  NAND2_X1 U5477 ( .A1(n6313), .A2(n6736), .ZN(n5827) );
  OAI211_X1 U5478 ( .C1(n4443), .C2(n6574), .A(n4448), .B(n5827), .ZN(U2788)
         );
  INV_X1 U5479 ( .A(n5827), .ZN(n4444) );
  NOR2_X1 U5480 ( .A1(n4444), .A2(READREQUEST_REG_SCAN_IN), .ZN(n4447) );
  OAI21_X1 U5481 ( .B1(n4445), .B2(n4497), .A(n6569), .ZN(n4446) );
  OAI21_X1 U5482 ( .B1(n4447), .B2(n6569), .A(n4446), .ZN(U3474) );
  INV_X1 U5483 ( .A(EAX_REG_15__SCAN_IN), .ZN(n4451) );
  INV_X1 U5484 ( .A(n4448), .ZN(n4449) );
  OAI21_X1 U5485 ( .B1(n4324), .B2(n6565), .A(n4449), .ZN(n6074) );
  INV_X1 U5486 ( .A(LWORD_REG_15__SCAN_IN), .ZN(n6814) );
  INV_X1 U5487 ( .A(DATAI_15_), .ZN(n4450) );
  OAI222_X1 U5488 ( .A1(n6045), .A2(n4451), .B1(n6044), .B2(n6814), .C1(n6081), 
        .C2(n4450), .ZN(U2954) );
  NAND2_X1 U5489 ( .A1(n4731), .A2(n4323), .ZN(n4454) );
  NAND2_X1 U5490 ( .A1(n4452), .A2(n6481), .ZN(n4453) );
  NAND3_X1 U5491 ( .A1(n4454), .A2(n4324), .A3(n4453), .ZN(n4455) );
  OR2_X1 U5492 ( .A1(n5364), .A2(n4455), .ZN(n4462) );
  OR2_X1 U5493 ( .A1(n5364), .A2(n4723), .ZN(n4461) );
  NAND2_X1 U5494 ( .A1(n5357), .A2(n5364), .ZN(n4460) );
  INV_X1 U5495 ( .A(n4719), .ZN(n4467) );
  AOI21_X1 U5496 ( .B1(n4467), .B2(n4531), .A(n4456), .ZN(n4458) );
  AND2_X1 U5497 ( .A1(n4458), .A2(n4457), .ZN(n4459) );
  NAND4_X1 U5498 ( .A1(n4462), .A2(n4461), .A3(n4460), .A4(n4459), .ZN(n4744)
         );
  INV_X1 U5499 ( .A(n4744), .ZN(n6433) );
  NOR2_X1 U5500 ( .A1(n6736), .A2(n4463), .ZN(n4760) );
  NAND2_X1 U5501 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4760), .ZN(n6545) );
  INV_X1 U5502 ( .A(FLUSH_REG_SCAN_IN), .ZN(n5832) );
  OAI22_X1 U5503 ( .A1(n6433), .A2(n6461), .B1(n6545), .B2(n5832), .ZN(n4466)
         );
  AOI21_X1 U5504 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n6567), .A(n4466), .ZN(
        n6553) );
  INV_X1 U5505 ( .A(n6553), .ZN(n4515) );
  INV_X1 U5506 ( .A(n6268), .ZN(n4691) );
  NOR2_X1 U5507 ( .A1(n4464), .A2(n4691), .ZN(n4465) );
  XNOR2_X1 U5508 ( .A(n4465), .B(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n5102)
         );
  INV_X1 U5509 ( .A(n5102), .ZN(n4468) );
  INV_X1 U5510 ( .A(n4512), .ZN(n6550) );
  NAND4_X1 U5511 ( .A1(n4468), .A2(n6550), .A3(n4467), .A4(n4466), .ZN(n4469)
         );
  OAI21_X1 U5512 ( .B1(n4515), .B2(n3436), .A(n4469), .ZN(U3455) );
  NOR2_X1 U5513 ( .A1(n4470), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4471)
         );
  OR2_X1 U5514 ( .A1(n4472), .A2(n4471), .ZN(n5108) );
  NAND3_X1 U5515 ( .A1(n5357), .A2(n5364), .A3(n6463), .ZN(n4478) );
  NAND4_X1 U5516 ( .A1(n3622), .A2(n3701), .A3(n4473), .A4(n6736), .ZN(n4532)
         );
  INV_X1 U5517 ( .A(n4532), .ZN(n4476) );
  NOR2_X1 U5518 ( .A1(n4474), .A2(n3196), .ZN(n4475) );
  NAND2_X1 U5519 ( .A1(n4476), .A2(n4475), .ZN(n4477) );
  INV_X1 U5520 ( .A(n3516), .ZN(n5468) );
  INV_X1 U5521 ( .A(n4479), .ZN(n4482) );
  OAI21_X1 U5522 ( .B1(n4482), .B2(n4481), .A(n4480), .ZN(n5114) );
  OAI222_X1 U5523 ( .A1(n5108), .A2(n5466), .B1(n5453), .B2(n5109), .C1(n3195), 
        .C2(n5114), .ZN(U2859) );
  XNOR2_X1 U5524 ( .A(n4483), .B(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4530)
         );
  INV_X1 U5525 ( .A(REIP_REG_0__SCAN_IN), .ZN(n4484) );
  NOR2_X1 U5526 ( .A1(n6175), .A2(n4484), .ZN(n4527) );
  INV_X1 U5527 ( .A(n4527), .ZN(n4485) );
  OAI211_X1 U5528 ( .C1(n6177), .C2(n5108), .A(n4486), .B(n4485), .ZN(n4490)
         );
  AOI21_X1 U5529 ( .B1(n5633), .B2(n4488), .A(n4487), .ZN(n4489) );
  NOR2_X1 U5530 ( .A1(n4490), .A2(n4489), .ZN(n4491) );
  OAI21_X1 U5531 ( .B1(n4530), .B2(n5815), .A(n4491), .ZN(U3018) );
  OR2_X1 U5532 ( .A1(n4493), .A2(n4492), .ZN(n4494) );
  NAND2_X1 U5533 ( .A1(n4495), .A2(n4494), .ZN(n5098) );
  OAI21_X1 U5534 ( .B1(n5093), .B2(n4497), .A(n4496), .ZN(n6226) );
  AOI22_X1 U5535 ( .A1(n5445), .A2(n6226), .B1(n5462), .B2(EBX_REG_1__SCAN_IN), 
        .ZN(n4498) );
  OAI21_X1 U5536 ( .B1(n5098), .B2(n3195), .A(n4498), .ZN(U2858) );
  INV_X1 U5537 ( .A(n5644), .ZN(n4767) );
  AND4_X1 U5538 ( .A1(n4719), .A2(n4323), .A3(n4533), .A4(n4500), .ZN(n4502)
         );
  AND3_X1 U5539 ( .A1(n4503), .A2(n4502), .A3(n4501), .ZN(n5326) );
  INV_X1 U5540 ( .A(n5326), .ZN(n4509) );
  INV_X1 U5541 ( .A(n5325), .ZN(n4506) );
  OAI21_X1 U5542 ( .B1(n4504), .B2(n4505), .A(n4506), .ZN(n4507) );
  OAI21_X1 U5543 ( .B1(n4731), .B2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(n4507), 
        .ZN(n4508) );
  AOI21_X1 U5544 ( .B1(n4767), .B2(n4509), .A(n4508), .ZN(n6432) );
  AOI22_X1 U5545 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n3214), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n6234), .ZN(n5335) );
  NAND2_X1 U5546 ( .A1(STATE2_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n5334) );
  INV_X1 U5547 ( .A(n5334), .ZN(n4510) );
  AOI22_X1 U5548 ( .A1(n5335), .A2(n4510), .B1(n4505), .B2(n6548), .ZN(n4511)
         );
  OAI21_X1 U5549 ( .B1(n6432), .B2(n4512), .A(n4511), .ZN(n4513) );
  AOI22_X1 U5550 ( .A1(n4515), .A2(n4513), .B1(n4504), .B2(n6548), .ZN(n4514)
         );
  OAI21_X1 U5551 ( .B1(n3394), .B2(n4515), .A(n4514), .ZN(U3460) );
  INV_X1 U5552 ( .A(EAX_REG_10__SCAN_IN), .ZN(n6023) );
  NAND2_X1 U5553 ( .A1(n6051), .A2(LWORD_REG_10__SCAN_IN), .ZN(n4516) );
  NAND2_X1 U5554 ( .A1(n6075), .A2(DATAI_10_), .ZN(n4520) );
  OAI211_X1 U5555 ( .C1(n6023), .C2(n6045), .A(n4516), .B(n4520), .ZN(U2949)
         );
  NAND2_X1 U5556 ( .A1(n6051), .A2(UWORD_REG_8__SCAN_IN), .ZN(n4517) );
  NAND2_X1 U5557 ( .A1(n6075), .A2(DATAI_8_), .ZN(n4518) );
  OAI211_X1 U5558 ( .C1(n4097), .C2(n6045), .A(n4517), .B(n4518), .ZN(U2932)
         );
  INV_X1 U5559 ( .A(EAX_REG_8__SCAN_IN), .ZN(n6026) );
  NAND2_X1 U5560 ( .A1(n6051), .A2(LWORD_REG_8__SCAN_IN), .ZN(n4519) );
  OAI211_X1 U5561 ( .C1(n6026), .C2(n6045), .A(n4519), .B(n4518), .ZN(U2947)
         );
  INV_X1 U5562 ( .A(EAX_REG_26__SCAN_IN), .ZN(n4566) );
  NAND2_X1 U5563 ( .A1(n6051), .A2(UWORD_REG_10__SCAN_IN), .ZN(n4521) );
  OAI211_X1 U5564 ( .C1(n4566), .C2(n6045), .A(n4521), .B(n4520), .ZN(U2934)
         );
  INV_X1 U5565 ( .A(EAX_REG_25__SCAN_IN), .ZN(n4564) );
  AOI22_X1 U5566 ( .A1(n6051), .A2(UWORD_REG_9__SCAN_IN), .B1(n6075), .B2(
        DATAI_9_), .ZN(n4522) );
  OAI21_X1 U5567 ( .B1(n4564), .B2(n6045), .A(n4522), .ZN(U2933) );
  INV_X1 U5568 ( .A(EAX_REG_27__SCAN_IN), .ZN(n4568) );
  AOI22_X1 U5569 ( .A1(n6051), .A2(UWORD_REG_11__SCAN_IN), .B1(n6075), .B2(
        DATAI_11_), .ZN(n4523) );
  OAI21_X1 U5570 ( .B1(n4568), .B2(n6045), .A(n4523), .ZN(U2935) );
  INV_X1 U5571 ( .A(EAX_REG_28__SCAN_IN), .ZN(n4570) );
  AOI22_X1 U5572 ( .A1(n6051), .A2(UWORD_REG_12__SCAN_IN), .B1(n6075), .B2(
        DATAI_12_), .ZN(n4524) );
  OAI21_X1 U5573 ( .B1(n4570), .B2(n6045), .A(n4524), .ZN(U2936) );
  NAND2_X1 U5574 ( .A1(n4525), .A2(n5791), .ZN(n4528) );
  NOR2_X1 U5575 ( .A1(n5114), .A2(n6138), .ZN(n4526) );
  AOI211_X1 U5576 ( .C1(PHYADDRPOINTER_REG_0__SCAN_IN), .C2(n4528), .A(n4527), 
        .B(n4526), .ZN(n4529) );
  OAI21_X1 U5577 ( .B1(n4530), .B2(n5831), .A(n4529), .ZN(U2986) );
  NAND2_X1 U5578 ( .A1(n6463), .A2(n4531), .ZN(n4534) );
  OAI22_X1 U5579 ( .A1(n4719), .A2(n4534), .B1(n4533), .B2(n4532), .ZN(n4535)
         );
  INV_X1 U5580 ( .A(n4535), .ZN(n4536) );
  NAND2_X1 U5581 ( .A1(n4537), .A2(n3516), .ZN(n4538) );
  INV_X1 U5582 ( .A(n4538), .ZN(n4539) );
  INV_X1 U5583 ( .A(DATAI_1_), .ZN(n6890) );
  OAI222_X1 U5584 ( .A1(n5098), .A2(n6970), .B1(n6969), .B2(n6890), .C1(n6967), 
        .C2(n3629), .ZN(U2890) );
  INV_X1 U5585 ( .A(DATAI_0_), .ZN(n6861) );
  INV_X1 U5586 ( .A(EAX_REG_0__SCAN_IN), .ZN(n6043) );
  OAI222_X1 U5587 ( .A1(n5114), .A2(n6970), .B1(n6969), .B2(n6861), .C1(n6967), 
        .C2(n6043), .ZN(U2891) );
  INV_X1 U5588 ( .A(n4540), .ZN(n4541) );
  OAI21_X1 U5589 ( .B1(n4543), .B2(n4542), .A(n4541), .ZN(n6148) );
  INV_X1 U5590 ( .A(n4575), .ZN(n4545) );
  XNOR2_X1 U5591 ( .A(n4544), .B(n4545), .ZN(n6209) );
  INV_X1 U5592 ( .A(EBX_REG_2__SCAN_IN), .ZN(n4546) );
  OAI222_X1 U5593 ( .A1(n6148), .A2(n3195), .B1(n5466), .B2(n6209), .C1(n5453), 
        .C2(n4546), .ZN(U2857) );
  INV_X1 U5594 ( .A(DATAI_2_), .ZN(n6060) );
  OAI222_X1 U5595 ( .A1(n6148), .A2(n6970), .B1(n6969), .B2(n6060), .C1(n6967), 
        .C2(n3649), .ZN(U2889) );
  XNOR2_X1 U5596 ( .A(n4548), .B(n4547), .ZN(n6222) );
  INV_X1 U5597 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6555) );
  NOR2_X1 U5598 ( .A1(n6175), .A2(n6555), .ZN(n6225) );
  OAI22_X1 U5599 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n6157), .B1(n6138), 
        .B2(n5098), .ZN(n4549) );
  AOI211_X1 U5600 ( .C1(n6147), .C2(PHYADDRPOINTER_REG_1__SCAN_IN), .A(n6225), 
        .B(n4549), .ZN(n4550) );
  OAI21_X1 U5601 ( .B1(n6222), .B2(n5831), .A(n4550), .ZN(U2985) );
  INV_X1 U5602 ( .A(EAX_REG_18__SCAN_IN), .ZN(n6841) );
  NAND2_X1 U5603 ( .A1(n6045), .A2(n4552), .ZN(n4554) );
  NAND2_X1 U5604 ( .A1(n6029), .A2(n4555), .ZN(n6009) );
  NAND2_X1 U5605 ( .A1(n6567), .A2(n4760), .ZN(n6033) );
  INV_X2 U5606 ( .A(n6033), .ZN(n6040) );
  AOI22_X1 U5607 ( .A1(UWORD_REG_2__SCAN_IN), .A2(n6040), .B1(n6039), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n4556) );
  OAI21_X1 U5608 ( .B1(n6841), .B2(n6009), .A(n4556), .ZN(U2905) );
  AOI22_X1 U5609 ( .A1(UWORD_REG_4__SCAN_IN), .A2(n6040), .B1(n6039), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n4557) );
  OAI21_X1 U5610 ( .B1(n3940), .B2(n6009), .A(n4557), .ZN(U2903) );
  INV_X1 U5611 ( .A(EAX_REG_16__SCAN_IN), .ZN(n6764) );
  AOI22_X1 U5612 ( .A1(UWORD_REG_0__SCAN_IN), .A2(n6040), .B1(n6039), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n4558) );
  OAI21_X1 U5613 ( .B1(n6764), .B2(n6009), .A(n4558), .ZN(U2907) );
  AOI22_X1 U5614 ( .A1(n6040), .A2(UWORD_REG_14__SCAN_IN), .B1(n6039), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n4559) );
  OAI21_X1 U5615 ( .B1(n4170), .B2(n6009), .A(n4559), .ZN(U2893) );
  AOI22_X1 U5616 ( .A1(n6040), .A2(UWORD_REG_7__SCAN_IN), .B1(n6039), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n4560) );
  OAI21_X1 U5617 ( .B1(n4561), .B2(n6009), .A(n4560), .ZN(U2900) );
  AOI22_X1 U5618 ( .A1(n6040), .A2(UWORD_REG_8__SCAN_IN), .B1(n6039), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n4562) );
  OAI21_X1 U5619 ( .B1(n4097), .B2(n6009), .A(n4562), .ZN(U2899) );
  AOI22_X1 U5620 ( .A1(n6040), .A2(UWORD_REG_9__SCAN_IN), .B1(n6039), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n4563) );
  OAI21_X1 U5621 ( .B1(n4564), .B2(n6009), .A(n4563), .ZN(U2898) );
  AOI22_X1 U5622 ( .A1(n6040), .A2(UWORD_REG_10__SCAN_IN), .B1(n6039), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n4565) );
  OAI21_X1 U5623 ( .B1(n4566), .B2(n6009), .A(n4565), .ZN(U2897) );
  AOI22_X1 U5624 ( .A1(n6040), .A2(UWORD_REG_11__SCAN_IN), .B1(n6039), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n4567) );
  OAI21_X1 U5625 ( .B1(n4568), .B2(n6009), .A(n4567), .ZN(U2896) );
  AOI22_X1 U5626 ( .A1(n6040), .A2(UWORD_REG_12__SCAN_IN), .B1(n6039), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n4569) );
  OAI21_X1 U5627 ( .B1(n4570), .B2(n6009), .A(n4569), .ZN(U2895) );
  INV_X1 U5628 ( .A(EAX_REG_29__SCAN_IN), .ZN(n4572) );
  AOI22_X1 U5629 ( .A1(n6040), .A2(UWORD_REG_13__SCAN_IN), .B1(n6039), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n4571) );
  OAI21_X1 U5630 ( .B1(n4572), .B2(n6009), .A(n4571), .ZN(U2894) );
  XOR2_X1 U5631 ( .A(n4540), .B(n4573), .Z(n6143) );
  INV_X1 U5632 ( .A(n6143), .ZN(n6971) );
  AOI21_X1 U5633 ( .B1(n3294), .B2(n4575), .A(n4574), .ZN(n4576) );
  INV_X1 U5634 ( .A(n4582), .ZN(n4639) );
  NOR2_X1 U5635 ( .A1(n4576), .A2(n4639), .ZN(n6203) );
  AOI22_X1 U5636 ( .A1(n5445), .A2(n6203), .B1(n5462), .B2(EBX_REG_3__SCAN_IN), 
        .ZN(n4577) );
  OAI21_X1 U5637 ( .B1(n6971), .B2(n3195), .A(n4577), .ZN(U2856) );
  NAND2_X1 U5638 ( .A1(n4580), .A2(n4579), .ZN(n4581) );
  NAND2_X1 U5639 ( .A1(n4578), .A2(n4581), .ZN(n6137) );
  XNOR2_X1 U5640 ( .A(n4582), .B(n4638), .ZN(n6196) );
  AOI22_X1 U5641 ( .A1(n5445), .A2(n6196), .B1(n5462), .B2(EBX_REG_4__SCAN_IN), 
        .ZN(n4583) );
  OAI21_X1 U5642 ( .B1(n6137), .B2(n3195), .A(n4583), .ZN(U2855) );
  INV_X1 U5643 ( .A(DATAI_4_), .ZN(n6063) );
  INV_X1 U5644 ( .A(EAX_REG_4__SCAN_IN), .ZN(n6034) );
  OAI222_X1 U5645 ( .A1(n6137), .A2(n6970), .B1(n6969), .B2(n6063), .C1(n6967), 
        .C2(n6034), .ZN(U2887) );
  OR3_X1 U5646 ( .A1(n4829), .A2(n4765), .A3(n4689), .ZN(n4597) );
  INV_X1 U5647 ( .A(n4597), .ZN(n4587) );
  AND2_X1 U5648 ( .A1(n6313), .A2(n6564), .ZN(n4980) );
  INV_X1 U5649 ( .A(n4980), .ZN(n6316) );
  OAI21_X1 U5650 ( .B1(n4587), .B2(n6138), .A(n6316), .ZN(n4590) );
  AND2_X1 U5651 ( .A1(n6311), .A2(n4860), .ZN(n4769) );
  INV_X1 U5652 ( .A(n4798), .ZN(n4705) );
  AOI21_X1 U5653 ( .B1(n4769), .B2(n4842), .A(n4705), .ZN(n4594) );
  NAND2_X1 U5654 ( .A1(n4590), .A2(n4594), .ZN(n4591) );
  OAI211_X1 U5655 ( .C1(n6313), .C2(n4595), .A(n4591), .B(n6272), .ZN(n4800)
         );
  INV_X1 U5656 ( .A(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4600) );
  NOR2_X2 U5657 ( .A1(n4703), .A2(n4593), .ZN(n6380) );
  INV_X1 U5658 ( .A(n4594), .ZN(n4596) );
  AOI22_X1 U5659 ( .A1(n4596), .A2(n6313), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4595), .ZN(n4803) );
  INV_X1 U5660 ( .A(n4803), .ZN(n4704) );
  AOI22_X1 U5661 ( .A1(n6380), .A2(n4705), .B1(n6383), .B2(n4704), .ZN(n4599)
         );
  INV_X1 U5662 ( .A(n6138), .ZN(n6124) );
  NAND2_X1 U5663 ( .A1(n6124), .A2(DATAI_24_), .ZN(n4900) );
  INV_X1 U5664 ( .A(n4900), .ZN(n6381) );
  NOR2_X2 U5665 ( .A1(n4597), .A2(n6276), .ZN(n4933) );
  NOR2_X2 U5666 ( .A1(n4597), .A2(n4866), .ZN(n5067) );
  NAND2_X1 U5667 ( .A1(n4403), .A2(DATAI_16_), .ZN(n6324) );
  INV_X1 U5668 ( .A(n6324), .ZN(n6382) );
  AOI22_X1 U5669 ( .A1(n6381), .A2(n4933), .B1(n5067), .B2(n6382), .ZN(n4598)
         );
  OAI211_X1 U5670 ( .C1(n4709), .C2(n4600), .A(n4599), .B(n4598), .ZN(U3140)
         );
  INV_X1 U5671 ( .A(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4604) );
  NOR2_X2 U5672 ( .A1(n4703), .A2(n4601), .ZN(n6358) );
  AOI22_X1 U5673 ( .A1(n6358), .A2(n4705), .B1(n6360), .B2(n4704), .ZN(n4603)
         );
  NAND2_X1 U5674 ( .A1(n6124), .A2(DATAI_28_), .ZN(n6363) );
  INV_X1 U5675 ( .A(n6363), .ZN(n6336) );
  NAND2_X1 U5676 ( .A1(n4403), .A2(DATAI_20_), .ZN(n6339) );
  INV_X1 U5677 ( .A(n6339), .ZN(n6359) );
  AOI22_X1 U5678 ( .A1(n6336), .A2(n4933), .B1(n5067), .B2(n6359), .ZN(n4602)
         );
  OAI211_X1 U5679 ( .C1(n4709), .C2(n4604), .A(n4603), .B(n4602), .ZN(U3144)
         );
  INV_X1 U5680 ( .A(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4608) );
  NOR2_X2 U5681 ( .A1(n4703), .A2(n4605), .ZN(n6407) );
  INV_X1 U5682 ( .A(DATAI_3_), .ZN(n6968) );
  AOI22_X1 U5683 ( .A1(n6407), .A2(n4705), .B1(n6408), .B2(n4704), .ZN(n4607)
         );
  NAND2_X1 U5684 ( .A1(n4403), .A2(DATAI_27_), .ZN(n6411) );
  INV_X1 U5685 ( .A(n6411), .ZN(n6332) );
  NAND2_X1 U5686 ( .A1(n6124), .A2(DATAI_19_), .ZN(n6335) );
  INV_X1 U5687 ( .A(n6335), .ZN(n6406) );
  AOI22_X1 U5688 ( .A1(n6332), .A2(n4933), .B1(n5067), .B2(n6406), .ZN(n4606)
         );
  OAI211_X1 U5689 ( .C1(n4709), .C2(n4608), .A(n4607), .B(n4606), .ZN(U3143)
         );
  INV_X1 U5690 ( .A(DATAI_7_), .ZN(n6069) );
  INV_X1 U5691 ( .A(n6373), .ZN(n5163) );
  NAND2_X1 U5692 ( .A1(n4403), .A2(DATAI_31_), .ZN(n6378) );
  INV_X1 U5693 ( .A(n6378), .ZN(n6351) );
  NAND2_X1 U5694 ( .A1(n4403), .A2(DATAI_23_), .ZN(n6355) );
  INV_X1 U5695 ( .A(n5067), .ZN(n5003) );
  OAI22_X1 U5696 ( .A1(n5010), .A2(n4798), .B1(n6355), .B2(n5003), .ZN(n4609)
         );
  AOI21_X1 U5697 ( .B1(n6351), .B2(n4933), .A(n4609), .ZN(n4611) );
  NAND2_X1 U5698 ( .A1(n4800), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4610)
         );
  OAI211_X1 U5699 ( .C1(n4803), .C2(n5163), .A(n4611), .B(n4610), .ZN(U3147)
         );
  AND2_X1 U5700 ( .A1(n5642), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5645) );
  AND2_X1 U5701 ( .A1(n5645), .A2(n4829), .ZN(n4947) );
  INV_X1 U5702 ( .A(n4947), .ZN(n4828) );
  INV_X1 U5703 ( .A(n4857), .ZN(n4756) );
  OAI21_X1 U5704 ( .B1(n4828), .B2(n4756), .A(n6313), .ZN(n4615) );
  AND2_X1 U5705 ( .A1(n3227), .A2(n6311), .ZN(n5150) );
  NOR2_X1 U5706 ( .A1(n6441), .A2(n4950), .ZN(n6420) );
  AOI21_X1 U5707 ( .B1(n5150), .B2(n4860), .A(n6420), .ZN(n4612) );
  NAND2_X1 U5708 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n4953), .ZN(n5149) );
  OAI22_X1 U5709 ( .A1(n4615), .A2(n4612), .B1(n5149), .B2(n4463), .ZN(n6422)
         );
  INV_X1 U5710 ( .A(n6422), .ZN(n4626) );
  INV_X1 U5711 ( .A(n4612), .ZN(n4614) );
  AOI21_X1 U5712 ( .B1(n6275), .B2(n5149), .A(n4958), .ZN(n4613) );
  OAI21_X1 U5713 ( .B1(n4615), .B2(n4614), .A(n4613), .ZN(n6424) );
  NAND2_X1 U5714 ( .A1(n4829), .A2(n5642), .ZN(n4646) );
  INV_X1 U5715 ( .A(n4646), .ZN(n4616) );
  NAND3_X1 U5716 ( .A1(n4616), .A2(n6276), .A3(n4857), .ZN(n5062) );
  AOI22_X1 U5717 ( .A1(n6358), .A2(n6420), .B1(n6419), .B2(n6359), .ZN(n4617)
         );
  OAI21_X1 U5718 ( .B1(n6363), .B2(n6427), .A(n4617), .ZN(n4618) );
  AOI21_X1 U5719 ( .B1(INSTQUEUE_REG_11__4__SCAN_IN), .B2(n6424), .A(n4618), 
        .ZN(n4619) );
  OAI21_X1 U5720 ( .B1(n4626), .B2(n5179), .A(n4619), .ZN(U3112) );
  INV_X1 U5721 ( .A(n6355), .ZN(n6371) );
  AOI22_X1 U5722 ( .A1(n6369), .A2(n6420), .B1(n6419), .B2(n6371), .ZN(n4620)
         );
  OAI21_X1 U5723 ( .B1(n6378), .B2(n6427), .A(n4620), .ZN(n4621) );
  AOI21_X1 U5724 ( .B1(INSTQUEUE_REG_11__7__SCAN_IN), .B2(n6424), .A(n4621), 
        .ZN(n4622) );
  OAI21_X1 U5725 ( .B1(n4626), .B2(n5163), .A(n4622), .ZN(U3115) );
  INV_X1 U5726 ( .A(n6383), .ZN(n5167) );
  AOI22_X1 U5727 ( .A1(n6380), .A2(n6420), .B1(n6419), .B2(n6382), .ZN(n4623)
         );
  OAI21_X1 U5728 ( .B1(n4900), .B2(n6427), .A(n4623), .ZN(n4624) );
  AOI21_X1 U5729 ( .B1(INSTQUEUE_REG_11__0__SCAN_IN), .B2(n6424), .A(n4624), 
        .ZN(n4625) );
  OAI21_X1 U5730 ( .B1(n4626), .B2(n5167), .A(n4625), .ZN(U3108) );
  OAI21_X1 U5731 ( .B1(n4627), .B2(n4630), .A(n4629), .ZN(n6122) );
  INV_X1 U5732 ( .A(n5239), .ZN(n5578) );
  OAI22_X1 U5733 ( .A1(n5578), .A2(n6213), .B1(n6212), .B2(n6235), .ZN(n6216)
         );
  NAND2_X1 U5734 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n4631), .ZN(n5209)
         );
  AND2_X1 U5735 ( .A1(n4632), .A2(n5209), .ZN(n4633) );
  OR2_X1 U5736 ( .A1(n6216), .A2(n4633), .ZN(n6189) );
  OAI211_X1 U5737 ( .C1(n5609), .C2(n4636), .A(n4635), .B(n4634), .ZN(n4644)
         );
  AOI21_X1 U5738 ( .B1(n4639), .B2(n4638), .A(n4637), .ZN(n4641) );
  CLKBUF_X1 U5739 ( .A(n4640), .Z(n5130) );
  OR2_X1 U5740 ( .A1(n4641), .A2(n5130), .ZN(n5968) );
  INV_X1 U5741 ( .A(REIP_REG_5__SCAN_IN), .ZN(n4642) );
  OAI22_X1 U5742 ( .A1(n6177), .A2(n5968), .B1(n6175), .B2(n4642), .ZN(n4643)
         );
  AOI21_X1 U5743 ( .B1(n6189), .B2(n4644), .A(n4643), .ZN(n4645) );
  OAI21_X1 U5744 ( .B1(n5815), .B2(n6122), .A(n4645), .ZN(U3013) );
  NOR2_X1 U5745 ( .A1(n5078), .A2(n4980), .ZN(n4650) );
  NAND2_X1 U5746 ( .A1(n5084), .A2(n5644), .ZN(n6269) );
  OR2_X1 U5747 ( .A1(n4829), .A2(n4586), .ZN(n4688) );
  AOI21_X1 U5748 ( .B1(n6277), .B2(STATEBS16_REG_SCAN_IN), .A(n6275), .ZN(
        n6279) );
  OAI21_X1 U5749 ( .B1(n6268), .B2(n6269), .A(n6279), .ZN(n4649) );
  NAND3_X1 U5750 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n6441), .A3(n6436), .ZN(n6281) );
  OR2_X1 U5751 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6281), .ZN(n5073)
         );
  AND2_X1 U5752 ( .A1(n4652), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6239) );
  INV_X1 U5753 ( .A(n4647), .ZN(n4806) );
  INV_X1 U5754 ( .A(n5146), .ZN(n6308) );
  NOR2_X1 U5755 ( .A1(n4806), .A2(n6308), .ZN(n4986) );
  OAI21_X1 U5756 ( .B1(n4986), .B2(n5155), .A(n4845), .ZN(n4983) );
  AOI211_X1 U5757 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5073), .A(n6239), .B(
        n4983), .ZN(n4648) );
  NAND2_X1 U5758 ( .A1(n5071), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4655) );
  INV_X1 U5759 ( .A(n6277), .ZN(n4651) );
  NOR2_X2 U5760 ( .A1(n4651), .A2(n6276), .ZN(n6302) );
  INV_X1 U5761 ( .A(n6407), .ZN(n4996) );
  NOR2_X1 U5762 ( .A1(n6269), .A2(n6275), .ZN(n4896) );
  INV_X1 U5763 ( .A(n6311), .ZN(n4949) );
  NOR2_X1 U5764 ( .A1(n4652), .A2(n5155), .ZN(n6309) );
  AOI22_X1 U5765 ( .A1(n4896), .A2(n4949), .B1(n4986), .B2(n6309), .ZN(n5072)
         );
  INV_X1 U5766 ( .A(n6408), .ZN(n5189) );
  OAI22_X1 U5767 ( .A1(n4996), .A2(n5073), .B1(n5072), .B2(n5189), .ZN(n4653)
         );
  AOI21_X1 U5768 ( .B1(n6406), .B2(n6302), .A(n4653), .ZN(n4654) );
  OAI211_X1 U5769 ( .C1(n5078), .C2(n6411), .A(n4655), .B(n4654), .ZN(U3055)
         );
  NAND2_X1 U5770 ( .A1(n5071), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4658) );
  INV_X1 U5771 ( .A(n6358), .ZN(n4992) );
  OAI22_X1 U5772 ( .A1(n4992), .A2(n5073), .B1(n5072), .B2(n5179), .ZN(n4656)
         );
  AOI21_X1 U5773 ( .B1(n6359), .B2(n6302), .A(n4656), .ZN(n4657) );
  OAI211_X1 U5774 ( .C1(n5078), .C2(n6363), .A(n4658), .B(n4657), .ZN(U3056)
         );
  NAND2_X1 U5775 ( .A1(n5071), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4661) );
  INV_X1 U5776 ( .A(n6380), .ZN(n4988) );
  OAI22_X1 U5777 ( .A1(n4988), .A2(n5073), .B1(n5072), .B2(n5167), .ZN(n4659)
         );
  AOI21_X1 U5778 ( .B1(n6382), .B2(n6302), .A(n4659), .ZN(n4660) );
  OAI211_X1 U5779 ( .C1(n5078), .C2(n4900), .A(n4661), .B(n4660), .ZN(U3052)
         );
  INV_X1 U5780 ( .A(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4664) );
  NOR2_X2 U5781 ( .A1(n4703), .A2(n3641), .ZN(n6421) );
  INV_X1 U5782 ( .A(DATAI_6_), .ZN(n6067) );
  AOI22_X1 U5783 ( .A1(n6421), .A2(n4705), .B1(n6423), .B2(n4704), .ZN(n4663)
         );
  NAND2_X1 U5784 ( .A1(n6124), .A2(DATAI_30_), .ZN(n6428) );
  INV_X1 U5785 ( .A(n6428), .ZN(n6344) );
  NAND2_X1 U5786 ( .A1(n6124), .A2(DATAI_22_), .ZN(n6347) );
  INV_X1 U5787 ( .A(n6347), .ZN(n6418) );
  AOI22_X1 U5788 ( .A1(n6344), .A2(n4933), .B1(n5067), .B2(n6418), .ZN(n4662)
         );
  OAI211_X1 U5789 ( .C1(n4709), .C2(n4664), .A(n4663), .B(n4662), .ZN(U3146)
         );
  INV_X1 U5790 ( .A(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4667) );
  NOR2_X2 U5791 ( .A1(n4703), .A2(n3205), .ZN(n6401) );
  AOI22_X1 U5792 ( .A1(n6401), .A2(n4705), .B1(n6402), .B2(n4704), .ZN(n4666)
         );
  NAND2_X1 U5793 ( .A1(n4403), .A2(DATAI_26_), .ZN(n6405) );
  INV_X1 U5794 ( .A(n6405), .ZN(n6328) );
  NAND2_X1 U5795 ( .A1(n6124), .A2(DATAI_18_), .ZN(n6331) );
  INV_X1 U5796 ( .A(n6331), .ZN(n6400) );
  AOI22_X1 U5797 ( .A1(n6328), .A2(n4933), .B1(n5067), .B2(n6400), .ZN(n4665)
         );
  OAI211_X1 U5798 ( .C1(n4709), .C2(n4667), .A(n4666), .B(n4665), .ZN(U3142)
         );
  OR3_X1 U5799 ( .A1(n4829), .A2(n4689), .A3(n5642), .ZN(n4673) );
  INV_X1 U5800 ( .A(n4673), .ZN(n4668) );
  INV_X1 U5801 ( .A(n6269), .ZN(n4888) );
  NAND3_X1 U5802 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n6436), .ZN(n4889) );
  NOR2_X1 U5803 ( .A1(n6430), .A2(n4889), .ZN(n4786) );
  AOI21_X1 U5804 ( .B1(n4769), .B2(n4888), .A(n4786), .ZN(n4672) );
  INV_X1 U5805 ( .A(n4672), .ZN(n4670) );
  NAND2_X1 U5806 ( .A1(n4668), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4753) );
  NAND2_X1 U5807 ( .A1(n6313), .A2(n4753), .ZN(n4671) );
  AOI21_X1 U5808 ( .B1(n6275), .B2(n4889), .A(n4958), .ZN(n4669) );
  OAI21_X1 U5809 ( .B1(n4670), .B2(n4671), .A(n4669), .ZN(n4785) );
  OAI22_X1 U5810 ( .A1(n4672), .A2(n4671), .B1(n5155), .B2(n4889), .ZN(n4784)
         );
  AOI22_X1 U5811 ( .A1(INSTQUEUE_REG_13__3__SCAN_IN), .A2(n4785), .B1(n6408), 
        .B2(n4784), .ZN(n4675) );
  NOR2_X2 U5812 ( .A1(n4673), .A2(n6276), .ZN(n5059) );
  AOI22_X1 U5813 ( .A1(n6407), .A2(n4786), .B1(n6332), .B2(n5059), .ZN(n4674)
         );
  OAI211_X1 U5814 ( .C1(n6335), .C2(n4851), .A(n4675), .B(n4674), .ZN(U3127)
         );
  AOI22_X1 U5815 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n4785), .B1(n6373), 
        .B2(n4784), .ZN(n4677) );
  AOI22_X1 U5816 ( .A1(n6369), .A2(n4786), .B1(n6351), .B2(n5059), .ZN(n4676)
         );
  OAI211_X1 U5817 ( .C1(n6355), .C2(n4851), .A(n4677), .B(n4676), .ZN(U3131)
         );
  NAND2_X1 U5818 ( .A1(n6124), .A2(DATAI_21_), .ZN(n6343) );
  INV_X1 U5819 ( .A(DATAI_5_), .ZN(n6065) );
  AOI22_X1 U5820 ( .A1(INSTQUEUE_REG_13__5__SCAN_IN), .A2(n4785), .B1(n6414), 
        .B2(n4784), .ZN(n4680) );
  NOR2_X1 U5821 ( .A1(n4703), .A2(n3208), .ZN(n6413) );
  NAND2_X1 U5822 ( .A1(n6124), .A2(DATAI_29_), .ZN(n6417) );
  INV_X1 U5823 ( .A(n6417), .ZN(n6340) );
  AOI22_X1 U5824 ( .A1(n6413), .A2(n4786), .B1(n6340), .B2(n5059), .ZN(n4679)
         );
  OAI211_X1 U5825 ( .C1(n6343), .C2(n4851), .A(n4680), .B(n4679), .ZN(U3129)
         );
  AOI22_X1 U5826 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n4785), .B1(n6360), 
        .B2(n4784), .ZN(n4682) );
  AOI22_X1 U5827 ( .A1(n6358), .A2(n4786), .B1(n6336), .B2(n5059), .ZN(n4681)
         );
  OAI211_X1 U5828 ( .C1(n6339), .C2(n4851), .A(n4682), .B(n4681), .ZN(U3128)
         );
  AOI22_X1 U5829 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n4785), .B1(n6383), 
        .B2(n4784), .ZN(n4684) );
  AOI22_X1 U5830 ( .A1(n6380), .A2(n4786), .B1(n6381), .B2(n5059), .ZN(n4683)
         );
  OAI211_X1 U5831 ( .C1(n6324), .C2(n4851), .A(n4684), .B(n4683), .ZN(U3124)
         );
  NAND2_X1 U5832 ( .A1(n5071), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4687) );
  INV_X1 U5833 ( .A(n5072), .ZN(n4791) );
  INV_X1 U5834 ( .A(n6302), .ZN(n4789) );
  OAI22_X1 U5835 ( .A1(n5010), .A2(n5073), .B1(n4789), .B2(n6355), .ZN(n4685)
         );
  AOI21_X1 U5836 ( .B1(n6373), .B2(n4791), .A(n4685), .ZN(n4686) );
  OAI211_X1 U5837 ( .C1(n5078), .C2(n6378), .A(n4687), .B(n4686), .ZN(U3059)
         );
  INV_X1 U5838 ( .A(n4829), .ZN(n4690) );
  NAND3_X1 U5839 ( .A1(n4690), .A2(n4689), .A3(n5645), .ZN(n4755) );
  NAND2_X1 U5840 ( .A1(n4755), .A2(n6313), .ZN(n4696) );
  AND2_X1 U5841 ( .A1(n4842), .A2(n4691), .ZN(n6315) );
  INV_X1 U5842 ( .A(n4692), .ZN(n6368) );
  AOI21_X1 U5843 ( .B1(n6315), .B2(n4860), .A(n6368), .ZN(n4693) );
  OAI22_X1 U5844 ( .A1(n4696), .A2(n4693), .B1(n6307), .B2(n5155), .ZN(n6372)
         );
  INV_X1 U5845 ( .A(n4693), .ZN(n4695) );
  AOI21_X1 U5846 ( .B1(n6275), .B2(n6307), .A(n4958), .ZN(n4694) );
  OAI21_X1 U5847 ( .B1(n4696), .B2(n4695), .A(n4694), .ZN(n6374) );
  AOI22_X1 U5848 ( .A1(n6383), .A2(n6372), .B1(n6374), .B2(
        INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4699) );
  AOI22_X1 U5849 ( .A1(n6382), .A2(n6370), .B1(n6380), .B2(n6368), .ZN(n4698)
         );
  OAI211_X1 U5850 ( .C1(n4900), .C2(n6377), .A(n4699), .B(n4698), .ZN(U3076)
         );
  AOI22_X1 U5851 ( .A1(n6408), .A2(n6372), .B1(n6374), .B2(
        INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4701) );
  AOI22_X1 U5852 ( .A1(n6406), .A2(n6370), .B1(n6407), .B2(n6368), .ZN(n4700)
         );
  OAI211_X1 U5853 ( .C1(n6411), .C2(n6377), .A(n4701), .B(n4700), .ZN(U3079)
         );
  INV_X1 U5854 ( .A(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4708) );
  AOI22_X1 U5855 ( .A1(n3193), .A2(n4705), .B1(n6396), .B2(n4704), .ZN(n4707)
         );
  NAND2_X1 U5856 ( .A1(n6124), .A2(DATAI_25_), .ZN(n6399) );
  INV_X1 U5857 ( .A(n6399), .ZN(n6387) );
  NAND2_X1 U5858 ( .A1(n6124), .A2(DATAI_17_), .ZN(n6327) );
  INV_X1 U5859 ( .A(n6327), .ZN(n6394) );
  AOI22_X1 U5860 ( .A1(n6387), .A2(n4933), .B1(n5067), .B2(n6394), .ZN(n4706)
         );
  OAI211_X1 U5861 ( .C1(n4709), .C2(n4708), .A(n4707), .B(n4706), .ZN(U3141)
         );
  AOI22_X1 U5862 ( .A1(INSTQUEUE_REG_13__6__SCAN_IN), .A2(n4785), .B1(n6423), 
        .B2(n4784), .ZN(n4711) );
  AOI22_X1 U5863 ( .A1(n6421), .A2(n4786), .B1(n6344), .B2(n5059), .ZN(n4710)
         );
  OAI211_X1 U5864 ( .C1(n6347), .C2(n4851), .A(n4711), .B(n4710), .ZN(U3130)
         );
  AOI22_X1 U5865 ( .A1(INSTQUEUE_REG_13__2__SCAN_IN), .A2(n4785), .B1(n6402), 
        .B2(n4784), .ZN(n4713) );
  AOI22_X1 U5866 ( .A1(n6401), .A2(n4786), .B1(n6328), .B2(n5059), .ZN(n4712)
         );
  OAI211_X1 U5867 ( .C1(n6331), .C2(n4851), .A(n4713), .B(n4712), .ZN(U3126)
         );
  AOI21_X1 U5868 ( .B1(n4716), .B2(n4715), .A(n5120), .ZN(n4717) );
  INV_X1 U5869 ( .A(n4717), .ZN(n6121) );
  XNOR2_X1 U5870 ( .A(n5130), .B(n5128), .ZN(n6190) );
  AOI22_X1 U5871 ( .A1(n5445), .A2(n6190), .B1(n5462), .B2(EBX_REG_6__SCAN_IN), 
        .ZN(n4718) );
  OAI21_X1 U5872 ( .B1(n6121), .B2(n3195), .A(n4718), .ZN(U2853) );
  OAI22_X1 U5873 ( .A1(n5102), .A2(n4719), .B1(n3436), .B2(n4744), .ZN(n4721)
         );
  NAND2_X1 U5874 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n5832), .ZN(n4748) );
  INV_X1 U5875 ( .A(n4748), .ZN(n4720) );
  AOI22_X1 U5876 ( .A1(n4721), .A2(n6736), .B1(n4720), .B2(
        INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4751) );
  INV_X1 U5877 ( .A(n4722), .ZN(n4747) );
  NAND2_X1 U5878 ( .A1(n4724), .A2(n4723), .ZN(n4741) );
  XNOR2_X1 U5879 ( .A(n5332), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4729)
         );
  XNOR2_X1 U5880 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4725) );
  OAI22_X1 U5881 ( .A1(n4731), .A2(n4725), .B1(n4733), .B2(n4729), .ZN(n4728)
         );
  INV_X1 U5882 ( .A(n5084), .ZN(n4726) );
  NOR2_X1 U5883 ( .A1(n4726), .A2(n5326), .ZN(n4727) );
  AOI211_X1 U5884 ( .C1(n4741), .C2(n4729), .A(n4728), .B(n4727), .ZN(n5331)
         );
  NAND2_X1 U5885 ( .A1(n5331), .A2(n4744), .ZN(n4730) );
  OAI21_X1 U5886 ( .B1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n4744), .A(n4730), 
        .ZN(n6439) );
  INV_X1 U5887 ( .A(n6439), .ZN(n4745) );
  INV_X1 U5888 ( .A(n4731), .ZN(n6431) );
  NAND2_X1 U5889 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4732) );
  XNOR2_X1 U5890 ( .A(n4732), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4737)
         );
  INV_X1 U5891 ( .A(n4733), .ZN(n4736) );
  INV_X1 U5892 ( .A(n5332), .ZN(n5338) );
  AOI211_X1 U5893 ( .C1(n4734), .C2(n5338), .A(n4738), .B(n4735), .ZN(n6549)
         );
  AOI22_X1 U5894 ( .A1(n6431), .A2(n4737), .B1(n4736), .B2(n6549), .ZN(n4743)
         );
  INV_X1 U5895 ( .A(n4738), .ZN(n4739) );
  MUX2_X1 U5896 ( .A(n4739), .B(n4734), .S(n5332), .Z(n4740) );
  NAND3_X1 U5897 ( .A1(n4741), .A2(n4747), .A3(n4740), .ZN(n4742) );
  OAI211_X1 U5898 ( .C1(n4949), .C2(n5326), .A(n4743), .B(n4742), .ZN(n6551)
         );
  MUX2_X1 U5899 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n6551), .S(n4744), 
        .Z(n6442) );
  NAND3_X1 U5900 ( .A1(n4745), .A2(n6442), .A3(n6736), .ZN(n4746) );
  OAI211_X1 U5901 ( .C1(n4748), .C2(n4747), .A(n4746), .B(n4751), .ZN(n6449)
         );
  INV_X1 U5902 ( .A(n6449), .ZN(n4749) );
  AOI21_X1 U5903 ( .B1(n4751), .B2(n4750), .A(n4749), .ZN(n4762) );
  NOR2_X1 U5904 ( .A1(n4762), .A2(FLUSH_REG_SCAN_IN), .ZN(n4752) );
  INV_X1 U5905 ( .A(n4753), .ZN(n4754) );
  AOI21_X1 U5906 ( .B1(n4857), .B2(n4829), .A(n4754), .ZN(n4948) );
  AOI21_X1 U5907 ( .B1(n4948), .B2(n4755), .A(n6275), .ZN(n4758) );
  NAND2_X1 U5908 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6547), .ZN(n4830) );
  INV_X1 U5909 ( .A(n4830), .ZN(n5643) );
  OAI22_X1 U5910 ( .A1(n4756), .A2(n6316), .B1(n4949), .B2(n5643), .ZN(n4757)
         );
  OAI21_X1 U5911 ( .B1(n4758), .B2(n4757), .A(n6236), .ZN(n4759) );
  OAI21_X1 U5912 ( .B1(n6236), .B2(n6441), .A(n4759), .ZN(U3462) );
  INV_X1 U5913 ( .A(n4760), .ZN(n4761) );
  NOR2_X1 U5914 ( .A1(n4762), .A2(n4761), .ZN(n6456) );
  OAI22_X1 U5915 ( .A1(n4866), .A2(n6275), .B1(n6267), .B2(n5643), .ZN(n4763)
         );
  OAI21_X1 U5916 ( .B1(n6456), .B2(n4763), .A(n6236), .ZN(n4764) );
  OAI21_X1 U5917 ( .B1(n6236), .B2(n6430), .A(n4764), .ZN(U3465) );
  NAND2_X1 U5918 ( .A1(n4765), .A2(n4829), .ZN(n4856) );
  INV_X1 U5919 ( .A(n4856), .ZN(n4766) );
  NAND2_X1 U5920 ( .A1(n4766), .A2(n4857), .ZN(n4775) );
  NAND3_X1 U5921 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n4859), .A3(n6436), .ZN(n4805) );
  INV_X1 U5922 ( .A(n4805), .ZN(n4772) );
  OAI21_X1 U5923 ( .B1(n4775), .B2(n6564), .A(n6313), .ZN(n4774) );
  INV_X1 U5924 ( .A(n4774), .ZN(n4770) );
  INV_X1 U5925 ( .A(n4858), .ZN(n4768) );
  NOR2_X1 U5926 ( .A1(n6430), .A2(n4805), .ZN(n6386) );
  AOI21_X1 U5927 ( .B1(n4769), .B2(n4768), .A(n6386), .ZN(n4773) );
  NAND2_X1 U5928 ( .A1(n4770), .A2(n4773), .ZN(n4771) );
  OAI211_X1 U5929 ( .C1(n6313), .C2(n4772), .A(n4771), .B(n6272), .ZN(n6379)
         );
  OAI22_X1 U5930 ( .A1(n4774), .A2(n4773), .B1(n4805), .B2(n5155), .ZN(n6390)
         );
  AOI22_X1 U5931 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n6379), .B1(n6414), 
        .B2(n6390), .ZN(n4777) );
  NOR2_X2 U5932 ( .A1(n4775), .A2(n6276), .ZN(n6388) );
  AOI22_X1 U5933 ( .A1(n6388), .A2(n6340), .B1(n6413), .B2(n6386), .ZN(n4776)
         );
  OAI211_X1 U5934 ( .C1(n6343), .C2(n5148), .A(n4777), .B(n4776), .ZN(U3097)
         );
  AOI22_X1 U5935 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n6379), .B1(n6360), 
        .B2(n6390), .ZN(n4779) );
  AOI22_X1 U5936 ( .A1(n6388), .A2(n6336), .B1(n6358), .B2(n6386), .ZN(n4778)
         );
  OAI211_X1 U5937 ( .C1(n6339), .C2(n5148), .A(n4779), .B(n4778), .ZN(U3096)
         );
  AOI22_X1 U5938 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n6379), .B1(n6373), 
        .B2(n6390), .ZN(n4781) );
  AOI22_X1 U5939 ( .A1(n6388), .A2(n6351), .B1(n6369), .B2(n6386), .ZN(n4780)
         );
  OAI211_X1 U5940 ( .C1(n6355), .C2(n5148), .A(n4781), .B(n4780), .ZN(U3099)
         );
  AOI22_X1 U5941 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n6379), .B1(n6408), 
        .B2(n6390), .ZN(n4783) );
  AOI22_X1 U5942 ( .A1(n6388), .A2(n6332), .B1(n6407), .B2(n6386), .ZN(n4782)
         );
  OAI211_X1 U5943 ( .C1(n6335), .C2(n5148), .A(n4783), .B(n4782), .ZN(U3095)
         );
  AOI22_X1 U5944 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(n4785), .B1(n6396), 
        .B2(n4784), .ZN(n4788) );
  AOI22_X1 U5945 ( .A1(n3193), .A2(n4786), .B1(n6387), .B2(n5059), .ZN(n4787)
         );
  OAI211_X1 U5946 ( .C1(n6327), .C2(n4851), .A(n4788), .B(n4787), .ZN(U3125)
         );
  NAND2_X1 U5947 ( .A1(n5071), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4793) );
  INV_X1 U5948 ( .A(n6413), .ZN(n5017) );
  OAI22_X1 U5949 ( .A1(n5017), .A2(n5073), .B1(n4789), .B2(n6343), .ZN(n4790)
         );
  AOI21_X1 U5950 ( .B1(n6414), .B2(n4791), .A(n4790), .ZN(n4792) );
  OAI211_X1 U5951 ( .C1(n5078), .C2(n6417), .A(n4793), .B(n4792), .ZN(U3057)
         );
  XNOR2_X1 U5952 ( .A(n4578), .B(n3726), .ZN(n6123) );
  INV_X1 U5953 ( .A(n6123), .ZN(n4797) );
  INV_X1 U5954 ( .A(EBX_REG_5__SCAN_IN), .ZN(n4795) );
  OAI222_X1 U5955 ( .A1(n5968), .A2(n5466), .B1(n3195), .B2(n4797), .C1(n5453), 
        .C2(n4795), .ZN(U2854) );
  OAI222_X1 U5956 ( .A1(n6065), .A2(n6969), .B1(n6970), .B2(n4797), .C1(n6967), 
        .C2(n4796), .ZN(U2886) );
  INV_X1 U5957 ( .A(n6414), .ZN(n5159) );
  OAI22_X1 U5958 ( .A1(n5017), .A2(n4798), .B1(n6343), .B2(n5003), .ZN(n4799)
         );
  AOI21_X1 U5959 ( .B1(n6340), .B2(n4933), .A(n4799), .ZN(n4802) );
  NAND2_X1 U5960 ( .A1(n4800), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4801)
         );
  OAI211_X1 U5961 ( .C1(n4803), .C2(n5159), .A(n4802), .B(n4801), .ZN(U3145)
         );
  INV_X1 U5962 ( .A(n6388), .ZN(n5022) );
  NAND3_X1 U5963 ( .A1(n5022), .A2(n6313), .A3(n5015), .ZN(n4804) );
  NOR2_X1 U5964 ( .A1(n4949), .A2(n4858), .ZN(n4810) );
  AOI21_X1 U5965 ( .B1(n4804), .B2(n6316), .A(n4810), .ZN(n4809) );
  NOR2_X1 U5966 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4805), .ZN(n5009)
         );
  INV_X1 U5967 ( .A(n6309), .ZN(n4837) );
  NAND2_X1 U5968 ( .A1(n4806), .A2(n5146), .ZN(n4894) );
  AOI21_X1 U5969 ( .B1(n4894), .B2(STATE2_REG_2__SCAN_IN), .A(n4807), .ZN(
        n4890) );
  OAI211_X1 U5970 ( .C1(n6547), .C2(n5009), .A(n4837), .B(n4890), .ZN(n4808)
         );
  INV_X1 U5971 ( .A(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4815) );
  INV_X1 U5972 ( .A(n4810), .ZN(n4811) );
  INV_X1 U5973 ( .A(n6239), .ZN(n6318) );
  OAI22_X1 U5974 ( .A1(n4811), .A2(n6275), .B1(n6318), .B2(n4894), .ZN(n5019)
         );
  AOI22_X1 U5975 ( .A1(n6380), .A2(n5009), .B1(n6383), .B2(n5019), .ZN(n4812)
         );
  OAI21_X1 U5976 ( .B1(n4900), .B2(n5015), .A(n4812), .ZN(n4813) );
  AOI21_X1 U5977 ( .B1(n6382), .B2(n6388), .A(n4813), .ZN(n4814) );
  OAI21_X1 U5978 ( .B1(n5008), .B2(n4815), .A(n4814), .ZN(U3084) );
  INV_X1 U5979 ( .A(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4819) );
  AOI22_X1 U5980 ( .A1(n6358), .A2(n5009), .B1(n6360), .B2(n5019), .ZN(n4816)
         );
  OAI21_X1 U5981 ( .B1(n6363), .B2(n5015), .A(n4816), .ZN(n4817) );
  AOI21_X1 U5982 ( .B1(n6359), .B2(n6388), .A(n4817), .ZN(n4818) );
  OAI21_X1 U5983 ( .B1(n5008), .B2(n4819), .A(n4818), .ZN(U3088) );
  INV_X1 U5984 ( .A(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4823) );
  AOI22_X1 U5985 ( .A1(n6407), .A2(n5009), .B1(n6408), .B2(n5019), .ZN(n4820)
         );
  OAI21_X1 U5986 ( .B1(n6411), .B2(n5015), .A(n4820), .ZN(n4821) );
  AOI21_X1 U5987 ( .B1(n6406), .B2(n6388), .A(n4821), .ZN(n4822) );
  OAI21_X1 U5988 ( .B1(n5008), .B2(n4823), .A(n4822), .ZN(U3087) );
  AOI22_X1 U5989 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n6379), .B1(n6402), 
        .B2(n6390), .ZN(n4825) );
  AOI22_X1 U5990 ( .A1(n6388), .A2(n6328), .B1(n6401), .B2(n6386), .ZN(n4824)
         );
  OAI211_X1 U5991 ( .C1(n6331), .C2(n5148), .A(n4825), .B(n4824), .ZN(U3094)
         );
  AOI22_X1 U5992 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n6379), .B1(n6423), 
        .B2(n6390), .ZN(n4827) );
  AOI22_X1 U5993 ( .A1(n6388), .A2(n6344), .B1(n6421), .B2(n6386), .ZN(n4826)
         );
  OAI211_X1 U5994 ( .C1(n6347), .C2(n5148), .A(n4827), .B(n4826), .ZN(U3098)
         );
  INV_X1 U5995 ( .A(n6236), .ZN(n4834) );
  OAI21_X1 U5996 ( .B1(n5645), .B2(n4829), .A(n4828), .ZN(n4831) );
  AOI22_X1 U5997 ( .A1(n4831), .A2(n6313), .B1(n4830), .B2(n5084), .ZN(n4833)
         );
  NAND2_X1 U5998 ( .A1(n4834), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4832) );
  OAI21_X1 U5999 ( .B1(n4834), .B2(n4833), .A(n4832), .ZN(U3463) );
  INV_X1 U6000 ( .A(EAX_REG_6__SCAN_IN), .ZN(n6900) );
  OAI222_X1 U6001 ( .A1(n6121), .A2(n6970), .B1(n6969), .B2(n6067), .C1(n6967), 
        .C2(n6900), .ZN(U2885) );
  AOI22_X1 U6002 ( .A1(n6396), .A2(n6372), .B1(n6374), .B2(
        INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4836) );
  AOI22_X1 U6003 ( .A1(n6394), .A2(n6370), .B1(n3193), .B2(n6368), .ZN(n4835)
         );
  OAI211_X1 U6004 ( .C1(n6399), .C2(n6377), .A(n4836), .B(n4835), .ZN(U3077)
         );
  NAND2_X1 U6005 ( .A1(n4842), .A2(n6313), .ZN(n6312) );
  INV_X1 U6006 ( .A(n6312), .ZN(n4839) );
  NOR3_X1 U6007 ( .A1(n4837), .A2(n6441), .A3(n5146), .ZN(n4838) );
  AOI21_X1 U6008 ( .B1(n4839), .B2(n6311), .A(n4838), .ZN(n4915) );
  NOR2_X1 U6009 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4840), .ZN(n4932)
         );
  INV_X1 U6010 ( .A(n4932), .ZN(n4852) );
  OAI22_X1 U6011 ( .A1(n5010), .A2(n4852), .B1(n6378), .B2(n4851), .ZN(n4841)
         );
  AOI21_X1 U6012 ( .B1(n6371), .B2(n4933), .A(n4841), .ZN(n4850) );
  INV_X1 U6013 ( .A(n4842), .ZN(n4844) );
  OAI21_X1 U6014 ( .B1(n4934), .B2(n4933), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n4843) );
  NAND3_X1 U6015 ( .A1(n4844), .A2(n6313), .A3(n4843), .ZN(n4848) );
  NAND2_X1 U6016 ( .A1(n5146), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4846) );
  NAND2_X1 U6017 ( .A1(n4846), .A2(n4845), .ZN(n6320) );
  NOR3_X1 U6018 ( .A1(n6320), .A2(n6441), .A3(n6239), .ZN(n4847) );
  OAI211_X1 U6019 ( .C1(n4932), .C2(n6547), .A(n4848), .B(n4847), .ZN(n4914)
         );
  NAND2_X1 U6020 ( .A1(n4914), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4849)
         );
  OAI211_X1 U6021 ( .C1(n4915), .C2(n5163), .A(n4850), .B(n4849), .ZN(U3139)
         );
  INV_X1 U6022 ( .A(n6343), .ZN(n6412) );
  OAI22_X1 U6023 ( .A1(n5017), .A2(n4852), .B1(n6417), .B2(n4851), .ZN(n4853)
         );
  AOI21_X1 U6024 ( .B1(n6412), .B2(n4933), .A(n4853), .ZN(n4855) );
  NAND2_X1 U6025 ( .A1(n4914), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4854)
         );
  OAI211_X1 U6026 ( .C1(n4915), .C2(n5159), .A(n4855), .B(n4854), .ZN(U3137)
         );
  NOR2_X1 U6027 ( .A1(n6311), .A2(n4858), .ZN(n4987) );
  NAND3_X1 U6028 ( .A1(n6441), .A2(n4859), .A3(n6436), .ZN(n4982) );
  NOR2_X1 U6029 ( .A1(n6430), .A2(n4982), .ZN(n4884) );
  AOI21_X1 U6030 ( .B1(n4987), .B2(n4860), .A(n4884), .ZN(n4864) );
  OR2_X1 U6031 ( .A1(n4867), .A2(n6564), .ZN(n4861) );
  AND2_X1 U6032 ( .A1(n4861), .A2(n6313), .ZN(n4863) );
  AOI22_X1 U6033 ( .A1(n4864), .A2(n4863), .B1(n6275), .B2(n4982), .ZN(n4862)
         );
  NAND2_X1 U6034 ( .A1(n6272), .A2(n4862), .ZN(n4883) );
  INV_X1 U6035 ( .A(n4863), .ZN(n4865) );
  OAI22_X1 U6036 ( .A1(n4865), .A2(n4864), .B1(n5155), .B2(n4982), .ZN(n4882)
         );
  AOI22_X1 U6037 ( .A1(INSTQUEUE_REG_1__3__SCAN_IN), .A2(n4883), .B1(n6408), 
        .B2(n4882), .ZN(n4869) );
  NOR2_X2 U6038 ( .A1(n4867), .A2(n4866), .ZN(n6262) );
  AOI22_X1 U6039 ( .A1(n4884), .A2(n6407), .B1(n6262), .B2(n6406), .ZN(n4868)
         );
  OAI211_X1 U6040 ( .C1(n5070), .C2(n6411), .A(n4869), .B(n4868), .ZN(U3031)
         );
  AOI22_X1 U6041 ( .A1(INSTQUEUE_REG_1__6__SCAN_IN), .A2(n4883), .B1(n6423), 
        .B2(n4882), .ZN(n4871) );
  AOI22_X1 U6042 ( .A1(n4884), .A2(n6421), .B1(n6262), .B2(n6418), .ZN(n4870)
         );
  OAI211_X1 U6043 ( .C1(n5070), .C2(n6428), .A(n4871), .B(n4870), .ZN(U3034)
         );
  AOI22_X1 U6044 ( .A1(INSTQUEUE_REG_1__7__SCAN_IN), .A2(n4883), .B1(n6373), 
        .B2(n4882), .ZN(n4873) );
  AOI22_X1 U6045 ( .A1(n4884), .A2(n6369), .B1(n6262), .B2(n6371), .ZN(n4872)
         );
  OAI211_X1 U6046 ( .C1(n5070), .C2(n6378), .A(n4873), .B(n4872), .ZN(U3035)
         );
  AOI22_X1 U6047 ( .A1(INSTQUEUE_REG_1__5__SCAN_IN), .A2(n4883), .B1(n6414), 
        .B2(n4882), .ZN(n4875) );
  AOI22_X1 U6048 ( .A1(n4884), .A2(n6413), .B1(n6262), .B2(n6412), .ZN(n4874)
         );
  OAI211_X1 U6049 ( .C1(n5070), .C2(n6417), .A(n4875), .B(n4874), .ZN(U3033)
         );
  AOI22_X1 U6050 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(n4883), .B1(n6383), 
        .B2(n4882), .ZN(n4877) );
  AOI22_X1 U6051 ( .A1(n6380), .A2(n4884), .B1(n6262), .B2(n6382), .ZN(n4876)
         );
  OAI211_X1 U6052 ( .C1(n5070), .C2(n4900), .A(n4877), .B(n4876), .ZN(U3028)
         );
  AOI22_X1 U6053 ( .A1(INSTQUEUE_REG_1__2__SCAN_IN), .A2(n4883), .B1(n6402), 
        .B2(n4882), .ZN(n4879) );
  AOI22_X1 U6054 ( .A1(n4884), .A2(n6401), .B1(n6262), .B2(n6400), .ZN(n4878)
         );
  OAI211_X1 U6055 ( .C1(n5070), .C2(n6405), .A(n4879), .B(n4878), .ZN(U3030)
         );
  AOI22_X1 U6056 ( .A1(INSTQUEUE_REG_1__1__SCAN_IN), .A2(n4883), .B1(n6396), 
        .B2(n4882), .ZN(n4881) );
  AOI22_X1 U6057 ( .A1(n4884), .A2(n3193), .B1(n6262), .B2(n6394), .ZN(n4880)
         );
  OAI211_X1 U6058 ( .C1(n5070), .C2(n6399), .A(n4881), .B(n4880), .ZN(U3029)
         );
  AOI22_X1 U6059 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n4883), .B1(n6360), 
        .B2(n4882), .ZN(n4886) );
  AOI22_X1 U6060 ( .A1(n4884), .A2(n6358), .B1(n6262), .B2(n6359), .ZN(n4885)
         );
  OAI211_X1 U6061 ( .C1(n5070), .C2(n6363), .A(n4886), .B(n4885), .ZN(U3032)
         );
  INV_X1 U6062 ( .A(n5059), .ZN(n4910) );
  AOI21_X1 U6063 ( .B1(n4910), .B2(n5062), .A(n6564), .ZN(n4887) );
  AOI211_X1 U6064 ( .C1(n4888), .C2(n6268), .A(n6275), .B(n4887), .ZN(n4892)
         );
  NOR2_X1 U6065 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4889), .ZN(n4893)
         );
  OAI211_X1 U6066 ( .C1(n6547), .C2(n4893), .A(n6318), .B(n4890), .ZN(n4891)
         );
  NAND2_X1 U6067 ( .A1(n5055), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n4899)
         );
  INV_X1 U6068 ( .A(n4893), .ZN(n5057) );
  INV_X1 U6069 ( .A(n4894), .ZN(n4895) );
  AOI22_X1 U6070 ( .A1(n4896), .A2(n6311), .B1(n6309), .B2(n4895), .ZN(n5056)
         );
  OAI22_X1 U6071 ( .A1(n4988), .A2(n5057), .B1(n5056), .B2(n5167), .ZN(n4897)
         );
  AOI21_X1 U6072 ( .B1(n6382), .B2(n5059), .A(n4897), .ZN(n4898) );
  OAI211_X1 U6073 ( .C1(n5062), .C2(n4900), .A(n4899), .B(n4898), .ZN(U3116)
         );
  NAND2_X1 U6074 ( .A1(n5055), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4903)
         );
  OAI22_X1 U6075 ( .A1(n4992), .A2(n5057), .B1(n5056), .B2(n5179), .ZN(n4901)
         );
  AOI21_X1 U6076 ( .B1(n6359), .B2(n5059), .A(n4901), .ZN(n4902) );
  OAI211_X1 U6077 ( .C1(n5062), .C2(n6363), .A(n4903), .B(n4902), .ZN(U3120)
         );
  NAND2_X1 U6078 ( .A1(n5055), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4906)
         );
  OAI22_X1 U6079 ( .A1(n4996), .A2(n5057), .B1(n5056), .B2(n5189), .ZN(n4904)
         );
  AOI21_X1 U6080 ( .B1(n6406), .B2(n5059), .A(n4904), .ZN(n4905) );
  OAI211_X1 U6081 ( .C1(n5062), .C2(n6411), .A(n4906), .B(n4905), .ZN(U3119)
         );
  NAND2_X1 U6082 ( .A1(n5055), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4909)
         );
  OAI22_X1 U6083 ( .A1(n5010), .A2(n5057), .B1(n6355), .B2(n4910), .ZN(n4907)
         );
  AOI21_X1 U6084 ( .B1(n6351), .B2(n6419), .A(n4907), .ZN(n4908) );
  OAI211_X1 U6085 ( .C1(n5056), .C2(n5163), .A(n4909), .B(n4908), .ZN(U3123)
         );
  NAND2_X1 U6086 ( .A1(n5055), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4913)
         );
  OAI22_X1 U6087 ( .A1(n5017), .A2(n5057), .B1(n6343), .B2(n4910), .ZN(n4911)
         );
  AOI21_X1 U6088 ( .B1(n6340), .B2(n6419), .A(n4911), .ZN(n4912) );
  OAI211_X1 U6089 ( .C1(n5056), .C2(n5159), .A(n4913), .B(n4912), .ZN(U3121)
         );
  INV_X1 U6090 ( .A(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4918) );
  INV_X1 U6091 ( .A(n4915), .ZN(n4931) );
  AOI22_X1 U6092 ( .A1(n6407), .A2(n4932), .B1(n6408), .B2(n4931), .ZN(n4917)
         );
  AOI22_X1 U6093 ( .A1(n4934), .A2(n6332), .B1(n4933), .B2(n6406), .ZN(n4916)
         );
  OAI211_X1 U6094 ( .C1(n4938), .C2(n4918), .A(n4917), .B(n4916), .ZN(U3135)
         );
  INV_X1 U6095 ( .A(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4921) );
  AOI22_X1 U6096 ( .A1(n6421), .A2(n4932), .B1(n6423), .B2(n4931), .ZN(n4920)
         );
  AOI22_X1 U6097 ( .A1(n4934), .A2(n6344), .B1(n4933), .B2(n6418), .ZN(n4919)
         );
  OAI211_X1 U6098 ( .C1(n4938), .C2(n4921), .A(n4920), .B(n4919), .ZN(U3138)
         );
  INV_X1 U6099 ( .A(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4924) );
  AOI22_X1 U6100 ( .A1(n6380), .A2(n4932), .B1(n6383), .B2(n4931), .ZN(n4923)
         );
  AOI22_X1 U6101 ( .A1(n4934), .A2(n6381), .B1(n4933), .B2(n6382), .ZN(n4922)
         );
  OAI211_X1 U6102 ( .C1(n4938), .C2(n4924), .A(n4923), .B(n4922), .ZN(U3132)
         );
  INV_X1 U6103 ( .A(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4927) );
  AOI22_X1 U6104 ( .A1(n3193), .A2(n4932), .B1(n6396), .B2(n4931), .ZN(n4926)
         );
  AOI22_X1 U6105 ( .A1(n4934), .A2(n6387), .B1(n4933), .B2(n6394), .ZN(n4925)
         );
  OAI211_X1 U6106 ( .C1(n4938), .C2(n4927), .A(n4926), .B(n4925), .ZN(U3133)
         );
  INV_X1 U6107 ( .A(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4930) );
  AOI22_X1 U6108 ( .A1(n6401), .A2(n4932), .B1(n6402), .B2(n4931), .ZN(n4929)
         );
  AOI22_X1 U6109 ( .A1(n4934), .A2(n6328), .B1(n4933), .B2(n6400), .ZN(n4928)
         );
  OAI211_X1 U6110 ( .C1(n4938), .C2(n4930), .A(n4929), .B(n4928), .ZN(U3134)
         );
  INV_X1 U6111 ( .A(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4937) );
  AOI22_X1 U6112 ( .A1(n6358), .A2(n4932), .B1(n6360), .B2(n4931), .ZN(n4936)
         );
  AOI22_X1 U6113 ( .A1(n4934), .A2(n6336), .B1(n4933), .B2(n6359), .ZN(n4935)
         );
  OAI211_X1 U6114 ( .C1(n4938), .C2(n4937), .A(n4936), .B(n4935), .ZN(U3136)
         );
  INV_X1 U6115 ( .A(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4942) );
  AOI22_X1 U6116 ( .A1(n6421), .A2(n5009), .B1(n6423), .B2(n5019), .ZN(n4939)
         );
  OAI21_X1 U6117 ( .B1(n6428), .B2(n5015), .A(n4939), .ZN(n4940) );
  AOI21_X1 U6118 ( .B1(n6418), .B2(n6388), .A(n4940), .ZN(n4941) );
  OAI21_X1 U6119 ( .B1(n5008), .B2(n4942), .A(n4941), .ZN(U3090) );
  INV_X1 U6120 ( .A(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4946) );
  AOI22_X1 U6121 ( .A1(n6401), .A2(n5009), .B1(n6402), .B2(n5019), .ZN(n4943)
         );
  OAI21_X1 U6122 ( .B1(n6405), .B2(n5015), .A(n4943), .ZN(n4944) );
  AOI21_X1 U6123 ( .B1(n6400), .B2(n6388), .A(n4944), .ZN(n4945) );
  OAI21_X1 U6124 ( .B1(n5008), .B2(n4946), .A(n4945), .ZN(U3086) );
  AOI21_X1 U6125 ( .B1(n4948), .B2(n4947), .A(n6275), .ZN(n4957) );
  NAND2_X1 U6126 ( .A1(n4949), .A2(n3227), .ZN(n6242) );
  OR2_X1 U6127 ( .A1(n6242), .A2(n6267), .ZN(n4952) );
  INV_X1 U6128 ( .A(n4950), .ZN(n4951) );
  NAND2_X1 U6129 ( .A1(n4951), .A2(n6441), .ZN(n5049) );
  NAND2_X1 U6130 ( .A1(n4952), .A2(n5049), .ZN(n4960) );
  NAND2_X1 U6131 ( .A1(n4953), .A2(n6441), .ZN(n6238) );
  INV_X1 U6132 ( .A(n6238), .ZN(n4954) );
  AOI22_X1 U6133 ( .A1(n4957), .A2(n4960), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4954), .ZN(n5054) );
  OAI22_X1 U6134 ( .A1(n5010), .A2(n5049), .B1(n6355), .B2(n5078), .ZN(n4956)
         );
  AOI21_X1 U6135 ( .B1(n6351), .B2(n6241), .A(n4956), .ZN(n4963) );
  INV_X1 U6136 ( .A(n4957), .ZN(n4961) );
  AOI21_X1 U6137 ( .B1(n6275), .B2(n6238), .A(n4958), .ZN(n4959) );
  NAND2_X1 U6138 ( .A1(n5051), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4962) );
  OAI211_X1 U6139 ( .C1(n5054), .C2(n5163), .A(n4963), .B(n4962), .ZN(U3051)
         );
  OAI22_X1 U6140 ( .A1(n4992), .A2(n5049), .B1(n6339), .B2(n5078), .ZN(n4964)
         );
  AOI21_X1 U6141 ( .B1(n6336), .B2(n6241), .A(n4964), .ZN(n4966) );
  NAND2_X1 U6142 ( .A1(n5051), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4965) );
  OAI211_X1 U6143 ( .C1(n5054), .C2(n5179), .A(n4966), .B(n4965), .ZN(U3048)
         );
  OAI22_X1 U6144 ( .A1(n4996), .A2(n5049), .B1(n6335), .B2(n5078), .ZN(n4967)
         );
  AOI21_X1 U6145 ( .B1(n6332), .B2(n6241), .A(n4967), .ZN(n4969) );
  NAND2_X1 U6146 ( .A1(n5051), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4968) );
  OAI211_X1 U6147 ( .C1(n5054), .C2(n5189), .A(n4969), .B(n4968), .ZN(U3047)
         );
  OAI22_X1 U6148 ( .A1(n4988), .A2(n5049), .B1(n6324), .B2(n5078), .ZN(n4970)
         );
  AOI21_X1 U6149 ( .B1(n6381), .B2(n6241), .A(n4970), .ZN(n4972) );
  NAND2_X1 U6150 ( .A1(n5051), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4971) );
  OAI211_X1 U6151 ( .C1(n5054), .C2(n5167), .A(n4972), .B(n4971), .ZN(U3044)
         );
  OAI22_X1 U6152 ( .A1(n5017), .A2(n5049), .B1(n6343), .B2(n5078), .ZN(n4973)
         );
  AOI21_X1 U6153 ( .B1(n6340), .B2(n6241), .A(n4973), .ZN(n4975) );
  NAND2_X1 U6154 ( .A1(n5051), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4974) );
  OAI211_X1 U6155 ( .C1(n5054), .C2(n5159), .A(n4975), .B(n4974), .ZN(U3049)
         );
  INV_X1 U6156 ( .A(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4979) );
  AOI22_X1 U6157 ( .A1(n3193), .A2(n5009), .B1(n6396), .B2(n5019), .ZN(n4976)
         );
  OAI21_X1 U6158 ( .B1(n6399), .B2(n5015), .A(n4976), .ZN(n4977) );
  AOI21_X1 U6159 ( .B1(n6394), .B2(n6388), .A(n4977), .ZN(n4978) );
  OAI21_X1 U6160 ( .B1(n5008), .B2(n4979), .A(n4978), .ZN(U3085) );
  NOR2_X1 U6161 ( .A1(n5067), .A2(n6275), .ZN(n4981) );
  AOI21_X1 U6162 ( .B1(n4981), .B2(n5070), .A(n4980), .ZN(n4985) );
  OR2_X1 U6163 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4982), .ZN(n5065)
         );
  AOI211_X1 U6164 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5065), .A(n6309), .B(
        n4983), .ZN(n4984) );
  NAND2_X1 U6165 ( .A1(n5063), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4991) );
  AOI22_X1 U6166 ( .A1(n4987), .A2(n6313), .B1(n6239), .B2(n4986), .ZN(n5064)
         );
  OAI22_X1 U6167 ( .A1(n4988), .A2(n5065), .B1(n5064), .B2(n5167), .ZN(n4989)
         );
  AOI21_X1 U6168 ( .B1(n6381), .B2(n5067), .A(n4989), .ZN(n4990) );
  OAI211_X1 U6169 ( .C1(n6324), .C2(n5070), .A(n4991), .B(n4990), .ZN(U3020)
         );
  NAND2_X1 U6170 ( .A1(n5063), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4995) );
  OAI22_X1 U6171 ( .A1(n4992), .A2(n5065), .B1(n5064), .B2(n5179), .ZN(n4993)
         );
  AOI21_X1 U6172 ( .B1(n6336), .B2(n5067), .A(n4993), .ZN(n4994) );
  OAI211_X1 U6173 ( .C1(n6339), .C2(n5070), .A(n4995), .B(n4994), .ZN(U3024)
         );
  NAND2_X1 U6174 ( .A1(n5063), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4999) );
  OAI22_X1 U6175 ( .A1(n4996), .A2(n5065), .B1(n5064), .B2(n5189), .ZN(n4997)
         );
  AOI21_X1 U6176 ( .B1(n6332), .B2(n5067), .A(n4997), .ZN(n4998) );
  OAI211_X1 U6177 ( .C1(n6335), .C2(n5070), .A(n4999), .B(n4998), .ZN(U3023)
         );
  NAND2_X1 U6178 ( .A1(n5063), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n5002) );
  INV_X1 U6179 ( .A(n5064), .ZN(n5005) );
  OAI22_X1 U6180 ( .A1(n5017), .A2(n5065), .B1(n6417), .B2(n5003), .ZN(n5000)
         );
  AOI21_X1 U6181 ( .B1(n6414), .B2(n5005), .A(n5000), .ZN(n5001) );
  OAI211_X1 U6182 ( .C1(n6343), .C2(n5070), .A(n5002), .B(n5001), .ZN(U3025)
         );
  NAND2_X1 U6183 ( .A1(n5063), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n5007) );
  OAI22_X1 U6184 ( .A1(n5010), .A2(n5065), .B1(n6378), .B2(n5003), .ZN(n5004)
         );
  AOI21_X1 U6185 ( .B1(n6373), .B2(n5005), .A(n5004), .ZN(n5006) );
  OAI211_X1 U6186 ( .C1(n6355), .C2(n5070), .A(n5007), .B(n5006), .ZN(U3027)
         );
  INV_X1 U6187 ( .A(n5008), .ZN(n5014) );
  NAND2_X1 U6188 ( .A1(n5014), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n5013) );
  INV_X1 U6189 ( .A(n5009), .ZN(n5016) );
  OAI22_X1 U6190 ( .A1(n5010), .A2(n5016), .B1(n6378), .B2(n5015), .ZN(n5011)
         );
  AOI21_X1 U6191 ( .B1(n6373), .B2(n5019), .A(n5011), .ZN(n5012) );
  OAI211_X1 U6192 ( .C1(n5022), .C2(n6355), .A(n5013), .B(n5012), .ZN(U3091)
         );
  NAND2_X1 U6193 ( .A1(n5014), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n5021) );
  OAI22_X1 U6194 ( .A1(n5017), .A2(n5016), .B1(n6417), .B2(n5015), .ZN(n5018)
         );
  AOI21_X1 U6195 ( .B1(n6414), .B2(n5019), .A(n5018), .ZN(n5020) );
  OAI211_X1 U6196 ( .C1(n5022), .C2(n6343), .A(n5021), .B(n5020), .ZN(U3089)
         );
  INV_X1 U6197 ( .A(n6423), .ZN(n5183) );
  INV_X1 U6198 ( .A(n6421), .ZN(n5045) );
  OAI22_X1 U6199 ( .A1(n5045), .A2(n5049), .B1(n6347), .B2(n5078), .ZN(n5023)
         );
  AOI21_X1 U6200 ( .B1(n6344), .B2(n6241), .A(n5023), .ZN(n5025) );
  NAND2_X1 U6201 ( .A1(n5051), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n5024) );
  OAI211_X1 U6202 ( .C1(n5054), .C2(n5183), .A(n5025), .B(n5024), .ZN(U3050)
         );
  INV_X1 U6203 ( .A(n6402), .ZN(n5175) );
  INV_X1 U6204 ( .A(n6401), .ZN(n5041) );
  OAI22_X1 U6205 ( .A1(n5041), .A2(n5049), .B1(n6331), .B2(n5078), .ZN(n5026)
         );
  AOI21_X1 U6206 ( .B1(n6328), .B2(n6241), .A(n5026), .ZN(n5028) );
  NAND2_X1 U6207 ( .A1(n5051), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n5027) );
  OAI211_X1 U6208 ( .C1(n5054), .C2(n5175), .A(n5028), .B(n5027), .ZN(U3046)
         );
  NAND2_X1 U6209 ( .A1(n5063), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n5031) );
  OAI22_X1 U6210 ( .A1(n5045), .A2(n5065), .B1(n5064), .B2(n5183), .ZN(n5029)
         );
  AOI21_X1 U6211 ( .B1(n6344), .B2(n5067), .A(n5029), .ZN(n5030) );
  OAI211_X1 U6212 ( .C1(n6347), .C2(n5070), .A(n5031), .B(n5030), .ZN(U3026)
         );
  NAND2_X1 U6213 ( .A1(n5063), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n5034) );
  OAI22_X1 U6214 ( .A1(n5041), .A2(n5065), .B1(n5064), .B2(n5175), .ZN(n5032)
         );
  AOI21_X1 U6215 ( .B1(n6328), .B2(n5067), .A(n5032), .ZN(n5033) );
  OAI211_X1 U6216 ( .C1(n6331), .C2(n5070), .A(n5034), .B(n5033), .ZN(U3022)
         );
  NAND2_X1 U6217 ( .A1(n5055), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n5037)
         );
  OAI22_X1 U6218 ( .A1(n5041), .A2(n5057), .B1(n5056), .B2(n5175), .ZN(n5035)
         );
  AOI21_X1 U6219 ( .B1(n6400), .B2(n5059), .A(n5035), .ZN(n5036) );
  OAI211_X1 U6220 ( .C1(n5062), .C2(n6405), .A(n5037), .B(n5036), .ZN(U3118)
         );
  NAND2_X1 U6221 ( .A1(n5055), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n5040)
         );
  OAI22_X1 U6222 ( .A1(n5045), .A2(n5057), .B1(n5056), .B2(n5183), .ZN(n5038)
         );
  AOI21_X1 U6223 ( .B1(n6418), .B2(n5059), .A(n5038), .ZN(n5039) );
  OAI211_X1 U6224 ( .C1(n5062), .C2(n6428), .A(n5040), .B(n5039), .ZN(U3122)
         );
  NAND2_X1 U6225 ( .A1(n5071), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n5044) );
  OAI22_X1 U6226 ( .A1(n5041), .A2(n5073), .B1(n5072), .B2(n5175), .ZN(n5042)
         );
  AOI21_X1 U6227 ( .B1(n6400), .B2(n6302), .A(n5042), .ZN(n5043) );
  OAI211_X1 U6228 ( .C1(n5078), .C2(n6405), .A(n5044), .B(n5043), .ZN(U3054)
         );
  NAND2_X1 U6229 ( .A1(n5071), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n5048) );
  OAI22_X1 U6230 ( .A1(n5045), .A2(n5073), .B1(n5072), .B2(n5183), .ZN(n5046)
         );
  AOI21_X1 U6231 ( .B1(n6418), .B2(n6302), .A(n5046), .ZN(n5047) );
  OAI211_X1 U6232 ( .C1(n5078), .C2(n6428), .A(n5048), .B(n5047), .ZN(U3058)
         );
  INV_X1 U6233 ( .A(n6396), .ZN(n5171) );
  OAI22_X1 U6235 ( .A1(n6974), .A2(n5049), .B1(n6327), .B2(n5078), .ZN(n5050)
         );
  AOI21_X1 U6236 ( .B1(n6387), .B2(n6241), .A(n5050), .ZN(n5053) );
  NAND2_X1 U6237 ( .A1(n5051), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n5052) );
  OAI211_X1 U6238 ( .C1(n5054), .C2(n5171), .A(n5053), .B(n5052), .ZN(U3045)
         );
  NAND2_X1 U6239 ( .A1(n5055), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n5061)
         );
  OAI22_X1 U6240 ( .A1(n6974), .A2(n5057), .B1(n5056), .B2(n5171), .ZN(n5058)
         );
  AOI21_X1 U6241 ( .B1(n6394), .B2(n5059), .A(n5058), .ZN(n5060) );
  OAI211_X1 U6242 ( .C1(n5062), .C2(n6399), .A(n5061), .B(n5060), .ZN(U3117)
         );
  NAND2_X1 U6243 ( .A1(n5063), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n5069) );
  OAI22_X1 U6244 ( .A1(n6974), .A2(n5065), .B1(n5064), .B2(n5171), .ZN(n5066)
         );
  AOI21_X1 U6245 ( .B1(n6387), .B2(n5067), .A(n5066), .ZN(n5068) );
  OAI211_X1 U6246 ( .C1(n6327), .C2(n5070), .A(n5069), .B(n5068), .ZN(U3021)
         );
  NAND2_X1 U6247 ( .A1(n5071), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n5077) );
  OAI22_X1 U6248 ( .A1(n6974), .A2(n5073), .B1(n5072), .B2(n5171), .ZN(n5075)
         );
  AOI21_X1 U6249 ( .B1(n6394), .B2(n6302), .A(n5075), .ZN(n5076) );
  OAI211_X1 U6250 ( .C1(n5078), .C2(n6399), .A(n5077), .B(n5076), .ZN(U3053)
         );
  OAI21_X1 U6251 ( .B1(n5080), .B2(n3524), .A(n5967), .ZN(n5992) );
  INV_X1 U6252 ( .A(n5992), .ZN(n5115) );
  INV_X1 U6253 ( .A(n6156), .ZN(n5088) );
  OR2_X1 U6254 ( .A1(n5976), .A2(REIP_REG_1__SCAN_IN), .ZN(n5090) );
  AND2_X1 U6255 ( .A1(n5090), .A2(REIP_REG_2__SCAN_IN), .ZN(n5079) );
  AND2_X1 U6256 ( .A1(n5953), .A2(n5079), .ZN(n5987) );
  AOI21_X1 U6257 ( .B1(n5986), .B2(REIP_REG_1__SCAN_IN), .A(
        REIP_REG_2__SCAN_IN), .ZN(n5086) );
  NOR2_X1 U6258 ( .A1(n5081), .A2(n5080), .ZN(n5984) );
  AOI22_X1 U6259 ( .A1(n5982), .A2(EBX_REG_2__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n5983), .ZN(n5082) );
  OAI21_X1 U6260 ( .B1(n6209), .B2(n5969), .A(n5082), .ZN(n5083) );
  AOI21_X1 U6261 ( .B1(n5084), .B2(n5984), .A(n5083), .ZN(n5085) );
  OAI21_X1 U6262 ( .B1(n5987), .B2(n5086), .A(n5085), .ZN(n5087) );
  AOI21_X1 U6263 ( .B1(n5964), .B2(n5088), .A(n5087), .ZN(n5089) );
  OAI21_X1 U6264 ( .B1(n5115), .B2(n6148), .A(n5089), .ZN(U2825) );
  INV_X1 U6265 ( .A(n5984), .ZN(n5107) );
  AOI22_X1 U6266 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n5983), .B1(n5103), 
        .B2(REIP_REG_1__SCAN_IN), .ZN(n5091) );
  OAI211_X1 U6267 ( .C1(n5961), .C2(n3275), .A(n5091), .B(n5090), .ZN(n5092)
         );
  AOI21_X1 U6268 ( .B1(n5093), .B2(n5981), .A(n5092), .ZN(n5094) );
  OAI21_X1 U6269 ( .B1(n5644), .B2(n5107), .A(n5094), .ZN(n5095) );
  AOI21_X1 U6270 ( .B1(n5964), .B2(n5096), .A(n5095), .ZN(n5097) );
  OAI21_X1 U6271 ( .B1(n5115), .B2(n5098), .A(n5097), .ZN(U2826) );
  NOR3_X1 U6272 ( .A1(n5976), .A2(n5985), .A3(REIP_REG_4__SCAN_IN), .ZN(n5099)
         );
  AOI211_X1 U6273 ( .C1(EBX_REG_4__SCAN_IN), .C2(n5982), .A(n5973), .B(n5099), 
        .ZN(n5101) );
  NAND2_X1 U6274 ( .A1(n6196), .A2(n5981), .ZN(n5100) );
  OAI211_X1 U6275 ( .C1(n5102), .C2(n5107), .A(n5101), .B(n5100), .ZN(n5105)
         );
  OAI21_X1 U6276 ( .B1(n5103), .B2(n5985), .A(n5894), .ZN(n5995) );
  OAI22_X1 U6277 ( .A1(n5995), .A2(n6719), .B1(n6897), .B2(n5970), .ZN(n5104)
         );
  AOI211_X1 U6278 ( .C1(n5964), .C2(n6133), .A(n5105), .B(n5104), .ZN(n5106)
         );
  OAI21_X1 U6279 ( .B1(n5115), .B2(n6137), .A(n5106), .ZN(U2823) );
  NOR2_X1 U6280 ( .A1(n6267), .A2(n5107), .ZN(n5111) );
  OAI22_X1 U6281 ( .A1(n5961), .A2(n5109), .B1(n5108), .B2(n5969), .ZN(n5110)
         );
  AOI211_X1 U6282 ( .C1(n5894), .C2(REIP_REG_0__SCAN_IN), .A(n5111), .B(n5110), 
        .ZN(n5113) );
  OAI21_X1 U6283 ( .B1(n5964), .B2(n5983), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n5112) );
  OAI211_X1 U6284 ( .C1(n5115), .C2(n5114), .A(n5113), .B(n5112), .ZN(U2827)
         );
  XNOR2_X1 U6285 ( .A(n5117), .B(n5116), .ZN(n6105) );
  AOI22_X1 U6286 ( .A1(n5479), .A2(DATAI_8_), .B1(n6005), .B2(
        EAX_REG_8__SCAN_IN), .ZN(n5118) );
  OAI21_X1 U6287 ( .B1(n6970), .B2(n6105), .A(n5118), .ZN(U2883) );
  XOR2_X1 U6288 ( .A(n5120), .B(n5119), .Z(n6110) );
  INV_X1 U6289 ( .A(n6110), .ZN(n5134) );
  AOI22_X1 U6290 ( .A1(n5479), .A2(DATAI_7_), .B1(n6005), .B2(
        EAX_REG_7__SCAN_IN), .ZN(n5121) );
  OAI21_X1 U6291 ( .B1(n5134), .B2(n6970), .A(n5121), .ZN(U2884) );
  OAI21_X1 U6292 ( .B1(n5124), .B2(n5123), .A(n5122), .ZN(n6097) );
  AOI22_X1 U6293 ( .A1(n5479), .A2(DATAI_9_), .B1(n6005), .B2(
        EAX_REG_9__SCAN_IN), .ZN(n5125) );
  OAI21_X1 U6294 ( .B1(n6097), .B2(n6970), .A(n5125), .ZN(U2882) );
  AOI21_X1 U6295 ( .B1(n5126), .B2(n5137), .A(n5200), .ZN(n6166) );
  AOI22_X1 U6296 ( .A1(n6166), .A2(n5445), .B1(n5462), .B2(EBX_REG_9__SCAN_IN), 
        .ZN(n5127) );
  OAI21_X1 U6297 ( .B1(n6097), .B2(n3195), .A(n5127), .ZN(U2850) );
  INV_X1 U6298 ( .A(n5128), .ZN(n5129) );
  NAND2_X1 U6299 ( .A1(n5130), .A2(n5129), .ZN(n5132) );
  INV_X1 U6300 ( .A(n5131), .ZN(n5139) );
  AOI21_X1 U6301 ( .B1(n5133), .B2(n5132), .A(n5139), .ZN(n6183) );
  INV_X1 U6302 ( .A(n6183), .ZN(n5135) );
  INV_X1 U6303 ( .A(EBX_REG_7__SCAN_IN), .ZN(n6743) );
  OAI222_X1 U6304 ( .A1(n5135), .A2(n5466), .B1(n5453), .B2(n6743), .C1(n3195), 
        .C2(n5134), .ZN(U2852) );
  INV_X1 U6305 ( .A(n5136), .ZN(n5138) );
  OAI21_X1 U6306 ( .B1(n5139), .B2(n5138), .A(n5137), .ZN(n6176) );
  INV_X1 U6307 ( .A(n6105), .ZN(n5140) );
  AOI22_X1 U6308 ( .A1(n6975), .A2(n5140), .B1(n5462), .B2(EBX_REG_8__SCAN_IN), 
        .ZN(n5141) );
  OAI21_X1 U6309 ( .B1(n6176), .B2(n5466), .A(n5141), .ZN(U2851) );
  AOI21_X1 U6310 ( .B1(n5122), .B2(n5143), .A(n5193), .ZN(n5925) );
  INV_X1 U6311 ( .A(n5925), .ZN(n5203) );
  AOI22_X1 U6312 ( .A1(n5479), .A2(DATAI_10_), .B1(n6005), .B2(
        EAX_REG_10__SCAN_IN), .ZN(n5144) );
  OAI21_X1 U6313 ( .B1(n5203), .B2(n6970), .A(n5144), .ZN(U2881) );
  NAND2_X1 U6314 ( .A1(n5148), .A2(n6427), .ZN(n5145) );
  AOI21_X1 U6315 ( .B1(n5145), .B2(STATEBS16_REG_SCAN_IN), .A(n6275), .ZN(
        n5153) );
  NOR3_X1 U6316 ( .A1(n6318), .A2(n6441), .A3(n5146), .ZN(n5147) );
  NOR2_X1 U6317 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5149), .ZN(n5185)
         );
  NOR2_X1 U6318 ( .A1(n6309), .A2(n6320), .ZN(n6244) );
  INV_X1 U6319 ( .A(n5150), .ZN(n5152) );
  INV_X1 U6320 ( .A(n5185), .ZN(n5151) );
  AOI22_X1 U6321 ( .A1(n5153), .A2(n5152), .B1(STATE2_REG_3__SCAN_IN), .B2(
        n5151), .ZN(n5154) );
  OAI211_X1 U6322 ( .C1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n5155), .A(n6244), .B(n5154), .ZN(n5184) );
  AOI22_X1 U6323 ( .A1(n6413), .A2(n5185), .B1(INSTQUEUE_REG_10__5__SCAN_IN), 
        .B2(n5184), .ZN(n5156) );
  OAI21_X1 U6324 ( .B1(n6343), .B2(n6427), .A(n5156), .ZN(n5157) );
  AOI21_X1 U6325 ( .B1(n6340), .B2(n6389), .A(n5157), .ZN(n5158) );
  OAI21_X1 U6326 ( .B1(n5190), .B2(n5159), .A(n5158), .ZN(U3105) );
  AOI22_X1 U6327 ( .A1(n6369), .A2(n5185), .B1(INSTQUEUE_REG_10__7__SCAN_IN), 
        .B2(n5184), .ZN(n5160) );
  OAI21_X1 U6328 ( .B1(n6355), .B2(n6427), .A(n5160), .ZN(n5161) );
  AOI21_X1 U6329 ( .B1(n6351), .B2(n6389), .A(n5161), .ZN(n5162) );
  OAI21_X1 U6330 ( .B1(n5190), .B2(n5163), .A(n5162), .ZN(U3107) );
  AOI22_X1 U6331 ( .A1(n6380), .A2(n5185), .B1(INSTQUEUE_REG_10__0__SCAN_IN), 
        .B2(n5184), .ZN(n5164) );
  OAI21_X1 U6332 ( .B1(n6324), .B2(n6427), .A(n5164), .ZN(n5165) );
  AOI21_X1 U6333 ( .B1(n6381), .B2(n6389), .A(n5165), .ZN(n5166) );
  OAI21_X1 U6334 ( .B1(n5190), .B2(n5167), .A(n5166), .ZN(U3100) );
  AOI22_X1 U6335 ( .A1(n3193), .A2(n5185), .B1(INSTQUEUE_REG_10__1__SCAN_IN), 
        .B2(n5184), .ZN(n5168) );
  OAI21_X1 U6336 ( .B1(n6327), .B2(n6427), .A(n5168), .ZN(n5169) );
  AOI21_X1 U6337 ( .B1(n6387), .B2(n6389), .A(n5169), .ZN(n5170) );
  OAI21_X1 U6338 ( .B1(n5190), .B2(n5171), .A(n5170), .ZN(U3101) );
  AOI22_X1 U6339 ( .A1(n6401), .A2(n5185), .B1(INSTQUEUE_REG_10__2__SCAN_IN), 
        .B2(n5184), .ZN(n5172) );
  OAI21_X1 U6340 ( .B1(n6331), .B2(n6427), .A(n5172), .ZN(n5173) );
  AOI21_X1 U6341 ( .B1(n6328), .B2(n6389), .A(n5173), .ZN(n5174) );
  OAI21_X1 U6342 ( .B1(n5190), .B2(n5175), .A(n5174), .ZN(U3102) );
  AOI22_X1 U6343 ( .A1(n6358), .A2(n5185), .B1(INSTQUEUE_REG_10__4__SCAN_IN), 
        .B2(n5184), .ZN(n5176) );
  OAI21_X1 U6344 ( .B1(n6339), .B2(n6427), .A(n5176), .ZN(n5177) );
  AOI21_X1 U6345 ( .B1(n6336), .B2(n6389), .A(n5177), .ZN(n5178) );
  OAI21_X1 U6346 ( .B1(n5190), .B2(n5179), .A(n5178), .ZN(U3104) );
  AOI22_X1 U6347 ( .A1(n6421), .A2(n5185), .B1(INSTQUEUE_REG_10__6__SCAN_IN), 
        .B2(n5184), .ZN(n5180) );
  OAI21_X1 U6348 ( .B1(n6347), .B2(n6427), .A(n5180), .ZN(n5181) );
  AOI21_X1 U6349 ( .B1(n6344), .B2(n6389), .A(n5181), .ZN(n5182) );
  OAI21_X1 U6350 ( .B1(n5190), .B2(n5183), .A(n5182), .ZN(U3106) );
  AOI22_X1 U6351 ( .A1(n6407), .A2(n5185), .B1(INSTQUEUE_REG_10__3__SCAN_IN), 
        .B2(n5184), .ZN(n5186) );
  OAI21_X1 U6352 ( .B1(n6335), .B2(n6427), .A(n5186), .ZN(n5187) );
  AOI21_X1 U6353 ( .B1(n6332), .B2(n6389), .A(n5187), .ZN(n5188) );
  OAI21_X1 U6354 ( .B1(n5190), .B2(n5189), .A(n5188), .ZN(U3103) );
  OAI21_X1 U6355 ( .B1(n5193), .B2(n5192), .A(n5191), .ZN(n6089) );
  AOI22_X1 U6356 ( .A1(n5479), .A2(DATAI_11_), .B1(n6005), .B2(
        EAX_REG_11__SCAN_IN), .ZN(n5194) );
  OAI21_X1 U6357 ( .B1(n6089), .B2(n6970), .A(n5194), .ZN(U2880) );
  OAI21_X1 U6358 ( .B1(n5202), .B2(n5196), .A(n5195), .ZN(n5197) );
  INV_X1 U6359 ( .A(n5197), .ZN(n6158) );
  AOI22_X1 U6360 ( .A1(n6158), .A2(n5445), .B1(n5462), .B2(EBX_REG_11__SCAN_IN), .ZN(n5198) );
  OAI21_X1 U6361 ( .B1(n6089), .B2(n3195), .A(n5198), .ZN(U2848) );
  NOR2_X1 U6362 ( .A1(n5200), .A2(n5199), .ZN(n5201) );
  OR2_X1 U6363 ( .A1(n5202), .A2(n5201), .ZN(n5922) );
  INV_X1 U6364 ( .A(EBX_REG_10__SCAN_IN), .ZN(n5923) );
  OAI222_X1 U6365 ( .A1(n5922), .A2(n5466), .B1(n5453), .B2(n5923), .C1(n3195), 
        .C2(n5203), .ZN(U2849) );
  NAND2_X1 U6366 ( .A1(n6082), .A2(n5204), .ZN(n5206) );
  XOR2_X1 U6367 ( .A(n5206), .B(n5205), .Z(n5220) );
  INV_X1 U6368 ( .A(n5210), .ZN(n6173) );
  OAI22_X1 U6369 ( .A1(n5578), .A2(n5208), .B1(n5573), .B2(n5207), .ZN(n6184)
         );
  INV_X1 U6370 ( .A(n6184), .ZN(n6182) );
  OAI21_X1 U6371 ( .B1(n6173), .B2(n5289), .A(n6182), .ZN(n6165) );
  INV_X1 U6372 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6501) );
  OAI22_X1 U6373 ( .A1(n5922), .A2(n6177), .B1(n6501), .B2(n6175), .ZN(n5214)
         );
  INV_X1 U6374 ( .A(n5609), .ZN(n6217) );
  AOI21_X1 U6375 ( .B1(n6213), .B2(n6217), .A(n6212), .ZN(n6198) );
  NOR2_X1 U6376 ( .A1(n6198), .A2(n5209), .ZN(n6191) );
  NAND2_X1 U6377 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n6191), .ZN(n6188)
         );
  NOR2_X1 U6378 ( .A1(n5210), .A2(n6188), .ZN(n6167) );
  OAI211_X1 U6379 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A(n6167), .B(n5211), .ZN(n5212) );
  INV_X1 U6380 ( .A(n5212), .ZN(n5213) );
  AOI211_X1 U6381 ( .C1(n6165), .C2(INSTADDRPOINTER_REG_10__SCAN_IN), .A(n5214), .B(n5213), .ZN(n5215) );
  OAI21_X1 U6382 ( .B1(n5220), .B2(n5815), .A(n5215), .ZN(U3008) );
  NAND2_X1 U6383 ( .A1(n5925), .A2(n6124), .ZN(n5219) );
  OAI22_X1 U6384 ( .A1(n5791), .A2(n5216), .B1(n6175), .B2(n6501), .ZN(n5217)
         );
  AOI21_X1 U6385 ( .B1(n6134), .B2(n5926), .A(n5217), .ZN(n5218) );
  OAI211_X1 U6386 ( .C1(n5220), .C2(n5831), .A(n5219), .B(n5218), .ZN(U2976)
         );
  AOI21_X1 U6387 ( .B1(n5191), .B2(n5222), .A(n5221), .ZN(n5908) );
  INV_X1 U6388 ( .A(n5908), .ZN(n5227) );
  AOI22_X1 U6389 ( .A1(n5479), .A2(DATAI_12_), .B1(n6005), .B2(
        EAX_REG_12__SCAN_IN), .ZN(n5223) );
  OAI21_X1 U6390 ( .B1(n5227), .B2(n6970), .A(n5223), .ZN(U2879) );
  INV_X1 U6391 ( .A(n5456), .ZN(n5224) );
  AOI21_X1 U6392 ( .B1(n5225), .B2(n5195), .A(n5224), .ZN(n5907) );
  AOI22_X1 U6393 ( .A1(n5907), .A2(n5445), .B1(n5462), .B2(EBX_REG_12__SCAN_IN), .ZN(n5226) );
  OAI21_X1 U6394 ( .B1(n5227), .B2(n3195), .A(n5226), .ZN(U2847) );
  INV_X1 U6395 ( .A(n5229), .ZN(n5230) );
  NOR2_X1 U6396 ( .A1(n5231), .A2(n5230), .ZN(n5232) );
  XNOR2_X1 U6397 ( .A(n5228), .B(n5232), .ZN(n5247) );
  NAND2_X1 U6398 ( .A1(n6134), .A2(n5909), .ZN(n5233) );
  NAND2_X1 U6399 ( .A1(n6210), .A2(REIP_REG_12__SCAN_IN), .ZN(n5240) );
  OAI211_X1 U6400 ( .C1(n5234), .C2(n5791), .A(n5233), .B(n5240), .ZN(n5235)
         );
  AOI21_X1 U6401 ( .B1(n5908), .B2(n4403), .A(n5235), .ZN(n5236) );
  OAI21_X1 U6402 ( .B1(n5247), .B2(n5831), .A(n5236), .ZN(U2974) );
  AOI22_X1 U6403 ( .A1(n5239), .A2(n5238), .B1(n5237), .B2(n5629), .ZN(n6164)
         );
  INV_X1 U6404 ( .A(n6164), .ZN(n5245) );
  INV_X1 U6405 ( .A(n5907), .ZN(n5241) );
  OAI21_X1 U6406 ( .B1(n5241), .B2(n6177), .A(n5240), .ZN(n5244) );
  INV_X1 U6407 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6163) );
  INV_X1 U6408 ( .A(n6159), .ZN(n5823) );
  INV_X1 U6409 ( .A(n5631), .ZN(n5817) );
  AOI211_X1 U6410 ( .C1(n6163), .C2(n5242), .A(n5823), .B(n5817), .ZN(n5243)
         );
  AOI211_X1 U6411 ( .C1(INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n5245), .A(n5244), .B(n5243), .ZN(n5246) );
  OAI21_X1 U6412 ( .B1(n5247), .B2(n5815), .A(n5246), .ZN(U3006) );
  OR2_X2 U6413 ( .A1(n5589), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5590)
         );
  INV_X1 U6414 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5595) );
  OAI21_X1 U6415 ( .B1(n5248), .B2(n5595), .A(n5604), .ZN(n5249) );
  INV_X1 U6416 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5250) );
  XNOR2_X1 U6417 ( .A(n5604), .B(n5250), .ZN(n5517) );
  OAI22_X1 U6418 ( .A1(n5496), .A2(n5517), .B1(n5604), .B2(n5250), .ZN(n5512)
         );
  INV_X1 U6419 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5251) );
  XNOR2_X1 U6420 ( .A(n5604), .B(n5251), .ZN(n5513) );
  NOR2_X1 U6421 ( .A1(n5604), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5505)
         );
  NAND2_X1 U6422 ( .A1(n5511), .A2(n5505), .ZN(n5498) );
  OAI21_X1 U6423 ( .B1(n5592), .B2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n5252), 
        .ZN(n5504) );
  NAND3_X1 U6424 ( .A1(n5604), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5253) );
  XNOR2_X1 U6425 ( .A(n5254), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5273)
         );
  NAND2_X1 U6426 ( .A1(n5255), .A2(n5256), .ZN(n5257) );
  NAND2_X1 U6427 ( .A1(n5392), .A2(n5257), .ZN(n5696) );
  INV_X1 U6428 ( .A(n5696), .ZN(n5262) );
  NAND2_X1 U6429 ( .A1(n6210), .A2(REIP_REG_24__SCAN_IN), .ZN(n5264) );
  INV_X1 U6430 ( .A(n5264), .ZN(n5261) );
  INV_X1 U6431 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5259) );
  NAND2_X1 U6432 ( .A1(n5560), .A2(n5497), .ZN(n5550) );
  AOI211_X1 U6433 ( .C1(n5259), .C2(n5550), .A(n5258), .B(n5808), .ZN(n5260)
         );
  AOI211_X1 U6434 ( .C1(n6227), .C2(n5262), .A(n5261), .B(n5260), .ZN(n5263)
         );
  OAI21_X1 U6435 ( .B1(n5273), .B2(n5815), .A(n5263), .ZN(U2994) );
  OAI21_X1 U6436 ( .B1(n5791), .B2(n5265), .A(n5264), .ZN(n5271) );
  INV_X1 U6437 ( .A(n5267), .ZN(n5269) );
  OR2_X2 U6438 ( .A1(n5268), .A2(n5267), .ZN(n5388) );
  NOR2_X1 U6439 ( .A1(n5692), .A2(n6138), .ZN(n5270) );
  AOI211_X1 U6440 ( .C1(n6134), .C2(n5689), .A(n5271), .B(n5270), .ZN(n5272)
         );
  OAI21_X1 U6441 ( .B1(n5273), .B2(n5831), .A(n5272), .ZN(U2962) );
  NOR3_X1 U6442 ( .A1(n6005), .A2(n5468), .A3(n3203), .ZN(n5274) );
  AOI22_X1 U6443 ( .A1(n6006), .A2(DATAI_8_), .B1(EAX_REG_24__SCAN_IN), .B2(
        n6005), .ZN(n5277) );
  NAND2_X1 U6444 ( .A1(n5996), .A2(DATAI_24_), .ZN(n5276) );
  OAI211_X1 U6445 ( .C1(n5692), .C2(n6970), .A(n5277), .B(n5276), .ZN(U2867)
         );
  INV_X1 U6446 ( .A(EBX_REG_24__SCAN_IN), .ZN(n5278) );
  OAI222_X1 U6447 ( .A1(n5696), .A2(n5466), .B1(n5453), .B2(n5278), .C1(n3195), 
        .C2(n5692), .ZN(U2835) );
  OR2_X2 U6448 ( .A1(n5388), .A2(n5389), .ZN(n5386) );
  AOI21_X2 U6449 ( .B1(n5280), .B2(n5386), .A(n5378), .ZN(n5281) );
  AOI22_X1 U6450 ( .A1(n6006), .A2(DATAI_10_), .B1(EAX_REG_26__SCAN_IN), .B2(
        n6005), .ZN(n5283) );
  NAND2_X1 U6451 ( .A1(n5996), .A2(DATAI_26_), .ZN(n5282) );
  OAI211_X1 U6452 ( .C1(n5768), .C2(n6970), .A(n5283), .B(n5282), .ZN(U2865)
         );
  OAI22_X1 U6453 ( .A1(n5673), .A2(n5466), .B1(n5679), .B2(n5453), .ZN(n5284)
         );
  INV_X1 U6454 ( .A(n5284), .ZN(n5285) );
  OAI21_X1 U6455 ( .B1(n5768), .B2(n3195), .A(n5285), .ZN(U2833) );
  XNOR2_X1 U6456 ( .A(n5604), .B(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5287)
         );
  XNOR2_X1 U6457 ( .A(n3201), .B(n5287), .ZN(n5308) );
  INV_X1 U6458 ( .A(n5617), .ZN(n5288) );
  OAI21_X1 U6459 ( .B1(n5289), .B2(n5288), .A(n6164), .ZN(n5615) );
  INV_X1 U6460 ( .A(n5290), .ZN(n5294) );
  INV_X1 U6461 ( .A(n5291), .ZN(n5449) );
  INV_X1 U6462 ( .A(n5292), .ZN(n5293) );
  AOI21_X1 U6463 ( .B1(n5294), .B2(n5449), .A(n5293), .ZN(n5881) );
  INV_X1 U6464 ( .A(n5881), .ZN(n5297) );
  NOR2_X1 U6465 ( .A1(n5823), .A2(n5617), .ZN(n5295) );
  NAND2_X1 U6466 ( .A1(n5295), .A2(n5618), .ZN(n5296) );
  NAND2_X1 U6467 ( .A1(n6210), .A2(REIP_REG_15__SCAN_IN), .ZN(n5303) );
  OAI211_X1 U6468 ( .C1(n6177), .C2(n5297), .A(n5296), .B(n5303), .ZN(n5298)
         );
  AOI21_X1 U6469 ( .B1(n5615), .B2(INSTADDRPOINTER_REG_15__SCAN_IN), .A(n5298), 
        .ZN(n5299) );
  OAI21_X1 U6470 ( .B1(n5308), .B2(n5815), .A(n5299), .ZN(U3003) );
  AOI21_X1 U6471 ( .B1(n5300), .B2(n5302), .A(n5301), .ZN(n5880) );
  NAND2_X1 U6472 ( .A1(n6134), .A2(n5882), .ZN(n5304) );
  OAI211_X1 U6473 ( .C1(n5791), .C2(n5305), .A(n5304), .B(n5303), .ZN(n5306)
         );
  AOI21_X1 U6474 ( .B1(n5880), .B2(n6124), .A(n5306), .ZN(n5307) );
  OAI21_X1 U6475 ( .B1(n5308), .B2(n5831), .A(n5307), .ZN(U2971) );
  AOI21_X1 U6476 ( .B1(INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n5310), .A(n5309), 
        .ZN(n5311) );
  INV_X1 U6477 ( .A(n5312), .ZN(n5316) );
  NOR2_X1 U6478 ( .A1(n6175), .A2(n6829), .ZN(n5322) );
  NOR4_X1 U6479 ( .A1(n5522), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .A3(n5314), 
        .A4(n5313), .ZN(n5315) );
  AOI211_X1 U6480 ( .C1(n5316), .C2(INSTADDRPOINTER_REG_31__SCAN_IN), .A(n5322), .B(n5315), .ZN(n5318) );
  NAND2_X1 U6481 ( .A1(n5367), .A2(n6227), .ZN(n5317) );
  OAI211_X1 U6482 ( .C1(n3222), .C2(n5815), .A(n5318), .B(n5317), .ZN(U2987)
         );
  NAND2_X1 U6483 ( .A1(n5319), .A2(n4403), .ZN(n5324) );
  NOR2_X1 U6484 ( .A1(n5320), .A2(n6157), .ZN(n5321) );
  AOI211_X1 U6485 ( .C1(n6147), .C2(PHYADDRPOINTER_REG_31__SCAN_IN), .A(n5322), 
        .B(n5321), .ZN(n5323) );
  OAI211_X1 U6486 ( .C1(n3222), .C2(n5831), .A(n5324), .B(n5323), .ZN(U2955)
         );
  AOI21_X1 U6487 ( .B1(n6431), .B2(n6550), .A(n6553), .ZN(n5330) );
  OAI22_X1 U6488 ( .A1(n6267), .A2(n5326), .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n5325), .ZN(n6429) );
  OAI22_X1 U6489 ( .A1(n6736), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n5327), .ZN(n5328) );
  AOI21_X1 U6490 ( .B1(n6429), .B2(n6550), .A(n5328), .ZN(n5329) );
  OAI22_X1 U6491 ( .A1(n5330), .A2(n3232), .B1(n6553), .B2(n5329), .ZN(U3461)
         );
  INV_X1 U6492 ( .A(n5331), .ZN(n5337) );
  NAND3_X1 U6493 ( .A1(n5332), .A2(n6548), .A3(n6876), .ZN(n5333) );
  OAI21_X1 U6494 ( .B1(n5335), .B2(n5334), .A(n5333), .ZN(n5336) );
  AOI21_X1 U6495 ( .B1(n5337), .B2(n6550), .A(n5336), .ZN(n5340) );
  AOI21_X1 U6496 ( .B1(n6548), .B2(n5338), .A(n6553), .ZN(n5339) );
  OAI22_X1 U6497 ( .A1(n5340), .A2(n6553), .B1(n5339), .B2(n6876), .ZN(U3459)
         );
  INV_X1 U6498 ( .A(n5489), .ZN(n5343) );
  XNOR2_X1 U6499 ( .A(n5344), .B(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5521)
         );
  NAND2_X1 U6500 ( .A1(n6210), .A2(REIP_REG_29__SCAN_IN), .ZN(n5525) );
  NAND2_X1 U6501 ( .A1(n6147), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5345)
         );
  OAI211_X1 U6502 ( .C1(n5346), .C2(n6157), .A(n5525), .B(n5345), .ZN(n5347)
         );
  AOI21_X1 U6503 ( .B1(n5521), .B2(n6152), .A(n5347), .ZN(n5348) );
  OAI21_X1 U6504 ( .B1(n5341), .B2(n6138), .A(n5348), .ZN(U2957) );
  OAI22_X1 U6505 ( .A1(n5526), .A2(n5466), .B1(n5349), .B2(n5453), .ZN(n5350)
         );
  INV_X1 U6506 ( .A(n5350), .ZN(n5351) );
  OAI21_X1 U6507 ( .B1(n5341), .B2(n3195), .A(n5351), .ZN(U2830) );
  INV_X1 U6508 ( .A(n5363), .ZN(n5352) );
  OR2_X1 U6509 ( .A1(n5353), .A2(n5352), .ZN(n5356) );
  AOI22_X1 U6510 ( .A1(n5364), .A2(n5356), .B1(n5355), .B2(n3528), .ZN(n5360)
         );
  INV_X1 U6511 ( .A(n5364), .ZN(n5358) );
  NAND2_X1 U6512 ( .A1(n5358), .A2(n5357), .ZN(n5359) );
  AND2_X1 U6513 ( .A1(n5360), .A2(n5359), .ZN(n6445) );
  INV_X1 U6514 ( .A(n6445), .ZN(n5366) );
  NAND2_X1 U6515 ( .A1(n5361), .A2(n3528), .ZN(n5362) );
  AOI22_X1 U6516 ( .A1(n5364), .A2(n3524), .B1(n5363), .B2(n5362), .ZN(n5824)
         );
  NAND3_X1 U6517 ( .A1(n3524), .A2(n3196), .A3(n6481), .ZN(n5365) );
  NAND2_X1 U6518 ( .A1(n5365), .A2(n4324), .ZN(n6563) );
  NAND2_X1 U6519 ( .A1(n5824), .A2(n6563), .ZN(n6447) );
  AND2_X1 U6520 ( .A1(n6447), .A2(n6463), .ZN(n5833) );
  MUX2_X1 U6521 ( .A(MORE_REG_SCAN_IN), .B(n5366), .S(n5833), .Z(U3471) );
  INV_X1 U6522 ( .A(n5367), .ZN(n5368) );
  OAI22_X1 U6523 ( .A1(n5368), .A2(n5466), .B1(n5453), .B2(n4415), .ZN(U2828)
         );
  INV_X1 U6524 ( .A(n5741), .ZN(n5370) );
  AOI22_X1 U6525 ( .A1(n5652), .A2(n5445), .B1(n5462), .B2(EBX_REG_30__SCAN_IN), .ZN(n5369) );
  OAI21_X1 U6526 ( .B1(n5370), .B2(n3195), .A(n5369), .ZN(U2829) );
  NAND2_X1 U6527 ( .A1(n5384), .A2(n5372), .ZN(n5373) );
  NAND2_X1 U6528 ( .A1(n5374), .A2(n5373), .ZN(n5660) );
  INV_X1 U6529 ( .A(EBX_REG_28__SCAN_IN), .ZN(n5376) );
  OAI222_X1 U6530 ( .A1(n5660), .A2(n5466), .B1(n5453), .B2(n5376), .C1(n3195), 
        .C2(n5661), .ZN(U2831) );
  OR2_X1 U6531 ( .A1(n5378), .A2(n5377), .ZN(n5379) );
  NAND2_X1 U6532 ( .A1(n5382), .A2(n5381), .ZN(n5383) );
  AND2_X1 U6533 ( .A1(n5384), .A2(n5383), .ZN(n5670) );
  AOI22_X1 U6534 ( .A1(n5670), .A2(n5445), .B1(n5462), .B2(EBX_REG_27__SCAN_IN), .ZN(n5385) );
  OAI21_X1 U6535 ( .B1(n5495), .B2(n3195), .A(n5385), .ZN(U2832) );
  INV_X1 U6536 ( .A(n5386), .ZN(n5387) );
  INV_X1 U6537 ( .A(n5773), .ZN(n5688) );
  AOI21_X1 U6538 ( .B1(n5392), .B2(n5391), .A(n5390), .ZN(n5803) );
  AOI22_X1 U6539 ( .A1(n5803), .A2(n5445), .B1(n5462), .B2(EBX_REG_25__SCAN_IN), .ZN(n5393) );
  OAI21_X1 U6540 ( .B1(n5688), .B2(n3195), .A(n5393), .ZN(U2834) );
  AOI21_X1 U6541 ( .B1(n5395), .B2(n3226), .A(n5266), .ZN(n5753) );
  OR2_X1 U6542 ( .A1(n5397), .A2(n5396), .ZN(n5398) );
  NAND2_X1 U6543 ( .A1(n5255), .A2(n5398), .ZN(n5704) );
  INV_X1 U6544 ( .A(EBX_REG_23__SCAN_IN), .ZN(n5698) );
  OAI22_X1 U6545 ( .A1(n5704), .A2(n5466), .B1(n5698), .B2(n5453), .ZN(n5399)
         );
  AOI21_X1 U6546 ( .B1(n5753), .B2(n6975), .A(n5399), .ZN(n5400) );
  INV_X1 U6547 ( .A(n5400), .ZN(U2836) );
  NAND2_X1 U6548 ( .A1(n5417), .A2(n5401), .ZN(n5406) );
  INV_X1 U6549 ( .A(n5406), .ZN(n5402) );
  XNOR2_X1 U6550 ( .A(n5409), .B(n5405), .ZN(n5710) );
  INV_X1 U6551 ( .A(EBX_REG_22__SCAN_IN), .ZN(n6910) );
  OAI222_X1 U6552 ( .A1(n5711), .A2(n3195), .B1(n5466), .B2(n5710), .C1(n5453), 
        .C2(n6910), .ZN(U2837) );
  AND2_X1 U6553 ( .A1(n5417), .A2(n5412), .ZN(n5408) );
  OAI21_X1 U6554 ( .B1(n5408), .B2(n5407), .A(n5406), .ZN(n5718) );
  AOI21_X1 U6555 ( .B1(n3220), .B2(n5410), .A(n5409), .ZN(n5716) );
  AOI22_X1 U6556 ( .A1(n5716), .A2(n5445), .B1(n5462), .B2(EBX_REG_21__SCAN_IN), .ZN(n5411) );
  OAI21_X1 U6557 ( .B1(n5718), .B2(n3195), .A(n5411), .ZN(U2838) );
  XOR2_X1 U6558 ( .A(n5417), .B(n5412), .Z(n5759) );
  INV_X1 U6559 ( .A(n5759), .ZN(n5726) );
  MUX2_X1 U6560 ( .A(n5421), .B(n3219), .S(n5413), .Z(n5415) );
  XNOR2_X1 U6561 ( .A(n5415), .B(n5414), .ZN(n5730) );
  INV_X1 U6562 ( .A(n5730), .ZN(n5585) );
  OAI222_X1 U6563 ( .A1(n5726), .A2(n3195), .B1(n5416), .B2(n5453), .C1(n5585), 
        .C2(n5466), .ZN(U2839) );
  AOI21_X1 U6564 ( .B1(n5430), .B2(n5418), .A(n5417), .ZN(n5778) );
  INV_X1 U6565 ( .A(n5778), .ZN(n5425) );
  MUX2_X1 U6566 ( .A(n5421), .B(n5420), .S(n5419), .Z(n5422) );
  INV_X1 U6567 ( .A(n5422), .ZN(n5426) );
  NAND2_X1 U6568 ( .A1(n5436), .A2(n5426), .ZN(n5428) );
  XNOR2_X1 U6569 ( .A(n5428), .B(n5423), .ZN(n5738) );
  AOI22_X1 U6570 ( .A1(n5738), .A2(n5445), .B1(n5462), .B2(EBX_REG_19__SCAN_IN), .ZN(n5424) );
  OAI21_X1 U6571 ( .B1(n5425), .B2(n3195), .A(n5424), .ZN(U2840) );
  OR2_X1 U6572 ( .A1(n5436), .A2(n5426), .ZN(n5427) );
  NAND2_X1 U6573 ( .A1(n5428), .A2(n5427), .ZN(n5848) );
  INV_X1 U6574 ( .A(EBX_REG_18__SCAN_IN), .ZN(n5432) );
  OAI21_X1 U6575 ( .B1(n5434), .B2(n5431), .A(n5430), .ZN(n5847) );
  OAI222_X1 U6576 ( .A1(n5848), .A2(n5466), .B1(n5453), .B2(n5432), .C1(n3195), 
        .C2(n5847), .ZN(U2841) );
  AOI21_X1 U6577 ( .B1(n5443), .B2(n5435), .A(n5434), .ZN(n5998) );
  INV_X1 U6578 ( .A(n5998), .ZN(n5439) );
  AOI21_X1 U6579 ( .B1(n5437), .B2(n5442), .A(n5436), .ZN(n5859) );
  AOI22_X1 U6580 ( .A1(n5859), .A2(n5445), .B1(n5462), .B2(EBX_REG_17__SCAN_IN), .ZN(n5438) );
  OAI21_X1 U6581 ( .B1(n5439), .B2(n3195), .A(n5438), .ZN(U2842) );
  NAND2_X1 U6582 ( .A1(n5292), .A2(n5440), .ZN(n5441) );
  NAND2_X1 U6583 ( .A1(n5442), .A2(n5441), .ZN(n5876) );
  INV_X1 U6584 ( .A(EBX_REG_16__SCAN_IN), .ZN(n6781) );
  OAI21_X1 U6585 ( .B1(n5301), .B2(n5444), .A(n5443), .ZN(n6003) );
  OAI222_X1 U6586 ( .A1(n5876), .A2(n5466), .B1(n5453), .B2(n6781), .C1(n3195), 
        .C2(n6003), .ZN(U2843) );
  INV_X1 U6587 ( .A(n5880), .ZN(n5478) );
  AOI22_X1 U6588 ( .A1(n5881), .A2(n5445), .B1(n5462), .B2(EBX_REG_15__SCAN_IN), .ZN(n5446) );
  OAI21_X1 U6589 ( .B1(n5478), .B2(n3195), .A(n5446), .ZN(U2844) );
  NAND2_X1 U6590 ( .A1(n5454), .A2(n5447), .ZN(n5448) );
  NAND2_X1 U6591 ( .A1(n5449), .A2(n5448), .ZN(n5886) );
  INV_X1 U6592 ( .A(EBX_REG_14__SCAN_IN), .ZN(n6946) );
  OAI21_X1 U6593 ( .B1(n5451), .B2(n5450), .A(n5300), .ZN(n5885) );
  OAI222_X1 U6594 ( .A1(n5886), .A2(n5466), .B1(n5453), .B2(n6946), .C1(n3195), 
        .C2(n5885), .ZN(U2845) );
  INV_X1 U6595 ( .A(n5454), .ZN(n5455) );
  AOI21_X1 U6596 ( .B1(n5457), .B2(n5456), .A(n5455), .ZN(n5895) );
  INV_X1 U6597 ( .A(n5895), .ZN(n5467) );
  OR2_X1 U6598 ( .A1(n5459), .A2(n5458), .ZN(n5461) );
  NAND2_X1 U6599 ( .A1(n5461), .A2(n5460), .ZN(n5904) );
  INV_X1 U6600 ( .A(n5904), .ZN(n5463) );
  AOI22_X1 U6601 ( .A1(n6975), .A2(n5463), .B1(n5462), .B2(EBX_REG_13__SCAN_IN), .ZN(n5465) );
  OAI21_X1 U6602 ( .B1(n5467), .B2(n5466), .A(n5465), .ZN(U2846) );
  NAND3_X1 U6603 ( .A1(n5319), .A2(n5468), .A3(n6967), .ZN(n5470) );
  AOI22_X1 U6604 ( .A1(n5996), .A2(DATAI_31_), .B1(n6005), .B2(
        EAX_REG_31__SCAN_IN), .ZN(n5469) );
  NAND2_X1 U6605 ( .A1(n5470), .A2(n5469), .ZN(U2860) );
  AOI22_X1 U6606 ( .A1(n6006), .A2(DATAI_12_), .B1(EAX_REG_28__SCAN_IN), .B2(
        n6005), .ZN(n5472) );
  NAND2_X1 U6607 ( .A1(n5996), .A2(DATAI_28_), .ZN(n5471) );
  OAI211_X1 U6608 ( .C1(n5661), .C2(n6970), .A(n5472), .B(n5471), .ZN(U2863)
         );
  AOI22_X1 U6609 ( .A1(n6006), .A2(DATAI_6_), .B1(EAX_REG_22__SCAN_IN), .B2(
        n6005), .ZN(n5474) );
  NAND2_X1 U6610 ( .A1(n5996), .A2(DATAI_22_), .ZN(n5473) );
  OAI211_X1 U6611 ( .C1(n5711), .C2(n6970), .A(n5474), .B(n5473), .ZN(U2869)
         );
  AOI22_X1 U6612 ( .A1(n6006), .A2(DATAI_2_), .B1(n6005), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n5476) );
  NAND2_X1 U6613 ( .A1(n5996), .A2(DATAI_18_), .ZN(n5475) );
  OAI211_X1 U6614 ( .C1(n5847), .C2(n6970), .A(n5476), .B(n5475), .ZN(U2873)
         );
  AOI22_X1 U6615 ( .A1(n5479), .A2(DATAI_15_), .B1(n6005), .B2(
        EAX_REG_15__SCAN_IN), .ZN(n5477) );
  OAI21_X1 U6616 ( .B1(n5478), .B2(n6970), .A(n5477), .ZN(U2876) );
  AOI22_X1 U6617 ( .A1(n5479), .A2(DATAI_14_), .B1(n6005), .B2(
        EAX_REG_14__SCAN_IN), .ZN(n5480) );
  OAI21_X1 U6618 ( .B1(n5885), .B2(n6970), .A(n5480), .ZN(U2877) );
  INV_X1 U6619 ( .A(DATAI_13_), .ZN(n6864) );
  OAI222_X1 U6620 ( .A1(n5904), .A2(n6970), .B1(n6969), .B2(n6864), .C1(n6967), 
        .C2(n6019), .ZN(U2878) );
  NAND3_X1 U6621 ( .A1(n5769), .A2(n5592), .A3(n6749), .ZN(n5481) );
  AOI22_X1 U6622 ( .A1(n5489), .A2(n5481), .B1(INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n6749), .ZN(n5483) );
  XNOR2_X1 U6623 ( .A(n5483), .B(n5482), .ZN(n5531) );
  NAND2_X1 U6624 ( .A1(n5656), .A2(n6134), .ZN(n5484) );
  NAND2_X1 U6625 ( .A1(n6210), .A2(REIP_REG_28__SCAN_IN), .ZN(n5536) );
  OAI211_X1 U6626 ( .C1(n5791), .C2(n5485), .A(n5484), .B(n5536), .ZN(n5486)
         );
  AOI21_X1 U6627 ( .B1(n5531), .B2(n6152), .A(n5486), .ZN(n5487) );
  OAI21_X1 U6628 ( .B1(n5661), .B2(n6138), .A(n5487), .ZN(U2958) );
  NAND2_X1 U6629 ( .A1(n5489), .A2(n5488), .ZN(n5490) );
  XNOR2_X1 U6630 ( .A(n5490), .B(n6749), .ZN(n5541) );
  NOR2_X1 U6631 ( .A1(n5667), .A2(n6157), .ZN(n5493) );
  NAND2_X1 U6632 ( .A1(n6210), .A2(REIP_REG_27__SCAN_IN), .ZN(n5542) );
  OAI21_X1 U6633 ( .B1(n5791), .B2(n5491), .A(n5542), .ZN(n5492) );
  AOI211_X1 U6634 ( .C1(n5541), .C2(n6152), .A(n5493), .B(n5492), .ZN(n5494)
         );
  OAI21_X1 U6635 ( .B1(n5495), .B2(n6138), .A(n5494), .ZN(U2959) );
  NAND3_X1 U6636 ( .A1(n5604), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .A3(n5497), .ZN(n5499) );
  OAI21_X1 U6637 ( .B1(n3215), .B2(n5499), .A(n5498), .ZN(n5500) );
  XNOR2_X1 U6638 ( .A(n5500), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5556)
         );
  NAND2_X1 U6639 ( .A1(n6210), .A2(REIP_REG_23__SCAN_IN), .ZN(n5551) );
  NAND2_X1 U6640 ( .A1(n6147), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5501)
         );
  OAI211_X1 U6641 ( .C1(n5697), .C2(n6157), .A(n5551), .B(n5501), .ZN(n5502)
         );
  AOI21_X1 U6642 ( .B1(n5753), .B2(n4403), .A(n5502), .ZN(n5503) );
  OAI21_X1 U6643 ( .B1(n5556), .B2(n5831), .A(n5503), .ZN(U2963) );
  AOI21_X1 U6644 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n5604), .A(n5505), 
        .ZN(n5506) );
  XNOR2_X1 U6645 ( .A(n5504), .B(n5506), .ZN(n5565) );
  NAND2_X1 U6646 ( .A1(n6210), .A2(REIP_REG_22__SCAN_IN), .ZN(n5561) );
  OAI21_X1 U6647 ( .B1(n5791), .B2(n5507), .A(n5561), .ZN(n5509) );
  NOR2_X1 U6648 ( .A1(n5711), .A2(n6138), .ZN(n5508) );
  AOI211_X1 U6649 ( .C1(n6134), .C2(n5707), .A(n5509), .B(n5508), .ZN(n5510)
         );
  OAI21_X1 U6650 ( .B1(n5565), .B2(n5831), .A(n5510), .ZN(U2964) );
  AOI21_X1 U6651 ( .B1(n5513), .B2(n5512), .A(n5511), .ZN(n5572) );
  INV_X1 U6652 ( .A(n5718), .ZN(n5756) );
  NAND2_X1 U6653 ( .A1(n6210), .A2(REIP_REG_21__SCAN_IN), .ZN(n5566) );
  NAND2_X1 U6654 ( .A1(n6147), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5514)
         );
  OAI211_X1 U6655 ( .C1(n5723), .C2(n6157), .A(n5566), .B(n5514), .ZN(n5515)
         );
  AOI21_X1 U6656 ( .B1(n5756), .B2(n6124), .A(n5515), .ZN(n5516) );
  OAI21_X1 U6657 ( .B1(n5572), .B2(n5831), .A(n5516), .ZN(U2965) );
  XNOR2_X1 U6658 ( .A(n3215), .B(n5517), .ZN(n5588) );
  NAND2_X1 U6659 ( .A1(n6210), .A2(REIP_REG_20__SCAN_IN), .ZN(n5584) );
  NAND2_X1 U6660 ( .A1(n6124), .A2(n5759), .ZN(n5518) );
  OAI211_X1 U6661 ( .C1(n5791), .C2(n5733), .A(n5584), .B(n5518), .ZN(n5519)
         );
  AOI21_X1 U6662 ( .B1(n5724), .B2(n6134), .A(n5519), .ZN(n5520) );
  OAI21_X1 U6663 ( .B1(n5588), .B2(n5831), .A(n5520), .ZN(U2966) );
  INV_X1 U6664 ( .A(n5521), .ZN(n5530) );
  INV_X1 U6665 ( .A(n5522), .ZN(n5545) );
  NAND3_X1 U6666 ( .A1(n5545), .A2(n5532), .A3(n5523), .ZN(n5524) );
  OAI211_X1 U6667 ( .C1(n5526), .C2(n6177), .A(n5525), .B(n5524), .ZN(n5527)
         );
  AOI21_X1 U6668 ( .B1(INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n5528), .A(n5527), 
        .ZN(n5529) );
  OAI21_X1 U6669 ( .B1(n5530), .B2(n5815), .A(n5529), .ZN(U2989) );
  INV_X1 U6670 ( .A(n5531), .ZN(n5540) );
  INV_X1 U6671 ( .A(n5548), .ZN(n5538) );
  INV_X1 U6672 ( .A(n5532), .ZN(n5533) );
  NAND3_X1 U6673 ( .A1(n5545), .A2(n5534), .A3(n5533), .ZN(n5535) );
  OAI211_X1 U6674 ( .C1(n5660), .C2(n6177), .A(n5536), .B(n5535), .ZN(n5537)
         );
  AOI21_X1 U6675 ( .B1(INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n5538), .A(n5537), 
        .ZN(n5539) );
  OAI21_X1 U6676 ( .B1(n5540), .B2(n5815), .A(n5539), .ZN(U2990) );
  NAND2_X1 U6677 ( .A1(n5541), .A2(n6231), .ZN(n5547) );
  INV_X1 U6678 ( .A(n5670), .ZN(n5543) );
  OAI21_X1 U6679 ( .B1(n5543), .B2(n6177), .A(n5542), .ZN(n5544) );
  AOI21_X1 U6680 ( .B1(n5545), .B2(n6749), .A(n5544), .ZN(n5546) );
  OAI211_X1 U6681 ( .C1(n5548), .C2(n6749), .A(n5547), .B(n5546), .ZN(U2991)
         );
  INV_X1 U6682 ( .A(n5549), .ZN(n5554) );
  NOR2_X1 U6683 ( .A1(n5550), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5553)
         );
  OAI21_X1 U6684 ( .B1(n5704), .B2(n6177), .A(n5551), .ZN(n5552) );
  AOI211_X1 U6685 ( .C1(INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n5554), .A(n5553), .B(n5552), .ZN(n5555) );
  OAI21_X1 U6686 ( .B1(n5556), .B2(n5815), .A(n5555), .ZN(U2995) );
  INV_X1 U6687 ( .A(n5557), .ZN(n5558) );
  NAND3_X1 U6688 ( .A1(n5560), .A2(n5559), .A3(n5558), .ZN(n5562) );
  OAI211_X1 U6689 ( .C1(n5710), .C2(n6177), .A(n5562), .B(n5561), .ZN(n5563)
         );
  AOI21_X1 U6690 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n5570), .A(n5563), 
        .ZN(n5564) );
  OAI21_X1 U6691 ( .B1(n5565), .B2(n5815), .A(n5564), .ZN(U2996) );
  NAND2_X1 U6692 ( .A1(n5716), .A2(n6227), .ZN(n5567) );
  OAI211_X1 U6693 ( .C1(n5568), .C2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n5567), .B(n5566), .ZN(n5569) );
  AOI21_X1 U6694 ( .B1(INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n5570), .A(n5569), 
        .ZN(n5571) );
  OAI21_X1 U6695 ( .B1(n5572), .B2(n5815), .A(n5571), .ZN(U2997) );
  AOI21_X1 U6696 ( .B1(n5574), .B2(INSTADDRPOINTER_REG_17__SCAN_IN), .A(n5573), 
        .ZN(n5576) );
  NOR2_X1 U6697 ( .A1(n5576), .A2(n5575), .ZN(n5810) );
  NAND2_X1 U6698 ( .A1(n6212), .A2(n5608), .ZN(n5577) );
  OAI211_X1 U6699 ( .C1(n5579), .C2(n5578), .A(n5810), .B(n5577), .ZN(n5600)
         );
  NOR3_X1 U6700 ( .A1(n5580), .A2(n5594), .A3(n5812), .ZN(n5581) );
  NAND2_X1 U6701 ( .A1(n5582), .A2(n5581), .ZN(n5583) );
  OAI211_X1 U6702 ( .C1(n5585), .C2(n6177), .A(n5584), .B(n5583), .ZN(n5586)
         );
  AOI21_X1 U6703 ( .B1(INSTADDRPOINTER_REG_20__SCAN_IN), .B2(n5600), .A(n5586), 
        .ZN(n5587) );
  OAI21_X1 U6704 ( .B1(n5588), .B2(n5815), .A(n5587), .ZN(U2998) );
  INV_X1 U6705 ( .A(n5589), .ZN(n5591) );
  OAI21_X1 U6706 ( .B1(n5591), .B2(n5595), .A(n5590), .ZN(n5593) );
  XNOR2_X1 U6707 ( .A(n5593), .B(n5592), .ZN(n5777) );
  INV_X1 U6708 ( .A(n5777), .ZN(n5602) );
  INV_X1 U6709 ( .A(n5738), .ZN(n5598) );
  NOR2_X1 U6710 ( .A1(n5594), .A2(n5812), .ZN(n5596) );
  AOI22_X1 U6711 ( .A1(n6210), .A2(REIP_REG_19__SCAN_IN), .B1(n5596), .B2(
        n5595), .ZN(n5597) );
  OAI21_X1 U6712 ( .B1(n5598), .B2(n6177), .A(n5597), .ZN(n5599) );
  AOI21_X1 U6713 ( .B1(n5600), .B2(INSTADDRPOINTER_REG_19__SCAN_IN), .A(n5599), 
        .ZN(n5601) );
  OAI21_X1 U6714 ( .B1(n5602), .B2(n5815), .A(n5601), .ZN(U2999) );
  NOR2_X1 U6715 ( .A1(n5592), .A2(n5625), .ZN(n5787) );
  NAND2_X1 U6716 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n5787), .ZN(n5606) );
  NOR2_X1 U6717 ( .A1(n5604), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5786)
         );
  NAND3_X1 U6718 ( .A1(n5786), .A2(n5811), .A3(n5785), .ZN(n5605) );
  OAI21_X1 U6719 ( .B1(n5606), .B2(n5785), .A(n5605), .ZN(n5607) );
  XNOR2_X1 U6720 ( .A(n5608), .B(n5607), .ZN(n5782) );
  OAI21_X1 U6721 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n5609), .A(n5810), 
        .ZN(n5611) );
  NOR3_X1 U6722 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n5811), .A3(n5812), 
        .ZN(n5610) );
  AOI21_X1 U6723 ( .B1(INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n5611), .A(n5610), 
        .ZN(n5612) );
  OAI21_X1 U6724 ( .B1(n6175), .B2(n6513), .A(n5612), .ZN(n5613) );
  AOI21_X1 U6725 ( .B1(n6231), .B2(n5782), .A(n5613), .ZN(n5614) );
  OAI21_X1 U6726 ( .B1(n5848), .B2(n6177), .A(n5614), .ZN(U3000) );
  INV_X1 U6727 ( .A(n5615), .ZN(n5626) );
  NOR2_X1 U6728 ( .A1(n5787), .A2(n5786), .ZN(n5616) );
  XOR2_X1 U6729 ( .A(n5616), .B(n5785), .Z(n5792) );
  NAND2_X1 U6730 ( .A1(n5792), .A2(n6231), .ZN(n5624) );
  AOI211_X1 U6731 ( .C1(n5618), .C2(n5625), .A(n5823), .B(n5617), .ZN(n5622)
         );
  INV_X1 U6732 ( .A(REIP_REG_16__SCAN_IN), .ZN(n5619) );
  OAI22_X1 U6733 ( .A1(n5876), .A2(n6177), .B1(n6175), .B2(n5619), .ZN(n5620)
         );
  AOI21_X1 U6734 ( .B1(n5622), .B2(n5621), .A(n5620), .ZN(n5623) );
  OAI211_X1 U6735 ( .C1(n5626), .C2(n5625), .A(n5624), .B(n5623), .ZN(U3002)
         );
  XNOR2_X1 U6736 ( .A(n5604), .B(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5628)
         );
  XNOR2_X1 U6737 ( .A(n3213), .B(n5628), .ZN(n5795) );
  INV_X1 U6738 ( .A(n5795), .ZN(n5641) );
  AOI21_X1 U6739 ( .B1(n5630), .B2(n5629), .A(INSTADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n5634) );
  NAND2_X1 U6740 ( .A1(n5631), .A2(n6224), .ZN(n5632) );
  OAI211_X1 U6741 ( .C1(n5635), .C2(n5633), .A(n6164), .B(n5632), .ZN(n5818)
         );
  OAI21_X1 U6742 ( .B1(n5634), .B2(n5818), .A(INSTADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n5640) );
  INV_X1 U6743 ( .A(n5635), .ZN(n5636) );
  NOR3_X1 U6744 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n5823), .A3(n5636), 
        .ZN(n5638) );
  INV_X1 U6745 ( .A(REIP_REG_14__SCAN_IN), .ZN(n6507) );
  OAI22_X1 U6746 ( .A1(n5886), .A2(n6177), .B1(n6507), .B2(n6175), .ZN(n5637)
         );
  NOR2_X1 U6747 ( .A1(n5638), .A2(n5637), .ZN(n5639) );
  OAI211_X1 U6748 ( .C1(n5641), .C2(n5815), .A(n5640), .B(n5639), .ZN(U3004)
         );
  OAI21_X1 U6749 ( .B1(n5642), .B2(STATEBS16_REG_SCAN_IN), .A(n6313), .ZN(
        n5646) );
  OAI22_X1 U6750 ( .A1(n5646), .A2(n5645), .B1(n5644), .B2(n5643), .ZN(n5647)
         );
  MUX2_X1 U6751 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n5647), .S(n6236), 
        .Z(U3464) );
  AND2_X1 U6752 ( .A1(DATAO_REG_31__SCAN_IN), .A2(n6039), .ZN(U2892) );
  AOI22_X1 U6753 ( .A1(EBX_REG_30__SCAN_IN), .A2(n5982), .B1(n5648), .B2(n6537), .ZN(n5649) );
  OAI21_X1 U6754 ( .B1(n6707), .B2(n5970), .A(n5649), .ZN(n5650) );
  AOI21_X1 U6755 ( .B1(n5651), .B2(n5964), .A(n5650), .ZN(n5654) );
  AOI22_X1 U6756 ( .A1(n5652), .A2(n5981), .B1(n5741), .B2(n5952), .ZN(n5653)
         );
  OAI211_X1 U6757 ( .C1(n6537), .C2(n5655), .A(n5654), .B(n5653), .ZN(U2797)
         );
  NAND2_X1 U6758 ( .A1(REIP_REG_27__SCAN_IN), .A2(n5669), .ZN(n5665) );
  INV_X1 U6759 ( .A(REIP_REG_28__SCAN_IN), .ZN(n5658) );
  AOI22_X1 U6760 ( .A1(PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n5983), .B1(n5656), 
        .B2(n5964), .ZN(n5657) );
  OAI21_X1 U6761 ( .B1(n5659), .B2(n5658), .A(n5657), .ZN(n5663) );
  OAI22_X1 U6762 ( .A1(n5661), .A2(n5967), .B1(n5660), .B2(n5969), .ZN(n5662)
         );
  AOI211_X1 U6763 ( .C1(EBX_REG_28__SCAN_IN), .C2(n5982), .A(n5663), .B(n5662), 
        .ZN(n5664) );
  OAI21_X1 U6764 ( .B1(REIP_REG_28__SCAN_IN), .B2(n5665), .A(n5664), .ZN(U2799) );
  INV_X1 U6765 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6528) );
  AOI22_X1 U6766 ( .A1(EBX_REG_27__SCAN_IN), .A2(n5982), .B1(
        PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n5983), .ZN(n5666) );
  OAI21_X1 U6767 ( .B1(n5667), .B2(n5990), .A(n5666), .ZN(n5668) );
  AOI221_X1 U6768 ( .B1(n5676), .B2(REIP_REG_27__SCAN_IN), .C1(n5669), .C2(
        n6528), .A(n5668), .ZN(n5672) );
  AOI22_X1 U6769 ( .A1(n5748), .A2(n5952), .B1(n5670), .B2(n5981), .ZN(n5671)
         );
  NAND2_X1 U6770 ( .A1(n5672), .A2(n5671), .ZN(U2800) );
  AOI22_X1 U6771 ( .A1(PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n5983), .B1(n5764), 
        .B2(n5964), .ZN(n5678) );
  OR2_X1 U6772 ( .A1(n6523), .A2(n5685), .ZN(n5681) );
  OAI21_X1 U6773 ( .B1(n6525), .B2(n5681), .A(n6526), .ZN(n5675) );
  OAI22_X1 U6774 ( .A1(n5768), .A2(n5967), .B1(n5673), .B2(n5969), .ZN(n5674)
         );
  AOI21_X1 U6775 ( .B1(n5676), .B2(n5675), .A(n5674), .ZN(n5677) );
  OAI211_X1 U6776 ( .C1(n5679), .C2(n5961), .A(n5678), .B(n5677), .ZN(U2801)
         );
  INV_X1 U6777 ( .A(EBX_REG_25__SCAN_IN), .ZN(n5680) );
  INV_X1 U6778 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n6893) );
  OAI22_X1 U6779 ( .A1(n5680), .A2(n5961), .B1(n6893), .B2(n5970), .ZN(n5683)
         );
  OAI22_X1 U6780 ( .A1(REIP_REG_25__SCAN_IN), .A2(n5681), .B1(n5776), .B2(
        n5990), .ZN(n5682) );
  AOI211_X1 U6781 ( .C1(n5981), .C2(n5803), .A(n5683), .B(n5682), .ZN(n5687)
         );
  NOR2_X1 U6782 ( .A1(n5865), .A2(n5684), .ZN(n5701) );
  NOR2_X1 U6783 ( .A1(REIP_REG_24__SCAN_IN), .A2(n5685), .ZN(n5693) );
  OAI21_X1 U6784 ( .B1(n5701), .B2(n5693), .A(REIP_REG_25__SCAN_IN), .ZN(n5686) );
  OAI211_X1 U6785 ( .C1(n5688), .C2(n5967), .A(n5687), .B(n5686), .ZN(U2802)
         );
  AOI22_X1 U6786 ( .A1(REIP_REG_24__SCAN_IN), .A2(n5701), .B1(
        PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n5983), .ZN(n5691) );
  AOI22_X1 U6787 ( .A1(EBX_REG_24__SCAN_IN), .A2(n5982), .B1(n5689), .B2(n5964), .ZN(n5690) );
  OAI211_X1 U6788 ( .C1(n5692), .C2(n5967), .A(n5691), .B(n5690), .ZN(n5694)
         );
  NOR2_X1 U6789 ( .A1(n5694), .A2(n5693), .ZN(n5695) );
  OAI21_X1 U6790 ( .B1(n5696), .B2(n5969), .A(n5695), .ZN(U2803) );
  OAI22_X1 U6791 ( .A1(n5698), .A2(n5961), .B1(n5697), .B2(n5990), .ZN(n5699)
         );
  AOI21_X1 U6792 ( .B1(PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n5983), .A(n5699), 
        .ZN(n5703) );
  INV_X1 U6793 ( .A(REIP_REG_22__SCAN_IN), .ZN(n6521) );
  NAND2_X1 U6794 ( .A1(REIP_REG_21__SCAN_IN), .A2(n5706), .ZN(n5709) );
  INV_X1 U6795 ( .A(REIP_REG_23__SCAN_IN), .ZN(n6519) );
  OAI21_X1 U6796 ( .B1(n6521), .B2(n5709), .A(n6519), .ZN(n5700) );
  AOI22_X1 U6797 ( .A1(n5753), .A2(n5952), .B1(n5701), .B2(n5700), .ZN(n5702)
         );
  OAI211_X1 U6798 ( .C1(n5704), .C2(n5969), .A(n5703), .B(n5702), .ZN(U2804)
         );
  NAND2_X1 U6799 ( .A1(n5894), .A2(n5705), .ZN(n5727) );
  INV_X1 U6800 ( .A(REIP_REG_21__SCAN_IN), .ZN(n6517) );
  NAND2_X1 U6801 ( .A1(n5706), .A2(n6517), .ZN(n5721) );
  AOI22_X1 U6802 ( .A1(PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n5983), .B1(n5707), 
        .B2(n5964), .ZN(n5708) );
  OAI21_X1 U6803 ( .B1(REIP_REG_22__SCAN_IN), .B2(n5709), .A(n5708), .ZN(n5713) );
  OAI22_X1 U6804 ( .A1(n5711), .A2(n5967), .B1(n5710), .B2(n5969), .ZN(n5712)
         );
  AOI211_X1 U6805 ( .C1(EBX_REG_22__SCAN_IN), .C2(n5982), .A(n5713), .B(n5712), 
        .ZN(n5714) );
  OAI221_X1 U6806 ( .B1(n6521), .B2(n5727), .C1(n6521), .C2(n5721), .A(n5714), 
        .ZN(U2805) );
  OAI22_X1 U6807 ( .A1(n5715), .A2(n5970), .B1(n6517), .B2(n5727), .ZN(n5720)
         );
  INV_X1 U6808 ( .A(n5716), .ZN(n5717) );
  OAI211_X1 U6809 ( .C1(n5990), .C2(n5723), .A(n5722), .B(n5721), .ZN(U2806)
         );
  AOI22_X1 U6810 ( .A1(EBX_REG_20__SCAN_IN), .A2(n5982), .B1(n5724), .B2(n5964), .ZN(n5732) );
  INV_X1 U6811 ( .A(n5736), .ZN(n5725) );
  AOI21_X1 U6812 ( .B1(REIP_REG_19__SCAN_IN), .B2(n5725), .A(
        REIP_REG_20__SCAN_IN), .ZN(n5728) );
  OAI22_X1 U6813 ( .A1(n5728), .A2(n5727), .B1(n5967), .B2(n5726), .ZN(n5729)
         );
  AOI21_X1 U6814 ( .B1(n5981), .B2(n5730), .A(n5729), .ZN(n5731) );
  OAI211_X1 U6815 ( .C1(n5733), .C2(n5970), .A(n5732), .B(n5731), .ZN(U2807)
         );
  NOR2_X1 U6816 ( .A1(n5865), .A2(n5734), .ZN(n5851) );
  AOI22_X1 U6817 ( .A1(EBX_REG_19__SCAN_IN), .A2(n5982), .B1(
        REIP_REG_19__SCAN_IN), .B2(n5851), .ZN(n5735) );
  OAI21_X1 U6818 ( .B1(REIP_REG_19__SCAN_IN), .B2(n5736), .A(n5735), .ZN(n5737) );
  AOI211_X1 U6819 ( .C1(n5983), .C2(PHYADDRPOINTER_REG_19__SCAN_IN), .A(n5973), 
        .B(n5737), .ZN(n5740) );
  AOI22_X1 U6820 ( .A1(n5981), .A2(n5738), .B1(n5952), .B2(n5778), .ZN(n5739)
         );
  OAI211_X1 U6821 ( .C1(n5781), .C2(n5990), .A(n5740), .B(n5739), .ZN(U2808)
         );
  AOI22_X1 U6822 ( .A1(n5741), .A2(n5997), .B1(n5996), .B2(DATAI_30_), .ZN(
        n5743) );
  AOI22_X1 U6823 ( .A1(n6006), .A2(DATAI_14_), .B1(EAX_REG_30__SCAN_IN), .B2(
        n6005), .ZN(n5742) );
  NAND2_X1 U6824 ( .A1(n5743), .A2(n5742), .ZN(U2861) );
  INV_X1 U6825 ( .A(n5996), .ZN(n6002) );
  INV_X1 U6826 ( .A(DATAI_29_), .ZN(n5744) );
  OAI22_X1 U6827 ( .A1(n5341), .A2(n6970), .B1(n6002), .B2(n5744), .ZN(n5745)
         );
  INV_X1 U6828 ( .A(n5745), .ZN(n5747) );
  AOI22_X1 U6829 ( .A1(n6006), .A2(DATAI_13_), .B1(n6005), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n5746) );
  NAND2_X1 U6830 ( .A1(n5747), .A2(n5746), .ZN(U2862) );
  AOI22_X1 U6831 ( .A1(n5748), .A2(n5997), .B1(n5996), .B2(DATAI_27_), .ZN(
        n5750) );
  AOI22_X1 U6832 ( .A1(n6006), .A2(DATAI_11_), .B1(EAX_REG_27__SCAN_IN), .B2(
        n6005), .ZN(n5749) );
  NAND2_X1 U6833 ( .A1(n5750), .A2(n5749), .ZN(U2864) );
  AOI22_X1 U6834 ( .A1(n5773), .A2(n5997), .B1(n5996), .B2(DATAI_25_), .ZN(
        n5752) );
  AOI22_X1 U6835 ( .A1(n6006), .A2(DATAI_9_), .B1(n6005), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n5751) );
  NAND2_X1 U6836 ( .A1(n5752), .A2(n5751), .ZN(U2866) );
  AOI22_X1 U6837 ( .A1(n5753), .A2(n5997), .B1(n5996), .B2(DATAI_23_), .ZN(
        n5755) );
  AOI22_X1 U6838 ( .A1(n6006), .A2(DATAI_7_), .B1(n6005), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n5754) );
  NAND2_X1 U6839 ( .A1(n5755), .A2(n5754), .ZN(U2868) );
  AOI22_X1 U6840 ( .A1(n5756), .A2(n5997), .B1(n5996), .B2(DATAI_21_), .ZN(
        n5758) );
  AOI22_X1 U6841 ( .A1(n6006), .A2(DATAI_5_), .B1(EAX_REG_21__SCAN_IN), .B2(
        n6005), .ZN(n5757) );
  NAND2_X1 U6842 ( .A1(n5758), .A2(n5757), .ZN(U2870) );
  AOI22_X1 U6843 ( .A1(n5996), .A2(DATAI_20_), .B1(n5997), .B2(n5759), .ZN(
        n5761) );
  AOI22_X1 U6844 ( .A1(n6006), .A2(DATAI_4_), .B1(EAX_REG_20__SCAN_IN), .B2(
        n6005), .ZN(n5760) );
  NAND2_X1 U6845 ( .A1(n5761), .A2(n5760), .ZN(U2871) );
  AOI22_X1 U6846 ( .A1(n5778), .A2(n5997), .B1(n5996), .B2(DATAI_19_), .ZN(
        n5763) );
  AOI22_X1 U6847 ( .A1(n6006), .A2(DATAI_3_), .B1(n6005), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n5762) );
  NAND2_X1 U6848 ( .A1(n5763), .A2(n5762), .ZN(U2872) );
  AOI22_X1 U6849 ( .A1(n6210), .A2(REIP_REG_26__SCAN_IN), .B1(n6147), .B2(
        PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5767) );
  AOI22_X1 U6850 ( .A1(n5765), .A2(n6152), .B1(n5764), .B2(n6134), .ZN(n5766)
         );
  OAI211_X1 U6851 ( .C1(n6138), .C2(n5768), .A(n5767), .B(n5766), .ZN(U2960)
         );
  AOI22_X1 U6852 ( .A1(n6210), .A2(REIP_REG_25__SCAN_IN), .B1(n6147), .B2(
        PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5775) );
  AOI21_X1 U6853 ( .B1(n5771), .B2(n5770), .A(n5769), .ZN(n5772) );
  INV_X1 U6854 ( .A(n5772), .ZN(n5804) );
  AOI22_X1 U6855 ( .A1(n5773), .A2(n4403), .B1(n6152), .B2(n5804), .ZN(n5774)
         );
  OAI211_X1 U6856 ( .C1(n6157), .C2(n5776), .A(n5775), .B(n5774), .ZN(U2961)
         );
  AOI22_X1 U6857 ( .A1(n6210), .A2(REIP_REG_19__SCAN_IN), .B1(n6147), .B2(
        PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5780) );
  AOI22_X1 U6858 ( .A1(n5778), .A2(n6124), .B1(n6152), .B2(n5777), .ZN(n5779)
         );
  OAI211_X1 U6859 ( .C1(n6157), .C2(n5781), .A(n5780), .B(n5779), .ZN(U2967)
         );
  AOI22_X1 U6860 ( .A1(n6210), .A2(REIP_REG_18__SCAN_IN), .B1(n6147), .B2(
        PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n5784) );
  AOI22_X1 U6861 ( .A1(n6152), .A2(n5782), .B1(n6134), .B2(n5850), .ZN(n5783)
         );
  OAI211_X1 U6862 ( .C1(n6138), .C2(n5847), .A(n5784), .B(n5783), .ZN(U2968)
         );
  INV_X1 U6863 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n6907) );
  MUX2_X1 U6864 ( .A(n5787), .B(n5786), .S(n5785), .Z(n5788) );
  XNOR2_X1 U6865 ( .A(n5788), .B(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5816)
         );
  OAI22_X1 U6866 ( .A1(n5816), .A2(n5831), .B1(n6157), .B2(n5857), .ZN(n5789)
         );
  AOI21_X1 U6867 ( .B1(n6124), .B2(n5998), .A(n5789), .ZN(n5790) );
  NAND2_X1 U6868 ( .A1(n6210), .A2(REIP_REG_17__SCAN_IN), .ZN(n5809) );
  OAI211_X1 U6869 ( .C1(n6907), .C2(n5791), .A(n5790), .B(n5809), .ZN(U2969)
         );
  AOI22_X1 U6870 ( .A1(n6210), .A2(REIP_REG_16__SCAN_IN), .B1(n6147), .B2(
        PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5794) );
  AOI22_X1 U6871 ( .A1(n5792), .A2(n6152), .B1(n6134), .B2(n5873), .ZN(n5793)
         );
  OAI211_X1 U6872 ( .C1(n6138), .C2(n6003), .A(n5794), .B(n5793), .ZN(U2970)
         );
  AOI22_X1 U6873 ( .A1(n6210), .A2(REIP_REG_14__SCAN_IN), .B1(n6147), .B2(
        PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5797) );
  AOI22_X1 U6874 ( .A1(n5795), .A2(n6152), .B1(n6134), .B2(n5888), .ZN(n5796)
         );
  OAI211_X1 U6875 ( .C1(n6138), .C2(n5885), .A(n5797), .B(n5796), .ZN(U2972)
         );
  AOI22_X1 U6876 ( .A1(n6210), .A2(REIP_REG_13__SCAN_IN), .B1(n6147), .B2(
        PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n5801) );
  XNOR2_X1 U6877 ( .A(n5798), .B(n5799), .ZN(n5819) );
  AOI22_X1 U6878 ( .A1(n5819), .A2(n6152), .B1(n6134), .B2(n5901), .ZN(n5800)
         );
  OAI211_X1 U6879 ( .C1(n6138), .C2(n5904), .A(n5801), .B(n5800), .ZN(U2973)
         );
  AOI22_X1 U6880 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6210), .B1(n5802), .B2(
        n5807), .ZN(n5806) );
  AOI22_X1 U6881 ( .A1(n5804), .A2(n6231), .B1(n6227), .B2(n5803), .ZN(n5805)
         );
  OAI211_X1 U6882 ( .C1(n5808), .C2(n5807), .A(n5806), .B(n5805), .ZN(U2993)
         );
  OAI221_X1 U6883 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n5812), .C1(
        n5811), .C2(n5810), .A(n5809), .ZN(n5813) );
  AOI21_X1 U6884 ( .B1(n5859), .B2(n6227), .A(n5813), .ZN(n5814) );
  OAI21_X1 U6885 ( .B1(n5816), .B2(n5815), .A(n5814), .ZN(U3001) );
  NAND2_X1 U6886 ( .A1(n5817), .A2(n4294), .ZN(n5822) );
  AOI22_X1 U6887 ( .A1(n5895), .A2(n6227), .B1(n6210), .B2(
        REIP_REG_13__SCAN_IN), .ZN(n5821) );
  AOI22_X1 U6888 ( .A1(n5819), .A2(n6231), .B1(INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n5818), .ZN(n5820) );
  OAI211_X1 U6889 ( .C1(n5823), .C2(n5822), .A(n5821), .B(n5820), .ZN(U3005)
         );
  INV_X1 U6890 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6475) );
  AOI21_X1 U6891 ( .B1(STATE_REG_1__SCAN_IN), .B2(n6475), .A(n6798), .ZN(n5829) );
  INV_X1 U6892 ( .A(ADS_N_REG_SCAN_IN), .ZN(n6913) );
  INV_X1 U6893 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6482) );
  NOR2_X2 U6894 ( .A1(STATE_REG_0__SCAN_IN), .A2(n6482), .ZN(n6575) );
  AOI21_X1 U6895 ( .B1(n5829), .B2(n6913), .A(n6575), .ZN(U2789) );
  INV_X1 U6896 ( .A(n5824), .ZN(n5825) );
  OAI21_X1 U6897 ( .B1(n5825), .B2(n6461), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n5826) );
  OAI21_X1 U6898 ( .B1(n5827), .B2(n6567), .A(n5826), .ZN(U2790) );
  INV_X2 U6899 ( .A(n6575), .ZN(n6573) );
  NOR2_X1 U6900 ( .A1(STATE_REG_0__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n5830) );
  OAI21_X1 U6901 ( .B1(D_C_N_REG_SCAN_IN), .B2(n5830), .A(n6573), .ZN(n5828)
         );
  OAI21_X1 U6902 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n6573), .A(n5828), .ZN(
        U2791) );
  NOR2_X1 U6903 ( .A1(n6575), .A2(n5829), .ZN(n6544) );
  OAI21_X1 U6904 ( .B1(n5830), .B2(BS16_N), .A(n6544), .ZN(n6542) );
  OAI21_X1 U6905 ( .B1(n6544), .B2(n6564), .A(n6542), .ZN(U2792) );
  OAI21_X1 U6906 ( .B1(n5833), .B2(n5832), .A(n5831), .ZN(U2793) );
  NOR4_X1 U6907 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(
        DATAWIDTH_REG_16__SCAN_IN), .A3(DATAWIDTH_REG_17__SCAN_IN), .A4(
        DATAWIDTH_REG_22__SCAN_IN), .ZN(n5837) );
  NOR4_X1 U6908 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(DATAWIDTH_REG_10__SCAN_IN), .A3(DATAWIDTH_REG_11__SCAN_IN), .A4(DATAWIDTH_REG_12__SCAN_IN), .ZN(n5836)
         );
  NOR4_X1 U6909 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(
        DATAWIDTH_REG_29__SCAN_IN), .A3(DATAWIDTH_REG_30__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n5835) );
  NOR4_X1 U6910 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(
        DATAWIDTH_REG_25__SCAN_IN), .A3(DATAWIDTH_REG_26__SCAN_IN), .A4(
        DATAWIDTH_REG_27__SCAN_IN), .ZN(n5834) );
  NAND4_X1 U6911 ( .A1(n5837), .A2(n5836), .A3(n5835), .A4(n5834), .ZN(n5843)
         );
  NOR4_X1 U6912 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(DATAWIDTH_REG_4__SCAN_IN), .A3(DATAWIDTH_REG_8__SCAN_IN), .A4(DATAWIDTH_REG_21__SCAN_IN), .ZN(n5841) );
  AOI211_X1 U6913 ( .C1(DATAWIDTH_REG_1__SCAN_IN), .C2(
        DATAWIDTH_REG_0__SCAN_IN), .A(DATAWIDTH_REG_19__SCAN_IN), .B(
        DATAWIDTH_REG_23__SCAN_IN), .ZN(n5840) );
  NOR4_X1 U6914 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(DATAWIDTH_REG_5__SCAN_IN), 
        .A3(DATAWIDTH_REG_6__SCAN_IN), .A4(DATAWIDTH_REG_7__SCAN_IN), .ZN(
        n5839) );
  NOR4_X1 U6915 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(
        DATAWIDTH_REG_13__SCAN_IN), .A3(DATAWIDTH_REG_20__SCAN_IN), .A4(
        DATAWIDTH_REG_2__SCAN_IN), .ZN(n5838) );
  NAND4_X1 U6916 ( .A1(n5841), .A2(n5840), .A3(n5839), .A4(n5838), .ZN(n5842)
         );
  NOR2_X1 U6917 ( .A1(n5843), .A2(n5842), .ZN(n6562) );
  INV_X1 U6918 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n6538) );
  NOR3_X1 U6919 ( .A1(REIP_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .A3(DATAWIDTH_REG_0__SCAN_IN), .ZN(n5845) );
  OAI21_X1 U6920 ( .B1(REIP_REG_1__SCAN_IN), .B2(n5845), .A(n6562), .ZN(n5844)
         );
  OAI21_X1 U6921 ( .B1(n6562), .B2(n6538), .A(n5844), .ZN(U2794) );
  INV_X1 U6922 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6543) );
  AOI21_X1 U6923 ( .B1(n6555), .B2(n6543), .A(n5845), .ZN(n5846) );
  INV_X1 U6924 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n6847) );
  INV_X1 U6925 ( .A(n6562), .ZN(n6557) );
  AOI22_X1 U6926 ( .A1(n6562), .A2(n5846), .B1(n6847), .B2(n6557), .ZN(U2795)
         );
  AOI22_X1 U6927 ( .A1(EBX_REG_18__SCAN_IN), .A2(n5982), .B1(
        PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n5983), .ZN(n5855) );
  OAI22_X1 U6928 ( .A1(n5969), .A2(n5848), .B1(n5967), .B2(n5847), .ZN(n5849)
         );
  AOI21_X1 U6929 ( .B1(n5850), .B2(n5964), .A(n5849), .ZN(n5854) );
  OAI21_X1 U6930 ( .B1(REIP_REG_18__SCAN_IN), .B2(n5852), .A(n5851), .ZN(n5853) );
  NAND4_X1 U6931 ( .A1(n5855), .A2(n5854), .A3(n5958), .A4(n5853), .ZN(U2809)
         );
  INV_X1 U6932 ( .A(REIP_REG_15__SCAN_IN), .ZN(n6811) );
  NOR2_X1 U6933 ( .A1(n6811), .A2(n5866), .ZN(n5863) );
  OAI221_X1 U6934 ( .B1(REIP_REG_17__SCAN_IN), .B2(REIP_REG_16__SCAN_IN), .C1(
        REIP_REG_17__SCAN_IN), .C2(n5863), .A(n5856), .ZN(n5862) );
  OAI22_X1 U6935 ( .A1(n6907), .A2(n5970), .B1(n5857), .B2(n5990), .ZN(n5858)
         );
  AOI211_X1 U6936 ( .C1(n5982), .C2(EBX_REG_17__SCAN_IN), .A(n5973), .B(n5858), 
        .ZN(n5861) );
  AOI22_X1 U6937 ( .A1(n5981), .A2(n5859), .B1(n5952), .B2(n5998), .ZN(n5860)
         );
  OAI211_X1 U6938 ( .C1(n5865), .C2(n5862), .A(n5861), .B(n5860), .ZN(U2810)
         );
  INV_X1 U6939 ( .A(n5863), .ZN(n5868) );
  NOR2_X1 U6940 ( .A1(n5865), .A2(n5864), .ZN(n5889) );
  NOR2_X1 U6941 ( .A1(REIP_REG_15__SCAN_IN), .A2(n5866), .ZN(n5879) );
  NOR2_X1 U6942 ( .A1(n5889), .A2(n5879), .ZN(n5867) );
  MUX2_X1 U6943 ( .A(n5868), .B(n5867), .S(REIP_REG_16__SCAN_IN), .Z(n5869) );
  OAI211_X1 U6944 ( .C1(n5970), .C2(n5870), .A(n5869), .B(n5958), .ZN(n5871)
         );
  AOI21_X1 U6945 ( .B1(EBX_REG_16__SCAN_IN), .B2(n5982), .A(n5871), .ZN(n5875)
         );
  INV_X1 U6946 ( .A(n6003), .ZN(n5872) );
  AOI22_X1 U6947 ( .A1(n5873), .A2(n5964), .B1(n5952), .B2(n5872), .ZN(n5874)
         );
  OAI211_X1 U6948 ( .C1(n5969), .C2(n5876), .A(n5875), .B(n5874), .ZN(U2811)
         );
  AOI22_X1 U6949 ( .A1(EBX_REG_15__SCAN_IN), .A2(n5982), .B1(
        REIP_REG_15__SCAN_IN), .B2(n5889), .ZN(n5877) );
  OAI211_X1 U6950 ( .C1(n5970), .C2(n5305), .A(n5877), .B(n5958), .ZN(n5878)
         );
  AOI211_X1 U6951 ( .C1(n5880), .C2(n5952), .A(n5879), .B(n5878), .ZN(n5884)
         );
  AOI22_X1 U6952 ( .A1(n5882), .A2(n5964), .B1(n5981), .B2(n5881), .ZN(n5883)
         );
  NAND2_X1 U6953 ( .A1(n5884), .A2(n5883), .ZN(U2812) );
  AOI22_X1 U6954 ( .A1(EBX_REG_14__SCAN_IN), .A2(n5982), .B1(
        PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n5983), .ZN(n5892) );
  OAI22_X1 U6955 ( .A1(n5969), .A2(n5886), .B1(n5967), .B2(n5885), .ZN(n5887)
         );
  AOI21_X1 U6956 ( .B1(n5888), .B2(n5964), .A(n5887), .ZN(n5891) );
  INV_X1 U6957 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6505) );
  INV_X1 U6958 ( .A(REIP_REG_12__SCAN_IN), .ZN(n5905) );
  NOR2_X1 U6959 ( .A1(n6505), .A2(n5905), .ZN(n5896) );
  OAI221_X1 U6960 ( .B1(REIP_REG_14__SCAN_IN), .B2(n5896), .C1(
        REIP_REG_14__SCAN_IN), .C2(n5906), .A(n5889), .ZN(n5890) );
  NAND4_X1 U6961 ( .A1(n5892), .A2(n5891), .A3(n5958), .A4(n5890), .ZN(U2813)
         );
  AND2_X1 U6962 ( .A1(n5894), .A2(n5893), .ZN(n5915) );
  AOI22_X1 U6963 ( .A1(n5981), .A2(n5895), .B1(REIP_REG_13__SCAN_IN), .B2(
        n5915), .ZN(n5903) );
  INV_X1 U6964 ( .A(EBX_REG_13__SCAN_IN), .ZN(n5899) );
  AOI21_X1 U6965 ( .B1(n6505), .B2(n5905), .A(n5896), .ZN(n5897) );
  AOI22_X1 U6966 ( .A1(PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n5983), .B1(n5906), 
        .B2(n5897), .ZN(n5898) );
  OAI211_X1 U6967 ( .C1(n5961), .C2(n5899), .A(n5898), .B(n5958), .ZN(n5900)
         );
  AOI21_X1 U6968 ( .B1(n5901), .B2(n5964), .A(n5900), .ZN(n5902) );
  OAI211_X1 U6969 ( .C1(n5967), .C2(n5904), .A(n5903), .B(n5902), .ZN(U2814)
         );
  AOI22_X1 U6970 ( .A1(n5981), .A2(n5907), .B1(n5906), .B2(n5905), .ZN(n5913)
         );
  AOI22_X1 U6971 ( .A1(EBX_REG_12__SCAN_IN), .A2(n5982), .B1(
        PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n5983), .ZN(n5912) );
  AOI21_X1 U6972 ( .B1(REIP_REG_12__SCAN_IN), .B2(n5915), .A(n5973), .ZN(n5911) );
  AOI22_X1 U6973 ( .A1(n5909), .A2(n5964), .B1(n5952), .B2(n5908), .ZN(n5910)
         );
  NAND4_X1 U6974 ( .A1(n5913), .A2(n5912), .A3(n5911), .A4(n5910), .ZN(U2815)
         );
  NOR2_X1 U6975 ( .A1(n5976), .A2(n5928), .ZN(n5929) );
  INV_X1 U6976 ( .A(n5929), .ZN(n5927) );
  NOR3_X1 U6977 ( .A1(n5927), .A2(REIP_REG_11__SCAN_IN), .A3(n5914), .ZN(n5919) );
  INV_X1 U6978 ( .A(EBX_REG_11__SCAN_IN), .ZN(n5917) );
  AOI22_X1 U6979 ( .A1(PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n5983), .B1(
        REIP_REG_11__SCAN_IN), .B2(n5915), .ZN(n5916) );
  OAI211_X1 U6980 ( .C1(n5961), .C2(n5917), .A(n5916), .B(n5958), .ZN(n5918)
         );
  AOI211_X1 U6981 ( .C1(n6158), .C2(n5981), .A(n5919), .B(n5918), .ZN(n5921)
         );
  NAND2_X1 U6982 ( .A1(n6086), .A2(n5964), .ZN(n5920) );
  OAI211_X1 U6983 ( .C1(n6089), .C2(n5967), .A(n5921), .B(n5920), .ZN(U2816)
         );
  OAI22_X1 U6984 ( .A1(n5923), .A2(n5961), .B1(n5969), .B2(n5922), .ZN(n5924)
         );
  AOI211_X1 U6985 ( .C1(n5983), .C2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n5973), 
        .B(n5924), .ZN(n5933) );
  AOI22_X1 U6986 ( .A1(n5926), .A2(n5964), .B1(n5952), .B2(n5925), .ZN(n5932)
         );
  NOR2_X1 U6987 ( .A1(n5927), .A2(REIP_REG_9__SCAN_IN), .ZN(n5937) );
  NAND2_X1 U6988 ( .A1(n5986), .A2(n5928), .ZN(n5940) );
  NAND2_X1 U6989 ( .A1(n5953), .A2(n5940), .ZN(n5942) );
  OAI21_X1 U6990 ( .B1(n5937), .B2(n5942), .A(REIP_REG_10__SCAN_IN), .ZN(n5931) );
  NAND3_X1 U6991 ( .A1(REIP_REG_9__SCAN_IN), .A2(n5929), .A3(n6501), .ZN(n5930) );
  NAND4_X1 U6992 ( .A1(n5933), .A2(n5932), .A3(n5931), .A4(n5930), .ZN(U2817)
         );
  AOI22_X1 U6993 ( .A1(EBX_REG_9__SCAN_IN), .A2(n5982), .B1(
        REIP_REG_9__SCAN_IN), .B2(n5942), .ZN(n5934) );
  OAI211_X1 U6994 ( .C1(n5970), .C2(n5935), .A(n5934), .B(n5958), .ZN(n5936)
         );
  AOI211_X1 U6995 ( .C1(n6166), .C2(n5981), .A(n5937), .B(n5936), .ZN(n5939)
         );
  NAND2_X1 U6996 ( .A1(n6094), .A2(n5964), .ZN(n5938) );
  OAI211_X1 U6997 ( .C1(n6097), .C2(n5967), .A(n5939), .B(n5938), .ZN(U2818)
         );
  OAI22_X1 U6998 ( .A1(n5969), .A2(n6176), .B1(n5941), .B2(n5940), .ZN(n5946)
         );
  AOI22_X1 U6999 ( .A1(PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n5983), .B1(
        REIP_REG_8__SCAN_IN), .B2(n5942), .ZN(n5943) );
  OAI211_X1 U7000 ( .C1(n5961), .C2(n5944), .A(n5943), .B(n5958), .ZN(n5945)
         );
  AOI211_X1 U7001 ( .C1(n6102), .C2(n5964), .A(n5946), .B(n5945), .ZN(n5947)
         );
  OAI21_X1 U7002 ( .B1(n5967), .B2(n6105), .A(n5947), .ZN(U2819) );
  INV_X1 U7003 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6496) );
  NAND3_X1 U7004 ( .A1(n5986), .A2(REIP_REG_5__SCAN_IN), .A3(n5974), .ZN(n5955) );
  NOR3_X1 U7005 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6496), .A3(n5955), .ZN(n5951)
         );
  INV_X1 U7006 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n5949) );
  AOI22_X1 U7007 ( .A1(EBX_REG_7__SCAN_IN), .A2(n5982), .B1(n5981), .B2(n6183), 
        .ZN(n5948) );
  OAI211_X1 U7008 ( .C1(n5970), .C2(n5949), .A(n5948), .B(n5958), .ZN(n5950)
         );
  AOI211_X1 U7009 ( .C1(n6110), .C2(n5952), .A(n5951), .B(n5950), .ZN(n5957)
         );
  OAI21_X1 U7010 ( .B1(n5954), .B2(n5976), .A(n5953), .ZN(n5978) );
  NOR2_X1 U7011 ( .A1(REIP_REG_6__SCAN_IN), .A2(n5955), .ZN(n5963) );
  OAI21_X1 U7012 ( .B1(n5978), .B2(n5963), .A(REIP_REG_7__SCAN_IN), .ZN(n5956)
         );
  OAI211_X1 U7013 ( .C1(n5990), .C2(n6113), .A(n5957), .B(n5956), .ZN(U2820)
         );
  INV_X1 U7014 ( .A(EBX_REG_6__SCAN_IN), .ZN(n5960) );
  AOI22_X1 U7015 ( .A1(PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n5983), .B1(n5981), 
        .B2(n6190), .ZN(n5959) );
  OAI211_X1 U7016 ( .C1(n5961), .C2(n5960), .A(n5959), .B(n5958), .ZN(n5962)
         );
  AOI211_X1 U7017 ( .C1(n5978), .C2(REIP_REG_6__SCAN_IN), .A(n5963), .B(n5962), 
        .ZN(n5966) );
  NAND2_X1 U7018 ( .A1(n6118), .A2(n5964), .ZN(n5965) );
  OAI211_X1 U7019 ( .C1(n6121), .C2(n5967), .A(n5966), .B(n5965), .ZN(U2821)
         );
  INV_X1 U7020 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n5971) );
  OAI22_X1 U7021 ( .A1(n5971), .A2(n5970), .B1(n5969), .B2(n5968), .ZN(n5972)
         );
  AOI211_X1 U7022 ( .C1(n5982), .C2(EBX_REG_5__SCAN_IN), .A(n5973), .B(n5972), 
        .ZN(n5980) );
  INV_X1 U7023 ( .A(n5974), .ZN(n5975) );
  OAI21_X1 U7024 ( .B1(n5976), .B2(n5975), .A(n4642), .ZN(n5977) );
  AOI22_X1 U7025 ( .A1(n5992), .A2(n6123), .B1(n5978), .B2(n5977), .ZN(n5979)
         );
  OAI211_X1 U7026 ( .C1(n6128), .C2(n5990), .A(n5980), .B(n5979), .ZN(U2822)
         );
  INV_X1 U7027 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6801) );
  AOI22_X1 U7028 ( .A1(EBX_REG_3__SCAN_IN), .A2(n5982), .B1(n5981), .B2(n6203), 
        .ZN(n5994) );
  AOI22_X1 U7029 ( .A1(n6311), .A2(n5984), .B1(PHYADDRPOINTER_REG_3__SCAN_IN), 
        .B2(n5983), .ZN(n5989) );
  NAND3_X1 U7030 ( .A1(n5987), .A2(n5986), .A3(n5985), .ZN(n5988) );
  OAI211_X1 U7031 ( .C1(n5990), .C2(n6146), .A(n5989), .B(n5988), .ZN(n5991)
         );
  AOI21_X1 U7032 ( .B1(n6143), .B2(n5992), .A(n5991), .ZN(n5993) );
  OAI211_X1 U7033 ( .C1(n5995), .C2(n6801), .A(n5994), .B(n5993), .ZN(U2824)
         );
  AOI22_X1 U7034 ( .A1(n5998), .A2(n5997), .B1(n5996), .B2(DATAI_17_), .ZN(
        n6000) );
  AOI22_X1 U7035 ( .A1(n6006), .A2(DATAI_1_), .B1(n6005), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n5999) );
  NAND2_X1 U7036 ( .A1(n6000), .A2(n5999), .ZN(U2874) );
  INV_X1 U7037 ( .A(DATAI_16_), .ZN(n6001) );
  OAI22_X1 U7038 ( .A1(n6003), .A2(n6970), .B1(n6002), .B2(n6001), .ZN(n6004)
         );
  INV_X1 U7039 ( .A(n6004), .ZN(n6008) );
  AOI22_X1 U7040 ( .A1(n6006), .A2(DATAI_0_), .B1(n6005), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n6007) );
  NAND2_X1 U7041 ( .A1(n6008), .A2(n6007), .ZN(U2875) );
  INV_X1 U7042 ( .A(DATAO_REG_22__SCAN_IN), .ZN(n6738) );
  INV_X1 U7043 ( .A(n6009), .ZN(n6013) );
  AOI22_X1 U7044 ( .A1(n6013), .A2(EAX_REG_22__SCAN_IN), .B1(n6040), .B2(
        UWORD_REG_6__SCAN_IN), .ZN(n6010) );
  OAI21_X1 U7045 ( .B1(n6738), .B2(n6035), .A(n6010), .ZN(U2901) );
  INV_X1 U7046 ( .A(UWORD_REG_5__SCAN_IN), .ZN(n6796) );
  AOI22_X1 U7047 ( .A1(n6039), .A2(DATAO_REG_21__SCAN_IN), .B1(n6013), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n6011) );
  OAI21_X1 U7048 ( .B1(n6796), .B2(n6033), .A(n6011), .ZN(U2902) );
  INV_X1 U7049 ( .A(DATAO_REG_19__SCAN_IN), .ZN(n6912) );
  AOI22_X1 U7050 ( .A1(n6013), .A2(EAX_REG_19__SCAN_IN), .B1(n6040), .B2(
        UWORD_REG_3__SCAN_IN), .ZN(n6012) );
  OAI21_X1 U7051 ( .B1(n6912), .B2(n6035), .A(n6012), .ZN(U2904) );
  INV_X1 U7052 ( .A(UWORD_REG_1__SCAN_IN), .ZN(n6721) );
  AOI22_X1 U7053 ( .A1(n6039), .A2(DATAO_REG_17__SCAN_IN), .B1(n6013), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n6014) );
  OAI21_X1 U7054 ( .B1(n6721), .B2(n6033), .A(n6014), .ZN(U2906) );
  AOI22_X1 U7055 ( .A1(EAX_REG_15__SCAN_IN), .A2(n6029), .B1(n6039), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n6015) );
  OAI21_X1 U7056 ( .B1(n6814), .B2(n6033), .A(n6015), .ZN(U2908) );
  INV_X1 U7057 ( .A(EAX_REG_14__SCAN_IN), .ZN(n6017) );
  AOI22_X1 U7058 ( .A1(n6040), .A2(LWORD_REG_14__SCAN_IN), .B1(n6039), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n6016) );
  OAI21_X1 U7059 ( .B1(n6017), .B2(n6042), .A(n6016), .ZN(U2909) );
  AOI22_X1 U7060 ( .A1(n6040), .A2(LWORD_REG_13__SCAN_IN), .B1(n6039), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n6018) );
  OAI21_X1 U7061 ( .B1(n6019), .B2(n6042), .A(n6018), .ZN(U2910) );
  INV_X1 U7062 ( .A(DATAO_REG_12__SCAN_IN), .ZN(n6891) );
  AOI22_X1 U7063 ( .A1(EAX_REG_12__SCAN_IN), .A2(n6029), .B1(n6040), .B2(
        LWORD_REG_12__SCAN_IN), .ZN(n6020) );
  OAI21_X1 U7064 ( .B1(n6891), .B2(n6035), .A(n6020), .ZN(U2911) );
  INV_X1 U7065 ( .A(DATAO_REG_11__SCAN_IN), .ZN(n6695) );
  AOI22_X1 U7066 ( .A1(EAX_REG_11__SCAN_IN), .A2(n6029), .B1(n6040), .B2(
        LWORD_REG_11__SCAN_IN), .ZN(n6021) );
  OAI21_X1 U7067 ( .B1(n6695), .B2(n6035), .A(n6021), .ZN(U2912) );
  AOI22_X1 U7068 ( .A1(DATAO_REG_10__SCAN_IN), .A2(n6039), .B1(n6040), .B2(
        LWORD_REG_10__SCAN_IN), .ZN(n6022) );
  OAI21_X1 U7069 ( .B1(n6023), .B2(n6042), .A(n6022), .ZN(U2913) );
  INV_X1 U7070 ( .A(DATAO_REG_9__SCAN_IN), .ZN(n6775) );
  AOI22_X1 U7071 ( .A1(EAX_REG_9__SCAN_IN), .A2(n6029), .B1(n6040), .B2(
        LWORD_REG_9__SCAN_IN), .ZN(n6024) );
  OAI21_X1 U7072 ( .B1(n6775), .B2(n6035), .A(n6024), .ZN(U2914) );
  AOI22_X1 U7073 ( .A1(n6040), .A2(LWORD_REG_8__SCAN_IN), .B1(n6039), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n6025) );
  OAI21_X1 U7074 ( .B1(n6026), .B2(n6042), .A(n6025), .ZN(U2915) );
  INV_X1 U7075 ( .A(EAX_REG_7__SCAN_IN), .ZN(n6028) );
  AOI22_X1 U7076 ( .A1(n6040), .A2(LWORD_REG_7__SCAN_IN), .B1(n6039), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n6027) );
  OAI21_X1 U7077 ( .B1(n6028), .B2(n6042), .A(n6027), .ZN(U2916) );
  INV_X1 U7078 ( .A(LWORD_REG_6__SCAN_IN), .ZN(n6840) );
  AOI22_X1 U7079 ( .A1(EAX_REG_6__SCAN_IN), .A2(n6029), .B1(n6039), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n6030) );
  OAI21_X1 U7080 ( .B1(n6840), .B2(n6033), .A(n6030), .ZN(U2917) );
  AOI22_X1 U7081 ( .A1(n6040), .A2(LWORD_REG_5__SCAN_IN), .B1(n6039), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n6031) );
  OAI21_X1 U7082 ( .B1(n4796), .B2(n6042), .A(n6031), .ZN(U2918) );
  INV_X1 U7083 ( .A(DATAO_REG_4__SCAN_IN), .ZN(n6826) );
  INV_X1 U7084 ( .A(LWORD_REG_4__SCAN_IN), .ZN(n6032) );
  OAI222_X1 U7085 ( .A1(n6035), .A2(n6826), .B1(n6042), .B2(n6034), .C1(n6033), 
        .C2(n6032), .ZN(U2919) );
  AOI22_X1 U7086 ( .A1(DATAO_REG_3__SCAN_IN), .A2(n6039), .B1(n6040), .B2(
        LWORD_REG_3__SCAN_IN), .ZN(n6036) );
  OAI21_X1 U7087 ( .B1(n3683), .B2(n6042), .A(n6036), .ZN(U2920) );
  AOI22_X1 U7088 ( .A1(n6040), .A2(LWORD_REG_2__SCAN_IN), .B1(n6039), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n6037) );
  OAI21_X1 U7089 ( .B1(n3649), .B2(n6042), .A(n6037), .ZN(U2921) );
  AOI22_X1 U7090 ( .A1(LWORD_REG_1__SCAN_IN), .A2(n6040), .B1(n6039), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n6038) );
  OAI21_X1 U7091 ( .B1(n3629), .B2(n6042), .A(n6038), .ZN(U2922) );
  AOI22_X1 U7092 ( .A1(LWORD_REG_0__SCAN_IN), .A2(n6040), .B1(n6039), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n6041) );
  OAI21_X1 U7093 ( .B1(n6043), .B2(n6042), .A(n6041), .ZN(U2923) );
  AOI22_X1 U7094 ( .A1(UWORD_REG_0__SCAN_IN), .A2(n6074), .B1(n6079), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n6046) );
  OAI21_X1 U7095 ( .B1(n6081), .B2(n6861), .A(n6046), .ZN(U2924) );
  AOI22_X1 U7096 ( .A1(UWORD_REG_1__SCAN_IN), .A2(n6051), .B1(n6079), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n6047) );
  OAI21_X1 U7097 ( .B1(n6081), .B2(n6890), .A(n6047), .ZN(U2925) );
  AOI22_X1 U7098 ( .A1(UWORD_REG_2__SCAN_IN), .A2(n6051), .B1(n6079), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n6048) );
  OAI21_X1 U7099 ( .B1(n6081), .B2(n6060), .A(n6048), .ZN(U2926) );
  AOI22_X1 U7100 ( .A1(UWORD_REG_3__SCAN_IN), .A2(n6051), .B1(n6079), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n6049) );
  OAI21_X1 U7101 ( .B1(n6081), .B2(n6968), .A(n6049), .ZN(U2927) );
  AOI22_X1 U7102 ( .A1(UWORD_REG_4__SCAN_IN), .A2(n6051), .B1(n6079), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n6050) );
  OAI21_X1 U7103 ( .B1(n6081), .B2(n6063), .A(n6050), .ZN(U2928) );
  AOI22_X1 U7104 ( .A1(UWORD_REG_5__SCAN_IN), .A2(n6051), .B1(n6079), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n6052) );
  OAI21_X1 U7105 ( .B1(n6081), .B2(n6065), .A(n6052), .ZN(U2929) );
  AOI22_X1 U7106 ( .A1(UWORD_REG_6__SCAN_IN), .A2(n6074), .B1(n6079), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n6053) );
  OAI21_X1 U7107 ( .B1(n6081), .B2(n6067), .A(n6053), .ZN(U2930) );
  AOI22_X1 U7108 ( .A1(UWORD_REG_7__SCAN_IN), .A2(n6074), .B1(n6079), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n6054) );
  OAI21_X1 U7109 ( .B1(n6081), .B2(n6069), .A(n6054), .ZN(U2931) );
  AOI22_X1 U7110 ( .A1(UWORD_REG_13__SCAN_IN), .A2(n6074), .B1(n6079), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n6055) );
  OAI21_X1 U7111 ( .B1(n6081), .B2(n6864), .A(n6055), .ZN(U2937) );
  INV_X1 U7112 ( .A(DATAI_14_), .ZN(n6896) );
  AOI22_X1 U7113 ( .A1(UWORD_REG_14__SCAN_IN), .A2(n6074), .B1(n6079), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n6056) );
  OAI21_X1 U7114 ( .B1(n6081), .B2(n6896), .A(n6056), .ZN(U2938) );
  AOI22_X1 U7115 ( .A1(LWORD_REG_0__SCAN_IN), .A2(n6074), .B1(n6079), .B2(
        EAX_REG_0__SCAN_IN), .ZN(n6057) );
  OAI21_X1 U7116 ( .B1(n6081), .B2(n6861), .A(n6057), .ZN(U2939) );
  AOI22_X1 U7117 ( .A1(LWORD_REG_1__SCAN_IN), .A2(n6074), .B1(n6079), .B2(
        EAX_REG_1__SCAN_IN), .ZN(n6058) );
  OAI21_X1 U7118 ( .B1(n6081), .B2(n6890), .A(n6058), .ZN(U2940) );
  AOI22_X1 U7119 ( .A1(LWORD_REG_2__SCAN_IN), .A2(n6051), .B1(n6079), .B2(
        EAX_REG_2__SCAN_IN), .ZN(n6059) );
  OAI21_X1 U7120 ( .B1(n6081), .B2(n6060), .A(n6059), .ZN(U2941) );
  AOI22_X1 U7121 ( .A1(LWORD_REG_3__SCAN_IN), .A2(n6051), .B1(n6079), .B2(
        EAX_REG_3__SCAN_IN), .ZN(n6061) );
  OAI21_X1 U7122 ( .B1(n6081), .B2(n6968), .A(n6061), .ZN(U2942) );
  AOI22_X1 U7123 ( .A1(LWORD_REG_4__SCAN_IN), .A2(n6051), .B1(n6079), .B2(
        EAX_REG_4__SCAN_IN), .ZN(n6062) );
  OAI21_X1 U7124 ( .B1(n6081), .B2(n6063), .A(n6062), .ZN(U2943) );
  AOI22_X1 U7125 ( .A1(LWORD_REG_5__SCAN_IN), .A2(n6051), .B1(n6079), .B2(
        EAX_REG_5__SCAN_IN), .ZN(n6064) );
  OAI21_X1 U7126 ( .B1(n6081), .B2(n6065), .A(n6064), .ZN(U2944) );
  AOI22_X1 U7127 ( .A1(LWORD_REG_6__SCAN_IN), .A2(n6051), .B1(n6079), .B2(
        EAX_REG_6__SCAN_IN), .ZN(n6066) );
  OAI21_X1 U7128 ( .B1(n6081), .B2(n6067), .A(n6066), .ZN(U2945) );
  AOI22_X1 U7129 ( .A1(LWORD_REG_7__SCAN_IN), .A2(n6051), .B1(n6079), .B2(
        EAX_REG_7__SCAN_IN), .ZN(n6068) );
  OAI21_X1 U7130 ( .B1(n6081), .B2(n6069), .A(n6068), .ZN(U2946) );
  AOI22_X1 U7131 ( .A1(LWORD_REG_9__SCAN_IN), .A2(n6051), .B1(n6079), .B2(
        EAX_REG_9__SCAN_IN), .ZN(n6071) );
  NAND2_X1 U7132 ( .A1(n6075), .A2(DATAI_9_), .ZN(n6070) );
  NAND2_X1 U7133 ( .A1(n6071), .A2(n6070), .ZN(U2948) );
  AOI22_X1 U7134 ( .A1(LWORD_REG_11__SCAN_IN), .A2(n6074), .B1(n6079), .B2(
        EAX_REG_11__SCAN_IN), .ZN(n6073) );
  NAND2_X1 U7135 ( .A1(n6075), .A2(DATAI_11_), .ZN(n6072) );
  NAND2_X1 U7136 ( .A1(n6073), .A2(n6072), .ZN(U2950) );
  AOI22_X1 U7137 ( .A1(LWORD_REG_12__SCAN_IN), .A2(n6074), .B1(n6079), .B2(
        EAX_REG_12__SCAN_IN), .ZN(n6077) );
  NAND2_X1 U7138 ( .A1(n6075), .A2(DATAI_12_), .ZN(n6076) );
  NAND2_X1 U7139 ( .A1(n6077), .A2(n6076), .ZN(U2951) );
  AOI22_X1 U7140 ( .A1(LWORD_REG_13__SCAN_IN), .A2(n6051), .B1(n6079), .B2(
        EAX_REG_13__SCAN_IN), .ZN(n6078) );
  OAI21_X1 U7141 ( .B1(n6081), .B2(n6864), .A(n6078), .ZN(U2952) );
  AOI22_X1 U7142 ( .A1(LWORD_REG_14__SCAN_IN), .A2(n6051), .B1(n6079), .B2(
        EAX_REG_14__SCAN_IN), .ZN(n6080) );
  OAI21_X1 U7143 ( .B1(n6081), .B2(n6896), .A(n6080), .ZN(U2953) );
  AOI22_X1 U7144 ( .A1(n6210), .A2(REIP_REG_11__SCAN_IN), .B1(n6147), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n6088) );
  NAND2_X1 U7145 ( .A1(n6083), .A2(n6082), .ZN(n6085) );
  XNOR2_X1 U7146 ( .A(n5604), .B(n6163), .ZN(n6084) );
  XNOR2_X1 U7147 ( .A(n6085), .B(n6084), .ZN(n6160) );
  AOI22_X1 U7148 ( .A1(n6152), .A2(n6160), .B1(n6134), .B2(n6086), .ZN(n6087)
         );
  OAI211_X1 U7149 ( .C1(n6138), .C2(n6089), .A(n6088), .B(n6087), .ZN(U2975)
         );
  AOI22_X1 U7150 ( .A1(n6210), .A2(REIP_REG_9__SCAN_IN), .B1(n6147), .B2(
        PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n6096) );
  NAND2_X1 U7151 ( .A1(n6091), .A2(n6090), .ZN(n6092) );
  XNOR2_X1 U7152 ( .A(n6093), .B(n6092), .ZN(n6168) );
  AOI22_X1 U7153 ( .A1(n6168), .A2(n6152), .B1(n6134), .B2(n6094), .ZN(n6095)
         );
  OAI211_X1 U7154 ( .C1(n6138), .C2(n6097), .A(n6096), .B(n6095), .ZN(U2977)
         );
  AOI22_X1 U7155 ( .A1(n6210), .A2(REIP_REG_8__SCAN_IN), .B1(n6147), .B2(
        PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n6104) );
  OAI21_X1 U7156 ( .B1(n3209), .B2(n6099), .A(n6098), .ZN(n6101) );
  INV_X1 U7157 ( .A(n6101), .ZN(n6180) );
  AOI22_X1 U7158 ( .A1(n6180), .A2(n6152), .B1(n6134), .B2(n6102), .ZN(n6103)
         );
  OAI211_X1 U7159 ( .C1(n6138), .C2(n6105), .A(n6104), .B(n6103), .ZN(U2978)
         );
  AOI22_X1 U7160 ( .A1(n6210), .A2(REIP_REG_7__SCAN_IN), .B1(n6147), .B2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n6112) );
  OAI21_X1 U7161 ( .B1(n6108), .B2(n6107), .A(n6106), .ZN(n6109) );
  INV_X1 U7162 ( .A(n6109), .ZN(n6185) );
  AOI22_X1 U7163 ( .A1(n6185), .A2(n6152), .B1(n6124), .B2(n6110), .ZN(n6111)
         );
  OAI211_X1 U7164 ( .C1(n6157), .C2(n6113), .A(n6112), .B(n6111), .ZN(U2979)
         );
  AOI22_X1 U7165 ( .A1(n6210), .A2(REIP_REG_6__SCAN_IN), .B1(n6147), .B2(
        PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n6120) );
  OAI21_X1 U7166 ( .B1(n6116), .B2(n6115), .A(n6114), .ZN(n6117) );
  INV_X1 U7167 ( .A(n6117), .ZN(n6192) );
  AOI22_X1 U7168 ( .A1(n6192), .A2(n6152), .B1(n6134), .B2(n6118), .ZN(n6119)
         );
  OAI211_X1 U7169 ( .C1(n6138), .C2(n6121), .A(n6120), .B(n6119), .ZN(U2980)
         );
  AOI22_X1 U7170 ( .A1(n6210), .A2(REIP_REG_5__SCAN_IN), .B1(n6147), .B2(
        PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n6127) );
  INV_X1 U7171 ( .A(n6122), .ZN(n6125) );
  AOI22_X1 U7172 ( .A1(n6125), .A2(n6152), .B1(n6124), .B2(n6123), .ZN(n6126)
         );
  OAI211_X1 U7173 ( .C1(n6157), .C2(n6128), .A(n6127), .B(n6126), .ZN(U2981)
         );
  AOI22_X1 U7174 ( .A1(n6210), .A2(REIP_REG_4__SCAN_IN), .B1(n6147), .B2(
        PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n6136) );
  OAI21_X1 U7175 ( .B1(n6131), .B2(n6129), .A(n3210), .ZN(n6132) );
  INV_X1 U7176 ( .A(n6132), .ZN(n6197) );
  AOI22_X1 U7177 ( .A1(n6197), .A2(n6152), .B1(n6134), .B2(n6133), .ZN(n6135)
         );
  OAI211_X1 U7178 ( .C1(n6138), .C2(n6137), .A(n6136), .B(n6135), .ZN(U2982)
         );
  AOI22_X1 U7179 ( .A1(n6210), .A2(REIP_REG_3__SCAN_IN), .B1(n6147), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n6145) );
  OAI21_X1 U7180 ( .B1(n6139), .B2(n6141), .A(n3216), .ZN(n6142) );
  INV_X1 U7181 ( .A(n6142), .ZN(n6204) );
  AOI22_X1 U7182 ( .A1(n6143), .A2(n4403), .B1(n6204), .B2(n6152), .ZN(n6144)
         );
  OAI211_X1 U7183 ( .C1(n6157), .C2(n6146), .A(n6145), .B(n6144), .ZN(U2983)
         );
  AOI22_X1 U7184 ( .A1(n6210), .A2(REIP_REG_2__SCAN_IN), .B1(n6147), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n6155) );
  INV_X1 U7185 ( .A(n6148), .ZN(n6153) );
  XOR2_X1 U7186 ( .A(n6150), .B(INSTADDRPOINTER_REG_2__SCAN_IN), .Z(n6151) );
  XNOR2_X1 U7187 ( .A(n6149), .B(n6151), .ZN(n6215) );
  AOI22_X1 U7188 ( .A1(n6124), .A2(n6153), .B1(n6215), .B2(n6152), .ZN(n6154)
         );
  OAI211_X1 U7189 ( .C1(n6157), .C2(n6156), .A(n6155), .B(n6154), .ZN(U2984)
         );
  AOI22_X1 U7190 ( .A1(n6158), .A2(n6227), .B1(n6210), .B2(
        REIP_REG_11__SCAN_IN), .ZN(n6162) );
  AOI22_X1 U7191 ( .A1(n6231), .A2(n6160), .B1(n6163), .B2(n6159), .ZN(n6161)
         );
  OAI211_X1 U7192 ( .C1(n6164), .C2(n6163), .A(n6162), .B(n6161), .ZN(U3007)
         );
  INV_X1 U7193 ( .A(n6165), .ZN(n6172) );
  AOI22_X1 U7194 ( .A1(n6166), .A2(n6227), .B1(n6210), .B2(REIP_REG_9__SCAN_IN), .ZN(n6170) );
  AOI22_X1 U7195 ( .A1(n6168), .A2(n6231), .B1(n6167), .B2(n6171), .ZN(n6169)
         );
  OAI211_X1 U7196 ( .C1(n6172), .C2(n6171), .A(n6170), .B(n6169), .ZN(U3009)
         );
  AOI211_X1 U7197 ( .C1(n6174), .C2(n6816), .A(n6173), .B(n6188), .ZN(n6179)
         );
  OAI22_X1 U7198 ( .A1(n6177), .A2(n6176), .B1(n6499), .B2(n6175), .ZN(n6178)
         );
  AOI211_X1 U7199 ( .C1(n6180), .C2(n6231), .A(n6179), .B(n6178), .ZN(n6181)
         );
  OAI21_X1 U7200 ( .B1(n6182), .B2(n6816), .A(n6181), .ZN(U3010) );
  AOI22_X1 U7201 ( .A1(n6227), .A2(n6183), .B1(n6210), .B2(REIP_REG_7__SCAN_IN), .ZN(n6187) );
  AOI22_X1 U7202 ( .A1(n6185), .A2(n6231), .B1(INSTADDRPOINTER_REG_7__SCAN_IN), 
        .B2(n6184), .ZN(n6186) );
  OAI211_X1 U7203 ( .C1(INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n6188), .A(n6187), 
        .B(n6186), .ZN(U3011) );
  INV_X1 U7204 ( .A(n6189), .ZN(n6195) );
  AOI22_X1 U7205 ( .A1(n6227), .A2(n6190), .B1(n6210), .B2(REIP_REG_6__SCAN_IN), .ZN(n6194) );
  AOI22_X1 U7206 ( .A1(n6192), .A2(n6231), .B1(n6191), .B2(n6752), .ZN(n6193)
         );
  OAI211_X1 U7207 ( .C1(n6195), .C2(n6752), .A(n6194), .B(n6193), .ZN(U3012)
         );
  AOI21_X1 U7208 ( .B1(n6212), .B2(n6214), .A(n6216), .ZN(n6208) );
  AOI222_X1 U7209 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6210), .B1(n6231), .B2(
        n6197), .C1(n6196), .C2(n6227), .ZN(n6201) );
  NOR2_X1 U7210 ( .A1(n6214), .A2(n6198), .ZN(n6205) );
  OAI211_X1 U7211 ( .C1(INSTADDRPOINTER_REG_3__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .A(n6205), .B(n6199), .ZN(n6200) );
  OAI211_X1 U7212 ( .C1(n6208), .C2(n6202), .A(n6201), .B(n6200), .ZN(U3014)
         );
  AOI22_X1 U7213 ( .A1(n6227), .A2(n6203), .B1(n6210), .B2(REIP_REG_3__SCAN_IN), .ZN(n6207) );
  AOI22_X1 U7214 ( .A1(n6205), .A2(n6802), .B1(n6204), .B2(n6231), .ZN(n6206)
         );
  OAI211_X1 U7215 ( .C1(n6208), .C2(n6802), .A(n6207), .B(n6206), .ZN(U3015)
         );
  INV_X1 U7216 ( .A(n6209), .ZN(n6211) );
  AOI22_X1 U7217 ( .A1(n6227), .A2(n6211), .B1(n6210), .B2(REIP_REG_2__SCAN_IN), .ZN(n6221) );
  OAI221_X1 U7218 ( .B1(n6214), .B2(n6213), .C1(n6214), .C2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .A(n6212), .ZN(n6220) );
  AOI22_X1 U7219 ( .A1(n6216), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .B1(n6231), 
        .B2(n6215), .ZN(n6219) );
  NAND3_X1 U7220 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n4230), .A3(n6217), 
        .ZN(n6218) );
  NAND4_X1 U7221 ( .A1(n6221), .A2(n6220), .A3(n6219), .A4(n6218), .ZN(U3016)
         );
  INV_X1 U7222 ( .A(n6222), .ZN(n6232) );
  AOI21_X1 U7223 ( .B1(n6224), .B2(INSTADDRPOINTER_REG_0__SCAN_IN), .A(n6223), 
        .ZN(n6229) );
  AOI21_X1 U7224 ( .B1(n6227), .B2(n6226), .A(n6225), .ZN(n6228) );
  OAI21_X1 U7225 ( .B1(n6229), .B2(INSTADDRPOINTER_REG_1__SCAN_IN), .A(n6228), 
        .ZN(n6230) );
  AOI21_X1 U7226 ( .B1(n6232), .B2(n6231), .A(n6230), .ZN(n6233) );
  OAI21_X1 U7227 ( .B1(n6235), .B2(n6234), .A(n6233), .ZN(U3017) );
  NOR2_X1 U7228 ( .A1(n6237), .A2(n6236), .ZN(U3019) );
  NOR2_X1 U7229 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6238), .ZN(n6260)
         );
  NAND3_X1 U7230 ( .A1(n6239), .A2(n6308), .A3(n6441), .ZN(n6240) );
  OAI21_X1 U7231 ( .B1(n6242), .B2(n6275), .A(n6240), .ZN(n6261) );
  AOI22_X1 U7232 ( .A1(n6380), .A2(n6260), .B1(n6383), .B2(n6261), .ZN(n6247)
         );
  OAI21_X1 U7233 ( .B1(n6241), .B2(n6262), .A(n6316), .ZN(n6243) );
  AOI21_X1 U7234 ( .B1(n6243), .B2(n6242), .A(STATE2_REG_3__SCAN_IN), .ZN(
        n6245) );
  AOI22_X1 U7235 ( .A1(n6263), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n6381), 
        .B2(n6262), .ZN(n6246) );
  OAI211_X1 U7236 ( .C1(n6324), .C2(n6266), .A(n6247), .B(n6246), .ZN(U3036)
         );
  AOI22_X1 U7237 ( .A1(n3193), .A2(n6260), .B1(n6396), .B2(n6261), .ZN(n6249)
         );
  AOI22_X1 U7238 ( .A1(n6263), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n6262), 
        .B2(n6387), .ZN(n6248) );
  OAI211_X1 U7239 ( .C1(n6266), .C2(n6327), .A(n6249), .B(n6248), .ZN(U3037)
         );
  AOI22_X1 U7240 ( .A1(n6401), .A2(n6260), .B1(n6402), .B2(n6261), .ZN(n6251)
         );
  AOI22_X1 U7241 ( .A1(n6263), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n6262), 
        .B2(n6328), .ZN(n6250) );
  OAI211_X1 U7242 ( .C1(n6266), .C2(n6331), .A(n6251), .B(n6250), .ZN(U3038)
         );
  AOI22_X1 U7243 ( .A1(n6407), .A2(n6260), .B1(n6408), .B2(n6261), .ZN(n6253)
         );
  AOI22_X1 U7244 ( .A1(n6263), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n6262), 
        .B2(n6332), .ZN(n6252) );
  OAI211_X1 U7245 ( .C1(n6266), .C2(n6335), .A(n6253), .B(n6252), .ZN(U3039)
         );
  AOI22_X1 U7246 ( .A1(n6358), .A2(n6260), .B1(n6360), .B2(n6261), .ZN(n6255)
         );
  AOI22_X1 U7247 ( .A1(n6263), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n6262), 
        .B2(n6336), .ZN(n6254) );
  OAI211_X1 U7248 ( .C1(n6266), .C2(n6339), .A(n6255), .B(n6254), .ZN(U3040)
         );
  AOI22_X1 U7249 ( .A1(n6414), .A2(n6261), .B1(n6413), .B2(n6260), .ZN(n6257)
         );
  AOI22_X1 U7250 ( .A1(n6263), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n6262), 
        .B2(n6340), .ZN(n6256) );
  OAI211_X1 U7251 ( .C1(n6266), .C2(n6343), .A(n6257), .B(n6256), .ZN(U3041)
         );
  AOI22_X1 U7252 ( .A1(n6421), .A2(n6260), .B1(n6423), .B2(n6261), .ZN(n6259)
         );
  AOI22_X1 U7253 ( .A1(n6263), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n6262), 
        .B2(n6344), .ZN(n6258) );
  OAI211_X1 U7254 ( .C1(n6266), .C2(n6347), .A(n6259), .B(n6258), .ZN(U3042)
         );
  AOI22_X1 U7255 ( .A1(n6373), .A2(n6261), .B1(n6369), .B2(n6260), .ZN(n6265)
         );
  AOI22_X1 U7256 ( .A1(n6263), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n6262), 
        .B2(n6351), .ZN(n6264) );
  OAI211_X1 U7257 ( .C1(n6266), .C2(n6355), .A(n6265), .B(n6264), .ZN(U3043)
         );
  INV_X1 U7258 ( .A(n6279), .ZN(n6273) );
  OR3_X1 U7259 ( .A1(n6269), .A2(n6268), .A3(n6267), .ZN(n6271) );
  NOR2_X1 U7260 ( .A1(n6430), .A2(n6281), .ZN(n6301) );
  INV_X1 U7261 ( .A(n6301), .ZN(n6270) );
  NAND2_X1 U7262 ( .A1(n6271), .A2(n6270), .ZN(n6278) );
  OAI21_X1 U7263 ( .B1(n6273), .B2(n6278), .A(n6272), .ZN(n6274) );
  INV_X1 U7264 ( .A(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n6805) );
  NAND2_X1 U7265 ( .A1(n6277), .A2(n6276), .ZN(n6314) );
  AOI22_X1 U7266 ( .A1(n6350), .A2(n6382), .B1(n6380), .B2(n6301), .ZN(n6283)
         );
  NAND2_X1 U7267 ( .A1(n6279), .A2(n6278), .ZN(n6280) );
  OAI21_X1 U7268 ( .B1(n6281), .B2(n4463), .A(n6280), .ZN(n6303) );
  AOI22_X1 U7269 ( .A1(n6303), .A2(n6383), .B1(n6381), .B2(n6302), .ZN(n6282)
         );
  OAI211_X1 U7270 ( .C1(n6306), .C2(n6805), .A(n6283), .B(n6282), .ZN(U3060)
         );
  INV_X1 U7271 ( .A(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n6286) );
  AOI22_X1 U7272 ( .A1(n6350), .A2(n6394), .B1(n3193), .B2(n6301), .ZN(n6285)
         );
  AOI22_X1 U7273 ( .A1(n6303), .A2(n6396), .B1(n6387), .B2(n6302), .ZN(n6284)
         );
  OAI211_X1 U7274 ( .C1(n6306), .C2(n6286), .A(n6285), .B(n6284), .ZN(U3061)
         );
  INV_X1 U7275 ( .A(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n6289) );
  AOI22_X1 U7276 ( .A1(n6350), .A2(n6400), .B1(n6401), .B2(n6301), .ZN(n6288)
         );
  AOI22_X1 U7277 ( .A1(n6303), .A2(n6402), .B1(n6328), .B2(n6302), .ZN(n6287)
         );
  OAI211_X1 U7278 ( .C1(n6306), .C2(n6289), .A(n6288), .B(n6287), .ZN(U3062)
         );
  INV_X1 U7279 ( .A(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n6724) );
  AOI22_X1 U7280 ( .A1(n6350), .A2(n6406), .B1(n6407), .B2(n6301), .ZN(n6291)
         );
  AOI22_X1 U7281 ( .A1(n6303), .A2(n6408), .B1(n6332), .B2(n6302), .ZN(n6290)
         );
  OAI211_X1 U7282 ( .C1(n6306), .C2(n6724), .A(n6291), .B(n6290), .ZN(U3063)
         );
  INV_X1 U7283 ( .A(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n6294) );
  AOI22_X1 U7284 ( .A1(n6350), .A2(n6359), .B1(n6358), .B2(n6301), .ZN(n6293)
         );
  AOI22_X1 U7285 ( .A1(n6303), .A2(n6360), .B1(n6336), .B2(n6302), .ZN(n6292)
         );
  OAI211_X1 U7286 ( .C1(n6306), .C2(n6294), .A(n6293), .B(n6292), .ZN(U3064)
         );
  INV_X1 U7287 ( .A(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n6297) );
  AOI22_X1 U7288 ( .A1(n6350), .A2(n6412), .B1(n6413), .B2(n6301), .ZN(n6296)
         );
  AOI22_X1 U7289 ( .A1(n6303), .A2(n6414), .B1(n6340), .B2(n6302), .ZN(n6295)
         );
  OAI211_X1 U7290 ( .C1(n6306), .C2(n6297), .A(n6296), .B(n6295), .ZN(U3065)
         );
  INV_X1 U7291 ( .A(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n6300) );
  AOI22_X1 U7292 ( .A1(n6350), .A2(n6418), .B1(n6421), .B2(n6301), .ZN(n6299)
         );
  AOI22_X1 U7293 ( .A1(n6303), .A2(n6423), .B1(n6344), .B2(n6302), .ZN(n6298)
         );
  OAI211_X1 U7294 ( .C1(n6306), .C2(n6300), .A(n6299), .B(n6298), .ZN(U3066)
         );
  INV_X1 U7295 ( .A(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n6763) );
  AOI22_X1 U7296 ( .A1(n6350), .A2(n6371), .B1(n6369), .B2(n6301), .ZN(n6305)
         );
  AOI22_X1 U7297 ( .A1(n6303), .A2(n6373), .B1(n6351), .B2(n6302), .ZN(n6304)
         );
  OAI211_X1 U7298 ( .C1(n6306), .C2(n6763), .A(n6305), .B(n6304), .ZN(U3067)
         );
  NOR2_X1 U7299 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6307), .ZN(n6348)
         );
  NAND3_X1 U7300 ( .A1(n6309), .A2(n6308), .A3(n6441), .ZN(n6310) );
  OAI21_X1 U7301 ( .B1(n6312), .B2(n6311), .A(n6310), .ZN(n6349) );
  AOI22_X1 U7302 ( .A1(n6380), .A2(n6348), .B1(n6383), .B2(n6349), .ZN(n6323)
         );
  NAND3_X1 U7303 ( .A1(n6377), .A2(n6314), .A3(n6313), .ZN(n6317) );
  AOI21_X1 U7304 ( .B1(n6317), .B2(n6316), .A(n6315), .ZN(n6321) );
  OAI211_X1 U7305 ( .C1(n6348), .C2(n6547), .A(n6318), .B(n6441), .ZN(n6319)
         );
  AOI22_X1 U7306 ( .A1(n6352), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n6381), 
        .B2(n6350), .ZN(n6322) );
  OAI211_X1 U7307 ( .C1(n6324), .C2(n6377), .A(n6323), .B(n6322), .ZN(U3068)
         );
  AOI22_X1 U7308 ( .A1(n3193), .A2(n6348), .B1(n6396), .B2(n6349), .ZN(n6326)
         );
  AOI22_X1 U7309 ( .A1(n6352), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n6387), 
        .B2(n6350), .ZN(n6325) );
  OAI211_X1 U7310 ( .C1(n6327), .C2(n6377), .A(n6326), .B(n6325), .ZN(U3069)
         );
  AOI22_X1 U7311 ( .A1(n6401), .A2(n6348), .B1(n6402), .B2(n6349), .ZN(n6330)
         );
  AOI22_X1 U7312 ( .A1(n6352), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n6328), 
        .B2(n6350), .ZN(n6329) );
  OAI211_X1 U7313 ( .C1(n6331), .C2(n6377), .A(n6330), .B(n6329), .ZN(U3070)
         );
  AOI22_X1 U7314 ( .A1(n6407), .A2(n6348), .B1(n6408), .B2(n6349), .ZN(n6334)
         );
  AOI22_X1 U7315 ( .A1(n6352), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n6332), 
        .B2(n6350), .ZN(n6333) );
  OAI211_X1 U7316 ( .C1(n6335), .C2(n6377), .A(n6334), .B(n6333), .ZN(U3071)
         );
  AOI22_X1 U7317 ( .A1(n6358), .A2(n6348), .B1(n6360), .B2(n6349), .ZN(n6338)
         );
  AOI22_X1 U7318 ( .A1(n6352), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n6336), 
        .B2(n6350), .ZN(n6337) );
  OAI211_X1 U7319 ( .C1(n6339), .C2(n6377), .A(n6338), .B(n6337), .ZN(U3072)
         );
  AOI22_X1 U7320 ( .A1(n6414), .A2(n6349), .B1(n6413), .B2(n6348), .ZN(n6342)
         );
  AOI22_X1 U7321 ( .A1(n6352), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n6340), 
        .B2(n6350), .ZN(n6341) );
  OAI211_X1 U7322 ( .C1(n6343), .C2(n6377), .A(n6342), .B(n6341), .ZN(U3073)
         );
  AOI22_X1 U7323 ( .A1(n6421), .A2(n6348), .B1(n6423), .B2(n6349), .ZN(n6346)
         );
  AOI22_X1 U7324 ( .A1(n6352), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n6344), 
        .B2(n6350), .ZN(n6345) );
  OAI211_X1 U7325 ( .C1(n6347), .C2(n6377), .A(n6346), .B(n6345), .ZN(U3074)
         );
  AOI22_X1 U7326 ( .A1(n6373), .A2(n6349), .B1(n6369), .B2(n6348), .ZN(n6354)
         );
  AOI22_X1 U7327 ( .A1(n6352), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n6351), 
        .B2(n6350), .ZN(n6353) );
  OAI211_X1 U7328 ( .C1(n6355), .C2(n6377), .A(n6354), .B(n6353), .ZN(U3075)
         );
  AOI22_X1 U7329 ( .A1(n6400), .A2(n6370), .B1(n6401), .B2(n6368), .ZN(n6357)
         );
  AOI22_X1 U7330 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n6374), .B1(n6402), 
        .B2(n6372), .ZN(n6356) );
  OAI211_X1 U7331 ( .C1(n6405), .C2(n6377), .A(n6357), .B(n6356), .ZN(U3078)
         );
  AOI22_X1 U7332 ( .A1(n6359), .A2(n6370), .B1(n6358), .B2(n6368), .ZN(n6362)
         );
  AOI22_X1 U7333 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n6374), .B1(n6360), 
        .B2(n6372), .ZN(n6361) );
  OAI211_X1 U7334 ( .C1(n6363), .C2(n6377), .A(n6362), .B(n6361), .ZN(U3080)
         );
  AOI22_X1 U7335 ( .A1(n6412), .A2(n6370), .B1(n6413), .B2(n6368), .ZN(n6365)
         );
  AOI22_X1 U7336 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n6374), .B1(n6414), 
        .B2(n6372), .ZN(n6364) );
  OAI211_X1 U7337 ( .C1(n6417), .C2(n6377), .A(n6365), .B(n6364), .ZN(U3081)
         );
  AOI22_X1 U7338 ( .A1(n6418), .A2(n6370), .B1(n6421), .B2(n6368), .ZN(n6367)
         );
  AOI22_X1 U7339 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n6374), .B1(n6423), 
        .B2(n6372), .ZN(n6366) );
  OAI211_X1 U7340 ( .C1(n6428), .C2(n6377), .A(n6367), .B(n6366), .ZN(U3082)
         );
  AOI22_X1 U7341 ( .A1(n6371), .A2(n6370), .B1(n6369), .B2(n6368), .ZN(n6376)
         );
  AOI22_X1 U7342 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n6374), .B1(n6373), 
        .B2(n6372), .ZN(n6375) );
  OAI211_X1 U7343 ( .C1(n6378), .C2(n6377), .A(n6376), .B(n6375), .ZN(U3083)
         );
  INV_X1 U7344 ( .A(n6379), .ZN(n6393) );
  INV_X1 U7345 ( .A(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n6863) );
  AOI22_X1 U7346 ( .A1(n6388), .A2(n6381), .B1(n6380), .B2(n6386), .ZN(n6385)
         );
  AOI22_X1 U7347 ( .A1(n6390), .A2(n6383), .B1(n6382), .B2(n6389), .ZN(n6384)
         );
  OAI211_X1 U7348 ( .C1(n6393), .C2(n6863), .A(n6385), .B(n6384), .ZN(U3092)
         );
  INV_X1 U7349 ( .A(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n6832) );
  AOI22_X1 U7350 ( .A1(n6388), .A2(n6387), .B1(n3193), .B2(n6386), .ZN(n6392)
         );
  AOI22_X1 U7351 ( .A1(n6390), .A2(n6396), .B1(n6394), .B2(n6389), .ZN(n6391)
         );
  OAI211_X1 U7352 ( .C1(n6393), .C2(n6832), .A(n6392), .B(n6391), .ZN(U3093)
         );
  AOI22_X1 U7353 ( .A1(n3193), .A2(n6420), .B1(n6419), .B2(n6394), .ZN(n6398)
         );
  AOI22_X1 U7354 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n6424), .B1(n6396), 
        .B2(n6422), .ZN(n6397) );
  OAI211_X1 U7355 ( .C1(n6399), .C2(n6427), .A(n6398), .B(n6397), .ZN(U3109)
         );
  AOI22_X1 U7356 ( .A1(n6401), .A2(n6420), .B1(n6419), .B2(n6400), .ZN(n6404)
         );
  AOI22_X1 U7357 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n6424), .B1(n6402), 
        .B2(n6422), .ZN(n6403) );
  OAI211_X1 U7358 ( .C1(n6405), .C2(n6427), .A(n6404), .B(n6403), .ZN(U3110)
         );
  AOI22_X1 U7359 ( .A1(n6407), .A2(n6420), .B1(n6419), .B2(n6406), .ZN(n6410)
         );
  AOI22_X1 U7360 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6424), .B1(n6408), 
        .B2(n6422), .ZN(n6409) );
  OAI211_X1 U7361 ( .C1(n6411), .C2(n6427), .A(n6410), .B(n6409), .ZN(U3111)
         );
  AOI22_X1 U7362 ( .A1(n6413), .A2(n6420), .B1(n6419), .B2(n6412), .ZN(n6416)
         );
  AOI22_X1 U7363 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6424), .B1(n6414), 
        .B2(n6422), .ZN(n6415) );
  OAI211_X1 U7364 ( .C1(n6417), .C2(n6427), .A(n6416), .B(n6415), .ZN(U3113)
         );
  AOI22_X1 U7365 ( .A1(n6421), .A2(n6420), .B1(n6419), .B2(n6418), .ZN(n6426)
         );
  AOI22_X1 U7366 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n6424), .B1(n6423), 
        .B2(n6422), .ZN(n6425) );
  OAI211_X1 U7367 ( .C1(n6428), .C2(n6427), .A(n6426), .B(n6425), .ZN(U3114)
         );
  AOI211_X1 U7368 ( .C1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n6431), .A(n6430), .B(n6429), .ZN(n6434) );
  INV_X1 U7369 ( .A(n6434), .ZN(n6437) );
  OAI22_X1 U7370 ( .A1(n6434), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(n6433), .B2(n6432), .ZN(n6435) );
  OAI21_X1 U7371 ( .B1(n6437), .B2(n6436), .A(n6435), .ZN(n6438) );
  AOI222_X1 U7372 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n6439), .B1(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n6438), .C1(n6439), .C2(n6438), 
        .ZN(n6440) );
  AOI222_X1 U7373 ( .A1(n6442), .A2(n6441), .B1(n6442), .B2(n6440), .C1(n6441), 
        .C2(n6440), .ZN(n6443) );
  NOR2_X1 U7374 ( .A1(n6443), .A2(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6450)
         );
  NOR2_X1 U7375 ( .A1(FLUSH_REG_SCAN_IN), .A2(MORE_REG_SCAN_IN), .ZN(n6446) );
  OAI211_X1 U7376 ( .C1(n6447), .C2(n6446), .A(n6445), .B(n6444), .ZN(n6448)
         );
  NOR3_X1 U7377 ( .A1(n6450), .A2(n6449), .A3(n6448), .ZN(n6462) );
  OAI21_X1 U7378 ( .B1(n6452), .B2(n6451), .A(STATE2_REG_2__SCAN_IN), .ZN(
        n6453) );
  AOI221_X1 U7379 ( .B1(n6736), .B2(n6567), .C1(n4324), .C2(n6567), .A(n6453), 
        .ZN(n6455) );
  AOI21_X1 U7380 ( .B1(n6471), .B2(n6548), .A(n6455), .ZN(n6454) );
  INV_X1 U7381 ( .A(n6454), .ZN(n6458) );
  OAI221_X1 U7382 ( .B1(n6567), .B2(n6462), .C1(n6567), .C2(n6736), .A(n6455), 
        .ZN(n6546) );
  OAI21_X1 U7383 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n4324), .A(n6546), .ZN(
        n6465) );
  NOR2_X1 U7384 ( .A1(n6456), .A2(n6465), .ZN(n6457) );
  MUX2_X1 U7385 ( .A(n6458), .B(n6457), .S(STATE2_REG_0__SCAN_IN), .Z(n6460)
         );
  OAI211_X1 U7386 ( .C1(n6462), .C2(n6461), .A(n6460), .B(n6459), .ZN(U3148)
         );
  INV_X1 U7387 ( .A(n6546), .ZN(n6470) );
  AOI21_X1 U7388 ( .B1(n6464), .B2(n4324), .A(n6463), .ZN(n6469) );
  NAND3_X1 U7389 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6466), .A3(n6465), .ZN(
        n6467) );
  OAI211_X1 U7390 ( .C1(n6470), .C2(n6469), .A(n6468), .B(n6467), .ZN(U3149)
         );
  INV_X1 U7391 ( .A(n6471), .ZN(n6566) );
  OAI211_X1 U7392 ( .C1(STATE2_REG_2__SCAN_IN), .C2(n4324), .A(n6545), .B(
        n6566), .ZN(n6473) );
  OAI21_X1 U7393 ( .B1(n6474), .B2(n6473), .A(n6472), .ZN(U3150) );
  AND2_X1 U7394 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6540), .ZN(U3151) );
  AND2_X1 U7395 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6540), .ZN(U3152) );
  AND2_X1 U7396 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6540), .ZN(U3153) );
  AND2_X1 U7397 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6540), .ZN(U3154) );
  AND2_X1 U7398 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6540), .ZN(U3155) );
  AND2_X1 U7399 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6540), .ZN(U3156) );
  AND2_X1 U7400 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6540), .ZN(U3157) );
  AND2_X1 U7401 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6540), .ZN(U3158) );
  INV_X1 U7402 ( .A(DATAWIDTH_REG_23__SCAN_IN), .ZN(n6740) );
  NOR2_X1 U7403 ( .A1(n6544), .A2(n6740), .ZN(U3159) );
  AND2_X1 U7404 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6540), .ZN(U3160) );
  INV_X1 U7405 ( .A(DATAWIDTH_REG_21__SCAN_IN), .ZN(n6767) );
  NOR2_X1 U7406 ( .A1(n6544), .A2(n6767), .ZN(U3161) );
  INV_X1 U7407 ( .A(DATAWIDTH_REG_20__SCAN_IN), .ZN(n6909) );
  NOR2_X1 U7408 ( .A1(n6544), .A2(n6909), .ZN(U3162) );
  AND2_X1 U7409 ( .A1(n6540), .A2(DATAWIDTH_REG_19__SCAN_IN), .ZN(U3163) );
  INV_X1 U7410 ( .A(DATAWIDTH_REG_18__SCAN_IN), .ZN(n6817) );
  NOR2_X1 U7411 ( .A1(n6544), .A2(n6817), .ZN(U3164) );
  AND2_X1 U7412 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n6540), .ZN(U3165) );
  AND2_X1 U7413 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6540), .ZN(U3166) );
  INV_X1 U7414 ( .A(DATAWIDTH_REG_15__SCAN_IN), .ZN(n6875) );
  NOR2_X1 U7415 ( .A1(n6544), .A2(n6875), .ZN(U3167) );
  AND2_X1 U7416 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6540), .ZN(U3168) );
  INV_X1 U7417 ( .A(DATAWIDTH_REG_13__SCAN_IN), .ZN(n6899) );
  NOR2_X1 U7418 ( .A1(n6544), .A2(n6899), .ZN(U3169) );
  AND2_X1 U7419 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(n6540), .ZN(U3170) );
  AND2_X1 U7420 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n6540), .ZN(U3171) );
  AND2_X1 U7421 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n6540), .ZN(U3172) );
  AND2_X1 U7422 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6540), .ZN(U3173) );
  INV_X1 U7423 ( .A(DATAWIDTH_REG_8__SCAN_IN), .ZN(n6867) );
  NOR2_X1 U7424 ( .A1(n6544), .A2(n6867), .ZN(U3174) );
  AND2_X1 U7425 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n6540), .ZN(U3175) );
  AND2_X1 U7426 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6540), .ZN(U3176) );
  AND2_X1 U7427 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(n6540), .ZN(U3177) );
  INV_X1 U7428 ( .A(DATAWIDTH_REG_4__SCAN_IN), .ZN(n6850) );
  NOR2_X1 U7429 ( .A1(n6544), .A2(n6850), .ZN(U3178) );
  AND2_X1 U7430 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n6540), .ZN(U3179) );
  AND2_X1 U7431 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6540), .ZN(U3180) );
  NOR2_X1 U7432 ( .A1(n6482), .A2(n6475), .ZN(n6483) );
  AOI22_X1 U7433 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .B1(
        STATE_REG_2__SCAN_IN), .B2(HOLD), .ZN(n6490) );
  AND2_X1 U7434 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n6479) );
  INV_X1 U7435 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6477) );
  INV_X1 U7436 ( .A(NA_N), .ZN(n6484) );
  AOI221_X1 U7437 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .C1(
        n6484), .C2(STATE_REG_2__SCAN_IN), .A(STATE_REG_0__SCAN_IN), .ZN(n6487) );
  AOI221_X1 U7438 ( .B1(n6479), .B2(n6573), .C1(n6477), .C2(n6573), .A(n6487), 
        .ZN(n6476) );
  OAI21_X1 U7439 ( .B1(n6483), .B2(n6490), .A(n6476), .ZN(U3181) );
  NOR2_X1 U7440 ( .A1(n6798), .A2(n6477), .ZN(n6485) );
  NAND2_X1 U7441 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n6478) );
  OAI21_X1 U7442 ( .B1(n6485), .B2(n6479), .A(n6478), .ZN(n6480) );
  OAI211_X1 U7443 ( .C1(n6482), .C2(n4324), .A(n6481), .B(n6480), .ZN(U3182)
         );
  AOI21_X1 U7444 ( .B1(n6485), .B2(n6484), .A(n6483), .ZN(n6489) );
  AOI221_X1 U7445 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n4324), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6486) );
  AOI221_X1 U7446 ( .B1(STATE_REG_2__SCAN_IN), .B2(HOLD), .C1(n6486), .C2(HOLD), .A(n6798), .ZN(n6488) );
  OAI22_X1 U7447 ( .A1(n6490), .A2(n6489), .B1(n6488), .B2(n6487), .ZN(U3183)
         );
  NAND2_X1 U7448 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6575), .ZN(n6536) );
  AOI22_X1 U7449 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6534), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n6573), .ZN(n6491) );
  OAI21_X1 U7450 ( .B1(n6555), .B2(n6536), .A(n6491), .ZN(U3184) );
  INV_X1 U7451 ( .A(n6536), .ZN(n6531) );
  AOI22_X1 U7452 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6531), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n6573), .ZN(n6492) );
  OAI21_X1 U7453 ( .B1(n6801), .B2(n6533), .A(n6492), .ZN(U3185) );
  AOI22_X1 U7454 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6534), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n6573), .ZN(n6493) );
  OAI21_X1 U7455 ( .B1(n6801), .B2(n6536), .A(n6493), .ZN(U3186) );
  AOI22_X1 U7456 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6531), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n6573), .ZN(n6494) );
  OAI21_X1 U7457 ( .B1(n4642), .B2(n6533), .A(n6494), .ZN(U3187) );
  AOI22_X1 U7458 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6534), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n6573), .ZN(n6495) );
  OAI21_X1 U7459 ( .B1(n4642), .B2(n6536), .A(n6495), .ZN(U3188) );
  INV_X1 U7460 ( .A(ADDRESS_REG_5__SCAN_IN), .ZN(n6769) );
  INV_X1 U7461 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6498) );
  OAI222_X1 U7462 ( .A1(n6536), .A2(n6496), .B1(n6769), .B2(n6575), .C1(n6498), 
        .C2(n6533), .ZN(U3189) );
  AOI22_X1 U7463 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6534), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n6573), .ZN(n6497) );
  OAI21_X1 U7464 ( .B1(n6498), .B2(n6536), .A(n6497), .ZN(U3190) );
  INV_X1 U7465 ( .A(REIP_REG_9__SCAN_IN), .ZN(n6500) );
  INV_X1 U7466 ( .A(ADDRESS_REG_7__SCAN_IN), .ZN(n6846) );
  OAI222_X1 U7467 ( .A1(n6533), .A2(n6500), .B1(n6846), .B2(n6575), .C1(n6499), 
        .C2(n6536), .ZN(U3191) );
  INV_X1 U7468 ( .A(ADDRESS_REG_8__SCAN_IN), .ZN(n6812) );
  OAI222_X1 U7469 ( .A1(n6533), .A2(n6501), .B1(n6812), .B2(n6575), .C1(n6500), 
        .C2(n6536), .ZN(U3192) );
  INV_X1 U7470 ( .A(ADDRESS_REG_9__SCAN_IN), .ZN(n6782) );
  OAI222_X1 U7471 ( .A1(n6536), .A2(n6501), .B1(n6782), .B2(n6575), .C1(n6503), 
        .C2(n6533), .ZN(U3193) );
  AOI22_X1 U7472 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6534), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n6573), .ZN(n6502) );
  OAI21_X1 U7473 ( .B1(n6503), .B2(n6536), .A(n6502), .ZN(U3194) );
  AOI22_X1 U7474 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6531), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n6573), .ZN(n6504) );
  OAI21_X1 U7475 ( .B1(n6505), .B2(n6533), .A(n6504), .ZN(U3195) );
  AOI22_X1 U7476 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6531), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n6573), .ZN(n6506) );
  OAI21_X1 U7477 ( .B1(n6507), .B2(n6533), .A(n6506), .ZN(U3196) );
  AOI22_X1 U7478 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6531), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6573), .ZN(n6508) );
  OAI21_X1 U7479 ( .B1(n6811), .B2(n6533), .A(n6508), .ZN(U3197) );
  AOI22_X1 U7480 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6531), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(n6573), .ZN(n6509) );
  OAI21_X1 U7481 ( .B1(n5619), .B2(n6533), .A(n6509), .ZN(U3198) );
  AOI22_X1 U7482 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6534), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n6573), .ZN(n6510) );
  OAI21_X1 U7483 ( .B1(n5619), .B2(n6536), .A(n6510), .ZN(U3199) );
  INV_X1 U7484 ( .A(REIP_REG_17__SCAN_IN), .ZN(n6511) );
  INV_X1 U7485 ( .A(ADDRESS_REG_16__SCAN_IN), .ZN(n6877) );
  OAI222_X1 U7486 ( .A1(n6536), .A2(n6511), .B1(n6877), .B2(n6575), .C1(n6513), 
        .C2(n6533), .ZN(U3200) );
  AOI22_X1 U7487 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6534), .B1(
        ADDRESS_REG_17__SCAN_IN), .B2(n6573), .ZN(n6512) );
  OAI21_X1 U7488 ( .B1(n6513), .B2(n6536), .A(n6512), .ZN(U3201) );
  INV_X1 U7489 ( .A(REIP_REG_19__SCAN_IN), .ZN(n6515) );
  AOI22_X1 U7490 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6534), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n6573), .ZN(n6514) );
  OAI21_X1 U7491 ( .B1(n6515), .B2(n6536), .A(n6514), .ZN(U3202) );
  AOI22_X1 U7492 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6531), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(n6573), .ZN(n6516) );
  OAI21_X1 U7493 ( .B1(n6517), .B2(n6533), .A(n6516), .ZN(U3203) );
  AOI22_X1 U7494 ( .A1(REIP_REG_21__SCAN_IN), .A2(n6531), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n6573), .ZN(n6518) );
  OAI21_X1 U7495 ( .B1(n6521), .B2(n6533), .A(n6518), .ZN(U3204) );
  INV_X1 U7496 ( .A(ADDRESS_REG_21__SCAN_IN), .ZN(n6520) );
  OAI222_X1 U7497 ( .A1(n6536), .A2(n6521), .B1(n6520), .B2(n6575), .C1(n6519), 
        .C2(n6533), .ZN(U3205) );
  AOI22_X1 U7498 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6531), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n6573), .ZN(n6522) );
  OAI21_X1 U7499 ( .B1(n6523), .B2(n6533), .A(n6522), .ZN(U3206) );
  INV_X1 U7500 ( .A(ADDRESS_REG_23__SCAN_IN), .ZN(n6524) );
  OAI222_X1 U7501 ( .A1(n6533), .A2(n6525), .B1(n6524), .B2(n6575), .C1(n6523), 
        .C2(n6536), .ZN(U3207) );
  INV_X1 U7502 ( .A(ADDRESS_REG_24__SCAN_IN), .ZN(n6709) );
  OAI222_X1 U7503 ( .A1(n6536), .A2(n6525), .B1(n6709), .B2(n6575), .C1(n6526), 
        .C2(n6533), .ZN(U3208) );
  INV_X1 U7504 ( .A(ADDRESS_REG_25__SCAN_IN), .ZN(n6882) );
  OAI222_X1 U7505 ( .A1(n6536), .A2(n6526), .B1(n6882), .B2(n6575), .C1(n6528), 
        .C2(n6533), .ZN(U3209) );
  AOI22_X1 U7506 ( .A1(REIP_REG_28__SCAN_IN), .A2(n6534), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(n6573), .ZN(n6527) );
  OAI21_X1 U7507 ( .B1(n6528), .B2(n6536), .A(n6527), .ZN(U3210) );
  AOI22_X1 U7508 ( .A1(REIP_REG_28__SCAN_IN), .A2(n6531), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(n6573), .ZN(n6529) );
  OAI21_X1 U7509 ( .B1(n6530), .B2(n6533), .A(n6529), .ZN(U3211) );
  AOI22_X1 U7510 ( .A1(REIP_REG_29__SCAN_IN), .A2(n6531), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n6573), .ZN(n6532) );
  OAI21_X1 U7511 ( .B1(n6537), .B2(n6533), .A(n6532), .ZN(U3212) );
  AOI22_X1 U7512 ( .A1(REIP_REG_31__SCAN_IN), .A2(n6534), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n6573), .ZN(n6535) );
  OAI21_X1 U7513 ( .B1(n6537), .B2(n6536), .A(n6535), .ZN(U3213) );
  MUX2_X1 U7514 ( .A(BE_N_REG_3__SCAN_IN), .B(BYTEENABLE_REG_3__SCAN_IN), .S(
        n6575), .Z(U3445) );
  MUX2_X1 U7515 ( .A(BE_N_REG_2__SCAN_IN), .B(BYTEENABLE_REG_2__SCAN_IN), .S(
        n6575), .Z(U3446) );
  INV_X1 U7516 ( .A(BE_N_REG_1__SCAN_IN), .ZN(n6799) );
  AOI22_X1 U7517 ( .A1(n6575), .A2(n6538), .B1(n6799), .B2(n6573), .ZN(U3447)
         );
  INV_X1 U7518 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6561) );
  INV_X1 U7519 ( .A(BE_N_REG_0__SCAN_IN), .ZN(n6779) );
  AOI22_X1 U7520 ( .A1(n6575), .A2(n6561), .B1(n6779), .B2(n6573), .ZN(U3448)
         );
  INV_X1 U7521 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6541) );
  INV_X1 U7522 ( .A(n6542), .ZN(n6539) );
  AOI21_X1 U7523 ( .B1(n6541), .B2(n6540), .A(n6539), .ZN(U3451) );
  OAI21_X1 U7524 ( .B1(n6544), .B2(n6543), .A(n6542), .ZN(U3452) );
  OAI221_X1 U7525 ( .B1(n6547), .B2(STATE2_REG_0__SCAN_IN), .C1(n6547), .C2(
        n6546), .A(n6545), .ZN(U3453) );
  AOI22_X1 U7526 ( .A1(n6551), .A2(n6550), .B1(n6549), .B2(n6548), .ZN(n6552)
         );
  INV_X1 U7527 ( .A(n6552), .ZN(n6554) );
  MUX2_X1 U7528 ( .A(n6554), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n6553), 
        .Z(U3456) );
  AOI21_X1 U7529 ( .B1(REIP_REG_0__SCAN_IN), .B2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6556) );
  AOI22_X1 U7530 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .B1(
        n6556), .B2(n6555), .ZN(n6559) );
  INV_X1 U7531 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6558) );
  AOI22_X1 U7532 ( .A1(n6562), .A2(n6559), .B1(n6558), .B2(n6557), .ZN(U3468)
         );
  OAI21_X1 U7533 ( .B1(REIP_REG_1__SCAN_IN), .B2(REIP_REG_0__SCAN_IN), .A(
        n6562), .ZN(n6560) );
  OAI21_X1 U7534 ( .B1(n6562), .B2(n6561), .A(n6560), .ZN(U3469) );
  INV_X1 U7535 ( .A(W_R_N_REG_SCAN_IN), .ZN(n6710) );
  AOI22_X1 U7536 ( .A1(n6575), .A2(READREQUEST_REG_SCAN_IN), .B1(n6710), .B2(
        n6573), .ZN(U3470) );
  AOI211_X1 U7537 ( .C1(n6565), .C2(n6564), .A(n5155), .B(n6563), .ZN(n6568)
         );
  OAI21_X1 U7538 ( .B1(n6568), .B2(n6567), .A(n6566), .ZN(n6572) );
  AOI211_X1 U7539 ( .C1(n6040), .C2(n4324), .A(n6570), .B(n6569), .ZN(n6571)
         );
  MUX2_X1 U7540 ( .A(n6572), .B(REQUESTPENDING_REG_SCAN_IN), .S(n6571), .Z(
        U3472) );
  INV_X1 U7541 ( .A(M_IO_N_REG_SCAN_IN), .ZN(n6885) );
  AOI22_X1 U7542 ( .A1(n6575), .A2(n6574), .B1(n6885), .B2(n6573), .ZN(U3473)
         );
  OAI22_X1 U7543 ( .A1(STATE2_REG_1__SCAN_IN), .A2(keyinput42), .B1(keyinput89), .B2(W_R_N_REG_SCAN_IN), .ZN(n6576) );
  AOI221_X1 U7544 ( .B1(STATE2_REG_1__SCAN_IN), .B2(keyinput42), .C1(
        W_R_N_REG_SCAN_IN), .C2(keyinput89), .A(n6576), .ZN(n6583) );
  OAI22_X1 U7545 ( .A1(ADDRESS_REG_23__SCAN_IN), .A2(keyinput29), .B1(
        DATAO_REG_22__SCAN_IN), .B2(keyinput91), .ZN(n6577) );
  AOI221_X1 U7546 ( .B1(ADDRESS_REG_23__SCAN_IN), .B2(keyinput29), .C1(
        keyinput91), .C2(DATAO_REG_22__SCAN_IN), .A(n6577), .ZN(n6582) );
  OAI22_X1 U7547 ( .A1(INSTQUEUE_REG_12__5__SCAN_IN), .A2(keyinput92), .B1(
        keyinput10), .B2(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n6578) );
  AOI221_X1 U7548 ( .B1(INSTQUEUE_REG_12__5__SCAN_IN), .B2(keyinput92), .C1(
        PHYADDRPOINTER_REG_2__SCAN_IN), .C2(keyinput10), .A(n6578), .ZN(n6581)
         );
  OAI22_X1 U7549 ( .A1(INSTQUEUE_REG_10__6__SCAN_IN), .A2(keyinput108), .B1(
        DATAWIDTH_REG_23__SCAN_IN), .B2(keyinput117), .ZN(n6579) );
  AOI221_X1 U7550 ( .B1(INSTQUEUE_REG_10__6__SCAN_IN), .B2(keyinput108), .C1(
        keyinput117), .C2(DATAWIDTH_REG_23__SCAN_IN), .A(n6579), .ZN(n6580) );
  NAND4_X1 U7551 ( .A1(n6583), .A2(n6582), .A3(n6581), .A4(n6580), .ZN(n6611)
         );
  OAI22_X1 U7552 ( .A1(INSTQUEUE_REG_12__7__SCAN_IN), .A2(keyinput109), .B1(
        keyinput82), .B2(REIP_REG_28__SCAN_IN), .ZN(n6584) );
  AOI221_X1 U7553 ( .B1(INSTQUEUE_REG_12__7__SCAN_IN), .B2(keyinput109), .C1(
        REIP_REG_28__SCAN_IN), .C2(keyinput82), .A(n6584), .ZN(n6591) );
  OAI22_X1 U7554 ( .A1(INSTQUEUE_REG_2__5__SCAN_IN), .A2(keyinput53), .B1(
        MEMORYFETCH_REG_SCAN_IN), .B2(keyinput115), .ZN(n6585) );
  AOI221_X1 U7555 ( .B1(INSTQUEUE_REG_2__5__SCAN_IN), .B2(keyinput53), .C1(
        keyinput115), .C2(MEMORYFETCH_REG_SCAN_IN), .A(n6585), .ZN(n6590) );
  OAI22_X1 U7556 ( .A1(INSTQUEUE_REG_5__7__SCAN_IN), .A2(keyinput56), .B1(
        DATAO_REG_31__SCAN_IN), .B2(keyinput65), .ZN(n6586) );
  AOI221_X1 U7557 ( .B1(INSTQUEUE_REG_5__7__SCAN_IN), .B2(keyinput56), .C1(
        keyinput65), .C2(DATAO_REG_31__SCAN_IN), .A(n6586), .ZN(n6589) );
  OAI22_X1 U7558 ( .A1(INSTQUEUE_REG_1__2__SCAN_IN), .A2(keyinput97), .B1(
        keyinput14), .B2(DATAO_REG_3__SCAN_IN), .ZN(n6587) );
  AOI221_X1 U7559 ( .B1(INSTQUEUE_REG_1__2__SCAN_IN), .B2(keyinput97), .C1(
        DATAO_REG_3__SCAN_IN), .C2(keyinput14), .A(n6587), .ZN(n6588) );
  NAND4_X1 U7560 ( .A1(n6591), .A2(n6590), .A3(n6589), .A4(n6588), .ZN(n6610)
         );
  OAI22_X1 U7561 ( .A1(INSTQUEUE_REG_2__3__SCAN_IN), .A2(keyinput72), .B1(
        keyinput24), .B2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n6592) );
  AOI221_X1 U7562 ( .B1(INSTQUEUE_REG_2__3__SCAN_IN), .B2(keyinput72), .C1(
        INSTADDRPOINTER_REG_6__SCAN_IN), .C2(keyinput24), .A(n6592), .ZN(n6599) );
  OAI22_X1 U7563 ( .A1(EBX_REG_4__SCAN_IN), .A2(keyinput47), .B1(keyinput16), 
        .B2(UWORD_REG_2__SCAN_IN), .ZN(n6593) );
  AOI221_X1 U7564 ( .B1(EBX_REG_4__SCAN_IN), .B2(keyinput47), .C1(
        UWORD_REG_2__SCAN_IN), .C2(keyinput16), .A(n6593), .ZN(n6598) );
  OAI22_X1 U7565 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(keyinput60), .B1(
        keyinput64), .B2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n6594) );
  AOI221_X1 U7566 ( .B1(INSTQUEUE_REG_13__0__SCAN_IN), .B2(keyinput60), .C1(
        PHYADDRPOINTER_REG_14__SCAN_IN), .C2(keyinput64), .A(n6594), .ZN(n6597) );
  OAI22_X1 U7567 ( .A1(READY_N), .A2(keyinput102), .B1(ADDRESS_REG_19__SCAN_IN), .B2(keyinput99), .ZN(n6595) );
  AOI221_X1 U7568 ( .B1(READY_N), .B2(keyinput102), .C1(keyinput99), .C2(
        ADDRESS_REG_19__SCAN_IN), .A(n6595), .ZN(n6596) );
  NAND4_X1 U7569 ( .A1(n6599), .A2(n6598), .A3(n6597), .A4(n6596), .ZN(n6609)
         );
  OAI22_X1 U7570 ( .A1(EBX_REG_1__SCAN_IN), .A2(keyinput84), .B1(
        EBX_REG_7__SCAN_IN), .B2(keyinput116), .ZN(n6600) );
  AOI221_X1 U7571 ( .B1(EBX_REG_1__SCAN_IN), .B2(keyinput84), .C1(keyinput116), 
        .C2(EBX_REG_7__SCAN_IN), .A(n6600), .ZN(n6607) );
  OAI22_X1 U7572 ( .A1(INSTQUEUE_REG_3__6__SCAN_IN), .A2(keyinput35), .B1(
        REIP_REG_18__SCAN_IN), .B2(keyinput77), .ZN(n6601) );
  AOI221_X1 U7573 ( .B1(INSTQUEUE_REG_3__6__SCAN_IN), .B2(keyinput35), .C1(
        keyinput77), .C2(REIP_REG_18__SCAN_IN), .A(n6601), .ZN(n6606) );
  OAI22_X1 U7574 ( .A1(INSTQUEUE_REG_10__7__SCAN_IN), .A2(keyinput112), .B1(
        INSTQUEUE_REG_5__3__SCAN_IN), .B2(keyinput107), .ZN(n6602) );
  AOI221_X1 U7575 ( .B1(INSTQUEUE_REG_10__7__SCAN_IN), .B2(keyinput112), .C1(
        keyinput107), .C2(INSTQUEUE_REG_5__3__SCAN_IN), .A(n6602), .ZN(n6605)
         );
  OAI22_X1 U7576 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(keyinput105), .B1(
        keyinput40), .B2(BE_N_REG_0__SCAN_IN), .ZN(n6603) );
  AOI221_X1 U7577 ( .B1(INSTQUEUE_REG_11__2__SCAN_IN), .B2(keyinput105), .C1(
        BE_N_REG_0__SCAN_IN), .C2(keyinput40), .A(n6603), .ZN(n6604) );
  NAND4_X1 U7578 ( .A1(n6607), .A2(n6606), .A3(n6605), .A4(n6604), .ZN(n6608)
         );
  NOR4_X1 U7579 ( .A1(n6611), .A2(n6610), .A3(n6609), .A4(n6608), .ZN(n6966)
         );
  AOI22_X1 U7580 ( .A1(BYTEENABLE_REG_1__SCAN_IN), .A2(keyinput183), .B1(
        EBX_REG_4__SCAN_IN), .B2(keyinput175), .ZN(n6612) );
  OAI221_X1 U7581 ( .B1(BYTEENABLE_REG_1__SCAN_IN), .B2(keyinput183), .C1(
        EBX_REG_4__SCAN_IN), .C2(keyinput175), .A(n6612), .ZN(n6619) );
  AOI22_X1 U7582 ( .A1(UWORD_REG_4__SCAN_IN), .A2(keyinput161), .B1(
        PHYADDRPOINTER_REG_14__SCAN_IN), .B2(keyinput192), .ZN(n6613) );
  OAI221_X1 U7583 ( .B1(UWORD_REG_4__SCAN_IN), .B2(keyinput161), .C1(
        PHYADDRPOINTER_REG_14__SCAN_IN), .C2(keyinput192), .A(n6613), .ZN(
        n6618) );
  AOI22_X1 U7584 ( .A1(ADDRESS_REG_23__SCAN_IN), .A2(keyinput157), .B1(
        EAX_REG_18__SCAN_IN), .B2(keyinput222), .ZN(n6614) );
  OAI221_X1 U7585 ( .B1(ADDRESS_REG_23__SCAN_IN), .B2(keyinput157), .C1(
        EAX_REG_18__SCAN_IN), .C2(keyinput222), .A(n6614), .ZN(n6617) );
  AOI22_X1 U7586 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(keyinput228), .B1(
        REIP_REG_3__SCAN_IN), .B2(keyinput139), .ZN(n6615) );
  OAI221_X1 U7587 ( .B1(DATAWIDTH_REG_15__SCAN_IN), .B2(keyinput228), .C1(
        REIP_REG_3__SCAN_IN), .C2(keyinput139), .A(n6615), .ZN(n6616) );
  NOR4_X1 U7588 ( .A1(n6619), .A2(n6618), .A3(n6617), .A4(n6616), .ZN(n6647)
         );
  AOI22_X1 U7589 ( .A1(ADDRESS_REG_25__SCAN_IN), .A2(keyinput202), .B1(
        DATAWIDTH_REG_13__SCAN_IN), .B2(keyinput211), .ZN(n6620) );
  OAI221_X1 U7590 ( .B1(ADDRESS_REG_25__SCAN_IN), .B2(keyinput202), .C1(
        DATAWIDTH_REG_13__SCAN_IN), .C2(keyinput211), .A(n6620), .ZN(n6627) );
  AOI22_X1 U7591 ( .A1(REIP_REG_9__SCAN_IN), .A2(keyinput155), .B1(READY_N), 
        .B2(keyinput230), .ZN(n6621) );
  OAI221_X1 U7592 ( .B1(REIP_REG_9__SCAN_IN), .B2(keyinput155), .C1(READY_N), 
        .C2(keyinput230), .A(n6621), .ZN(n6626) );
  AOI22_X1 U7593 ( .A1(REIP_REG_15__SCAN_IN), .A2(keyinput194), .B1(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(keyinput224), .ZN(n6622) );
  OAI221_X1 U7594 ( .B1(REIP_REG_15__SCAN_IN), .B2(keyinput194), .C1(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C2(keyinput224), .A(n6622), .ZN(
        n6625) );
  AOI22_X1 U7595 ( .A1(DATAI_1_), .A2(keyinput231), .B1(REIP_REG_18__SCAN_IN), 
        .B2(keyinput205), .ZN(n6623) );
  OAI221_X1 U7596 ( .B1(DATAI_1_), .B2(keyinput231), .C1(REIP_REG_18__SCAN_IN), 
        .C2(keyinput205), .A(n6623), .ZN(n6624) );
  NOR4_X1 U7597 ( .A1(n6627), .A2(n6626), .A3(n6625), .A4(n6624), .ZN(n6646)
         );
  AOI22_X1 U7598 ( .A1(PHYADDRPOINTER_REG_15__SCAN_IN), .A2(keyinput182), .B1(
        INSTQUEUE_REG_4__0__SCAN_IN), .B2(keyinput216), .ZN(n6628) );
  OAI221_X1 U7599 ( .B1(PHYADDRPOINTER_REG_15__SCAN_IN), .B2(keyinput182), 
        .C1(INSTQUEUE_REG_4__0__SCAN_IN), .C2(keyinput216), .A(n6628), .ZN(
        n6635) );
  AOI22_X1 U7600 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(keyinput186), .B1(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(keyinput166), .ZN(n6629) );
  OAI221_X1 U7601 ( .B1(INSTQUEUE_REG_9__6__SCAN_IN), .B2(keyinput186), .C1(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C2(keyinput166), .A(n6629), .ZN(
        n6634) );
  AOI22_X1 U7602 ( .A1(DATAI_29_), .A2(keyinput159), .B1(EAX_REG_24__SCAN_IN), 
        .B2(keyinput201), .ZN(n6630) );
  OAI221_X1 U7603 ( .B1(DATAI_29_), .B2(keyinput159), .C1(EAX_REG_24__SCAN_IN), 
        .C2(keyinput201), .A(n6630), .ZN(n6633) );
  AOI22_X1 U7604 ( .A1(EAX_REG_20__SCAN_IN), .A2(keyinput173), .B1(
        EAX_REG_3__SCAN_IN), .B2(keyinput215), .ZN(n6631) );
  OAI221_X1 U7605 ( .B1(EAX_REG_20__SCAN_IN), .B2(keyinput173), .C1(
        EAX_REG_3__SCAN_IN), .C2(keyinput215), .A(n6631), .ZN(n6632) );
  NOR4_X1 U7606 ( .A1(n6635), .A2(n6634), .A3(n6633), .A4(n6632), .ZN(n6645)
         );
  AOI22_X1 U7607 ( .A1(UWORD_REG_5__SCAN_IN), .A2(keyinput187), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(keyinput140), .ZN(n6636) );
  OAI221_X1 U7608 ( .B1(UWORD_REG_5__SCAN_IN), .B2(keyinput187), .C1(
        ADDRESS_REG_7__SCAN_IN), .C2(keyinput140), .A(n6636), .ZN(n6643) );
  AOI22_X1 U7609 ( .A1(DATAO_REG_10__SCAN_IN), .A2(keyinput226), .B1(
        INSTQUEUE_REG_3__4__SCAN_IN), .B2(keyinput179), .ZN(n6637) );
  OAI221_X1 U7610 ( .B1(DATAO_REG_10__SCAN_IN), .B2(keyinput226), .C1(
        INSTQUEUE_REG_3__4__SCAN_IN), .C2(keyinput179), .A(n6637), .ZN(n6642)
         );
  AOI22_X1 U7611 ( .A1(M_IO_N_REG_SCAN_IN), .A2(keyinput145), .B1(
        PHYADDRPOINTER_REG_4__SCAN_IN), .B2(keyinput198), .ZN(n6638) );
  OAI221_X1 U7612 ( .B1(M_IO_N_REG_SCAN_IN), .B2(keyinput145), .C1(
        PHYADDRPOINTER_REG_4__SCAN_IN), .C2(keyinput198), .A(n6638), .ZN(n6641) );
  AOI22_X1 U7613 ( .A1(BE_N_REG_1__SCAN_IN), .A2(keyinput254), .B1(
        DATAO_REG_3__SCAN_IN), .B2(keyinput142), .ZN(n6639) );
  OAI221_X1 U7614 ( .B1(BE_N_REG_1__SCAN_IN), .B2(keyinput254), .C1(
        DATAO_REG_3__SCAN_IN), .C2(keyinput142), .A(n6639), .ZN(n6640) );
  NOR4_X1 U7615 ( .A1(n6643), .A2(n6642), .A3(n6641), .A4(n6640), .ZN(n6644)
         );
  NAND4_X1 U7616 ( .A1(n6647), .A2(n6646), .A3(n6645), .A4(n6644), .ZN(n6794)
         );
  AOI22_X1 U7617 ( .A1(PHYADDRPOINTER_REG_29__SCAN_IN), .A2(keyinput130), .B1(
        EBX_REG_14__SCAN_IN), .B2(keyinput133), .ZN(n6648) );
  OAI221_X1 U7618 ( .B1(PHYADDRPOINTER_REG_29__SCAN_IN), .B2(keyinput130), 
        .C1(EBX_REG_14__SCAN_IN), .C2(keyinput133), .A(n6648), .ZN(n6655) );
  AOI22_X1 U7619 ( .A1(PHYADDRPOINTER_REG_25__SCAN_IN), .A2(keyinput147), .B1(
        INSTQUEUE_REG_0__7__SCAN_IN), .B2(keyinput174), .ZN(n6649) );
  OAI221_X1 U7620 ( .B1(PHYADDRPOINTER_REG_25__SCAN_IN), .B2(keyinput147), 
        .C1(INSTQUEUE_REG_0__7__SCAN_IN), .C2(keyinput174), .A(n6649), .ZN(
        n6654) );
  AOI22_X1 U7621 ( .A1(ADDRESS_REG_8__SCAN_IN), .A2(keyinput213), .B1(
        MEMORYFETCH_REG_SCAN_IN), .B2(keyinput243), .ZN(n6650) );
  OAI221_X1 U7622 ( .B1(ADDRESS_REG_8__SCAN_IN), .B2(keyinput213), .C1(
        MEMORYFETCH_REG_SCAN_IN), .C2(keyinput243), .A(n6650), .ZN(n6653) );
  AOI22_X1 U7623 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(keyinput188), .B1(
        INSTQUEUE_REG_12__7__SCAN_IN), .B2(keyinput237), .ZN(n6651) );
  OAI221_X1 U7624 ( .B1(INSTQUEUE_REG_13__0__SCAN_IN), .B2(keyinput188), .C1(
        INSTQUEUE_REG_12__7__SCAN_IN), .C2(keyinput237), .A(n6651), .ZN(n6652)
         );
  NOR4_X1 U7625 ( .A1(n6655), .A2(n6654), .A3(n6653), .A4(n6652), .ZN(n6683)
         );
  AOI22_X1 U7626 ( .A1(DATAO_REG_19__SCAN_IN), .A2(keyinput223), .B1(
        EAX_REG_25__SCAN_IN), .B2(keyinput238), .ZN(n6656) );
  OAI221_X1 U7627 ( .B1(DATAO_REG_19__SCAN_IN), .B2(keyinput223), .C1(
        EAX_REG_25__SCAN_IN), .C2(keyinput238), .A(n6656), .ZN(n6663) );
  AOI22_X1 U7628 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(keyinput209), .B1(
        PHYADDRPOINTER_REG_2__SCAN_IN), .B2(keyinput138), .ZN(n6657) );
  OAI221_X1 U7629 ( .B1(DATAWIDTH_REG_19__SCAN_IN), .B2(keyinput209), .C1(
        PHYADDRPOINTER_REG_2__SCAN_IN), .C2(keyinput138), .A(n6657), .ZN(n6662) );
  AOI22_X1 U7630 ( .A1(BYTEENABLE_REG_3__SCAN_IN), .A2(keyinput199), .B1(
        DATAWIDTH_REG_18__SCAN_IN), .B2(keyinput164), .ZN(n6658) );
  OAI221_X1 U7631 ( .B1(BYTEENABLE_REG_3__SCAN_IN), .B2(keyinput199), .C1(
        DATAWIDTH_REG_18__SCAN_IN), .C2(keyinput164), .A(n6658), .ZN(n6661) );
  AOI22_X1 U7632 ( .A1(LWORD_REG_6__SCAN_IN), .A2(keyinput252), .B1(
        DATAO_REG_31__SCAN_IN), .B2(keyinput193), .ZN(n6659) );
  OAI221_X1 U7633 ( .B1(LWORD_REG_6__SCAN_IN), .B2(keyinput252), .C1(
        DATAO_REG_31__SCAN_IN), .C2(keyinput193), .A(n6659), .ZN(n6660) );
  NOR4_X1 U7634 ( .A1(n6663), .A2(n6662), .A3(n6661), .A4(n6660), .ZN(n6682)
         );
  AOI22_X1 U7635 ( .A1(DATAI_14_), .A2(keyinput148), .B1(REIP_REG_1__SCAN_IN), 
        .B2(keyinput134), .ZN(n6664) );
  OAI221_X1 U7636 ( .B1(DATAI_14_), .B2(keyinput148), .C1(REIP_REG_1__SCAN_IN), 
        .C2(keyinput134), .A(n6664), .ZN(n6671) );
  AOI22_X1 U7637 ( .A1(ADDRESS_REG_19__SCAN_IN), .A2(keyinput227), .B1(
        REIP_REG_31__SCAN_IN), .B2(keyinput162), .ZN(n6665) );
  OAI221_X1 U7638 ( .B1(ADDRESS_REG_19__SCAN_IN), .B2(keyinput227), .C1(
        REIP_REG_31__SCAN_IN), .C2(keyinput162), .A(n6665), .ZN(n6670) );
  AOI22_X1 U7639 ( .A1(REIP_REG_28__SCAN_IN), .A2(keyinput210), .B1(
        INSTQUEUE_REG_2__4__SCAN_IN), .B2(keyinput180), .ZN(n6666) );
  OAI221_X1 U7640 ( .B1(REIP_REG_28__SCAN_IN), .B2(keyinput210), .C1(
        INSTQUEUE_REG_2__4__SCAN_IN), .C2(keyinput180), .A(n6666), .ZN(n6669)
         );
  AOI22_X1 U7641 ( .A1(ADS_N_REG_SCAN_IN), .A2(keyinput165), .B1(
        INSTQUEUE_REG_15__1__SCAN_IN), .B2(keyinput190), .ZN(n6667) );
  OAI221_X1 U7642 ( .B1(ADS_N_REG_SCAN_IN), .B2(keyinput165), .C1(
        INSTQUEUE_REG_15__1__SCAN_IN), .C2(keyinput190), .A(n6667), .ZN(n6668)
         );
  NOR4_X1 U7643 ( .A1(n6671), .A2(n6670), .A3(n6669), .A4(n6668), .ZN(n6681)
         );
  AOI22_X1 U7644 ( .A1(ADDRESS_REG_21__SCAN_IN), .A2(keyinput153), .B1(
        INSTQUEUE_REG_15__2__SCAN_IN), .B2(keyinput131), .ZN(n6672) );
  OAI221_X1 U7645 ( .B1(ADDRESS_REG_21__SCAN_IN), .B2(keyinput153), .C1(
        INSTQUEUE_REG_15__2__SCAN_IN), .C2(keyinput131), .A(n6672), .ZN(n6679)
         );
  AOI22_X1 U7646 ( .A1(LWORD_REG_1__SCAN_IN), .A2(keyinput203), .B1(
        INSTADDRPOINTER_REG_3__SCAN_IN), .B2(keyinput239), .ZN(n6673) );
  OAI221_X1 U7647 ( .B1(LWORD_REG_1__SCAN_IN), .B2(keyinput203), .C1(
        INSTADDRPOINTER_REG_3__SCAN_IN), .C2(keyinput239), .A(n6673), .ZN(
        n6678) );
  AOI22_X1 U7648 ( .A1(DATAI_13_), .A2(keyinput177), .B1(EAX_REG_27__SCAN_IN), 
        .B2(keyinput136), .ZN(n6674) );
  OAI221_X1 U7649 ( .B1(DATAI_13_), .B2(keyinput177), .C1(EAX_REG_27__SCAN_IN), 
        .C2(keyinput136), .A(n6674), .ZN(n6677) );
  AOI22_X1 U7650 ( .A1(PHYADDRPOINTER_REG_17__SCAN_IN), .A2(keyinput178), .B1(
        EBX_REG_1__SCAN_IN), .B2(keyinput212), .ZN(n6675) );
  OAI221_X1 U7651 ( .B1(PHYADDRPOINTER_REG_17__SCAN_IN), .B2(keyinput178), 
        .C1(EBX_REG_1__SCAN_IN), .C2(keyinput212), .A(n6675), .ZN(n6676) );
  NOR4_X1 U7652 ( .A1(n6679), .A2(n6678), .A3(n6677), .A4(n6676), .ZN(n6680)
         );
  NAND4_X1 U7653 ( .A1(n6683), .A2(n6682), .A3(n6681), .A4(n6680), .ZN(n6793)
         );
  AOI22_X1 U7654 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(keyinput129), .B1(
        INSTQUEUE_REG_14__2__SCAN_IN), .B2(keyinput247), .ZN(n6684) );
  OAI221_X1 U7655 ( .B1(DATAWIDTH_REG_4__SCAN_IN), .B2(keyinput129), .C1(
        INSTQUEUE_REG_14__2__SCAN_IN), .C2(keyinput247), .A(n6684), .ZN(n6693)
         );
  AOI22_X1 U7656 ( .A1(PHYADDRPOINTER_REG_31__SCAN_IN), .A2(keyinput253), .B1(
        EBX_REG_13__SCAN_IN), .B2(keyinput171), .ZN(n6685) );
  OAI221_X1 U7657 ( .B1(PHYADDRPOINTER_REG_31__SCAN_IN), .B2(keyinput253), 
        .C1(EBX_REG_13__SCAN_IN), .C2(keyinput171), .A(n6685), .ZN(n6692) );
  INV_X1 U7658 ( .A(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n6894) );
  INV_X1 U7659 ( .A(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n6687) );
  AOI22_X1 U7660 ( .A1(n6894), .A2(keyinput135), .B1(n6687), .B2(keyinput181), 
        .ZN(n6686) );
  OAI221_X1 U7661 ( .B1(n6894), .B2(keyinput135), .C1(n6687), .C2(keyinput181), 
        .A(n6686), .ZN(n6691) );
  INV_X1 U7662 ( .A(EBX_REG_17__SCAN_IN), .ZN(n6844) );
  INV_X1 U7663 ( .A(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n6689) );
  AOI22_X1 U7664 ( .A1(n6844), .A2(keyinput137), .B1(n6689), .B2(keyinput149), 
        .ZN(n6688) );
  OAI221_X1 U7665 ( .B1(n6844), .B2(keyinput137), .C1(n6689), .C2(keyinput149), 
        .A(n6688), .ZN(n6690) );
  NOR4_X1 U7666 ( .A1(n6693), .A2(n6692), .A3(n6691), .A4(n6690), .ZN(n6733)
         );
  AOI22_X1 U7667 ( .A1(n6909), .A2(keyinput197), .B1(keyinput206), .B2(n6695), 
        .ZN(n6694) );
  OAI221_X1 U7668 ( .B1(n6909), .B2(keyinput197), .C1(n6695), .C2(keyinput206), 
        .A(n6694), .ZN(n6703) );
  AOI22_X1 U7669 ( .A1(n6900), .A2(keyinput156), .B1(n4924), .B2(keyinput248), 
        .ZN(n6696) );
  OAI221_X1 U7670 ( .B1(n6900), .B2(keyinput156), .C1(n4924), .C2(keyinput248), 
        .A(n6696), .ZN(n6702) );
  INV_X1 U7671 ( .A(UWORD_REG_0__SCAN_IN), .ZN(n6698) );
  AOI22_X1 U7672 ( .A1(n6861), .A2(keyinput196), .B1(keyinput249), .B2(n6698), 
        .ZN(n6697) );
  OAI221_X1 U7673 ( .B1(n6861), .B2(keyinput196), .C1(n6698), .C2(keyinput249), 
        .A(n6697), .ZN(n6701) );
  AOI22_X1 U7674 ( .A1(n3629), .A2(keyinput234), .B1(n6798), .B2(keyinput207), 
        .ZN(n6699) );
  OAI221_X1 U7675 ( .B1(n3629), .B2(keyinput234), .C1(n6798), .C2(keyinput207), 
        .A(n6699), .ZN(n6700) );
  NOR4_X1 U7676 ( .A1(n6703), .A2(n6702), .A3(n6701), .A4(n6700), .ZN(n6732)
         );
  INV_X1 U7677 ( .A(LWORD_REG_0__SCAN_IN), .ZN(n6705) );
  AOI22_X1 U7678 ( .A1(n6826), .A2(keyinput132), .B1(keyinput172), .B2(n6705), 
        .ZN(n6704) );
  OAI221_X1 U7679 ( .B1(n6826), .B2(keyinput132), .C1(n6705), .C2(keyinput172), 
        .A(n6704), .ZN(n6716) );
  INV_X1 U7680 ( .A(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n6860) );
  AOI22_X1 U7681 ( .A1(n6707), .A2(keyinput221), .B1(n6860), .B2(keyinput151), 
        .ZN(n6706) );
  OAI221_X1 U7682 ( .B1(n6707), .B2(keyinput221), .C1(n6860), .C2(keyinput151), 
        .A(n6706), .ZN(n6715) );
  AOI22_X1 U7683 ( .A1(n6710), .A2(keyinput217), .B1(keyinput250), .B2(n6709), 
        .ZN(n6708) );
  OAI221_X1 U7684 ( .B1(n6710), .B2(keyinput217), .C1(n6709), .C2(keyinput250), 
        .A(n6708), .ZN(n6714) );
  INV_X1 U7685 ( .A(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n6712) );
  AOI22_X1 U7686 ( .A1(n6712), .A2(keyinput141), .B1(keyinput185), .B2(n6814), 
        .ZN(n6711) );
  OAI221_X1 U7687 ( .B1(n6712), .B2(keyinput141), .C1(n6814), .C2(keyinput185), 
        .A(n6711), .ZN(n6713) );
  NOR4_X1 U7688 ( .A1(n6716), .A2(n6715), .A3(n6714), .A4(n6713), .ZN(n6731)
         );
  INV_X1 U7689 ( .A(UWORD_REG_2__SCAN_IN), .ZN(n6718) );
  AOI22_X1 U7690 ( .A1(n6719), .A2(keyinput191), .B1(keyinput144), .B2(n6718), 
        .ZN(n6717) );
  OAI221_X1 U7691 ( .B1(n6719), .B2(keyinput191), .C1(n6718), .C2(keyinput144), 
        .A(n6717), .ZN(n6729) );
  AOI22_X1 U7692 ( .A1(n6721), .A2(keyinput241), .B1(n5491), .B2(keyinput154), 
        .ZN(n6720) );
  OAI221_X1 U7693 ( .B1(n6721), .B2(keyinput241), .C1(n5491), .C2(keyinput154), 
        .A(n6720), .ZN(n6728) );
  AOI22_X1 U7694 ( .A1(n6724), .A2(keyinput235), .B1(n6723), .B2(keyinput229), 
        .ZN(n6722) );
  OAI221_X1 U7695 ( .B1(n6724), .B2(keyinput235), .C1(n6723), .C2(keyinput229), 
        .A(n6722), .ZN(n6727) );
  INV_X1 U7696 ( .A(DATAI_24_), .ZN(n6843) );
  INV_X1 U7697 ( .A(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n6906) );
  AOI22_X1 U7698 ( .A1(n6843), .A2(keyinput208), .B1(n6906), .B2(keyinput143), 
        .ZN(n6725) );
  OAI221_X1 U7699 ( .B1(n6843), .B2(keyinput208), .C1(n6906), .C2(keyinput143), 
        .A(n6725), .ZN(n6726) );
  NOR4_X1 U7700 ( .A1(n6729), .A2(n6728), .A3(n6727), .A4(n6726), .ZN(n6730)
         );
  NAND4_X1 U7701 ( .A1(n6733), .A2(n6732), .A3(n6731), .A4(n6730), .ZN(n6792)
         );
  INV_X1 U7702 ( .A(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n6735) );
  AOI22_X1 U7703 ( .A1(n6736), .A2(keyinput170), .B1(keyinput200), .B2(n6735), 
        .ZN(n6734) );
  OAI221_X1 U7704 ( .B1(n6736), .B2(keyinput170), .C1(n6735), .C2(keyinput200), 
        .A(n6734), .ZN(n6747) );
  INV_X1 U7705 ( .A(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n6818) );
  AOI22_X1 U7706 ( .A1(n6818), .A2(keyinput146), .B1(keyinput219), .B2(n6738), 
        .ZN(n6737) );
  OAI221_X1 U7707 ( .B1(n6818), .B2(keyinput146), .C1(n6738), .C2(keyinput219), 
        .A(n6737), .ZN(n6746) );
  AOI22_X1 U7708 ( .A1(n6877), .A2(keyinput128), .B1(keyinput245), .B2(n6740), 
        .ZN(n6739) );
  OAI221_X1 U7709 ( .B1(n6877), .B2(keyinput128), .C1(n6740), .C2(keyinput245), 
        .A(n6739), .ZN(n6745) );
  INV_X1 U7710 ( .A(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n6742) );
  AOI22_X1 U7711 ( .A1(n6743), .A2(keyinput244), .B1(n6742), .B2(keyinput233), 
        .ZN(n6741) );
  OAI221_X1 U7712 ( .B1(n6743), .B2(keyinput244), .C1(n6742), .C2(keyinput233), 
        .A(n6741), .ZN(n6744) );
  NOR4_X1 U7713 ( .A1(n6747), .A2(n6746), .A3(n6745), .A4(n6744), .ZN(n6790)
         );
  AOI22_X1 U7714 ( .A1(n6749), .A2(keyinput255), .B1(n6804), .B2(keyinput214), 
        .ZN(n6748) );
  OAI221_X1 U7715 ( .B1(n6749), .B2(keyinput255), .C1(n6804), .C2(keyinput214), 
        .A(n6748), .ZN(n6760) );
  INV_X1 U7716 ( .A(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n6751) );
  AOI22_X1 U7717 ( .A1(n6752), .A2(keyinput152), .B1(n6751), .B2(keyinput220), 
        .ZN(n6750) );
  OAI221_X1 U7718 ( .B1(n6752), .B2(keyinput152), .C1(n6751), .C2(keyinput220), 
        .A(n6750), .ZN(n6759) );
  INV_X1 U7719 ( .A(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n6834) );
  AOI22_X1 U7720 ( .A1(n6832), .A2(keyinput167), .B1(n6834), .B2(keyinput251), 
        .ZN(n6753) );
  OAI221_X1 U7721 ( .B1(n6832), .B2(keyinput167), .C1(n6834), .C2(keyinput251), 
        .A(n6753), .ZN(n6758) );
  INV_X1 U7722 ( .A(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n6756) );
  INV_X1 U7723 ( .A(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n6755) );
  AOI22_X1 U7724 ( .A1(n6756), .A2(keyinput236), .B1(n6755), .B2(keyinput225), 
        .ZN(n6754) );
  OAI221_X1 U7725 ( .B1(n6756), .B2(keyinput236), .C1(n6755), .C2(keyinput225), 
        .A(n6754), .ZN(n6757) );
  NOR4_X1 U7726 ( .A1(n6760), .A2(n6759), .A3(n6758), .A4(n6757), .ZN(n6789)
         );
  AOI22_X1 U7727 ( .A1(n6910), .A2(keyinput242), .B1(keyinput246), .B2(n6867), 
        .ZN(n6761) );
  OAI221_X1 U7728 ( .B1(n6910), .B2(keyinput242), .C1(n6867), .C2(keyinput246), 
        .A(n6761), .ZN(n6773) );
  AOI22_X1 U7729 ( .A1(n6764), .A2(keyinput218), .B1(n6763), .B2(keyinput184), 
        .ZN(n6762) );
  OAI221_X1 U7730 ( .B1(n6764), .B2(keyinput218), .C1(n6763), .C2(keyinput184), 
        .A(n6762), .ZN(n6772) );
  INV_X1 U7731 ( .A(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n6766) );
  AOI22_X1 U7732 ( .A1(n6767), .A2(keyinput189), .B1(n6766), .B2(keyinput163), 
        .ZN(n6765) );
  OAI221_X1 U7733 ( .B1(n6767), .B2(keyinput189), .C1(n6766), .C2(keyinput163), 
        .A(n6765), .ZN(n6771) );
  AOI22_X1 U7734 ( .A1(n6816), .A2(keyinput150), .B1(keyinput158), .B2(n6769), 
        .ZN(n6768) );
  OAI221_X1 U7735 ( .B1(n6816), .B2(keyinput150), .C1(n6769), .C2(keyinput158), 
        .A(n6768), .ZN(n6770) );
  NOR4_X1 U7736 ( .A1(n6773), .A2(n6772), .A3(n6771), .A4(n6770), .ZN(n6788)
         );
  AOI22_X1 U7737 ( .A1(n6775), .A2(keyinput160), .B1(keyinput169), .B2(n6891), 
        .ZN(n6774) );
  OAI221_X1 U7738 ( .B1(n6775), .B2(keyinput160), .C1(n6891), .C2(keyinput169), 
        .A(n6774), .ZN(n6786) );
  INV_X1 U7739 ( .A(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n6777) );
  AOI22_X1 U7740 ( .A1(n6777), .A2(keyinput240), .B1(keyinput204), .B2(n6863), 
        .ZN(n6776) );
  OAI221_X1 U7741 ( .B1(n6777), .B2(keyinput240), .C1(n6863), .C2(keyinput204), 
        .A(n6776), .ZN(n6785) );
  AOI22_X1 U7742 ( .A1(n6779), .A2(keyinput168), .B1(n6805), .B2(keyinput232), 
        .ZN(n6778) );
  OAI221_X1 U7743 ( .B1(n6779), .B2(keyinput168), .C1(n6805), .C2(keyinput232), 
        .A(n6778), .ZN(n6784) );
  AOI22_X1 U7744 ( .A1(n6782), .A2(keyinput176), .B1(n6781), .B2(keyinput195), 
        .ZN(n6780) );
  OAI221_X1 U7745 ( .B1(n6782), .B2(keyinput176), .C1(n6781), .C2(keyinput195), 
        .A(n6780), .ZN(n6783) );
  NOR4_X1 U7746 ( .A1(n6786), .A2(n6785), .A3(n6784), .A4(n6783), .ZN(n6787)
         );
  NAND4_X1 U7747 ( .A1(n6790), .A2(n6789), .A3(n6788), .A4(n6787), .ZN(n6791)
         );
  NOR4_X1 U7748 ( .A1(n6794), .A2(n6793), .A3(n6792), .A4(n6791), .ZN(n6926)
         );
  AOI22_X1 U7749 ( .A1(n4708), .A2(keyinput62), .B1(keyinput59), .B2(n6796), 
        .ZN(n6795) );
  OAI221_X1 U7750 ( .B1(n4708), .B2(keyinput62), .C1(n6796), .C2(keyinput59), 
        .A(n6795), .ZN(n6809) );
  AOI22_X1 U7751 ( .A1(n6799), .A2(keyinput126), .B1(n6798), .B2(keyinput79), 
        .ZN(n6797) );
  OAI221_X1 U7752 ( .B1(n6799), .B2(keyinput126), .C1(n6798), .C2(keyinput79), 
        .A(n6797), .ZN(n6808) );
  AOI22_X1 U7753 ( .A1(n6802), .A2(keyinput111), .B1(keyinput11), .B2(n6801), 
        .ZN(n6800) );
  OAI221_X1 U7754 ( .B1(n6802), .B2(keyinput111), .C1(n6801), .C2(keyinput11), 
        .A(n6800), .ZN(n6807) );
  AOI22_X1 U7755 ( .A1(n6805), .A2(keyinput104), .B1(n6804), .B2(keyinput86), 
        .ZN(n6803) );
  OAI221_X1 U7756 ( .B1(n6805), .B2(keyinput104), .C1(n6804), .C2(keyinput86), 
        .A(n6803), .ZN(n6806) );
  NOR4_X1 U7757 ( .A1(n6809), .A2(n6808), .A3(n6807), .A4(n6806), .ZN(n6858)
         );
  AOI22_X1 U7758 ( .A1(n6812), .A2(keyinput85), .B1(n6811), .B2(keyinput66), 
        .ZN(n6810) );
  OAI221_X1 U7759 ( .B1(n6812), .B2(keyinput85), .C1(n6811), .C2(keyinput66), 
        .A(n6810), .ZN(n6824) );
  AOI22_X1 U7760 ( .A1(n6814), .A2(keyinput57), .B1(n5744), .B2(keyinput31), 
        .ZN(n6813) );
  OAI221_X1 U7761 ( .B1(n6814), .B2(keyinput57), .C1(n5744), .C2(keyinput31), 
        .A(n6813), .ZN(n6823) );
  AOI22_X1 U7762 ( .A1(n6817), .A2(keyinput36), .B1(n6816), .B2(keyinput22), 
        .ZN(n6815) );
  OAI221_X1 U7763 ( .B1(n6817), .B2(keyinput36), .C1(n6816), .C2(keyinput22), 
        .A(n6815), .ZN(n6822) );
  XOR2_X1 U7764 ( .A(n6818), .B(keyinput18), .Z(n6820) );
  XNOR2_X1 U7765 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(keyinput96), .ZN(
        n6819) );
  NAND2_X1 U7766 ( .A1(n6820), .A2(n6819), .ZN(n6821) );
  NOR4_X1 U7767 ( .A1(n6824), .A2(n6823), .A3(n6822), .A4(n6821), .ZN(n6857)
         );
  INV_X1 U7768 ( .A(LWORD_REG_1__SCAN_IN), .ZN(n6827) );
  AOI22_X1 U7769 ( .A1(n6827), .A2(keyinput75), .B1(keyinput4), .B2(n6826), 
        .ZN(n6825) );
  OAI221_X1 U7770 ( .B1(n6827), .B2(keyinput75), .C1(n6826), .C2(keyinput4), 
        .A(n6825), .ZN(n6838) );
  AOI22_X1 U7771 ( .A1(n3940), .A2(keyinput45), .B1(keyinput34), .B2(n6829), 
        .ZN(n6828) );
  OAI221_X1 U7772 ( .B1(n3940), .B2(keyinput45), .C1(n6829), .C2(keyinput34), 
        .A(n6828), .ZN(n6837) );
  AOI22_X1 U7773 ( .A1(n6832), .A2(keyinput39), .B1(n6831), .B2(keyinput46), 
        .ZN(n6830) );
  OAI221_X1 U7774 ( .B1(n6832), .B2(keyinput39), .C1(n6831), .C2(keyinput46), 
        .A(n6830), .ZN(n6836) );
  AOI22_X1 U7775 ( .A1(n6834), .A2(keyinput123), .B1(keyinput125), .B2(n4182), 
        .ZN(n6833) );
  OAI221_X1 U7776 ( .B1(n6834), .B2(keyinput123), .C1(n4182), .C2(keyinput125), 
        .A(n6833), .ZN(n6835) );
  NOR4_X1 U7777 ( .A1(n6838), .A2(n6837), .A3(n6836), .A4(n6835), .ZN(n6856)
         );
  AOI22_X1 U7778 ( .A1(n6841), .A2(keyinput94), .B1(keyinput124), .B2(n6840), 
        .ZN(n6839) );
  OAI221_X1 U7779 ( .B1(n6841), .B2(keyinput94), .C1(n6840), .C2(keyinput124), 
        .A(n6839), .ZN(n6854) );
  AOI22_X1 U7780 ( .A1(n6844), .A2(keyinput9), .B1(keyinput80), .B2(n6843), 
        .ZN(n6842) );
  OAI221_X1 U7781 ( .B1(n6844), .B2(keyinput9), .C1(n6843), .C2(keyinput80), 
        .A(n6842), .ZN(n6853) );
  AOI22_X1 U7782 ( .A1(n6847), .A2(keyinput71), .B1(n6846), .B2(keyinput12), 
        .ZN(n6845) );
  OAI221_X1 U7783 ( .B1(n6847), .B2(keyinput71), .C1(n6846), .C2(keyinput12), 
        .A(n6845), .ZN(n6852) );
  INV_X1 U7784 ( .A(UWORD_REG_4__SCAN_IN), .ZN(n6849) );
  AOI22_X1 U7785 ( .A1(n6850), .A2(keyinput1), .B1(n6849), .B2(keyinput33), 
        .ZN(n6848) );
  OAI221_X1 U7786 ( .B1(n6850), .B2(keyinput1), .C1(n6849), .C2(keyinput33), 
        .A(n6848), .ZN(n6851) );
  NOR4_X1 U7787 ( .A1(n6854), .A2(n6853), .A3(n6852), .A4(n6851), .ZN(n6855)
         );
  NAND4_X1 U7788 ( .A1(n6858), .A2(n6857), .A3(n6856), .A4(n6855), .ZN(n6925)
         );
  AOI22_X1 U7789 ( .A1(n6861), .A2(keyinput68), .B1(n6860), .B2(keyinput23), 
        .ZN(n6859) );
  OAI221_X1 U7790 ( .B1(n6861), .B2(keyinput68), .C1(n6860), .C2(keyinput23), 
        .A(n6859), .ZN(n6873) );
  AOI22_X1 U7791 ( .A1(n6864), .A2(keyinput49), .B1(n6863), .B2(keyinput76), 
        .ZN(n6862) );
  OAI221_X1 U7792 ( .B1(n6864), .B2(keyinput49), .C1(n6863), .C2(keyinput76), 
        .A(n6862), .ZN(n6872) );
  INV_X1 U7793 ( .A(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n6866) );
  AOI22_X1 U7794 ( .A1(n6867), .A2(keyinput118), .B1(n6866), .B2(keyinput52), 
        .ZN(n6865) );
  OAI221_X1 U7795 ( .B1(n6867), .B2(keyinput118), .C1(n6866), .C2(keyinput52), 
        .A(n6865), .ZN(n6871) );
  XOR2_X1 U7796 ( .A(n3629), .B(keyinput106), .Z(n6869) );
  XNOR2_X1 U7797 ( .A(INSTQUEUE_REG_4__0__SCAN_IN), .B(keyinput88), .ZN(n6868)
         );
  NAND2_X1 U7798 ( .A1(n6869), .A2(n6868), .ZN(n6870) );
  NOR4_X1 U7799 ( .A1(n6873), .A2(n6872), .A3(n6871), .A4(n6870), .ZN(n6923)
         );
  AOI22_X1 U7800 ( .A1(n6875), .A2(keyinput100), .B1(n4097), .B2(keyinput73), 
        .ZN(n6874) );
  OAI221_X1 U7801 ( .B1(n6875), .B2(keyinput100), .C1(n4097), .C2(keyinput73), 
        .A(n6874), .ZN(n6880) );
  XNOR2_X1 U7802 ( .A(n6876), .B(keyinput38), .ZN(n6879) );
  XNOR2_X1 U7803 ( .A(n6877), .B(keyinput0), .ZN(n6878) );
  OR3_X1 U7804 ( .A1(n6880), .A2(n6879), .A3(n6878), .ZN(n6888) );
  AOI22_X1 U7805 ( .A1(n3683), .A2(keyinput87), .B1(keyinput74), .B2(n6882), 
        .ZN(n6881) );
  OAI221_X1 U7806 ( .B1(n3683), .B2(keyinput87), .C1(n6882), .C2(keyinput74), 
        .A(n6881), .ZN(n6887) );
  AOI22_X1 U7807 ( .A1(n6885), .A2(keyinput17), .B1(n6884), .B2(keyinput2), 
        .ZN(n6883) );
  OAI221_X1 U7808 ( .B1(n6885), .B2(keyinput17), .C1(n6884), .C2(keyinput2), 
        .A(n6883), .ZN(n6886) );
  NOR3_X1 U7809 ( .A1(n6888), .A2(n6887), .A3(n6886), .ZN(n6922) );
  AOI22_X1 U7810 ( .A1(n6891), .A2(keyinput41), .B1(n6890), .B2(keyinput103), 
        .ZN(n6889) );
  OAI221_X1 U7811 ( .B1(n6891), .B2(keyinput41), .C1(n6890), .C2(keyinput103), 
        .A(n6889), .ZN(n6904) );
  AOI22_X1 U7812 ( .A1(n6894), .A2(keyinput7), .B1(keyinput19), .B2(n6893), 
        .ZN(n6892) );
  OAI221_X1 U7813 ( .B1(n6894), .B2(keyinput7), .C1(n6893), .C2(keyinput19), 
        .A(n6892), .ZN(n6903) );
  AOI22_X1 U7814 ( .A1(n6897), .A2(keyinput70), .B1(keyinput20), .B2(n6896), 
        .ZN(n6895) );
  OAI221_X1 U7815 ( .B1(n6897), .B2(keyinput70), .C1(n6896), .C2(keyinput20), 
        .A(n6895), .ZN(n6902) );
  AOI22_X1 U7816 ( .A1(n6900), .A2(keyinput28), .B1(keyinput83), .B2(n6899), 
        .ZN(n6898) );
  OAI221_X1 U7817 ( .B1(n6900), .B2(keyinput28), .C1(n6899), .C2(keyinput83), 
        .A(n6898), .ZN(n6901) );
  NOR4_X1 U7818 ( .A1(n6904), .A2(n6903), .A3(n6902), .A4(n6901), .ZN(n6921)
         );
  AOI22_X1 U7819 ( .A1(n6907), .A2(keyinput50), .B1(n6906), .B2(keyinput15), 
        .ZN(n6905) );
  OAI221_X1 U7820 ( .B1(n6907), .B2(keyinput50), .C1(n6906), .C2(keyinput15), 
        .A(n6905), .ZN(n6919) );
  AOI22_X1 U7821 ( .A1(n6910), .A2(keyinput114), .B1(keyinput69), .B2(n6909), 
        .ZN(n6908) );
  OAI221_X1 U7822 ( .B1(n6910), .B2(keyinput114), .C1(n6909), .C2(keyinput69), 
        .A(n6908), .ZN(n6918) );
  AOI22_X1 U7823 ( .A1(n6913), .A2(keyinput37), .B1(n6912), .B2(keyinput95), 
        .ZN(n6911) );
  OAI221_X1 U7824 ( .B1(n6913), .B2(keyinput37), .C1(n6912), .C2(keyinput95), 
        .A(n6911), .ZN(n6917) );
  INV_X1 U7825 ( .A(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n6915) );
  AOI22_X1 U7826 ( .A1(n5491), .A2(keyinput26), .B1(n6915), .B2(keyinput58), 
        .ZN(n6914) );
  OAI221_X1 U7827 ( .B1(n5491), .B2(keyinput26), .C1(n6915), .C2(keyinput58), 
        .A(n6914), .ZN(n6916) );
  NOR4_X1 U7828 ( .A1(n6919), .A2(n6918), .A3(n6917), .A4(n6916), .ZN(n6920)
         );
  NAND4_X1 U7829 ( .A1(n6923), .A2(n6922), .A3(n6921), .A4(n6920), .ZN(n6924)
         );
  NOR3_X1 U7830 ( .A1(n6926), .A2(n6925), .A3(n6924), .ZN(n6965) );
  OAI22_X1 U7831 ( .A1(REIP_REG_9__SCAN_IN), .A2(keyinput27), .B1(keyinput25), 
        .B2(ADDRESS_REG_21__SCAN_IN), .ZN(n6927) );
  AOI221_X1 U7832 ( .B1(REIP_REG_9__SCAN_IN), .B2(keyinput27), .C1(
        ADDRESS_REG_21__SCAN_IN), .C2(keyinput25), .A(n6927), .ZN(n6934) );
  OAI22_X1 U7833 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(keyinput51), .B1(
        keyinput81), .B2(DATAWIDTH_REG_19__SCAN_IN), .ZN(n6928) );
  AOI221_X1 U7834 ( .B1(INSTQUEUE_REG_3__4__SCAN_IN), .B2(keyinput51), .C1(
        DATAWIDTH_REG_19__SCAN_IN), .C2(keyinput81), .A(n6928), .ZN(n6933) );
  OAI22_X1 U7835 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(keyinput127), 
        .B1(keyinput48), .B2(ADDRESS_REG_9__SCAN_IN), .ZN(n6929) );
  AOI221_X1 U7836 ( .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(keyinput127), 
        .C1(ADDRESS_REG_9__SCAN_IN), .C2(keyinput48), .A(n6929), .ZN(n6932) );
  OAI22_X1 U7837 ( .A1(EAX_REG_25__SCAN_IN), .A2(keyinput110), .B1(
        EAX_REG_27__SCAN_IN), .B2(keyinput8), .ZN(n6930) );
  AOI221_X1 U7838 ( .B1(EAX_REG_25__SCAN_IN), .B2(keyinput110), .C1(keyinput8), 
        .C2(EAX_REG_27__SCAN_IN), .A(n6930), .ZN(n6931) );
  NAND4_X1 U7839 ( .A1(n6934), .A2(n6933), .A3(n6932), .A4(n6931), .ZN(n6963)
         );
  OAI22_X1 U7840 ( .A1(INSTQUEUE_REG_15__2__SCAN_IN), .A2(keyinput3), .B1(
        keyinput93), .B2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n6935) );
  AOI221_X1 U7841 ( .B1(INSTQUEUE_REG_15__2__SCAN_IN), .B2(keyinput3), .C1(
        PHYADDRPOINTER_REG_30__SCAN_IN), .C2(keyinput93), .A(n6935), .ZN(n6942) );
  OAI22_X1 U7842 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(keyinput101), .B1(
        keyinput63), .B2(REIP_REG_4__SCAN_IN), .ZN(n6936) );
  AOI221_X1 U7843 ( .B1(INSTQUEUE_REG_11__5__SCAN_IN), .B2(keyinput101), .C1(
        REIP_REG_4__SCAN_IN), .C2(keyinput63), .A(n6936), .ZN(n6941) );
  OAI22_X1 U7844 ( .A1(INSTQUEUE_REG_4__7__SCAN_IN), .A2(keyinput13), .B1(
        keyinput21), .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n6937) );
  AOI221_X1 U7845 ( .B1(INSTQUEUE_REG_4__7__SCAN_IN), .B2(keyinput13), .C1(
        INSTQUEUE_REG_1__4__SCAN_IN), .C2(keyinput21), .A(n6937), .ZN(n6940)
         );
  OAI22_X1 U7846 ( .A1(INSTQUEUE_REG_14__2__SCAN_IN), .A2(keyinput119), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(keyinput122), .ZN(n6938) );
  AOI221_X1 U7847 ( .B1(INSTQUEUE_REG_14__2__SCAN_IN), .B2(keyinput119), .C1(
        keyinput122), .C2(ADDRESS_REG_24__SCAN_IN), .A(n6938), .ZN(n6939) );
  NAND4_X1 U7848 ( .A1(n6942), .A2(n6941), .A3(n6940), .A4(n6939), .ZN(n6962)
         );
  OAI22_X1 U7849 ( .A1(LWORD_REG_0__SCAN_IN), .A2(keyinput44), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(keyinput30), .ZN(n6943) );
  AOI221_X1 U7850 ( .B1(LWORD_REG_0__SCAN_IN), .B2(keyinput44), .C1(keyinput30), .C2(ADDRESS_REG_5__SCAN_IN), .A(n6943), .ZN(n6951) );
  OAI22_X1 U7851 ( .A1(EBX_REG_13__SCAN_IN), .A2(keyinput43), .B1(keyinput55), 
        .B2(BYTEENABLE_REG_1__SCAN_IN), .ZN(n6944) );
  AOI221_X1 U7852 ( .B1(EBX_REG_13__SCAN_IN), .B2(keyinput43), .C1(
        BYTEENABLE_REG_1__SCAN_IN), .C2(keyinput55), .A(n6944), .ZN(n6950) );
  OAI22_X1 U7853 ( .A1(n6946), .A2(keyinput5), .B1(keyinput6), .B2(
        REIP_REG_1__SCAN_IN), .ZN(n6945) );
  AOI221_X1 U7854 ( .B1(n6946), .B2(keyinput5), .C1(REIP_REG_1__SCAN_IN), .C2(
        keyinput6), .A(n6945), .ZN(n6949) );
  OAI22_X1 U7855 ( .A1(DATAO_REG_11__SCAN_IN), .A2(keyinput78), .B1(
        keyinput113), .B2(UWORD_REG_1__SCAN_IN), .ZN(n6947) );
  AOI221_X1 U7856 ( .B1(DATAO_REG_11__SCAN_IN), .B2(keyinput78), .C1(
        UWORD_REG_1__SCAN_IN), .C2(keyinput113), .A(n6947), .ZN(n6948) );
  NAND4_X1 U7857 ( .A1(n6951), .A2(n6950), .A3(n6949), .A4(n6948), .ZN(n6961)
         );
  OAI22_X1 U7858 ( .A1(UWORD_REG_0__SCAN_IN), .A2(keyinput121), .B1(
        DATAO_REG_9__SCAN_IN), .B2(keyinput32), .ZN(n6952) );
  AOI221_X1 U7859 ( .B1(UWORD_REG_0__SCAN_IN), .B2(keyinput121), .C1(
        keyinput32), .C2(DATAO_REG_9__SCAN_IN), .A(n6952), .ZN(n6959) );
  OAI22_X1 U7860 ( .A1(EBX_REG_16__SCAN_IN), .A2(keyinput67), .B1(keyinput54), 
        .B2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n6953) );
  AOI221_X1 U7861 ( .B1(EBX_REG_16__SCAN_IN), .B2(keyinput67), .C1(
        PHYADDRPOINTER_REG_15__SCAN_IN), .C2(keyinput54), .A(n6953), .ZN(n6958) );
  OAI22_X1 U7862 ( .A1(EAX_REG_16__SCAN_IN), .A2(keyinput90), .B1(keyinput98), 
        .B2(DATAO_REG_10__SCAN_IN), .ZN(n6954) );
  AOI221_X1 U7863 ( .B1(EAX_REG_16__SCAN_IN), .B2(keyinput90), .C1(
        DATAO_REG_10__SCAN_IN), .C2(keyinput98), .A(n6954), .ZN(n6957) );
  OAI22_X1 U7864 ( .A1(INSTQUEUE_REG_14__0__SCAN_IN), .A2(keyinput120), .B1(
        DATAWIDTH_REG_21__SCAN_IN), .B2(keyinput61), .ZN(n6955) );
  AOI221_X1 U7865 ( .B1(INSTQUEUE_REG_14__0__SCAN_IN), .B2(keyinput120), .C1(
        keyinput61), .C2(DATAWIDTH_REG_21__SCAN_IN), .A(n6955), .ZN(n6956) );
  NAND4_X1 U7866 ( .A1(n6959), .A2(n6958), .A3(n6957), .A4(n6956), .ZN(n6960)
         );
  NOR4_X1 U7867 ( .A1(n6963), .A2(n6962), .A3(n6961), .A4(n6960), .ZN(n6964)
         );
  NAND3_X1 U7868 ( .A1(n6966), .A2(n6965), .A3(n6964), .ZN(n6973) );
  OAI222_X1 U7869 ( .A1(n6971), .A2(n6970), .B1(n6969), .B2(n6968), .C1(n6967), 
        .C2(n3683), .ZN(n6972) );
  XNOR2_X1 U7870 ( .A(n6973), .B(n6972), .ZN(U2888) );
  AND2_X2 U4183 ( .A1(n4505), .A2(n3238), .ZN(n4050) );
  AND4_X1 U3658 ( .A1(n3451), .A2(n3450), .A3(n3449), .A4(n3448), .ZN(n3452)
         );
  CLKBUF_X1 U3660 ( .A(n4427), .Z(n3212) );
  OR2_X1 U3670 ( .A1(n5512), .A2(n5513), .ZN(n5252) );
  CLKBUF_X1 U3672 ( .A(n5627), .Z(n3213) );
  NAND2_X1 U3673 ( .A1(n5205), .A2(n5204), .ZN(n6083) );
  NAND2_X1 U3674 ( .A1(n6098), .A2(n4288), .ZN(n6093) );
  CLKBUF_X1 U3678 ( .A(n3643), .Z(n6267) );
  CLKBUF_X1 U3682 ( .A(n4584), .Z(n4829) );
  CLKBUF_X1 U3748 ( .A(n4234), .Z(n3202) );
  CLKBUF_X1 U3769 ( .A(n5404), .Z(n5409) );
  NAND2_X2 U3770 ( .A1(n3274), .A2(n3273), .ZN(n3401) );
  CLKBUF_X1 U3797 ( .A(n5433), .Z(n5443) );
  CLKBUF_X1 U3915 ( .A(n4589), .Z(n5084) );
  OR2_X1 U3939 ( .A1(n4703), .A2(n4702), .ZN(n6974) );
  AND2_X1 U3950 ( .A1(n5453), .A2(n3516), .ZN(n6975) );
endmodule

