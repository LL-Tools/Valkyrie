

module b21_C_2inp_gates_syn ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, 
        ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, 
        ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, 
        ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, 
        ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, P1_U3352, P1_U3351, 
        P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, 
        P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, 
        P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, 
        P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, 
        P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, 
        P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, 
        P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, 
        P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, 
        P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, 
        P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, 
        P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, 
        P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, 
        P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, 
        P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, 
        P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, 
        P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, 
        P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, 
        P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, 
        P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, 
        P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, 
        P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, 
        P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, 
        P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, 
        P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, 
        P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, 
        P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, 
        P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, 
        P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, 
        P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, 
        P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, 
        P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, 
        P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, 
        P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, 
        P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, 
        P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, 
        P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, 
        P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, 
        P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, 
        P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, 
        P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, 
        P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, 
        P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, 
        P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, 
        P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, 
        P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, 
        P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, 
        P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, 
        P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3152, P2_U3151, P2_U3966, keyinput127, keyinput126, 
        keyinput125, keyinput124, keyinput123, keyinput122, keyinput121, 
        keyinput120, keyinput119, keyinput118, keyinput117, keyinput116, 
        keyinput115, keyinput114, keyinput113, keyinput112, keyinput111, 
        keyinput110, keyinput109, keyinput108, keyinput107, keyinput106, 
        keyinput105, keyinput104, keyinput103, keyinput102, keyinput101, 
        keyinput100, keyinput99, keyinput98, keyinput97, keyinput96, 
        keyinput95, keyinput94, keyinput93, keyinput92, keyinput91, keyinput90, 
        keyinput89, keyinput88, keyinput87, keyinput86, keyinput85, keyinput84, 
        keyinput83, keyinput82, keyinput81, keyinput80, keyinput79, keyinput78, 
        keyinput77, keyinput76, keyinput75, keyinput74, keyinput73, keyinput72, 
        keyinput71, keyinput70, keyinput69, keyinput68, keyinput67, keyinput66, 
        keyinput65, keyinput64, keyinput63, keyinput62, keyinput61, keyinput60, 
        keyinput59, keyinput58, keyinput57, keyinput56, keyinput55, keyinput54, 
        keyinput53, keyinput52, keyinput51, keyinput50, keyinput49, keyinput48, 
        keyinput47, keyinput46, keyinput45, keyinput44, keyinput43, keyinput42, 
        keyinput41, keyinput40, keyinput39, keyinput38, keyinput37, keyinput36, 
        keyinput35, keyinput34, keyinput33, keyinput32, keyinput31, keyinput30, 
        keyinput29, keyinput28, keyinput27, keyinput26, keyinput25, keyinput24, 
        keyinput23, keyinput22, keyinput21, keyinput20, keyinput19, keyinput18, 
        keyinput17, keyinput16, keyinput15, keyinput14, keyinput13, keyinput12, 
        keyinput11, keyinput10, keyinput9, keyinput8, keyinput7, keyinput6, 
        keyinput5, keyinput4, keyinput3, keyinput2, keyinput1, keyinput0 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput127, keyinput126, keyinput125,
         keyinput124, keyinput123, keyinput122, keyinput121, keyinput120,
         keyinput119, keyinput118, keyinput117, keyinput116, keyinput115,
         keyinput114, keyinput113, keyinput112, keyinput111, keyinput110,
         keyinput109, keyinput108, keyinput107, keyinput106, keyinput105,
         keyinput104, keyinput103, keyinput102, keyinput101, keyinput100,
         keyinput99, keyinput98, keyinput97, keyinput96, keyinput95,
         keyinput94, keyinput93, keyinput92, keyinput91, keyinput90,
         keyinput89, keyinput88, keyinput87, keyinput86, keyinput85,
         keyinput84, keyinput83, keyinput82, keyinput81, keyinput80,
         keyinput79, keyinput78, keyinput77, keyinput76, keyinput75,
         keyinput74, keyinput73, keyinput72, keyinput71, keyinput70,
         keyinput69, keyinput68, keyinput67, keyinput66, keyinput65,
         keyinput64, keyinput63, keyinput62, keyinput61, keyinput60,
         keyinput59, keyinput58, keyinput57, keyinput56, keyinput55,
         keyinput54, keyinput53, keyinput52, keyinput51, keyinput50,
         keyinput49, keyinput48, keyinput47, keyinput46, keyinput45,
         keyinput44, keyinput43, keyinput42, keyinput41, keyinput40,
         keyinput39, keyinput38, keyinput37, keyinput36, keyinput35,
         keyinput34, keyinput33, keyinput32, keyinput31, keyinput30,
         keyinput29, keyinput28, keyinput27, keyinput26, keyinput25,
         keyinput24, keyinput23, keyinput22, keyinput21, keyinput20,
         keyinput19, keyinput18, keyinput17, keyinput16, keyinput15,
         keyinput14, keyinput13, keyinput12, keyinput11, keyinput10, keyinput9,
         keyinput8, keyinput7, keyinput6, keyinput5, keyinput4, keyinput3,
         keyinput2, keyinput1, keyinput0;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395,
         n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405,
         n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415,
         n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425,
         n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435,
         n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445,
         n4446, n4447, n4448, n4449, n4450, n4451, n4453, n4454, n4455, n4456,
         n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466,
         n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476,
         n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486,
         n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496,
         n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506,
         n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516,
         n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526,
         n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536,
         n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546,
         n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556,
         n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566,
         n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576,
         n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586,
         n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596,
         n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606,
         n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616,
         n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626,
         n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636,
         n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646,
         n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656,
         n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666,
         n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676,
         n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686,
         n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696,
         n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706,
         n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716,
         n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726,
         n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736,
         n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746,
         n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756,
         n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766,
         n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776,
         n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786,
         n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796,
         n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806,
         n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816,
         n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826,
         n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836,
         n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846,
         n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856,
         n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866,
         n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876,
         n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886,
         n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896,
         n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906,
         n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916,
         n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926,
         n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936,
         n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946,
         n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956,
         n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966,
         n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976,
         n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986,
         n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996,
         n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006,
         n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016,
         n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026,
         n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036,
         n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046,
         n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056,
         n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066,
         n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076,
         n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086,
         n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096,
         n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106,
         n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116,
         n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126,
         n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136,
         n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146,
         n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156,
         n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166,
         n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176,
         n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186,
         n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196,
         n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206,
         n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216,
         n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226,
         n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236,
         n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246,
         n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256,
         n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266,
         n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276,
         n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286,
         n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296,
         n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306,
         n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316,
         n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326,
         n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336,
         n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346,
         n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356,
         n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366,
         n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376,
         n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386,
         n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396,
         n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406,
         n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416,
         n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426,
         n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436,
         n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446,
         n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456,
         n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466,
         n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476,
         n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486,
         n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496,
         n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506,
         n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516,
         n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526,
         n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536,
         n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546,
         n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556,
         n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566,
         n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576,
         n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586,
         n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596,
         n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606,
         n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616,
         n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626,
         n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636,
         n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646,
         n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656,
         n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666,
         n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676,
         n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686,
         n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696,
         n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706,
         n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716,
         n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726,
         n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736,
         n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746,
         n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756,
         n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766,
         n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776,
         n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786,
         n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796,
         n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806,
         n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816,
         n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826,
         n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836,
         n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846,
         n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856,
         n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866,
         n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876,
         n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886,
         n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896,
         n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906,
         n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916,
         n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926,
         n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936,
         n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946,
         n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956,
         n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966,
         n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976,
         n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986,
         n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996,
         n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006,
         n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016,
         n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026,
         n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036,
         n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046,
         n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056,
         n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066,
         n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076,
         n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086,
         n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096,
         n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106,
         n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116,
         n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126,
         n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136,
         n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146,
         n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156,
         n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166,
         n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176,
         n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186,
         n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196,
         n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206,
         n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216,
         n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226,
         n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236,
         n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246,
         n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256,
         n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266,
         n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276,
         n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286,
         n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296,
         n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306,
         n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316,
         n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326,
         n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336,
         n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346,
         n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356,
         n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366,
         n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376,
         n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386,
         n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396,
         n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406,
         n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416,
         n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426,
         n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436,
         n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446,
         n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456,
         n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466,
         n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476,
         n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486,
         n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496,
         n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506,
         n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516,
         n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526,
         n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536,
         n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546,
         n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556,
         n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566,
         n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576,
         n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586,
         n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596,
         n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606,
         n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616,
         n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626,
         n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636,
         n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646,
         n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656,
         n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666,
         n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676,
         n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686,
         n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696,
         n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706,
         n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716,
         n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726,
         n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736,
         n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746,
         n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756,
         n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766,
         n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776,
         n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786,
         n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796,
         n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806,
         n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816,
         n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826,
         n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836,
         n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846,
         n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856,
         n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866,
         n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876,
         n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886,
         n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896,
         n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906,
         n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916,
         n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926,
         n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936,
         n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946,
         n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956,
         n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966,
         n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976,
         n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986,
         n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996,
         n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006,
         n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016,
         n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026,
         n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036,
         n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046,
         n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056,
         n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066,
         n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076,
         n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086,
         n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096,
         n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106,
         n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116,
         n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126,
         n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136,
         n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146,
         n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156,
         n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166,
         n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176,
         n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186,
         n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196,
         n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206,
         n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216,
         n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226,
         n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236,
         n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246,
         n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256,
         n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266,
         n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276,
         n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286,
         n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296,
         n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306,
         n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316,
         n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326,
         n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336,
         n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346,
         n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356,
         n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366,
         n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376,
         n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386,
         n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396,
         n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406,
         n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416,
         n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426,
         n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436,
         n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446,
         n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456,
         n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466,
         n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476,
         n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486,
         n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496,
         n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506,
         n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516,
         n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526,
         n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7536, n7537,
         n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547,
         n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557,
         n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567,
         n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577,
         n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587,
         n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597,
         n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607,
         n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617,
         n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627,
         n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637,
         n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647,
         n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657,
         n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667,
         n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677,
         n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687,
         n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697,
         n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707,
         n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717,
         n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727,
         n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737,
         n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747,
         n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757,
         n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767,
         n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777,
         n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787,
         n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797,
         n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807,
         n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817,
         n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827,
         n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837,
         n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847,
         n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857,
         n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867,
         n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877,
         n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887,
         n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897,
         n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907,
         n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917,
         n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927,
         n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937,
         n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947,
         n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957,
         n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967,
         n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977,
         n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987,
         n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997,
         n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007,
         n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017,
         n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027,
         n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037,
         n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047,
         n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057,
         n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067,
         n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077,
         n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087,
         n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097,
         n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107,
         n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117,
         n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127,
         n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137,
         n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147,
         n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157,
         n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167,
         n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177,
         n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187,
         n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197,
         n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207,
         n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217,
         n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227,
         n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237,
         n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247,
         n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257,
         n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267,
         n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277,
         n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287,
         n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297,
         n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307,
         n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317,
         n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327,
         n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337,
         n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347,
         n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357,
         n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367,
         n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377,
         n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387,
         n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397,
         n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407,
         n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417,
         n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427,
         n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437,
         n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447,
         n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457,
         n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467,
         n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477,
         n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487,
         n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497,
         n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507,
         n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517,
         n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527,
         n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537,
         n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547,
         n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557,
         n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567,
         n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577,
         n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587,
         n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597,
         n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607,
         n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617,
         n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627,
         n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637,
         n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647,
         n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657,
         n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667,
         n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677,
         n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8688,
         n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698,
         n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708,
         n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718,
         n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728,
         n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738,
         n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748,
         n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758,
         n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768,
         n8769, n8770, n8771, n8772, n8774, n8775, n8776, n8777, n8778, n8779,
         n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789,
         n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799,
         n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809,
         n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819,
         n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829,
         n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839,
         n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849,
         n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859,
         n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869,
         n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879,
         n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889,
         n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899,
         n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909,
         n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919,
         n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929,
         n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939,
         n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949,
         n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959,
         n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969,
         n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979,
         n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989,
         n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999,
         n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009,
         n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019,
         n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029,
         n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039,
         n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049,
         n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059,
         n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069,
         n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079,
         n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089,
         n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099,
         n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109,
         n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119,
         n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129,
         n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139,
         n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149,
         n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159,
         n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169,
         n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179,
         n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189,
         n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199,
         n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209,
         n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219,
         n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229,
         n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239,
         n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249,
         n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259,
         n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269,
         n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279,
         n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289,
         n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299,
         n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309,
         n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319,
         n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329,
         n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339,
         n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349,
         n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359,
         n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369,
         n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379,
         n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389,
         n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399,
         n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409,
         n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419,
         n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429,
         n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439,
         n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449,
         n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459,
         n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469,
         n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479,
         n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489,
         n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499,
         n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509,
         n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519,
         n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529,
         n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539,
         n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549,
         n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559,
         n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569,
         n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579,
         n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589,
         n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599,
         n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609,
         n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619,
         n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629,
         n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639,
         n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649,
         n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659,
         n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669,
         n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679,
         n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689,
         n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699,
         n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709,
         n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719,
         n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729,
         n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739,
         n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749,
         n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759,
         n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769,
         n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779,
         n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789,
         n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799,
         n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809,
         n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819,
         n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829,
         n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839,
         n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849,
         n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859,
         n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869,
         n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879,
         n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889,
         n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899,
         n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909,
         n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919,
         n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929,
         n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939,
         n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949,
         n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959,
         n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969,
         n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979,
         n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989,
         n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999,
         n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190;

  NAND2_X1 U4891 ( .A1(n6257), .A2(n6256), .ZN(n9306) );
  INV_X1 U4892 ( .A(n7887), .ZN(n7890) );
  NAND2_X1 U4894 ( .A1(n5754), .A2(n5756), .ZN(n8693) );
  CLKBUF_X1 U4895 ( .A(n5152), .Z(n7593) );
  NAND4_X2 U4896 ( .A1(n5078), .A2(n5077), .A3(n5076), .A4(n5075), .ZN(n7965)
         );
  AND2_X1 U4898 ( .A1(n5042), .A2(n5041), .ZN(n5152) );
  NAND2_X1 U4899 ( .A1(n5042), .A2(n7526), .ZN(n5129) );
  CLKBUF_X2 U4900 ( .A(n7875), .Z(n4478) );
  AND2_X1 U4901 ( .A1(n5824), .A2(n6829), .ZN(n8689) );
  OR2_X1 U4902 ( .A1(n6102), .A2(n6101), .ZN(n6133) );
  NAND2_X1 U4903 ( .A1(n7050), .A2(n9048), .ZN(n8889) );
  CLKBUF_X2 U4904 ( .A(n5088), .Z(n4387) );
  NAND2_X1 U4905 ( .A1(n6896), .A2(n4907), .ZN(n7117) );
  BUF_X1 U4906 ( .A(n5035), .Z(n5011) );
  INV_X1 U4907 ( .A(n9358), .ZN(n9210) );
  AND2_X1 U4908 ( .A1(n4555), .A2(n4553), .ZN(n8752) );
  INV_X1 U4909 ( .A(n8689), .ZN(n6278) );
  INV_X1 U4910 ( .A(n9387), .ZN(n9388) );
  BUF_X1 U4911 ( .A(n5129), .Z(n7598) );
  AOI21_X1 U4912 ( .B1(n6990), .B2(n8639), .A(n8638), .ZN(n8641) );
  INV_X1 U4913 ( .A(n5955), .ZN(n8866) );
  AND3_X1 U4914 ( .A1(n5188), .A2(n5187), .A3(n5186), .ZN(n10075) );
  XNOR2_X1 U4915 ( .A(n5752), .B(n5751), .ZN(n7565) );
  INV_X2 U4916 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  NAND2_X2 U4917 ( .A1(n7529), .A2(n7528), .ZN(n7527) );
  INV_X2 U4918 ( .A(n6824), .ZN(n9846) );
  NAND2_X1 U4919 ( .A1(n5754), .A2(n5756), .ZN(n4386) );
  NAND2_X1 U4920 ( .A1(n4592), .A2(n4771), .ZN(n9298) );
  AOI21_X2 U4921 ( .B1(n8091), .B2(n8092), .A(n7848), .ZN(n8073) );
  OAI21_X2 U4922 ( .B1(n8233), .B2(n4941), .A(n4939), .ZN(n8199) );
  AOI21_X2 U4923 ( .B1(n7570), .B2(n7910), .A(n7569), .ZN(n8233) );
  INV_X1 U4924 ( .A(n5639), .ZN(n5724) );
  CLKBUF_X3 U4925 ( .A(n5117), .Z(n5639) );
  XNOR2_X1 U4926 ( .A(n7962), .B(n7736), .ZN(n7899) );
  INV_X2 U4927 ( .A(n5845), .ZN(n6279) );
  NAND2_X1 U4928 ( .A1(n4477), .A2(n5570), .ZN(n7657) );
  NAND2_X1 U4929 ( .A1(n4733), .A2(n4422), .ZN(n9599) );
  OAI22_X1 U4930 ( .A1(n8106), .A2(n7844), .B1(n8134), .B2(n8294), .ZN(n8089)
         );
  NAND2_X1 U4931 ( .A1(n9270), .A2(n9277), .ZN(n4788) );
  NAND2_X1 U4932 ( .A1(n4895), .A2(n4894), .ZN(n5541) );
  MUX2_X1 U4933 ( .A(n8987), .B(n8986), .S(n8996), .Z(n8989) );
  OR2_X1 U4934 ( .A1(n8145), .A2(n8144), .ZN(n8148) );
  NAND2_X1 U4935 ( .A1(n6203), .A2(n6202), .ZN(n8770) );
  NAND2_X1 U4936 ( .A1(n7642), .A2(n5418), .ZN(n7652) );
  NAND2_X1 U4937 ( .A1(n4811), .A2(n4809), .ZN(n8239) );
  OAI21_X1 U4938 ( .B1(n9357), .B2(n9363), .A(n9233), .ZN(n9348) );
  AND2_X1 U4939 ( .A1(n8729), .A2(n6021), .ZN(n7488) );
  NAND2_X1 U4940 ( .A1(n7117), .A2(n4906), .ZN(n9911) );
  OR2_X1 U4941 ( .A1(n5615), .A2(n7704), .ZN(n5637) );
  AOI21_X1 U4942 ( .B1(n4585), .B2(n4957), .A(n4980), .ZN(n4584) );
  NAND2_X1 U4943 ( .A1(n7135), .A2(n7134), .ZN(n7136) );
  AND2_X2 U4944 ( .A1(n6887), .A2(n10028), .ZN(n8208) );
  NAND2_X1 U4945 ( .A1(n5987), .A2(n5986), .ZN(n9589) );
  OR2_X1 U4946 ( .A1(n7191), .A2(n4964), .ZN(n4961) );
  NAND2_X2 U4947 ( .A1(n7138), .A2(n9407), .ZN(n9425) );
  AND2_X1 U4948 ( .A1(n7078), .A2(n6826), .ZN(n7013) );
  INV_X1 U4949 ( .A(n7736), .ZN(n10070) );
  INV_X1 U4950 ( .A(n7082), .ZN(n9015) );
  OR2_X1 U4951 ( .A1(n5472), .A2(n8438), .ZN(n5495) );
  INV_X2 U4952 ( .A(n5825), .ZN(n8684) );
  NAND2_X1 U4953 ( .A1(n6747), .A2(n10055), .ZN(n7751) );
  AND3_X1 U4954 ( .A1(n5100), .A2(n5099), .A3(n5098), .ZN(n6773) );
  NOR2_X2 U4955 ( .A1(n6440), .A2(n7087), .ZN(n7081) );
  AND3_X1 U4956 ( .A1(n5073), .A2(n5072), .A3(n5071), .ZN(n6750) );
  NAND2_X1 U4957 ( .A1(n5797), .A2(n4996), .ZN(n9104) );
  INV_X1 U4958 ( .A(n5152), .ZN(n5619) );
  NAND3_X1 U4959 ( .A1(n5759), .A2(n5758), .A3(n5757), .ZN(n6677) );
  NAND4_X2 U4960 ( .A1(n5852), .A2(n5851), .A3(n5850), .A4(n5849), .ZN(n9103)
         );
  INV_X2 U4961 ( .A(n5129), .ZN(n5725) );
  NAND2_X1 U4962 ( .A1(n4908), .A2(n7526), .ZN(n5118) );
  CLKBUF_X1 U4963 ( .A(n5047), .Z(n7923) );
  OR2_X1 U4964 ( .A1(n5042), .A2(n7526), .ZN(n5117) );
  NAND2_X1 U4965 ( .A1(n7522), .A2(n7565), .ZN(n6162) );
  NAND2_X1 U4966 ( .A1(n5097), .A2(n5096), .ZN(n5109) );
  NAND2_X4 U4967 ( .A1(n6323), .A2(n9723), .ZN(n5838) );
  NAND2_X1 U4968 ( .A1(n8625), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5037) );
  CLKBUF_X1 U4969 ( .A(n6323), .Z(n9726) );
  AND2_X2 U4970 ( .A1(n5755), .A2(n7565), .ZN(n8814) );
  OR2_X1 U4971 ( .A1(n5038), .A2(n4613), .ZN(n5039) );
  OR2_X1 U4972 ( .A1(n5011), .A2(n4611), .ZN(n4610) );
  XNOR2_X1 U4973 ( .A(n5110), .B(n4674), .ZN(n5108) );
  AND2_X1 U4974 ( .A1(n5035), .A2(n5034), .ZN(n5038) );
  XNOR2_X1 U4975 ( .A(n5136), .B(SI_4_), .ZN(n5135) );
  NAND2_X1 U4976 ( .A1(n6085), .A2(n5761), .ZN(n6097) );
  OR2_X1 U4977 ( .A1(n5750), .A2(n6084), .ZN(n5752) );
  AND2_X1 U4978 ( .A1(n6043), .A2(n5760), .ZN(n6085) );
  INV_X2 U4979 ( .A(n9622), .ZN(n7433) );
  OAI21_X1 U4980 ( .B1(n7515), .B2(P1_DATAO_REG_4__SCAN_IN), .A(n4483), .ZN(
        n5136) );
  OR2_X1 U4981 ( .A1(n4478), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n4483) );
  AND2_X1 U4982 ( .A1(n5879), .A2(n4589), .ZN(n6043) );
  INV_X4 U4983 ( .A(n7875), .ZN(n7515) );
  AND2_X1 U4984 ( .A1(n5747), .A2(n4442), .ZN(n4796) );
  AND2_X2 U4985 ( .A1(n4990), .A2(n4982), .ZN(n4797) );
  AND2_X1 U4986 ( .A1(n4966), .A2(n5738), .ZN(n4965) );
  AND3_X1 U4987 ( .A1(n4790), .A2(n4789), .A3(n5742), .ZN(n4990) );
  AND2_X1 U4988 ( .A1(n4868), .A2(n4869), .ZN(n5230) );
  AND4_X1 U4989 ( .A1(n4870), .A2(n4998), .A3(n4871), .A4(n4867), .ZN(n4866)
         );
  INV_X1 U4990 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n6059) );
  INV_X1 U4991 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5781) );
  INV_X1 U4992 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5685) );
  INV_X1 U4993 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5682) );
  NOR2_X1 U4994 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n4790) );
  NOR2_X1 U4995 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n4789) );
  INV_X1 U4996 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n6125) );
  INV_X1 U4997 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5766) );
  INV_X1 U4998 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5345) );
  INV_X1 U4999 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5296) );
  NOR2_X1 U5000 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n4868) );
  NOR2_X1 U5001 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n4869) );
  INV_X1 U5002 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n4871) );
  INV_X1 U5003 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n4997) );
  INV_X1 U5004 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n4912) );
  OAI22_X2 U5005 ( .A1(n8199), .A2(n7571), .B1(n8211), .B2(n8229), .ZN(n8184)
         );
  INV_X1 U5006 ( .A(n6462), .ZN(n5088) );
  AOI21_X4 U5007 ( .B1(n9284), .B2(n9216), .A(n9215), .ZN(n9270) );
  AOI22_X2 U5008 ( .A1(n9298), .A2(n9305), .B1(n9288), .B2(n9302), .ZN(n9284)
         );
  NAND2_X1 U5009 ( .A1(n8143), .A2(n7628), .ZN(n4934) );
  INV_X1 U5010 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5742) );
  INV_X1 U5011 ( .A(n4517), .ZN(n4516) );
  INV_X1 U5012 ( .A(n4515), .ZN(n4514) );
  OAI21_X1 U5013 ( .B1(n4518), .B2(n4516), .A(n7826), .ZN(n4515) );
  AOI21_X1 U5014 ( .B1(n4851), .B2(n7851), .A(n7887), .ZN(n4845) );
  NAND2_X1 U5015 ( .A1(n7847), .A2(n4843), .ZN(n4851) );
  INV_X1 U5016 ( .A(n7848), .ZN(n4843) );
  NAND2_X1 U5017 ( .A1(n7854), .A2(n7853), .ZN(n4849) );
  INV_X1 U5018 ( .A(n5252), .ZN(n5002) );
  NAND2_X1 U5019 ( .A1(n7676), .A2(n5542), .ZN(n5571) );
  OR2_X1 U5020 ( .A1(n5541), .A2(n5540), .ZN(n5542) );
  OR2_X1 U5021 ( .A1(n8314), .A2(n7951), .ZN(n7827) );
  OR2_X1 U5022 ( .A1(n7495), .A2(n7910), .ZN(n4811) );
  OR2_X1 U5023 ( .A1(n7568), .A2(n8242), .ZN(n7807) );
  NAND2_X1 U5024 ( .A1(n4997), .A2(n4912), .ZN(n4911) );
  OR2_X1 U5025 ( .A1(n5825), .A2(n9850), .ZN(n5805) );
  NAND2_X1 U5026 ( .A1(n9433), .A2(n9423), .ZN(n4769) );
  AND2_X1 U5027 ( .A1(n4757), .A2(n4759), .ZN(n4755) );
  NAND2_X1 U5028 ( .A1(n4758), .A2(n9200), .ZN(n4757) );
  NOR2_X1 U5029 ( .A1(n9027), .A2(n4732), .ZN(n4731) );
  INV_X1 U5030 ( .A(n8826), .ZN(n4732) );
  NAND2_X1 U5031 ( .A1(n4437), .A2(n4391), .ZN(n4778) );
  NAND2_X1 U5032 ( .A1(n4405), .A2(n7338), .ZN(n4779) );
  NAND2_X1 U5033 ( .A1(n9855), .A2(n9103), .ZN(n8887) );
  NAND2_X1 U5034 ( .A1(n7019), .A2(n6836), .ZN(n9046) );
  NAND2_X1 U5035 ( .A1(n5628), .A2(n5627), .ZN(n5650) );
  INV_X1 U5036 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5771) );
  OAI21_X1 U5037 ( .B1(n5584), .B2(n5583), .A(n5587), .ZN(n5608) );
  NAND2_X1 U5038 ( .A1(n4686), .A2(n5509), .ZN(n5523) );
  NAND2_X1 U5039 ( .A1(n5507), .A2(n5508), .ZN(n4686) );
  NAND2_X1 U5040 ( .A1(n5464), .A2(n5463), .ZN(n5487) );
  AND2_X1 U5041 ( .A1(n5421), .A2(n5400), .ZN(n5419) );
  NOR2_X1 U5042 ( .A1(n4983), .A2(n4590), .ZN(n4589) );
  NAND2_X1 U5043 ( .A1(n5741), .A2(n4591), .ZN(n4590) );
  INV_X1 U5044 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n4591) );
  NAND2_X1 U5045 ( .A1(n4687), .A2(n4691), .ZN(n5343) );
  AOI21_X1 U5046 ( .B1(n4693), .B2(n4856), .A(n4692), .ZN(n4691) );
  INV_X1 U5047 ( .A(n4993), .ZN(n4692) );
  INV_X1 U5048 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5740) );
  AND2_X1 U5049 ( .A1(n4676), .A2(n4675), .ZN(n5110) );
  NAND2_X1 U5050 ( .A1(n7515), .A2(n6394), .ZN(n4675) );
  AND2_X1 U5051 ( .A1(n9912), .A2(n5244), .ZN(n4906) );
  NAND2_X1 U5052 ( .A1(n5512), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n5534) );
  OR3_X1 U5053 ( .A1(n7435), .A2(n7301), .A3(n7456), .ZN(n6342) );
  NAND2_X1 U5054 ( .A1(n7536), .A2(n8020), .ZN(n6761) );
  AND3_X1 U5055 ( .A1(n5538), .A2(n5537), .A3(n5536), .ZN(n7628) );
  CLKBUF_X1 U5057 ( .A(n5118), .Z(n5406) );
  NAND2_X1 U5058 ( .A1(n7974), .A2(n7975), .ZN(n7973) );
  NOR2_X1 U5059 ( .A1(n7929), .A2(n7862), .ZN(n7930) );
  AND2_X1 U5060 ( .A1(n5564), .A2(n5563), .ZN(n8094) );
  OR2_X1 U5061 ( .A1(n8302), .A2(n7628), .ZN(n7836) );
  INV_X1 U5062 ( .A(n4931), .ZN(n4930) );
  OAI21_X1 U5063 ( .B1(n8201), .B2(n7911), .A(n7826), .ZN(n8192) );
  AND2_X1 U5064 ( .A1(n8333), .A2(n7955), .ZN(n4945) );
  NAND2_X1 U5065 ( .A1(n6342), .A2(n10048), .ZN(n10037) );
  NAND2_X1 U5066 ( .A1(n5703), .A2(n5702), .ZN(n5705) );
  NAND2_X1 U5067 ( .A1(n5705), .A2(n5704), .ZN(n6423) );
  OR2_X1 U5068 ( .A1(n5703), .A2(n5702), .ZN(n5704) );
  INV_X1 U5069 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5031) );
  NAND2_X1 U5070 ( .A1(n5027), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5032) );
  INV_X1 U5071 ( .A(n4575), .ZN(n4571) );
  INV_X1 U5072 ( .A(n4976), .ZN(n4975) );
  AND2_X1 U5073 ( .A1(n4568), .A2(n4972), .ZN(n4567) );
  AOI21_X1 U5074 ( .B1(n4976), .B2(n4974), .A(n4973), .ZN(n4972) );
  NAND2_X1 U5075 ( .A1(n4570), .A2(n4576), .ZN(n4568) );
  INV_X1 U5076 ( .A(n6155), .ZN(n4974) );
  NAND2_X1 U5077 ( .A1(n6733), .A2(n5867), .ZN(n6987) );
  AND2_X1 U5078 ( .A1(n7000), .A2(n9321), .ZN(n6313) );
  INV_X1 U5079 ( .A(n7565), .ZN(n5756) );
  NAND2_X1 U5080 ( .A1(n4785), .A2(n4783), .ZN(n4782) );
  NAND2_X1 U5081 ( .A1(n4786), .A2(n9244), .ZN(n4783) );
  NAND2_X1 U5082 ( .A1(n4596), .A2(n4760), .ZN(n9386) );
  AOI21_X1 U5083 ( .B1(n4762), .B2(n4765), .A(n4425), .ZN(n4760) );
  NAND2_X1 U5084 ( .A1(n9442), .A2(n4762), .ZN(n4596) );
  AND2_X1 U5085 ( .A1(n4763), .A2(n9418), .ZN(n4762) );
  NAND2_X1 U5086 ( .A1(n4764), .A2(n4766), .ZN(n4763) );
  INV_X1 U5087 ( .A(n4767), .ZN(n4764) );
  INV_X1 U5088 ( .A(n4766), .ZN(n4765) );
  INV_X1 U5089 ( .A(n8869), .ZN(n6140) );
  OR2_X1 U5090 ( .A1(n8841), .A2(n8897), .ZN(n4725) );
  NAND2_X1 U5091 ( .A1(n6316), .A2(n9841), .ZN(n8710) );
  NAND2_X1 U5092 ( .A1(n6290), .A2(n5778), .ZN(n6315) );
  AND2_X1 U5093 ( .A1(n6288), .A2(n6287), .ZN(n5778) );
  NOR2_X1 U5094 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n4982) );
  AND2_X1 U5095 ( .A1(n5555), .A2(n5550), .ZN(n5553) );
  NAND2_X1 U5096 ( .A1(n4524), .A2(n5196), .ZN(n4522) );
  INV_X1 U5097 ( .A(n5838), .ZN(n6346) );
  INV_X1 U5098 ( .A(n8937), .ZN(n4488) );
  INV_X1 U5099 ( .A(n7819), .ZN(n4520) );
  AOI21_X1 U5100 ( .B1(n4514), .B2(n4516), .A(n4428), .ZN(n4512) );
  AOI21_X1 U5101 ( .B1(n7803), .B2(n7799), .A(n4814), .ZN(n7800) );
  AOI21_X1 U5102 ( .B1(n4506), .B2(n4505), .A(n7846), .ZN(n7850) );
  NAND2_X1 U5103 ( .A1(n7845), .A2(n7887), .ZN(n4505) );
  NAND2_X1 U5104 ( .A1(n4507), .A2(n8092), .ZN(n4506) );
  NOR2_X1 U5105 ( .A1(n4842), .A2(n4840), .ZN(n4839) );
  AND2_X1 U5106 ( .A1(n4845), .A2(n8059), .ZN(n4842) );
  NAND2_X1 U5107 ( .A1(n7849), .A2(n7887), .ZN(n4844) );
  NAND2_X1 U5108 ( .A1(n4850), .A2(n4848), .ZN(n4847) );
  NAND2_X1 U5109 ( .A1(n7855), .A2(n7887), .ZN(n4850) );
  INV_X1 U5110 ( .A(n4898), .ZN(n4897) );
  OAI21_X1 U5111 ( .B1(n4900), .B2(n4899), .A(n7627), .ZN(n4898) );
  INV_X1 U5112 ( .A(n4402), .ZN(n4899) );
  INV_X1 U5113 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n4867) );
  INV_X1 U5114 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n4998) );
  INV_X1 U5115 ( .A(n8060), .ZN(n7857) );
  OR2_X1 U5116 ( .A1(n9512), .A2(n9217), .ZN(n9002) );
  INV_X1 U5117 ( .A(n4682), .ZN(n4681) );
  OAI21_X1 U5118 ( .B1(n4684), .B2(n4683), .A(n5553), .ZN(n4682) );
  INV_X1 U5119 ( .A(n5545), .ZN(n4683) );
  INV_X1 U5120 ( .A(n5419), .ZN(n4831) );
  OAI21_X1 U5121 ( .B1(n7592), .B2(n8072), .A(n7853), .ZN(n4829) );
  OR2_X1 U5122 ( .A1(n5660), .A2(n5721), .ZN(n5723) );
  INV_X1 U5123 ( .A(n4829), .ZN(n4828) );
  AND2_X1 U5124 ( .A1(n4934), .A2(n7573), .ZN(n4932) );
  AOI21_X1 U5125 ( .B1(n7805), .B2(n4814), .A(n4813), .ZN(n4812) );
  INV_X1 U5126 ( .A(n7807), .ZN(n4813) );
  NAND2_X1 U5127 ( .A1(n7416), .A2(n4937), .ZN(n4936) );
  NOR2_X1 U5128 ( .A1(n7907), .A2(n4938), .ZN(n4937) );
  NOR2_X1 U5129 ( .A1(n9956), .A2(n7414), .ZN(n4542) );
  OR2_X1 U5130 ( .A1(n9993), .A2(n10075), .ZN(n7769) );
  INV_X1 U5131 ( .A(n6409), .ZN(n4481) );
  NOR2_X1 U5132 ( .A1(n6950), .A2(n7736), .ZN(n6949) );
  NAND2_X1 U5133 ( .A1(n4613), .A2(n5034), .ZN(n4608) );
  NAND2_X1 U5134 ( .A1(n5011), .A2(n5034), .ZN(n4609) );
  INV_X1 U5135 ( .A(n4947), .ZN(n4946) );
  NAND2_X1 U5136 ( .A1(n5684), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5703) );
  OR2_X1 U5137 ( .A1(n5401), .A2(n4947), .ZN(n5025) );
  INV_X1 U5138 ( .A(n5830), .ZN(n6260) );
  NAND2_X1 U5139 ( .A1(n4655), .A2(n4654), .ZN(n7260) );
  NAND2_X1 U5140 ( .A1(n9128), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4654) );
  INV_X1 U5141 ( .A(n9124), .ZN(n4655) );
  OR2_X1 U5142 ( .A1(n9507), .A2(n9261), .ZN(n8978) );
  AND2_X1 U5143 ( .A1(n9521), .A2(n9306), .ZN(n9215) );
  OR2_X1 U5144 ( .A1(n9524), .A2(n9288), .ZN(n9238) );
  NOR2_X1 U5145 ( .A1(n9539), .A2(n9368), .ZN(n4659) );
  NOR2_X1 U5146 ( .A1(n9199), .A2(n9574), .ZN(n4657) );
  INV_X1 U5147 ( .A(n8847), .ZN(n4707) );
  AND2_X1 U5148 ( .A1(n8929), .A2(n7459), .ZN(n8847) );
  OR2_X1 U5149 ( .A1(n9586), .A2(n7402), .ZN(n8929) );
  INV_X1 U5150 ( .A(n9026), .ZN(n8920) );
  OR2_X1 U5151 ( .A1(n9103), .A2(n9855), .ZN(n9049) );
  OAI21_X1 U5152 ( .B1(n9379), .B2(n9232), .A(n9231), .ZN(n9357) );
  NAND2_X1 U5153 ( .A1(n7521), .A2(n7520), .ZN(n7872) );
  NAND2_X1 U5154 ( .A1(n7514), .A2(n7513), .ZN(n7524) );
  NAND2_X1 U5155 ( .A1(n7512), .A2(n7511), .ZN(n7514) );
  NAND2_X1 U5156 ( .A1(n5652), .A2(n5651), .ZN(n7512) );
  NAND2_X1 U5157 ( .A1(n5650), .A2(n5649), .ZN(n5652) );
  OAI21_X1 U5158 ( .B1(n5608), .B2(n5607), .A(n5606), .ZN(n5626) );
  AND2_X1 U5159 ( .A1(n5877), .A2(n4795), .ZN(n4794) );
  AND2_X1 U5160 ( .A1(n5740), .A2(n6305), .ZN(n4795) );
  NAND2_X1 U5161 ( .A1(n5765), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5767) );
  AOI21_X1 U5162 ( .B1(n6097), .B2(P1_IR_REG_31__SCAN_IN), .A(n4578), .ZN(
        n4577) );
  NAND2_X1 U5163 ( .A1(n4579), .A2(n5769), .ZN(n4578) );
  OAI21_X1 U5164 ( .B1(n5487), .B2(n5486), .A(n5488), .ZN(n5507) );
  OAI21_X1 U5165 ( .B1(n5442), .B2(n5441), .A(n5440), .ZN(n5461) );
  INV_X1 U5166 ( .A(n5368), .ZN(n4835) );
  INV_X1 U5167 ( .A(n4834), .ZN(n4833) );
  OAI21_X1 U5168 ( .B1(n4837), .B2(n4398), .A(n5394), .ZN(n4834) );
  NAND2_X1 U5169 ( .A1(n5269), .A2(n4994), .ZN(n5271) );
  OAI21_X1 U5170 ( .B1(n7515), .B2(P1_DATAO_REG_6__SCAN_IN), .A(n4479), .ZN(
        n5182) );
  NAND2_X1 U5171 ( .A1(n7515), .A2(n8574), .ZN(n4479) );
  OAI21_X1 U5172 ( .B1(n7515), .B2(P1_DATAO_REG_5__SCAN_IN), .A(n4471), .ZN(
        n5164) );
  NAND2_X1 U5173 ( .A1(n7515), .A2(n6402), .ZN(n4471) );
  INV_X2 U5174 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5738) );
  NAND2_X2 U5175 ( .A1(n4605), .A2(n4604), .ZN(n7875) );
  NOR2_X1 U5176 ( .A1(n4887), .A2(n4883), .ZN(n4882) );
  INV_X1 U5177 ( .A(n7634), .ZN(n4883) );
  INV_X1 U5178 ( .A(n7701), .ZN(n4887) );
  NAND2_X1 U5179 ( .A1(n7701), .A2(n4886), .ZN(n4885) );
  INV_X1 U5180 ( .A(n7633), .ZN(n4886) );
  AND3_X1 U5181 ( .A1(n5116), .A2(n5115), .A3(n5114), .ZN(n6756) );
  AND2_X1 U5182 ( .A1(n9944), .A2(n9941), .ZN(n5123) );
  NAND2_X1 U5183 ( .A1(n5107), .A2(n5106), .ZN(n9942) );
  AND2_X1 U5184 ( .A1(n6705), .A2(n5127), .ZN(n4905) );
  AND2_X1 U5185 ( .A1(n5383), .A2(n5393), .ZN(n7713) );
  NAND2_X1 U5186 ( .A1(n7713), .A2(n7712), .ZN(n7711) );
  NAND2_X1 U5187 ( .A1(n5047), .A2(n7921), .ZN(n7939) );
  NAND2_X1 U5188 ( .A1(n5673), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5683) );
  AOI21_X1 U5189 ( .B1(n8130), .B2(n5724), .A(n5578), .ZN(n7840) );
  AND3_X1 U5190 ( .A1(n5519), .A2(n5518), .A3(n5517), .ZN(n7589) );
  AND4_X1 U5191 ( .A1(n5502), .A2(n5501), .A3(n5500), .A4(n5499), .ZN(n7951)
         );
  AND4_X1 U5192 ( .A1(n5161), .A2(n5160), .A3(n5159), .A4(n5158), .ZN(n7737)
         );
  NOR2_X1 U5193 ( .A1(n9644), .A2(n9645), .ZN(n9643) );
  NOR2_X1 U5194 ( .A1(n9643), .A2(n4501), .ZN(n9656) );
  NOR2_X1 U5195 ( .A1(n6482), .A2(n6465), .ZN(n4501) );
  OR2_X1 U5196 ( .A1(n9656), .A2(n9655), .ZN(n4500) );
  NOR2_X1 U5197 ( .A1(n6493), .A2(n4504), .ZN(n6474) );
  AND2_X1 U5198 ( .A1(n6469), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n4504) );
  OR2_X1 U5199 ( .A1(n6474), .A2(n6473), .ZN(n4503) );
  NAND2_X1 U5200 ( .A1(n7973), .A2(n6666), .ZN(n6668) );
  NAND2_X1 U5201 ( .A1(n6668), .A2(n6667), .ZN(n4496) );
  OR2_X1 U5202 ( .A1(n5324), .A2(P2_IR_REG_13__SCAN_IN), .ZN(n5344) );
  NOR2_X1 U5203 ( .A1(n8030), .A2(n4535), .ZN(n4534) );
  INV_X1 U5204 ( .A(n4536), .ZN(n4535) );
  NAND2_X1 U5205 ( .A1(n4702), .A2(n7854), .ZN(n4827) );
  OAI21_X1 U5206 ( .B1(n4829), .B2(n4703), .A(n8038), .ZN(n4702) );
  INV_X1 U5207 ( .A(n7592), .ZN(n4703) );
  AND2_X1 U5208 ( .A1(n8073), .A2(n8072), .ZN(n8075) );
  NAND2_X1 U5209 ( .A1(n8140), .A2(n4423), .ZN(n8077) );
  INV_X1 U5210 ( .A(n8282), .ZN(n4543) );
  NOR2_X1 U5211 ( .A1(n8077), .A2(n8274), .ZN(n8055) );
  AOI21_X1 U5212 ( .B1(n7591), .B2(n4805), .A(n4804), .ZN(n4803) );
  INV_X1 U5213 ( .A(n7727), .ZN(n4804) );
  NAND2_X1 U5214 ( .A1(n4439), .A2(n4934), .ZN(n4931) );
  NAND2_X1 U5215 ( .A1(n4476), .A2(n4932), .ZN(n4926) );
  AOI21_X1 U5216 ( .B1(n4931), .B2(n4929), .A(n4928), .ZN(n4927) );
  INV_X1 U5217 ( .A(n4932), .ZN(n4929) );
  AOI21_X1 U5218 ( .B1(n7588), .B2(n4820), .A(n4819), .ZN(n4818) );
  INV_X1 U5219 ( .A(n7827), .ZN(n4819) );
  INV_X1 U5220 ( .A(n8193), .ZN(n4820) );
  OR2_X1 U5221 ( .A1(n8192), .A2(n4821), .ZN(n4817) );
  INV_X1 U5222 ( .A(n7588), .ZN(n4821) );
  AOI21_X1 U5224 ( .B1(n8190), .B2(n8203), .A(n7572), .ZN(n8170) );
  NAND2_X1 U5225 ( .A1(n8192), .A2(n8193), .ZN(n8191) );
  NAND2_X1 U5226 ( .A1(n8239), .A2(n7587), .ZN(n4621) );
  NAND2_X1 U5227 ( .A1(n8224), .A2(n4942), .ZN(n4941) );
  INV_X1 U5228 ( .A(n4945), .ZN(n4942) );
  AND2_X1 U5229 ( .A1(n8233), .A2(n8236), .ZN(n8235) );
  OAI21_X1 U5230 ( .B1(n7302), .B2(n4636), .A(n4633), .ZN(n7495) );
  INV_X1 U5231 ( .A(n4637), .ZN(n4636) );
  AOI21_X1 U5232 ( .B1(n4637), .B2(n4635), .A(n4634), .ZN(n4633) );
  INV_X1 U5233 ( .A(n7791), .ZN(n4635) );
  OR2_X1 U5234 ( .A1(n5304), .A2(n5303), .ZN(n5331) );
  NAND2_X1 U5235 ( .A1(n5329), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5352) );
  INV_X1 U5236 ( .A(n5331), .ZN(n5329) );
  OR2_X1 U5237 ( .A1(n7414), .A2(n9953), .ZN(n7794) );
  AOI21_X1 U5238 ( .B1(n4618), .B2(n4620), .A(n4616), .ZN(n4615) );
  INV_X1 U5239 ( .A(n7784), .ZN(n4616) );
  NAND2_X1 U5240 ( .A1(n4617), .A2(n7779), .ZN(n7209) );
  NAND2_X1 U5241 ( .A1(n7147), .A2(n7900), .ZN(n4617) );
  CLKBUF_X1 U5242 ( .A(n7146), .Z(n4480) );
  OR2_X1 U5243 ( .A1(n10070), .A2(n7737), .ZN(n4922) );
  NAND2_X1 U5244 ( .A1(n7737), .A2(n10070), .ZN(n4921) );
  NAND2_X1 U5245 ( .A1(n7769), .A2(n7768), .ZN(n7099) );
  CLKBUF_X1 U5246 ( .A(n6948), .Z(n4482) );
  NAND3_X1 U5247 ( .A1(n5023), .A2(n5022), .A3(n5021), .ZN(n6748) );
  NAND2_X1 U5248 ( .A1(n7725), .A2(n7932), .ZN(n7925) );
  INV_X1 U5249 ( .A(n9995), .ZN(n9935) );
  INV_X1 U5250 ( .A(n7585), .ZN(n8265) );
  NAND2_X1 U5251 ( .A1(n5533), .A2(n5532), .ZN(n8302) );
  NAND2_X1 U5252 ( .A1(n5404), .A2(n5403), .ZN(n8333) );
  OR2_X1 U5253 ( .A1(n7925), .A2(n7923), .ZN(n10102) );
  AND2_X1 U5254 ( .A1(n5690), .A2(n5689), .ZN(n10036) );
  CLKBUF_X1 U5255 ( .A(n5732), .Z(n5733) );
  NOR2_X1 U5256 ( .A1(n5673), .A2(n5672), .ZN(n5677) );
  NAND2_X1 U5257 ( .A1(n5025), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5443) );
  AND2_X1 U5258 ( .A1(n5298), .A2(n5324), .ZN(n6815) );
  INV_X1 U5259 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5140) );
  NAND2_X1 U5260 ( .A1(n4955), .A2(n5965), .ZN(n4954) );
  INV_X1 U5261 ( .A(n4959), .ZN(n4955) );
  OR2_X1 U5262 ( .A1(n7541), .A2(n7540), .ZN(n4575) );
  INV_X1 U5263 ( .A(n4567), .ZN(n4566) );
  AOI21_X1 U5264 ( .B1(n4567), .B2(n4569), .A(n4565), .ZN(n4564) );
  INV_X1 U5265 ( .A(n8715), .ZN(n4565) );
  OR2_X1 U5266 ( .A1(n6215), .A2(n4562), .ZN(n4561) );
  INV_X1 U5267 ( .A(n8665), .ZN(n4562) );
  INV_X1 U5268 ( .A(n6725), .ZN(n4953) );
  AOI21_X1 U5269 ( .B1(n8684), .B2(n7030), .A(n5827), .ZN(n5828) );
  NAND2_X1 U5270 ( .A1(n8674), .A2(n6155), .ZN(n4978) );
  INV_X1 U5271 ( .A(n4963), .ZN(n4958) );
  AND2_X1 U5272 ( .A1(n4954), .A2(n4586), .ZN(n4585) );
  INV_X1 U5273 ( .A(n7329), .ZN(n4586) );
  OAI21_X1 U5274 ( .B1(n6714), .B2(n6715), .A(n6712), .ZN(n6675) );
  OR2_X1 U5275 ( .A1(n5907), .A2(n7003), .ZN(n4991) );
  NAND2_X1 U5276 ( .A1(n4560), .A2(n4554), .ZN(n4553) );
  INV_X1 U5277 ( .A(n8755), .ZN(n4554) );
  INV_X1 U5278 ( .A(n8736), .ZN(n4971) );
  NAND2_X1 U5279 ( .A1(n8736), .A2(n4970), .ZN(n4969) );
  INV_X1 U5280 ( .A(n6232), .ZN(n4970) );
  NAND2_X1 U5281 ( .A1(n5767), .A2(n5766), .ZN(n5789) );
  INV_X1 U5282 ( .A(n8693), .ZN(n6276) );
  INV_X1 U5283 ( .A(n5868), .ZN(n6446) );
  AND4_X1 U5284 ( .A1(n6095), .A2(n6094), .A3(n6093), .A4(n6092), .ZN(n8852)
         );
  OAI22_X1 U5285 ( .A1(n6162), .A2(n4949), .B1(n6007), .B2(n6366), .ZN(n4948)
         );
  OR2_X1 U5286 ( .A1(n8693), .A2(n7027), .ZN(n5816) );
  NAND2_X1 U5287 ( .A1(n6310), .A2(n6309), .ZN(n9043) );
  AOI21_X1 U5288 ( .B1(n9784), .B2(n4648), .A(n6592), .ZN(n4647) );
  INV_X1 U5289 ( .A(n6591), .ZN(n4648) );
  OR2_X1 U5290 ( .A1(n6590), .A2(n4649), .ZN(n4646) );
  NOR2_X1 U5291 ( .A1(n9159), .A2(n4470), .ZN(n9163) );
  OR2_X1 U5292 ( .A1(n9163), .A2(n9162), .ZN(n4642) );
  NAND2_X1 U5293 ( .A1(n4667), .A2(n4666), .ZN(n4665) );
  AOI21_X1 U5294 ( .B1(n4787), .B2(n9269), .A(n4434), .ZN(n4785) );
  AOI21_X1 U5295 ( .B1(n9286), .B2(n9242), .A(n9241), .ZN(n9278) );
  AND2_X1 U5296 ( .A1(n9299), .A2(n9295), .ZN(n9290) );
  NOR2_X1 U5297 ( .A1(n9318), .A2(n9524), .ZN(n9299) );
  NAND2_X1 U5298 ( .A1(n9312), .A2(n9214), .ZN(n4771) );
  NAND2_X1 U5299 ( .A1(n9393), .A2(n9230), .ZN(n9379) );
  NOR2_X1 U5300 ( .A1(n9387), .A2(n9551), .ZN(n9373) );
  AND2_X1 U5301 ( .A1(n9554), .A2(n9205), .ZN(n4595) );
  AOI22_X1 U5302 ( .A1(n9449), .A2(n9229), .B1(n9228), .B2(n9227), .ZN(n9394)
         );
  INV_X1 U5303 ( .A(n9561), .ZN(n9406) );
  AND2_X1 U5304 ( .A1(n4769), .A2(n9441), .ZN(n4767) );
  NAND2_X1 U5305 ( .A1(n4438), .A2(n4769), .ZN(n4766) );
  NAND2_X1 U5306 ( .A1(n4729), .A2(n4727), .ZN(n4726) );
  AND2_X1 U5307 ( .A1(n4731), .A2(n9226), .ZN(n4730) );
  NAND2_X1 U5308 ( .A1(n4728), .A2(n9226), .ZN(n4727) );
  AOI21_X1 U5309 ( .B1(n4751), .B2(n4754), .A(n4459), .ZN(n4749) );
  OR2_X1 U5310 ( .A1(n9199), .A2(n9200), .ZN(n9223) );
  NAND2_X1 U5311 ( .A1(n7461), .A2(n4731), .ZN(n9224) );
  NOR2_X1 U5312 ( .A1(n8827), .A2(n4709), .ZN(n4708) );
  AOI21_X1 U5313 ( .B1(n4775), .B2(n4777), .A(n4431), .ZN(n4772) );
  NOR2_X1 U5314 ( .A1(n7232), .A2(n4724), .ZN(n4723) );
  INV_X1 U5315 ( .A(n8900), .ZN(n4724) );
  INV_X1 U5316 ( .A(n8887), .ZN(n4742) );
  OR2_X1 U5317 ( .A1(n9043), .A2(n9087), .ZN(n9422) );
  AND2_X1 U5318 ( .A1(n6309), .A2(n7000), .ZN(n6916) );
  AND2_X1 U5319 ( .A1(n6440), .A2(n7030), .ZN(n7079) );
  NAND2_X1 U5320 ( .A1(n7082), .A2(n7081), .ZN(n7080) );
  INV_X1 U5321 ( .A(n9422), .ZN(n9484) );
  INV_X1 U5322 ( .A(n9510), .ZN(n4734) );
  NAND2_X1 U5323 ( .A1(n6271), .A2(n6270), .ZN(n9514) );
  AND3_X1 U5324 ( .A1(n5924), .A2(n5923), .A3(n5922), .ZN(n9876) );
  INV_X1 U5325 ( .A(n9892), .ZN(n9881) );
  NOR2_X1 U5326 ( .A1(n8710), .A2(n6648), .ZN(n6908) );
  NAND2_X1 U5327 ( .A1(n6308), .A2(n9069), .ZN(n6910) );
  XNOR2_X1 U5328 ( .A(n5749), .B(P1_IR_REG_30__SCAN_IN), .ZN(n5755) );
  NAND2_X1 U5329 ( .A1(n9620), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5749) );
  NOR2_X1 U5330 ( .A1(n4711), .A2(n4400), .ZN(n4710) );
  NAND2_X1 U5331 ( .A1(n4981), .A2(n4712), .ZN(n4711) );
  NAND2_X1 U5332 ( .A1(n4794), .A2(n4796), .ZN(n4716) );
  INV_X1 U5333 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5751) );
  XNOR2_X1 U5334 ( .A(n7524), .B(n7523), .ZN(n8867) );
  XNOR2_X1 U5335 ( .A(n4792), .B(n5779), .ZN(n6323) );
  NAND2_X1 U5336 ( .A1(n4793), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4792) );
  NAND2_X1 U5337 ( .A1(n5780), .A2(n5781), .ZN(n4793) );
  XNOR2_X1 U5338 ( .A(n5773), .B(P1_IR_REG_26__SCAN_IN), .ZN(n6290) );
  NOR2_X1 U5339 ( .A1(n5543), .A2(n4685), .ZN(n4684) );
  INV_X1 U5340 ( .A(n5528), .ZN(n4685) );
  NAND2_X1 U5341 ( .A1(n5525), .A2(n5524), .ZN(n4862) );
  XNOR2_X1 U5342 ( .A(n6306), .B(n6305), .ZN(n7274) );
  NAND2_X1 U5343 ( .A1(n4836), .A2(n5368), .ZN(n5396) );
  NAND2_X1 U5344 ( .A1(n5343), .A2(n4837), .ZN(n4836) );
  NAND2_X1 U5345 ( .A1(n4990), .A2(n4984), .ZN(n4983) );
  XNOR2_X1 U5346 ( .A(n5269), .B(n4994), .ZN(n6427) );
  NAND2_X1 U5347 ( .A1(n4853), .A2(n4852), .ZN(n5163) );
  AOI21_X1 U5348 ( .B1(n5135), .B2(n4854), .A(n4406), .ZN(n4853) );
  NAND2_X1 U5349 ( .A1(n6084), .A2(n4653), .ZN(n4652) );
  INV_X1 U5350 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n4653) );
  NOR2_X1 U5351 ( .A1(n9680), .A2(n10164), .ZN(n9681) );
  NOR2_X1 U5352 ( .A1(n9685), .A2(n10161), .ZN(n9686) );
  AND2_X1 U5353 ( .A1(n5194), .A2(n5173), .ZN(n4889) );
  NAND2_X1 U5354 ( .A1(n5349), .A2(n5348), .ZN(n7497) );
  AND2_X1 U5355 ( .A1(n7117), .A2(n5244), .ZN(n9913) );
  NAND2_X1 U5356 ( .A1(n6851), .A2(n5195), .ZN(n6898) );
  NAND2_X1 U5357 ( .A1(n6898), .A2(n6897), .ZN(n6896) );
  INV_X1 U5358 ( .A(n8159), .ZN(n8307) );
  NAND2_X1 U5359 ( .A1(n5581), .A2(n5580), .ZN(n7635) );
  NAND2_X1 U5360 ( .A1(n5592), .A2(n5591), .ZN(n8289) );
  AND4_X1 U5361 ( .A1(n5414), .A2(n5413), .A3(n5412), .A4(n5411), .ZN(n8228)
         );
  AND4_X1 U5362 ( .A1(n5357), .A2(n5356), .A3(n5355), .A4(n5354), .ZN(n7716)
         );
  NAND2_X1 U5363 ( .A1(n5720), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9966) );
  INV_X1 U5364 ( .A(n9949), .ZN(n7709) );
  AND2_X1 U5365 ( .A1(n5708), .A2(n10024), .ZN(n9957) );
  INV_X1 U5366 ( .A(n7568), .ZN(n9697) );
  INV_X1 U5367 ( .A(n10037), .ZN(n7943) );
  AND2_X1 U5368 ( .A1(n6762), .A2(n5735), .ZN(n9992) );
  OAI21_X1 U5369 ( .B1(n7922), .B2(n7923), .A(n4530), .ZN(n4529) );
  OR2_X1 U5370 ( .A1(n7920), .A2(n7921), .ZN(n4530) );
  XNOR2_X1 U5371 ( .A(n4801), .B(n8020), .ZN(n4800) );
  AOI21_X1 U5372 ( .B1(n4698), .B2(n4697), .A(n7937), .ZN(n4801) );
  NAND2_X1 U5373 ( .A1(n7936), .A2(n7935), .ZN(n4697) );
  AOI21_X1 U5374 ( .B1(n4700), .B2(n4699), .A(n7934), .ZN(n4698) );
  XNOR2_X1 U5375 ( .A(n5683), .B(P2_IR_REG_22__SCAN_IN), .ZN(n5048) );
  AND2_X1 U5376 ( .A1(n4500), .A2(n4499), .ZN(n6539) );
  NAND2_X1 U5377 ( .A1(n9658), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n4499) );
  OAI22_X1 U5378 ( .A1(n8018), .A2(n9972), .B1(n8019), .B2(n9970), .ZN(n4494)
         );
  OAI21_X1 U5379 ( .B1(n8017), .B2(n9972), .A(n4411), .ZN(n4492) );
  OAI21_X1 U5380 ( .B1(n8022), .B2(n4864), .A(n8021), .ZN(n4490) );
  INV_X1 U5381 ( .A(n10001), .ZN(n8071) );
  NAND2_X1 U5382 ( .A1(n5008), .A2(n4613), .ZN(n4612) );
  OR2_X1 U5383 ( .A1(n5010), .A2(n5008), .ZN(n4607) );
  INV_X1 U5384 ( .A(n9096), .ZN(n7411) );
  INV_X1 U5385 ( .A(n7380), .ZN(n7351) );
  INV_X1 U5386 ( .A(n9392), .ZN(n9554) );
  OR2_X1 U5387 ( .A1(n8728), .A2(n4979), .ZN(n8729) );
  OR2_X1 U5388 ( .A1(n8726), .A2(n8727), .ZN(n4979) );
  NAND2_X1 U5389 ( .A1(n6025), .A2(n6024), .ZN(n9579) );
  INV_X1 U5390 ( .A(n6313), .ZN(n9085) );
  INV_X1 U5391 ( .A(n8852), .ZN(n9467) );
  AND2_X1 U5392 ( .A1(n4748), .A2(n4747), .ZN(n4746) );
  NAND2_X1 U5393 ( .A1(n4745), .A2(n5756), .ZN(n4748) );
  AOI21_X1 U5394 ( .B1(n9623), .B2(n8866), .A(n8808), .ZN(n9498) );
  NAND2_X1 U5395 ( .A1(n4738), .A2(n4735), .ZN(n9510) );
  AOI21_X1 U5396 ( .B1(n9486), .B2(n4737), .A(n4736), .ZN(n4735) );
  OAI21_X1 U5397 ( .B1(n9259), .B2(n9260), .A(n9489), .ZN(n4738) );
  NOR2_X1 U5398 ( .A1(n9261), .A2(n9422), .ZN(n4736) );
  NAND2_X1 U5399 ( .A1(n9253), .A2(n4593), .ZN(n9513) );
  NAND2_X1 U5400 ( .A1(n4788), .A2(n4787), .ZN(n9253) );
  NAND2_X1 U5401 ( .A1(n4788), .A2(n4407), .ZN(n4594) );
  AND2_X1 U5402 ( .A1(n6205), .A2(n6204), .ZN(n9333) );
  OR2_X1 U5403 ( .A1(n9843), .A2(n6909), .ZN(n9407) );
  XNOR2_X1 U5404 ( .A(n5791), .B(n5764), .ZN(n9321) );
  NOR2_X1 U5405 ( .A1(n10163), .A2(n10162), .ZN(n10161) );
  NOR2_X1 U5406 ( .A1(n10181), .A2(n10180), .ZN(n10179) );
  NAND2_X1 U5407 ( .A1(n4488), .A2(n4409), .ZN(n4487) );
  NAND2_X1 U5408 ( .A1(n7792), .A2(n4526), .ZN(n4525) );
  AND2_X1 U5409 ( .A1(n7794), .A2(n7887), .ZN(n4526) );
  AND2_X1 U5410 ( .A1(n4520), .A2(n4447), .ZN(n4518) );
  NAND2_X1 U5411 ( .A1(n4520), .A2(n4414), .ZN(n4517) );
  INV_X1 U5412 ( .A(n4510), .ZN(n4509) );
  OAI21_X1 U5413 ( .B1(n4512), .B2(n7828), .A(n7827), .ZN(n4510) );
  INV_X1 U5414 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5000) );
  INV_X1 U5415 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n4999) );
  AOI21_X1 U5416 ( .B1(n8924), .B2(n9223), .A(n4472), .ZN(n8844) );
  INV_X1 U5417 ( .A(n8843), .ZN(n4472) );
  AND2_X1 U5418 ( .A1(n4390), .A2(n7930), .ZN(n4826) );
  INV_X1 U5419 ( .A(n7930), .ZN(n4825) );
  AND2_X1 U5420 ( .A1(n4846), .A2(n4841), .ZN(n7859) );
  NOR2_X1 U5421 ( .A1(n7856), .A2(n4847), .ZN(n4846) );
  INV_X1 U5422 ( .A(n4922), .ZN(n4919) );
  INV_X1 U5423 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n8351) );
  INV_X1 U5424 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n8349) );
  NOR2_X1 U5425 ( .A1(n8297), .A2(n8294), .ZN(n4544) );
  NAND2_X1 U5426 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_28__SCAN_IN), 
        .ZN(n4611) );
  AND3_X1 U5427 ( .A1(n4872), .A2(n5682), .A3(n5685), .ZN(n5007) );
  NAND2_X1 U5428 ( .A1(n5003), .A2(n8493), .ZN(n4947) );
  INV_X1 U5429 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5003) );
  NAND2_X1 U5430 ( .A1(n4580), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4579) );
  INV_X1 U5431 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n5423) );
  INV_X1 U5432 ( .A(SI_15_), .ZN(n5371) );
  NOR2_X1 U5433 ( .A1(n4857), .A2(n4689), .ZN(n4688) );
  INV_X1 U5434 ( .A(n5246), .ZN(n4689) );
  INV_X1 U5435 ( .A(n4694), .ZN(n4693) );
  NAND2_X1 U5436 ( .A1(n4859), .A2(n5287), .ZN(n4858) );
  INV_X1 U5437 ( .A(n5315), .ZN(n4859) );
  NAND2_X1 U5438 ( .A1(n5245), .A2(n4992), .ZN(n5247) );
  AOI21_X1 U5439 ( .B1(n4897), .B2(n4899), .A(n4458), .ZN(n4894) );
  NAND2_X1 U5440 ( .A1(n7618), .A2(n4897), .ZN(n4895) );
  XNOR2_X1 U5441 ( .A(n5669), .B(n6750), .ZN(n5079) );
  INV_X1 U5442 ( .A(n5669), .ZN(n5635) );
  AND2_X1 U5443 ( .A1(n5082), .A2(n5062), .ZN(n4878) );
  NOR2_X1 U5444 ( .A1(n4701), .A2(n4823), .ZN(n7933) );
  OAI21_X1 U5445 ( .B1(n4827), .B2(n4825), .A(n4824), .ZN(n4823) );
  AND2_X1 U5446 ( .A1(n4826), .A2(n8073), .ZN(n4701) );
  INV_X1 U5447 ( .A(n7929), .ZN(n4824) );
  INV_X1 U5448 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n4870) );
  NOR2_X1 U5449 ( .A1(n8265), .A2(n8272), .ZN(n4536) );
  NAND2_X1 U5450 ( .A1(n5634), .A2(n4419), .ZN(n7853) );
  OR2_X1 U5451 ( .A1(n8294), .A2(n8094), .ZN(n7727) );
  INV_X1 U5452 ( .A(n7591), .ZN(n4806) );
  INV_X1 U5453 ( .A(n4807), .ZN(n4805) );
  AND2_X1 U5454 ( .A1(n7727), .A2(n7726), .ZN(n7844) );
  NOR2_X1 U5455 ( .A1(n8126), .A2(n4808), .ZN(n4807) );
  INV_X1 U5456 ( .A(n7836), .ZN(n4808) );
  OR2_X1 U5457 ( .A1(n5534), .A2(n7681), .ZN(n5572) );
  NAND2_X1 U5458 ( .A1(n4548), .A2(n8190), .ZN(n4547) );
  INV_X1 U5459 ( .A(n4549), .ZN(n4548) );
  NAND2_X1 U5460 ( .A1(n8211), .A2(n4944), .ZN(n4549) );
  INV_X1 U5461 ( .A(n7799), .ZN(n4634) );
  AND2_X1 U5462 ( .A1(n7907), .A2(n7794), .ZN(n4637) );
  NAND2_X1 U5463 ( .A1(n7302), .A2(n7791), .ZN(n7419) );
  INV_X1 U5464 ( .A(n4619), .ZN(n4618) );
  OAI21_X1 U5465 ( .B1(n7900), .B2(n4620), .A(n7786), .ZN(n4619) );
  AND2_X1 U5466 ( .A1(n7099), .A2(n4918), .ZN(n4916) );
  AND2_X1 U5467 ( .A1(n4918), .A2(n4920), .ZN(n4914) );
  INV_X1 U5468 ( .A(n4921), .ZN(n4920) );
  AND3_X1 U5469 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .A3(P2_REG3_REG_5__SCAN_IN), .ZN(n5153) );
  NAND2_X1 U5470 ( .A1(n8140), .A2(n4404), .ZN(n8096) );
  AND2_X1 U5471 ( .A1(n8140), .A2(n4544), .ZN(n8116) );
  AOI21_X1 U5472 ( .B1(n10036), .B2(n10046), .A(n10047), .ZN(n6745) );
  NAND2_X1 U5473 ( .A1(n5028), .A2(n5024), .ZN(n5673) );
  INV_X1 U5474 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5024) );
  INV_X1 U5475 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5026) );
  OR2_X1 U5476 ( .A1(n5184), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n5206) );
  AOI21_X1 U5477 ( .B1(n7488), .B2(n7484), .A(n7485), .ZN(n6076) );
  OR2_X1 U5478 ( .A1(n5825), .A2(n9846), .ZN(n5842) );
  INV_X1 U5479 ( .A(n6170), .ZN(n4973) );
  INV_X1 U5480 ( .A(n5945), .ZN(n4964) );
  OR2_X1 U5481 ( .A1(n8671), .A2(n8672), .ZN(n6155) );
  NAND2_X1 U5482 ( .A1(n7191), .A2(n4964), .ZN(n4963) );
  OR2_X1 U5483 ( .A1(n6986), .A2(n5906), .ZN(n5889) );
  NOR2_X1 U5484 ( .A1(n5904), .A2(n5903), .ZN(n5910) );
  NOR2_X1 U5485 ( .A1(n8755), .A2(n4557), .ZN(n4556) );
  INV_X1 U5486 ( .A(n4561), .ZN(n4557) );
  INV_X1 U5487 ( .A(n6315), .ZN(n6344) );
  NOR2_X1 U5488 ( .A1(n9809), .A2(n9810), .ZN(n9811) );
  OR2_X1 U5489 ( .A1(n9514), .A2(n9289), .ZN(n9257) );
  INV_X1 U5490 ( .A(n9223), .ZN(n4728) );
  AOI21_X1 U5491 ( .B1(n4778), .B2(n4776), .A(n4426), .ZN(n4775) );
  INV_X1 U5492 ( .A(n4401), .ZN(n4776) );
  INV_X1 U5493 ( .A(n4778), .ZN(n4777) );
  NAND2_X1 U5494 ( .A1(n4741), .A2(n8887), .ZN(n4740) );
  INV_X1 U5495 ( .A(n4743), .ZN(n4741) );
  NOR2_X1 U5496 ( .A1(n7133), .A2(n7184), .ZN(n4661) );
  NOR2_X1 U5497 ( .A1(n7070), .A2(n7074), .ZN(n7069) );
  NOR2_X1 U5498 ( .A1(n8892), .A2(n4744), .ZN(n4743) );
  INV_X1 U5499 ( .A(n9048), .ZN(n4744) );
  NOR2_X1 U5500 ( .A1(n7086), .A2(n7018), .ZN(n6843) );
  NAND2_X1 U5501 ( .A1(n7037), .A2(n4598), .ZN(n4597) );
  AND2_X1 U5502 ( .A1(n7061), .A2(n4599), .ZN(n4598) );
  NAND2_X1 U5503 ( .A1(n6308), .A2(n9356), .ZN(n8995) );
  XNOR2_X1 U5504 ( .A(n7872), .B(n7871), .ZN(n7869) );
  AND2_X1 U5505 ( .A1(n7520), .A2(n7519), .ZN(n7523) );
  INV_X1 U5506 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5779) );
  AND2_X1 U5507 ( .A1(n5651), .A2(n5632), .ZN(n5649) );
  AND2_X1 U5508 ( .A1(n5627), .A2(n5612), .ZN(n5625) );
  NAND2_X1 U5509 ( .A1(n4797), .A2(n4712), .ZN(n4714) );
  NAND2_X1 U5510 ( .A1(n4679), .A2(n4677), .ZN(n5584) );
  AOI21_X1 U5511 ( .B1(n4681), .B2(n4683), .A(n4678), .ZN(n4677) );
  INV_X1 U5512 ( .A(n5555), .ZN(n4678) );
  NAND2_X1 U5513 ( .A1(n5422), .A2(n5421), .ZN(n5442) );
  NAND2_X1 U5514 ( .A1(n4832), .A2(n4830), .ZN(n5422) );
  AOI21_X1 U5515 ( .B1(n4833), .B2(n4398), .A(n4831), .ZN(n4830) );
  NOR2_X1 U5516 ( .A1(n5369), .A2(n4838), .ZN(n4837) );
  INV_X1 U5517 ( .A(n5342), .ZN(n4838) );
  NOR2_X1 U5518 ( .A1(n4858), .A2(n4695), .ZN(n4694) );
  INV_X1 U5519 ( .A(n4994), .ZN(n4695) );
  NOR2_X1 U5520 ( .A1(n5288), .A2(n4861), .ZN(n4860) );
  INV_X1 U5521 ( .A(n5270), .ZN(n4861) );
  OR2_X1 U5522 ( .A1(n4412), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n5967) );
  INV_X1 U5523 ( .A(n5111), .ZN(n4854) );
  OAI21_X2 U5524 ( .B1(P1_ADDR_REG_19__SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        n4864), .ZN(n4604) );
  NAND2_X1 U5525 ( .A1(n4863), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n4605) );
  INV_X1 U5526 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5013) );
  AND2_X1 U5527 ( .A1(n5153), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5174) );
  NAND2_X1 U5528 ( .A1(n4891), .A2(n4890), .ZN(n7473) );
  AND2_X1 U5529 ( .A1(n5363), .A2(n5340), .ZN(n4890) );
  NAND2_X1 U5530 ( .A1(n7371), .A2(n7372), .ZN(n4891) );
  NAND2_X1 U5531 ( .A1(n6760), .A2(n7932), .ZN(n5033) );
  NOR2_X1 U5532 ( .A1(n7670), .A2(n4901), .ZN(n4900) );
  INV_X1 U5533 ( .A(n5485), .ZN(n4901) );
  NOR2_X1 U5534 ( .A1(n5210), .A2(n6899), .ZN(n5235) );
  INV_X1 U5535 ( .A(n5495), .ZN(n5494) );
  XNOR2_X1 U5536 ( .A(n5079), .B(n5080), .ZN(n7689) );
  INV_X1 U5537 ( .A(n5448), .ZN(n5446) );
  NAND2_X1 U5538 ( .A1(n7933), .A2(n8264), .ZN(n4700) );
  NOR2_X1 U5539 ( .A1(n8025), .A2(n7932), .ZN(n4699) );
  AND2_X1 U5540 ( .A1(n5601), .A2(n5600), .ZN(n7702) );
  INV_X1 U5541 ( .A(n6342), .ZN(n6460) );
  NAND2_X1 U5542 ( .A1(n5152), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5045) );
  OR2_X1 U5543 ( .A1(n5118), .A2(n5051), .ZN(n5052) );
  AND2_X1 U5544 ( .A1(n4503), .A2(n4502), .ZN(n6560) );
  NAND2_X1 U5545 ( .A1(n6505), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n4502) );
  NOR2_X1 U5546 ( .A1(n6560), .A2(n6559), .ZN(n6558) );
  CLKBUF_X1 U5547 ( .A(n5252), .Z(n5253) );
  NAND2_X1 U5548 ( .A1(n6684), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n4495) );
  NAND2_X1 U5549 ( .A1(n7984), .A2(n4498), .ZN(n7987) );
  OR2_X1 U5550 ( .A1(n7985), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n4498) );
  NOR2_X1 U5551 ( .A1(n7987), .A2(n7986), .ZN(n7995) );
  NOR2_X1 U5552 ( .A1(n7995), .A2(n4497), .ZN(n7997) );
  AND2_X1 U5553 ( .A1(n7996), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n4497) );
  NAND2_X1 U5554 ( .A1(n7997), .A2(n7998), .ZN(n8007) );
  AND2_X1 U5555 ( .A1(n5723), .A2(n5661), .ZN(n8046) );
  OAI21_X1 U5556 ( .B1(n8073), .B2(n7592), .A(n4828), .ZN(n8039) );
  NOR2_X1 U5557 ( .A1(n8042), .A2(n8241), .ZN(n4629) );
  NAND2_X1 U5558 ( .A1(n7852), .A2(n7853), .ZN(n8060) );
  NAND2_X1 U5559 ( .A1(n8133), .A2(n7591), .ZN(n8110) );
  NAND2_X1 U5560 ( .A1(n4923), .A2(n4925), .ZN(n8106) );
  AOI21_X1 U5561 ( .B1(n4927), .B2(n4930), .A(n4432), .ZN(n4925) );
  NAND2_X1 U5562 ( .A1(n8153), .A2(n4927), .ZN(n4923) );
  INV_X1 U5563 ( .A(n7844), .ZN(n8107) );
  NAND2_X1 U5564 ( .A1(n8148), .A2(n4807), .ZN(n8133) );
  AND2_X1 U5565 ( .A1(n8140), .A2(n8132), .ZN(n8128) );
  NOR2_X1 U5566 ( .A1(n4816), .A2(n8160), .ZN(n4815) );
  INV_X1 U5567 ( .A(n4818), .ZN(n4816) );
  NOR2_X1 U5568 ( .A1(n8154), .A2(n8302), .ZN(n8140) );
  OR2_X1 U5569 ( .A1(n8176), .A2(n8307), .ZN(n8154) );
  NOR2_X1 U5570 ( .A1(n8248), .A2(n4549), .ZN(n8204) );
  INV_X1 U5571 ( .A(n4940), .ZN(n4939) );
  OAI21_X1 U5572 ( .B1(n4941), .B2(n8236), .A(n4943), .ZN(n4940) );
  NAND2_X1 U5573 ( .A1(n4944), .A2(n8240), .ZN(n4943) );
  NOR2_X1 U5574 ( .A1(n8248), .A2(n8329), .ZN(n8217) );
  OR2_X1 U5575 ( .A1(n8246), .A2(n8333), .ZN(n8248) );
  AND2_X1 U5576 ( .A1(n4812), .A2(n4810), .ZN(n4809) );
  NAND2_X1 U5577 ( .A1(n4811), .A2(n4812), .ZN(n8237) );
  AND3_X1 U5578 ( .A1(n4394), .A2(n7215), .A3(n9700), .ZN(n7502) );
  NAND2_X1 U5579 ( .A1(n7419), .A2(n4637), .ZN(n7444) );
  AND2_X1 U5580 ( .A1(n7794), .A2(n7796), .ZN(n7906) );
  NAND2_X1 U5581 ( .A1(n7215), .A2(n4542), .ZN(n7425) );
  NAND2_X1 U5582 ( .A1(n7215), .A2(n10101), .ZN(n7308) );
  AND4_X1 U5583 ( .A1(n5262), .A2(n5261), .A3(n5260), .A4(n5259), .ZN(n9958)
         );
  AND2_X1 U5584 ( .A1(n7153), .A2(n10093), .ZN(n7215) );
  NOR2_X1 U5585 ( .A1(n9985), .A2(n7144), .ZN(n7153) );
  NAND2_X1 U5586 ( .A1(n7102), .A2(n7772), .ZN(n7147) );
  OR2_X1 U5587 ( .A1(n9983), .A2(n9982), .ZN(n9985) );
  AND4_X1 U5588 ( .A1(n5240), .A2(n5239), .A3(n5238), .A4(n5237), .ZN(n9996)
         );
  NAND2_X1 U5589 ( .A1(n4798), .A2(n4421), .ZN(n7736) );
  NAND2_X1 U5590 ( .A1(n4481), .A2(n7879), .ZN(n4798) );
  NAND2_X1 U5591 ( .A1(n4539), .A2(n6890), .ZN(n6950) );
  INV_X1 U5592 ( .A(n10023), .ZN(n4539) );
  NAND2_X1 U5593 ( .A1(n4540), .A2(n6756), .ZN(n10023) );
  INV_X1 U5594 ( .A(n9992), .ZN(n8241) );
  OR2_X1 U5595 ( .A1(n5734), .A2(n5735), .ZN(n9995) );
  INV_X1 U5596 ( .A(n10012), .ZN(n8226) );
  NOR2_X1 U5597 ( .A1(n6971), .A2(n7686), .ZN(n6973) );
  CLKBUF_X1 U5598 ( .A(n6766), .Z(n7752) );
  INV_X1 U5599 ( .A(n6765), .ZN(n7895) );
  OR2_X1 U5600 ( .A1(n6764), .A2(n7554), .ZN(n7746) );
  INV_X1 U5601 ( .A(n8271), .ZN(n4627) );
  NAND2_X1 U5602 ( .A1(n8272), .A2(n10024), .ZN(n4626) );
  OR2_X1 U5603 ( .A1(n8075), .A2(n8074), .ZN(n8076) );
  AND2_X1 U5604 ( .A1(n10050), .A2(n6761), .ZN(n10024) );
  INV_X1 U5605 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5678) );
  XNOR2_X1 U5606 ( .A(n5030), .B(P2_IR_REG_21__SCAN_IN), .ZN(n7921) );
  AND2_X1 U5607 ( .A1(n5375), .A2(n5347), .ZN(n7248) );
  INV_X1 U5608 ( .A(n5089), .ZN(n4910) );
  NAND2_X1 U5609 ( .A1(n5946), .A2(n4956), .ZN(n4587) );
  INV_X1 U5610 ( .A(n9396), .ZN(n9207) );
  INV_X1 U5611 ( .A(n6090), .ZN(n6089) );
  AND2_X1 U5612 ( .A1(n6229), .A2(n6228), .ZN(n6230) );
  NOR2_X1 U5613 ( .A1(n7222), .A2(n4960), .ZN(n4959) );
  INV_X1 U5614 ( .A(n4961), .ZN(n4960) );
  NAND2_X1 U5615 ( .A1(n5946), .A2(n4963), .ZN(n4962) );
  NOR2_X1 U5616 ( .A1(n8762), .A2(n4977), .ZN(n4976) );
  INV_X1 U5617 ( .A(n6156), .ZN(n4977) );
  INV_X1 U5618 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n6026) );
  NAND2_X1 U5619 ( .A1(n8793), .A2(n8796), .ZN(n4968) );
  NOR2_X1 U5620 ( .A1(n5910), .A2(n5905), .ZN(n6988) );
  AND2_X1 U5621 ( .A1(n5904), .A2(n5903), .ZN(n5905) );
  NAND2_X1 U5622 ( .A1(n8734), .A2(n8736), .ZN(n8735) );
  INV_X1 U5623 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n6064) );
  OR2_X1 U5624 ( .A1(n6065), .A2(n6064), .ZN(n6090) );
  NAND2_X1 U5625 ( .A1(n6047), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n6065) );
  INV_X1 U5626 ( .A(n6048), .ZN(n6047) );
  NAND2_X1 U5627 ( .A1(n6083), .A2(n6082), .ZN(n8794) );
  AND2_X1 U5628 ( .A1(n6334), .A2(n6333), .ZN(n9217) );
  AND2_X1 U5629 ( .A1(n6226), .A2(n6225), .ZN(n9214) );
  NOR2_X1 U5630 ( .A1(n5754), .A2(n6361), .ZN(n4745) );
  NAND2_X1 U5631 ( .A1(n6624), .A2(n6625), .ZN(n6623) );
  NAND2_X1 U5632 ( .A1(n9628), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n4638) );
  NOR2_X1 U5633 ( .A1(n6381), .A2(n4410), .ZN(n6576) );
  NAND2_X1 U5634 ( .A1(n6576), .A2(n6577), .ZN(n6575) );
  NOR2_X1 U5635 ( .A1(n4645), .A2(n4650), .ZN(n4644) );
  INV_X1 U5636 ( .A(n6593), .ZN(n4650) );
  INV_X1 U5637 ( .A(n4647), .ZN(n4645) );
  NOR2_X1 U5638 ( .A1(n9111), .A2(n4656), .ZN(n9126) );
  AND2_X1 U5639 ( .A1(n9115), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n4656) );
  NOR2_X1 U5640 ( .A1(n9126), .A2(n9125), .ZN(n9124) );
  INV_X1 U5641 ( .A(n7260), .ZN(n7259) );
  AND2_X1 U5642 ( .A1(n4642), .A2(n4641), .ZN(n9809) );
  NAND2_X1 U5643 ( .A1(n9175), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n4641) );
  OR2_X1 U5644 ( .A1(n9271), .A2(n9512), .ZN(n9262) );
  NOR2_X1 U5645 ( .A1(n9271), .A2(n4665), .ZN(n9219) );
  AND2_X1 U5646 ( .A1(n8699), .A2(n8698), .ZN(n9261) );
  INV_X1 U5647 ( .A(n9289), .ZN(n4737) );
  AND2_X1 U5648 ( .A1(n8876), .A2(n9216), .ZN(n9285) );
  NAND2_X1 U5649 ( .A1(n9373), .A2(n4393), .ZN(n9318) );
  NAND2_X1 U5650 ( .A1(n9238), .A2(n9004), .ZN(n9305) );
  AOI21_X1 U5651 ( .B1(n9348), .B2(n9235), .A(n9234), .ZN(n9335) );
  NAND2_X1 U5652 ( .A1(n9373), .A2(n4389), .ZN(n9327) );
  OR2_X1 U5653 ( .A1(n9539), .A2(n9358), .ZN(n9209) );
  AND2_X1 U5654 ( .A1(n9373), .A2(n4659), .ZN(n9342) );
  NAND2_X1 U5655 ( .A1(n6144), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n6159) );
  AND4_X1 U5656 ( .A1(n6179), .A2(n6178), .A3(n6177), .A4(n6176), .ZN(n9382)
         );
  NAND2_X1 U5657 ( .A1(n9394), .A2(n9395), .ZN(n9393) );
  OR2_X1 U5658 ( .A1(n9403), .A2(n9554), .ZN(n9387) );
  NAND2_X1 U5659 ( .A1(n6131), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n6146) );
  INV_X1 U5660 ( .A(n6133), .ZN(n6131) );
  AND4_X1 U5661 ( .A1(n6151), .A2(n6150), .A3(n6149), .A4(n6148), .ZN(n9421)
         );
  INV_X1 U5662 ( .A(n9453), .ZN(n9423) );
  AND2_X1 U5663 ( .A1(n9474), .A2(n4397), .ZN(n9429) );
  NAND2_X1 U5664 ( .A1(n9450), .A2(n9451), .ZN(n9449) );
  NAND2_X1 U5665 ( .A1(n9474), .A2(n4396), .ZN(n9444) );
  AND2_X1 U5666 ( .A1(n4752), .A2(n4443), .ZN(n4751) );
  NAND2_X1 U5667 ( .A1(n4755), .A2(n4753), .ZN(n4752) );
  INV_X1 U5668 ( .A(n7458), .ZN(n4753) );
  INV_X1 U5669 ( .A(n4755), .ZN(n4754) );
  NAND2_X1 U5670 ( .A1(n9474), .A2(n4758), .ZN(n9460) );
  NAND2_X1 U5671 ( .A1(n7461), .A2(n8826), .ZN(n7462) );
  AOI21_X1 U5672 ( .B1(n4706), .B2(n8847), .A(n8846), .ZN(n4705) );
  INV_X1 U5673 ( .A(n4708), .ZN(n4706) );
  AND2_X1 U5674 ( .A1(n9473), .A2(n9481), .ZN(n9474) );
  NOR2_X1 U5675 ( .A1(n7403), .A2(n9586), .ZN(n9473) );
  OR2_X1 U5676 ( .A1(n5971), .A2(n7331), .ZN(n5991) );
  NAND2_X1 U5677 ( .A1(n5989), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n6009) );
  INV_X1 U5678 ( .A(n5991), .ZN(n5989) );
  OR2_X1 U5679 ( .A1(n7363), .A2(n9589), .ZN(n7403) );
  AND4_X1 U5680 ( .A1(n6014), .A2(n6013), .A3(n6012), .A4(n6011), .ZN(n7402)
         );
  NAND2_X1 U5681 ( .A1(n4774), .A2(n4778), .ZN(n7400) );
  NAND2_X1 U5682 ( .A1(n7339), .A2(n4401), .ZN(n4774) );
  NAND2_X1 U5683 ( .A1(n7357), .A2(n8829), .ZN(n7408) );
  AND2_X1 U5684 ( .A1(n4661), .A2(n7069), .ZN(n7137) );
  NAND2_X1 U5685 ( .A1(n7069), .A2(n9863), .ZN(n7178) );
  NAND2_X1 U5686 ( .A1(n4739), .A2(n8887), .ZN(n7173) );
  NAND2_X1 U5687 ( .A1(n7050), .A2(n4743), .ZN(n4739) );
  NAND2_X1 U5688 ( .A1(n4603), .A2(n9014), .ZN(n7060) );
  INV_X1 U5689 ( .A(n7058), .ZN(n4603) );
  NAND2_X1 U5690 ( .A1(n6249), .A2(n6248), .ZN(n9521) );
  NAND2_X1 U5691 ( .A1(n6234), .A2(n6233), .ZN(n9524) );
  AND3_X1 U5692 ( .A1(n5901), .A2(n5900), .A3(n5899), .ZN(n9868) );
  AND3_X1 U5693 ( .A1(n5857), .A2(n5856), .A3(n5855), .ZN(n9855) );
  OR2_X1 U5694 ( .A1(n8995), .A2(n9080), .ZN(n9843) );
  AND2_X1 U5695 ( .A1(n6641), .A2(n9085), .ZN(n9892) );
  INV_X1 U5696 ( .A(n9883), .ZN(n9590) );
  OR2_X1 U5697 ( .A1(n6910), .A2(n9080), .ZN(n9883) );
  NAND2_X1 U5698 ( .A1(n6304), .A2(n6303), .ZN(n6907) );
  AND2_X1 U5699 ( .A1(n5779), .A2(n5781), .ZN(n4981) );
  XNOR2_X1 U5700 ( .A(n7869), .B(SI_30_), .ZN(n8810) );
  XNOR2_X1 U5701 ( .A(n7512), .B(n7511), .ZN(n8680) );
  NAND2_X1 U5702 ( .A1(n4797), .A2(n4715), .ZN(n4640) );
  NOR2_X1 U5703 ( .A1(n4400), .A2(P1_IR_REG_24__SCAN_IN), .ZN(n4715) );
  XNOR2_X1 U5704 ( .A(n5650), .B(n5649), .ZN(n7508) );
  XNOR2_X1 U5705 ( .A(n5608), .B(n5607), .ZN(n7431) );
  NAND2_X1 U5706 ( .A1(n4862), .A2(n5528), .ZN(n5544) );
  OR2_X1 U5707 ( .A1(n5767), .A2(n5766), .ZN(n5768) );
  NAND2_X1 U5708 ( .A1(n4581), .A2(n5764), .ZN(n4580) );
  INV_X1 U5709 ( .A(n5763), .ZN(n4581) );
  INV_X1 U5710 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5761) );
  OAI21_X1 U5711 ( .B1(n5343), .B2(n4398), .A(n4833), .ZN(n5420) );
  XNOR2_X1 U5712 ( .A(n5341), .B(n4993), .ZN(n6452) );
  NAND2_X1 U5713 ( .A1(n4690), .A2(n4856), .ZN(n5341) );
  NAND2_X1 U5714 ( .A1(n5269), .A2(n4694), .ZN(n4690) );
  NAND2_X1 U5715 ( .A1(n5271), .A2(n5270), .ZN(n5289) );
  AOI21_X1 U5716 ( .B1(n5180), .B2(n4671), .A(n4433), .ZN(n4670) );
  INV_X1 U5717 ( .A(n5166), .ZN(n4671) );
  NOR2_X1 U5718 ( .A1(n4672), .A2(n4669), .ZN(n4668) );
  INV_X1 U5719 ( .A(SI_3_), .ZN(n4674) );
  XNOR2_X1 U5720 ( .A(n5068), .B(n5020), .ZN(n5067) );
  NOR2_X1 U5721 ( .A1(n9683), .A2(n10172), .ZN(n9684) );
  NAND2_X1 U5722 ( .A1(n6795), .A2(n5173), .ZN(n6850) );
  AND2_X1 U5723 ( .A1(n4885), .A2(n5624), .ZN(n4884) );
  NAND2_X1 U5724 ( .A1(n4891), .A2(n5340), .ZN(n7475) );
  NAND2_X1 U5725 ( .A1(n5470), .A2(n5469), .ZN(n8318) );
  INV_X1 U5726 ( .A(n5715), .ZN(n4474) );
  NAND2_X1 U5727 ( .A1(n4896), .A2(n4402), .ZN(n7626) );
  NAND2_X1 U5728 ( .A1(n7618), .A2(n4900), .ZN(n4896) );
  AND4_X1 U5729 ( .A1(n5279), .A2(n5278), .A3(n5277), .A4(n5276), .ZN(n7324)
         );
  AND4_X1 U5730 ( .A1(n5336), .A2(n5335), .A3(n5334), .A4(n5333), .ZN(n7479)
         );
  AND4_X1 U5731 ( .A1(n5392), .A2(n5391), .A3(n5390), .A4(n5389), .ZN(n8242)
         );
  NAND2_X1 U5732 ( .A1(n7711), .A2(n5393), .ZN(n7643) );
  AND2_X1 U5733 ( .A1(n9943), .A2(n5127), .ZN(n6706) );
  NAND2_X1 U5734 ( .A1(n9943), .A2(n4905), .ZN(n6704) );
  NAND2_X1 U5735 ( .A1(n9942), .A2(n5123), .ZN(n9943) );
  INV_X1 U5736 ( .A(n6756), .ZN(n10025) );
  AND2_X1 U5737 ( .A1(n7119), .A2(n5222), .ZN(n4907) );
  AND2_X1 U5738 ( .A1(n6896), .A2(n5222), .ZN(n7118) );
  NAND2_X1 U5739 ( .A1(n7618), .A2(n5485), .ZN(n7669) );
  NAND2_X1 U5740 ( .A1(n5493), .A2(n5492), .ZN(n8314) );
  AND4_X1 U5741 ( .A1(n5309), .A2(n5308), .A3(n5307), .A4(n5306), .ZN(n9953)
         );
  OR2_X1 U5742 ( .A1(n7705), .A2(n9995), .ZN(n9954) );
  OR2_X1 U5743 ( .A1(n7705), .A2(n8241), .ZN(n9959) );
  NAND2_X1 U5744 ( .A1(n5731), .A2(n7941), .ZN(n7705) );
  INV_X1 U5745 ( .A(n6750), .ZN(n7686) );
  NAND2_X1 U5746 ( .A1(n5445), .A2(n5444), .ZN(n8324) );
  INV_X1 U5747 ( .A(n5151), .ZN(n4904) );
  AND2_X1 U5748 ( .A1(n5123), .A2(n5151), .ZN(n4902) );
  NAND2_X1 U5749 ( .A1(n4888), .A2(n7633), .ZN(n7700) );
  NAND2_X1 U5750 ( .A1(n7635), .A2(n7634), .ZN(n4888) );
  AND2_X1 U5751 ( .A1(n5637), .A2(n5616), .ZN(n8079) );
  NAND2_X1 U5752 ( .A1(n7938), .A2(n7939), .ZN(n4799) );
  INV_X1 U5753 ( .A(n7702), .ZN(n8113) );
  INV_X1 U5754 ( .A(P2_U3966), .ZN(n7967) );
  INV_X1 U5755 ( .A(n4500), .ZN(n9654) );
  INV_X1 U5756 ( .A(n4503), .ZN(n6504) );
  INV_X1 U5757 ( .A(n4496), .ZN(n6683) );
  AND2_X1 U5758 ( .A1(n5325), .A2(n5344), .ZN(n6866) );
  AND2_X1 U5759 ( .A1(n6488), .A2(n6487), .ZN(n9968) );
  OAI211_X1 U5760 ( .C1(n4534), .C2(n7886), .A(n4533), .B(n4531), .ZN(n8259)
         );
  AND2_X1 U5761 ( .A1(n7886), .A2(n4534), .ZN(n4532) );
  AOI222_X1 U5762 ( .A1(n7600), .A2(n10012), .B1(n8062), .B2(n9992), .C1(n7948), .C2(n8024), .ZN(n8268) );
  NAND2_X1 U5763 ( .A1(n4822), .A2(n4827), .ZN(n7931) );
  NAND2_X1 U5764 ( .A1(n8073), .A2(n4390), .ZN(n4822) );
  AND2_X1 U5765 ( .A1(n7581), .A2(n7580), .ZN(n7585) );
  XNOR2_X1 U5766 ( .A(n7582), .B(n7930), .ZN(n8269) );
  NAND2_X1 U5767 ( .A1(n4631), .A2(n4628), .ZN(n8270) );
  NOR2_X1 U5768 ( .A1(n4630), .A2(n4629), .ZN(n4628) );
  OR2_X1 U5769 ( .A1(n8040), .A2(n8226), .ZN(n4631) );
  NOR2_X1 U5770 ( .A1(n8041), .A2(n9995), .ZN(n4630) );
  NAND2_X1 U5771 ( .A1(n5614), .A2(n5613), .ZN(n8282) );
  NAND2_X1 U5772 ( .A1(n4924), .A2(n4927), .ZN(n8125) );
  NAND2_X1 U5773 ( .A1(n4926), .A2(n4931), .ZN(n8127) );
  OR2_X1 U5774 ( .A1(n4476), .A2(n4930), .ZN(n4924) );
  AND2_X1 U5775 ( .A1(n4933), .A2(n4408), .ZN(n8139) );
  NAND2_X1 U5776 ( .A1(n4476), .A2(n7573), .ZN(n4933) );
  NAND2_X1 U5777 ( .A1(n4817), .A2(n4818), .ZN(n8161) );
  AND2_X1 U5778 ( .A1(n5511), .A2(n5510), .ZN(n8159) );
  NAND2_X1 U5779 ( .A1(n8191), .A2(n7588), .ZN(n8171) );
  NOR2_X1 U5780 ( .A1(n8235), .A2(n4945), .ZN(n8215) );
  OR2_X1 U5781 ( .A1(n8235), .A2(n4941), .ZN(n8214) );
  NOR2_X1 U5782 ( .A1(n7503), .A2(n10102), .ZN(n8254) );
  NAND2_X1 U5783 ( .A1(n7495), .A2(n7798), .ZN(n7586) );
  NAND2_X1 U5784 ( .A1(n5378), .A2(n5377), .ZN(n7568) );
  NAND2_X1 U5785 ( .A1(n5300), .A2(n5299), .ZN(n7414) );
  NAND2_X1 U5786 ( .A1(n4528), .A2(n5255), .ZN(n9916) );
  NAND2_X1 U5787 ( .A1(n6427), .A2(n7879), .ZN(n4528) );
  NAND2_X1 U5788 ( .A1(n4480), .A2(n7145), .ZN(n7205) );
  CLKBUF_X1 U5789 ( .A(n9978), .Z(n9979) );
  NAND2_X1 U5790 ( .A1(n4917), .A2(n4921), .ZN(n7092) );
  NAND2_X1 U5791 ( .A1(n4922), .A2(n4482), .ZN(n4917) );
  INV_X1 U5792 ( .A(n7503), .ZN(n8222) );
  NAND2_X1 U5793 ( .A1(n10035), .A2(n6888), .ZN(n10001) );
  NAND2_X1 U5794 ( .A1(n6939), .A2(n4606), .ZN(n10059) );
  NAND2_X1 U5795 ( .A1(n7895), .A2(n5057), .ZN(n4606) );
  INV_X1 U5796 ( .A(n10049), .ZN(n7554) );
  NAND2_X1 U5797 ( .A1(n7943), .A2(n6884), .ZN(n10028) );
  NAND2_X1 U5798 ( .A1(n4632), .A2(n4624), .ZN(n8612) );
  NOR2_X1 U5799 ( .A1(n8270), .A2(n4625), .ZN(n4624) );
  NAND2_X1 U5800 ( .A1(n8037), .A2(n10114), .ZN(n4632) );
  NAND2_X1 U5801 ( .A1(n4627), .A2(n4626), .ZN(n4625) );
  AND2_X1 U5802 ( .A1(n6423), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10048) );
  INV_X1 U5803 ( .A(n10042), .ZN(n10045) );
  NAND2_X1 U5804 ( .A1(n5676), .A2(n5675), .ZN(n7456) );
  NAND2_X1 U5805 ( .A1(n5705), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5686) );
  INV_X1 U5806 ( .A(n5048), .ZN(n7725) );
  INV_X1 U5807 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7128) );
  INV_X1 U5808 ( .A(n7921), .ZN(n7932) );
  INV_X1 U5809 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n8578) );
  INV_X1 U5810 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n8340) );
  INV_X1 U5811 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n8587) );
  INV_X1 U5812 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6653) );
  INV_X1 U5813 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6458) );
  INV_X1 U5814 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6455) );
  INV_X1 U5815 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n8556) );
  INV_X1 U5816 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6439) );
  INV_X1 U5817 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n8552) );
  INV_X1 U5818 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6410) );
  OR2_X1 U5819 ( .A1(n5142), .A2(n5141), .ZN(n6503) );
  XNOR2_X1 U5820 ( .A(n5064), .B(P2_IR_REG_2__SCAN_IN), .ZN(n9658) );
  NAND2_X1 U5821 ( .A1(n4558), .A2(n6216), .ZN(n8663) );
  NAND2_X1 U5822 ( .A1(n6214), .A2(n8770), .ZN(n4558) );
  INV_X1 U5823 ( .A(n9333), .ZN(n9534) );
  AND2_X1 U5824 ( .A1(n4587), .A2(n4585), .ZN(n7389) );
  NAND2_X1 U5825 ( .A1(n4587), .A2(n4954), .ZN(n7330) );
  NAND2_X1 U5826 ( .A1(n4572), .A2(n4575), .ZN(n8674) );
  NAND2_X1 U5827 ( .A1(n4574), .A2(n4573), .ZN(n4572) );
  INV_X1 U5828 ( .A(n7539), .ZN(n4574) );
  OAI22_X1 U5829 ( .A1(n8752), .A2(n4427), .B1(n4388), .B2(n4392), .ZN(n8692)
         );
  NAND2_X1 U5830 ( .A1(n5946), .A2(n5945), .ZN(n7190) );
  NAND2_X1 U5831 ( .A1(n7539), .A2(n4570), .ZN(n4563) );
  NAND2_X1 U5832 ( .A1(n4968), .A2(n8794), .ZN(n7555) );
  AND3_X1 U5833 ( .A1(n6212), .A2(n6211), .A3(n6210), .ZN(n9212) );
  AND2_X1 U5834 ( .A1(n4552), .A2(n4559), .ZN(n8754) );
  AND2_X1 U5835 ( .A1(n6734), .A2(n6735), .ZN(n4950) );
  NAND2_X1 U5836 ( .A1(n4962), .A2(n4961), .ZN(n7221) );
  NAND2_X1 U5837 ( .A1(n4978), .A2(n6156), .ZN(n8761) );
  NAND2_X1 U5838 ( .A1(n6158), .A2(n6157), .ZN(n9551) );
  INV_X1 U5839 ( .A(n4585), .ZN(n4582) );
  OR2_X1 U5840 ( .A1(n7388), .A2(n7387), .ZN(n4980) );
  NAND2_X1 U5841 ( .A1(n6335), .A2(n9726), .ZN(n8786) );
  NAND2_X1 U5842 ( .A1(n6130), .A2(n6129), .ZN(n9561) );
  INV_X1 U5843 ( .A(n8786), .ZN(n8800) );
  AND2_X1 U5844 ( .A1(n6319), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8789) );
  OAI21_X1 U5845 ( .B1(n8752), .B2(n4971), .A(n4388), .ZN(n6286) );
  INV_X1 U5846 ( .A(n8806), .ZN(n8783) );
  OR3_X1 U5847 ( .A1(n6320), .A2(n9892), .A3(n6832), .ZN(n8806) );
  NAND2_X1 U5848 ( .A1(n6063), .A2(n6062), .ZN(n9574) );
  INV_X1 U5849 ( .A(n8792), .ZN(n8804) );
  NAND2_X1 U5850 ( .A1(n5789), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5790) );
  INV_X1 U5851 ( .A(n9288), .ZN(n9316) );
  INV_X1 U5852 ( .A(n9212), .ZN(n9349) );
  INV_X1 U5853 ( .A(n4948), .ZN(n5757) );
  AND3_X1 U5854 ( .A1(n5796), .A2(n5795), .A3(n5794), .ZN(n4996) );
  OR2_X1 U5855 ( .A1(n4386), .A2(n6682), .ZN(n5797) );
  OR2_X1 U5856 ( .A1(n6376), .A2(P1_U3084), .ZN(n9105) );
  OR2_X1 U5857 ( .A1(n6050), .A2(n5813), .ZN(n5814) );
  NAND2_X1 U5858 ( .A1(n6623), .A2(n6352), .ZN(n9626) );
  NAND2_X1 U5859 ( .A1(n4967), .A2(n5739), .ZN(n5853) );
  INV_X1 U5860 ( .A(n5782), .ZN(n4967) );
  OAI21_X1 U5861 ( .B1(n9748), .B2(n9749), .A(n4643), .ZN(n6382) );
  OR2_X1 U5862 ( .A1(n9746), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n4643) );
  NOR2_X1 U5863 ( .A1(n6382), .A2(n6383), .ZN(n6381) );
  AND2_X1 U5864 ( .A1(n9783), .A2(n9784), .ZN(n9785) );
  NAND2_X1 U5865 ( .A1(n6590), .A2(n6591), .ZN(n9783) );
  INV_X1 U5866 ( .A(n4642), .ZN(n9167) );
  AND2_X1 U5867 ( .A1(n9171), .A2(n9726), .ZN(n9815) );
  NOR2_X1 U5868 ( .A1(n9193), .A2(n4663), .ZN(n4662) );
  NAND2_X1 U5869 ( .A1(n4664), .A2(n9276), .ZN(n4663) );
  INV_X1 U5870 ( .A(n4665), .ZN(n4664) );
  NAND2_X1 U5871 ( .A1(n4787), .A2(n9218), .ZN(n4784) );
  OAI21_X1 U5872 ( .B1(n4785), .B2(n9218), .A(n4782), .ZN(n4781) );
  INV_X1 U5873 ( .A(n9514), .ZN(n9276) );
  INV_X1 U5874 ( .A(n9521), .ZN(n9295) );
  AND2_X1 U5875 ( .A1(n6326), .A2(n6251), .ZN(n9292) );
  NAND2_X1 U5876 ( .A1(n9364), .A2(n9363), .ZN(n9365) );
  AND2_X1 U5877 ( .A1(n6142), .A2(n6141), .ZN(n9392) );
  OAI21_X1 U5878 ( .B1(n9442), .B2(n4765), .A(n4762), .ZN(n9401) );
  NAND2_X1 U5879 ( .A1(n4761), .A2(n4766), .ZN(n9402) );
  NAND2_X1 U5880 ( .A1(n9442), .A2(n4767), .ZN(n4761) );
  AND2_X1 U5881 ( .A1(n4768), .A2(n4770), .ZN(n9428) );
  NAND2_X1 U5882 ( .A1(n9442), .A2(n9441), .ZN(n4768) );
  NAND2_X1 U5883 ( .A1(n9224), .A2(n9223), .ZN(n9465) );
  INV_X1 U5884 ( .A(n9574), .ZN(n9464) );
  AND2_X1 U5885 ( .A1(n4756), .A2(n4759), .ZN(n9198) );
  NAND2_X1 U5886 ( .A1(n9472), .A2(n7458), .ZN(n4756) );
  NAND2_X1 U5887 ( .A1(n7357), .A2(n4708), .ZN(n7460) );
  AND2_X1 U5888 ( .A1(n5970), .A2(n5969), .ZN(n7380) );
  OAI21_X1 U5889 ( .B1(n7339), .B2(n4405), .A(n7338), .ZN(n7352) );
  NAND2_X1 U5890 ( .A1(n4725), .A2(n4723), .ZN(n7341) );
  NAND2_X1 U5891 ( .A1(n4725), .A2(n8900), .ZN(n7233) );
  INV_X1 U5892 ( .A(n9868), .ZN(n7133) );
  INV_X1 U5893 ( .A(n9855), .ZN(n7074) );
  NAND2_X1 U5894 ( .A1(n9425), .A2(n7010), .ZN(n9495) );
  AND2_X1 U5895 ( .A1(n7009), .A2(n5830), .ZN(n7010) );
  INV_X1 U5896 ( .A(n9321), .ZN(n9356) );
  INV_X1 U5897 ( .A(n9480), .ZN(n9367) );
  AND2_X1 U5898 ( .A1(n9425), .A2(n6911), .ZN(n9493) );
  NOR2_X1 U5899 ( .A1(n9511), .A2(n4456), .ZN(n4602) );
  AND2_X1 U5900 ( .A1(n6292), .A2(n6291), .ZN(n9616) );
  AND2_X1 U5901 ( .A1(n6315), .A2(n6307), .ZN(n9841) );
  XNOR2_X1 U5902 ( .A(n7878), .B(n7877), .ZN(n9623) );
  NOR2_X1 U5903 ( .A1(n4716), .A2(n4713), .ZN(n5750) );
  NAND2_X1 U5904 ( .A1(n4797), .A2(n4710), .ZN(n4713) );
  INV_X1 U5905 ( .A(n6287), .ZN(n7298) );
  INV_X1 U5906 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n8411) );
  NAND2_X1 U5907 ( .A1(n4680), .A2(n5545), .ZN(n5554) );
  NAND2_X1 U5908 ( .A1(n4862), .A2(n4684), .ZN(n4680) );
  INV_X1 U5909 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7204) );
  INV_X1 U5910 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7116) );
  INV_X1 U5911 ( .A(n6309), .ZN(n9069) );
  INV_X1 U5912 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n6999) );
  XNOR2_X1 U5913 ( .A(n5770), .B(n5769), .ZN(n7000) );
  OAI21_X1 U5914 ( .B1(n6097), .B2(n4580), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5770) );
  INV_X1 U5915 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n6700) );
  INV_X1 U5916 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6655) );
  INV_X1 U5917 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n6457) );
  NAND2_X1 U5918 ( .A1(n5879), .A2(n4588), .ZN(n6022) );
  NOR2_X1 U5919 ( .A1(n4983), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n4588) );
  INV_X1 U5920 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6429) );
  INV_X1 U5921 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n8588) );
  INV_X1 U5922 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6419) );
  INV_X1 U5923 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6413) );
  XNOR2_X1 U5924 ( .A(n5181), .B(n5180), .ZN(n6409) );
  NAND2_X1 U5925 ( .A1(n4673), .A2(n5166), .ZN(n5181) );
  NAND2_X1 U5926 ( .A1(n5163), .A2(n5162), .ZN(n4673) );
  INV_X1 U5927 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n8574) );
  INV_X1 U5928 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6402) );
  INV_X1 U5929 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6400) );
  XNOR2_X1 U5930 ( .A(n4537), .B(n5135), .ZN(n6399) );
  NAND2_X1 U5931 ( .A1(n4538), .A2(n5111), .ZN(n4537) );
  NAND2_X1 U5932 ( .A1(n5109), .A2(n5108), .ZN(n4538) );
  NAND2_X1 U5933 ( .A1(n4435), .A2(n4651), .ZN(n6391) );
  NAND2_X1 U5934 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n4424), .ZN(n4651) );
  NOR2_X1 U5935 ( .A1(n10166), .A2(n10165), .ZN(n10164) );
  NOR2_X1 U5936 ( .A1(n10174), .A2(n10173), .ZN(n10172) );
  NOR2_X1 U5937 ( .A1(n9688), .A2(n10179), .ZN(n10160) );
  AOI21_X1 U5938 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10158), .ZN(n10157) );
  NOR2_X1 U5939 ( .A1(n10157), .A2(n10156), .ZN(n10155) );
  AOI21_X1 U5940 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10155), .ZN(n10154) );
  OAI21_X1 U5941 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10152), .ZN(n10150) );
  OAI21_X1 U5942 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n10146), .ZN(n10144) );
  AOI211_X1 U5943 ( .C1(n8289), .C2(n9957), .A(n7639), .B(n7638), .ZN(n7640)
         );
  AOI22_X1 U5944 ( .A1(n4529), .A2(n7940), .B1(n4799), .B2(n4800), .ZN(n7947)
         );
  INV_X1 U5945 ( .A(n4490), .ZN(n4489) );
  NAND2_X1 U5946 ( .A1(n4492), .A2(n8081), .ZN(n4491) );
  NAND2_X1 U5947 ( .A1(n4494), .A2(n8020), .ZN(n4493) );
  NAND2_X1 U5948 ( .A1(n4623), .A2(n4622), .ZN(P2_U3516) );
  NAND2_X1 U5949 ( .A1(n10115), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n4622) );
  NAND2_X1 U5950 ( .A1(n8612), .A2(n10117), .ZN(n4623) );
  INV_X1 U5951 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n9184) );
  NAND2_X1 U5952 ( .A1(n4601), .A2(n4600), .ZN(P1_U3551) );
  NAND2_X1 U5953 ( .A1(n9908), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n4600) );
  NAND2_X1 U5954 ( .A1(n9599), .A2(n9910), .ZN(n4601) );
  AND2_X1 U5955 ( .A1(n6265), .A2(n4969), .ZN(n4388) );
  NOR2_X1 U5956 ( .A1(n6916), .A2(n6344), .ZN(n5824) );
  INV_X1 U5957 ( .A(n8126), .ZN(n4928) );
  INV_X1 U5958 ( .A(n9199), .ZN(n4758) );
  INV_X1 U5959 ( .A(n6310), .ZN(n6308) );
  AND2_X1 U5960 ( .A1(n4659), .A2(n9333), .ZN(n4389) );
  AND2_X1 U5961 ( .A1(n4828), .A2(n7854), .ZN(n4390) );
  OR2_X1 U5962 ( .A1(n9097), .A2(n7351), .ZN(n4391) );
  OR2_X1 U5963 ( .A1(n6285), .A2(n6284), .ZN(n4392) );
  NAND2_X1 U5964 ( .A1(n5552), .A2(n5551), .ZN(n8297) );
  AND2_X1 U5965 ( .A1(n4389), .A2(n9312), .ZN(n4393) );
  NAND2_X1 U5966 ( .A1(n4910), .A2(n4997), .ZN(n5112) );
  INV_X1 U5967 ( .A(n9539), .ZN(n9346) );
  NAND2_X1 U5968 ( .A1(n6189), .A2(n6188), .ZN(n9539) );
  INV_X1 U5969 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5034) );
  AND2_X1 U5970 ( .A1(n4542), .A2(n4541), .ZN(n4394) );
  NAND2_X1 U5971 ( .A1(n7786), .A2(n7784), .ZN(n4395) );
  AND2_X1 U5972 ( .A1(n9570), .A2(n9467), .ZN(n9203) );
  INV_X1 U5973 ( .A(n9882), .ZN(n7229) );
  AND3_X1 U5974 ( .A1(n5943), .A2(n5942), .A3(n5941), .ZN(n9882) );
  INV_X1 U5975 ( .A(n9990), .ZN(n7094) );
  INV_X1 U5976 ( .A(n8042), .ZN(n4696) );
  AND2_X1 U5977 ( .A1(n4657), .A2(n9187), .ZN(n4396) );
  NAND2_X1 U5978 ( .A1(n8683), .A2(n8682), .ZN(n9512) );
  INV_X1 U5979 ( .A(n9512), .ZN(n4666) );
  NAND2_X1 U5980 ( .A1(n5634), .A2(n5633), .ZN(n8274) );
  AND2_X1 U5981 ( .A1(n4396), .A2(n9433), .ZN(n4397) );
  OR2_X1 U5982 ( .A1(n5395), .A2(n4835), .ZN(n4398) );
  NOR2_X1 U5983 ( .A1(n5089), .A2(n4911), .ZN(n5138) );
  INV_X1 U5984 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5036) );
  NAND2_X1 U5985 ( .A1(n5756), .A2(n7522), .ZN(n6007) );
  NAND2_X1 U5987 ( .A1(n9706), .A2(n7958), .ZN(n4399) );
  NAND2_X1 U5988 ( .A1(n5748), .A2(n5771), .ZN(n4400) );
  AOI21_X1 U5989 ( .B1(n8810), .B2(n7879), .A(n7867), .ZN(n8264) );
  AND2_X1 U5990 ( .A1(n4391), .A2(n7338), .ZN(n4401) );
  OR2_X1 U5991 ( .A1(n5506), .A2(n5505), .ZN(n4402) );
  NAND3_X1 U5992 ( .A1(n4872), .A2(n5026), .A3(n5031), .ZN(n4403) );
  AND2_X1 U5993 ( .A1(n4544), .A2(n8103), .ZN(n4404) );
  NOR2_X1 U5994 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5015) );
  AND2_X1 U5995 ( .A1(n9098), .A2(n9891), .ZN(n4405) );
  AND2_X1 U5996 ( .A1(n5137), .A2(SI_4_), .ZN(n4406) );
  NAND2_X1 U5997 ( .A1(n6045), .A2(n6044), .ZN(n9199) );
  INV_X2 U5998 ( .A(n8814), .ZN(n6050) );
  INV_X1 U5999 ( .A(n7779), .ZN(n4620) );
  NAND2_X1 U6000 ( .A1(n9276), .A2(n9289), .ZN(n4407) );
  NAND2_X1 U6001 ( .A1(n8307), .A2(n7950), .ZN(n4408) );
  AND2_X1 U6002 ( .A1(n8978), .A2(n9065), .ZN(n9218) );
  INV_X1 U6003 ( .A(n8236), .ZN(n4810) );
  AND2_X1 U6004 ( .A1(n5877), .A2(n5740), .ZN(n5879) );
  AND4_X1 U6005 ( .A1(n8929), .A2(n8996), .A3(n8917), .A4(n8920), .ZN(n4409)
         );
  AND2_X1 U6006 ( .A1(n6359), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n4410) );
  AND2_X1 U6007 ( .A1(n8016), .A2(n9971), .ZN(n4411) );
  NAND2_X1 U6008 ( .A1(n7881), .A2(n7880), .ZN(n8257) );
  NAND2_X1 U6009 ( .A1(n9481), .A2(n8842), .ZN(n4759) );
  OR2_X1 U6010 ( .A1(n7497), .A2(n7716), .ZN(n7798) );
  INV_X1 U6011 ( .A(n7798), .ZN(n4814) );
  AND2_X1 U6012 ( .A1(n8884), .A2(n8891), .ZN(n8888) );
  OR2_X1 U6013 ( .A1(n5920), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n4412) );
  AND2_X1 U6014 ( .A1(n4496), .A2(n4495), .ZN(n4413) );
  OR2_X1 U6015 ( .A1(n7814), .A2(n8224), .ZN(n4414) );
  INV_X1 U6016 ( .A(n5755), .ZN(n7522) );
  NAND2_X1 U6018 ( .A1(n5879), .A2(n5741), .ZN(n5920) );
  AND2_X1 U6019 ( .A1(n4639), .A2(n4638), .ZN(n4415) );
  NAND2_X1 U6020 ( .A1(n5659), .A2(n5658), .ZN(n8272) );
  AND2_X1 U6021 ( .A1(n9564), .A2(n9453), .ZN(n4416) );
  AND3_X1 U6022 ( .A1(n5883), .A2(n5882), .A3(n5881), .ZN(n9863) );
  AND2_X1 U6023 ( .A1(n8148), .A2(n7836), .ZN(n4417) );
  INV_X1 U6024 ( .A(n4857), .ZN(n4856) );
  OAI21_X1 U6025 ( .B1(n4860), .B2(n4858), .A(n5317), .ZN(n4857) );
  AND2_X1 U6026 ( .A1(n4978), .A2(n4976), .ZN(n4418) );
  AND2_X1 U6027 ( .A1(n4696), .A2(n5633), .ZN(n4419) );
  AND2_X1 U6028 ( .A1(n4513), .A2(n4517), .ZN(n4420) );
  AND2_X1 U6029 ( .A1(n5168), .A2(n5169), .ZN(n4421) );
  INV_X1 U6030 ( .A(n4957), .ZN(n4956) );
  OR2_X1 U6031 ( .A1(n5966), .A2(n4958), .ZN(n4957) );
  OR2_X1 U6032 ( .A1(n8272), .A2(n7606), .ZN(n7854) );
  INV_X1 U6033 ( .A(n9193), .ZN(n9503) );
  NAND2_X1 U6034 ( .A1(n8813), .A2(n8812), .ZN(n9193) );
  AND2_X1 U6035 ( .A1(n4734), .A2(n4602), .ZN(n4422) );
  AND2_X1 U6036 ( .A1(n4404), .A2(n4543), .ZN(n4423) );
  INV_X1 U6037 ( .A(n9368), .ZN(n9355) );
  NAND2_X1 U6038 ( .A1(n6172), .A2(n6171), .ZN(n9368) );
  INV_X1 U6039 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n4712) );
  NAND2_X1 U6040 ( .A1(n5836), .A2(n4746), .ZN(n9106) );
  AND2_X1 U6041 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n4424) );
  NOR2_X1 U6042 ( .A1(n9406), .A2(n9204), .ZN(n4425) );
  AND2_X1 U6043 ( .A1(n7401), .A2(n7411), .ZN(n4426) );
  OR2_X1 U6044 ( .A1(n4392), .A2(n4971), .ZN(n4427) );
  INV_X1 U6045 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n4984) );
  OR2_X1 U6046 ( .A1(n7824), .A2(n7825), .ZN(n4428) );
  OR2_X1 U6047 ( .A1(n6097), .A2(n5763), .ZN(n4429) );
  AND4_X1 U6048 ( .A1(n5007), .A2(n5006), .A3(n5005), .A4(n5004), .ZN(n4430)
         );
  NAND2_X1 U6049 ( .A1(n4871), .A2(n5015), .ZN(n5089) );
  NOR2_X1 U6050 ( .A1(n7401), .A2(n7411), .ZN(n4431) );
  NOR2_X1 U6051 ( .A1(n8132), .A2(n7840), .ZN(n4432) );
  NAND2_X1 U6052 ( .A1(n5798), .A2(n5738), .ZN(n5782) );
  AND2_X1 U6053 ( .A1(n5183), .A2(SI_6_), .ZN(n4433) );
  INV_X1 U6054 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6407) );
  INV_X1 U6055 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6397) );
  INV_X1 U6056 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n8436) );
  NOR2_X1 U6057 ( .A1(n4666), .A2(n9217), .ZN(n4434) );
  INV_X1 U6058 ( .A(n4787), .ZN(n4786) );
  AND2_X1 U6059 ( .A1(n9254), .A2(n4407), .ZN(n4787) );
  AND2_X1 U6060 ( .A1(n5837), .A2(n4652), .ZN(n4435) );
  AND2_X1 U6061 ( .A1(n9534), .A2(n9349), .ZN(n4436) );
  NAND2_X1 U6062 ( .A1(n4779), .A2(n9023), .ZN(n4437) );
  INV_X1 U6063 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5741) );
  OR2_X1 U6064 ( .A1(n9203), .A2(n4416), .ZN(n4438) );
  NAND2_X1 U6065 ( .A1(n8144), .A2(n4408), .ZN(n4439) );
  AND4_X1 U6066 ( .A1(n4999), .A2(n5000), .A3(n8363), .A4(n5345), .ZN(n4440)
         );
  AND2_X1 U6067 ( .A1(n4785), .A2(n9244), .ZN(n4441) );
  AND3_X1 U6068 ( .A1(n5745), .A2(n5744), .A3(n5746), .ZN(n4442) );
  INV_X1 U6069 ( .A(n9225), .ZN(n4729) );
  OR2_X1 U6070 ( .A1(n4758), .A2(n9200), .ZN(n4443) );
  NOR2_X1 U6071 ( .A1(n9993), .A2(n7093), .ZN(n4444) );
  AND2_X1 U6072 ( .A1(n7442), .A2(n4399), .ZN(n4445) );
  AND3_X1 U6073 ( .A1(n5786), .A2(n5785), .A3(n5784), .ZN(n6915) );
  NOR2_X1 U6074 ( .A1(n4845), .A2(n7887), .ZN(n4446) );
  AND2_X1 U6075 ( .A1(n4810), .A2(n7809), .ZN(n4447) );
  AND2_X1 U6076 ( .A1(n7802), .A2(n7443), .ZN(n7907) );
  AND2_X1 U6077 ( .A1(n7129), .A2(n4740), .ZN(n4448) );
  AND2_X1 U6078 ( .A1(n4981), .A2(n5751), .ZN(n4449) );
  AND2_X1 U6079 ( .A1(n4514), .A2(n4519), .ZN(n4450) );
  AND2_X1 U6080 ( .A1(n4395), .A2(n7145), .ZN(n4451) );
  INV_X1 U6081 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n4613) );
  INV_X1 U6082 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5739) );
  OR2_X1 U6083 ( .A1(n4716), .A2(n4714), .ZN(n4717) );
  OR2_X1 U6084 ( .A1(n9186), .A2(n9185), .ZN(P1_U3260) );
  INV_X1 U6085 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n4551) );
  NAND2_X1 U6086 ( .A1(n9202), .A2(n4988), .ZN(n9442) );
  INV_X1 U6087 ( .A(n9485), .ZN(n9200) );
  AND2_X1 U6088 ( .A1(n5789), .A2(n5768), .ZN(n6309) );
  INV_X1 U6089 ( .A(n7828), .ZN(n4519) );
  NAND2_X1 U6090 ( .A1(n9373), .A2(n9355), .ZN(n4453) );
  XNOR2_X1 U6091 ( .A(n5790), .B(P1_IR_REG_22__SCAN_IN), .ZN(n6310) );
  OAI21_X1 U6092 ( .B1(n7652), .B2(n7651), .A(n5436), .ZN(n7694) );
  NAND2_X1 U6093 ( .A1(n6099), .A2(n6098), .ZN(n9564) );
  INV_X1 U6094 ( .A(n8829), .ZN(n4709) );
  NAND2_X1 U6095 ( .A1(n8871), .A2(n8870), .ZN(n9507) );
  INV_X1 U6096 ( .A(n9507), .ZN(n4667) );
  OR2_X1 U6097 ( .A1(n5401), .A2(P2_IR_REG_16__SCAN_IN), .ZN(n4454) );
  INV_X1 U6098 ( .A(n7606), .ZN(n8062) );
  NOR3_X1 U6099 ( .A1(n8248), .A2(n8314), .A3(n4547), .ZN(n4545) );
  NOR2_X1 U6100 ( .A1(n7557), .A2(n6116), .ZN(n4455) );
  AND2_X1 U6101 ( .A1(n5644), .A2(n5643), .ZN(n8042) );
  INV_X1 U6102 ( .A(n9214), .ZN(n9336) );
  AND2_X1 U6103 ( .A1(n9512), .A2(n9892), .ZN(n4456) );
  NAND2_X1 U6104 ( .A1(n4563), .A2(n4567), .ZN(n8713) );
  INV_X1 U6105 ( .A(n4570), .ZN(n4569) );
  NOR2_X1 U6106 ( .A1(n4975), .A2(n4571), .ZN(n4570) );
  NAND2_X1 U6107 ( .A1(n9474), .A2(n4657), .ZN(n4658) );
  AND2_X1 U6108 ( .A1(n7419), .A2(n7794), .ZN(n4457) );
  INV_X1 U6109 ( .A(n6890), .ZN(n6933) );
  AND3_X1 U6110 ( .A1(n5145), .A2(n5144), .A3(n5143), .ZN(n6890) );
  NAND2_X1 U6111 ( .A1(n5557), .A2(n5556), .ZN(n8294) );
  INV_X1 U6112 ( .A(n4546), .ZN(n8185) );
  NOR2_X1 U6113 ( .A1(n8248), .A2(n4547), .ZN(n4546) );
  NAND2_X1 U6114 ( .A1(n6088), .A2(n6087), .ZN(n9570) );
  INV_X1 U6115 ( .A(n4576), .ZN(n4573) );
  AND2_X1 U6116 ( .A1(n7541), .A2(n7540), .ZN(n4576) );
  AND2_X1 U6117 ( .A1(n5522), .A2(n5521), .ZN(n4458) );
  NOR2_X1 U6118 ( .A1(n9574), .A2(n9452), .ZN(n4459) );
  INV_X1 U6119 ( .A(n9312), .ZN(n9530) );
  AND2_X1 U6120 ( .A1(n6218), .A2(n6217), .ZN(n9312) );
  INV_X1 U6121 ( .A(n4560), .ZN(n4559) );
  NOR2_X1 U6122 ( .A1(n6216), .A2(n8665), .ZN(n4560) );
  NOR2_X1 U6123 ( .A1(n5736), .A2(n5737), .ZN(n4460) );
  OR2_X1 U6124 ( .A1(n8181), .A2(n7951), .ZN(n4461) );
  AND2_X1 U6125 ( .A1(n4935), .A2(n4399), .ZN(n4462) );
  OR2_X1 U6126 ( .A1(n9312), .A2(n9214), .ZN(n4463) );
  AND2_X1 U6127 ( .A1(n4952), .A2(n4951), .ZN(n4464) );
  INV_X2 U6128 ( .A(n10115), .ZN(n10117) );
  AND2_X1 U6129 ( .A1(n4394), .A2(n7215), .ZN(n4465) );
  OR2_X1 U6130 ( .A1(n5946), .A2(n5945), .ZN(n4466) );
  AND2_X1 U6131 ( .A1(n4646), .A2(n4647), .ZN(n4467) );
  AND2_X1 U6132 ( .A1(n7781), .A2(n7779), .ZN(n7900) );
  OAI21_X1 U6133 ( .B1(n5946), .B2(n4582), .A(n4584), .ZN(n4583) );
  NAND3_X1 U6134 ( .A1(n5879), .A2(n4797), .A3(n4796), .ZN(n4468) );
  AND2_X1 U6135 ( .A1(n4962), .A2(n4959), .ZN(n4469) );
  INV_X1 U6136 ( .A(n9203), .ZN(n4770) );
  INV_X1 U6137 ( .A(n9784), .ZN(n4649) );
  AND2_X2 U6138 ( .A1(n6649), .A2(n6640), .ZN(n9910) );
  AND2_X1 U6139 ( .A1(n6832), .A2(n9087), .ZN(n9486) );
  AND2_X1 U6140 ( .A1(n9160), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n4470) );
  NAND2_X1 U6141 ( .A1(n5426), .A2(n5425), .ZN(n8329) );
  INV_X1 U6142 ( .A(n8329), .ZN(n4944) );
  AND2_X1 U6143 ( .A1(n9989), .A2(n10080), .ZN(n8331) );
  NAND2_X1 U6144 ( .A1(n5327), .A2(n5326), .ZN(n9706) );
  INV_X1 U6145 ( .A(n9706), .ZN(n4541) );
  NAND2_X1 U6146 ( .A1(n6973), .A2(n6773), .ZN(n10020) );
  INV_X1 U6147 ( .A(n10020), .ZN(n4540) );
  INV_X1 U6148 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n4966) );
  NAND2_X1 U6149 ( .A1(n9626), .A2(n9627), .ZN(n4639) );
  INV_X1 U6150 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4864) );
  INV_X1 U6151 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n4949) );
  NAND2_X1 U6152 ( .A1(n6766), .A2(n7751), .ZN(n6765) );
  NAND2_X1 U6153 ( .A1(n7208), .A2(n7903), .ZN(n7313) );
  NAND2_X1 U6154 ( .A1(n6935), .A2(n6934), .ZN(n6948) );
  NAND2_X1 U6155 ( .A1(n10017), .A2(n6757), .ZN(n6758) );
  NAND2_X1 U6156 ( .A1(n6752), .A2(n6751), .ZN(n6782) );
  NAND2_X1 U6157 ( .A1(n10015), .A2(n10014), .ZN(n10017) );
  AND2_X2 U6158 ( .A1(n7313), .A2(n7312), .ZN(n7315) );
  INV_X1 U6159 ( .A(n5042), .ZN(n4908) );
  BUF_X1 U6160 ( .A(n6747), .Z(n7966) );
  NAND2_X1 U6161 ( .A1(n6746), .A2(n6748), .ZN(n6766) );
  NAND2_X1 U6162 ( .A1(n7499), .A2(n7498), .ZN(n7570) );
  NAND2_X1 U6163 ( .A1(n8034), .A2(n7578), .ZN(n7582) );
  NAND2_X1 U6164 ( .A1(n8170), .A2(n8169), .ZN(n8168) );
  AOI21_X1 U6165 ( .B1(n7952), .B2(n8318), .A(n8184), .ZN(n7572) );
  INV_X1 U6166 ( .A(n4909), .ZN(n5046) );
  NAND2_X1 U6167 ( .A1(n8068), .A2(n7575), .ZN(n8053) );
  NAND3_X1 U6168 ( .A1(n5046), .A2(n5045), .A3(n5044), .ZN(n6747) );
  OAI22_X1 U6169 ( .A1(n5040), .A2(n5118), .B1(n5117), .B2(n6943), .ZN(n4909)
         );
  NAND2_X1 U6170 ( .A1(n8168), .A2(n4461), .ZN(n8153) );
  OR2_X1 U6171 ( .A1(n8938), .A2(n8995), .ZN(n4485) );
  MUX2_X2 U6172 ( .A(n8896), .B(n8895), .S(n8995), .Z(n8898) );
  MUX2_X2 U6173 ( .A(n9082), .B(n9081), .S(n9080), .Z(n9093) );
  NOR2_X1 U6174 ( .A1(n8967), .A2(n8966), .ZN(n8969) );
  MUX2_X2 U6175 ( .A(n8957), .B(n8956), .S(n8995), .Z(n8961) );
  MUX2_X1 U6176 ( .A(n9075), .B(n9074), .S(n9321), .Z(n9079) );
  NAND2_X2 U6177 ( .A1(n9046), .A2(n9012), .ZN(n7050) );
  INV_X1 U6178 ( .A(n5162), .ZN(n4669) );
  AOI21_X1 U6179 ( .B1(n8959), .B2(n8960), .A(n9234), .ZN(n8965) );
  NAND2_X1 U6180 ( .A1(n4876), .A2(n5082), .ZN(n4875) );
  NAND2_X1 U6181 ( .A1(n7473), .A2(n5364), .ZN(n5382) );
  NAND2_X1 U6182 ( .A1(n4881), .A2(n4884), .ZN(n7605) );
  INV_X1 U6183 ( .A(n5571), .ZN(n4477) );
  NAND2_X1 U6184 ( .A1(n5002), .A2(n4985), .ZN(n5401) );
  NAND2_X1 U6185 ( .A1(n9952), .A2(n9951), .ZN(n9950) );
  OAI21_X1 U6186 ( .B1(n5714), .B2(n4473), .A(n4460), .ZN(P2_U3222) );
  NAND2_X1 U6187 ( .A1(n4475), .A2(n4474), .ZN(n4473) );
  NAND2_X1 U6188 ( .A1(n5717), .A2(n5716), .ZN(n4475) );
  OAI21_X1 U6189 ( .B1(n4905), .B2(n4904), .A(n4903), .ZN(n6796) );
  AOI21_X2 U6190 ( .B1(n9326), .B2(n9213), .A(n4436), .ZN(n9311) );
  OR2_X1 U6191 ( .A1(n6162), .A2(n5833), .ZN(n5835) );
  NAND2_X1 U6192 ( .A1(n4594), .A2(n9256), .ZN(n4593) );
  NAND2_X1 U6193 ( .A1(n4597), .A2(n7039), .ZN(n7040) );
  NAND2_X2 U6194 ( .A1(n7163), .A2(n9021), .ZN(n7231) );
  NAND2_X2 U6195 ( .A1(n7231), .A2(n7230), .ZN(n7339) );
  NAND2_X1 U6196 ( .A1(n7013), .A2(n7012), .ZN(n7011) );
  NAND2_X1 U6197 ( .A1(n4773), .A2(n4772), .ZN(n7457) );
  NAND3_X1 U6198 ( .A1(n4866), .A2(n5230), .A3(n4865), .ZN(n5252) );
  NAND2_X1 U6199 ( .A1(n4621), .A2(n7815), .ZN(n8201) );
  AOI222_X2 U6200 ( .A1(n10012), .A2(n8064), .B1(n8063), .B2(n9992), .C1(n8062), .C2(n9935), .ZN(n8277) );
  NAND2_X1 U6201 ( .A1(n4802), .A2(n4803), .ZN(n8091) );
  NAND2_X1 U6202 ( .A1(n7207), .A2(n7206), .ZN(n7208) );
  NAND2_X1 U6203 ( .A1(n8070), .A2(n8069), .ZN(n8068) );
  MUX2_X1 U6204 ( .A(n8995), .B(n8994), .S(n9071), .Z(n9001) );
  OAI21_X1 U6205 ( .B1(n5224), .B2(n5223), .A(n5225), .ZN(n5245) );
  INV_X1 U6206 ( .A(n5180), .ZN(n4672) );
  NAND2_X1 U6207 ( .A1(n5271), .A2(n4860), .ZN(n4855) );
  NAND2_X1 U6208 ( .A1(n8936), .A2(n4487), .ZN(n4486) );
  NAND2_X1 U6209 ( .A1(n4486), .A2(n4484), .ZN(n8940) );
  NAND2_X1 U6210 ( .A1(n6782), .A2(n6784), .ZN(n6781) );
  NAND2_X1 U6211 ( .A1(n6781), .A2(n6755), .ZN(n10015) );
  INV_X1 U6212 ( .A(n4911), .ZN(n4865) );
  NAND2_X1 U6213 ( .A1(n7098), .A2(n7097), .ZN(n7146) );
  NAND2_X1 U6214 ( .A1(n7635), .A2(n4882), .ZN(n4881) );
  NAND2_X1 U6215 ( .A1(n5380), .A2(n5379), .ZN(n5383) );
  NAND2_X1 U6216 ( .A1(n4919), .A2(n4921), .ZN(n4918) );
  NAND2_X1 U6217 ( .A1(n5013), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n4863) );
  AND4_X2 U6218 ( .A1(n5002), .A2(n4430), .A3(n4946), .A4(n4985), .ZN(n5009)
         );
  OR2_X1 U6219 ( .A1(n5118), .A2(n6981), .ZN(n5075) );
  NAND2_X2 U6220 ( .A1(n7315), .A2(n7314), .ZN(n7416) );
  NAND2_X1 U6221 ( .A1(n4915), .A2(n4913), .ZN(n9980) );
  NAND2_X1 U6222 ( .A1(n8971), .A2(n9036), .ZN(n8974) );
  NAND3_X1 U6223 ( .A1(n4521), .A2(n4522), .A3(n5200), .ZN(n5224) );
  NAND2_X1 U6224 ( .A1(n4855), .A2(n5287), .ZN(n5316) );
  OR2_X1 U6225 ( .A1(n8847), .A2(n8846), .ZN(n8925) );
  MUX2_X1 U6226 ( .A(n8965), .B(n8964), .S(n8995), .Z(n8967) );
  AND2_X1 U6227 ( .A1(n4485), .A2(n9226), .ZN(n4484) );
  NAND2_X1 U6228 ( .A1(n4877), .A2(n4875), .ZN(n5107) );
  NAND2_X1 U6229 ( .A1(n5458), .A2(n5457), .ZN(n7621) );
  NAND3_X1 U6230 ( .A1(n4493), .A2(n4491), .A3(n4489), .ZN(P2_U3264) );
  MUX2_X1 U6231 ( .A(n6466), .B(P2_REG1_REG_2__SCAN_IN), .S(n9658), .Z(n9655)
         );
  NAND3_X1 U6232 ( .A1(n4508), .A2(n7843), .A3(n7844), .ZN(n4507) );
  NAND3_X1 U6233 ( .A1(n7839), .A2(n7838), .A3(n4928), .ZN(n4508) );
  NAND2_X1 U6234 ( .A1(n7810), .A2(n4450), .ZN(n4511) );
  NAND2_X1 U6235 ( .A1(n4511), .A2(n4509), .ZN(n7831) );
  NAND2_X1 U6236 ( .A1(n7810), .A2(n4518), .ZN(n4513) );
  NAND3_X1 U6237 ( .A1(n5163), .A2(n4668), .A3(n5196), .ZN(n4521) );
  NAND2_X1 U6238 ( .A1(n4523), .A2(n4670), .ZN(n5197) );
  NAND2_X1 U6239 ( .A1(n4668), .A2(n5163), .ZN(n4523) );
  INV_X1 U6240 ( .A(n4670), .ZN(n4524) );
  NAND3_X1 U6241 ( .A1(n5109), .A2(n5108), .A3(n5135), .ZN(n4852) );
  NAND3_X1 U6242 ( .A1(n4527), .A2(n4525), .A3(n7907), .ZN(n7803) );
  NAND3_X1 U6243 ( .A1(n7797), .A2(n7890), .A3(n7796), .ZN(n4527) );
  NAND2_X1 U6244 ( .A1(n4478), .A2(n6396), .ZN(n4676) );
  AND2_X1 U6245 ( .A1(n8055), .A2(n4536), .ZN(n8028) );
  NAND2_X1 U6246 ( .A1(n8055), .A2(n4532), .ZN(n4531) );
  NAND2_X1 U6247 ( .A1(n8055), .A2(n8049), .ZN(n8043) );
  NAND2_X1 U6248 ( .A1(n8055), .A2(n4534), .ZN(n8260) );
  OR2_X1 U6249 ( .A1(n8055), .A2(n7886), .ZN(n4533) );
  INV_X1 U6250 ( .A(n4545), .ZN(n8176) );
  NAND2_X1 U6251 ( .A1(n5067), .A2(n5066), .ZN(n5070) );
  OAI21_X1 U6252 ( .B1(n7875), .B2(n4551), .A(n4550), .ZN(n5066) );
  NAND2_X1 U6253 ( .A1(n7875), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n4550) );
  NAND3_X1 U6254 ( .A1(n6214), .A2(n8770), .A3(n4561), .ZN(n4552) );
  NAND3_X1 U6255 ( .A1(n6214), .A2(n8770), .A3(n4556), .ZN(n4555) );
  NAND3_X1 U6256 ( .A1(n6214), .A2(n8770), .A3(n6215), .ZN(n8662) );
  OAI21_X1 U6257 ( .B1(n7539), .B2(n4566), .A(n4564), .ZN(n8714) );
  INV_X1 U6258 ( .A(n4577), .ZN(n5765) );
  INV_X1 U6259 ( .A(n4583), .ZN(n8728) );
  NAND2_X1 U6260 ( .A1(n5824), .A2(n7033), .ZN(n5787) );
  NAND2_X1 U6261 ( .A1(n9311), .A2(n4463), .ZN(n4592) );
  NAND2_X1 U6262 ( .A1(n9211), .A2(n4986), .ZN(n9326) );
  AOI21_X2 U6263 ( .B1(n9386), .B2(n9206), .A(n4595), .ZN(n9372) );
  NAND2_X1 U6264 ( .A1(n7037), .A2(n7061), .ZN(n7180) );
  INV_X1 U6265 ( .A(n4597), .ZN(n7038) );
  INV_X1 U6266 ( .A(n8888), .ZN(n4599) );
  NAND2_X1 U6267 ( .A1(n9049), .A2(n8887), .ZN(n9014) );
  NAND3_X1 U6268 ( .A1(n4605), .A2(n4604), .A3(n5018), .ZN(n5820) );
  NAND3_X2 U6269 ( .A1(n4607), .A2(n5012), .A3(n4612), .ZN(n7599) );
  NAND3_X1 U6270 ( .A1(n4610), .A2(n4609), .A3(n4608), .ZN(n5732) );
  NAND2_X2 U6271 ( .A1(n5732), .A2(n7599), .ZN(n6462) );
  NAND2_X1 U6272 ( .A1(n7147), .A2(n4618), .ZN(n4614) );
  NAND2_X1 U6273 ( .A1(n4614), .A2(n4615), .ZN(n7211) );
  NOR2_X2 U6274 ( .A1(n4716), .A2(n4640), .ZN(n5780) );
  AND3_X2 U6275 ( .A1(n4965), .A2(n5739), .A3(n5798), .ZN(n5877) );
  NAND2_X1 U6276 ( .A1(n4646), .A2(n4644), .ZN(n7257) );
  MUX2_X1 U6277 ( .A(n6349), .B(P1_REG2_REG_1__SCAN_IN), .S(n6391), .Z(n6607)
         );
  INV_X1 U6278 ( .A(n4658), .ZN(n9443) );
  NAND3_X1 U6279 ( .A1(n4661), .A2(n9876), .A3(n7069), .ZN(n7166) );
  INV_X1 U6280 ( .A(n7166), .ZN(n4660) );
  NAND2_X1 U6281 ( .A1(n4660), .A2(n9882), .ZN(n7237) );
  NAND2_X1 U6282 ( .A1(n9290), .A2(n4662), .ZN(n9499) );
  NAND2_X1 U6283 ( .A1(n9290), .A2(n9276), .ZN(n9271) );
  NAND2_X1 U6284 ( .A1(n4862), .A2(n4681), .ZN(n4679) );
  NAND2_X1 U6285 ( .A1(n5247), .A2(n5246), .ZN(n5269) );
  NAND2_X1 U6286 ( .A1(n5247), .A2(n4688), .ZN(n4687) );
  NAND2_X1 U6287 ( .A1(n7080), .A2(n6835), .ZN(n7020) );
  AND2_X2 U6288 ( .A1(n6835), .A2(n8836), .ZN(n7082) );
  OR2_X1 U6289 ( .A1(n7357), .A2(n4707), .ZN(n4704) );
  NAND2_X1 U6290 ( .A1(n4704), .A2(n4705), .ZN(n9483) );
  NAND3_X1 U6291 ( .A1(n4794), .A2(n4796), .A3(n4797), .ZN(n5775) );
  NAND3_X1 U6292 ( .A1(n4720), .A2(n8914), .A3(n4718), .ZN(n7356) );
  NAND3_X1 U6293 ( .A1(n4722), .A2(n8909), .A3(n4719), .ZN(n4718) );
  INV_X1 U6294 ( .A(n4723), .ZN(n4719) );
  NAND3_X1 U6295 ( .A1(n4721), .A2(n8909), .A3(n4722), .ZN(n4720) );
  INV_X1 U6296 ( .A(n8841), .ZN(n4721) );
  NAND2_X1 U6297 ( .A1(n4723), .A2(n8897), .ZN(n4722) );
  AOI21_X1 U6298 ( .B1(n7461), .B2(n4730), .A(n4726), .ZN(n9450) );
  OR2_X2 U6299 ( .A1(n9513), .A2(n9894), .ZN(n4733) );
  OAI21_X1 U6300 ( .B1(n7050), .B2(n4742), .A(n4448), .ZN(n7131) );
  INV_X1 U6301 ( .A(n9106), .ZN(n6825) );
  NAND3_X1 U6302 ( .A1(n5754), .A2(n5756), .A3(P1_REG3_REG_1__SCAN_IN), .ZN(
        n4747) );
  OAI21_X2 U6303 ( .B1(n9335), .B2(n9237), .A(n9236), .ZN(n9315) );
  AOI21_X2 U6304 ( .B1(n9313), .B2(n9240), .A(n9239), .ZN(n9286) );
  NAND2_X1 U6305 ( .A1(n7131), .A2(n8833), .ZN(n8841) );
  OR2_X2 U6306 ( .A1(n8869), .A2(n4551), .ZN(n5841) );
  AOI211_X2 U6307 ( .C1(n9892), .C2(n9507), .A(n9506), .B(n9505), .ZN(n9508)
         );
  NAND2_X1 U6308 ( .A1(n9278), .A2(n9269), .ZN(n9258) );
  NAND2_X1 U6309 ( .A1(n6825), .A2(n6824), .ZN(n6835) );
  NAND3_X2 U6310 ( .A1(n5841), .A2(n5839), .A3(n5840), .ZN(n6824) );
  OAI21_X1 U6311 ( .B1(n9472), .B2(n4754), .A(n4751), .ZN(n9459) );
  NAND2_X1 U6312 ( .A1(n4750), .A2(n4749), .ZN(n9202) );
  NAND2_X1 U6313 ( .A1(n9472), .A2(n4751), .ZN(n4750) );
  NAND2_X1 U6314 ( .A1(n7339), .A2(n4775), .ZN(n4773) );
  OAI211_X1 U6315 ( .C1(n9270), .C2(n4784), .A(n4781), .B(n4780), .ZN(n9504)
         );
  NAND2_X1 U6316 ( .A1(n9270), .A2(n4441), .ZN(n4780) );
  XNOR2_X2 U6317 ( .A(n4791), .B(n5781), .ZN(n9723) );
  OR2_X2 U6318 ( .A1(n5780), .A2(n6084), .ZN(n4791) );
  OR2_X1 U6319 ( .A1(n8148), .A2(n4806), .ZN(n4802) );
  NAND2_X1 U6320 ( .A1(n4817), .A2(n4815), .ZN(n7590) );
  NAND2_X1 U6321 ( .A1(n5343), .A2(n4833), .ZN(n4832) );
  NAND2_X1 U6322 ( .A1(n5343), .A2(n5342), .ZN(n5370) );
  NAND2_X1 U6323 ( .A1(n7857), .A2(n4844), .ZN(n4840) );
  OAI21_X1 U6324 ( .B1(n7850), .B2(n4446), .A(n4839), .ZN(n4841) );
  NAND2_X1 U6325 ( .A1(n4849), .A2(n7890), .ZN(n4848) );
  MUX2_X1 U6326 ( .A(n6392), .B(n5063), .S(n7875), .Z(n5094) );
  XNOR2_X1 U6327 ( .A(n4873), .B(n4872), .ZN(n5047) );
  INV_X1 U6328 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n4872) );
  AOI21_X1 U6329 ( .B1(n5032), .B2(n5031), .A(n4613), .ZN(n4873) );
  INV_X1 U6330 ( .A(n7689), .ZN(n4876) );
  INV_X1 U6331 ( .A(n5062), .ZN(n4880) );
  OAI21_X1 U6332 ( .B1(n4876), .B2(n7527), .A(n4874), .ZN(n9928) );
  AOI21_X1 U6333 ( .B1(n7689), .B2(n4880), .A(n4879), .ZN(n4874) );
  NAND2_X1 U6334 ( .A1(n7527), .A2(n4878), .ZN(n4877) );
  INV_X1 U6335 ( .A(n5082), .ZN(n4879) );
  NAND2_X1 U6336 ( .A1(n7688), .A2(n7689), .ZN(n7687) );
  NAND2_X1 U6337 ( .A1(n7527), .A2(n5062), .ZN(n7688) );
  NAND2_X1 U6338 ( .A1(n6795), .A2(n4889), .ZN(n6851) );
  NAND2_X1 U6339 ( .A1(n4892), .A2(n5393), .ZN(n4893) );
  NAND2_X1 U6340 ( .A1(n5383), .A2(n7712), .ZN(n4892) );
  NAND2_X1 U6341 ( .A1(n4893), .A2(n7644), .ZN(n7642) );
  NAND2_X1 U6342 ( .A1(n9942), .A2(n4902), .ZN(n4903) );
  INV_X1 U6343 ( .A(n7526), .ZN(n5041) );
  NAND2_X1 U6344 ( .A1(n7146), .A2(n4451), .ZN(n7207) );
  AOI21_X1 U6345 ( .B1(n7099), .B2(n4914), .A(n4444), .ZN(n4913) );
  NAND2_X1 U6346 ( .A1(n6948), .A2(n4916), .ZN(n4915) );
  NAND2_X1 U6347 ( .A1(n4936), .A2(n4445), .ZN(n7499) );
  CLKBUF_X1 U6348 ( .A(n4936), .Z(n4935) );
  NAND2_X1 U6349 ( .A1(n7416), .A2(n7415), .ZN(n7417) );
  INV_X1 U6350 ( .A(n7415), .ZN(n4938) );
  INV_X2 U6351 ( .A(n6162), .ZN(n5868) );
  NAND3_X1 U6352 ( .A1(n4952), .A2(n4951), .A3(n4950), .ZN(n6733) );
  NAND2_X1 U6353 ( .A1(n6724), .A2(n4953), .ZN(n4952) );
  NAND3_X1 U6354 ( .A1(n6675), .A2(n4995), .A3(n6724), .ZN(n4951) );
  NAND3_X1 U6355 ( .A1(n4968), .A2(n8794), .A3(n4455), .ZN(n6124) );
  NAND2_X1 U6356 ( .A1(n8752), .A2(n6232), .ZN(n8734) );
  NAND2_X1 U6357 ( .A1(n5780), .A2(n4449), .ZN(n9620) );
  NAND2_X1 U6358 ( .A1(n5461), .A2(n5460), .ZN(n5464) );
  INV_X1 U6359 ( .A(n6940), .ZN(n5057) );
  INV_X1 U6360 ( .A(n5011), .ZN(n5012) );
  OR2_X1 U6361 ( .A1(n8282), .A2(n8063), .ZN(n7575) );
  NAND2_X1 U6362 ( .A1(n6796), .A2(n6797), .ZN(n6795) );
  NAND4_X2 U6363 ( .A1(n5817), .A2(n5816), .A3(n5815), .A4(n5814), .ZN(n6440)
         );
  OR3_X1 U6364 ( .A1(n5048), .A2(n7923), .A3(n8020), .ZN(n10080) );
  OR2_X1 U6365 ( .A1(n10102), .A2(n8020), .ZN(n6883) );
  NAND2_X1 U6366 ( .A1(n7939), .A2(n7924), .ZN(n10012) );
  OR2_X1 U6367 ( .A1(n8289), .A2(n8113), .ZN(n7574) );
  NAND2_X1 U6368 ( .A1(n9341), .A2(n9209), .ZN(n9211) );
  INV_X1 U6369 ( .A(n6200), .ZN(n6203) );
  INV_X1 U6370 ( .A(n5047), .ZN(n7536) );
  XNOR2_X1 U6371 ( .A(n5792), .B(n5830), .ZN(n5861) );
  INV_X1 U6372 ( .A(n5523), .ZN(n5525) );
  OAI22_X1 U6373 ( .A1(n7885), .A2(n7884), .B1(n7917), .B2(n7887), .ZN(n7889)
         );
  AND2_X1 U6374 ( .A1(n4440), .A2(n4989), .ZN(n4985) );
  OR2_X1 U6375 ( .A1(n9346), .A2(n9210), .ZN(n4986) );
  OR2_X1 U6376 ( .A1(n9355), .A2(n9382), .ZN(n4987) );
  OR2_X1 U6377 ( .A1(n9464), .A2(n9201), .ZN(n4988) );
  AND2_X1 U6378 ( .A1(n5296), .A2(n5001), .ZN(n4989) );
  AND2_X1 U6379 ( .A1(n5246), .A2(n5229), .ZN(n4992) );
  AND2_X1 U6380 ( .A1(n5342), .A2(n5322), .ZN(n4993) );
  AND2_X1 U6381 ( .A1(n5270), .A2(n5251), .ZN(n4994) );
  INV_X1 U6382 ( .A(n9570), .ZN(n9187) );
  INV_X1 U6383 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5764) );
  AND2_X1 U6384 ( .A1(n6725), .A2(n5812), .ZN(n4995) );
  INV_X2 U6385 ( .A(n8208), .ZN(n10035) );
  OR2_X1 U6386 ( .A1(n6778), .A2(n6880), .ZN(n10131) );
  INV_X1 U6387 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5001) );
  INV_X1 U6388 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n8363) );
  INV_X1 U6389 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5748) );
  NAND2_X1 U6390 ( .A1(n6677), .A2(n5845), .ZN(n5788) );
  INV_X1 U6391 ( .A(n5865), .ZN(n5866) );
  INV_X1 U6392 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n5318) );
  INV_X1 U6393 ( .A(n5409), .ZN(n5407) );
  INV_X1 U6394 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n8438) );
  INV_X1 U6395 ( .A(n9937), .ZN(n6753) );
  INV_X1 U6396 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5008) );
  NAND2_X1 U6397 ( .A1(n5864), .A2(n5866), .ZN(n5867) );
  INV_X1 U6398 ( .A(n6192), .ZN(n6190) );
  OR2_X1 U6399 ( .A1(n6220), .A2(n6219), .ZN(n6237) );
  INV_X1 U6400 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5947) );
  INV_X1 U6401 ( .A(SI_25_), .ZN(n8456) );
  INV_X1 U6402 ( .A(SI_22_), .ZN(n8457) );
  INV_X1 U6403 ( .A(SI_13_), .ZN(n5319) );
  INV_X1 U6404 ( .A(n7476), .ZN(n5363) );
  INV_X1 U6405 ( .A(n9927), .ZN(n5106) );
  INV_X1 U6406 ( .A(n7620), .ZN(n5483) );
  XNOR2_X1 U6407 ( .A(n10055), .B(n5669), .ZN(n5059) );
  NAND2_X1 U6408 ( .A1(n5407), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5427) );
  NAND2_X1 U6409 ( .A1(n5494), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5513) );
  OR2_X1 U6410 ( .A1(n5091), .A2(n5063), .ZN(n5073) );
  OR2_X1 U6411 ( .A1(n5572), .A2(n7612), .ZN(n5574) );
  NAND2_X1 U6412 ( .A1(n5446), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5472) );
  NAND2_X1 U6413 ( .A1(n6462), .A2(n7515), .ZN(n5091) );
  OR2_X1 U6414 ( .A1(n5427), .A2(n8406), .ZN(n5448) );
  OR2_X1 U6415 ( .A1(n5386), .A2(n5385), .ZN(n5409) );
  INV_X1 U6416 ( .A(n7900), .ZN(n7097) );
  NAND2_X1 U6417 ( .A1(n6926), .A2(n7741), .ZN(n6956) );
  OR2_X2 U6418 ( .A1(n7965), .A2(n6750), .ZN(n7753) );
  INV_X1 U6419 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5702) );
  AND2_X1 U6420 ( .A1(n6988), .A2(n4991), .ZN(n5908) );
  XNOR2_X1 U6421 ( .A(n5861), .B(n5862), .ZN(n6724) );
  NAND2_X1 U6422 ( .A1(n6089), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n6102) );
  INV_X1 U6423 ( .A(n6201), .ZN(n6202) );
  NAND2_X1 U6424 ( .A1(n6190), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n6208) );
  OR2_X1 U6425 ( .A1(n6027), .A2(n6026), .ZN(n6048) );
  OR2_X1 U6426 ( .A1(n6159), .A2(n8763), .ZN(n6174) );
  OR2_X1 U6427 ( .A1(n5948), .A2(n5947), .ZN(n5971) );
  INV_X1 U6428 ( .A(n9863), .ZN(n7184) );
  AND2_X1 U6429 ( .A1(n8901), .A2(n9050), .ZN(n9018) );
  INV_X1 U6430 ( .A(n7069), .ZN(n7177) );
  OR2_X1 U6431 ( .A1(n7872), .A2(n7871), .ZN(n7873) );
  INV_X1 U6432 ( .A(n6849), .ZN(n5194) );
  INV_X1 U6433 ( .A(n7938), .ZN(n5668) );
  AND2_X1 U6434 ( .A1(n7548), .A2(n5058), .ZN(n7528) );
  OR2_X1 U6435 ( .A1(n8056), .A2(n5639), .ZN(n5644) );
  INV_X1 U6436 ( .A(n6430), .ZN(n7594) );
  INV_X1 U6437 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n6899) );
  INV_X1 U6438 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n8562) );
  INV_X1 U6439 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8406) );
  INV_X1 U6440 ( .A(n7953), .ZN(n8229) );
  AND2_X1 U6441 ( .A1(n5048), .A2(n7921), .ZN(n6762) );
  INV_X1 U6442 ( .A(n10102), .ZN(n10022) );
  INV_X1 U6443 ( .A(n7456), .ZN(n5690) );
  INV_X1 U6444 ( .A(n8789), .ZN(n8802) );
  INV_X1 U6445 ( .A(n7009), .ZN(n9088) );
  OR2_X1 U6446 ( .A1(n6250), .A2(n8785), .ZN(n6326) );
  INV_X1 U6447 ( .A(n6254), .ZN(n8694) );
  INV_X1 U6448 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n7331) );
  OR2_X1 U6449 ( .A1(n9521), .A2(n9306), .ZN(n9216) );
  OR2_X1 U6450 ( .A1(n6174), .A2(n6173), .ZN(n6192) );
  AND2_X1 U6451 ( .A1(n9009), .A2(n9230), .ZN(n9395) );
  NOR2_X1 U6452 ( .A1(n7237), .A2(n9891), .ZN(n7343) );
  INV_X1 U6453 ( .A(n9726), .ZN(n9087) );
  INV_X1 U6454 ( .A(n9486), .ZN(n9424) );
  AND2_X1 U6455 ( .A1(n6838), .A2(n6837), .ZN(n9420) );
  NAND2_X1 U6456 ( .A1(n7874), .A2(n7873), .ZN(n7878) );
  AND2_X1 U6457 ( .A1(n7513), .A2(n5657), .ZN(n7511) );
  INV_X1 U6458 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n6305) );
  AND2_X1 U6459 ( .A1(n5509), .A2(n5491), .ZN(n5508) );
  OR2_X1 U6460 ( .A1(n5256), .A2(n8562), .ZN(n5304) );
  AND2_X1 U6461 ( .A1(n5731), .A2(n5710), .ZN(n9949) );
  AND2_X1 U6462 ( .A1(n5667), .A2(n5666), .ZN(n7606) );
  AND4_X1 U6463 ( .A1(n5433), .A2(n5432), .A3(n5431), .A4(n5430), .ZN(n8240)
         );
  INV_X1 U6464 ( .A(n9972), .ZN(n9967) );
  INV_X2 U6465 ( .A(n5065), .ZN(n7879) );
  INV_X1 U6466 ( .A(n8232), .ZN(n7500) );
  NAND2_X1 U6467 ( .A1(n5701), .A2(n5700), .ZN(n6880) );
  INV_X1 U6468 ( .A(n10024), .ZN(n10110) );
  INV_X1 U6469 ( .A(n8331), .ZN(n10114) );
  INV_X1 U6470 ( .A(n6880), .ZN(n6777) );
  OAI21_X1 U6471 ( .B1(n9276), .B2(n8792), .A(n6338), .ZN(n6339) );
  INV_X1 U6472 ( .A(n8798), .ZN(n8774) );
  INV_X1 U6473 ( .A(n7000), .ZN(n9080) );
  AND2_X1 U6474 ( .A1(n6244), .A2(n6243), .ZN(n9288) );
  AND4_X1 U6475 ( .A1(n6138), .A2(n6137), .A3(n6136), .A4(n6135), .ZN(n9204)
         );
  INV_X1 U6476 ( .A(n9819), .ZN(n9765) );
  OR2_X1 U6477 ( .A1(n6375), .A2(n9726), .ZN(n9819) );
  INV_X1 U6478 ( .A(n9828), .ZN(n9778) );
  NAND2_X1 U6479 ( .A1(n9365), .A2(n4987), .ZN(n9341) );
  INV_X1 U6480 ( .A(n9031), .ZN(n9434) );
  INV_X1 U6481 ( .A(n9420), .ZN(n9489) );
  INV_X1 U6482 ( .A(n9850), .ZN(n7018) );
  NOR2_X1 U6483 ( .A1(n8710), .A2(n6639), .ZN(n6640) );
  INV_X1 U6484 ( .A(n9887), .ZN(n9894) );
  NAND2_X1 U6485 ( .A1(n7340), .A2(n9843), .ZN(n9887) );
  AND2_X1 U6486 ( .A1(n6638), .A2(n6907), .ZN(n6649) );
  OAI211_X1 U6487 ( .C1(P1_B_REG_SCAN_IN), .C2(n7298), .A(n6290), .B(n6289), 
        .ZN(n9829) );
  INV_X1 U6488 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5769) );
  INV_X1 U6489 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n9678) );
  OAI21_X1 U6490 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10137), .ZN(n10176) );
  INV_X1 U6491 ( .A(n8022), .ZN(n9969) );
  AND4_X1 U6492 ( .A1(n9963), .A2(n9962), .A3(n9961), .A4(n9960), .ZN(n9964)
         );
  INV_X1 U6493 ( .A(n9957), .ZN(n7723) );
  NAND2_X1 U6494 ( .A1(n6460), .A2(n10048), .ZN(n7963) );
  NAND2_X1 U6495 ( .A1(n6472), .A2(n7599), .ZN(n9972) );
  AND2_X1 U6496 ( .A1(n6426), .A2(n6425), .ZN(n8022) );
  OR2_X1 U6497 ( .A1(n8235), .A2(n8234), .ZN(n8336) );
  NAND2_X1 U6498 ( .A1(n10035), .A2(n10018), .ZN(n8232) );
  OR2_X1 U6499 ( .A1(n6778), .A2(n6777), .ZN(n10115) );
  NOR2_X1 U6500 ( .A1(n10037), .A2(n10036), .ZN(n10042) );
  AND2_X1 U6501 ( .A1(n7301), .A2(n7456), .ZN(n10044) );
  XNOR2_X1 U6502 ( .A(n5686), .B(n5685), .ZN(n7301) );
  INV_X1 U6503 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n8594) );
  INV_X1 U6504 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6422) );
  OR4_X1 U6505 ( .A1(n8692), .A2(n8704), .A3(n8705), .A4(n8806), .ZN(n8709) );
  INV_X1 U6506 ( .A(n9524), .ZN(n9302) );
  NAND2_X1 U6507 ( .A1(n8712), .A2(n6314), .ZN(n8792) );
  INV_X1 U6508 ( .A(n9217), .ZN(n9279) );
  INV_X1 U6509 ( .A(n9204), .ZN(n9436) );
  INV_X1 U6510 ( .A(n7402), .ZN(n9487) );
  INV_X1 U6511 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n9682) );
  OR2_X1 U6512 ( .A1(P1_U3083), .A2(n6635), .ZN(n9828) );
  NAND2_X1 U6513 ( .A1(n9425), .A2(n6912), .ZN(n9480) );
  INV_X1 U6514 ( .A(n9425), .ZN(n9490) );
  INV_X1 U6515 ( .A(n9910), .ZN(n9908) );
  OR2_X1 U6516 ( .A1(n9595), .A2(n9594), .ZN(n9615) );
  INV_X1 U6517 ( .A(n9900), .ZN(n9898) );
  AND2_X2 U6518 ( .A1(n6908), .A2(n6649), .ZN(n9900) );
  AND2_X1 U6519 ( .A1(n9841), .A2(n9829), .ZN(n9837) );
  INV_X1 U6520 ( .A(n9837), .ZN(n9838) );
  INV_X1 U6521 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n8681) );
  INV_X1 U6522 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7276) );
  INV_X1 U6523 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n6878) );
  INV_X1 U6524 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6444) );
  INV_X1 U6525 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6415) );
  INV_X1 U6526 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n10171) );
  NOR2_X1 U6527 ( .A1(n10160), .A2(n10159), .ZN(n10158) );
  OAI21_X1 U6528 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10149), .ZN(n10147) );
  INV_X1 U6529 ( .A(n7963), .ZN(P2_U3966) );
  INV_X1 U6530 ( .A(n9105), .ZN(P1_U4006) );
  NOR2_X1 U6531 ( .A1(P2_IR_REG_26__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n5006) );
  NOR2_X1 U6532 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n5005) );
  NOR2_X1 U6533 ( .A1(P2_IR_REG_23__SCAN_IN), .A2(P2_IR_REG_25__SCAN_IN), .ZN(
        n5004) );
  AND2_X2 U6534 ( .A1(n5009), .A2(n5008), .ZN(n5035) );
  INV_X1 U6535 ( .A(n5009), .ZN(n5675) );
  NAND2_X1 U6536 ( .A1(n5675), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5010) );
  INV_X1 U6537 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n8590) );
  OR2_X1 U6538 ( .A1(n5091), .A2(n8590), .ZN(n5023) );
  NAND2_X1 U6539 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5014) );
  MUX2_X1 U6540 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5014), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n5017) );
  INV_X1 U6541 ( .A(n5015), .ZN(n5016) );
  NAND2_X1 U6542 ( .A1(n5017), .A2(n5016), .ZN(n6482) );
  INV_X1 U6543 ( .A(n6482), .ZN(n9647) );
  NAND2_X1 U6544 ( .A1(n5088), .A2(n9647), .ZN(n5022) );
  NAND2_X1 U6545 ( .A1(n6462), .A2(n4478), .ZN(n5065) );
  AND2_X1 U6546 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5018) );
  NAND3_X1 U6547 ( .A1(n7875), .A2(SI_0_), .A3(P1_DATAO_REG_0__SCAN_IN), .ZN(
        n5019) );
  NAND2_X1 U6548 ( .A1(n5820), .A2(n5019), .ZN(n5068) );
  INV_X1 U6549 ( .A(SI_1_), .ZN(n5020) );
  XNOR2_X1 U6550 ( .A(n5067), .B(n5066), .ZN(n6406) );
  OR2_X1 U6551 ( .A1(n5065), .A2(n6406), .ZN(n5021) );
  INV_X2 U6552 ( .A(n6748), .ZN(n10055) );
  NOR2_X2 U6553 ( .A1(n5025), .A2(n4403), .ZN(n5028) );
  NAND2_X1 U6554 ( .A1(n5443), .A2(n5026), .ZN(n5027) );
  XNOR2_X2 U6555 ( .A(n5032), .B(n5031), .ZN(n8020) );
  NAND2_X1 U6556 ( .A1(n5048), .A2(n8020), .ZN(n6760) );
  INV_X1 U6557 ( .A(n5028), .ZN(n5029) );
  NAND2_X1 U6558 ( .A1(n5029), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5030) );
  NAND2_X4 U6559 ( .A1(n5033), .A2(n7939), .ZN(n5669) );
  NAND2_X1 U6560 ( .A1(n5038), .A2(n5036), .ZN(n8625) );
  INV_X1 U6561 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n8626) );
  XNOR2_X2 U6562 ( .A(n5037), .B(n8626), .ZN(n5042) );
  INV_X1 U6564 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n6943) );
  INV_X1 U6565 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n5040) );
  INV_X1 U6566 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n5043) );
  OR2_X1 U6567 ( .A1(n5129), .A2(n5043), .ZN(n5044) );
  OR2_X2 U6568 ( .A1(n6761), .A2(n7925), .ZN(n7938) );
  NAND2_X1 U6569 ( .A1(n7966), .A2(n7938), .ZN(n5060) );
  XNOR2_X1 U6570 ( .A(n5059), .B(n5060), .ZN(n7529) );
  NAND2_X1 U6571 ( .A1(n5152), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5055) );
  INV_X1 U6572 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n5049) );
  OR2_X1 U6573 ( .A1(n5117), .A2(n5049), .ZN(n5054) );
  INV_X1 U6574 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n5050) );
  OR2_X1 U6575 ( .A1(n5129), .A2(n5050), .ZN(n5053) );
  INV_X1 U6576 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n5051) );
  NAND4_X1 U6577 ( .A1(n5055), .A2(n5054), .A3(n5053), .A4(n5052), .ZN(n6764)
         );
  NAND2_X1 U6578 ( .A1(n4478), .A2(SI_0_), .ZN(n5056) );
  XNOR2_X1 U6579 ( .A(n5056), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n8637) );
  MUX2_X1 U6580 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8637), .S(n6462), .Z(n10049)
         );
  NAND2_X1 U6581 ( .A1(n6764), .A2(n10049), .ZN(n6940) );
  NAND2_X1 U6582 ( .A1(n5057), .A2(n7938), .ZN(n7548) );
  NAND2_X1 U6583 ( .A1(n7554), .A2(n5669), .ZN(n5058) );
  INV_X1 U6584 ( .A(n5059), .ZN(n5061) );
  NAND2_X1 U6585 ( .A1(n5061), .A2(n5060), .ZN(n5062) );
  INV_X1 U6586 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n5063) );
  OR2_X1 U6587 ( .A1(n5015), .A2(n4613), .ZN(n5064) );
  NAND2_X1 U6588 ( .A1(n5088), .A2(n9658), .ZN(n5072) );
  NAND2_X1 U6589 ( .A1(n5068), .A2(SI_1_), .ZN(n5069) );
  NAND2_X1 U6590 ( .A1(n5070), .A2(n5069), .ZN(n5093) );
  INV_X1 U6591 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6392) );
  XNOR2_X1 U6592 ( .A(n5094), .B(SI_2_), .ZN(n5092) );
  XNOR2_X1 U6593 ( .A(n5093), .B(n5092), .ZN(n6405) );
  OR2_X1 U6594 ( .A1(n5065), .A2(n6405), .ZN(n5071) );
  NAND2_X1 U6595 ( .A1(n5152), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5078) );
  NAND2_X1 U6596 ( .A1(n5725), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5077) );
  INV_X1 U6597 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n5074) );
  OR2_X1 U6598 ( .A1(n5117), .A2(n5074), .ZN(n5076) );
  INV_X1 U6599 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6981) );
  NAND2_X1 U6600 ( .A1(n7965), .A2(n7938), .ZN(n5080) );
  INV_X1 U6601 ( .A(n5079), .ZN(n5081) );
  NAND2_X1 U6602 ( .A1(n5081), .A2(n5080), .ZN(n5082) );
  NAND2_X1 U6603 ( .A1(n5152), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5087) );
  OR2_X1 U6604 ( .A1(n5117), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5086) );
  INV_X1 U6605 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n5083) );
  OR2_X1 U6606 ( .A1(n5129), .A2(n5083), .ZN(n5085) );
  INV_X1 U6607 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6480) );
  OR2_X1 U6608 ( .A1(n5118), .A2(n6480), .ZN(n5084) );
  NAND4_X1 U6609 ( .A1(n5087), .A2(n5086), .A3(n5085), .A4(n5084), .ZN(n9937)
         );
  AND2_X1 U6610 ( .A1(n9937), .A2(n7938), .ZN(n5102) );
  NAND2_X1 U6611 ( .A1(n5089), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5090) );
  XNOR2_X1 U6612 ( .A(n5090), .B(P2_IR_REG_3__SCAN_IN), .ZN(n6479) );
  NAND2_X1 U6613 ( .A1(n4387), .A2(n6479), .ZN(n5100) );
  INV_X4 U6614 ( .A(n5091), .ZN(n7579) );
  NAND2_X1 U6615 ( .A1(n7579), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n5099) );
  NAND2_X1 U6616 ( .A1(n5093), .A2(n5092), .ZN(n5097) );
  INV_X1 U6617 ( .A(n5094), .ZN(n5095) );
  NAND2_X1 U6618 ( .A1(n5095), .A2(SI_2_), .ZN(n5096) );
  INV_X1 U6619 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6396) );
  INV_X1 U6620 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6394) );
  XNOR2_X1 U6621 ( .A(n5109), .B(n5108), .ZN(n6395) );
  OR2_X1 U6622 ( .A1(n5065), .A2(n6395), .ZN(n5098) );
  XNOR2_X1 U6623 ( .A(n6773), .B(n5669), .ZN(n5101) );
  NAND2_X1 U6624 ( .A1(n5102), .A2(n5101), .ZN(n9941) );
  INV_X1 U6625 ( .A(n5101), .ZN(n5104) );
  INV_X1 U6626 ( .A(n5102), .ZN(n5103) );
  NAND2_X1 U6627 ( .A1(n5104), .A2(n5103), .ZN(n5105) );
  NAND2_X1 U6628 ( .A1(n9941), .A2(n5105), .ZN(n9927) );
  NAND2_X1 U6629 ( .A1(n7579), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n5116) );
  NAND2_X1 U6630 ( .A1(n5110), .A2(SI_3_), .ZN(n5111) );
  OR2_X1 U6631 ( .A1(n5065), .A2(n6399), .ZN(n5115) );
  NAND2_X1 U6632 ( .A1(n5112), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5113) );
  XNOR2_X1 U6633 ( .A(n5113), .B(P2_IR_REG_4__SCAN_IN), .ZN(n6477) );
  NAND2_X1 U6634 ( .A1(n4387), .A2(n6477), .ZN(n5114) );
  XNOR2_X1 U6635 ( .A(n6756), .B(n5669), .ZN(n5124) );
  NAND2_X1 U6636 ( .A1(n5725), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5122) );
  XNOR2_X1 U6637 ( .A(P2_REG3_REG_4__SCAN_IN), .B(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n10029) );
  OR2_X1 U6638 ( .A1(n5639), .A2(n10029), .ZN(n5121) );
  INV_X1 U6639 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6468) );
  OR2_X1 U6640 ( .A1(n5619), .A2(n6468), .ZN(n5120) );
  INV_X1 U6641 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6478) );
  OR2_X1 U6642 ( .A1(n5406), .A2(n6478), .ZN(n5119) );
  NAND4_X1 U6643 ( .A1(n5122), .A2(n5121), .A3(n5120), .A4(n5119), .ZN(n7964)
         );
  NAND2_X1 U6644 ( .A1(n7964), .A2(n7938), .ZN(n5125) );
  XNOR2_X1 U6645 ( .A(n5124), .B(n5125), .ZN(n9944) );
  INV_X1 U6646 ( .A(n5124), .ZN(n5126) );
  NAND2_X1 U6647 ( .A1(n5126), .A2(n5125), .ZN(n5127) );
  AOI21_X1 U6648 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(P2_REG3_REG_4__SCAN_IN), 
        .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5128) );
  NOR2_X1 U6649 ( .A1(n5128), .A2(n5153), .ZN(n6701) );
  NAND2_X1 U6650 ( .A1(n5724), .A2(n6701), .ZN(n5134) );
  INV_X1 U6651 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n6886) );
  OR2_X1 U6652 ( .A1(n5406), .A2(n6886), .ZN(n5133) );
  INV_X1 U6653 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6464) );
  OR2_X1 U6654 ( .A1(n5619), .A2(n6464), .ZN(n5132) );
  INV_X1 U6655 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n5130) );
  OR2_X1 U6656 ( .A1(n7598), .A2(n5130), .ZN(n5131) );
  NAND4_X1 U6657 ( .A1(n5134), .A2(n5133), .A3(n5132), .A4(n5131), .ZN(n9936)
         );
  AND2_X1 U6658 ( .A1(n9936), .A2(n7938), .ZN(n5147) );
  INV_X1 U6659 ( .A(n5136), .ZN(n5137) );
  XNOR2_X1 U6660 ( .A(n5164), .B(SI_5_), .ZN(n5162) );
  XNOR2_X1 U6661 ( .A(n5163), .B(n5162), .ZN(n6403) );
  OR2_X1 U6662 ( .A1(n5065), .A2(n6403), .ZN(n5145) );
  OR2_X1 U6663 ( .A1(n5091), .A2(n8436), .ZN(n5144) );
  NOR2_X1 U6664 ( .A1(n5138), .A2(n4613), .ZN(n5139) );
  MUX2_X1 U6665 ( .A(n4613), .B(n5139), .S(P2_IR_REG_5__SCAN_IN), .Z(n5142) );
  NAND2_X1 U6666 ( .A1(n5138), .A2(n5140), .ZN(n5184) );
  INV_X1 U6667 ( .A(n5184), .ZN(n5141) );
  INV_X1 U6668 ( .A(n6503), .ZN(n6469) );
  NAND2_X1 U6669 ( .A1(n4387), .A2(n6469), .ZN(n5143) );
  XNOR2_X1 U6670 ( .A(n6890), .B(n5669), .ZN(n5146) );
  NAND2_X1 U6671 ( .A1(n5147), .A2(n5146), .ZN(n5151) );
  INV_X1 U6672 ( .A(n5146), .ZN(n5149) );
  INV_X1 U6673 ( .A(n5147), .ZN(n5148) );
  NAND2_X1 U6674 ( .A1(n5149), .A2(n5148), .ZN(n5150) );
  AND2_X1 U6675 ( .A1(n5151), .A2(n5150), .ZN(n6705) );
  NAND2_X1 U6676 ( .A1(n7593), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5161) );
  INV_X1 U6677 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6486) );
  OR2_X1 U6678 ( .A1(n6430), .A2(n6486), .ZN(n5160) );
  INV_X1 U6679 ( .A(n5174), .ZN(n5156) );
  INV_X1 U6680 ( .A(n5153), .ZN(n5154) );
  INV_X1 U6681 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n6802) );
  NAND2_X1 U6682 ( .A1(n5154), .A2(n6802), .ZN(n5155) );
  NAND2_X1 U6683 ( .A1(n5156), .A2(n5155), .ZN(n6799) );
  OR2_X1 U6684 ( .A1(n5639), .A2(n6799), .ZN(n5159) );
  INV_X1 U6685 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n5157) );
  OR2_X1 U6686 ( .A1(n7598), .A2(n5157), .ZN(n5158) );
  OR2_X1 U6687 ( .A1(n7737), .A2(n5668), .ZN(n5172) );
  NAND2_X1 U6688 ( .A1(n7579), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n5169) );
  INV_X1 U6689 ( .A(n5164), .ZN(n5165) );
  NAND2_X1 U6690 ( .A1(n5165), .A2(SI_5_), .ZN(n5166) );
  XNOR2_X1 U6691 ( .A(n5182), .B(SI_6_), .ZN(n5180) );
  NAND2_X1 U6692 ( .A1(n5184), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5167) );
  XNOR2_X1 U6693 ( .A(n5167), .B(P2_IR_REG_6__SCAN_IN), .ZN(n6505) );
  NAND2_X1 U6694 ( .A1(n4387), .A2(n6505), .ZN(n5168) );
  XNOR2_X1 U6695 ( .A(n10070), .B(n5669), .ZN(n5170) );
  XNOR2_X1 U6696 ( .A(n5172), .B(n5170), .ZN(n6797) );
  INV_X1 U6697 ( .A(n5170), .ZN(n5171) );
  NAND2_X1 U6698 ( .A1(n5172), .A2(n5171), .ZN(n5173) );
  NAND2_X1 U6699 ( .A1(n7593), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5179) );
  INV_X1 U6700 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6512) );
  OR2_X1 U6701 ( .A1(n5406), .A2(n6512), .ZN(n5178) );
  NAND2_X1 U6702 ( .A1(n5174), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5210) );
  OAI21_X1 U6703 ( .B1(n5174), .B2(P2_REG3_REG_7__SCAN_IN), .A(n5210), .ZN(
        n6930) );
  OR2_X1 U6704 ( .A1(n5639), .A2(n6930), .ZN(n5177) );
  INV_X1 U6705 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n5175) );
  OR2_X1 U6706 ( .A1(n7598), .A2(n5175), .ZN(n5176) );
  NAND4_X1 U6707 ( .A1(n5179), .A2(n5178), .A3(n5177), .A4(n5176), .ZN(n9993)
         );
  AND2_X1 U6708 ( .A1(n9993), .A2(n7938), .ZN(n5190) );
  NAND2_X1 U6709 ( .A1(n7579), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n5188) );
  INV_X1 U6710 ( .A(n5182), .ZN(n5183) );
  MUX2_X1 U6711 ( .A(n6410), .B(n6413), .S(n7515), .Z(n5198) );
  XNOR2_X1 U6712 ( .A(n5198), .B(SI_7_), .ZN(n5196) );
  XNOR2_X1 U6713 ( .A(n5197), .B(n5196), .ZN(n6412) );
  OR2_X1 U6714 ( .A1(n5065), .A2(n6412), .ZN(n5187) );
  NAND2_X1 U6715 ( .A1(n5206), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5185) );
  XNOR2_X1 U6716 ( .A(n5185), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6511) );
  NAND2_X1 U6717 ( .A1(n4387), .A2(n6511), .ZN(n5186) );
  XNOR2_X1 U6718 ( .A(n10075), .B(n5669), .ZN(n5189) );
  NAND2_X1 U6719 ( .A1(n5190), .A2(n5189), .ZN(n5195) );
  INV_X1 U6720 ( .A(n5189), .ZN(n5192) );
  INV_X1 U6721 ( .A(n5190), .ZN(n5191) );
  NAND2_X1 U6722 ( .A1(n5192), .A2(n5191), .ZN(n5193) );
  NAND2_X1 U6723 ( .A1(n5195), .A2(n5193), .ZN(n6849) );
  INV_X1 U6724 ( .A(n5198), .ZN(n5199) );
  NAND2_X1 U6725 ( .A1(n5199), .A2(SI_7_), .ZN(n5200) );
  INV_X1 U6726 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6417) );
  MUX2_X1 U6727 ( .A(n6417), .B(n6415), .S(n7515), .Z(n5202) );
  INV_X1 U6728 ( .A(SI_8_), .ZN(n5201) );
  NAND2_X1 U6729 ( .A1(n5202), .A2(n5201), .ZN(n5225) );
  INV_X1 U6730 ( .A(n5202), .ZN(n5203) );
  NAND2_X1 U6731 ( .A1(n5203), .A2(SI_8_), .ZN(n5204) );
  NAND2_X1 U6732 ( .A1(n5225), .A2(n5204), .ZN(n5223) );
  INV_X1 U6733 ( .A(n5223), .ZN(n5205) );
  XNOR2_X1 U6734 ( .A(n5224), .B(n5205), .ZN(n6416) );
  OR2_X1 U6735 ( .A1(n6416), .A2(n5065), .ZN(n5209) );
  OAI21_X1 U6736 ( .B1(n5206), .B2(P2_IR_REG_7__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5207) );
  XNOR2_X1 U6737 ( .A(n5207), .B(P2_IR_REG_8__SCAN_IN), .ZN(n6528) );
  AOI22_X1 U6738 ( .A1(n7579), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n4387), .B2(
        n6528), .ZN(n5208) );
  NAND2_X1 U6739 ( .A1(n5209), .A2(n5208), .ZN(n9982) );
  XNOR2_X1 U6740 ( .A(n9982), .B(n5635), .ZN(n5217) );
  NAND2_X1 U6741 ( .A1(n7593), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5216) );
  INV_X1 U6742 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n10003) );
  OR2_X1 U6743 ( .A1(n6430), .A2(n10003), .ZN(n5215) );
  AND2_X1 U6744 ( .A1(n5210), .A2(n6899), .ZN(n5211) );
  OR2_X1 U6745 ( .A1(n5211), .A2(n5235), .ZN(n10002) );
  OR2_X1 U6746 ( .A1(n5639), .A2(n10002), .ZN(n5214) );
  INV_X1 U6747 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n5212) );
  OR2_X1 U6748 ( .A1(n7598), .A2(n5212), .ZN(n5213) );
  NAND4_X1 U6749 ( .A1(n5216), .A2(n5215), .A3(n5214), .A4(n5213), .ZN(n7961)
         );
  AND2_X1 U6750 ( .A1(n7961), .A2(n7938), .ZN(n5218) );
  NAND2_X1 U6751 ( .A1(n5217), .A2(n5218), .ZN(n5222) );
  INV_X1 U6752 ( .A(n5217), .ZN(n5220) );
  INV_X1 U6753 ( .A(n5218), .ZN(n5219) );
  NAND2_X1 U6754 ( .A1(n5220), .A2(n5219), .ZN(n5221) );
  AND2_X1 U6755 ( .A1(n5222), .A2(n5221), .ZN(n6897) );
  MUX2_X1 U6756 ( .A(n6422), .B(n6419), .S(n7515), .Z(n5227) );
  INV_X1 U6757 ( .A(SI_9_), .ZN(n5226) );
  NAND2_X1 U6758 ( .A1(n5227), .A2(n5226), .ZN(n5246) );
  INV_X1 U6759 ( .A(n5227), .ZN(n5228) );
  NAND2_X1 U6760 ( .A1(n5228), .A2(SI_9_), .ZN(n5229) );
  XNOR2_X1 U6761 ( .A(n5245), .B(n4992), .ZN(n6418) );
  NAND2_X1 U6762 ( .A1(n6418), .A2(n7879), .ZN(n5234) );
  AND2_X1 U6763 ( .A1(n5230), .A2(n5138), .ZN(n5231) );
  OR2_X1 U6764 ( .A1(n5231), .A2(n4613), .ZN(n5232) );
  XNOR2_X1 U6765 ( .A(n5232), .B(P2_IR_REG_9__SCAN_IN), .ZN(n6662) );
  AOI22_X1 U6766 ( .A1(n7579), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n4387), .B2(
        n6662), .ZN(n5233) );
  NAND2_X1 U6767 ( .A1(n5234), .A2(n5233), .ZN(n7144) );
  XNOR2_X1 U6768 ( .A(n7144), .B(n5635), .ZN(n5241) );
  NAND2_X1 U6769 ( .A1(n7593), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5240) );
  INV_X1 U6770 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7109) );
  OR2_X1 U6771 ( .A1(n6430), .A2(n7109), .ZN(n5239) );
  NAND2_X1 U6772 ( .A1(n5235), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5256) );
  OR2_X1 U6773 ( .A1(n5235), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5236) );
  NAND2_X1 U6774 ( .A1(n5256), .A2(n5236), .ZN(n7123) );
  OR2_X1 U6775 ( .A1(n5639), .A2(n7123), .ZN(n5238) );
  OR2_X1 U6776 ( .A1(n7598), .A2(n10092), .ZN(n5237) );
  OR2_X1 U6777 ( .A1(n9996), .A2(n5668), .ZN(n5242) );
  XNOR2_X1 U6778 ( .A(n5241), .B(n5242), .ZN(n7119) );
  INV_X1 U6779 ( .A(n5241), .ZN(n5243) );
  NAND2_X1 U6780 ( .A1(n5243), .A2(n5242), .ZN(n5244) );
  MUX2_X1 U6781 ( .A(n8552), .B(n8588), .S(n7515), .Z(n5249) );
  INV_X1 U6782 ( .A(SI_10_), .ZN(n5248) );
  NAND2_X1 U6783 ( .A1(n5249), .A2(n5248), .ZN(n5270) );
  INV_X1 U6784 ( .A(n5249), .ZN(n5250) );
  NAND2_X1 U6785 ( .A1(n5250), .A2(SI_10_), .ZN(n5251) );
  NAND2_X1 U6786 ( .A1(n5253), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5254) );
  XNOR2_X1 U6787 ( .A(n5254), .B(P2_IR_REG_10__SCAN_IN), .ZN(n7968) );
  AOI22_X1 U6788 ( .A1(n7579), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n4387), .B2(
        n7968), .ZN(n5255) );
  XNOR2_X1 U6789 ( .A(n9916), .B(n5635), .ZN(n5263) );
  NAND2_X1 U6790 ( .A1(n7593), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5262) );
  INV_X1 U6791 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7155) );
  OR2_X1 U6792 ( .A1(n6430), .A2(n7155), .ZN(n5261) );
  NAND2_X1 U6793 ( .A1(n5256), .A2(n8562), .ZN(n5257) );
  NAND2_X1 U6794 ( .A1(n5304), .A2(n5257), .ZN(n9923) );
  OR2_X1 U6795 ( .A1(n5639), .A2(n9923), .ZN(n5260) );
  INV_X1 U6796 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n5258) );
  OR2_X1 U6797 ( .A1(n7598), .A2(n5258), .ZN(n5259) );
  NOR2_X1 U6798 ( .A1(n9958), .A2(n5668), .ZN(n5264) );
  NAND2_X1 U6799 ( .A1(n5263), .A2(n5264), .ZN(n5268) );
  INV_X1 U6800 ( .A(n5263), .ZN(n5266) );
  INV_X1 U6801 ( .A(n5264), .ZN(n5265) );
  NAND2_X1 U6802 ( .A1(n5266), .A2(n5265), .ZN(n5267) );
  AND2_X1 U6803 ( .A1(n5268), .A2(n5267), .ZN(n9912) );
  NAND2_X1 U6804 ( .A1(n9911), .A2(n5268), .ZN(n9952) );
  MUX2_X1 U6805 ( .A(n6439), .B(n6429), .S(n7515), .Z(n5285) );
  XNOR2_X1 U6806 ( .A(n5285), .B(SI_11_), .ZN(n5284) );
  XNOR2_X1 U6807 ( .A(n5289), .B(n5284), .ZN(n6428) );
  NAND2_X1 U6808 ( .A1(n6428), .A2(n7879), .ZN(n5274) );
  OR2_X1 U6809 ( .A1(n5253), .A2(P2_IR_REG_10__SCAN_IN), .ZN(n5294) );
  NAND2_X1 U6810 ( .A1(n5294), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5272) );
  XNOR2_X1 U6811 ( .A(n5272), .B(P2_IR_REG_11__SCAN_IN), .ZN(n6684) );
  AOI22_X1 U6812 ( .A1(n7579), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n4387), .B2(
        n6684), .ZN(n5273) );
  NAND2_X1 U6813 ( .A1(n5274), .A2(n5273), .ZN(n9956) );
  XNOR2_X1 U6814 ( .A(n9956), .B(n5669), .ZN(n5280) );
  NAND2_X1 U6815 ( .A1(n5725), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5279) );
  INV_X1 U6816 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n5302) );
  XNOR2_X1 U6817 ( .A(n5304), .B(n5302), .ZN(n9965) );
  OR2_X1 U6818 ( .A1(n5639), .A2(n9965), .ZN(n5278) );
  INV_X1 U6819 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n5275) );
  OR2_X1 U6820 ( .A1(n5619), .A2(n5275), .ZN(n5277) );
  INV_X1 U6821 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7216) );
  OR2_X1 U6822 ( .A1(n6430), .A2(n7216), .ZN(n5276) );
  NOR2_X1 U6823 ( .A1(n7324), .A2(n5668), .ZN(n5281) );
  XNOR2_X1 U6824 ( .A(n5280), .B(n5281), .ZN(n9951) );
  INV_X1 U6825 ( .A(n5280), .ZN(n5282) );
  NAND2_X1 U6826 ( .A1(n5282), .A2(n5281), .ZN(n5283) );
  NAND2_X1 U6827 ( .A1(n9950), .A2(n5283), .ZN(n7320) );
  INV_X1 U6828 ( .A(n5284), .ZN(n5288) );
  INV_X1 U6829 ( .A(n5285), .ZN(n5286) );
  NAND2_X1 U6830 ( .A1(n5286), .A2(SI_11_), .ZN(n5287) );
  MUX2_X1 U6831 ( .A(n8556), .B(n6444), .S(n7515), .Z(n5291) );
  INV_X1 U6832 ( .A(SI_12_), .ZN(n5290) );
  NAND2_X1 U6833 ( .A1(n5291), .A2(n5290), .ZN(n5317) );
  INV_X1 U6834 ( .A(n5291), .ZN(n5292) );
  NAND2_X1 U6835 ( .A1(n5292), .A2(SI_12_), .ZN(n5293) );
  NAND2_X1 U6836 ( .A1(n5317), .A2(n5293), .ZN(n5315) );
  XNOR2_X1 U6837 ( .A(n5316), .B(n5315), .ZN(n6443) );
  NAND2_X1 U6838 ( .A1(n6443), .A2(n7879), .ZN(n5300) );
  NOR2_X1 U6839 ( .A1(n5294), .A2(P2_IR_REG_11__SCAN_IN), .ZN(n5297) );
  OR2_X1 U6840 ( .A1(n5297), .A2(n4613), .ZN(n5295) );
  MUX2_X1 U6841 ( .A(n5295), .B(P2_IR_REG_31__SCAN_IN), .S(n5296), .Z(n5298)
         );
  NAND2_X1 U6842 ( .A1(n5297), .A2(n5296), .ZN(n5324) );
  AOI22_X1 U6843 ( .A1(n7579), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n4387), .B2(
        n6815), .ZN(n5299) );
  XNOR2_X1 U6844 ( .A(n7414), .B(n5669), .ZN(n5310) );
  NAND2_X1 U6845 ( .A1(n5725), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5309) );
  INV_X1 U6846 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7307) );
  OR2_X1 U6847 ( .A1(n6430), .A2(n7307), .ZN(n5308) );
  INV_X1 U6848 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n6685) );
  OR2_X1 U6849 ( .A1(n5619), .A2(n6685), .ZN(n5307) );
  INV_X1 U6850 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n5301) );
  OAI21_X1 U6851 ( .B1(n5304), .B2(n5302), .A(n5301), .ZN(n5305) );
  NAND2_X1 U6852 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_REG3_REG_11__SCAN_IN), 
        .ZN(n5303) );
  NAND2_X1 U6853 ( .A1(n5305), .A2(n5331), .ZN(n7323) );
  OR2_X1 U6854 ( .A1(n5639), .A2(n7323), .ZN(n5306) );
  OR2_X1 U6855 ( .A1(n9953), .A2(n5668), .ZN(n5311) );
  NAND2_X1 U6856 ( .A1(n5310), .A2(n5311), .ZN(n7319) );
  NAND2_X1 U6857 ( .A1(n7320), .A2(n7319), .ZN(n5314) );
  INV_X1 U6858 ( .A(n5310), .ZN(n5313) );
  INV_X1 U6859 ( .A(n5311), .ZN(n5312) );
  NAND2_X1 U6860 ( .A1(n5313), .A2(n5312), .ZN(n7318) );
  NAND2_X1 U6861 ( .A1(n5314), .A2(n7318), .ZN(n7371) );
  MUX2_X1 U6862 ( .A(n6455), .B(n5318), .S(n7515), .Z(n5320) );
  NAND2_X1 U6863 ( .A1(n5320), .A2(n5319), .ZN(n5342) );
  INV_X1 U6864 ( .A(n5320), .ZN(n5321) );
  NAND2_X1 U6865 ( .A1(n5321), .A2(SI_13_), .ZN(n5322) );
  NAND2_X1 U6866 ( .A1(n6452), .A2(n7879), .ZN(n5327) );
  NAND2_X1 U6867 ( .A1(n5324), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5323) );
  MUX2_X1 U6868 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5323), .S(
        P2_IR_REG_13__SCAN_IN), .Z(n5325) );
  AOI22_X1 U6869 ( .A1(n7579), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n4387), .B2(
        n6866), .ZN(n5326) );
  XNOR2_X1 U6870 ( .A(n9706), .B(n5669), .ZN(n5337) );
  NAND2_X1 U6871 ( .A1(n5725), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5336) );
  INV_X1 U6872 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n5328) );
  OR2_X1 U6873 ( .A1(n5619), .A2(n5328), .ZN(n5335) );
  INV_X1 U6874 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n7424) );
  OR2_X1 U6875 ( .A1(n5406), .A2(n7424), .ZN(n5334) );
  INV_X1 U6876 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5330) );
  NAND2_X1 U6877 ( .A1(n5331), .A2(n5330), .ZN(n5332) );
  NAND2_X1 U6878 ( .A1(n5352), .A2(n5332), .ZN(n7423) );
  OR2_X1 U6879 ( .A1(n5639), .A2(n7423), .ZN(n5333) );
  NOR2_X1 U6880 ( .A1(n7479), .A2(n5668), .ZN(n5338) );
  XNOR2_X1 U6881 ( .A(n5337), .B(n5338), .ZN(n7372) );
  INV_X1 U6882 ( .A(n5337), .ZN(n5339) );
  NAND2_X1 U6883 ( .A1(n5339), .A2(n5338), .ZN(n5340) );
  MUX2_X1 U6884 ( .A(n6458), .B(n6457), .S(n7515), .Z(n5366) );
  XNOR2_X1 U6885 ( .A(n5366), .B(SI_14_), .ZN(n5365) );
  XNOR2_X1 U6886 ( .A(n5370), .B(n5365), .ZN(n6456) );
  NAND2_X1 U6887 ( .A1(n6456), .A2(n7879), .ZN(n5349) );
  NAND2_X1 U6888 ( .A1(n5344), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5346) );
  NAND2_X1 U6889 ( .A1(n5346), .A2(n5345), .ZN(n5375) );
  OR2_X1 U6890 ( .A1(n5346), .A2(n5345), .ZN(n5347) );
  AOI22_X1 U6891 ( .A1(n7579), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n4387), .B2(
        n7248), .ZN(n5348) );
  XNOR2_X1 U6892 ( .A(n7497), .B(n5669), .ZN(n5358) );
  NAND2_X1 U6893 ( .A1(n5725), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5357) );
  INV_X1 U6894 ( .A(n5352), .ZN(n5350) );
  NAND2_X1 U6895 ( .A1(n5350), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5386) );
  INV_X1 U6896 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n5351) );
  NAND2_X1 U6897 ( .A1(n5352), .A2(n5351), .ZN(n5353) );
  NAND2_X1 U6898 ( .A1(n5386), .A2(n5353), .ZN(n7478) );
  OR2_X1 U6899 ( .A1(n5639), .A2(n7478), .ZN(n5356) );
  INV_X1 U6900 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n6867) );
  OR2_X1 U6901 ( .A1(n5619), .A2(n6867), .ZN(n5355) );
  INV_X1 U6902 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n7449) );
  OR2_X1 U6903 ( .A1(n6430), .A2(n7449), .ZN(n5354) );
  OR2_X1 U6904 ( .A1(n7716), .A2(n5668), .ZN(n5359) );
  NAND2_X1 U6905 ( .A1(n5358), .A2(n5359), .ZN(n5364) );
  INV_X1 U6906 ( .A(n5358), .ZN(n5361) );
  INV_X1 U6907 ( .A(n5359), .ZN(n5360) );
  NAND2_X1 U6908 ( .A1(n5361), .A2(n5360), .ZN(n5362) );
  NAND2_X1 U6909 ( .A1(n5364), .A2(n5362), .ZN(n7476) );
  INV_X1 U6910 ( .A(n5382), .ZN(n5380) );
  INV_X1 U6911 ( .A(n5365), .ZN(n5369) );
  INV_X1 U6912 ( .A(n5366), .ZN(n5367) );
  NAND2_X1 U6913 ( .A1(n5367), .A2(SI_14_), .ZN(n5368) );
  MUX2_X1 U6914 ( .A(n6653), .B(n6655), .S(n7515), .Z(n5372) );
  NAND2_X1 U6915 ( .A1(n5372), .A2(n5371), .ZN(n5394) );
  INV_X1 U6916 ( .A(n5372), .ZN(n5373) );
  NAND2_X1 U6917 ( .A1(n5373), .A2(SI_15_), .ZN(n5374) );
  NAND2_X1 U6918 ( .A1(n5394), .A2(n5374), .ZN(n5395) );
  XNOR2_X1 U6919 ( .A(n5396), .B(n5395), .ZN(n6652) );
  NAND2_X1 U6920 ( .A1(n6652), .A2(n7879), .ZN(n5378) );
  NAND2_X1 U6921 ( .A1(n5375), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5376) );
  XNOR2_X1 U6922 ( .A(n5376), .B(P2_IR_REG_15__SCAN_IN), .ZN(n7287) );
  AOI22_X1 U6923 ( .A1(n7579), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n4387), .B2(
        n7287), .ZN(n5377) );
  XNOR2_X1 U6924 ( .A(n7568), .B(n5669), .ZN(n5381) );
  INV_X1 U6925 ( .A(n5381), .ZN(n5379) );
  NAND2_X1 U6926 ( .A1(n5382), .A2(n5381), .ZN(n5393) );
  NAND2_X1 U6927 ( .A1(n7594), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n5392) );
  INV_X1 U6928 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n5384) );
  OR2_X1 U6929 ( .A1(n5619), .A2(n5384), .ZN(n5391) );
  INV_X1 U6930 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n5385) );
  NAND2_X1 U6931 ( .A1(n5386), .A2(n5385), .ZN(n5387) );
  NAND2_X1 U6932 ( .A1(n5409), .A2(n5387), .ZN(n7715) );
  OR2_X1 U6933 ( .A1(n5639), .A2(n7715), .ZN(n5390) );
  INV_X1 U6934 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n5388) );
  OR2_X1 U6935 ( .A1(n7598), .A2(n5388), .ZN(n5389) );
  OR2_X1 U6936 ( .A1(n8242), .A2(n5668), .ZN(n7712) );
  MUX2_X1 U6937 ( .A(n8594), .B(n6700), .S(n7515), .Z(n5398) );
  INV_X1 U6938 ( .A(SI_16_), .ZN(n5397) );
  NAND2_X1 U6939 ( .A1(n5398), .A2(n5397), .ZN(n5421) );
  INV_X1 U6940 ( .A(n5398), .ZN(n5399) );
  NAND2_X1 U6941 ( .A1(n5399), .A2(SI_16_), .ZN(n5400) );
  XNOR2_X1 U6942 ( .A(n5420), .B(n5419), .ZN(n6656) );
  NAND2_X1 U6943 ( .A1(n6656), .A2(n7879), .ZN(n5404) );
  NAND2_X1 U6944 ( .A1(n5401), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5402) );
  XNOR2_X1 U6945 ( .A(n5402), .B(P2_IR_REG_16__SCAN_IN), .ZN(n7985) );
  AOI22_X1 U6946 ( .A1(n7579), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n4387), .B2(
        n7985), .ZN(n5403) );
  XNOR2_X1 U6947 ( .A(n8333), .B(n5669), .ZN(n5417) );
  NAND2_X1 U6948 ( .A1(n5725), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5414) );
  INV_X1 U6949 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n7281) );
  OR2_X1 U6950 ( .A1(n5619), .A2(n7281), .ZN(n5413) );
  INV_X1 U6951 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n5405) );
  OR2_X1 U6952 ( .A1(n6430), .A2(n5405), .ZN(n5412) );
  INV_X1 U6953 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n5408) );
  NAND2_X1 U6954 ( .A1(n5409), .A2(n5408), .ZN(n5410) );
  NAND2_X1 U6955 ( .A1(n5427), .A2(n5410), .ZN(n7646) );
  OR2_X1 U6956 ( .A1(n5639), .A2(n7646), .ZN(n5411) );
  NOR2_X1 U6957 ( .A1(n8228), .A2(n5668), .ZN(n5415) );
  XNOR2_X1 U6958 ( .A(n5417), .B(n5415), .ZN(n7644) );
  INV_X1 U6959 ( .A(n5415), .ZN(n5416) );
  NAND2_X1 U6960 ( .A1(n5417), .A2(n5416), .ZN(n5418) );
  MUX2_X1 U6961 ( .A(n8587), .B(n5423), .S(n7515), .Z(n5438) );
  XNOR2_X1 U6962 ( .A(n5438), .B(SI_17_), .ZN(n5437) );
  XNOR2_X1 U6963 ( .A(n5442), .B(n5437), .ZN(n6709) );
  NAND2_X1 U6964 ( .A1(n6709), .A2(n7879), .ZN(n5426) );
  NAND2_X1 U6965 ( .A1(n4454), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5424) );
  XNOR2_X1 U6966 ( .A(n5424), .B(P2_IR_REG_17__SCAN_IN), .ZN(n7996) );
  AOI22_X1 U6967 ( .A1(n7579), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n4387), .B2(
        n7996), .ZN(n5425) );
  XNOR2_X1 U6968 ( .A(n8329), .B(n5635), .ZN(n5435) );
  NAND2_X1 U6969 ( .A1(n7593), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n5433) );
  INV_X1 U6970 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8219) );
  OR2_X1 U6971 ( .A1(n6430), .A2(n8219), .ZN(n5432) );
  NAND2_X1 U6972 ( .A1(n5427), .A2(n8406), .ZN(n5428) );
  NAND2_X1 U6973 ( .A1(n5448), .A2(n5428), .ZN(n8218) );
  OR2_X1 U6974 ( .A1(n5639), .A2(n8218), .ZN(n5431) );
  INV_X1 U6975 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n5429) );
  OR2_X1 U6976 ( .A1(n7598), .A2(n5429), .ZN(n5430) );
  NOR2_X1 U6977 ( .A1(n8240), .A2(n5668), .ZN(n5434) );
  XNOR2_X1 U6978 ( .A(n5435), .B(n5434), .ZN(n7651) );
  NAND2_X1 U6979 ( .A1(n5435), .A2(n5434), .ZN(n5436) );
  INV_X1 U6980 ( .A(n5437), .ZN(n5441) );
  INV_X1 U6981 ( .A(n5438), .ZN(n5439) );
  NAND2_X1 U6982 ( .A1(n5439), .A2(SI_17_), .ZN(n5440) );
  MUX2_X1 U6983 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n7515), .Z(n5462) );
  XNOR2_X1 U6984 ( .A(n5462), .B(SI_18_), .ZN(n5459) );
  XNOR2_X1 U6985 ( .A(n5461), .B(n5459), .ZN(n6806) );
  NAND2_X1 U6986 ( .A1(n6806), .A2(n7879), .ZN(n5445) );
  XNOR2_X1 U6987 ( .A(n5443), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8011) );
  AOI22_X1 U6988 ( .A1(n7579), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n4387), .B2(
        n8011), .ZN(n5444) );
  XNOR2_X1 U6989 ( .A(n8324), .B(n5635), .ZN(n5456) );
  NAND2_X1 U6990 ( .A1(n5725), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n5453) );
  INV_X1 U6991 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n7994) );
  OR2_X1 U6992 ( .A1(n5619), .A2(n7994), .ZN(n5452) );
  INV_X1 U6993 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n5447) );
  NAND2_X1 U6994 ( .A1(n5448), .A2(n5447), .ZN(n5449) );
  NAND2_X1 U6995 ( .A1(n5472), .A2(n5449), .ZN(n8206) );
  OR2_X1 U6996 ( .A1(n5639), .A2(n8206), .ZN(n5451) );
  INV_X1 U6997 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8009) );
  OR2_X1 U6998 ( .A1(n6430), .A2(n8009), .ZN(n5450) );
  NAND4_X1 U6999 ( .A1(n5453), .A2(n5452), .A3(n5451), .A4(n5450), .ZN(n7953)
         );
  NAND2_X1 U7000 ( .A1(n7953), .A2(n7938), .ZN(n5454) );
  XNOR2_X1 U7001 ( .A(n5456), .B(n5454), .ZN(n7695) );
  NAND2_X1 U7002 ( .A1(n7694), .A2(n7695), .ZN(n5458) );
  INV_X1 U7003 ( .A(n5454), .ZN(n5455) );
  NAND2_X1 U7004 ( .A1(n5456), .A2(n5455), .ZN(n5457) );
  INV_X1 U7005 ( .A(n7621), .ZN(n5484) );
  INV_X1 U7006 ( .A(n5459), .ZN(n5460) );
  NAND2_X1 U7007 ( .A1(n5462), .A2(SI_18_), .ZN(n5463) );
  MUX2_X1 U7008 ( .A(n8340), .B(n6878), .S(n7515), .Z(n5466) );
  INV_X1 U7009 ( .A(SI_19_), .ZN(n5465) );
  NAND2_X1 U7010 ( .A1(n5466), .A2(n5465), .ZN(n5488) );
  INV_X1 U7011 ( .A(n5466), .ZN(n5467) );
  NAND2_X1 U7012 ( .A1(n5467), .A2(SI_19_), .ZN(n5468) );
  NAND2_X1 U7013 ( .A1(n5488), .A2(n5468), .ZN(n5486) );
  XNOR2_X1 U7014 ( .A(n5487), .B(n5486), .ZN(n6877) );
  NAND2_X1 U7015 ( .A1(n6877), .A2(n7879), .ZN(n5470) );
  INV_X1 U7016 ( .A(n8020), .ZN(n8081) );
  AOI22_X1 U7017 ( .A1(n7579), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n5088), .B2(
        n8081), .ZN(n5469) );
  XNOR2_X1 U7018 ( .A(n8318), .B(n5669), .ZN(n5478) );
  NAND2_X1 U7019 ( .A1(n7594), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n5477) );
  INV_X1 U7020 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n5471) );
  OR2_X1 U7021 ( .A1(n5619), .A2(n5471), .ZN(n5476) );
  NAND2_X1 U7022 ( .A1(n5472), .A2(n8438), .ZN(n5473) );
  NAND2_X1 U7023 ( .A1(n5495), .A2(n5473), .ZN(n8187) );
  OR2_X1 U7024 ( .A1(n5639), .A2(n8187), .ZN(n5475) );
  INV_X1 U7025 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n8516) );
  OR2_X1 U7026 ( .A1(n7598), .A2(n8516), .ZN(n5474) );
  NAND4_X1 U7027 ( .A1(n5477), .A2(n5476), .A3(n5475), .A4(n5474), .ZN(n7952)
         );
  NAND2_X1 U7028 ( .A1(n7952), .A2(n7938), .ZN(n5479) );
  NAND2_X1 U7029 ( .A1(n5478), .A2(n5479), .ZN(n5485) );
  INV_X1 U7030 ( .A(n5478), .ZN(n5481) );
  INV_X1 U7031 ( .A(n5479), .ZN(n5480) );
  NAND2_X1 U7032 ( .A1(n5481), .A2(n5480), .ZN(n5482) );
  NAND2_X1 U7033 ( .A1(n5485), .A2(n5482), .ZN(n7620) );
  NAND2_X2 U7034 ( .A1(n5484), .A2(n5483), .ZN(n7618) );
  MUX2_X1 U7035 ( .A(n8578), .B(n6999), .S(n7515), .Z(n5489) );
  INV_X1 U7036 ( .A(SI_20_), .ZN(n8511) );
  NAND2_X1 U7037 ( .A1(n5489), .A2(n8511), .ZN(n5509) );
  INV_X1 U7038 ( .A(n5489), .ZN(n5490) );
  NAND2_X1 U7039 ( .A1(n5490), .A2(SI_20_), .ZN(n5491) );
  XNOR2_X1 U7040 ( .A(n5507), .B(n5508), .ZN(n6998) );
  NAND2_X1 U7041 ( .A1(n6998), .A2(n7879), .ZN(n5493) );
  NAND2_X1 U7042 ( .A1(n7579), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n5492) );
  XNOR2_X1 U7043 ( .A(n8314), .B(n5635), .ZN(n5503) );
  INV_X1 U7044 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n7671) );
  NAND2_X1 U7045 ( .A1(n5495), .A2(n7671), .ZN(n5496) );
  NAND2_X1 U7046 ( .A1(n5513), .A2(n5496), .ZN(n8177) );
  OR2_X1 U7047 ( .A1(n8177), .A2(n5639), .ZN(n5502) );
  NAND2_X1 U7048 ( .A1(n7594), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n5501) );
  INV_X1 U7049 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n5497) );
  OR2_X1 U7050 ( .A1(n5619), .A2(n5497), .ZN(n5500) );
  INV_X1 U7051 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n5498) );
  OR2_X1 U7052 ( .A1(n7598), .A2(n5498), .ZN(n5499) );
  NOR2_X1 U7053 ( .A1(n7951), .A2(n5668), .ZN(n5504) );
  XNOR2_X1 U7054 ( .A(n5503), .B(n5504), .ZN(n7670) );
  INV_X1 U7055 ( .A(n5503), .ZN(n5506) );
  INV_X1 U7056 ( .A(n5504), .ZN(n5505) );
  MUX2_X1 U7057 ( .A(n7128), .B(n7116), .S(n7515), .Z(n5526) );
  XNOR2_X1 U7058 ( .A(n5526), .B(SI_21_), .ZN(n5524) );
  XNOR2_X1 U7059 ( .A(n5523), .B(n5524), .ZN(n7115) );
  NAND2_X1 U7060 ( .A1(n7115), .A2(n7879), .ZN(n5511) );
  NAND2_X1 U7061 ( .A1(n7579), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n5510) );
  XNOR2_X1 U7062 ( .A(n8159), .B(n5635), .ZN(n5520) );
  INV_X1 U7063 ( .A(n5513), .ZN(n5512) );
  INV_X1 U7064 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n8501) );
  NAND2_X1 U7065 ( .A1(n5513), .A2(n8501), .ZN(n5514) );
  NAND2_X1 U7066 ( .A1(n5534), .A2(n5514), .ZN(n8156) );
  OR2_X1 U7067 ( .A1(n8156), .A2(n5639), .ZN(n5519) );
  NAND2_X1 U7068 ( .A1(n7593), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n5516) );
  NAND2_X1 U7069 ( .A1(n5725), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n5515) );
  AND2_X1 U7070 ( .A1(n5516), .A2(n5515), .ZN(n5518) );
  NAND2_X1 U7071 ( .A1(n7594), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n5517) );
  NOR2_X1 U7072 ( .A1(n7589), .A2(n5668), .ZN(n5521) );
  XNOR2_X1 U7073 ( .A(n5520), .B(n5521), .ZN(n7627) );
  INV_X1 U7074 ( .A(n5520), .ZN(n5522) );
  INV_X1 U7075 ( .A(n5526), .ZN(n5527) );
  NAND2_X1 U7076 ( .A1(n5527), .A2(SI_21_), .ZN(n5528) );
  INV_X1 U7077 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7202) );
  MUX2_X1 U7078 ( .A(n7202), .B(n7204), .S(n7515), .Z(n5529) );
  NAND2_X1 U7079 ( .A1(n5529), .A2(n8457), .ZN(n5545) );
  INV_X1 U7080 ( .A(n5529), .ZN(n5530) );
  NAND2_X1 U7081 ( .A1(n5530), .A2(SI_22_), .ZN(n5531) );
  NAND2_X1 U7082 ( .A1(n5545), .A2(n5531), .ZN(n5543) );
  XNOR2_X1 U7083 ( .A(n5544), .B(n5543), .ZN(n7201) );
  NAND2_X1 U7084 ( .A1(n7201), .A2(n7879), .ZN(n5533) );
  NAND2_X1 U7085 ( .A1(n7579), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n5532) );
  XNOR2_X1 U7086 ( .A(n8302), .B(n5669), .ZN(n5539) );
  XNOR2_X1 U7087 ( .A(n5541), .B(n5539), .ZN(n7678) );
  INV_X1 U7088 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n7681) );
  NAND2_X1 U7089 ( .A1(n5534), .A2(n7681), .ZN(n5535) );
  NAND2_X1 U7090 ( .A1(n5572), .A2(n5535), .ZN(n7680) );
  OR2_X1 U7091 ( .A1(n7680), .A2(n5639), .ZN(n5538) );
  AOI22_X1 U7092 ( .A1(n7593), .A2(P2_REG1_REG_22__SCAN_IN), .B1(n7594), .B2(
        P2_REG2_REG_22__SCAN_IN), .ZN(n5537) );
  NAND2_X1 U7093 ( .A1(n5725), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n5536) );
  INV_X1 U7094 ( .A(n7628), .ZN(n8163) );
  NAND2_X1 U7095 ( .A1(n8163), .A2(n7938), .ZN(n7677) );
  NAND2_X1 U7096 ( .A1(n7678), .A2(n7677), .ZN(n7676) );
  INV_X1 U7097 ( .A(n5539), .ZN(n5540) );
  INV_X1 U7098 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n5546) );
  MUX2_X1 U7099 ( .A(n5546), .B(n7276), .S(n7515), .Z(n5548) );
  INV_X1 U7100 ( .A(SI_23_), .ZN(n5547) );
  NAND2_X1 U7101 ( .A1(n5548), .A2(n5547), .ZN(n5555) );
  INV_X1 U7102 ( .A(n5548), .ZN(n5549) );
  NAND2_X1 U7103 ( .A1(n5549), .A2(SI_23_), .ZN(n5550) );
  XNOR2_X1 U7104 ( .A(n5554), .B(n5553), .ZN(n7273) );
  NAND2_X1 U7105 ( .A1(n7273), .A2(n7879), .ZN(n5552) );
  NAND2_X1 U7106 ( .A1(n7579), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n5551) );
  XNOR2_X1 U7107 ( .A(n8297), .B(n5635), .ZN(n5570) );
  INV_X1 U7108 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7299) );
  MUX2_X1 U7109 ( .A(n7299), .B(n8411), .S(n7515), .Z(n5585) );
  XNOR2_X1 U7110 ( .A(n5585), .B(SI_24_), .ZN(n5582) );
  XNOR2_X1 U7111 ( .A(n5584), .B(n5582), .ZN(n7297) );
  NAND2_X1 U7112 ( .A1(n7297), .A2(n7879), .ZN(n5557) );
  NAND2_X1 U7113 ( .A1(n7579), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n5556) );
  XNOR2_X1 U7114 ( .A(n8294), .B(n5669), .ZN(n7661) );
  INV_X1 U7115 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n7612) );
  INV_X1 U7116 ( .A(n5574), .ZN(n5558) );
  NAND2_X1 U7117 ( .A1(n5558), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5594) );
  INV_X1 U7118 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n7664) );
  NAND2_X1 U7119 ( .A1(n5574), .A2(n7664), .ZN(n5559) );
  NAND2_X1 U7120 ( .A1(n5594), .A2(n5559), .ZN(n8118) );
  OR2_X1 U7121 ( .A1(n8118), .A2(n5639), .ZN(n5564) );
  INV_X1 U7122 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n8568) );
  NAND2_X1 U7123 ( .A1(n7594), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n5561) );
  NAND2_X1 U7124 ( .A1(n5725), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n5560) );
  OAI211_X1 U7125 ( .C1(n5619), .C2(n8568), .A(n5561), .B(n5560), .ZN(n5562)
         );
  INV_X1 U7126 ( .A(n5562), .ZN(n5563) );
  INV_X1 U7127 ( .A(n8094), .ZN(n8134) );
  NAND2_X1 U7128 ( .A1(n8134), .A2(n7938), .ZN(n5565) );
  AND2_X1 U7129 ( .A1(n7661), .A2(n5565), .ZN(n5568) );
  INV_X1 U7130 ( .A(n7661), .ZN(n5566) );
  INV_X1 U7131 ( .A(n5565), .ZN(n7660) );
  NAND2_X1 U7132 ( .A1(n5566), .A2(n7660), .ZN(n5567) );
  OAI21_X1 U7133 ( .B1(n7657), .B2(n5568), .A(n5567), .ZN(n5569) );
  INV_X1 U7134 ( .A(n5569), .ZN(n5581) );
  XNOR2_X1 U7135 ( .A(n5571), .B(n5570), .ZN(n7611) );
  NAND2_X1 U7136 ( .A1(n5572), .A2(n7612), .ZN(n5573) );
  AND2_X1 U7137 ( .A1(n5574), .A2(n5573), .ZN(n8130) );
  INV_X1 U7138 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n5577) );
  NAND2_X1 U7139 ( .A1(n7593), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n5576) );
  NAND2_X1 U7140 ( .A1(n7594), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n5575) );
  OAI211_X1 U7141 ( .C1(n5577), .C2(n7598), .A(n5576), .B(n5575), .ZN(n5578)
         );
  OR2_X1 U7142 ( .A1(n7840), .A2(n5668), .ZN(n7658) );
  AOI21_X1 U7143 ( .B1(n7661), .B2(n8094), .A(n7658), .ZN(n5579) );
  NAND2_X1 U7144 ( .A1(n7611), .A2(n5579), .ZN(n5580) );
  INV_X1 U7145 ( .A(n5582), .ZN(n5583) );
  INV_X1 U7146 ( .A(n5585), .ZN(n5586) );
  NAND2_X1 U7147 ( .A1(n5586), .A2(SI_24_), .ZN(n5587) );
  INV_X1 U7148 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7437) );
  INV_X1 U7149 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7434) );
  MUX2_X1 U7150 ( .A(n7437), .B(n7434), .S(n7515), .Z(n5588) );
  NAND2_X1 U7151 ( .A1(n5588), .A2(n8456), .ZN(n5606) );
  INV_X1 U7152 ( .A(n5588), .ZN(n5589) );
  NAND2_X1 U7153 ( .A1(n5589), .A2(SI_25_), .ZN(n5590) );
  NAND2_X1 U7154 ( .A1(n5606), .A2(n5590), .ZN(n5607) );
  NAND2_X1 U7155 ( .A1(n7431), .A2(n7879), .ZN(n5592) );
  NAND2_X1 U7156 ( .A1(n7579), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n5591) );
  XNOR2_X1 U7157 ( .A(n8289), .B(n5669), .ZN(n5602) );
  INV_X1 U7158 ( .A(n5594), .ZN(n5593) );
  NAND2_X1 U7159 ( .A1(n5593), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n5615) );
  INV_X1 U7160 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n7637) );
  NAND2_X1 U7161 ( .A1(n5594), .A2(n7637), .ZN(n5595) );
  NAND2_X1 U7162 ( .A1(n5615), .A2(n5595), .ZN(n8099) );
  OR2_X1 U7163 ( .A1(n8099), .A2(n5639), .ZN(n5601) );
  INV_X1 U7164 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n5598) );
  NAND2_X1 U7165 ( .A1(n7594), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n5597) );
  NAND2_X1 U7166 ( .A1(n7593), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n5596) );
  OAI211_X1 U7167 ( .C1(n5598), .C2(n7598), .A(n5597), .B(n5596), .ZN(n5599)
         );
  INV_X1 U7168 ( .A(n5599), .ZN(n5600) );
  NAND2_X1 U7169 ( .A1(n8113), .A2(n7938), .ZN(n5603) );
  NAND2_X1 U7170 ( .A1(n5602), .A2(n5603), .ZN(n7634) );
  INV_X1 U7171 ( .A(n5602), .ZN(n5605) );
  INV_X1 U7172 ( .A(n5603), .ZN(n5604) );
  NAND2_X1 U7173 ( .A1(n5605), .A2(n5604), .ZN(n7633) );
  INV_X1 U7174 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n8409) );
  INV_X1 U7175 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7439) );
  MUX2_X1 U7176 ( .A(n8409), .B(n7439), .S(n7515), .Z(n5610) );
  INV_X1 U7177 ( .A(SI_26_), .ZN(n5609) );
  NAND2_X1 U7178 ( .A1(n5610), .A2(n5609), .ZN(n5627) );
  INV_X1 U7179 ( .A(n5610), .ZN(n5611) );
  NAND2_X1 U7180 ( .A1(n5611), .A2(SI_26_), .ZN(n5612) );
  XNOR2_X1 U7181 ( .A(n5626), .B(n5625), .ZN(n7438) );
  NAND2_X1 U7182 ( .A1(n7438), .A2(n7879), .ZN(n5614) );
  NAND2_X1 U7183 ( .A1(n7579), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n5613) );
  XNOR2_X1 U7184 ( .A(n8282), .B(n5669), .ZN(n5621) );
  INV_X1 U7185 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n7704) );
  NAND2_X1 U7186 ( .A1(n5615), .A2(n7704), .ZN(n5616) );
  INV_X1 U7187 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8398) );
  NAND2_X1 U7188 ( .A1(n5725), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n5618) );
  NAND2_X1 U7189 ( .A1(n7594), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n5617) );
  OAI211_X1 U7190 ( .C1(n5619), .C2(n8398), .A(n5618), .B(n5617), .ZN(n5620)
         );
  AOI21_X1 U7191 ( .B1(n8079), .B2(n5724), .A(n5620), .ZN(n8095) );
  NOR2_X1 U7192 ( .A1(n8095), .A2(n5668), .ZN(n5622) );
  XNOR2_X1 U7193 ( .A(n5621), .B(n5622), .ZN(n7701) );
  INV_X1 U7194 ( .A(n5621), .ZN(n5623) );
  NAND2_X1 U7195 ( .A1(n5623), .A2(n5622), .ZN(n5624) );
  NAND2_X1 U7196 ( .A1(n5626), .A2(n5625), .ZN(n5628) );
  INV_X1 U7197 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n7510) );
  INV_X1 U7198 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n8476) );
  MUX2_X1 U7199 ( .A(n7510), .B(n8476), .S(n7515), .Z(n5630) );
  INV_X1 U7200 ( .A(SI_27_), .ZN(n5629) );
  NAND2_X1 U7201 ( .A1(n5630), .A2(n5629), .ZN(n5651) );
  INV_X1 U7202 ( .A(n5630), .ZN(n5631) );
  NAND2_X1 U7203 ( .A1(n5631), .A2(SI_27_), .ZN(n5632) );
  NAND2_X1 U7204 ( .A1(n7508), .A2(n7879), .ZN(n5634) );
  NAND2_X1 U7205 ( .A1(n7579), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n5633) );
  XNOR2_X1 U7206 ( .A(n8274), .B(n5635), .ZN(n5647) );
  INV_X1 U7207 ( .A(n5637), .ZN(n5636) );
  NAND2_X1 U7208 ( .A1(n5636), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n5660) );
  INV_X1 U7209 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n8421) );
  NAND2_X1 U7210 ( .A1(n5637), .A2(n8421), .ZN(n5638) );
  NAND2_X1 U7211 ( .A1(n5660), .A2(n5638), .ZN(n8056) );
  INV_X1 U7212 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n8490) );
  NAND2_X1 U7213 ( .A1(n7593), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n5641) );
  NAND2_X1 U7214 ( .A1(n7594), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n5640) );
  OAI211_X1 U7215 ( .C1(n8490), .C2(n7598), .A(n5641), .B(n5640), .ZN(n5642)
         );
  INV_X1 U7216 ( .A(n5642), .ZN(n5643) );
  NAND2_X1 U7217 ( .A1(n4696), .A2(n7938), .ZN(n5645) );
  XNOR2_X1 U7218 ( .A(n5647), .B(n5645), .ZN(n7604) );
  INV_X1 U7219 ( .A(n5645), .ZN(n5646) );
  AND2_X1 U7220 ( .A1(n5647), .A2(n5646), .ZN(n5648) );
  AOI21_X1 U7221 ( .B1(n7605), .B2(n7604), .A(n5648), .ZN(n5717) );
  INV_X1 U7222 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n5653) );
  MUX2_X1 U7223 ( .A(n5653), .B(n8681), .S(n7515), .Z(n5655) );
  INV_X1 U7224 ( .A(SI_28_), .ZN(n5654) );
  NAND2_X1 U7225 ( .A1(n5655), .A2(n5654), .ZN(n7513) );
  INV_X1 U7226 ( .A(n5655), .ZN(n5656) );
  NAND2_X1 U7227 ( .A1(n5656), .A2(SI_28_), .ZN(n5657) );
  NAND2_X1 U7228 ( .A1(n8680), .A2(n7879), .ZN(n5659) );
  NAND2_X1 U7229 ( .A1(n7579), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n5658) );
  INV_X1 U7230 ( .A(n7925), .ZN(n10050) );
  NAND2_X1 U7231 ( .A1(n8272), .A2(n10110), .ZN(n5712) );
  INV_X1 U7232 ( .A(n5712), .ZN(n5671) );
  INV_X1 U7233 ( .A(n8272), .ZN(n8049) );
  INV_X1 U7234 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n5721) );
  NAND2_X1 U7235 ( .A1(n5660), .A2(n5721), .ZN(n5661) );
  NAND2_X1 U7236 ( .A1(n8046), .A2(n5724), .ZN(n5667) );
  INV_X1 U7237 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n5664) );
  NAND2_X1 U7238 ( .A1(n7594), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n5663) );
  NAND2_X1 U7239 ( .A1(n7593), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n5662) );
  OAI211_X1 U7240 ( .C1(n5664), .C2(n7598), .A(n5663), .B(n5662), .ZN(n5665)
         );
  INV_X1 U7241 ( .A(n5665), .ZN(n5666) );
  NOR2_X1 U7242 ( .A1(n7606), .A2(n5668), .ZN(n5670) );
  XNOR2_X1 U7243 ( .A(n5670), .B(n5669), .ZN(n5711) );
  MUX2_X1 U7244 ( .A(n5671), .B(n8049), .S(n5711), .Z(n5716) );
  NAND3_X1 U7245 ( .A1(n5702), .A2(n5682), .A3(n5685), .ZN(n5672) );
  NAND2_X1 U7246 ( .A1(n5677), .A2(n5678), .ZN(n5680) );
  NAND2_X1 U7247 ( .A1(n5680), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5674) );
  MUX2_X1 U7248 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5674), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n5676) );
  OR2_X1 U7249 ( .A1(n5677), .A2(n4613), .ZN(n5679) );
  MUX2_X1 U7250 ( .A(n5679), .B(P2_IR_REG_31__SCAN_IN), .S(n5678), .Z(n5681)
         );
  NAND2_X1 U7251 ( .A1(n5681), .A2(n5680), .ZN(n7435) );
  NAND2_X1 U7252 ( .A1(n5683), .A2(n5682), .ZN(n5684) );
  INV_X1 U7253 ( .A(P2_B_REG_SCAN_IN), .ZN(n5687) );
  XOR2_X1 U7254 ( .A(n7301), .B(n5687), .Z(n5688) );
  NAND2_X1 U7255 ( .A1(n7435), .A2(n5688), .ZN(n5689) );
  INV_X1 U7256 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n10046) );
  AND2_X1 U7257 ( .A1(n7456), .A2(n7435), .ZN(n10047) );
  NOR4_X1 U7258 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_16__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n5694) );
  NOR4_X1 U7259 ( .A1(P2_D_REG_12__SCAN_IN), .A2(P2_D_REG_13__SCAN_IN), .A3(
        P2_D_REG_14__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n5693) );
  NOR4_X1 U7260 ( .A1(P2_D_REG_24__SCAN_IN), .A2(P2_D_REG_29__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n5692) );
  NOR4_X1 U7261 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_23__SCAN_IN), .ZN(n5691) );
  NAND4_X1 U7262 ( .A1(n5694), .A2(n5693), .A3(n5692), .A4(n5691), .ZN(n5699)
         );
  NOR4_X1 U7263 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_19__SCAN_IN), .A4(P2_D_REG_26__SCAN_IN), .ZN(n8391) );
  NOR2_X1 U7264 ( .A1(P2_D_REG_30__SCAN_IN), .A2(P2_D_REG_31__SCAN_IN), .ZN(
        n5697) );
  NOR4_X1 U7265 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_7__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n5696) );
  NOR4_X1 U7266 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n5695) );
  NAND4_X1 U7267 ( .A1(n8391), .A2(n5697), .A3(n5696), .A4(n5695), .ZN(n5698)
         );
  OAI21_X1 U7268 ( .B1(n5699), .B2(n5698), .A(n10036), .ZN(n6742) );
  AND2_X1 U7269 ( .A1(n6745), .A2(n6742), .ZN(n6882) );
  INV_X1 U7270 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n10043) );
  NAND2_X1 U7271 ( .A1(n10036), .A2(n10043), .ZN(n5701) );
  INV_X1 U7272 ( .A(n10044), .ZN(n5700) );
  NAND2_X1 U7273 ( .A1(n6882), .A2(n6777), .ZN(n5718) );
  INV_X1 U7274 ( .A(n5718), .ZN(n5706) );
  NAND2_X1 U7275 ( .A1(n5706), .A2(n7943), .ZN(n5709) );
  NAND2_X1 U7276 ( .A1(n7943), .A2(n7536), .ZN(n5707) );
  NAND2_X1 U7277 ( .A1(n5709), .A2(n5707), .ZN(n5708) );
  INV_X1 U7278 ( .A(n5709), .ZN(n5731) );
  NOR2_X1 U7279 ( .A1(n10024), .A2(n6762), .ZN(n5710) );
  AOI21_X1 U7280 ( .B1(n8272), .B2(n9957), .A(n9949), .ZN(n5715) );
  MUX2_X1 U7281 ( .A(n8272), .B(n5712), .S(n5711), .Z(n5713) );
  NOR2_X1 U7282 ( .A1(n5717), .A2(n5713), .ZN(n5714) );
  INV_X1 U7283 ( .A(n8046), .ZN(n5722) );
  NAND2_X1 U7284 ( .A1(n5718), .A2(n6883), .ZN(n7531) );
  AND2_X1 U7285 ( .A1(n6762), .A2(n6761), .ZN(n6741) );
  INV_X1 U7286 ( .A(n6741), .ZN(n5719) );
  NAND4_X1 U7287 ( .A1(n7531), .A2(n6342), .A3(n6423), .A4(n5719), .ZN(n5720)
         );
  OAI22_X1 U7288 ( .A1(n5722), .A2(n9966), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5721), .ZN(n5737) );
  INV_X1 U7289 ( .A(n5723), .ZN(n7583) );
  NAND2_X1 U7290 ( .A1(n7583), .A2(n5724), .ZN(n5730) );
  INV_X1 U7291 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n8566) );
  NAND2_X1 U7292 ( .A1(n7593), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n5727) );
  NAND2_X1 U7293 ( .A1(n5725), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n5726) );
  OAI211_X1 U7294 ( .C1(n8566), .C2(n6430), .A(n5727), .B(n5726), .ZN(n5728)
         );
  INV_X1 U7295 ( .A(n5728), .ZN(n5729) );
  NAND2_X1 U7296 ( .A1(n5730), .A2(n5729), .ZN(n7949) );
  INV_X1 U7297 ( .A(n7949), .ZN(n8041) );
  INV_X1 U7298 ( .A(n6761), .ZN(n7941) );
  INV_X1 U7299 ( .A(n6762), .ZN(n5734) );
  INV_X1 U7300 ( .A(n5733), .ZN(n5735) );
  OAI22_X1 U7301 ( .A1(n8041), .A2(n9954), .B1(n9959), .B2(n8042), .ZN(n5736)
         );
  NOR2_X4 U7302 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n5798) );
  NAND4_X1 U7303 ( .A1(n5764), .A2(n6059), .A3(n6125), .A4(n5766), .ZN(n5743)
         );
  INV_X1 U7304 ( .A(n5743), .ZN(n5747) );
  NOR2_X1 U7305 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n5746) );
  NOR2_X1 U7306 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n5745) );
  NOR2_X1 U7307 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n5744) );
  INV_X1 U7308 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n5753) );
  OR2_X1 U7309 ( .A1(n6050), .A2(n5753), .ZN(n5759) );
  OR2_X1 U7310 ( .A1(n8693), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n5758) );
  INV_X1 U7311 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6366) );
  NOR2_X1 U7312 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n5760) );
  INV_X1 U7313 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5762) );
  NAND2_X1 U7314 ( .A1(n6125), .A2(n5762), .ZN(n5763) );
  NAND2_X1 U7315 ( .A1(n4717), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5774) );
  NAND2_X1 U7316 ( .A1(n5774), .A2(n5771), .ZN(n5772) );
  NAND2_X1 U7317 ( .A1(n5772), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5773) );
  XNOR2_X1 U7318 ( .A(n5774), .B(P1_IR_REG_25__SCAN_IN), .ZN(n6288) );
  NAND2_X1 U7319 ( .A1(n5775), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5776) );
  MUX2_X1 U7320 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5776), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n5777) );
  AND2_X1 U7321 ( .A1(n5777), .A2(n4717), .ZN(n6287) );
  AND2_X2 U7322 ( .A1(n6916), .A2(n6315), .ZN(n5845) );
  NAND2_X4 U7323 ( .A1(n5838), .A2(n4478), .ZN(n8869) );
  OR2_X1 U7324 ( .A1(n8869), .A2(n6394), .ZN(n5786) );
  NAND2_X2 U7325 ( .A1(n5838), .A2(n7515), .ZN(n5955) );
  OR2_X1 U7326 ( .A1(n5955), .A2(n6395), .ZN(n5785) );
  NAND2_X1 U7327 ( .A1(n5782), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5783) );
  XNOR2_X1 U7328 ( .A(n5783), .B(n5739), .ZN(n6393) );
  OR2_X1 U7329 ( .A1(n5838), .A2(n6393), .ZN(n5784) );
  NAND2_X1 U7330 ( .A1(n5788), .A2(n5787), .ZN(n5792) );
  NAND2_X1 U7331 ( .A1(n4429), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5791) );
  NAND2_X1 U7332 ( .A1(n6310), .A2(n9321), .ZN(n6828) );
  INV_X1 U7333 ( .A(n6916), .ZN(n6321) );
  NAND2_X1 U7335 ( .A1(n6308), .A2(n6313), .ZN(n6829) );
  INV_X1 U7336 ( .A(n6915), .ZN(n7033) );
  AOI22_X1 U7337 ( .A1(n8689), .A2(n6677), .B1(n5845), .B2(n7033), .ZN(n5862)
         );
  INV_X1 U7338 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n6682) );
  INV_X1 U7339 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6364) );
  OR2_X1 U7340 ( .A1(n6007), .A2(n6364), .ZN(n5796) );
  INV_X1 U7341 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n5793) );
  OR2_X1 U7342 ( .A1(n6162), .A2(n5793), .ZN(n5795) );
  NAND2_X1 U7343 ( .A1(n8814), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5794) );
  NAND2_X1 U7344 ( .A1(n9104), .A2(n5845), .ZN(n5806) );
  OR2_X1 U7345 ( .A1(n8869), .A2(n6392), .ZN(n5804) );
  OR2_X1 U7346 ( .A1(n5955), .A2(n6405), .ZN(n5803) );
  NOR2_X1 U7347 ( .A1(n5798), .A2(n6084), .ZN(n5799) );
  MUX2_X1 U7348 ( .A(n6084), .B(n5799), .S(P1_IR_REG_2__SCAN_IN), .Z(n5800) );
  INV_X1 U7349 ( .A(n5800), .ZN(n5801) );
  NAND2_X1 U7350 ( .A1(n5801), .A2(n5782), .ZN(n6627) );
  OR2_X1 U7351 ( .A1(n5838), .A2(n6627), .ZN(n5802) );
  AND3_X2 U7352 ( .A1(n5804), .A2(n5803), .A3(n5802), .ZN(n9850) );
  NAND2_X1 U7353 ( .A1(n5806), .A2(n5805), .ZN(n5807) );
  XNOR2_X1 U7354 ( .A(n5807), .B(n6260), .ZN(n5808) );
  AOI22_X1 U7355 ( .A1(n8689), .A2(n9104), .B1(n5845), .B2(n7018), .ZN(n5809)
         );
  NAND2_X1 U7356 ( .A1(n5808), .A2(n5809), .ZN(n6725) );
  INV_X1 U7357 ( .A(n5808), .ZN(n5811) );
  INV_X1 U7358 ( .A(n5809), .ZN(n5810) );
  NAND2_X1 U7359 ( .A1(n5811), .A2(n5810), .ZN(n5812) );
  NAND2_X1 U7360 ( .A1(n5868), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5817) );
  INV_X1 U7361 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n7027) );
  INV_X1 U7362 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n5826) );
  OR2_X1 U7363 ( .A1(n6007), .A2(n5826), .ZN(n5815) );
  INV_X1 U7364 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n5813) );
  NAND2_X1 U7365 ( .A1(n8689), .A2(n6440), .ZN(n5823) );
  INV_X1 U7366 ( .A(SI_0_), .ZN(n5819) );
  INV_X1 U7367 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5818) );
  OAI21_X1 U7368 ( .B1(n4478), .B2(n5819), .A(n5818), .ZN(n5821) );
  AND2_X1 U7369 ( .A1(n5821), .A2(n5820), .ZN(n9625) );
  MUX2_X1 U7370 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9625), .S(n5838), .Z(n7030) );
  AOI22_X1 U7371 ( .A1(n5845), .A2(n7030), .B1(n6344), .B2(
        P1_IR_REG_0__SCAN_IN), .ZN(n5822) );
  AND2_X1 U7372 ( .A1(n5823), .A2(n5822), .ZN(n6572) );
  NAND2_X1 U7373 ( .A1(n6440), .A2(n5845), .ZN(n5829) );
  INV_X2 U7374 ( .A(n5824), .ZN(n5825) );
  NOR2_X1 U7375 ( .A1(n6315), .A2(n5826), .ZN(n5827) );
  NAND2_X1 U7376 ( .A1(n5829), .A2(n5828), .ZN(n6571) );
  NAND2_X1 U7377 ( .A1(n6572), .A2(n6571), .ZN(n6570) );
  INV_X1 U7378 ( .A(n6571), .ZN(n5831) );
  NAND2_X1 U7379 ( .A1(n5831), .A2(n5830), .ZN(n5832) );
  NAND2_X1 U7380 ( .A1(n6570), .A2(n5832), .ZN(n5847) );
  INV_X1 U7381 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n5833) );
  NAND2_X1 U7382 ( .A1(n8814), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5834) );
  AND2_X1 U7383 ( .A1(n5835), .A2(n5834), .ZN(n5836) );
  INV_X1 U7384 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n7088) );
  INV_X1 U7385 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6361) );
  NAND2_X1 U7386 ( .A1(n9106), .A2(n5845), .ZN(n5843) );
  OR2_X1 U7387 ( .A1(n5955), .A2(n6406), .ZN(n5840) );
  INV_X1 U7388 ( .A(n5798), .ZN(n5837) );
  OR2_X1 U7389 ( .A1(n5838), .A2(n6391), .ZN(n5839) );
  NAND2_X1 U7390 ( .A1(n5843), .A2(n5842), .ZN(n5844) );
  XNOR2_X1 U7391 ( .A(n5844), .B(n6260), .ZN(n5846) );
  NOR2_X1 U7392 ( .A1(n5847), .A2(n5846), .ZN(n6714) );
  OAI22_X1 U7393 ( .A1(n6825), .A2(n6278), .B1(n9846), .B2(n6279), .ZN(n6715)
         );
  NAND2_X1 U7394 ( .A1(n5847), .A2(n5846), .ZN(n6712) );
  NAND2_X1 U7395 ( .A1(n5868), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5852) );
  INV_X1 U7396 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n5848) );
  OR2_X1 U7397 ( .A1(n6007), .A2(n5848), .ZN(n5851) );
  XNOR2_X1 U7398 ( .A(P1_REG3_REG_3__SCAN_IN), .B(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n7067) );
  OR2_X1 U7399 ( .A1(n8693), .A2(n7067), .ZN(n5850) );
  INV_X1 U7400 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n7068) );
  OR2_X1 U7401 ( .A1(n6050), .A2(n7068), .ZN(n5849) );
  NAND2_X1 U7402 ( .A1(n9103), .A2(n5845), .ZN(n5859) );
  OR2_X1 U7403 ( .A1(n8869), .A2(n6400), .ZN(n5857) );
  OR2_X1 U7404 ( .A1(n5955), .A2(n6399), .ZN(n5856) );
  NAND2_X1 U7405 ( .A1(n5853), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5854) );
  XNOR2_X1 U7406 ( .A(n5854), .B(P1_IR_REG_4__SCAN_IN), .ZN(n9735) );
  INV_X1 U7407 ( .A(n9735), .ZN(n6398) );
  OR2_X1 U7408 ( .A1(n5838), .A2(n6398), .ZN(n5855) );
  OR2_X1 U7409 ( .A1(n5825), .A2(n9855), .ZN(n5858) );
  NAND2_X1 U7410 ( .A1(n5859), .A2(n5858), .ZN(n5860) );
  XNOR2_X1 U7411 ( .A(n5860), .B(n5830), .ZN(n5864) );
  AOI22_X1 U7412 ( .A1(n8689), .A2(n9103), .B1(n5845), .B2(n7074), .ZN(n5865)
         );
  XNOR2_X1 U7413 ( .A(n5864), .B(n5865), .ZN(n6734) );
  INV_X1 U7414 ( .A(n5861), .ZN(n5863) );
  NAND2_X1 U7415 ( .A1(n5863), .A2(n5862), .ZN(n6735) );
  NAND2_X1 U7416 ( .A1(n5868), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5876) );
  INV_X1 U7417 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n5869) );
  OR2_X1 U7418 ( .A1(n6007), .A2(n5869), .ZN(n5875) );
  NAND3_X1 U7419 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n5892) );
  INV_X1 U7420 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5871) );
  NAND2_X1 U7421 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n5870) );
  NAND2_X1 U7422 ( .A1(n5871), .A2(n5870), .ZN(n5872) );
  NAND2_X1 U7423 ( .A1(n5892), .A2(n5872), .ZN(n7181) );
  OR2_X1 U7424 ( .A1(n8693), .A2(n7181), .ZN(n5874) );
  INV_X1 U7425 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n7182) );
  OR2_X1 U7426 ( .A1(n6050), .A2(n7182), .ZN(n5873) );
  NAND4_X1 U7427 ( .A1(n5876), .A2(n5875), .A3(n5874), .A4(n5873), .ZN(n9102)
         );
  NAND2_X1 U7428 ( .A1(n9102), .A2(n5845), .ZN(n5885) );
  OR2_X1 U7429 ( .A1(n5955), .A2(n6403), .ZN(n5883) );
  OR2_X1 U7430 ( .A1(n8869), .A2(n6402), .ZN(n5882) );
  NOR2_X1 U7431 ( .A1(n5877), .A2(n6084), .ZN(n5878) );
  MUX2_X1 U7432 ( .A(n6084), .B(n5878), .S(P1_IR_REG_5__SCAN_IN), .Z(n5880) );
  OR2_X1 U7433 ( .A1(n5880), .A2(n5879), .ZN(n6401) );
  OR2_X1 U7434 ( .A1(n5838), .A2(n6401), .ZN(n5881) );
  OR2_X1 U7435 ( .A1(n5825), .A2(n9863), .ZN(n5884) );
  NAND2_X1 U7436 ( .A1(n5885), .A2(n5884), .ZN(n5886) );
  XNOR2_X1 U7437 ( .A(n5886), .B(n5830), .ZN(n6986) );
  NAND2_X1 U7438 ( .A1(n8689), .A2(n9102), .ZN(n5888) );
  OR2_X1 U7439 ( .A1(n6279), .A2(n9863), .ZN(n5887) );
  NAND2_X1 U7440 ( .A1(n5888), .A2(n5887), .ZN(n5906) );
  NAND2_X1 U7441 ( .A1(n6987), .A2(n5889), .ZN(n5909) );
  NAND2_X1 U7442 ( .A1(n5868), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5897) );
  INV_X1 U7443 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n5890) );
  OR2_X1 U7444 ( .A1(n6007), .A2(n5890), .ZN(n5896) );
  INV_X1 U7445 ( .A(n5892), .ZN(n5891) );
  NAND2_X1 U7446 ( .A1(n5891), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5914) );
  INV_X1 U7447 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6380) );
  NAND2_X1 U7448 ( .A1(n5892), .A2(n6380), .ZN(n5893) );
  NAND2_X1 U7449 ( .A1(n5914), .A2(n5893), .ZN(n7043) );
  OR2_X1 U7450 ( .A1(n8693), .A2(n7043), .ZN(n5895) );
  INV_X1 U7451 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n7044) );
  OR2_X1 U7452 ( .A1(n6050), .A2(n7044), .ZN(n5894) );
  NAND4_X1 U7453 ( .A1(n5897), .A2(n5896), .A3(n5895), .A4(n5894), .ZN(n9101)
         );
  OR2_X1 U7454 ( .A1(n5955), .A2(n6409), .ZN(n5901) );
  OR2_X1 U7455 ( .A1(n8869), .A2(n8574), .ZN(n5900) );
  OR2_X1 U7456 ( .A1(n5879), .A2(n6084), .ZN(n5898) );
  XNOR2_X1 U7457 ( .A(n5898), .B(P1_IR_REG_6__SCAN_IN), .ZN(n6359) );
  INV_X1 U7458 ( .A(n6359), .ZN(n6408) );
  OR2_X1 U7459 ( .A1(n5838), .A2(n6408), .ZN(n5899) );
  AOI22_X1 U7460 ( .A1(n9101), .A2(n5845), .B1(n7133), .B2(n8684), .ZN(n5902)
         );
  XOR2_X1 U7461 ( .A(n5830), .B(n5902), .Z(n5904) );
  INV_X1 U7462 ( .A(n9101), .ZN(n8642) );
  OAI22_X1 U7463 ( .A1(n8642), .A2(n6278), .B1(n9868), .B2(n6279), .ZN(n5903)
         );
  INV_X1 U7464 ( .A(n6986), .ZN(n5907) );
  INV_X1 U7465 ( .A(n5906), .ZN(n7003) );
  NAND2_X1 U7466 ( .A1(n5909), .A2(n5908), .ZN(n6990) );
  INV_X1 U7467 ( .A(n5910), .ZN(n8639) );
  NAND2_X1 U7468 ( .A1(n5868), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5919) );
  INV_X1 U7469 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n5911) );
  OR2_X1 U7470 ( .A1(n6254), .A2(n5911), .ZN(n5918) );
  INV_X1 U7471 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n7139) );
  OR2_X1 U7472 ( .A1(n6050), .A2(n7139), .ZN(n5917) );
  INV_X1 U7473 ( .A(n5914), .ZN(n5912) );
  NAND2_X1 U7474 ( .A1(n5912), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5934) );
  INV_X1 U7475 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5913) );
  NAND2_X1 U7476 ( .A1(n5914), .A2(n5913), .ZN(n5915) );
  NAND2_X1 U7477 ( .A1(n5934), .A2(n5915), .ZN(n8645) );
  OR2_X1 U7478 ( .A1(n4386), .A2(n8645), .ZN(n5916) );
  NAND4_X1 U7479 ( .A1(n5919), .A2(n5918), .A3(n5917), .A4(n5916), .ZN(n9100)
         );
  NAND2_X1 U7480 ( .A1(n9100), .A2(n5845), .ZN(n5926) );
  OR2_X1 U7481 ( .A1(n5955), .A2(n6412), .ZN(n5924) );
  OR2_X1 U7482 ( .A1(n8869), .A2(n6413), .ZN(n5923) );
  NAND2_X1 U7483 ( .A1(n5920), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5921) );
  XNOR2_X1 U7484 ( .A(n5921), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6578) );
  INV_X1 U7485 ( .A(n6578), .ZN(n6411) );
  OR2_X1 U7486 ( .A1(n5838), .A2(n6411), .ZN(n5922) );
  OR2_X1 U7487 ( .A1(n5825), .A2(n9876), .ZN(n5925) );
  NAND2_X1 U7488 ( .A1(n5926), .A2(n5925), .ZN(n5927) );
  XNOR2_X1 U7489 ( .A(n5927), .B(n6260), .ZN(n5929) );
  INV_X1 U7490 ( .A(n9876), .ZN(n8646) );
  AOI22_X1 U7491 ( .A1(n8689), .A2(n9100), .B1(n5845), .B2(n8646), .ZN(n5928)
         );
  NAND2_X1 U7492 ( .A1(n5929), .A2(n5928), .ZN(n5931) );
  OR2_X1 U7493 ( .A1(n5929), .A2(n5928), .ZN(n5930) );
  NAND2_X1 U7494 ( .A1(n5931), .A2(n5930), .ZN(n8638) );
  INV_X1 U7495 ( .A(n5931), .ZN(n5932) );
  NOR2_X2 U7496 ( .A1(n8641), .A2(n5932), .ZN(n5946) );
  NAND2_X1 U7497 ( .A1(n5868), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5939) );
  INV_X1 U7498 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6369) );
  OR2_X1 U7499 ( .A1(n6254), .A2(n6369), .ZN(n5938) );
  INV_X1 U7500 ( .A(n5934), .ZN(n5933) );
  NAND2_X1 U7501 ( .A1(n5933), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5948) );
  INV_X1 U7502 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n8499) );
  NAND2_X1 U7503 ( .A1(n5934), .A2(n8499), .ZN(n5935) );
  NAND2_X1 U7504 ( .A1(n5948), .A2(n5935), .ZN(n7193) );
  OR2_X1 U7505 ( .A1(n8693), .A2(n7193), .ZN(n5937) );
  INV_X1 U7506 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n7167) );
  OR2_X1 U7507 ( .A1(n6050), .A2(n7167), .ZN(n5936) );
  NAND4_X1 U7508 ( .A1(n5939), .A2(n5938), .A3(n5937), .A4(n5936), .ZN(n9099)
         );
  INV_X1 U7509 ( .A(n9099), .ZN(n7236) );
  OR2_X1 U7510 ( .A1(n5955), .A2(n6416), .ZN(n5943) );
  OR2_X1 U7511 ( .A1(n8869), .A2(n6415), .ZN(n5942) );
  NAND2_X1 U7512 ( .A1(n4412), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5940) );
  XNOR2_X1 U7513 ( .A(n5940), .B(P1_IR_REG_8__SCAN_IN), .ZN(n9774) );
  INV_X1 U7514 ( .A(n9774), .ZN(n6414) );
  OR2_X1 U7515 ( .A1(n5838), .A2(n6414), .ZN(n5941) );
  OAI22_X1 U7516 ( .A1(n7236), .A2(n6278), .B1(n9882), .B2(n6279), .ZN(n5945)
         );
  AOI22_X1 U7517 ( .A1(n9099), .A2(n5845), .B1(n7229), .B2(n8684), .ZN(n5944)
         );
  XNOR2_X1 U7518 ( .A(n5944), .B(n5830), .ZN(n7191) );
  NAND2_X1 U7519 ( .A1(n5868), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5953) );
  INV_X1 U7520 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n6370) );
  OR2_X1 U7521 ( .A1(n6007), .A2(n6370), .ZN(n5952) );
  NAND2_X1 U7522 ( .A1(n5948), .A2(n5947), .ZN(n5949) );
  NAND2_X1 U7523 ( .A1(n5971), .A2(n5949), .ZN(n7239) );
  OR2_X1 U7524 ( .A1(n8693), .A2(n7239), .ZN(n5951) );
  INV_X1 U7525 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n6356) );
  OR2_X1 U7526 ( .A1(n6050), .A2(n6356), .ZN(n5950) );
  NAND4_X1 U7527 ( .A1(n5953), .A2(n5952), .A3(n5951), .A4(n5950), .ZN(n9098)
         );
  NAND2_X1 U7528 ( .A1(n9098), .A2(n5845), .ZN(n5959) );
  NAND2_X1 U7529 ( .A1(n5967), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5954) );
  XNOR2_X1 U7530 ( .A(n5954), .B(P1_IR_REG_9__SCAN_IN), .ZN(n6597) );
  INV_X1 U7531 ( .A(n6597), .ZN(n6420) );
  NAND2_X1 U7532 ( .A1(n6418), .A2(n8866), .ZN(n5957) );
  OR2_X1 U7533 ( .A1(n8869), .A2(n6419), .ZN(n5956) );
  OAI211_X1 U7534 ( .C1(n5838), .C2(n6420), .A(n5957), .B(n5956), .ZN(n9891)
         );
  NAND2_X1 U7535 ( .A1(n8684), .A2(n9891), .ZN(n5958) );
  NAND2_X1 U7536 ( .A1(n5959), .A2(n5958), .ZN(n5960) );
  XNOR2_X1 U7537 ( .A(n5960), .B(n6260), .ZN(n5964) );
  NAND2_X1 U7538 ( .A1(n8689), .A2(n9098), .ZN(n5962) );
  NAND2_X1 U7539 ( .A1(n9891), .A2(n5845), .ZN(n5961) );
  AND2_X1 U7540 ( .A1(n5962), .A2(n5961), .ZN(n5963) );
  NAND2_X1 U7541 ( .A1(n5964), .A2(n5963), .ZN(n5965) );
  OAI21_X1 U7542 ( .B1(n5964), .B2(n5963), .A(n5965), .ZN(n7222) );
  INV_X1 U7543 ( .A(n5965), .ZN(n5966) );
  NAND2_X1 U7544 ( .A1(n6427), .A2(n8866), .ZN(n5970) );
  NOR2_X1 U7545 ( .A1(n5967), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n5984) );
  OR2_X1 U7546 ( .A1(n5984), .A2(n6084), .ZN(n5968) );
  XNOR2_X1 U7547 ( .A(n5968), .B(P1_IR_REG_10__SCAN_IN), .ZN(n9779) );
  AOI22_X1 U7548 ( .A1(n6140), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6346), .B2(
        n9779), .ZN(n5969) );
  OR2_X1 U7549 ( .A1(n7380), .A2(n6279), .ZN(n5978) );
  NAND2_X1 U7550 ( .A1(n5868), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5976) );
  INV_X1 U7551 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6595) );
  OR2_X1 U7552 ( .A1(n6254), .A2(n6595), .ZN(n5975) );
  NAND2_X1 U7553 ( .A1(n5971), .A2(n7331), .ZN(n5972) );
  NAND2_X1 U7554 ( .A1(n5991), .A2(n5972), .ZN(n7332) );
  OR2_X1 U7555 ( .A1(n8693), .A2(n7332), .ZN(n5974) );
  INV_X1 U7556 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n6588) );
  OR2_X1 U7557 ( .A1(n6050), .A2(n6588), .ZN(n5973) );
  NAND4_X1 U7558 ( .A1(n5976), .A2(n5975), .A3(n5974), .A4(n5973), .ZN(n9097)
         );
  NAND2_X1 U7559 ( .A1(n8689), .A2(n9097), .ZN(n5977) );
  NAND2_X1 U7560 ( .A1(n5978), .A2(n5977), .ZN(n5981) );
  AOI22_X1 U7561 ( .A1(n7351), .A2(n8684), .B1(n5845), .B2(n9097), .ZN(n5979)
         );
  XNOR2_X1 U7562 ( .A(n5979), .B(n5830), .ZN(n5980) );
  XOR2_X1 U7563 ( .A(n5981), .B(n5980), .Z(n7329) );
  INV_X1 U7564 ( .A(n5980), .ZN(n5982) );
  NOR2_X1 U7565 ( .A1(n5982), .A2(n5981), .ZN(n7388) );
  NAND2_X1 U7566 ( .A1(n6428), .A2(n8866), .ZN(n5987) );
  INV_X1 U7567 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5983) );
  NAND2_X1 U7568 ( .A1(n5984), .A2(n5983), .ZN(n6002) );
  NAND2_X1 U7569 ( .A1(n6002), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5985) );
  XNOR2_X1 U7570 ( .A(n5985), .B(P1_IR_REG_11__SCAN_IN), .ZN(n7267) );
  AOI22_X1 U7571 ( .A1(n6140), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n6346), .B2(
        n7267), .ZN(n5986) );
  NAND2_X1 U7572 ( .A1(n9589), .A2(n8684), .ZN(n5998) );
  NAND2_X1 U7573 ( .A1(n5868), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5996) );
  INV_X1 U7574 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n5988) );
  OR2_X1 U7575 ( .A1(n6254), .A2(n5988), .ZN(n5995) );
  INV_X1 U7576 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5990) );
  NAND2_X1 U7577 ( .A1(n5991), .A2(n5990), .ZN(n5992) );
  NAND2_X1 U7578 ( .A1(n6009), .A2(n5992), .ZN(n7392) );
  OR2_X1 U7579 ( .A1(n4386), .A2(n7392), .ZN(n5994) );
  INV_X1 U7580 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7365) );
  OR2_X1 U7581 ( .A1(n6050), .A2(n7365), .ZN(n5993) );
  NAND4_X1 U7582 ( .A1(n5996), .A2(n5995), .A3(n5994), .A4(n5993), .ZN(n9096)
         );
  NAND2_X1 U7583 ( .A1(n9096), .A2(n5845), .ZN(n5997) );
  NAND2_X1 U7584 ( .A1(n5998), .A2(n5997), .ZN(n5999) );
  XNOR2_X1 U7585 ( .A(n5999), .B(n6260), .ZN(n6001) );
  AOI22_X1 U7586 ( .A1(n9589), .A2(n5845), .B1(n8689), .B2(n9096), .ZN(n6000)
         );
  XNOR2_X1 U7587 ( .A(n6001), .B(n6000), .ZN(n7387) );
  NOR2_X1 U7588 ( .A1(n6001), .A2(n6000), .ZN(n8727) );
  NAND2_X1 U7589 ( .A1(n6443), .A2(n8866), .ZN(n6005) );
  OAI21_X1 U7590 ( .B1(n6002), .B2(P1_IR_REG_11__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6003) );
  XNOR2_X1 U7591 ( .A(n6003), .B(P1_IR_REG_12__SCAN_IN), .ZN(n9115) );
  AOI22_X1 U7592 ( .A1(n6140), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n6346), .B2(
        n9115), .ZN(n6004) );
  NAND2_X2 U7593 ( .A1(n6005), .A2(n6004), .ZN(n9586) );
  NAND2_X1 U7594 ( .A1(n9586), .A2(n8684), .ZN(n6016) );
  NAND2_X1 U7595 ( .A1(n5868), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n6014) );
  INV_X1 U7596 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n6006) );
  OR2_X1 U7597 ( .A1(n6007), .A2(n6006), .ZN(n6013) );
  INV_X1 U7598 ( .A(n6009), .ZN(n6008) );
  NAND2_X1 U7599 ( .A1(n6008), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n6027) );
  INV_X1 U7600 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n8722) );
  NAND2_X1 U7601 ( .A1(n6009), .A2(n8722), .ZN(n6010) );
  NAND2_X1 U7602 ( .A1(n6027), .A2(n6010), .ZN(n8725) );
  OR2_X1 U7603 ( .A1(n8693), .A2(n8725), .ZN(n6012) );
  INV_X1 U7604 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7405) );
  OR2_X1 U7605 ( .A1(n6050), .A2(n7405), .ZN(n6011) );
  OR2_X1 U7606 ( .A1(n7402), .A2(n6279), .ZN(n6015) );
  NAND2_X1 U7607 ( .A1(n6016), .A2(n6015), .ZN(n6017) );
  XNOR2_X1 U7608 ( .A(n6017), .B(n6260), .ZN(n6020) );
  NOR2_X1 U7609 ( .A1(n7402), .A2(n6278), .ZN(n6018) );
  AOI21_X1 U7610 ( .B1(n9586), .B2(n5845), .A(n6018), .ZN(n6019) );
  XNOR2_X1 U7611 ( .A(n6020), .B(n6019), .ZN(n8726) );
  NAND2_X1 U7612 ( .A1(n6020), .A2(n6019), .ZN(n6021) );
  NAND2_X1 U7613 ( .A1(n6452), .A2(n8866), .ZN(n6025) );
  NAND2_X1 U7614 ( .A1(n6022), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6023) );
  XNOR2_X1 U7615 ( .A(n6023), .B(P1_IR_REG_13__SCAN_IN), .ZN(n9128) );
  AOI22_X1 U7616 ( .A1(n6140), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n6346), .B2(
        n9128), .ZN(n6024) );
  NAND2_X1 U7617 ( .A1(n9579), .A2(n8684), .ZN(n6035) );
  NAND2_X1 U7618 ( .A1(n5868), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n6033) );
  INV_X1 U7619 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n7264) );
  OR2_X1 U7620 ( .A1(n6254), .A2(n7264), .ZN(n6032) );
  NAND2_X1 U7621 ( .A1(n6027), .A2(n6026), .ZN(n6028) );
  NAND2_X1 U7622 ( .A1(n6048), .A2(n6028), .ZN(n9476) );
  OR2_X1 U7623 ( .A1(n4386), .A2(n9476), .ZN(n6031) );
  INV_X1 U7624 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n6029) );
  OR2_X1 U7625 ( .A1(n6050), .A2(n6029), .ZN(n6030) );
  NAND4_X1 U7626 ( .A1(n6033), .A2(n6032), .A3(n6031), .A4(n6030), .ZN(n9095)
         );
  NAND2_X1 U7627 ( .A1(n9095), .A2(n5845), .ZN(n6034) );
  NAND2_X1 U7628 ( .A1(n6035), .A2(n6034), .ZN(n6036) );
  XNOR2_X1 U7629 ( .A(n6036), .B(n5830), .ZN(n6042) );
  INV_X1 U7630 ( .A(n6042), .ZN(n6040) );
  NAND2_X1 U7631 ( .A1(n9579), .A2(n5845), .ZN(n6038) );
  NAND2_X1 U7632 ( .A1(n8689), .A2(n9095), .ZN(n6037) );
  NAND2_X1 U7633 ( .A1(n6038), .A2(n6037), .ZN(n6041) );
  INV_X1 U7634 ( .A(n6041), .ZN(n6039) );
  NAND2_X1 U7635 ( .A1(n6040), .A2(n6039), .ZN(n7484) );
  AND2_X1 U7636 ( .A1(n6042), .A2(n6041), .ZN(n7485) );
  NAND2_X1 U7637 ( .A1(n6456), .A2(n8866), .ZN(n6045) );
  OR2_X1 U7638 ( .A1(n6043), .A2(n6084), .ZN(n6057) );
  XNOR2_X1 U7639 ( .A(n6057), .B(P1_IR_REG_14__SCAN_IN), .ZN(n9796) );
  AOI22_X1 U7640 ( .A1(n6140), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n6346), .B2(
        n9796), .ZN(n6044) );
  NAND2_X1 U7641 ( .A1(n5868), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n6054) );
  INV_X1 U7642 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n6046) );
  OR2_X1 U7643 ( .A1(n6254), .A2(n6046), .ZN(n6053) );
  INV_X1 U7644 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n8655) );
  NAND2_X1 U7645 ( .A1(n6048), .A2(n8655), .ZN(n6049) );
  NAND2_X1 U7646 ( .A1(n6065), .A2(n6049), .ZN(n8658) );
  OR2_X1 U7647 ( .A1(n8693), .A2(n8658), .ZN(n6052) );
  INV_X1 U7648 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7466) );
  OR2_X1 U7649 ( .A1(n6050), .A2(n7466), .ZN(n6051) );
  NAND4_X1 U7650 ( .A1(n6054), .A2(n6053), .A3(n6052), .A4(n6051), .ZN(n9485)
         );
  OAI22_X1 U7651 ( .A1(n4758), .A2(n5825), .B1(n9200), .B2(n6279), .ZN(n6055)
         );
  XOR2_X1 U7652 ( .A(n5830), .B(n6055), .Z(n6077) );
  NAND2_X1 U7653 ( .A1(n6076), .A2(n6077), .ZN(n8652) );
  OAI22_X1 U7654 ( .A1(n4758), .A2(n6279), .B1(n9200), .B2(n6278), .ZN(n8654)
         );
  NAND2_X1 U7655 ( .A1(n8652), .A2(n8654), .ZN(n6080) );
  NAND2_X1 U7656 ( .A1(n6652), .A2(n8866), .ZN(n6063) );
  INV_X1 U7657 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n6056) );
  NAND2_X1 U7658 ( .A1(n6057), .A2(n6056), .ZN(n6058) );
  NAND2_X1 U7659 ( .A1(n6058), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6060) );
  XNOR2_X1 U7660 ( .A(n6060), .B(n6059), .ZN(n9141) );
  INV_X1 U7661 ( .A(n9141), .ZN(n6061) );
  AOI22_X1 U7662 ( .A1(n6140), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n6346), .B2(
        n6061), .ZN(n6062) );
  NAND2_X1 U7663 ( .A1(n9574), .A2(n8684), .ZN(n6074) );
  NAND2_X1 U7664 ( .A1(n5868), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n6072) );
  NAND2_X1 U7665 ( .A1(n6065), .A2(n6064), .ZN(n6066) );
  NAND2_X1 U7666 ( .A1(n6090), .A2(n6066), .ZN(n9461) );
  OR2_X1 U7667 ( .A1(n4386), .A2(n9461), .ZN(n6071) );
  INV_X1 U7668 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n6067) );
  OR2_X1 U7669 ( .A1(n6254), .A2(n6067), .ZN(n6070) );
  INV_X1 U7670 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n6068) );
  OR2_X1 U7671 ( .A1(n6050), .A2(n6068), .ZN(n6069) );
  NAND4_X1 U7672 ( .A1(n6072), .A2(n6071), .A3(n6070), .A4(n6069), .ZN(n9452)
         );
  NAND2_X1 U7673 ( .A1(n9452), .A2(n5845), .ZN(n6073) );
  NAND2_X1 U7674 ( .A1(n6074), .A2(n6073), .ZN(n6075) );
  XNOR2_X1 U7675 ( .A(n6075), .B(n6260), .ZN(n6081) );
  INV_X1 U7676 ( .A(n6076), .ZN(n6079) );
  INV_X1 U7677 ( .A(n6077), .ZN(n6078) );
  NAND2_X1 U7678 ( .A1(n6079), .A2(n6078), .ZN(n8651) );
  NAND3_X1 U7679 ( .A1(n6080), .A2(n6081), .A3(n8651), .ZN(n8793) );
  INV_X1 U7680 ( .A(n9452), .ZN(n9201) );
  OAI22_X1 U7681 ( .A1(n9464), .A2(n6279), .B1(n9201), .B2(n6278), .ZN(n8796)
         );
  NAND2_X1 U7682 ( .A1(n6080), .A2(n8651), .ZN(n6083) );
  INV_X1 U7683 ( .A(n6081), .ZN(n6082) );
  NAND2_X1 U7684 ( .A1(n6656), .A2(n8866), .ZN(n6088) );
  OR2_X1 U7685 ( .A1(n6085), .A2(n6084), .ZN(n6086) );
  XNOR2_X1 U7686 ( .A(n6086), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9160) );
  AOI22_X1 U7687 ( .A1(n6140), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n6346), .B2(
        n9160), .ZN(n6087) );
  NAND2_X1 U7688 ( .A1(n5868), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n6095) );
  INV_X1 U7689 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n8487) );
  OR2_X1 U7690 ( .A1(n6254), .A2(n8487), .ZN(n6094) );
  INV_X1 U7691 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n7559) );
  NAND2_X1 U7692 ( .A1(n6090), .A2(n7559), .ZN(n6091) );
  NAND2_X1 U7693 ( .A1(n6102), .A2(n6091), .ZN(n7558) );
  OR2_X1 U7694 ( .A1(n4386), .A2(n7558), .ZN(n6093) );
  INV_X1 U7695 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n9136) );
  OR2_X1 U7696 ( .A1(n6050), .A2(n9136), .ZN(n6092) );
  AOI22_X1 U7697 ( .A1(n9570), .A2(n8684), .B1(n5845), .B2(n9467), .ZN(n6096)
         );
  XNOR2_X1 U7698 ( .A(n6096), .B(n5830), .ZN(n6113) );
  AOI22_X1 U7699 ( .A1(n9570), .A2(n5845), .B1(n8689), .B2(n9467), .ZN(n6112)
         );
  XNOR2_X1 U7700 ( .A(n6113), .B(n6112), .ZN(n7557) );
  NAND2_X1 U7701 ( .A1(n6709), .A2(n8866), .ZN(n6099) );
  NAND2_X1 U7702 ( .A1(n6097), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6126) );
  XNOR2_X1 U7703 ( .A(n6126), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9175) );
  AOI22_X1 U7704 ( .A1(n6140), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n6346), .B2(
        n9175), .ZN(n6098) );
  INV_X1 U7705 ( .A(n9564), .ZN(n9433) );
  NAND2_X1 U7706 ( .A1(n8814), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n6108) );
  INV_X1 U7707 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n6100) );
  OR2_X1 U7708 ( .A1(n6254), .A2(n6100), .ZN(n6107) );
  INV_X1 U7709 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n6101) );
  NAND2_X1 U7710 ( .A1(n6102), .A2(n6101), .ZN(n6103) );
  NAND2_X1 U7711 ( .A1(n6133), .A2(n6103), .ZN(n9430) );
  OR2_X1 U7712 ( .A1(n8693), .A2(n9430), .ZN(n6106) );
  INV_X1 U7713 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n6104) );
  OR2_X1 U7714 ( .A1(n6162), .A2(n6104), .ZN(n6105) );
  NAND4_X1 U7715 ( .A1(n6108), .A2(n6107), .A3(n6106), .A4(n6105), .ZN(n9453)
         );
  OAI22_X1 U7716 ( .A1(n9433), .A2(n6279), .B1(n9423), .B2(n6278), .ZN(n6118)
         );
  NAND2_X1 U7717 ( .A1(n9564), .A2(n8684), .ZN(n6110) );
  NAND2_X1 U7718 ( .A1(n9453), .A2(n5845), .ZN(n6109) );
  NAND2_X1 U7719 ( .A1(n6110), .A2(n6109), .ZN(n6111) );
  XNOR2_X1 U7720 ( .A(n6111), .B(n5830), .ZN(n6117) );
  XOR2_X1 U7721 ( .A(n6118), .B(n6117), .Z(n8746) );
  INV_X1 U7722 ( .A(n8746), .ZN(n6116) );
  INV_X1 U7723 ( .A(n6112), .ZN(n6115) );
  INV_X1 U7724 ( .A(n6113), .ZN(n6114) );
  OR2_X1 U7725 ( .A1(n6115), .A2(n6114), .ZN(n8744) );
  OR2_X1 U7726 ( .A1(n6116), .A2(n8744), .ZN(n6122) );
  INV_X1 U7727 ( .A(n6117), .ZN(n6120) );
  INV_X1 U7728 ( .A(n6118), .ZN(n6119) );
  NAND2_X1 U7729 ( .A1(n6120), .A2(n6119), .ZN(n6121) );
  AND2_X1 U7730 ( .A1(n6122), .A2(n6121), .ZN(n6123) );
  NAND2_X1 U7731 ( .A1(n6124), .A2(n6123), .ZN(n7539) );
  NAND2_X1 U7732 ( .A1(n6806), .A2(n8866), .ZN(n6130) );
  NAND2_X1 U7733 ( .A1(n6126), .A2(n6125), .ZN(n6127) );
  NAND2_X1 U7734 ( .A1(n6127), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6128) );
  XNOR2_X1 U7735 ( .A(n6128), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9814) );
  AOI22_X1 U7736 ( .A1(n6140), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n6346), .B2(
        n9814), .ZN(n6129) );
  INV_X1 U7737 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n8508) );
  OR2_X1 U7738 ( .A1(n6162), .A2(n8508), .ZN(n6138) );
  INV_X1 U7739 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9173) );
  OR2_X1 U7740 ( .A1(n6254), .A2(n9173), .ZN(n6137) );
  INV_X1 U7741 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n6132) );
  NAND2_X1 U7742 ( .A1(n6133), .A2(n6132), .ZN(n6134) );
  NAND2_X1 U7743 ( .A1(n6146), .A2(n6134), .ZN(n9408) );
  OR2_X1 U7744 ( .A1(n8693), .A2(n9408), .ZN(n6136) );
  INV_X1 U7745 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9409) );
  OR2_X1 U7746 ( .A1(n6050), .A2(n9409), .ZN(n6135) );
  OAI22_X1 U7747 ( .A1(n9406), .A2(n5825), .B1(n9204), .B2(n6279), .ZN(n6139)
         );
  XOR2_X1 U7748 ( .A(n5830), .B(n6139), .Z(n7541) );
  AOI22_X1 U7749 ( .A1(n9561), .A2(n5845), .B1(n8689), .B2(n9436), .ZN(n7540)
         );
  NAND2_X1 U7750 ( .A1(n6877), .A2(n8866), .ZN(n6142) );
  AOI22_X1 U7751 ( .A1(n6140), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9356), .B2(
        n6346), .ZN(n6141) );
  NAND2_X1 U7752 ( .A1(n8694), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n6151) );
  INV_X1 U7753 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n6143) );
  OR2_X1 U7754 ( .A1(n6050), .A2(n6143), .ZN(n6150) );
  INV_X1 U7755 ( .A(n6146), .ZN(n6144) );
  INV_X1 U7756 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n6145) );
  NAND2_X1 U7757 ( .A1(n6146), .A2(n6145), .ZN(n6147) );
  NAND2_X1 U7758 ( .A1(n6159), .A2(n6147), .ZN(n9389) );
  OR2_X1 U7759 ( .A1(n8693), .A2(n9389), .ZN(n6149) );
  INV_X1 U7760 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n8489) );
  OR2_X1 U7761 ( .A1(n6446), .A2(n8489), .ZN(n6148) );
  OAI22_X1 U7762 ( .A1(n9392), .A2(n5825), .B1(n9421), .B2(n6279), .ZN(n6152)
         );
  XNOR2_X1 U7763 ( .A(n6152), .B(n5830), .ZN(n8671) );
  OR2_X1 U7764 ( .A1(n9392), .A2(n6279), .ZN(n6154) );
  OR2_X1 U7765 ( .A1(n9421), .A2(n6278), .ZN(n6153) );
  NAND2_X1 U7766 ( .A1(n6154), .A2(n6153), .ZN(n8672) );
  NAND2_X1 U7767 ( .A1(n8671), .A2(n8672), .ZN(n6156) );
  NAND2_X1 U7768 ( .A1(n6998), .A2(n8866), .ZN(n6158) );
  OR2_X1 U7769 ( .A1(n8869), .A2(n6999), .ZN(n6157) );
  INV_X1 U7770 ( .A(n9551), .ZN(n9374) );
  NAND2_X1 U7771 ( .A1(n8694), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n6166) );
  INV_X1 U7772 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n9376) );
  OR2_X1 U7773 ( .A1(n6050), .A2(n9376), .ZN(n6165) );
  INV_X1 U7774 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n8763) );
  NAND2_X1 U7775 ( .A1(n6159), .A2(n8763), .ZN(n6160) );
  NAND2_X1 U7776 ( .A1(n6174), .A2(n6160), .ZN(n9375) );
  OR2_X1 U7777 ( .A1(n4386), .A2(n9375), .ZN(n6164) );
  INV_X1 U7778 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n6161) );
  OR2_X1 U7779 ( .A1(n6162), .A2(n6161), .ZN(n6163) );
  NAND4_X1 U7780 ( .A1(n6166), .A2(n6165), .A3(n6164), .A4(n6163), .ZN(n9396)
         );
  OAI22_X1 U7781 ( .A1(n9374), .A2(n5825), .B1(n9207), .B2(n6279), .ZN(n6167)
         );
  XOR2_X1 U7782 ( .A(n5830), .B(n6167), .Z(n6169) );
  AOI22_X1 U7783 ( .A1(n9551), .A2(n5845), .B1(n8689), .B2(n9396), .ZN(n6168)
         );
  NAND2_X1 U7784 ( .A1(n6169), .A2(n6168), .ZN(n6170) );
  OAI21_X1 U7785 ( .B1(n6169), .B2(n6168), .A(n6170), .ZN(n8762) );
  NAND2_X1 U7786 ( .A1(n7115), .A2(n8866), .ZN(n6172) );
  OR2_X1 U7787 ( .A1(n8869), .A2(n7116), .ZN(n6171) );
  INV_X1 U7788 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n6173) );
  NAND2_X1 U7789 ( .A1(n6174), .A2(n6173), .ZN(n6175) );
  AND2_X1 U7790 ( .A1(n6192), .A2(n6175), .ZN(n9362) );
  NAND2_X1 U7791 ( .A1(n6276), .A2(n9362), .ZN(n6179) );
  INV_X1 U7792 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n8554) );
  OR2_X1 U7793 ( .A1(n6446), .A2(n8554), .ZN(n6178) );
  INV_X1 U7794 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n8492) );
  OR2_X1 U7795 ( .A1(n6254), .A2(n8492), .ZN(n6177) );
  INV_X1 U7796 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n8426) );
  OR2_X1 U7797 ( .A1(n6050), .A2(n8426), .ZN(n6176) );
  OAI22_X1 U7798 ( .A1(n9355), .A2(n6279), .B1(n9382), .B2(n6278), .ZN(n6184)
         );
  NAND2_X1 U7799 ( .A1(n9368), .A2(n8684), .ZN(n6181) );
  OR2_X1 U7800 ( .A1(n9382), .A2(n6279), .ZN(n6180) );
  NAND2_X1 U7801 ( .A1(n6181), .A2(n6180), .ZN(n6182) );
  XNOR2_X1 U7802 ( .A(n6182), .B(n5830), .ZN(n6183) );
  XOR2_X1 U7803 ( .A(n6184), .B(n6183), .Z(n8715) );
  INV_X1 U7804 ( .A(n6183), .ZN(n6186) );
  INV_X1 U7805 ( .A(n6184), .ZN(n6185) );
  NAND2_X1 U7806 ( .A1(n6186), .A2(n6185), .ZN(n6187) );
  NAND2_X1 U7807 ( .A1(n8714), .A2(n6187), .ZN(n6200) );
  NAND2_X1 U7808 ( .A1(n7201), .A2(n8866), .ZN(n6189) );
  OR2_X1 U7809 ( .A1(n8869), .A2(n7204), .ZN(n6188) );
  INV_X1 U7810 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n6198) );
  INV_X1 U7811 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n6191) );
  NAND2_X1 U7812 ( .A1(n6192), .A2(n6191), .ZN(n6193) );
  NAND2_X1 U7813 ( .A1(n6208), .A2(n6193), .ZN(n9343) );
  OR2_X1 U7814 ( .A1(n9343), .A2(n8693), .ZN(n6197) );
  NAND2_X1 U7815 ( .A1(n8694), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n6195) );
  NAND2_X1 U7816 ( .A1(n8814), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n6194) );
  AND2_X1 U7817 ( .A1(n6195), .A2(n6194), .ZN(n6196) );
  OAI211_X1 U7818 ( .C1(n6446), .C2(n6198), .A(n6197), .B(n6196), .ZN(n9358)
         );
  AOI22_X1 U7819 ( .A1(n9539), .A2(n5845), .B1(n8689), .B2(n9358), .ZN(n6201)
         );
  NAND2_X1 U7820 ( .A1(n6200), .A2(n6201), .ZN(n8769) );
  OAI22_X1 U7821 ( .A1(n9346), .A2(n5825), .B1(n9210), .B2(n6279), .ZN(n6199)
         );
  XNOR2_X1 U7822 ( .A(n6199), .B(n5830), .ZN(n8772) );
  NAND2_X1 U7823 ( .A1(n8769), .A2(n8772), .ZN(n6214) );
  NAND2_X1 U7824 ( .A1(n7273), .A2(n8866), .ZN(n6205) );
  OR2_X1 U7825 ( .A1(n8869), .A2(n7276), .ZN(n6204) );
  INV_X1 U7826 ( .A(n6208), .ZN(n6206) );
  NAND2_X1 U7827 ( .A1(n6206), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n6220) );
  INV_X1 U7828 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n6207) );
  NAND2_X1 U7829 ( .A1(n6208), .A2(n6207), .ZN(n6209) );
  NAND2_X1 U7830 ( .A1(n6220), .A2(n6209), .ZN(n9330) );
  OR2_X1 U7831 ( .A1(n9330), .A2(n4386), .ZN(n6212) );
  AOI22_X1 U7832 ( .A1(n8694), .A2(P1_REG1_REG_23__SCAN_IN), .B1(n5868), .B2(
        P1_REG0_REG_23__SCAN_IN), .ZN(n6211) );
  NAND2_X1 U7833 ( .A1(n8814), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n6210) );
  OAI22_X1 U7834 ( .A1(n9333), .A2(n5825), .B1(n9212), .B2(n6279), .ZN(n6213)
         );
  XNOR2_X1 U7835 ( .A(n6213), .B(n6260), .ZN(n6215) );
  OAI22_X1 U7836 ( .A1(n9333), .A2(n6279), .B1(n9212), .B2(n6278), .ZN(n8665)
         );
  INV_X1 U7837 ( .A(n6215), .ZN(n6216) );
  NAND2_X1 U7838 ( .A1(n7297), .A2(n8866), .ZN(n6218) );
  OR2_X1 U7839 ( .A1(n8869), .A2(n8411), .ZN(n6217) );
  INV_X1 U7840 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n6219) );
  NAND2_X1 U7841 ( .A1(n6220), .A2(n6219), .ZN(n6221) );
  AND2_X1 U7842 ( .A1(n6237), .A2(n6221), .ZN(n9320) );
  NAND2_X1 U7843 ( .A1(n9320), .A2(n6276), .ZN(n6226) );
  INV_X1 U7844 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n8412) );
  NAND2_X1 U7845 ( .A1(n8694), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n6223) );
  INV_X1 U7846 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n8581) );
  OR2_X1 U7847 ( .A1(n6446), .A2(n8581), .ZN(n6222) );
  OAI211_X1 U7848 ( .C1(n8412), .C2(n6050), .A(n6223), .B(n6222), .ZN(n6224)
         );
  INV_X1 U7849 ( .A(n6224), .ZN(n6225) );
  OAI22_X1 U7850 ( .A1(n9312), .A2(n5825), .B1(n9214), .B2(n6279), .ZN(n6227)
         );
  XNOR2_X1 U7851 ( .A(n6227), .B(n6260), .ZN(n6231) );
  OR2_X1 U7852 ( .A1(n9312), .A2(n6279), .ZN(n6229) );
  NAND2_X1 U7853 ( .A1(n9336), .A2(n8689), .ZN(n6228) );
  NAND2_X1 U7854 ( .A1(n6231), .A2(n6230), .ZN(n6232) );
  OAI21_X1 U7855 ( .B1(n6231), .B2(n6230), .A(n6232), .ZN(n8755) );
  NAND2_X1 U7856 ( .A1(n7431), .A2(n8866), .ZN(n6234) );
  OR2_X1 U7857 ( .A1(n8869), .A2(n7434), .ZN(n6233) );
  INV_X1 U7858 ( .A(n6237), .ZN(n6235) );
  NAND2_X1 U7859 ( .A1(n6235), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n6250) );
  INV_X1 U7860 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n6236) );
  NAND2_X1 U7861 ( .A1(n6237), .A2(n6236), .ZN(n6238) );
  NAND2_X1 U7862 ( .A1(n6250), .A2(n6238), .ZN(n8738) );
  OR2_X1 U7863 ( .A1(n8738), .A2(n8693), .ZN(n6244) );
  INV_X1 U7864 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n6241) );
  NAND2_X1 U7865 ( .A1(n8814), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n6240) );
  NAND2_X1 U7866 ( .A1(n5868), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n6239) );
  OAI211_X1 U7867 ( .C1(n6254), .C2(n6241), .A(n6240), .B(n6239), .ZN(n6242)
         );
  INV_X1 U7868 ( .A(n6242), .ZN(n6243) );
  OAI22_X1 U7869 ( .A1(n9302), .A2(n6279), .B1(n9288), .B2(n6278), .ZN(n6263)
         );
  NAND2_X1 U7870 ( .A1(n9524), .A2(n8684), .ZN(n6246) );
  NAND2_X1 U7871 ( .A1(n9316), .A2(n5845), .ZN(n6245) );
  NAND2_X1 U7872 ( .A1(n6246), .A2(n6245), .ZN(n6247) );
  XNOR2_X1 U7873 ( .A(n6247), .B(n5830), .ZN(n6264) );
  XOR2_X1 U7874 ( .A(n6263), .B(n6264), .Z(n8736) );
  NAND2_X1 U7875 ( .A1(n7438), .A2(n8866), .ZN(n6249) );
  OR2_X1 U7876 ( .A1(n8869), .A2(n7439), .ZN(n6248) );
  NAND2_X1 U7877 ( .A1(n9521), .A2(n8684), .ZN(n6259) );
  INV_X1 U7878 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n8785) );
  NAND2_X1 U7879 ( .A1(n6250), .A2(n8785), .ZN(n6251) );
  NAND2_X1 U7880 ( .A1(n9292), .A2(n6276), .ZN(n6257) );
  INV_X1 U7881 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n8506) );
  NAND2_X1 U7882 ( .A1(n8814), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n6253) );
  INV_X1 U7883 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n8592) );
  OR2_X1 U7884 ( .A1(n6446), .A2(n8592), .ZN(n6252) );
  OAI211_X1 U7885 ( .C1(n6254), .C2(n8506), .A(n6253), .B(n6252), .ZN(n6255)
         );
  INV_X1 U7886 ( .A(n6255), .ZN(n6256) );
  NAND2_X1 U7887 ( .A1(n9306), .A2(n5845), .ZN(n6258) );
  NAND2_X1 U7888 ( .A1(n6259), .A2(n6258), .ZN(n6261) );
  XNOR2_X1 U7889 ( .A(n6261), .B(n6260), .ZN(n6266) );
  AND2_X1 U7890 ( .A1(n9306), .A2(n8689), .ZN(n6262) );
  AOI21_X1 U7891 ( .B1(n9521), .B2(n5845), .A(n6262), .ZN(n6267) );
  XNOR2_X1 U7892 ( .A(n6266), .B(n6267), .ZN(n8780) );
  NOR2_X1 U7893 ( .A1(n6264), .A2(n6263), .ZN(n8781) );
  NOR2_X1 U7894 ( .A1(n8780), .A2(n8781), .ZN(n6265) );
  INV_X1 U7895 ( .A(n6266), .ZN(n6269) );
  INV_X1 U7896 ( .A(n6267), .ZN(n6268) );
  NAND2_X1 U7897 ( .A1(n6269), .A2(n6268), .ZN(n6283) );
  NAND2_X1 U7898 ( .A1(n7508), .A2(n8866), .ZN(n6271) );
  OR2_X1 U7899 ( .A1(n8869), .A2(n8476), .ZN(n6270) );
  XNOR2_X1 U7900 ( .A(n6326), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n9274) );
  INV_X1 U7901 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n6274) );
  NAND2_X1 U7902 ( .A1(n8694), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n6273) );
  NAND2_X1 U7903 ( .A1(n5868), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n6272) );
  OAI211_X1 U7904 ( .C1(n6050), .C2(n6274), .A(n6273), .B(n6272), .ZN(n6275)
         );
  AOI21_X2 U7905 ( .B1(n9274), .B2(n6276), .A(n6275), .ZN(n9289) );
  OAI22_X1 U7906 ( .A1(n9276), .A2(n5825), .B1(n9289), .B2(n6279), .ZN(n6277)
         );
  XNOR2_X1 U7907 ( .A(n6277), .B(n5830), .ZN(n6281) );
  OAI22_X1 U7908 ( .A1(n9276), .A2(n6279), .B1(n9289), .B2(n6278), .ZN(n6280)
         );
  NOR2_X1 U7909 ( .A1(n6281), .A2(n6280), .ZN(n8704) );
  AOI21_X1 U7910 ( .B1(n6281), .B2(n6280), .A(n8704), .ZN(n6282) );
  AOI21_X1 U7911 ( .B1(n6286), .B2(n6283), .A(n6282), .ZN(n6311) );
  INV_X1 U7912 ( .A(n6282), .ZN(n6285) );
  INV_X1 U7913 ( .A(n6283), .ZN(n6284) );
  INV_X1 U7914 ( .A(n6288), .ZN(n7432) );
  NAND3_X1 U7915 ( .A1(n7432), .A2(P1_B_REG_SCAN_IN), .A3(n7298), .ZN(n6289)
         );
  OR2_X1 U7916 ( .A1(n9829), .A2(P1_D_REG_0__SCAN_IN), .ZN(n6292) );
  INV_X1 U7917 ( .A(n6290), .ZN(n7440) );
  NAND2_X1 U7918 ( .A1(n7440), .A2(n7298), .ZN(n6291) );
  NOR4_X1 U7919 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_17__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n8392) );
  NOR2_X1 U7920 ( .A1(P1_D_REG_30__SCAN_IN), .A2(P1_D_REG_31__SCAN_IN), .ZN(
        n6295) );
  NOR4_X1 U7921 ( .A1(P1_D_REG_5__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_6__SCAN_IN), .ZN(n6294) );
  NOR4_X1 U7922 ( .A1(P1_D_REG_24__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_25__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n6293) );
  NAND4_X1 U7923 ( .A1(n8392), .A2(n6295), .A3(n6294), .A4(n6293), .ZN(n6301)
         );
  NOR4_X1 U7924 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), .A3(
        P1_D_REG_14__SCAN_IN), .A4(P1_D_REG_15__SCAN_IN), .ZN(n6299) );
  NOR4_X1 U7925 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_8__SCAN_IN), .A3(
        P1_D_REG_10__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n6298) );
  NOR4_X1 U7926 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_29__SCAN_IN), .A3(
        P1_D_REG_26__SCAN_IN), .A4(P1_D_REG_28__SCAN_IN), .ZN(n6297) );
  NOR4_X1 U7927 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .A3(
        P1_D_REG_23__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n6296) );
  NAND4_X1 U7928 ( .A1(n6299), .A2(n6298), .A3(n6297), .A4(n6296), .ZN(n6300)
         );
  NOR2_X1 U7929 ( .A1(n6301), .A2(n6300), .ZN(n6302) );
  OR2_X1 U7930 ( .A1(n9829), .A2(n6302), .ZN(n6646) );
  NAND2_X1 U7931 ( .A1(n9616), .A2(n6646), .ZN(n6639) );
  OR2_X1 U7932 ( .A1(n9829), .A2(P1_D_REG_1__SCAN_IN), .ZN(n6304) );
  NAND2_X1 U7933 ( .A1(n7440), .A2(n7432), .ZN(n6303) );
  NOR2_X1 U7934 ( .A1(n6639), .A2(n6907), .ZN(n6312) );
  NAND2_X1 U7935 ( .A1(n4468), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6306) );
  AND2_X1 U7936 ( .A1(n7274), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6307) );
  NAND2_X1 U7937 ( .A1(n6312), .A2(n9841), .ZN(n6320) );
  INV_X1 U7938 ( .A(n6910), .ZN(n6641) );
  INV_X1 U7939 ( .A(n9043), .ZN(n6832) );
  OAI21_X1 U7940 ( .B1(n6311), .B2(n8692), .A(n8783), .ZN(n6341) );
  INV_X1 U7941 ( .A(n6312), .ZN(n6569) );
  NOR2_X1 U7942 ( .A1(n6910), .A2(n7000), .ZN(n6912) );
  NAND2_X1 U7943 ( .A1(n6569), .A2(n6912), .ZN(n8712) );
  OR2_X1 U7944 ( .A1(n9043), .A2(n6313), .ZN(n6316) );
  NOR2_X1 U7945 ( .A1(n9881), .A2(n8710), .ZN(n6314) );
  NAND3_X1 U7946 ( .A1(n6316), .A2(n6315), .A3(n7274), .ZN(n6317) );
  AOI21_X1 U7947 ( .B1(n9881), .B2(n6569), .A(n6317), .ZN(n6318) );
  NAND2_X1 U7948 ( .A1(n8712), .A2(n6318), .ZN(n6319) );
  INV_X1 U7949 ( .A(n9306), .ZN(n8859) );
  INV_X1 U7950 ( .A(n6320), .ZN(n6322) );
  OR2_X1 U7951 ( .A1(n6321), .A2(n6828), .ZN(n7009) );
  AND2_X1 U7952 ( .A1(n6322), .A2(n9088), .ZN(n6335) );
  NAND2_X1 U7953 ( .A1(n6335), .A2(n9087), .ZN(n8798) );
  INV_X1 U7954 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n6325) );
  OAI22_X1 U7955 ( .A1(n8859), .A2(n8798), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6325), .ZN(n6337) );
  INV_X1 U7956 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n6324) );
  OAI21_X1 U7957 ( .B1(n6326), .B2(n6325), .A(n6324), .ZN(n6329) );
  INV_X1 U7958 ( .A(n6326), .ZN(n6328) );
  AND2_X1 U7959 ( .A1(P1_REG3_REG_28__SCAN_IN), .A2(P1_REG3_REG_27__SCAN_IN), 
        .ZN(n6327) );
  NAND2_X1 U7960 ( .A1(n6328), .A2(n6327), .ZN(n9220) );
  NAND2_X1 U7961 ( .A1(n6329), .A2(n9220), .ZN(n8700) );
  OR2_X1 U7962 ( .A1(n8700), .A2(n4386), .ZN(n6334) );
  INV_X1 U7963 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n8474) );
  NAND2_X1 U7964 ( .A1(n8694), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n6331) );
  NAND2_X1 U7965 ( .A1(n8814), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n6330) );
  OAI211_X1 U7966 ( .C1(n6446), .C2(n8474), .A(n6331), .B(n6330), .ZN(n6332)
         );
  INV_X1 U7967 ( .A(n6332), .ZN(n6333) );
  NOR2_X1 U7968 ( .A1(n9217), .A2(n8786), .ZN(n6336) );
  AOI211_X1 U7969 ( .C1(n9274), .C2(n8789), .A(n6337), .B(n6336), .ZN(n6338)
         );
  INV_X1 U7970 ( .A(n6339), .ZN(n6340) );
  NAND2_X1 U7971 ( .A1(n6341), .A2(n6340), .ZN(P1_U3212) );
  INV_X2 U7972 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  INV_X1 U7973 ( .A(n7274), .ZN(n6343) );
  OR2_X1 U7974 ( .A1(n9043), .A2(n6343), .ZN(n6345) );
  NAND2_X1 U7975 ( .A1(n6344), .A2(n7274), .ZN(n6376) );
  NAND2_X1 U7976 ( .A1(n6345), .A2(n6376), .ZN(n9728) );
  OAI21_X1 U7977 ( .B1(n9728), .B2(n6346), .A(P1_STATE_REG_SCAN_IN), .ZN(
        P1_U3083) );
  AND2_X1 U7978 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7224) );
  NOR2_X1 U7979 ( .A1(n9774), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6347) );
  AOI21_X1 U7980 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n9774), .A(n6347), .ZN(
        n9760) );
  NOR2_X1 U7981 ( .A1(P1_REG2_REG_7__SCAN_IN), .A2(n6578), .ZN(n6348) );
  AOI21_X1 U7982 ( .B1(n6578), .B2(P1_REG2_REG_7__SCAN_IN), .A(n6348), .ZN(
        n6577) );
  XNOR2_X1 U7983 ( .A(n6401), .B(n7182), .ZN(n9749) );
  INV_X1 U7984 ( .A(n6393), .ZN(n9628) );
  INV_X1 U7985 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6349) );
  NAND2_X1 U7986 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n6631) );
  INV_X1 U7987 ( .A(n6631), .ZN(n9722) );
  NAND2_X1 U7988 ( .A1(n6607), .A2(n9722), .ZN(n6606) );
  INV_X1 U7989 ( .A(n6391), .ZN(n6615) );
  NAND2_X1 U7990 ( .A1(n6615), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6350) );
  NAND2_X1 U7991 ( .A1(n6606), .A2(n6350), .ZN(n6624) );
  INV_X1 U7992 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n8350) );
  OR2_X1 U7993 ( .A1(n6627), .A2(n8350), .ZN(n6352) );
  NAND2_X1 U7994 ( .A1(n6627), .A2(n8350), .ZN(n6351) );
  AND2_X1 U7995 ( .A1(n6352), .A2(n6351), .ZN(n6625) );
  XNOR2_X1 U7996 ( .A(n6393), .B(P1_REG2_REG_3__SCAN_IN), .ZN(n9627) );
  NOR2_X1 U7997 ( .A1(n9735), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6353) );
  AOI21_X1 U7998 ( .B1(n9735), .B2(P1_REG2_REG_4__SCAN_IN), .A(n6353), .ZN(
        n9734) );
  NAND2_X1 U7999 ( .A1(n4415), .A2(n9734), .ZN(n9733) );
  OAI21_X1 U8000 ( .B1(n9735), .B2(P1_REG2_REG_4__SCAN_IN), .A(n9733), .ZN(
        n6354) );
  INV_X1 U8001 ( .A(n6354), .ZN(n9748) );
  INV_X1 U8002 ( .A(n6401), .ZN(n9746) );
  NAND2_X1 U8003 ( .A1(n6359), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6355) );
  OAI21_X1 U8004 ( .B1(n6359), .B2(P1_REG2_REG_6__SCAN_IN), .A(n6355), .ZN(
        n6383) );
  OAI21_X1 U8005 ( .B1(P1_REG2_REG_7__SCAN_IN), .B2(n6578), .A(n6575), .ZN(
        n9759) );
  NAND2_X1 U8006 ( .A1(n9760), .A2(n9759), .ZN(n9758) );
  OAI21_X1 U8007 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n9774), .A(n9758), .ZN(
        n6358) );
  MUX2_X1 U8008 ( .A(n6356), .B(P1_REG2_REG_9__SCAN_IN), .S(n6597), .Z(n6357)
         );
  NOR2_X1 U8009 ( .A1(n6358), .A2(n6357), .ZN(n6589) );
  NOR2_X1 U8010 ( .A1(n9728), .A2(P1_U3084), .ZN(n6373) );
  INV_X1 U8011 ( .A(n9723), .ZN(n9188) );
  NAND2_X1 U8012 ( .A1(n6373), .A2(n9188), .ZN(n6375) );
  AOI211_X1 U8013 ( .C1(n6358), .C2(n6357), .A(n6589), .B(n9819), .ZN(n6379)
         );
  AOI22_X1 U8014 ( .A1(n6359), .A2(n5890), .B1(P1_REG1_REG_6__SCAN_IN), .B2(
        n6408), .ZN(n6386) );
  NAND2_X1 U8015 ( .A1(n9746), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6367) );
  INV_X1 U8016 ( .A(n6367), .ZN(n6360) );
  AOI21_X1 U8017 ( .B1(n5869), .B2(n6401), .A(n6360), .ZN(n9753) );
  AOI22_X1 U8018 ( .A1(n9735), .A2(n5848), .B1(P1_REG1_REG_4__SCAN_IN), .B2(
        n6398), .ZN(n9738) );
  MUX2_X1 U8019 ( .A(n6364), .B(P1_REG1_REG_2__SCAN_IN), .S(n6627), .Z(n6363)
         );
  MUX2_X1 U8020 ( .A(n6361), .B(P1_REG1_REG_1__SCAN_IN), .S(n6391), .Z(n6610)
         );
  AND2_X1 U8021 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n6611) );
  NAND2_X1 U8022 ( .A1(n6610), .A2(n6611), .ZN(n6617) );
  NAND2_X1 U8023 ( .A1(n6615), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6618) );
  NAND2_X1 U8024 ( .A1(n6617), .A2(n6618), .ZN(n6362) );
  NAND2_X1 U8025 ( .A1(n6363), .A2(n6362), .ZN(n9631) );
  OR2_X1 U8026 ( .A1(n6627), .A2(n6364), .ZN(n9630) );
  MUX2_X1 U8027 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n6366), .S(n6393), .Z(n9629)
         );
  AOI21_X1 U8028 ( .B1(n9631), .B2(n9630), .A(n9629), .ZN(n9633) );
  INV_X1 U8029 ( .A(n9633), .ZN(n6365) );
  OAI21_X1 U8030 ( .B1(n6366), .B2(n6393), .A(n6365), .ZN(n9739) );
  NOR2_X1 U8031 ( .A1(n9738), .A2(n9739), .ZN(n9737) );
  AOI21_X1 U8032 ( .B1(n6398), .B2(n5848), .A(n9737), .ZN(n9752) );
  NAND2_X1 U8033 ( .A1(n9753), .A2(n9752), .ZN(n9751) );
  NAND2_X1 U8034 ( .A1(n6367), .A2(n9751), .ZN(n6385) );
  NOR2_X1 U8035 ( .A1(n6386), .A2(n6385), .ZN(n6384) );
  AOI21_X1 U8036 ( .B1(n6408), .B2(n5890), .A(n6384), .ZN(n6582) );
  AOI22_X1 U8037 ( .A1(P1_REG1_REG_7__SCAN_IN), .A2(n6411), .B1(n6578), .B2(
        n5911), .ZN(n6581) );
  NOR2_X1 U8038 ( .A1(n6582), .A2(n6581), .ZN(n6580) );
  NOR2_X1 U8039 ( .A1(n6578), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6368) );
  OR2_X1 U8040 ( .A1(n6580), .A2(n6368), .ZN(n9770) );
  INV_X1 U8041 ( .A(n9770), .ZN(n9761) );
  NOR2_X1 U8042 ( .A1(n6414), .A2(n6369), .ZN(n9762) );
  NAND2_X1 U8043 ( .A1(n6414), .A2(n6369), .ZN(n9766) );
  OAI21_X1 U8044 ( .B1(n9761), .B2(n9762), .A(n9766), .ZN(n9767) );
  MUX2_X1 U8045 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n6370), .S(n6597), .Z(n6371)
         );
  NAND2_X1 U8046 ( .A1(n6371), .A2(n9767), .ZN(n6596) );
  OAI21_X1 U8047 ( .B1(n9767), .B2(n6371), .A(n6596), .ZN(n6374) );
  NOR2_X1 U8048 ( .A1(n9726), .A2(n9188), .ZN(n6372) );
  NAND2_X1 U8049 ( .A1(n6373), .A2(n6372), .ZN(n9769) );
  INV_X1 U8050 ( .A(n9769), .ZN(n9824) );
  AND2_X1 U8051 ( .A1(n6374), .A2(n9824), .ZN(n6378) );
  INV_X1 U8052 ( .A(n6375), .ZN(n9171) );
  INV_X1 U8053 ( .A(n9815), .ZN(n9149) );
  INV_X1 U8054 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10181) );
  INV_X1 U8055 ( .A(n6376), .ZN(n6635) );
  OAI22_X1 U8056 ( .A1(n9149), .A2(n6420), .B1(n10181), .B2(n9828), .ZN(n6377)
         );
  OR4_X1 U8057 ( .A1(n7224), .A2(n6379), .A3(n6378), .A4(n6377), .ZN(P1_U3250)
         );
  NOR2_X1 U8058 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6380), .ZN(n6994) );
  AOI211_X1 U8059 ( .C1(n6383), .C2(n6382), .A(n6381), .B(n9819), .ZN(n6390)
         );
  AOI21_X1 U8060 ( .B1(n6386), .B2(n6385), .A(n6384), .ZN(n6387) );
  NOR2_X1 U8061 ( .A1(n9769), .A2(n6387), .ZN(n6389) );
  OAI22_X1 U8062 ( .A1(n9149), .A2(n6408), .B1(n9678), .B2(n9828), .ZN(n6388)
         );
  OR4_X1 U8063 ( .A1(n6994), .A2(n6390), .A3(n6389), .A4(n6388), .ZN(P1_U3247)
         );
  AND2_X1 U8064 ( .A1(n4478), .A2(P1_U3084), .ZN(n6710) );
  INV_X2 U8065 ( .A(n6710), .ZN(n9618) );
  NOR2_X1 U8066 ( .A1(n4478), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9622) );
  OAI222_X1 U8067 ( .A1(n9618), .A2(n4551), .B1(n7433), .B2(n6406), .C1(
        P1_U3084), .C2(n6391), .ZN(P1_U3352) );
  OAI222_X1 U8068 ( .A1(n9618), .A2(n6392), .B1(n7433), .B2(n6405), .C1(
        P1_U3084), .C2(n6627), .ZN(P1_U3351) );
  OAI222_X1 U8069 ( .A1(n9618), .A2(n6394), .B1(n7433), .B2(n6395), .C1(
        P1_U3084), .C2(n6393), .ZN(P1_U3350) );
  AND2_X1 U8070 ( .A1(n7515), .A2(P2_U3152), .ZN(n8633) );
  INV_X2 U8071 ( .A(n8633), .ZN(n8627) );
  NAND2_X1 U8072 ( .A1(n4478), .A2(P2_U3152), .ZN(n8635) );
  INV_X1 U8073 ( .A(n6479), .ZN(n6546) );
  OAI222_X1 U8074 ( .A1(n8627), .A2(n6396), .B1(n8635), .B2(n6395), .C1(
        P2_U3152), .C2(n6546), .ZN(P2_U3355) );
  INV_X1 U8075 ( .A(n6477), .ZN(n6557) );
  OAI222_X1 U8076 ( .A1(n8627), .A2(n6397), .B1(n8635), .B2(n6399), .C1(
        P2_U3152), .C2(n6557), .ZN(P2_U3354) );
  OAI222_X1 U8077 ( .A1(n9618), .A2(n6400), .B1(n7433), .B2(n6399), .C1(
        P1_U3084), .C2(n6398), .ZN(P1_U3349) );
  OAI222_X1 U8078 ( .A1(n9618), .A2(n6402), .B1(n7433), .B2(n6403), .C1(
        P1_U3084), .C2(n6401), .ZN(P1_U3348) );
  OAI222_X1 U8079 ( .A1(n8627), .A2(n8436), .B1(n8635), .B2(n6403), .C1(
        P2_U3152), .C2(n6503), .ZN(P2_U3353) );
  INV_X1 U8080 ( .A(n8635), .ZN(n8630) );
  INV_X1 U8081 ( .A(n8630), .ZN(n7538) );
  AOI22_X1 U8082 ( .A1(n8633), .A2(P1_DATAO_REG_2__SCAN_IN), .B1(n9658), .B2(
        P2_STATE_REG_SCAN_IN), .ZN(n6404) );
  OAI21_X1 U8083 ( .B1(n6405), .B2(n7538), .A(n6404), .ZN(P2_U3356) );
  OAI222_X1 U8084 ( .A1(n8627), .A2(n8590), .B1(n7538), .B2(n6406), .C1(
        P2_U3152), .C2(n6482), .ZN(P2_U3357) );
  INV_X1 U8085 ( .A(n6505), .ZN(n6514) );
  OAI222_X1 U8086 ( .A1(n8627), .A2(n6407), .B1(n8635), .B2(n6409), .C1(
        P2_U3152), .C2(n6514), .ZN(P2_U3352) );
  OAI222_X1 U8087 ( .A1(n9618), .A2(n8574), .B1(n7433), .B2(n6409), .C1(
        P1_U3084), .C2(n6408), .ZN(P1_U3347) );
  INV_X1 U8088 ( .A(n6511), .ZN(n6568) );
  OAI222_X1 U8089 ( .A1(n8627), .A2(n6410), .B1(n8635), .B2(n6412), .C1(
        P2_U3152), .C2(n6568), .ZN(P2_U3351) );
  OAI222_X1 U8090 ( .A1(n9618), .A2(n6413), .B1(n7433), .B2(n6412), .C1(
        P1_U3084), .C2(n6411), .ZN(P1_U3346) );
  OAI222_X1 U8091 ( .A1(n9618), .A2(n6415), .B1(n7433), .B2(n6416), .C1(
        P1_U3084), .C2(n6414), .ZN(P1_U3345) );
  INV_X1 U8092 ( .A(n6528), .ZN(n6521) );
  OAI222_X1 U8093 ( .A1(n8627), .A2(n6417), .B1(n8635), .B2(n6416), .C1(
        P2_U3152), .C2(n6521), .ZN(P2_U3350) );
  INV_X1 U8094 ( .A(n6418), .ZN(n6421) );
  OAI222_X1 U8095 ( .A1(n7433), .A2(n6421), .B1(n6420), .B2(P1_U3084), .C1(
        n6419), .C2(n9618), .ZN(P1_U3344) );
  INV_X1 U8096 ( .A(n6662), .ZN(n6536) );
  OAI222_X1 U8097 ( .A1(n8627), .A2(n6422), .B1(n8635), .B2(n6421), .C1(n6536), 
        .C2(P2_U3152), .ZN(P2_U3349) );
  NAND2_X1 U8098 ( .A1(n7943), .A2(n6762), .ZN(n6426) );
  OR2_X1 U8099 ( .A1(n6423), .A2(P2_U3152), .ZN(n7946) );
  NAND2_X1 U8100 ( .A1(n10037), .A2(n7946), .ZN(n6424) );
  NAND2_X1 U8101 ( .A1(n6424), .A2(n4387), .ZN(n6425) );
  NOR2_X1 U8102 ( .A1(n9969), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U8103 ( .A(n7968), .ZN(n6659) );
  INV_X1 U8104 ( .A(n6427), .ZN(n6436) );
  OAI222_X1 U8105 ( .A1(P2_U3152), .A2(n6659), .B1(n7538), .B2(n6436), .C1(
        n8552), .C2(n8627), .ZN(P2_U3348) );
  INV_X1 U8106 ( .A(n6428), .ZN(n6438) );
  INV_X1 U8107 ( .A(n7267), .ZN(n6598) );
  OAI222_X1 U8108 ( .A1(n7433), .A2(n6438), .B1(n6598), .B2(P1_U3084), .C1(
        n6429), .C2(n9618), .ZN(P1_U3342) );
  INV_X1 U8109 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n6435) );
  INV_X1 U8110 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n6433) );
  INV_X1 U8111 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n8023) );
  OR2_X1 U8112 ( .A1(n6430), .A2(n8023), .ZN(n6432) );
  NAND2_X1 U8113 ( .A1(n7593), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n6431) );
  OAI211_X1 U8114 ( .C1(n7598), .C2(n6433), .A(n6432), .B(n6431), .ZN(n8025)
         );
  NAND2_X1 U8115 ( .A1(n8025), .A2(P2_U3966), .ZN(n6434) );
  OAI21_X1 U8116 ( .B1(n6435), .B2(P2_U3966), .A(n6434), .ZN(P2_U3583) );
  INV_X1 U8117 ( .A(n9779), .ZN(n6437) );
  OAI222_X1 U8118 ( .A1(n9618), .A2(n8588), .B1(n6437), .B2(P1_U3084), .C1(
        n7433), .C2(n6436), .ZN(P1_U3343) );
  INV_X1 U8119 ( .A(n6684), .ZN(n6690) );
  OAI222_X1 U8120 ( .A1(n8627), .A2(n6439), .B1(n7538), .B2(n6438), .C1(n6690), 
        .C2(P2_U3152), .ZN(P2_U3347) );
  INV_X1 U8121 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n6442) );
  NAND2_X1 U8122 ( .A1(n6440), .A2(P1_U4006), .ZN(n6441) );
  OAI21_X1 U8123 ( .B1(P1_U4006), .B2(n6442), .A(n6441), .ZN(P1_U3555) );
  INV_X1 U8124 ( .A(n6443), .ZN(n6445) );
  INV_X1 U8125 ( .A(n9115), .ZN(n7265) );
  OAI222_X1 U8126 ( .A1(n9618), .A2(n6444), .B1(n7433), .B2(n6445), .C1(
        P1_U3084), .C2(n7265), .ZN(P1_U3341) );
  INV_X1 U8127 ( .A(n6815), .ZN(n6698) );
  OAI222_X1 U8128 ( .A1(n8627), .A2(n8556), .B1(n7538), .B2(n6445), .C1(
        P2_U3152), .C2(n6698), .ZN(P2_U3346) );
  INV_X1 U8129 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6451) );
  INV_X1 U8130 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n6449) );
  NAND2_X1 U8131 ( .A1(n8814), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6448) );
  INV_X1 U8132 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n8576) );
  OR2_X1 U8133 ( .A1(n6446), .A2(n8576), .ZN(n6447) );
  OAI211_X1 U8134 ( .C1(n6254), .C2(n6449), .A(n6448), .B(n6447), .ZN(n9190)
         );
  NAND2_X1 U8135 ( .A1(n9190), .A2(P1_U4006), .ZN(n6450) );
  OAI21_X1 U8136 ( .B1(P1_U4006), .B2(n6451), .A(n6450), .ZN(P1_U3586) );
  INV_X1 U8137 ( .A(n6452), .ZN(n6454) );
  AOI22_X1 U8138 ( .A1(n9128), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n6710), .ZN(n6453) );
  OAI21_X1 U8139 ( .B1(n6454), .B2(n7433), .A(n6453), .ZN(P1_U3340) );
  INV_X1 U8140 ( .A(n6866), .ZN(n6861) );
  OAI222_X1 U8141 ( .A1(n8627), .A2(n6455), .B1(n7538), .B2(n6454), .C1(n6861), 
        .C2(P2_U3152), .ZN(P2_U3345) );
  INV_X1 U8142 ( .A(n6456), .ZN(n6459) );
  INV_X1 U8143 ( .A(n9796), .ZN(n7263) );
  OAI222_X1 U8144 ( .A1(n7433), .A2(n6459), .B1(n7263), .B2(P1_U3084), .C1(
        n6457), .C2(n9618), .ZN(P1_U3339) );
  INV_X1 U8145 ( .A(n7248), .ZN(n6871) );
  OAI222_X1 U8146 ( .A1(P2_U3152), .A2(n6871), .B1(n7538), .B2(n6459), .C1(
        n6458), .C2(n8627), .ZN(P2_U3344) );
  NOR2_X1 U8147 ( .A1(n5733), .A2(P2_U3152), .ZN(n8632) );
  NAND2_X1 U8148 ( .A1(n6460), .A2(n8632), .ZN(n6461) );
  OAI211_X1 U8149 ( .C1(n10037), .C2(n6762), .A(n7946), .B(n6461), .ZN(n6463)
         );
  NAND2_X1 U8150 ( .A1(n6463), .A2(n6462), .ZN(n6471) );
  NAND2_X1 U8151 ( .A1(n6471), .A2(n7967), .ZN(n6488) );
  NAND2_X1 U8152 ( .A1(n6488), .A2(n5733), .ZN(n9971) );
  NOR2_X1 U8153 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6802), .ZN(n6476) );
  XNOR2_X1 U8154 ( .A(n6503), .B(n6464), .ZN(n6494) );
  NAND2_X1 U8155 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n9645) );
  INV_X1 U8156 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6465) );
  MUX2_X1 U8157 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n6465), .S(n6482), .Z(n9644)
         );
  INV_X1 U8158 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6466) );
  NAND2_X1 U8159 ( .A1(n6479), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6467) );
  OAI21_X1 U8160 ( .B1(n6479), .B2(P2_REG1_REG_3__SCAN_IN), .A(n6467), .ZN(
        n6538) );
  NOR2_X1 U8161 ( .A1(n6539), .A2(n6538), .ZN(n6537) );
  AOI21_X1 U8162 ( .B1(n6479), .B2(P2_REG1_REG_3__SCAN_IN), .A(n6537), .ZN(
        n6549) );
  MUX2_X1 U8163 ( .A(n6468), .B(P2_REG1_REG_4__SCAN_IN), .S(n6477), .Z(n6548)
         );
  NOR2_X1 U8164 ( .A1(n6549), .A2(n6548), .ZN(n6547) );
  AOI21_X1 U8165 ( .B1(n6477), .B2(P2_REG1_REG_4__SCAN_IN), .A(n6547), .ZN(
        n6495) );
  NOR2_X1 U8166 ( .A1(n6494), .A2(n6495), .ZN(n6493) );
  INV_X1 U8167 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6470) );
  MUX2_X1 U8168 ( .A(n6470), .B(P2_REG1_REG_6__SCAN_IN), .S(n6505), .Z(n6473)
         );
  INV_X1 U8169 ( .A(n6471), .ZN(n6472) );
  AOI211_X1 U8170 ( .C1(n6474), .C2(n6473), .A(n6504), .B(n9972), .ZN(n6475)
         );
  AOI211_X1 U8171 ( .C1(P2_ADDR_REG_6__SCAN_IN), .C2(n9969), .A(n6476), .B(
        n6475), .ZN(n6492) );
  NAND2_X1 U8172 ( .A1(P2_REG2_REG_4__SCAN_IN), .A2(n6477), .ZN(n6485) );
  MUX2_X1 U8173 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n6478), .S(n6477), .Z(n6553)
         );
  NAND2_X1 U8174 ( .A1(n6479), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6484) );
  MUX2_X1 U8175 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n6480), .S(n6479), .Z(n6542)
         );
  NAND2_X1 U8176 ( .A1(P2_REG2_REG_2__SCAN_IN), .A2(n9658), .ZN(n6483) );
  MUX2_X1 U8177 ( .A(n6981), .B(P2_REG2_REG_2__SCAN_IN), .S(n9658), .Z(n6481)
         );
  INV_X1 U8178 ( .A(n6481), .ZN(n9661) );
  MUX2_X1 U8179 ( .A(n5040), .B(P2_REG2_REG_1__SCAN_IN), .S(n6482), .Z(n9649)
         );
  NAND3_X1 U8180 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .A3(n9649), .ZN(n9648) );
  OAI21_X1 U8181 ( .B1(n6482), .B2(n5040), .A(n9648), .ZN(n9662) );
  NAND2_X1 U8182 ( .A1(n9661), .A2(n9662), .ZN(n9660) );
  NAND2_X1 U8183 ( .A1(n6483), .A2(n9660), .ZN(n6543) );
  NAND2_X1 U8184 ( .A1(n6542), .A2(n6543), .ZN(n6541) );
  NAND2_X1 U8185 ( .A1(n6484), .A2(n6541), .ZN(n6554) );
  NAND2_X1 U8186 ( .A1(n6553), .A2(n6554), .ZN(n6552) );
  NAND2_X1 U8187 ( .A1(n6485), .A2(n6552), .ZN(n6500) );
  MUX2_X1 U8188 ( .A(n6886), .B(P2_REG2_REG_5__SCAN_IN), .S(n6503), .Z(n6499)
         );
  NAND2_X1 U8189 ( .A1(n6500), .A2(n6499), .ZN(n6498) );
  OAI21_X1 U8190 ( .B1(n6886), .B2(n6503), .A(n6498), .ZN(n6490) );
  MUX2_X1 U8191 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n6486), .S(n6505), .Z(n6489)
         );
  NOR2_X1 U8192 ( .A1(n5733), .A2(n7599), .ZN(n6487) );
  NAND2_X1 U8193 ( .A1(n6489), .A2(n6490), .ZN(n6513) );
  OAI211_X1 U8194 ( .C1(n6490), .C2(n6489), .A(n9968), .B(n6513), .ZN(n6491)
         );
  OAI211_X1 U8195 ( .C1(n9971), .C2(n6514), .A(n6492), .B(n6491), .ZN(P2_U3251) );
  INV_X1 U8196 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n8579) );
  NOR2_X1 U8197 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8579), .ZN(n6497) );
  AOI211_X1 U8198 ( .C1(n6495), .C2(n6494), .A(n6493), .B(n9972), .ZN(n6496)
         );
  AOI211_X1 U8199 ( .C1(P2_ADDR_REG_5__SCAN_IN), .C2(n9969), .A(n6497), .B(
        n6496), .ZN(n6502) );
  OAI211_X1 U8200 ( .C1(n6500), .C2(n6499), .A(n9968), .B(n6498), .ZN(n6501)
         );
  OAI211_X1 U8201 ( .C1(n9971), .C2(n6503), .A(n6502), .B(n6501), .ZN(P2_U3250) );
  NOR2_X1 U8202 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6899), .ZN(n6510) );
  INV_X1 U8203 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6506) );
  MUX2_X1 U8204 ( .A(n6506), .B(P2_REG1_REG_7__SCAN_IN), .S(n6511), .Z(n6559)
         );
  AOI21_X1 U8205 ( .B1(n6511), .B2(P2_REG1_REG_7__SCAN_IN), .A(n6558), .ZN(
        n6508) );
  INV_X1 U8206 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n8362) );
  MUX2_X1 U8207 ( .A(n8362), .B(P2_REG1_REG_8__SCAN_IN), .S(n6528), .Z(n6507)
         );
  NOR2_X1 U8208 ( .A1(n6508), .A2(n6507), .ZN(n6522) );
  AOI211_X1 U8209 ( .C1(n6508), .C2(n6507), .A(n6522), .B(n9972), .ZN(n6509)
         );
  AOI211_X1 U8210 ( .C1(P2_ADDR_REG_8__SCAN_IN), .C2(n9969), .A(n6510), .B(
        n6509), .ZN(n6520) );
  NAND2_X1 U8211 ( .A1(n6511), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6515) );
  MUX2_X1 U8212 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n6512), .S(n6511), .Z(n6565)
         );
  OAI21_X1 U8213 ( .B1(n6514), .B2(n6486), .A(n6513), .ZN(n6564) );
  NAND2_X1 U8214 ( .A1(n6565), .A2(n6564), .ZN(n6563) );
  NAND2_X1 U8215 ( .A1(n6515), .A2(n6563), .ZN(n6518) );
  MUX2_X1 U8216 ( .A(n10003), .B(P2_REG2_REG_8__SCAN_IN), .S(n6528), .Z(n6516)
         );
  INV_X1 U8217 ( .A(n6516), .ZN(n6517) );
  NAND2_X1 U8218 ( .A1(n6517), .A2(n6518), .ZN(n6529) );
  OAI211_X1 U8219 ( .C1(n6518), .C2(n6517), .A(n9968), .B(n6529), .ZN(n6519)
         );
  OAI211_X1 U8220 ( .C1(n9971), .C2(n6521), .A(n6520), .B(n6519), .ZN(P2_U3253) );
  INV_X1 U8221 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n8407) );
  NOR2_X1 U8222 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8407), .ZN(n6527) );
  AOI21_X1 U8223 ( .B1(n6528), .B2(P2_REG1_REG_8__SCAN_IN), .A(n6522), .ZN(
        n6525) );
  INV_X1 U8224 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n6523) );
  MUX2_X1 U8225 ( .A(n6523), .B(P2_REG1_REG_9__SCAN_IN), .S(n6662), .Z(n6524)
         );
  NOR2_X1 U8226 ( .A1(n6525), .A2(n6524), .ZN(n6663) );
  AOI211_X1 U8227 ( .C1(n6525), .C2(n6524), .A(n6663), .B(n9972), .ZN(n6526)
         );
  AOI211_X1 U8228 ( .C1(P2_ADDR_REG_9__SCAN_IN), .C2(n9969), .A(n6527), .B(
        n6526), .ZN(n6535) );
  NAND2_X1 U8229 ( .A1(n6528), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n6530) );
  NAND2_X1 U8230 ( .A1(n6530), .A2(n6529), .ZN(n6533) );
  MUX2_X1 U8231 ( .A(n7109), .B(P2_REG2_REG_9__SCAN_IN), .S(n6662), .Z(n6531)
         );
  INV_X1 U8232 ( .A(n6531), .ZN(n6532) );
  NAND2_X1 U8233 ( .A1(n6532), .A2(n6533), .ZN(n6657) );
  OAI211_X1 U8234 ( .C1(n6533), .C2(n6532), .A(n9968), .B(n6657), .ZN(n6534)
         );
  OAI211_X1 U8235 ( .C1(n9971), .C2(n6536), .A(n6535), .B(n6534), .ZN(P2_U3254) );
  INV_X1 U8236 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n8468) );
  NOR2_X1 U8237 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8468), .ZN(n9926) );
  AOI211_X1 U8238 ( .C1(n6539), .C2(n6538), .A(n6537), .B(n9972), .ZN(n6540)
         );
  AOI211_X1 U8239 ( .C1(P2_ADDR_REG_3__SCAN_IN), .C2(n9969), .A(n9926), .B(
        n6540), .ZN(n6545) );
  OAI211_X1 U8240 ( .C1(n6543), .C2(n6542), .A(n9968), .B(n6541), .ZN(n6544)
         );
  OAI211_X1 U8241 ( .C1(n9971), .C2(n6546), .A(n6545), .B(n6544), .ZN(P2_U3248) );
  AND2_X1 U8242 ( .A1(P2_U3152), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n6551) );
  AOI211_X1 U8243 ( .C1(n6549), .C2(n6548), .A(n6547), .B(n9972), .ZN(n6550)
         );
  AOI211_X1 U8244 ( .C1(P2_ADDR_REG_4__SCAN_IN), .C2(n9969), .A(n6551), .B(
        n6550), .ZN(n6556) );
  OAI211_X1 U8245 ( .C1(n6554), .C2(n6553), .A(n9968), .B(n6552), .ZN(n6555)
         );
  OAI211_X1 U8246 ( .C1(n9971), .C2(n6557), .A(n6556), .B(n6555), .ZN(P2_U3249) );
  AND2_X1 U8247 ( .A1(P2_U3152), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6562) );
  AOI211_X1 U8248 ( .C1(n6560), .C2(n6559), .A(n6558), .B(n9972), .ZN(n6561)
         );
  AOI211_X1 U8249 ( .C1(P2_ADDR_REG_7__SCAN_IN), .C2(n9969), .A(n6562), .B(
        n6561), .ZN(n6567) );
  OAI211_X1 U8250 ( .C1(n6565), .C2(n6564), .A(n9968), .B(n6563), .ZN(n6566)
         );
  OAI211_X1 U8251 ( .C1(n9971), .C2(n6568), .A(n6567), .B(n6566), .ZN(P2_U3252) );
  OAI21_X1 U8252 ( .B1(n6569), .B2(n8710), .A(n8792), .ZN(n6718) );
  OAI21_X1 U8253 ( .B1(n6572), .B2(n6571), .A(n6570), .ZN(n6630) );
  INV_X1 U8254 ( .A(n7030), .ZN(n7087) );
  OAI22_X1 U8255 ( .A1(n8792), .A2(n7087), .B1(n8786), .B2(n6825), .ZN(n6573)
         );
  AOI21_X1 U8256 ( .B1(n8783), .B2(n6630), .A(n6573), .ZN(n6574) );
  OAI21_X1 U8257 ( .B1(n7027), .B2(n6718), .A(n6574), .ZN(P1_U3230) );
  OAI21_X1 U8258 ( .B1(n6577), .B2(n6576), .A(n6575), .ZN(n6579) );
  AOI22_X1 U8259 ( .A1(n9765), .A2(n6579), .B1(n9815), .B2(n6578), .ZN(n6587)
         );
  AOI21_X1 U8260 ( .B1(n6582), .B2(n6581), .A(n6580), .ZN(n6584) );
  NOR2_X1 U8261 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n5913), .ZN(n8644) );
  INV_X1 U8262 ( .A(n8644), .ZN(n6583) );
  OAI21_X1 U8263 ( .B1(n9769), .B2(n6584), .A(n6583), .ZN(n6585) );
  INV_X1 U8264 ( .A(n6585), .ZN(n6586) );
  OAI211_X1 U8265 ( .C1(n9682), .C2(n9828), .A(n6587), .B(n6586), .ZN(P1_U3248) );
  INV_X1 U8266 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n6604) );
  XNOR2_X1 U8267 ( .A(n9779), .B(n6588), .ZN(n9784) );
  NAND2_X1 U8268 ( .A1(n6597), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6591) );
  INV_X1 U8269 ( .A(n6589), .ZN(n6590) );
  AND2_X1 U8270 ( .A1(n9779), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6592) );
  AOI22_X1 U8271 ( .A1(P1_REG2_REG_11__SCAN_IN), .A2(n7267), .B1(n6598), .B2(
        n7365), .ZN(n6593) );
  OAI21_X1 U8272 ( .B1(n4467), .B2(n6593), .A(n7257), .ZN(n6594) );
  AOI22_X1 U8273 ( .A1(n9765), .A2(n6594), .B1(n9815), .B2(n7267), .ZN(n6603)
         );
  MUX2_X1 U8274 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n6595), .S(n9779), .Z(n9781)
         );
  OAI21_X1 U8275 ( .B1(n6597), .B2(P1_REG1_REG_9__SCAN_IN), .A(n6596), .ZN(
        n9782) );
  NAND2_X1 U8276 ( .A1(n9781), .A2(n9782), .ZN(n9780) );
  OAI21_X1 U8277 ( .B1(n9779), .B2(P1_REG1_REG_10__SCAN_IN), .A(n9780), .ZN(
        n6600) );
  AOI22_X1 U8278 ( .A1(P1_REG1_REG_11__SCAN_IN), .A2(n7267), .B1(n6598), .B2(
        n5988), .ZN(n6599) );
  NAND2_X1 U8279 ( .A1(n6599), .A2(n6600), .ZN(n7266) );
  OAI21_X1 U8280 ( .B1(n6600), .B2(n6599), .A(n7266), .ZN(n6601) );
  NOR2_X1 U8281 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n5990), .ZN(n7391) );
  AOI21_X1 U8282 ( .B1(n9824), .B2(n6601), .A(n7391), .ZN(n6602) );
  OAI211_X1 U8283 ( .C1(n9828), .C2(n6604), .A(n6603), .B(n6602), .ZN(P1_U3252) );
  NAND2_X1 U8284 ( .A1(n9105), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n6605) );
  OAI21_X1 U8285 ( .B1(n9289), .B2(n9105), .A(n6605), .ZN(P1_U3582) );
  OAI21_X1 U8286 ( .B1(n6607), .B2(n9722), .A(n6606), .ZN(n6609) );
  INV_X1 U8287 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n6608) );
  OAI22_X1 U8288 ( .A1(n9819), .A2(n6609), .B1(n9828), .B2(n6608), .ZN(n6614)
         );
  OAI211_X1 U8289 ( .C1(n6611), .C2(n6610), .A(n9824), .B(n6617), .ZN(n6612)
         );
  OAI21_X1 U8290 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n7088), .A(n6612), .ZN(n6613) );
  AOI211_X1 U8291 ( .C1(n9815), .C2(n6615), .A(n6614), .B(n6613), .ZN(n6616)
         );
  INV_X1 U8292 ( .A(n6616), .ZN(P1_U3242) );
  INV_X1 U8293 ( .A(n6617), .ZN(n6621) );
  MUX2_X1 U8294 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n6364), .S(n6627), .Z(n6619)
         );
  NAND2_X1 U8295 ( .A1(n6619), .A2(n6618), .ZN(n6620) );
  OAI211_X1 U8296 ( .C1(n6621), .C2(n6620), .A(n9824), .B(n9631), .ZN(n6622)
         );
  OAI21_X1 U8297 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n6682), .A(n6622), .ZN(n6629) );
  OAI21_X1 U8298 ( .B1(n6625), .B2(n6624), .A(n6623), .ZN(n6626) );
  OAI22_X1 U8299 ( .A1(n9149), .A2(n6627), .B1(n9819), .B2(n6626), .ZN(n6628)
         );
  AOI211_X1 U8300 ( .C1(n9778), .C2(P1_ADDR_REG_2__SCAN_IN), .A(n6629), .B(
        n6628), .ZN(n6637) );
  MUX2_X1 U8301 ( .A(n6631), .B(n6630), .S(n9723), .Z(n6636) );
  NOR2_X1 U8302 ( .A1(n9723), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6632) );
  OR2_X1 U8303 ( .A1(n6632), .A2(n9726), .ZN(n6634) );
  INV_X1 U8304 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n6633) );
  AOI21_X1 U8305 ( .B1(n6634), .B2(n6633), .A(P1_U3084), .ZN(n9724) );
  OAI211_X1 U8306 ( .C1(n6636), .C2(n9726), .A(n6635), .B(n9724), .ZN(n9743)
         );
  NAND2_X1 U8307 ( .A1(n6637), .A2(n9743), .ZN(P1_U3243) );
  OR2_X1 U8308 ( .A1(n9843), .A2(n6309), .ZN(n6638) );
  AND2_X1 U8309 ( .A1(n6440), .A2(n7087), .ZN(n8834) );
  NOR2_X1 U8310 ( .A1(n7081), .A2(n8834), .ZN(n9013) );
  OR3_X1 U8311 ( .A1(n9013), .A2(n9088), .A3(n6641), .ZN(n6643) );
  NAND2_X1 U8312 ( .A1(n9106), .A2(n9484), .ZN(n6642) );
  NAND2_X1 U8313 ( .A1(n6643), .A2(n6642), .ZN(n7029) );
  INV_X1 U8314 ( .A(n7029), .ZN(n6644) );
  OAI21_X1 U8315 ( .B1(n7087), .B2(n6910), .A(n6644), .ZN(n6650) );
  NAND2_X1 U8316 ( .A1(n6650), .A2(n9910), .ZN(n6645) );
  OAI21_X1 U8317 ( .B1(n9910), .B2(n5826), .A(n6645), .ZN(P1_U3523) );
  INV_X1 U8318 ( .A(n9616), .ZN(n6647) );
  NAND2_X1 U8319 ( .A1(n6647), .A2(n6646), .ZN(n6648) );
  INV_X1 U8320 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n8394) );
  NAND2_X1 U8321 ( .A1(n6650), .A2(n9900), .ZN(n6651) );
  OAI21_X1 U8322 ( .B1(n9900), .B2(n8394), .A(n6651), .ZN(P1_U3454) );
  INV_X1 U8323 ( .A(n6652), .ZN(n6654) );
  INV_X1 U8324 ( .A(n7287), .ZN(n7278) );
  OAI222_X1 U8325 ( .A1(n8627), .A2(n6653), .B1(n7538), .B2(n6654), .C1(
        P2_U3152), .C2(n7278), .ZN(P2_U3343) );
  OAI222_X1 U8326 ( .A1(n9618), .A2(n6655), .B1(n7433), .B2(n6654), .C1(
        P1_U3084), .C2(n9141), .ZN(P1_U3338) );
  INV_X1 U8327 ( .A(n6656), .ZN(n6699) );
  INV_X1 U8328 ( .A(n7985), .ZN(n7291) );
  OAI222_X1 U8329 ( .A1(n8627), .A2(n8594), .B1(n7538), .B2(n6699), .C1(n7291), 
        .C2(P2_U3152), .ZN(P2_U3342) );
  NAND2_X1 U8330 ( .A1(P2_REG2_REG_9__SCAN_IN), .A2(n6662), .ZN(n6658) );
  NAND2_X1 U8331 ( .A1(n6658), .A2(n6657), .ZN(n7971) );
  MUX2_X1 U8332 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n7155), .S(n7968), .Z(n7970)
         );
  NAND2_X1 U8333 ( .A1(n7971), .A2(n7970), .ZN(n7969) );
  OAI21_X1 U8334 ( .B1(n7155), .B2(n6659), .A(n7969), .ZN(n6661) );
  MUX2_X1 U8335 ( .A(n7216), .B(P2_REG2_REG_11__SCAN_IN), .S(n6684), .Z(n6660)
         );
  NOR2_X1 U8336 ( .A1(n6660), .A2(n6661), .ZN(n6689) );
  AOI21_X1 U8337 ( .B1(n6661), .B2(n6660), .A(n6689), .ZN(n6674) );
  INV_X1 U8338 ( .A(n9968), .ZN(n9970) );
  NOR2_X1 U8339 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5302), .ZN(n6671) );
  INV_X1 U8340 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n10128) );
  MUX2_X1 U8341 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n10128), .S(n7968), .Z(n7975) );
  NAND2_X1 U8342 ( .A1(n6662), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n6665) );
  INV_X1 U8343 ( .A(n6663), .ZN(n6664) );
  NAND2_X1 U8344 ( .A1(n6665), .A2(n6664), .ZN(n7974) );
  NAND2_X1 U8345 ( .A1(n7968), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n6666) );
  MUX2_X1 U8346 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n5275), .S(n6684), .Z(n6667)
         );
  NOR2_X1 U8347 ( .A1(n6668), .A2(n6667), .ZN(n6669) );
  NOR3_X1 U8348 ( .A1(n9972), .A2(n6683), .A3(n6669), .ZN(n6670) );
  AOI211_X1 U8349 ( .C1(P2_ADDR_REG_11__SCAN_IN), .C2(n9969), .A(n6671), .B(
        n6670), .ZN(n6673) );
  INV_X1 U8350 ( .A(n9971), .ZN(n9659) );
  NAND2_X1 U8351 ( .A1(n9659), .A2(n6684), .ZN(n6672) );
  OAI211_X1 U8352 ( .C1(n6674), .C2(n9970), .A(n6673), .B(n6672), .ZN(P2_U3256) );
  NAND2_X1 U8353 ( .A1(n6675), .A2(n4995), .ZN(n6726) );
  OAI21_X1 U8354 ( .B1(n4995), .B2(n6675), .A(n6726), .ZN(n6676) );
  NAND2_X1 U8355 ( .A1(n6676), .A2(n8783), .ZN(n6681) );
  INV_X1 U8356 ( .A(n6677), .ZN(n6678) );
  OAI22_X1 U8357 ( .A1(n6825), .A2(n8798), .B1(n8786), .B2(n6678), .ZN(n6679)
         );
  AOI21_X1 U8358 ( .B1(n8804), .B2(n7018), .A(n6679), .ZN(n6680) );
  OAI211_X1 U8359 ( .C1(n6718), .C2(n6682), .A(n6681), .B(n6680), .ZN(P1_U3235) );
  MUX2_X1 U8360 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n6685), .S(n6815), .Z(n6686)
         );
  NAND2_X1 U8361 ( .A1(n6686), .A2(n4413), .ZN(n6814) );
  OAI21_X1 U8362 ( .B1(n4413), .B2(n6686), .A(n6814), .ZN(n6688) );
  INV_X1 U8363 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n8423) );
  NAND2_X1 U8364 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3152), .ZN(n7322) );
  OAI21_X1 U8365 ( .B1(n8022), .B2(n8423), .A(n7322), .ZN(n6687) );
  AOI21_X1 U8366 ( .B1(n9967), .B2(n6688), .A(n6687), .ZN(n6697) );
  MUX2_X1 U8367 ( .A(n7307), .B(P2_REG2_REG_12__SCAN_IN), .S(n6815), .Z(n6691)
         );
  AOI21_X1 U8368 ( .B1(n6690), .B2(n7216), .A(n6689), .ZN(n6692) );
  NOR2_X1 U8369 ( .A1(n6691), .A2(n6692), .ZN(n6811) );
  INV_X1 U8370 ( .A(n6691), .ZN(n6694) );
  INV_X1 U8371 ( .A(n6692), .ZN(n6693) );
  NOR2_X1 U8372 ( .A1(n6694), .A2(n6693), .ZN(n6695) );
  OAI21_X1 U8373 ( .B1(n6811), .B2(n6695), .A(n9968), .ZN(n6696) );
  OAI211_X1 U8374 ( .C1(n9971), .C2(n6698), .A(n6697), .B(n6696), .ZN(P2_U3257) );
  INV_X1 U8375 ( .A(n9160), .ZN(n9148) );
  OAI222_X1 U8376 ( .A1(n9618), .A2(n6700), .B1(n9148), .B2(P1_U3084), .C1(
        n7433), .C2(n6699), .ZN(P1_U3337) );
  INV_X1 U8377 ( .A(n6701), .ZN(n6889) );
  INV_X1 U8378 ( .A(n7705), .ZN(n9940) );
  INV_X1 U8379 ( .A(n7964), .ZN(n9924) );
  OAI22_X1 U8380 ( .A1(n9924), .A2(n8241), .B1(n7737), .B2(n9995), .ZN(n6771)
         );
  AOI22_X1 U8381 ( .A1(n9940), .A2(n6771), .B1(P2_REG3_REG_5__SCAN_IN), .B2(
        P2_U3152), .ZN(n6702) );
  OAI21_X1 U8382 ( .B1(n6889), .B2(n9966), .A(n6702), .ZN(n6703) );
  AOI21_X1 U8383 ( .B1(n9957), .B2(n6933), .A(n6703), .ZN(n6708) );
  OAI211_X1 U8384 ( .C1(n6706), .C2(n6705), .A(n6704), .B(n9949), .ZN(n6707)
         );
  NAND2_X1 U8385 ( .A1(n6708), .A2(n6707), .ZN(P2_U3229) );
  INV_X1 U8386 ( .A(n6709), .ZN(n6723) );
  AOI22_X1 U8387 ( .A1(n9175), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n6710), .ZN(n6711) );
  OAI21_X1 U8388 ( .B1(n6723), .B2(n7433), .A(n6711), .ZN(P1_U3336) );
  INV_X1 U8389 ( .A(n6712), .ZN(n6713) );
  NOR2_X1 U8390 ( .A1(n6714), .A2(n6713), .ZN(n6716) );
  XNOR2_X1 U8391 ( .A(n6716), .B(n6715), .ZN(n6722) );
  INV_X1 U8392 ( .A(n6440), .ZN(n6717) );
  INV_X1 U8393 ( .A(n9104), .ZN(n6834) );
  OAI22_X1 U8394 ( .A1(n6717), .A2(n8798), .B1(n8786), .B2(n6834), .ZN(n6720)
         );
  NOR2_X1 U8395 ( .A1(n6718), .A2(n7088), .ZN(n6719) );
  AOI211_X1 U8396 ( .C1(n8804), .C2(n6824), .A(n6720), .B(n6719), .ZN(n6721)
         );
  OAI21_X1 U8397 ( .B1(n6722), .B2(n8806), .A(n6721), .ZN(P1_U3220) );
  INV_X1 U8398 ( .A(n7996), .ZN(n7993) );
  OAI222_X1 U8399 ( .A1(P2_U3152), .A2(n7993), .B1(n7538), .B2(n6723), .C1(
        n8587), .C2(n8627), .ZN(P2_U3341) );
  NAND2_X1 U8400 ( .A1(n6726), .A2(n6725), .ZN(n6727) );
  OAI21_X1 U8401 ( .B1(n6724), .B2(n6727), .A(n4464), .ZN(n6731) );
  AOI22_X1 U8402 ( .A1(n8804), .A2(n7033), .B1(n8800), .B2(n9103), .ZN(n6729)
         );
  INV_X1 U8403 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n6913) );
  NOR2_X1 U8404 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6913), .ZN(n9634) );
  AOI21_X1 U8405 ( .B1(n8774), .B2(n9104), .A(n9634), .ZN(n6728) );
  OAI211_X1 U8406 ( .C1(n8802), .C2(P1_REG3_REG_3__SCAN_IN), .A(n6729), .B(
        n6728), .ZN(n6730) );
  AOI21_X1 U8407 ( .B1(n6731), .B2(n8783), .A(n6730), .ZN(n6732) );
  INV_X1 U8408 ( .A(n6732), .ZN(P1_U3216) );
  NAND2_X1 U8409 ( .A1(n6733), .A2(n8783), .ZN(n6740) );
  AOI21_X1 U8410 ( .B1(n4464), .B2(n6735), .A(n6734), .ZN(n6739) );
  AOI22_X1 U8411 ( .A1(n8804), .A2(n7074), .B1(n8800), .B2(n9102), .ZN(n6738)
         );
  AND2_X1 U8412 ( .A1(P1_U3084), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n9742) );
  NOR2_X1 U8413 ( .A1(n8802), .A2(n7067), .ZN(n6736) );
  AOI211_X1 U8414 ( .C1(n8774), .C2(n6677), .A(n9742), .B(n6736), .ZN(n6737)
         );
  OAI211_X1 U8415 ( .C1(n6740), .C2(n6739), .A(n6738), .B(n6737), .ZN(P1_U3228) );
  NOR2_X1 U8416 ( .A1(n10037), .A2(n6741), .ZN(n7530) );
  AND2_X1 U8417 ( .A1(n7530), .A2(n6883), .ZN(n6743) );
  NAND2_X1 U8418 ( .A1(n6743), .A2(n6742), .ZN(n6744) );
  OR2_X1 U8419 ( .A1(n6745), .A2(n6744), .ZN(n6778) );
  INV_X2 U8420 ( .A(n10131), .ZN(n10124) );
  INV_X1 U8421 ( .A(n6747), .ZN(n6746) );
  NAND2_X1 U8422 ( .A1(n6765), .A2(n6940), .ZN(n6939) );
  OR2_X1 U8423 ( .A1(n6747), .A2(n6748), .ZN(n6749) );
  NAND2_X1 U8424 ( .A1(n6939), .A2(n6749), .ZN(n6982) );
  NAND2_X1 U8425 ( .A1(n7965), .A2(n6750), .ZN(n7755) );
  NAND2_X1 U8426 ( .A1(n7753), .A2(n7755), .ZN(n6983) );
  NAND2_X1 U8427 ( .A1(n6982), .A2(n6983), .ZN(n6752) );
  OR2_X1 U8428 ( .A1(n7965), .A2(n7686), .ZN(n6751) );
  INV_X1 U8429 ( .A(n6773), .ZN(n6754) );
  NAND2_X1 U8430 ( .A1(n6754), .A2(n6753), .ZN(n10008) );
  NAND2_X1 U8431 ( .A1(n9937), .A2(n6773), .ZN(n7734) );
  NAND2_X1 U8432 ( .A1(n10008), .A2(n7734), .ZN(n6784) );
  OR2_X1 U8433 ( .A1(n9937), .A2(n6754), .ZN(n6755) );
  OR2_X1 U8434 ( .A1(n7964), .A2(n6756), .ZN(n7730) );
  NAND2_X1 U8435 ( .A1(n7964), .A2(n6756), .ZN(n6924) );
  NAND2_X1 U8436 ( .A1(n7730), .A2(n6924), .ZN(n10014) );
  OR2_X1 U8437 ( .A1(n7964), .A2(n10025), .ZN(n6757) );
  OR2_X1 U8438 ( .A1(n9936), .A2(n6890), .ZN(n7741) );
  NAND2_X1 U8439 ( .A1(n9936), .A2(n6890), .ZN(n7733) );
  NAND2_X1 U8440 ( .A1(n7741), .A2(n7733), .ZN(n7897) );
  NAND2_X1 U8441 ( .A1(n6758), .A2(n7897), .ZN(n6935) );
  OAI21_X1 U8442 ( .B1(n6758), .B2(n7897), .A(n6935), .ZN(n6759) );
  INV_X1 U8443 ( .A(n6759), .ZN(n6895) );
  OAI22_X1 U8444 ( .A1(n6762), .A2(n6761), .B1(n6760), .B2(n7536), .ZN(n6763)
         );
  NAND2_X1 U8445 ( .A1(n6763), .A2(n7925), .ZN(n9989) );
  INV_X1 U8446 ( .A(n7746), .ZN(n6941) );
  NAND2_X1 U8447 ( .A1(n6941), .A2(n7895), .ZN(n6977) );
  NAND2_X1 U8448 ( .A1(n6977), .A2(n7752), .ZN(n6767) );
  INV_X1 U8449 ( .A(n6983), .ZN(n7896) );
  NAND2_X1 U8450 ( .A1(n6767), .A2(n7896), .ZN(n6979) );
  NAND2_X1 U8451 ( .A1(n6979), .A2(n7753), .ZN(n6768) );
  INV_X1 U8452 ( .A(n6784), .ZN(n7894) );
  NAND2_X1 U8453 ( .A1(n6768), .A2(n7894), .ZN(n6783) );
  NAND2_X1 U8454 ( .A1(n7730), .A2(n10008), .ZN(n7743) );
  INV_X1 U8455 ( .A(n7743), .ZN(n6769) );
  NAND2_X1 U8456 ( .A1(n6783), .A2(n6769), .ZN(n6925) );
  NAND2_X1 U8457 ( .A1(n6925), .A2(n6924), .ZN(n6770) );
  XNOR2_X1 U8458 ( .A(n6770), .B(n7897), .ZN(n6772) );
  NAND2_X1 U8459 ( .A1(n5048), .A2(n8081), .ZN(n7924) );
  AOI21_X1 U8460 ( .B1(n6772), .B2(n10012), .A(n6771), .ZN(n6885) );
  NAND2_X1 U8461 ( .A1(n10055), .A2(n7554), .ZN(n6971) );
  INV_X1 U8462 ( .A(n6950), .ZN(n6774) );
  AOI211_X1 U8463 ( .C1(n6933), .C2(n10023), .A(n10102), .B(n6774), .ZN(n6892)
         );
  AOI21_X1 U8464 ( .B1(n10024), .B2(n6933), .A(n6892), .ZN(n6775) );
  OAI211_X1 U8465 ( .C1(n6895), .C2(n8331), .A(n6885), .B(n6775), .ZN(n6779)
         );
  NAND2_X1 U8466 ( .A1(n6779), .A2(n10124), .ZN(n6776) );
  OAI21_X1 U8467 ( .B1(n10124), .B2(n6464), .A(n6776), .ZN(P2_U3525) );
  NAND2_X1 U8468 ( .A1(n6779), .A2(n10117), .ZN(n6780) );
  OAI21_X1 U8469 ( .B1(n10117), .B2(n5130), .A(n6780), .ZN(P2_U3466) );
  OAI21_X1 U8470 ( .B1(n6782), .B2(n6784), .A(n6781), .ZN(n6964) );
  INV_X1 U8471 ( .A(n6964), .ZN(n6790) );
  INV_X1 U8472 ( .A(n9989), .ZN(n7152) );
  INV_X1 U8473 ( .A(n7965), .ZN(n9925) );
  OAI22_X1 U8474 ( .A1(n9925), .A2(n8241), .B1(n9924), .B2(n9995), .ZN(n6787)
         );
  NAND3_X1 U8475 ( .A1(n6979), .A2(n6784), .A3(n7753), .ZN(n6785) );
  AOI21_X1 U8476 ( .B1(n6783), .B2(n6785), .A(n8226), .ZN(n6786) );
  AOI211_X1 U8477 ( .C1(n7152), .C2(n6964), .A(n6787), .B(n6786), .ZN(n6970)
         );
  INV_X1 U8478 ( .A(n6973), .ZN(n6788) );
  AOI211_X1 U8479 ( .C1(n6754), .C2(n6788), .A(n10102), .B(n4540), .ZN(n6965)
         );
  AOI21_X1 U8480 ( .B1(n10024), .B2(n6754), .A(n6965), .ZN(n6789) );
  OAI211_X1 U8481 ( .C1(n6790), .C2(n10080), .A(n6970), .B(n6789), .ZN(n6792)
         );
  NAND2_X1 U8482 ( .A1(n6792), .A2(n10117), .ZN(n6791) );
  OAI21_X1 U8483 ( .B1(n10117), .B2(n5083), .A(n6791), .ZN(P2_U3460) );
  INV_X1 U8484 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6794) );
  NAND2_X1 U8485 ( .A1(n6792), .A2(n10124), .ZN(n6793) );
  OAI21_X1 U8486 ( .B1(n10124), .B2(n6794), .A(n6793), .ZN(P2_U3523) );
  OAI21_X1 U8487 ( .B1(n6797), .B2(n6796), .A(n6795), .ZN(n6798) );
  NAND2_X1 U8488 ( .A1(n6798), .A2(n9949), .ZN(n6805) );
  INV_X1 U8489 ( .A(n6799), .ZN(n6953) );
  INV_X1 U8490 ( .A(n9966), .ZN(n7719) );
  NAND2_X1 U8491 ( .A1(n9993), .A2(n9935), .ZN(n6801) );
  NAND2_X1 U8492 ( .A1(n9936), .A2(n9992), .ZN(n6800) );
  AND2_X1 U8493 ( .A1(n6801), .A2(n6800), .ZN(n6957) );
  OAI22_X1 U8494 ( .A1(n7705), .A2(n6957), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6802), .ZN(n6803) );
  AOI21_X1 U8495 ( .B1(n6953), .B2(n7719), .A(n6803), .ZN(n6804) );
  OAI211_X1 U8496 ( .C1(n10070), .C2(n7723), .A(n6805), .B(n6804), .ZN(
        P2_U3241) );
  INV_X1 U8497 ( .A(n6806), .ZN(n6808) );
  AOI22_X1 U8498 ( .A1(n8011), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n8633), .ZN(n6807) );
  OAI21_X1 U8499 ( .B1(n6808), .B2(n8635), .A(n6807), .ZN(P2_U3340) );
  INV_X1 U8500 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n6809) );
  INV_X1 U8501 ( .A(n9814), .ZN(n9172) );
  OAI222_X1 U8502 ( .A1(n9618), .A2(n6809), .B1(n7433), .B2(n6808), .C1(
        P1_U3084), .C2(n9172), .ZN(P1_U3335) );
  NOR2_X1 U8503 ( .A1(n6815), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n6810) );
  NOR2_X1 U8504 ( .A1(n6811), .A2(n6810), .ZN(n6813) );
  AOI22_X1 U8505 ( .A1(n6866), .A2(n7424), .B1(P2_REG2_REG_13__SCAN_IN), .B2(
        n6861), .ZN(n6812) );
  NOR2_X1 U8506 ( .A1(n6813), .A2(n6812), .ZN(n6860) );
  AOI21_X1 U8507 ( .B1(n6813), .B2(n6812), .A(n6860), .ZN(n6823) );
  INV_X1 U8508 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n6820) );
  AOI22_X1 U8509 ( .A1(n6866), .A2(P2_REG1_REG_13__SCAN_IN), .B1(n5328), .B2(
        n6861), .ZN(n6817) );
  OAI21_X1 U8510 ( .B1(P2_REG1_REG_12__SCAN_IN), .B2(n6815), .A(n6814), .ZN(
        n6816) );
  NAND2_X1 U8511 ( .A1(n6817), .A2(n6816), .ZN(n6865) );
  OAI21_X1 U8512 ( .B1(n6817), .B2(n6816), .A(n6865), .ZN(n6818) );
  NAND2_X1 U8513 ( .A1(n9967), .A2(n6818), .ZN(n6819) );
  NAND2_X1 U8514 ( .A1(P2_U3152), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n7373) );
  OAI211_X1 U8515 ( .C1(n8022), .C2(n6820), .A(n6819), .B(n7373), .ZN(n6821)
         );
  AOI21_X1 U8516 ( .B1(n6866), .B2(n9659), .A(n6821), .ZN(n6822) );
  OAI21_X1 U8517 ( .B1(n6823), .B2(n9970), .A(n6822), .ZN(P2_U3258) );
  NAND2_X1 U8518 ( .A1(n9106), .A2(n9846), .ZN(n8836) );
  NAND2_X1 U8519 ( .A1(n9015), .A2(n7079), .ZN(n7078) );
  NAND2_X1 U8520 ( .A1(n9106), .A2(n6824), .ZN(n6826) );
  XNOR2_X1 U8521 ( .A(n9104), .B(n9850), .ZN(n7012) );
  OR2_X1 U8522 ( .A1(n9104), .A2(n7018), .ZN(n6827) );
  NAND2_X1 U8523 ( .A1(n7011), .A2(n6827), .ZN(n7036) );
  OR2_X1 U8524 ( .A1(n6677), .A2(n6915), .ZN(n9048) );
  NAND2_X1 U8525 ( .A1(n6677), .A2(n6915), .ZN(n9044) );
  NAND2_X1 U8526 ( .A1(n9048), .A2(n9044), .ZN(n7049) );
  NAND2_X1 U8527 ( .A1(n7036), .A2(n7049), .ZN(n7059) );
  OAI21_X1 U8528 ( .B1(n7036), .B2(n7049), .A(n7059), .ZN(n6842) );
  INV_X1 U8529 ( .A(n6842), .ZN(n6918) );
  OR2_X1 U8530 ( .A1(n6916), .A2(n6828), .ZN(n6831) );
  OR2_X1 U8531 ( .A1(n6829), .A2(n9069), .ZN(n6830) );
  AND2_X1 U8532 ( .A1(n6831), .A2(n6830), .ZN(n7340) );
  INV_X1 U8533 ( .A(n7340), .ZN(n7353) );
  INV_X1 U8534 ( .A(n9103), .ZN(n6833) );
  OAI22_X1 U8535 ( .A1(n6834), .A2(n9424), .B1(n6833), .B2(n9422), .ZN(n6841)
         );
  INV_X1 U8536 ( .A(n7012), .ZN(n9017) );
  NAND2_X1 U8537 ( .A1(n7020), .A2(n9017), .ZN(n7019) );
  OR2_X1 U8538 ( .A1(n9104), .A2(n9850), .ZN(n6836) );
  XNOR2_X1 U8539 ( .A(n9046), .B(n7049), .ZN(n6839) );
  NAND2_X1 U8540 ( .A1(n6310), .A2(n9356), .ZN(n6838) );
  NAND2_X1 U8541 ( .A1(n6309), .A2(n9080), .ZN(n6837) );
  NOR2_X1 U8542 ( .A1(n6839), .A2(n9420), .ZN(n6840) );
  AOI211_X1 U8543 ( .C1(n7353), .C2(n6842), .A(n6841), .B(n6840), .ZN(n6923)
         );
  OR2_X1 U8544 ( .A1(n6824), .A2(n7030), .ZN(n7086) );
  INV_X1 U8545 ( .A(n6843), .ZN(n7014) );
  NAND2_X1 U8546 ( .A1(n6843), .A2(n6915), .ZN(n7070) );
  INV_X1 U8547 ( .A(n7070), .ZN(n6844) );
  AOI21_X1 U8548 ( .B1(n7033), .B2(n7014), .A(n6844), .ZN(n6921) );
  AOI22_X1 U8549 ( .A1(n6921), .A2(n9590), .B1(n9892), .B2(n7033), .ZN(n6845)
         );
  OAI211_X1 U8550 ( .C1(n6918), .C2(n9843), .A(n6923), .B(n6845), .ZN(n6847)
         );
  NAND2_X1 U8551 ( .A1(n6847), .A2(n9910), .ZN(n6846) );
  OAI21_X1 U8552 ( .B1(n9910), .B2(n6366), .A(n6846), .ZN(P1_U3526) );
  NAND2_X1 U8553 ( .A1(n6847), .A2(n9900), .ZN(n6848) );
  OAI21_X1 U8554 ( .B1(n9900), .B2(n4949), .A(n6848), .ZN(P1_U3463) );
  AOI21_X1 U8555 ( .B1(n6850), .B2(n6849), .A(n7709), .ZN(n6852) );
  NAND2_X1 U8556 ( .A1(n6852), .A2(n6851), .ZN(n6859) );
  INV_X1 U8557 ( .A(n6930), .ZN(n6857) );
  OR2_X1 U8558 ( .A1(n7737), .A2(n8241), .ZN(n6854) );
  NAND2_X1 U8559 ( .A1(n7961), .A2(n9935), .ZN(n6853) );
  AND2_X1 U8560 ( .A1(n6854), .A2(n6853), .ZN(n6928) );
  INV_X1 U8561 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n6855) );
  OAI22_X1 U8562 ( .A1(n7705), .A2(n6928), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6855), .ZN(n6856) );
  AOI21_X1 U8563 ( .B1(n6857), .B2(n7719), .A(n6856), .ZN(n6858) );
  OAI211_X1 U8564 ( .C1(n10075), .C2(n7723), .A(n6859), .B(n6858), .ZN(
        P2_U3215) );
  AOI21_X1 U8565 ( .B1(n6861), .B2(n7424), .A(n6860), .ZN(n6864) );
  NOR2_X1 U8566 ( .A1(n7248), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n7245) );
  INV_X1 U8567 ( .A(n7245), .ZN(n6862) );
  OAI21_X1 U8568 ( .B1(n7449), .B2(n6871), .A(n6862), .ZN(n6863) );
  NOR2_X1 U8569 ( .A1(n6864), .A2(n6863), .ZN(n7244) );
  AOI21_X1 U8570 ( .B1(n6864), .B2(n6863), .A(n7244), .ZN(n6876) );
  OAI21_X1 U8571 ( .B1(n6866), .B2(P2_REG1_REG_13__SCAN_IN), .A(n6865), .ZN(
        n6869) );
  MUX2_X1 U8572 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n6867), .S(n7248), .Z(n6868)
         );
  NAND2_X1 U8573 ( .A1(n6868), .A2(n6869), .ZN(n7247) );
  OAI21_X1 U8574 ( .B1(n6869), .B2(n6868), .A(n7247), .ZN(n6874) );
  INV_X1 U8575 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n6870) );
  NAND2_X1 U8576 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3152), .ZN(n7477) );
  OAI21_X1 U8577 ( .B1(n8022), .B2(n6870), .A(n7477), .ZN(n6873) );
  NOR2_X1 U8578 ( .A1(n9971), .A2(n6871), .ZN(n6872) );
  AOI211_X1 U8579 ( .C1(n9967), .C2(n6874), .A(n6873), .B(n6872), .ZN(n6875)
         );
  OAI21_X1 U8580 ( .B1(n6876), .B2(n9970), .A(n6875), .ZN(P2_U3259) );
  INV_X1 U8581 ( .A(n6877), .ZN(n6879) );
  OAI222_X1 U8582 ( .A1(n9618), .A2(n6878), .B1(n7433), .B2(n6879), .C1(n9321), 
        .C2(P1_U3084), .ZN(P1_U3334) );
  OAI222_X1 U8583 ( .A1(n8627), .A2(n8340), .B1(n7538), .B2(n6879), .C1(
        P2_U3152), .C2(n8020), .ZN(P2_U3339) );
  AND2_X1 U8584 ( .A1(n7530), .A2(n6880), .ZN(n6881) );
  NAND2_X1 U8585 ( .A1(n6882), .A2(n6881), .ZN(n6887) );
  INV_X1 U8586 ( .A(n6883), .ZN(n6884) );
  NOR2_X1 U8587 ( .A1(n7932), .A2(n8020), .ZN(n7724) );
  NAND2_X1 U8588 ( .A1(n7724), .A2(n7536), .ZN(n6962) );
  NAND2_X1 U8589 ( .A1(n9989), .A2(n6962), .ZN(n10018) );
  MUX2_X1 U8590 ( .A(n6886), .B(n6885), .S(n10035), .Z(n6894) );
  OR2_X1 U8591 ( .A1(n6887), .A2(n8081), .ZN(n7503) );
  NOR2_X1 U8592 ( .A1(n7925), .A2(n7536), .ZN(n6888) );
  OAI22_X1 U8593 ( .A1(n10001), .A2(n6890), .B1(n10028), .B2(n6889), .ZN(n6891) );
  AOI21_X1 U8594 ( .B1(n6892), .B2(n8222), .A(n6891), .ZN(n6893) );
  OAI211_X1 U8595 ( .C1(n6895), .C2(n8232), .A(n6894), .B(n6893), .ZN(P2_U3291) );
  OAI211_X1 U8596 ( .C1(n6898), .C2(n6897), .A(n6896), .B(n9949), .ZN(n6903)
         );
  INV_X1 U8597 ( .A(n9959), .ZN(n9918) );
  OAI22_X1 U8598 ( .A1(n9966), .A2(n10002), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6899), .ZN(n6901) );
  INV_X1 U8599 ( .A(n9982), .ZN(n10082) );
  OAI22_X1 U8600 ( .A1(n7723), .A2(n10082), .B1(n9954), .B2(n9996), .ZN(n6900)
         );
  AOI211_X1 U8601 ( .C1(n9918), .C2(n9993), .A(n6901), .B(n6900), .ZN(n6902)
         );
  NAND2_X1 U8602 ( .A1(n6903), .A2(n6902), .ZN(P2_U3223) );
  NOR2_X1 U8603 ( .A1(n8254), .A2(n8071), .ZN(n10031) );
  NAND2_X1 U8604 ( .A1(n6764), .A2(n7554), .ZN(n7750) );
  NAND2_X1 U8605 ( .A1(n7746), .A2(n7750), .ZN(n10051) );
  AOI22_X1 U8606 ( .A1(n10051), .A2(n10012), .B1(n9935), .B2(n7966), .ZN(
        n10053) );
  OAI21_X1 U8607 ( .B1(n5049), .B2(n10028), .A(n10053), .ZN(n6904) );
  MUX2_X1 U8608 ( .A(P2_REG2_REG_0__SCAN_IN), .B(n6904), .S(n10035), .Z(n6905)
         );
  AOI21_X1 U8609 ( .B1(n7500), .B2(n10051), .A(n6905), .ZN(n6906) );
  OAI21_X1 U8610 ( .B1(n10031), .B2(n7554), .A(n6906), .ZN(P2_U3296) );
  INV_X1 U8611 ( .A(n6907), .ZN(n9839) );
  NAND2_X1 U8612 ( .A1(n6908), .A2(n9839), .ZN(n7138) );
  NAND2_X1 U8613 ( .A1(n9069), .A2(n9841), .ZN(n6909) );
  NOR2_X1 U8614 ( .A1(n6910), .A2(n9085), .ZN(n6911) );
  INV_X1 U8615 ( .A(n9407), .ZN(n9477) );
  AOI22_X1 U8616 ( .A1(n9447), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n9477), .B2(
        n6913), .ZN(n6914) );
  OAI21_X1 U8617 ( .B1(n6915), .B2(n9480), .A(n6914), .ZN(n6920) );
  AND2_X1 U8618 ( .A1(n6916), .A2(n9356), .ZN(n6917) );
  NAND2_X1 U8619 ( .A1(n9425), .A2(n6917), .ZN(n7370) );
  NOR2_X1 U8620 ( .A1(n6918), .A2(n7370), .ZN(n6919) );
  AOI211_X1 U8621 ( .C1(n6921), .C2(n9493), .A(n6920), .B(n6919), .ZN(n6922)
         );
  OAI21_X1 U8622 ( .B1(n6923), .B2(n9490), .A(n6922), .ZN(P1_U3288) );
  AND2_X1 U8623 ( .A1(n7733), .A2(n6924), .ZN(n7735) );
  NAND2_X1 U8624 ( .A1(n6925), .A2(n7735), .ZN(n6926) );
  INV_X1 U8625 ( .A(n7737), .ZN(n7962) );
  NAND2_X1 U8626 ( .A1(n6956), .A2(n7899), .ZN(n6927) );
  OR2_X1 U8627 ( .A1(n7962), .A2(n10070), .ZN(n7762) );
  NAND2_X1 U8628 ( .A1(n6927), .A2(n7762), .ZN(n7100) );
  NAND2_X1 U8629 ( .A1(n9993), .A2(n10075), .ZN(n7768) );
  XNOR2_X1 U8630 ( .A(n7100), .B(n7099), .ZN(n6929) );
  OAI21_X1 U8631 ( .B1(n6929), .B2(n8226), .A(n6928), .ZN(n10077) );
  INV_X1 U8632 ( .A(n10077), .ZN(n6938) );
  INV_X1 U8633 ( .A(n10075), .ZN(n7093) );
  OAI22_X1 U8634 ( .A1(n10035), .A2(n6512), .B1(n6930), .B2(n10028), .ZN(n6932) );
  INV_X1 U8635 ( .A(n8254), .ZN(n9986) );
  NAND2_X1 U8636 ( .A1(n6949), .A2(n10075), .ZN(n9983) );
  OAI21_X1 U8637 ( .B1(n6949), .B2(n10075), .A(n9983), .ZN(n10076) );
  NOR2_X1 U8638 ( .A1(n9986), .A2(n10076), .ZN(n6931) );
  AOI211_X1 U8639 ( .C1(n8071), .C2(n7093), .A(n6932), .B(n6931), .ZN(n6937)
         );
  OR2_X1 U8640 ( .A1(n9936), .A2(n6933), .ZN(n6934) );
  XNOR2_X1 U8641 ( .A(n7092), .B(n7099), .ZN(n10079) );
  NAND2_X1 U8642 ( .A1(n10079), .A2(n7500), .ZN(n6936) );
  OAI211_X1 U8643 ( .C1(n6938), .C2(n8208), .A(n6937), .B(n6936), .ZN(P2_U3289) );
  OAI211_X1 U8644 ( .C1(n7554), .C2(n10055), .A(n10022), .B(n6971), .ZN(n10054) );
  OAI22_X1 U8645 ( .A1(n10001), .A2(n10055), .B1(n10054), .B2(n7503), .ZN(
        n6946) );
  OAI21_X1 U8646 ( .B1(n7895), .B2(n6941), .A(n6977), .ZN(n6942) );
  AOI222_X1 U8647 ( .A1(n10012), .A2(n6942), .B1(n7965), .B2(n9935), .C1(n6764), .C2(n9992), .ZN(n10056) );
  OAI21_X1 U8648 ( .B1(n6943), .B2(n10028), .A(n10056), .ZN(n6944) );
  MUX2_X1 U8649 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n6944), .S(n10035), .Z(n6945)
         );
  AOI211_X1 U8650 ( .C1(n7500), .C2(n10059), .A(n6946), .B(n6945), .ZN(n6947)
         );
  INV_X1 U8651 ( .A(n6947), .ZN(P2_U3295) );
  XOR2_X1 U8652 ( .A(n4482), .B(n7899), .Z(n10074) );
  INV_X1 U8653 ( .A(n6949), .ZN(n6952) );
  NAND2_X1 U8654 ( .A1(n6950), .A2(n7736), .ZN(n6951) );
  NAND2_X1 U8655 ( .A1(n6952), .A2(n6951), .ZN(n10071) );
  INV_X1 U8656 ( .A(n10071), .ZN(n6954) );
  INV_X1 U8657 ( .A(n10028), .ZN(n8249) );
  AOI22_X1 U8658 ( .A1(n6954), .A2(n8254), .B1(n6953), .B2(n8249), .ZN(n6955)
         );
  OAI21_X1 U8659 ( .B1(n10070), .B2(n10001), .A(n6955), .ZN(n6960) );
  XOR2_X1 U8660 ( .A(n7899), .B(n6956), .Z(n6958) );
  OAI21_X1 U8661 ( .B1(n6958), .B2(n8226), .A(n6957), .ZN(n10072) );
  MUX2_X1 U8662 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n10072), .S(n10035), .Z(n6959) );
  AOI211_X1 U8663 ( .C1(n7500), .C2(n10074), .A(n6960), .B(n6959), .ZN(n6961)
         );
  INV_X1 U8664 ( .A(n6961), .ZN(P2_U3290) );
  INV_X1 U8665 ( .A(n6962), .ZN(n6963) );
  NAND2_X1 U8666 ( .A1(n10035), .A2(n6963), .ZN(n9987) );
  INV_X1 U8667 ( .A(n9987), .ZN(n7159) );
  AOI22_X1 U8668 ( .A1(n7159), .A2(n6964), .B1(n8071), .B2(n6754), .ZN(n6969)
         );
  INV_X1 U8669 ( .A(n6965), .ZN(n6966) );
  OAI22_X1 U8670 ( .A1(n6966), .A2(n7503), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n10028), .ZN(n6967) );
  AOI21_X1 U8671 ( .B1(n8208), .B2(P2_REG2_REG_3__SCAN_IN), .A(n6967), .ZN(
        n6968) );
  OAI211_X1 U8672 ( .C1(n6970), .C2(n8208), .A(n6969), .B(n6968), .ZN(P2_U3293) );
  NAND2_X1 U8673 ( .A1(n7686), .A2(n6971), .ZN(n6972) );
  NAND2_X1 U8674 ( .A1(n6972), .A2(n10022), .ZN(n6974) );
  OR2_X1 U8675 ( .A1(n6974), .A2(n6973), .ZN(n6976) );
  NAND2_X1 U8676 ( .A1(n7686), .A2(n10024), .ZN(n6975) );
  AND2_X1 U8677 ( .A1(n6976), .A2(n6975), .ZN(n10060) );
  NAND3_X1 U8678 ( .A1(n6977), .A2(n6983), .A3(n7752), .ZN(n6978) );
  NAND2_X1 U8679 ( .A1(n6979), .A2(n6978), .ZN(n6980) );
  AOI222_X1 U8680 ( .A1(n10012), .A2(n6980), .B1(n9937), .B2(n9935), .C1(n7966), .C2(n9992), .ZN(n10061) );
  MUX2_X1 U8681 ( .A(n6981), .B(n10061), .S(n10035), .Z(n6985) );
  XNOR2_X1 U8682 ( .A(n6983), .B(n6982), .ZN(n10063) );
  AOI22_X1 U8683 ( .A1(n7500), .A2(n10063), .B1(P2_REG3_REG_2__SCAN_IN), .B2(
        n8249), .ZN(n6984) );
  OAI211_X1 U8684 ( .C1(n10031), .C2(n10060), .A(n6985), .B(n6984), .ZN(
        P2_U3294) );
  NOR2_X1 U8685 ( .A1(n6987), .A2(n6986), .ZN(n6989) );
  AOI21_X1 U8686 ( .B1(n6987), .B2(n6986), .A(n6989), .ZN(n7002) );
  NAND2_X1 U8687 ( .A1(n7002), .A2(n7003), .ZN(n7001) );
  NOR2_X1 U8688 ( .A1(n6989), .A2(n6988), .ZN(n6992) );
  INV_X1 U8689 ( .A(n6990), .ZN(n6991) );
  AOI21_X1 U8690 ( .B1(n7001), .B2(n6992), .A(n6991), .ZN(n6997) );
  AOI22_X1 U8691 ( .A1(n8804), .A2(n7133), .B1(n8800), .B2(n9100), .ZN(n6996)
         );
  NOR2_X1 U8692 ( .A1(n8802), .A2(n7043), .ZN(n6993) );
  AOI211_X1 U8693 ( .C1(n8774), .C2(n9102), .A(n6994), .B(n6993), .ZN(n6995)
         );
  OAI211_X1 U8694 ( .C1(n6997), .C2(n8806), .A(n6996), .B(n6995), .ZN(P1_U3237) );
  INV_X1 U8695 ( .A(n6998), .ZN(n7537) );
  OAI222_X1 U8696 ( .A1(n7433), .A2(n7537), .B1(P1_U3084), .B2(n7000), .C1(
        n6999), .C2(n9618), .ZN(P1_U3333) );
  OAI21_X1 U8697 ( .B1(n7003), .B2(n7002), .A(n7001), .ZN(n7007) );
  AOI22_X1 U8698 ( .A1(n8804), .A2(n7184), .B1(n8800), .B2(n9101), .ZN(n7005)
         );
  NOR2_X1 U8699 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n5871), .ZN(n9747) );
  AOI21_X1 U8700 ( .B1(n8774), .B2(n9103), .A(n9747), .ZN(n7004) );
  OAI211_X1 U8701 ( .C1(n8802), .C2(n7181), .A(n7005), .B(n7004), .ZN(n7006)
         );
  AOI21_X1 U8702 ( .B1(n7007), .B2(n8783), .A(n7006), .ZN(n7008) );
  INV_X1 U8703 ( .A(n7008), .ZN(P1_U3225) );
  OAI21_X1 U8704 ( .B1(n7013), .B2(n7012), .A(n7011), .ZN(n9854) );
  INV_X1 U8705 ( .A(n9854), .ZN(n7026) );
  INV_X1 U8706 ( .A(n9493), .ZN(n7170) );
  INV_X1 U8707 ( .A(n7086), .ZN(n7015) );
  OAI21_X1 U8708 ( .B1(n9850), .B2(n7015), .A(n7014), .ZN(n9851) );
  AOI22_X1 U8709 ( .A1(n9447), .A2(P1_REG2_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n9477), .ZN(n7016) );
  OAI21_X1 U8710 ( .B1(n7170), .B2(n9851), .A(n7016), .ZN(n7017) );
  AOI21_X1 U8711 ( .B1(n9367), .B2(n7018), .A(n7017), .ZN(n7025) );
  OAI21_X1 U8712 ( .B1(n7020), .B2(n9017), .A(n7019), .ZN(n7021) );
  NAND2_X1 U8713 ( .A1(n7021), .A2(n9489), .ZN(n7023) );
  AOI22_X1 U8714 ( .A1(n9486), .A2(n9106), .B1(n6677), .B2(n9484), .ZN(n7022)
         );
  NAND2_X1 U8715 ( .A1(n7023), .A2(n7022), .ZN(n9852) );
  NAND2_X1 U8716 ( .A1(n9852), .A2(n9425), .ZN(n7024) );
  OAI211_X1 U8717 ( .C1(n9495), .C2(n7026), .A(n7025), .B(n7024), .ZN(P1_U3289) );
  NOR2_X1 U8718 ( .A1(n9407), .A2(n7027), .ZN(n7028) );
  OAI21_X1 U8719 ( .B1(n7029), .B2(n7028), .A(n9425), .ZN(n7032) );
  OAI21_X1 U8720 ( .B1(n9367), .B2(n9493), .A(n7030), .ZN(n7031) );
  OAI211_X1 U8721 ( .C1(n5813), .C2(n9425), .A(n7032), .B(n7031), .ZN(P1_U3291) );
  OR2_X1 U8722 ( .A1(n9103), .A2(n7074), .ZN(n7034) );
  OR2_X1 U8723 ( .A1(n6677), .A2(n7033), .ZN(n7058) );
  AND2_X1 U8724 ( .A1(n7034), .A2(n7060), .ZN(n7037) );
  AND2_X1 U8725 ( .A1(n7049), .A2(n9014), .ZN(n7035) );
  NAND2_X1 U8726 ( .A1(n7036), .A2(n7035), .ZN(n7061) );
  OR2_X1 U8727 ( .A1(n9102), .A2(n9863), .ZN(n8884) );
  NAND2_X1 U8728 ( .A1(n9102), .A2(n9863), .ZN(n8891) );
  NAND2_X1 U8729 ( .A1(n9102), .A2(n7184), .ZN(n7039) );
  INV_X1 U8730 ( .A(n7040), .ZN(n7042) );
  OR2_X1 U8731 ( .A1(n9101), .A2(n9868), .ZN(n8901) );
  NAND2_X1 U8732 ( .A1(n9101), .A2(n9868), .ZN(n9050) );
  INV_X1 U8733 ( .A(n9018), .ZN(n7041) );
  OR2_X2 U8734 ( .A1(n7040), .A2(n9018), .ZN(n7135) );
  OAI21_X1 U8735 ( .B1(n7042), .B2(n7041), .A(n7135), .ZN(n9872) );
  INV_X1 U8736 ( .A(n9872), .ZN(n7057) );
  OAI22_X1 U8737 ( .A1(n9425), .A2(n7044), .B1(n7043), .B2(n9407), .ZN(n7048)
         );
  INV_X1 U8738 ( .A(n7178), .ZN(n7046) );
  INV_X1 U8739 ( .A(n7137), .ZN(n7045) );
  OAI21_X1 U8740 ( .B1(n9868), .B2(n7046), .A(n7045), .ZN(n9869) );
  NOR2_X1 U8741 ( .A1(n9869), .A2(n7170), .ZN(n7047) );
  AOI211_X1 U8742 ( .C1(n9367), .C2(n7133), .A(n7048), .B(n7047), .ZN(n7056)
         );
  INV_X1 U8743 ( .A(n7049), .ZN(n9012) );
  INV_X1 U8744 ( .A(n9049), .ZN(n8892) );
  OAI21_X1 U8745 ( .B1(n7173), .B2(n4599), .A(n8884), .ZN(n7051) );
  XNOR2_X1 U8746 ( .A(n7051), .B(n9018), .ZN(n7052) );
  NAND2_X1 U8747 ( .A1(n7052), .A2(n9489), .ZN(n7054) );
  AOI22_X1 U8748 ( .A1(n9486), .A2(n9102), .B1(n9100), .B2(n9484), .ZN(n7053)
         );
  NAND2_X1 U8749 ( .A1(n7054), .A2(n7053), .ZN(n9870) );
  NAND2_X1 U8750 ( .A1(n9870), .A2(n9425), .ZN(n7055) );
  OAI211_X1 U8751 ( .C1(n7057), .C2(n9495), .A(n7056), .B(n7055), .ZN(P1_U3285) );
  NAND2_X1 U8752 ( .A1(n7059), .A2(n7058), .ZN(n7063) );
  AND2_X1 U8753 ( .A1(n7061), .A2(n7060), .ZN(n7062) );
  OAI21_X1 U8754 ( .B1(n7063), .B2(n9014), .A(n7062), .ZN(n9859) );
  INV_X1 U8755 ( .A(n9859), .ZN(n7077) );
  XNOR2_X1 U8756 ( .A(n9014), .B(n8889), .ZN(n7066) );
  NAND2_X1 U8757 ( .A1(n9859), .A2(n7353), .ZN(n7065) );
  AOI22_X1 U8758 ( .A1(n9486), .A2(n6677), .B1(n9102), .B2(n9484), .ZN(n7064)
         );
  OAI211_X1 U8759 ( .C1(n9420), .C2(n7066), .A(n7065), .B(n7064), .ZN(n9857)
         );
  NAND2_X1 U8760 ( .A1(n9857), .A2(n9425), .ZN(n7076) );
  OAI22_X1 U8761 ( .A1(n9425), .A2(n7068), .B1(n7067), .B2(n9407), .ZN(n7073)
         );
  NAND2_X1 U8762 ( .A1(n7070), .A2(n7074), .ZN(n7071) );
  NAND2_X1 U8763 ( .A1(n7177), .A2(n7071), .ZN(n9856) );
  NOR2_X1 U8764 ( .A1(n7170), .A2(n9856), .ZN(n7072) );
  AOI211_X1 U8765 ( .C1(n9367), .C2(n7074), .A(n7073), .B(n7072), .ZN(n7075)
         );
  OAI211_X1 U8766 ( .C1(n7077), .C2(n7370), .A(n7076), .B(n7075), .ZN(P1_U3287) );
  OAI21_X1 U8767 ( .B1(n9015), .B2(n7079), .A(n7078), .ZN(n9844) );
  AOI22_X1 U8768 ( .A1(n9486), .A2(n6440), .B1(n9104), .B2(n9484), .ZN(n7085)
         );
  OAI21_X1 U8769 ( .B1(n7082), .B2(n7081), .A(n7080), .ZN(n7083) );
  NAND2_X1 U8770 ( .A1(n7083), .A2(n9489), .ZN(n7084) );
  OAI211_X1 U8771 ( .C1(n9844), .C2(n7340), .A(n7085), .B(n7084), .ZN(n9847)
         );
  OAI211_X1 U8772 ( .C1(n7087), .C2(n9846), .A(n9590), .B(n7086), .ZN(n9845)
         );
  OAI22_X1 U8773 ( .A1(n9845), .A2(n9356), .B1(n9407), .B2(n7088), .ZN(n7089)
         );
  OAI21_X1 U8774 ( .B1(n9847), .B2(n7089), .A(n9425), .ZN(n7091) );
  AOI22_X1 U8775 ( .A1(n9367), .A2(n6824), .B1(n9490), .B2(
        P1_REG2_REG_1__SCAN_IN), .ZN(n7090) );
  OAI211_X1 U8776 ( .C1(n9844), .C2(n7370), .A(n7091), .B(n7090), .ZN(P1_U3290) );
  INV_X1 U8777 ( .A(n9980), .ZN(n7095) );
  XNOR2_X1 U8778 ( .A(n7961), .B(n9982), .ZN(n9990) );
  NAND2_X1 U8779 ( .A1(n7095), .A2(n7094), .ZN(n9978) );
  NAND2_X1 U8780 ( .A1(n7961), .A2(n9982), .ZN(n7096) );
  AND2_X2 U8781 ( .A1(n9978), .A2(n7096), .ZN(n7098) );
  OR2_X1 U8782 ( .A1(n9996), .A2(n7144), .ZN(n7781) );
  NAND2_X1 U8783 ( .A1(n9996), .A2(n7144), .ZN(n7779) );
  OAI21_X1 U8784 ( .B1(n7098), .B2(n7097), .A(n4480), .ZN(n10091) );
  INV_X1 U8785 ( .A(n10091), .ZN(n7114) );
  INV_X1 U8786 ( .A(n7099), .ZN(n7901) );
  NAND2_X1 U8787 ( .A1(n7100), .A2(n7901), .ZN(n7101) );
  NAND2_X1 U8788 ( .A1(n7101), .A2(n7769), .ZN(n9991) );
  NAND2_X1 U8789 ( .A1(n9991), .A2(n9990), .ZN(n7102) );
  OR2_X1 U8790 ( .A1(n7961), .A2(n10082), .ZN(n7772) );
  XOR2_X1 U8791 ( .A(n7900), .B(n7147), .Z(n7106) );
  OR2_X1 U8792 ( .A1(n9958), .A2(n9995), .ZN(n7104) );
  NAND2_X1 U8793 ( .A1(n7961), .A2(n9992), .ZN(n7103) );
  NAND2_X1 U8794 ( .A1(n7104), .A2(n7103), .ZN(n7120) );
  INV_X1 U8795 ( .A(n7120), .ZN(n7105) );
  OAI21_X1 U8796 ( .B1(n7106), .B2(n8226), .A(n7105), .ZN(n10089) );
  INV_X1 U8797 ( .A(n7144), .ZN(n10087) );
  INV_X1 U8798 ( .A(n9985), .ZN(n7108) );
  INV_X1 U8799 ( .A(n7153), .ZN(n7107) );
  OAI21_X1 U8800 ( .B1(n10087), .B2(n7108), .A(n7107), .ZN(n10088) );
  OAI22_X1 U8801 ( .A1(n10035), .A2(n7109), .B1(n7123), .B2(n10028), .ZN(n7110) );
  AOI21_X1 U8802 ( .B1(n8071), .B2(n7144), .A(n7110), .ZN(n7111) );
  OAI21_X1 U8803 ( .B1(n10088), .B2(n9986), .A(n7111), .ZN(n7112) );
  AOI21_X1 U8804 ( .B1(n10089), .B2(n10035), .A(n7112), .ZN(n7113) );
  OAI21_X1 U8805 ( .B1(n7114), .B2(n8232), .A(n7113), .ZN(P2_U3287) );
  INV_X1 U8806 ( .A(n7115), .ZN(n7127) );
  OAI222_X1 U8807 ( .A1(n7433), .A2(n7127), .B1(P1_U3084), .B2(n9069), .C1(
        n7116), .C2(n9618), .ZN(P1_U3332) );
  OAI21_X1 U8808 ( .B1(n7119), .B2(n7118), .A(n7117), .ZN(n7125) );
  AOI22_X1 U8809 ( .A1(n9940), .A2(n7120), .B1(P2_REG3_REG_9__SCAN_IN), .B2(
        P2_U3152), .ZN(n7122) );
  NAND2_X1 U8810 ( .A1(n9957), .A2(n7144), .ZN(n7121) );
  OAI211_X1 U8811 ( .C1(n9966), .C2(n7123), .A(n7122), .B(n7121), .ZN(n7124)
         );
  AOI21_X1 U8812 ( .B1(n7125), .B2(n9949), .A(n7124), .ZN(n7126) );
  INV_X1 U8813 ( .A(n7126), .ZN(P2_U3233) );
  OAI222_X1 U8814 ( .A1(n8627), .A2(n7128), .B1(n7538), .B2(n7127), .C1(n7932), 
        .C2(P2_U3152), .ZN(P2_U3337) );
  NAND2_X1 U8815 ( .A1(n8901), .A2(n8884), .ZN(n9051) );
  INV_X1 U8816 ( .A(n9051), .ZN(n7129) );
  NAND2_X1 U8817 ( .A1(n9050), .A2(n8891), .ZN(n7130) );
  NAND2_X1 U8818 ( .A1(n7130), .A2(n8901), .ZN(n8833) );
  OR2_X1 U8819 ( .A1(n9100), .A2(n9876), .ZN(n8900) );
  NAND2_X1 U8820 ( .A1(n9100), .A2(n9876), .ZN(n8902) );
  NAND2_X1 U8821 ( .A1(n8900), .A2(n8902), .ZN(n8897) );
  XNOR2_X1 U8822 ( .A(n8841), .B(n8897), .ZN(n7132) );
  AOI222_X1 U8823 ( .A1(n9489), .A2(n7132), .B1(n9099), .B2(n9484), .C1(n9101), 
        .C2(n9486), .ZN(n9875) );
  OR2_X1 U8824 ( .A1(n9101), .A2(n7133), .ZN(n7134) );
  NAND2_X1 U8825 ( .A1(n7136), .A2(n8897), .ZN(n7162) );
  OAI21_X1 U8826 ( .B1(n7136), .B2(n8897), .A(n7162), .ZN(n9878) );
  INV_X1 U8827 ( .A(n9495), .ZN(n9366) );
  OAI211_X1 U8828 ( .C1(n7137), .C2(n9876), .A(n7166), .B(n9590), .ZN(n9874)
         );
  NOR2_X1 U8829 ( .A1(n7138), .A2(n9356), .ZN(n9457) );
  INV_X1 U8830 ( .A(n9457), .ZN(n7469) );
  OAI22_X1 U8831 ( .A1(n9425), .A2(n7139), .B1(n8645), .B2(n9407), .ZN(n7140)
         );
  AOI21_X1 U8832 ( .B1(n9367), .B2(n8646), .A(n7140), .ZN(n7141) );
  OAI21_X1 U8833 ( .B1(n9874), .B2(n7469), .A(n7141), .ZN(n7142) );
  AOI21_X1 U8834 ( .B1(n9878), .B2(n9366), .A(n7142), .ZN(n7143) );
  OAI21_X1 U8835 ( .B1(n9875), .B2(n9490), .A(n7143), .ZN(P1_U3284) );
  INV_X1 U8836 ( .A(n9996), .ZN(n9917) );
  OR2_X1 U8837 ( .A1(n7144), .A2(n9917), .ZN(n7145) );
  OR2_X1 U8838 ( .A1(n9916), .A2(n9958), .ZN(n7786) );
  NAND2_X1 U8839 ( .A1(n9916), .A2(n9958), .ZN(n7784) );
  XNOR2_X1 U8840 ( .A(n7205), .B(n4395), .ZN(n10097) );
  XNOR2_X1 U8841 ( .A(n7209), .B(n4395), .ZN(n7150) );
  OAI22_X1 U8842 ( .A1(n7324), .A2(n9995), .B1(n9996), .B2(n8241), .ZN(n7148)
         );
  INV_X1 U8843 ( .A(n7148), .ZN(n7149) );
  OAI21_X1 U8844 ( .B1(n7150), .B2(n8226), .A(n7149), .ZN(n7151) );
  AOI21_X1 U8845 ( .B1(n10097), .B2(n7152), .A(n7151), .ZN(n10099) );
  INV_X1 U8846 ( .A(n9916), .ZN(n10093) );
  NOR2_X1 U8847 ( .A1(n7153), .A2(n10093), .ZN(n7154) );
  OR2_X1 U8848 ( .A1(n7215), .A2(n7154), .ZN(n10094) );
  OAI22_X1 U8849 ( .A1(n10035), .A2(n7155), .B1(n9923), .B2(n10028), .ZN(n7156) );
  AOI21_X1 U8850 ( .B1(n8071), .B2(n9916), .A(n7156), .ZN(n7157) );
  OAI21_X1 U8851 ( .B1(n10094), .B2(n9986), .A(n7157), .ZN(n7158) );
  AOI21_X1 U8852 ( .B1(n10097), .B2(n7159), .A(n7158), .ZN(n7160) );
  OAI21_X1 U8853 ( .B1(n10099), .B2(n8208), .A(n7160), .ZN(P2_U3286) );
  OR2_X1 U8854 ( .A1(n9100), .A2(n8646), .ZN(n7161) );
  AND2_X2 U8855 ( .A1(n7162), .A2(n7161), .ZN(n7163) );
  OR2_X1 U8856 ( .A1(n9099), .A2(n9882), .ZN(n8913) );
  NAND2_X1 U8857 ( .A1(n9099), .A2(n9882), .ZN(n8911) );
  NAND2_X1 U8858 ( .A1(n8913), .A2(n8911), .ZN(n9021) );
  OAI21_X1 U8859 ( .B1(n7163), .B2(n9021), .A(n7231), .ZN(n9880) );
  INV_X1 U8860 ( .A(n9098), .ZN(n7197) );
  INV_X1 U8861 ( .A(n9100), .ZN(n7165) );
  XNOR2_X1 U8862 ( .A(n7233), .B(n9021), .ZN(n7164) );
  OAI222_X1 U8863 ( .A1(n9422), .A2(n7197), .B1(n9424), .B2(n7165), .C1(n7164), 
        .C2(n9420), .ZN(n9885) );
  OAI21_X1 U8864 ( .B1(n4660), .B2(n9882), .A(n7237), .ZN(n9884) );
  OAI22_X1 U8865 ( .A1(n9425), .A2(n7167), .B1(n7193), .B2(n9407), .ZN(n7168)
         );
  AOI21_X1 U8866 ( .B1(n9367), .B2(n7229), .A(n7168), .ZN(n7169) );
  OAI21_X1 U8867 ( .B1(n9884), .B2(n7170), .A(n7169), .ZN(n7171) );
  AOI21_X1 U8868 ( .B1(n9885), .B2(n9425), .A(n7171), .ZN(n7172) );
  OAI21_X1 U8869 ( .B1(n9495), .B2(n9880), .A(n7172), .ZN(P1_U3283) );
  XNOR2_X1 U8870 ( .A(n7173), .B(n4599), .ZN(n7174) );
  NAND2_X1 U8871 ( .A1(n7174), .A2(n9489), .ZN(n7176) );
  AOI22_X1 U8872 ( .A1(n9486), .A2(n9103), .B1(n9101), .B2(n9484), .ZN(n7175)
         );
  NAND2_X1 U8873 ( .A1(n7176), .A2(n7175), .ZN(n9864) );
  AND2_X1 U8874 ( .A1(n9425), .A2(n9321), .ZN(n9412) );
  INV_X1 U8875 ( .A(n9412), .ZN(n7187) );
  AOI21_X1 U8876 ( .B1(n7177), .B2(n7184), .A(n9883), .ZN(n7179) );
  NAND2_X1 U8877 ( .A1(n7179), .A2(n7178), .ZN(n9862) );
  AOI21_X1 U8878 ( .B1(n8888), .B2(n7180), .A(n7038), .ZN(n9866) );
  NAND2_X1 U8879 ( .A1(n9866), .A2(n9366), .ZN(n7186) );
  OAI22_X1 U8880 ( .A1(n9425), .A2(n7182), .B1(n7181), .B2(n9407), .ZN(n7183)
         );
  AOI21_X1 U8881 ( .B1(n9367), .B2(n7184), .A(n7183), .ZN(n7185) );
  OAI211_X1 U8882 ( .C1(n7187), .C2(n9862), .A(n7186), .B(n7185), .ZN(n7188)
         );
  AOI21_X1 U8883 ( .B1(n9425), .B2(n9864), .A(n7188), .ZN(n7189) );
  INV_X1 U8884 ( .A(n7189), .ZN(P1_U3286) );
  NAND2_X1 U8885 ( .A1(n4466), .A2(n7190), .ZN(n7192) );
  XNOR2_X1 U8886 ( .A(n7192), .B(n7191), .ZN(n7200) );
  NOR2_X1 U8887 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8499), .ZN(n9773) );
  AOI21_X1 U8888 ( .B1(n8774), .B2(n9100), .A(n9773), .ZN(n7196) );
  INV_X1 U8889 ( .A(n7193), .ZN(n7194) );
  NAND2_X1 U8890 ( .A1(n8789), .A2(n7194), .ZN(n7195) );
  OAI211_X1 U8891 ( .C1(n7197), .C2(n8786), .A(n7196), .B(n7195), .ZN(n7198)
         );
  AOI21_X1 U8892 ( .B1(n8804), .B2(n7229), .A(n7198), .ZN(n7199) );
  OAI21_X1 U8893 ( .B1(n7200), .B2(n8806), .A(n7199), .ZN(P1_U3219) );
  INV_X1 U8894 ( .A(n7201), .ZN(n7203) );
  OAI222_X1 U8895 ( .A1(n8627), .A2(n7202), .B1(n7538), .B2(n7203), .C1(
        P2_U3152), .C2(n7725), .ZN(P2_U3336) );
  OAI222_X1 U8896 ( .A1(n9618), .A2(n7204), .B1(n7433), .B2(n7203), .C1(n6308), 
        .C2(P1_U3084), .ZN(P1_U3331) );
  INV_X1 U8897 ( .A(n9958), .ZN(n7960) );
  NAND2_X1 U8898 ( .A1(n9916), .A2(n7960), .ZN(n7206) );
  OR2_X1 U8899 ( .A1(n9956), .A2(n7324), .ZN(n7793) );
  NAND2_X1 U8900 ( .A1(n9956), .A2(n7324), .ZN(n7785) );
  NAND2_X1 U8901 ( .A1(n7793), .A2(n7785), .ZN(n7903) );
  OAI21_X1 U8902 ( .B1(n7208), .B2(n7903), .A(n7313), .ZN(n10100) );
  INV_X1 U8903 ( .A(n7211), .ZN(n7213) );
  INV_X1 U8904 ( .A(n7903), .ZN(n7210) );
  NAND2_X1 U8905 ( .A1(n7211), .A2(n7210), .ZN(n7302) );
  INV_X1 U8906 ( .A(n7302), .ZN(n7212) );
  AOI21_X1 U8907 ( .B1(n7213), .B2(n7903), .A(n7212), .ZN(n7214) );
  OAI222_X1 U8908 ( .A1(n8241), .A2(n9958), .B1(n9995), .B2(n9953), .C1(n8226), 
        .C2(n7214), .ZN(n10104) );
  INV_X1 U8909 ( .A(n9956), .ZN(n10101) );
  OAI21_X1 U8910 ( .B1(n7215), .B2(n10101), .A(n7308), .ZN(n10103) );
  OAI22_X1 U8911 ( .A1(n10035), .A2(n7216), .B1(n9965), .B2(n10028), .ZN(n7217) );
  AOI21_X1 U8912 ( .B1(n8071), .B2(n9956), .A(n7217), .ZN(n7218) );
  OAI21_X1 U8913 ( .B1(n10103), .B2(n9986), .A(n7218), .ZN(n7219) );
  AOI21_X1 U8914 ( .B1(n10104), .B2(n10035), .A(n7219), .ZN(n7220) );
  OAI21_X1 U8915 ( .B1(n8232), .B2(n10100), .A(n7220), .ZN(P2_U3285) );
  AOI21_X1 U8916 ( .B1(n7222), .B2(n7221), .A(n4469), .ZN(n7228) );
  NOR2_X1 U8917 ( .A1(n8798), .A2(n7236), .ZN(n7223) );
  AOI211_X1 U8918 ( .C1(n8800), .C2(n9097), .A(n7224), .B(n7223), .ZN(n7225)
         );
  OAI21_X1 U8919 ( .B1(n7239), .B2(n8802), .A(n7225), .ZN(n7226) );
  AOI21_X1 U8920 ( .B1(n8804), .B2(n9891), .A(n7226), .ZN(n7227) );
  OAI21_X1 U8921 ( .B1(n7228), .B2(n8806), .A(n7227), .ZN(P1_U3229) );
  NAND2_X1 U8922 ( .A1(n9099), .A2(n7229), .ZN(n7230) );
  INV_X1 U8923 ( .A(n9891), .ZN(n7238) );
  OR2_X1 U8924 ( .A1(n9098), .A2(n7238), .ZN(n8914) );
  NAND2_X1 U8925 ( .A1(n9098), .A2(n7238), .ZN(n8916) );
  NAND2_X1 U8926 ( .A1(n8914), .A2(n8916), .ZN(n9022) );
  XNOR2_X1 U8927 ( .A(n7339), .B(n9022), .ZN(n9895) );
  INV_X1 U8928 ( .A(n9097), .ZN(n7396) );
  INV_X1 U8929 ( .A(n8913), .ZN(n7232) );
  NAND2_X1 U8930 ( .A1(n7341), .A2(n8911), .ZN(n7234) );
  XOR2_X1 U8931 ( .A(n9022), .B(n7234), .Z(n7235) );
  OAI222_X1 U8932 ( .A1(n9422), .A2(n7396), .B1(n9424), .B2(n7236), .C1(n9420), 
        .C2(n7235), .ZN(n9897) );
  NAND2_X1 U8933 ( .A1(n9897), .A2(n9425), .ZN(n7243) );
  AOI211_X1 U8934 ( .C1(n9891), .C2(n7237), .A(n9883), .B(n7343), .ZN(n9890)
         );
  NOR2_X1 U8935 ( .A1(n9480), .A2(n7238), .ZN(n7241) );
  OAI22_X1 U8936 ( .A1(n9425), .A2(n6356), .B1(n7239), .B2(n9407), .ZN(n7240)
         );
  AOI211_X1 U8937 ( .C1(n9890), .C2(n9412), .A(n7241), .B(n7240), .ZN(n7242)
         );
  OAI211_X1 U8938 ( .C1(n9495), .C2(n9895), .A(n7243), .B(n7242), .ZN(P1_U3282) );
  NOR2_X1 U8939 ( .A1(n7245), .A2(n7244), .ZN(n7286) );
  XNOR2_X1 U8940 ( .A(n7287), .B(n7286), .ZN(n7246) );
  NOR2_X1 U8941 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n7246), .ZN(n7288) );
  AOI21_X1 U8942 ( .B1(n7246), .B2(P2_REG2_REG_15__SCAN_IN), .A(n7288), .ZN(
        n7253) );
  AND2_X1 U8943 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(P2_U3152), .ZN(n7718) );
  OAI21_X1 U8944 ( .B1(P2_REG1_REG_14__SCAN_IN), .B2(n7248), .A(n7247), .ZN(
        n7277) );
  XNOR2_X1 U8945 ( .A(n7277), .B(n7278), .ZN(n7249) );
  NOR2_X1 U8946 ( .A1(n5384), .A2(n7249), .ZN(n7279) );
  AOI211_X1 U8947 ( .C1(n5384), .C2(n7249), .A(n7279), .B(n9972), .ZN(n7250)
         );
  AOI211_X1 U8948 ( .C1(P2_ADDR_REG_15__SCAN_IN), .C2(n9969), .A(n7718), .B(
        n7250), .ZN(n7252) );
  NAND2_X1 U8949 ( .A1(n9659), .A2(n7287), .ZN(n7251) );
  OAI211_X1 U8950 ( .C1(n7253), .C2(n9970), .A(n7252), .B(n7251), .ZN(P2_U3260) );
  INV_X1 U8951 ( .A(n7273), .ZN(n7255) );
  NAND2_X1 U8952 ( .A1(n8633), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n7254) );
  OAI211_X1 U8953 ( .C1(n7255), .C2(n8635), .A(n7946), .B(n7254), .ZN(P2_U3335) );
  NAND2_X1 U8954 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n9115), .ZN(n7256) );
  OAI21_X1 U8955 ( .B1(n9115), .B2(P1_REG2_REG_12__SCAN_IN), .A(n7256), .ZN(
        n9112) );
  OAI21_X1 U8956 ( .B1(n7267), .B2(P1_REG2_REG_11__SCAN_IN), .A(n7257), .ZN(
        n9113) );
  NOR2_X1 U8957 ( .A1(n9112), .A2(n9113), .ZN(n9111) );
  MUX2_X1 U8958 ( .A(P1_REG2_REG_13__SCAN_IN), .B(n6029), .S(n9128), .Z(n7258)
         );
  INV_X1 U8959 ( .A(n7258), .ZN(n9125) );
  NOR2_X1 U8960 ( .A1(n7259), .A2(n7263), .ZN(n7261) );
  XNOR2_X1 U8961 ( .A(n9796), .B(n7260), .ZN(n9792) );
  NOR2_X1 U8962 ( .A1(n7466), .A2(n9792), .ZN(n9793) );
  NOR2_X1 U8963 ( .A1(n7261), .A2(n9793), .ZN(n9133) );
  XNOR2_X1 U8964 ( .A(n9133), .B(n9141), .ZN(n7262) );
  NOR2_X1 U8965 ( .A1(n6068), .A2(n7262), .ZN(n9134) );
  AOI211_X1 U8966 ( .C1(n7262), .C2(n6068), .A(n9134), .B(n9819), .ZN(n7272)
         );
  AOI22_X1 U8967 ( .A1(n9796), .A2(P1_REG1_REG_14__SCAN_IN), .B1(n6046), .B2(
        n7263), .ZN(n9803) );
  MUX2_X1 U8968 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n7264), .S(n9128), .Z(n9121)
         );
  AOI22_X1 U8969 ( .A1(P1_REG1_REG_12__SCAN_IN), .A2(n9115), .B1(n7265), .B2(
        n6006), .ZN(n9108) );
  OAI21_X1 U8970 ( .B1(P1_REG1_REG_11__SCAN_IN), .B2(n7267), .A(n7266), .ZN(
        n9109) );
  NAND2_X1 U8971 ( .A1(n9108), .A2(n9109), .ZN(n9107) );
  OAI21_X1 U8972 ( .B1(P1_REG1_REG_12__SCAN_IN), .B2(n9115), .A(n9107), .ZN(
        n9122) );
  NAND2_X1 U8973 ( .A1(n9121), .A2(n9122), .ZN(n9120) );
  OAI21_X1 U8974 ( .B1(P1_REG1_REG_13__SCAN_IN), .B2(n9128), .A(n9120), .ZN(
        n9804) );
  NAND2_X1 U8975 ( .A1(n9803), .A2(n9804), .ZN(n9802) );
  OAI21_X1 U8976 ( .B1(n9796), .B2(P1_REG1_REG_14__SCAN_IN), .A(n9802), .ZN(
        n9140) );
  XNOR2_X1 U8977 ( .A(n9140), .B(n9141), .ZN(n7268) );
  NOR2_X1 U8978 ( .A1(n6067), .A2(n7268), .ZN(n9142) );
  AOI211_X1 U8979 ( .C1(n7268), .C2(n6067), .A(n9142), .B(n9769), .ZN(n7271)
         );
  NAND2_X1 U8980 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n8797) );
  NAND2_X1 U8981 ( .A1(n9778), .A2(P1_ADDR_REG_15__SCAN_IN), .ZN(n7269) );
  OAI211_X1 U8982 ( .C1(n9149), .C2(n9141), .A(n8797), .B(n7269), .ZN(n7270)
         );
  OR3_X1 U8983 ( .A1(n7272), .A2(n7271), .A3(n7270), .ZN(P1_U3256) );
  NAND2_X1 U8984 ( .A1(n7273), .A2(n9622), .ZN(n7275) );
  OR2_X1 U8985 ( .A1(n7274), .A2(P1_U3084), .ZN(n9090) );
  OAI211_X1 U8986 ( .C1(n7276), .C2(n9618), .A(n7275), .B(n9090), .ZN(P1_U3330) );
  NOR2_X1 U8987 ( .A1(n7278), .A2(n7277), .ZN(n7280) );
  NOR2_X1 U8988 ( .A1(n7280), .A2(n7279), .ZN(n7283) );
  XNOR2_X1 U8989 ( .A(n7985), .B(n7281), .ZN(n7282) );
  NAND2_X1 U8990 ( .A1(n7282), .A2(n7283), .ZN(n7984) );
  OAI21_X1 U8991 ( .B1(n7283), .B2(n7282), .A(n7984), .ZN(n7284) );
  INV_X1 U8992 ( .A(n7284), .ZN(n7296) );
  AND2_X1 U8993 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3152), .ZN(n7648) );
  NOR2_X1 U8994 ( .A1(n9971), .A2(n7291), .ZN(n7285) );
  AOI211_X1 U8995 ( .C1(P2_ADDR_REG_16__SCAN_IN), .C2(n9969), .A(n7648), .B(
        n7285), .ZN(n7295) );
  NOR2_X1 U8996 ( .A1(n7287), .A2(n7286), .ZN(n7289) );
  NOR2_X1 U8997 ( .A1(n7289), .A2(n7288), .ZN(n7293) );
  NAND2_X1 U8998 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n7985), .ZN(n7981) );
  INV_X1 U8999 ( .A(n7981), .ZN(n7290) );
  AOI21_X1 U9000 ( .B1(n5405), .B2(n7291), .A(n7290), .ZN(n7292) );
  NAND2_X1 U9001 ( .A1(n7292), .A2(n7293), .ZN(n7980) );
  OAI211_X1 U9002 ( .C1(n7293), .C2(n7292), .A(n9968), .B(n7980), .ZN(n7294)
         );
  OAI211_X1 U9003 ( .C1(n7296), .C2(n9972), .A(n7295), .B(n7294), .ZN(P2_U3261) );
  INV_X1 U9004 ( .A(n7297), .ZN(n7300) );
  OAI222_X1 U9005 ( .A1(n7433), .A2(n7300), .B1(P1_U3084), .B2(n7298), .C1(
        n8411), .C2(n9618), .ZN(P1_U3329) );
  OAI222_X1 U9006 ( .A1(P2_U3152), .A2(n7301), .B1(n8635), .B2(n7300), .C1(
        n7299), .C2(n8627), .ZN(P2_U3334) );
  NAND2_X1 U9007 ( .A1(n7414), .A2(n9953), .ZN(n7796) );
  AND2_X1 U9008 ( .A1(n7796), .A2(n7785), .ZN(n7791) );
  INV_X1 U9009 ( .A(n7419), .ZN(n7304) );
  AOI21_X1 U9010 ( .B1(n7302), .B2(n7785), .A(n7906), .ZN(n7303) );
  AOI211_X1 U9011 ( .C1(n7304), .C2(n7794), .A(n8226), .B(n7303), .ZN(n7306)
         );
  OAI22_X1 U9012 ( .A1(n7324), .A2(n8241), .B1(n7479), .B2(n9995), .ZN(n7305)
         );
  NOR2_X1 U9013 ( .A1(n7306), .A2(n7305), .ZN(n10109) );
  OAI22_X1 U9014 ( .A1(n10035), .A2(n7307), .B1(n7323), .B2(n10028), .ZN(n7311) );
  INV_X1 U9015 ( .A(n7308), .ZN(n7309) );
  INV_X1 U9016 ( .A(n7414), .ZN(n10111) );
  OAI211_X1 U9017 ( .C1(n7309), .C2(n10111), .A(n10022), .B(n7425), .ZN(n10108) );
  NOR2_X1 U9018 ( .A1(n10108), .A2(n7503), .ZN(n7310) );
  AOI211_X1 U9019 ( .C1(n8071), .C2(n7414), .A(n7311), .B(n7310), .ZN(n7317)
         );
  INV_X1 U9020 ( .A(n7324), .ZN(n9914) );
  NAND2_X1 U9021 ( .A1(n9956), .A2(n9914), .ZN(n7312) );
  INV_X1 U9022 ( .A(n7906), .ZN(n7314) );
  OAI21_X1 U9023 ( .B1(n7315), .B2(n7314), .A(n7416), .ZN(n10113) );
  NAND2_X1 U9024 ( .A1(n10113), .A2(n7500), .ZN(n7316) );
  OAI211_X1 U9025 ( .C1(n10109), .C2(n8208), .A(n7317), .B(n7316), .ZN(
        P2_U3284) );
  NAND2_X1 U9026 ( .A1(n7319), .A2(n7318), .ZN(n7321) );
  XOR2_X1 U9027 ( .A(n7321), .B(n7320), .Z(n7328) );
  OAI21_X1 U9028 ( .B1(n9966), .B2(n7323), .A(n7322), .ZN(n7326) );
  OAI22_X1 U9029 ( .A1(n7324), .A2(n9959), .B1(n9954), .B2(n7479), .ZN(n7325)
         );
  AOI211_X1 U9030 ( .C1(n9957), .C2(n7414), .A(n7326), .B(n7325), .ZN(n7327)
         );
  OAI21_X1 U9031 ( .B1(n7328), .B2(n7709), .A(n7327), .ZN(P2_U3226) );
  AOI21_X1 U9032 ( .B1(n7330), .B2(n7329), .A(n7389), .ZN(n7337) );
  NOR2_X1 U9033 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7331), .ZN(n9788) );
  AOI21_X1 U9034 ( .B1(n8774), .B2(n9098), .A(n9788), .ZN(n7334) );
  INV_X1 U9035 ( .A(n7332), .ZN(n7378) );
  NAND2_X1 U9036 ( .A1(n8789), .A2(n7378), .ZN(n7333) );
  OAI211_X1 U9037 ( .C1(n7411), .C2(n8786), .A(n7334), .B(n7333), .ZN(n7335)
         );
  AOI21_X1 U9038 ( .B1(n8804), .B2(n7351), .A(n7335), .ZN(n7336) );
  OAI21_X1 U9039 ( .B1(n7337), .B2(n8806), .A(n7336), .ZN(P1_U3215) );
  OR2_X1 U9040 ( .A1(n9098), .A2(n9891), .ZN(n7338) );
  OR2_X1 U9041 ( .A1(n9097), .A2(n7380), .ZN(n8921) );
  NAND2_X1 U9042 ( .A1(n7380), .A2(n9097), .ZN(n8917) );
  NAND2_X1 U9043 ( .A1(n8921), .A2(n8917), .ZN(n9023) );
  INV_X1 U9044 ( .A(n9023), .ZN(n7355) );
  XNOR2_X1 U9045 ( .A(n7352), .B(n7355), .ZN(n7386) );
  AND2_X1 U9046 ( .A1(n8911), .A2(n8916), .ZN(n8909) );
  XNOR2_X1 U9047 ( .A(n7356), .B(n7355), .ZN(n7342) );
  AOI222_X1 U9048 ( .A1(n9489), .A2(n7342), .B1(n9098), .B2(n9486), .C1(n9096), 
        .C2(n9484), .ZN(n7381) );
  INV_X1 U9049 ( .A(n7343), .ZN(n7345) );
  NAND2_X1 U9050 ( .A1(n7343), .A2(n7380), .ZN(n7363) );
  INV_X1 U9051 ( .A(n7363), .ZN(n7344) );
  AOI211_X1 U9052 ( .C1(n7351), .C2(n7345), .A(n9883), .B(n7344), .ZN(n7384)
         );
  AOI21_X1 U9053 ( .B1(n9892), .B2(n7351), .A(n7384), .ZN(n7346) );
  OAI211_X1 U9054 ( .C1(n7386), .C2(n9894), .A(n7381), .B(n7346), .ZN(n7348)
         );
  NAND2_X1 U9055 ( .A1(n7348), .A2(n9910), .ZN(n7347) );
  OAI21_X1 U9056 ( .B1(n9910), .B2(n6595), .A(n7347), .ZN(P1_U3533) );
  INV_X1 U9057 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n7350) );
  NAND2_X1 U9058 ( .A1(n7348), .A2(n9900), .ZN(n7349) );
  OAI21_X1 U9059 ( .B1(n9900), .B2(n7350), .A(n7349), .ZN(P1_U3484) );
  XNOR2_X1 U9060 ( .A(n9589), .B(n7411), .ZN(n9026) );
  XNOR2_X1 U9061 ( .A(n7400), .B(n8920), .ZN(n7354) );
  INV_X1 U9062 ( .A(n7354), .ZN(n9593) );
  NAND2_X1 U9063 ( .A1(n7354), .A2(n7353), .ZN(n7362) );
  NAND2_X1 U9064 ( .A1(n7356), .A2(n7355), .ZN(n7357) );
  NAND2_X1 U9065 ( .A1(n8921), .A2(n8914), .ZN(n8908) );
  NAND2_X1 U9066 ( .A1(n8908), .A2(n8917), .ZN(n8829) );
  XNOR2_X1 U9067 ( .A(n7408), .B(n8920), .ZN(n7360) );
  NAND2_X1 U9068 ( .A1(n9097), .A2(n9486), .ZN(n7358) );
  OAI21_X1 U9069 ( .B1(n7402), .B2(n9422), .A(n7358), .ZN(n7359) );
  AOI21_X1 U9070 ( .B1(n7360), .B2(n9489), .A(n7359), .ZN(n7361) );
  NAND2_X1 U9071 ( .A1(n7362), .A2(n7361), .ZN(n9595) );
  NAND2_X1 U9072 ( .A1(n9595), .A2(n9425), .ZN(n7369) );
  NAND2_X1 U9073 ( .A1(n7363), .A2(n9589), .ZN(n7364) );
  AND2_X1 U9074 ( .A1(n7403), .A2(n7364), .ZN(n9591) );
  INV_X1 U9075 ( .A(n9589), .ZN(n7401) );
  NOR2_X1 U9076 ( .A1(n9480), .A2(n7401), .ZN(n7367) );
  OAI22_X1 U9077 ( .A1(n9425), .A2(n7365), .B1(n7392), .B2(n9407), .ZN(n7366)
         );
  AOI211_X1 U9078 ( .C1(n9591), .C2(n9493), .A(n7367), .B(n7366), .ZN(n7368)
         );
  OAI211_X1 U9079 ( .C1(n9593), .C2(n7370), .A(n7369), .B(n7368), .ZN(P1_U3280) );
  XNOR2_X1 U9080 ( .A(n7371), .B(n7372), .ZN(n7377) );
  OAI21_X1 U9081 ( .B1(n9966), .B2(n7423), .A(n7373), .ZN(n7375) );
  OAI22_X1 U9082 ( .A1(n9953), .A2(n9959), .B1(n9954), .B2(n7716), .ZN(n7374)
         );
  AOI211_X1 U9083 ( .C1(n9957), .C2(n9706), .A(n7375), .B(n7374), .ZN(n7376)
         );
  OAI21_X1 U9084 ( .B1(n7377), .B2(n7709), .A(n7376), .ZN(P2_U3236) );
  AOI22_X1 U9085 ( .A1(n9447), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n7378), .B2(
        n9477), .ZN(n7379) );
  OAI21_X1 U9086 ( .B1(n7380), .B2(n9480), .A(n7379), .ZN(n7383) );
  NOR2_X1 U9087 ( .A1(n7381), .A2(n9490), .ZN(n7382) );
  AOI211_X1 U9088 ( .C1(n7384), .C2(n9457), .A(n7383), .B(n7382), .ZN(n7385)
         );
  OAI21_X1 U9089 ( .B1(n9495), .B2(n7386), .A(n7385), .ZN(P1_U3281) );
  OAI21_X1 U9090 ( .B1(n7389), .B2(n7388), .A(n7387), .ZN(n7390) );
  NAND3_X1 U9091 ( .A1(n4583), .A2(n8783), .A3(n7390), .ZN(n7399) );
  AOI21_X1 U9092 ( .B1(n8800), .B2(n9487), .A(n7391), .ZN(n7395) );
  INV_X1 U9093 ( .A(n7392), .ZN(n7393) );
  NAND2_X1 U9094 ( .A1(n8789), .A2(n7393), .ZN(n7394) );
  OAI211_X1 U9095 ( .C1(n7396), .C2(n8798), .A(n7395), .B(n7394), .ZN(n7397)
         );
  INV_X1 U9096 ( .A(n7397), .ZN(n7398) );
  OAI211_X1 U9097 ( .C1(n7401), .C2(n8792), .A(n7399), .B(n7398), .ZN(P1_U3234) );
  NAND2_X1 U9098 ( .A1(n9586), .A2(n7402), .ZN(n8922) );
  NAND2_X1 U9099 ( .A1(n8929), .A2(n8922), .ZN(n9025) );
  XNOR2_X1 U9100 ( .A(n7457), .B(n9025), .ZN(n9588) );
  AOI211_X1 U9101 ( .C1(n9586), .C2(n7403), .A(n9883), .B(n9473), .ZN(n9585)
         );
  INV_X1 U9102 ( .A(n9586), .ZN(n7404) );
  NOR2_X1 U9103 ( .A1(n9480), .A2(n7404), .ZN(n7407) );
  OAI22_X1 U9104 ( .A1(n9425), .A2(n7405), .B1(n8725), .B2(n9407), .ZN(n7406)
         );
  AOI211_X1 U9105 ( .C1(n9585), .C2(n9457), .A(n7407), .B(n7406), .ZN(n7413)
         );
  INV_X1 U9106 ( .A(n9095), .ZN(n8842) );
  AND2_X1 U9107 ( .A1(n9589), .A2(n7411), .ZN(n8827) );
  OR2_X1 U9108 ( .A1(n9589), .A2(n7411), .ZN(n7459) );
  NAND2_X1 U9109 ( .A1(n7460), .A2(n7459), .ZN(n7409) );
  XOR2_X1 U9110 ( .A(n9025), .B(n7409), .Z(n7410) );
  OAI222_X1 U9111 ( .A1(n9424), .A2(n7411), .B1(n9422), .B2(n8842), .C1(n9420), 
        .C2(n7410), .ZN(n9584) );
  NAND2_X1 U9112 ( .A1(n9584), .A2(n9425), .ZN(n7412) );
  OAI211_X1 U9113 ( .C1(n9588), .C2(n9495), .A(n7413), .B(n7412), .ZN(P1_U3279) );
  INV_X1 U9114 ( .A(n9953), .ZN(n7959) );
  OR2_X1 U9115 ( .A1(n7414), .A2(n7959), .ZN(n7415) );
  OR2_X1 U9116 ( .A1(n9706), .A2(n7479), .ZN(n7802) );
  NAND2_X1 U9117 ( .A1(n9706), .A2(n7479), .ZN(n7443) );
  NAND2_X1 U9118 ( .A1(n7417), .A2(n7907), .ZN(n7418) );
  NAND2_X1 U9119 ( .A1(n4935), .A2(n7418), .ZN(n9705) );
  OAI21_X1 U9120 ( .B1(n4457), .B2(n7907), .A(n7444), .ZN(n7421) );
  OAI22_X1 U9121 ( .A1(n9953), .A2(n8241), .B1(n7716), .B2(n9995), .ZN(n7420)
         );
  AOI21_X1 U9122 ( .B1(n7421), .B2(n10012), .A(n7420), .ZN(n7422) );
  OAI21_X1 U9123 ( .B1(n9705), .B2(n9989), .A(n7422), .ZN(n9708) );
  NAND2_X1 U9124 ( .A1(n9708), .A2(n10035), .ZN(n7430) );
  OAI22_X1 U9125 ( .A1(n10035), .A2(n7424), .B1(n7423), .B2(n10028), .ZN(n7428) );
  AND2_X1 U9126 ( .A1(n7425), .A2(n9706), .ZN(n7426) );
  OR2_X1 U9127 ( .A1(n7426), .A2(n4465), .ZN(n9707) );
  NOR2_X1 U9128 ( .A1(n9707), .A2(n9986), .ZN(n7427) );
  AOI211_X1 U9129 ( .C1(n8071), .C2(n9706), .A(n7428), .B(n7427), .ZN(n7429)
         );
  OAI211_X1 U9130 ( .C1(n9705), .C2(n9987), .A(n7430), .B(n7429), .ZN(P2_U3283) );
  INV_X1 U9131 ( .A(n7431), .ZN(n7436) );
  OAI222_X1 U9132 ( .A1(n9618), .A2(n7434), .B1(n7433), .B2(n7436), .C1(n7432), 
        .C2(P1_U3084), .ZN(P1_U3328) );
  OAI222_X1 U9133 ( .A1(n8627), .A2(n7437), .B1(n7538), .B2(n7436), .C1(
        P2_U3152), .C2(n7435), .ZN(P2_U3333) );
  INV_X1 U9134 ( .A(n7438), .ZN(n7455) );
  OAI222_X1 U9135 ( .A1(n7433), .A2(n7455), .B1(P1_U3084), .B2(n7440), .C1(
        n7439), .C2(n9618), .ZN(P1_U3327) );
  INV_X1 U9136 ( .A(n7479), .ZN(n7958) );
  NAND2_X1 U9137 ( .A1(n7497), .A2(n7716), .ZN(n7801) );
  NAND2_X1 U9138 ( .A1(n7798), .A2(n7801), .ZN(n7442) );
  OAI21_X1 U9139 ( .B1(n4462), .B2(n7442), .A(n7499), .ZN(n9704) );
  INV_X1 U9140 ( .A(n9704), .ZN(n7454) );
  INV_X1 U9141 ( .A(n7443), .ZN(n7441) );
  NOR2_X1 U9142 ( .A1(n7442), .A2(n7441), .ZN(n7799) );
  NAND2_X1 U9143 ( .A1(n7495), .A2(n10012), .ZN(n7447) );
  INV_X1 U9144 ( .A(n7442), .ZN(n7908) );
  AOI21_X1 U9145 ( .B1(n7444), .B2(n7443), .A(n7908), .ZN(n7446) );
  INV_X1 U9146 ( .A(n8242), .ZN(n7956) );
  AOI22_X1 U9147 ( .A1(n9935), .A2(n7956), .B1(n7958), .B2(n9992), .ZN(n7445)
         );
  OAI21_X1 U9148 ( .B1(n7447), .B2(n7446), .A(n7445), .ZN(n9703) );
  INV_X1 U9149 ( .A(n7497), .ZN(n9700) );
  INV_X1 U9150 ( .A(n7502), .ZN(n7448) );
  OAI21_X1 U9151 ( .B1(n9700), .B2(n4465), .A(n7448), .ZN(n9701) );
  OAI22_X1 U9152 ( .A1(n10035), .A2(n7449), .B1(n7478), .B2(n10028), .ZN(n7450) );
  AOI21_X1 U9153 ( .B1(n7497), .B2(n8071), .A(n7450), .ZN(n7451) );
  OAI21_X1 U9154 ( .B1(n9701), .B2(n9986), .A(n7451), .ZN(n7452) );
  AOI21_X1 U9155 ( .B1(n9703), .B2(n10035), .A(n7452), .ZN(n7453) );
  OAI21_X1 U9156 ( .B1(n7454), .B2(n8232), .A(n7453), .ZN(P2_U3282) );
  OAI222_X1 U9157 ( .A1(P2_U3152), .A2(n7456), .B1(n8635), .B2(n7455), .C1(
        n8409), .C2(n8627), .ZN(P2_U3332) );
  AOI22_X2 U9158 ( .A1(n7457), .A2(n9025), .B1(n9487), .B2(n9586), .ZN(n9472)
         );
  NAND2_X1 U9159 ( .A1(n9579), .A2(n9095), .ZN(n7458) );
  INV_X1 U9160 ( .A(n9579), .ZN(n9481) );
  NAND2_X1 U9161 ( .A1(n9199), .A2(n9200), .ZN(n8843) );
  NAND2_X1 U9162 ( .A1(n9223), .A2(n8843), .ZN(n9027) );
  XOR2_X1 U9163 ( .A(n9198), .B(n9027), .Z(n9719) );
  INV_X1 U9164 ( .A(n9719), .ZN(n7472) );
  XNOR2_X1 U9165 ( .A(n9579), .B(n9095), .ZN(n9482) );
  NAND2_X1 U9166 ( .A1(n9483), .A2(n9482), .ZN(n7461) );
  NAND2_X1 U9167 ( .A1(n9579), .A2(n8842), .ZN(n8826) );
  NAND2_X1 U9168 ( .A1(n7462), .A2(n9027), .ZN(n7463) );
  NAND3_X1 U9169 ( .A1(n9224), .A2(n9489), .A3(n7463), .ZN(n7465) );
  AOI22_X1 U9170 ( .A1(n9486), .A2(n9095), .B1(n9452), .B2(n9484), .ZN(n7464)
         );
  NAND2_X1 U9171 ( .A1(n7465), .A2(n7464), .ZN(n9718) );
  OAI211_X1 U9172 ( .C1(n9474), .C2(n4758), .A(n9590), .B(n9460), .ZN(n9716)
         );
  OAI22_X1 U9173 ( .A1(n9425), .A2(n7466), .B1(n8658), .B2(n9407), .ZN(n7467)
         );
  AOI21_X1 U9174 ( .B1(n9199), .B2(n9367), .A(n7467), .ZN(n7468) );
  OAI21_X1 U9175 ( .B1(n9716), .B2(n7469), .A(n7468), .ZN(n7470) );
  AOI21_X1 U9176 ( .B1(n9718), .B2(n9425), .A(n7470), .ZN(n7471) );
  OAI21_X1 U9177 ( .B1(n7472), .B2(n9495), .A(n7471), .ZN(P1_U3277) );
  INV_X1 U9178 ( .A(n7473), .ZN(n7474) );
  AOI21_X1 U9179 ( .B1(n7476), .B2(n7475), .A(n7474), .ZN(n7483) );
  OAI21_X1 U9180 ( .B1(n9966), .B2(n7478), .A(n7477), .ZN(n7481) );
  OAI22_X1 U9181 ( .A1(n8242), .A2(n9954), .B1(n9959), .B2(n7479), .ZN(n7480)
         );
  AOI211_X1 U9182 ( .C1(n9957), .C2(n7497), .A(n7481), .B(n7480), .ZN(n7482)
         );
  OAI21_X1 U9183 ( .B1(n7483), .B2(n7709), .A(n7482), .ZN(P2_U3217) );
  INV_X1 U9184 ( .A(n7484), .ZN(n7486) );
  NOR2_X1 U9185 ( .A1(n7486), .A2(n7485), .ZN(n7487) );
  XNOR2_X1 U9186 ( .A(n7488), .B(n7487), .ZN(n7494) );
  NAND2_X1 U9187 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9131) );
  INV_X1 U9188 ( .A(n9131), .ZN(n7490) );
  NOR2_X1 U9189 ( .A1(n8786), .A2(n9200), .ZN(n7489) );
  AOI211_X1 U9190 ( .C1(n8774), .C2(n9487), .A(n7490), .B(n7489), .ZN(n7491)
         );
  OAI21_X1 U9191 ( .B1(n9476), .B2(n8802), .A(n7491), .ZN(n7492) );
  AOI21_X1 U9192 ( .B1(n8804), .B2(n9579), .A(n7492), .ZN(n7493) );
  OAI21_X1 U9193 ( .B1(n7494), .B2(n8806), .A(n7493), .ZN(P1_U3232) );
  NAND2_X1 U9194 ( .A1(n7568), .A2(n8242), .ZN(n7808) );
  NAND2_X1 U9195 ( .A1(n7807), .A2(n7808), .ZN(n7910) );
  XNOR2_X1 U9196 ( .A(n7586), .B(n7910), .ZN(n7496) );
  INV_X1 U9197 ( .A(n7716), .ZN(n7957) );
  INV_X1 U9198 ( .A(n8228), .ZN(n7955) );
  AOI222_X1 U9199 ( .A1(n10012), .A2(n7496), .B1(n7957), .B2(n9992), .C1(n7955), .C2(n9935), .ZN(n9696) );
  OR2_X1 U9200 ( .A1(n7497), .A2(n7957), .ZN(n7498) );
  XNOR2_X1 U9201 ( .A(n7570), .B(n7910), .ZN(n9699) );
  NAND2_X1 U9202 ( .A1(n9699), .A2(n7500), .ZN(n7507) );
  INV_X1 U9203 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n7501) );
  OAI22_X1 U9204 ( .A1(n10035), .A2(n7501), .B1(n7715), .B2(n10028), .ZN(n7505) );
  NAND2_X1 U9205 ( .A1(n7502), .A2(n9697), .ZN(n8246) );
  OAI211_X1 U9206 ( .C1(n7502), .C2(n9697), .A(n10022), .B(n8246), .ZN(n9695)
         );
  NOR2_X1 U9207 ( .A1(n9695), .A2(n7503), .ZN(n7504) );
  AOI211_X1 U9208 ( .C1(n8071), .C2(n7568), .A(n7505), .B(n7504), .ZN(n7506)
         );
  OAI211_X1 U9209 ( .C1(n8208), .C2(n9696), .A(n7507), .B(n7506), .ZN(P2_U3281) );
  INV_X1 U9210 ( .A(n7508), .ZN(n7509) );
  OAI222_X1 U9211 ( .A1(n7433), .A2(n7509), .B1(n9723), .B2(P1_U3084), .C1(
        n8476), .C2(n9618), .ZN(P1_U3326) );
  OAI222_X1 U9212 ( .A1(n8627), .A2(n7510), .B1(n8635), .B2(n7509), .C1(n7599), 
        .C2(P2_U3152), .ZN(P2_U3331) );
  INV_X1 U9213 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n7525) );
  INV_X1 U9214 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n8868) );
  MUX2_X1 U9215 ( .A(n7525), .B(n8868), .S(n7515), .Z(n7517) );
  INV_X1 U9216 ( .A(SI_29_), .ZN(n7516) );
  NAND2_X1 U9217 ( .A1(n7517), .A2(n7516), .ZN(n7520) );
  INV_X1 U9218 ( .A(n7517), .ZN(n7518) );
  NAND2_X1 U9219 ( .A1(n7518), .A2(SI_29_), .ZN(n7519) );
  NAND2_X1 U9220 ( .A1(n7524), .A2(n7523), .ZN(n7521) );
  INV_X1 U9221 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8811) );
  INV_X1 U9222 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n7866) );
  MUX2_X1 U9223 ( .A(n8811), .B(n7866), .S(n4478), .Z(n7871) );
  INV_X1 U9224 ( .A(n8810), .ZN(n7567) );
  OAI222_X1 U9225 ( .A1(n7433), .A2(n7567), .B1(n7522), .B2(P1_U3084), .C1(
        n8811), .C2(n9618), .ZN(P1_U3323) );
  INV_X1 U9226 ( .A(n8867), .ZN(n7566) );
  OAI222_X1 U9227 ( .A1(n7526), .A2(P2_U3152), .B1(n8635), .B2(n7566), .C1(
        n7525), .C2(n8627), .ZN(P2_U3329) );
  INV_X1 U9228 ( .A(n9954), .ZN(n9915) );
  AOI22_X1 U9229 ( .A1(n9918), .A2(n6764), .B1(n9915), .B2(n7965), .ZN(n7534)
         );
  OAI21_X1 U9230 ( .B1(n7529), .B2(n7528), .A(n7527), .ZN(n7532) );
  NAND2_X1 U9231 ( .A1(n7531), .A2(n7530), .ZN(n7685) );
  AOI22_X1 U9232 ( .A1(n9949), .A2(n7532), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n7685), .ZN(n7533) );
  OAI211_X1 U9233 ( .C1(n10055), .C2(n7723), .A(n7534), .B(n7533), .ZN(
        P2_U3224) );
  OAI222_X1 U9234 ( .A1(n8627), .A2(n8578), .B1(n7538), .B2(n7537), .C1(n7536), 
        .C2(P2_U3152), .ZN(P2_U3338) );
  XNOR2_X1 U9235 ( .A(n7541), .B(n7540), .ZN(n7542) );
  XNOR2_X1 U9236 ( .A(n7539), .B(n7542), .ZN(n7547) );
  NAND2_X1 U9237 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9816) );
  OAI21_X1 U9238 ( .B1(n8786), .B2(n9421), .A(n9816), .ZN(n7543) );
  AOI21_X1 U9239 ( .B1(n8774), .B2(n9453), .A(n7543), .ZN(n7544) );
  OAI21_X1 U9240 ( .B1(n9408), .B2(n8802), .A(n7544), .ZN(n7545) );
  AOI21_X1 U9241 ( .B1(n9561), .B2(n8804), .A(n7545), .ZN(n7546) );
  OAI21_X1 U9242 ( .B1(n7547), .B2(n8806), .A(n7546), .ZN(P1_U3236) );
  INV_X1 U9243 ( .A(n7548), .ZN(n7550) );
  AOI21_X1 U9244 ( .B1(n6764), .B2(n7938), .A(n10049), .ZN(n7549) );
  NOR3_X1 U9245 ( .A1(n7709), .A2(n7550), .A3(n7549), .ZN(n7551) );
  AOI21_X1 U9246 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(n7685), .A(n7551), .ZN(
        n7553) );
  NAND2_X1 U9247 ( .A1(n9915), .A2(n7966), .ZN(n7552) );
  OAI211_X1 U9248 ( .C1(n7723), .C2(n7554), .A(n7553), .B(n7552), .ZN(P2_U3234) );
  OR2_X1 U9249 ( .A1(n7555), .A2(n7557), .ZN(n8743) );
  INV_X1 U9250 ( .A(n8743), .ZN(n7556) );
  AOI21_X1 U9251 ( .B1(n7557), .B2(n7555), .A(n7556), .ZN(n7564) );
  INV_X1 U9252 ( .A(n7558), .ZN(n9446) );
  NOR2_X1 U9253 ( .A1(n8798), .A2(n9201), .ZN(n7561) );
  OAI22_X1 U9254 ( .A1(n8786), .A2(n9423), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7559), .ZN(n7560) );
  AOI211_X1 U9255 ( .C1(n8789), .C2(n9446), .A(n7561), .B(n7560), .ZN(n7563)
         );
  NAND2_X1 U9256 ( .A1(n9570), .A2(n8804), .ZN(n7562) );
  OAI211_X1 U9257 ( .C1(n7564), .C2(n8806), .A(n7563), .B(n7562), .ZN(P1_U3224) );
  OAI222_X1 U9258 ( .A1(n7433), .A2(n7566), .B1(n7565), .B2(P1_U3084), .C1(
        n8868), .C2(n9618), .ZN(P1_U3324) );
  INV_X1 U9259 ( .A(n8680), .ZN(n8636) );
  OAI222_X1 U9260 ( .A1(n7433), .A2(n8636), .B1(n9726), .B2(P1_U3084), .C1(
        n8681), .C2(n9618), .ZN(P1_U3325) );
  OAI222_X1 U9261 ( .A1(n5042), .A2(P2_U3152), .B1(n8635), .B2(n7567), .C1(
        n7866), .C2(n8627), .ZN(P2_U3328) );
  INV_X1 U9262 ( .A(n8297), .ZN(n8132) );
  INV_X1 U9263 ( .A(n8314), .ZN(n8181) );
  INV_X1 U9264 ( .A(n8318), .ZN(n8190) );
  INV_X1 U9265 ( .A(n7952), .ZN(n8203) );
  INV_X1 U9266 ( .A(n8240), .ZN(n7954) );
  NOR2_X1 U9267 ( .A1(n7568), .A2(n7956), .ZN(n7569) );
  OR2_X1 U9268 ( .A1(n8333), .A2(n8228), .ZN(n7811) );
  NAND2_X1 U9269 ( .A1(n8333), .A2(n8228), .ZN(n8223) );
  NAND2_X1 U9270 ( .A1(n7811), .A2(n8223), .ZN(n8236) );
  OR2_X1 U9271 ( .A1(n8329), .A2(n8240), .ZN(n7815) );
  NAND2_X1 U9272 ( .A1(n8329), .A2(n8240), .ZN(n7816) );
  NAND2_X1 U9273 ( .A1(n7815), .A2(n7816), .ZN(n8224) );
  NOR2_X1 U9274 ( .A1(n8324), .A2(n7953), .ZN(n7571) );
  INV_X1 U9275 ( .A(n8324), .ZN(n8211) );
  NAND2_X1 U9276 ( .A1(n8314), .A2(n7951), .ZN(n7830) );
  NAND2_X1 U9277 ( .A1(n7827), .A2(n7830), .ZN(n8169) );
  NAND2_X1 U9278 ( .A1(n8159), .A2(n7589), .ZN(n7573) );
  INV_X1 U9279 ( .A(n7589), .ZN(n7950) );
  NAND2_X1 U9280 ( .A1(n8302), .A2(n7628), .ZN(n7837) );
  NAND2_X1 U9281 ( .A1(n7836), .A2(n7837), .ZN(n8144) );
  INV_X1 U9282 ( .A(n8302), .ZN(n8143) );
  XNOR2_X1 U9283 ( .A(n8297), .B(n7840), .ZN(n8126) );
  NAND2_X1 U9284 ( .A1(n8294), .A2(n8094), .ZN(n7726) );
  XNOR2_X1 U9285 ( .A(n8289), .B(n7702), .ZN(n8088) );
  NAND2_X1 U9286 ( .A1(n8089), .A2(n8088), .ZN(n8087) );
  NAND2_X1 U9287 ( .A1(n8087), .A2(n7574), .ZN(n8070) );
  OR2_X1 U9288 ( .A1(n8282), .A2(n8095), .ZN(n7847) );
  NAND2_X1 U9289 ( .A1(n8282), .A2(n8095), .ZN(n7851) );
  NAND2_X1 U9290 ( .A1(n7847), .A2(n7851), .ZN(n8069) );
  INV_X1 U9291 ( .A(n8095), .ZN(n8063) );
  NAND2_X1 U9292 ( .A1(n8274), .A2(n8042), .ZN(n7852) );
  NAND2_X1 U9293 ( .A1(n8053), .A2(n8060), .ZN(n8052) );
  INV_X1 U9294 ( .A(n8274), .ZN(n7576) );
  NAND2_X1 U9295 ( .A1(n7576), .A2(n8042), .ZN(n7577) );
  NAND2_X1 U9296 ( .A1(n8052), .A2(n7577), .ZN(n8036) );
  NAND2_X1 U9297 ( .A1(n8272), .A2(n7606), .ZN(n7860) );
  NAND2_X1 U9298 ( .A1(n7854), .A2(n7860), .ZN(n8035) );
  NAND2_X1 U9299 ( .A1(n8036), .A2(n8035), .ZN(n8034) );
  NAND2_X1 U9300 ( .A1(n8049), .A2(n7606), .ZN(n7578) );
  NAND2_X1 U9301 ( .A1(n8867), .A2(n7879), .ZN(n7581) );
  NAND2_X1 U9302 ( .A1(n7579), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n7580) );
  NOR2_X1 U9303 ( .A1(n7585), .A2(n7949), .ZN(n7929) );
  NOR2_X1 U9304 ( .A1(n8265), .A2(n8041), .ZN(n7862) );
  INV_X1 U9305 ( .A(n8294), .ZN(n8122) );
  INV_X1 U9306 ( .A(n8289), .ZN(n8103) );
  AOI21_X1 U9307 ( .B1(n8265), .B2(n8043), .A(n8028), .ZN(n8266) );
  AOI22_X1 U9308 ( .A1(P2_REG2_REG_29__SCAN_IN), .A2(n8208), .B1(n7583), .B2(
        n8249), .ZN(n7584) );
  OAI21_X1 U9309 ( .B1(n7585), .B2(n10001), .A(n7584), .ZN(n7602) );
  INV_X1 U9310 ( .A(n7910), .ZN(n7805) );
  INV_X1 U9311 ( .A(n8223), .ZN(n7813) );
  NOR2_X1 U9312 ( .A1(n8224), .A2(n7813), .ZN(n7587) );
  XNOR2_X1 U9313 ( .A(n8324), .B(n8229), .ZN(n7911) );
  NAND2_X1 U9314 ( .A1(n8324), .A2(n8229), .ZN(n7826) );
  XNOR2_X1 U9315 ( .A(n8318), .B(n7952), .ZN(n8193) );
  AND2_X1 U9316 ( .A1(n8318), .A2(n8203), .ZN(n7828) );
  NOR2_X1 U9317 ( .A1(n8169), .A2(n7828), .ZN(n7588) );
  OR2_X1 U9318 ( .A1(n8307), .A2(n7589), .ZN(n7832) );
  NAND2_X1 U9319 ( .A1(n8307), .A2(n7589), .ZN(n7829) );
  NAND2_X1 U9320 ( .A1(n7832), .A2(n7829), .ZN(n8160) );
  NAND2_X1 U9321 ( .A1(n7590), .A2(n7829), .ZN(n8145) );
  AND2_X1 U9322 ( .A1(n8297), .A2(n7840), .ZN(n8108) );
  NOR2_X1 U9323 ( .A1(n8107), .A2(n8108), .ZN(n7591) );
  INV_X1 U9324 ( .A(n8088), .ZN(n8092) );
  NOR2_X1 U9325 ( .A1(n8289), .A2(n7702), .ZN(n7848) );
  INV_X1 U9326 ( .A(n8069), .ZN(n8072) );
  NAND2_X1 U9327 ( .A1(n7857), .A2(n7851), .ZN(n7592) );
  INV_X1 U9328 ( .A(n8035), .ZN(n8038) );
  XNOR2_X1 U9329 ( .A(n7931), .B(n7930), .ZN(n7600) );
  INV_X1 U9330 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n7597) );
  NAND2_X1 U9331 ( .A1(n7593), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n7596) );
  NAND2_X1 U9332 ( .A1(n7594), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n7595) );
  OAI211_X1 U9333 ( .C1(n7598), .C2(n7597), .A(n7596), .B(n7595), .ZN(n7948)
         );
  INV_X1 U9334 ( .A(n7599), .ZN(n7942) );
  AOI21_X1 U9335 ( .B1(n7942), .B2(P2_B_REG_SCAN_IN), .A(n9995), .ZN(n8024) );
  NOR2_X1 U9336 ( .A1(n8268), .A2(n8208), .ZN(n7601) );
  AOI211_X1 U9337 ( .C1(n8266), .C2(n8254), .A(n7602), .B(n7601), .ZN(n7603)
         );
  OAI21_X1 U9338 ( .B1(n8269), .B2(n8232), .A(n7603), .ZN(P2_U3267) );
  XNOR2_X1 U9339 ( .A(n7605), .B(n7604), .ZN(n7610) );
  OAI22_X1 U9340 ( .A1(n9966), .A2(n8056), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8421), .ZN(n7608) );
  OAI22_X1 U9341 ( .A1(n7606), .A2(n9954), .B1(n9959), .B2(n8095), .ZN(n7607)
         );
  AOI211_X1 U9342 ( .C1(n8274), .C2(n9957), .A(n7608), .B(n7607), .ZN(n7609)
         );
  OAI21_X1 U9343 ( .B1(n7610), .B2(n7709), .A(n7609), .ZN(P2_U3216) );
  INV_X1 U9344 ( .A(n7611), .ZN(n7659) );
  XNOR2_X1 U9345 ( .A(n7659), .B(n7658), .ZN(n7617) );
  INV_X1 U9346 ( .A(n8130), .ZN(n7613) );
  OAI22_X1 U9347 ( .A1(n9966), .A2(n7613), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7612), .ZN(n7615) );
  OAI22_X1 U9348 ( .A1(n8094), .A2(n9954), .B1(n9959), .B2(n7628), .ZN(n7614)
         );
  AOI211_X1 U9349 ( .C1(n8297), .C2(n9957), .A(n7615), .B(n7614), .ZN(n7616)
         );
  OAI21_X1 U9350 ( .B1(n7617), .B2(n7709), .A(n7616), .ZN(P2_U3218) );
  INV_X1 U9351 ( .A(n7618), .ZN(n7619) );
  AOI21_X1 U9352 ( .B1(n7621), .B2(n7620), .A(n7619), .ZN(n7625) );
  OAI22_X1 U9353 ( .A1(n7951), .A2(n9995), .B1(n8229), .B2(n8241), .ZN(n8194)
         );
  NAND2_X1 U9354 ( .A1(n9940), .A2(n8194), .ZN(n7622) );
  NAND2_X1 U9355 ( .A1(P2_U3152), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8021) );
  OAI211_X1 U9356 ( .C1(n9966), .C2(n8187), .A(n7622), .B(n8021), .ZN(n7623)
         );
  AOI21_X1 U9357 ( .B1(n8318), .B2(n9957), .A(n7623), .ZN(n7624) );
  OAI21_X1 U9358 ( .B1(n7625), .B2(n7709), .A(n7624), .ZN(P2_U3221) );
  XNOR2_X1 U9359 ( .A(n7626), .B(n7627), .ZN(n7632) );
  OAI22_X1 U9360 ( .A1(n9966), .A2(n8156), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8501), .ZN(n7630) );
  OAI22_X1 U9361 ( .A1(n7951), .A2(n9959), .B1(n9954), .B2(n7628), .ZN(n7629)
         );
  AOI211_X1 U9362 ( .C1(n8307), .C2(n9957), .A(n7630), .B(n7629), .ZN(n7631)
         );
  OAI21_X1 U9363 ( .B1(n7632), .B2(n7709), .A(n7631), .ZN(P2_U3225) );
  NAND2_X1 U9364 ( .A1(n7634), .A2(n7633), .ZN(n7636) );
  XOR2_X1 U9365 ( .A(n7636), .B(n7635), .Z(n7641) );
  OAI22_X1 U9366 ( .A1(n9966), .A2(n8099), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7637), .ZN(n7639) );
  OAI22_X1 U9367 ( .A1(n8094), .A2(n9959), .B1(n9954), .B2(n8095), .ZN(n7638)
         );
  OAI21_X1 U9368 ( .B1(n7641), .B2(n7709), .A(n7640), .ZN(P2_U3227) );
  INV_X1 U9369 ( .A(n8333), .ZN(n8252) );
  OAI21_X1 U9370 ( .B1(n7644), .B2(n7643), .A(n7642), .ZN(n7645) );
  NAND2_X1 U9371 ( .A1(n7645), .A2(n9949), .ZN(n7650) );
  INV_X1 U9372 ( .A(n7646), .ZN(n8250) );
  OAI22_X1 U9373 ( .A1(n8242), .A2(n9959), .B1(n9954), .B2(n8240), .ZN(n7647)
         );
  AOI211_X1 U9374 ( .C1(n8250), .C2(n7719), .A(n7648), .B(n7647), .ZN(n7649)
         );
  OAI211_X1 U9375 ( .C1(n8252), .C2(n7723), .A(n7650), .B(n7649), .ZN(P2_U3228) );
  XNOR2_X1 U9376 ( .A(n7652), .B(n7651), .ZN(n7656) );
  OAI22_X1 U9377 ( .A1(n9966), .A2(n8218), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8406), .ZN(n7654) );
  OAI22_X1 U9378 ( .A1(n8228), .A2(n9959), .B1(n9954), .B2(n8229), .ZN(n7653)
         );
  AOI211_X1 U9379 ( .C1(n8329), .C2(n9957), .A(n7654), .B(n7653), .ZN(n7655)
         );
  OAI21_X1 U9380 ( .B1(n7656), .B2(n7709), .A(n7655), .ZN(P2_U3230) );
  OAI21_X1 U9381 ( .B1(n7659), .B2(n7658), .A(n7657), .ZN(n7663) );
  XNOR2_X1 U9382 ( .A(n7661), .B(n7660), .ZN(n7662) );
  XNOR2_X1 U9383 ( .A(n7663), .B(n7662), .ZN(n7668) );
  OAI22_X1 U9384 ( .A1(n9966), .A2(n8118), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7664), .ZN(n7666) );
  OAI22_X1 U9385 ( .A1(n7702), .A2(n9954), .B1(n9959), .B2(n7840), .ZN(n7665)
         );
  AOI211_X1 U9386 ( .C1(n8294), .C2(n9957), .A(n7666), .B(n7665), .ZN(n7667)
         );
  OAI21_X1 U9387 ( .B1(n7668), .B2(n7709), .A(n7667), .ZN(P2_U3231) );
  XNOR2_X1 U9388 ( .A(n7669), .B(n7670), .ZN(n7675) );
  NOR2_X1 U9389 ( .A1(n9966), .A2(n8177), .ZN(n7673) );
  AOI22_X1 U9390 ( .A1(n7950), .A2(n9935), .B1(n9992), .B2(n7952), .ZN(n8173)
         );
  OAI22_X1 U9391 ( .A1(n7705), .A2(n8173), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7671), .ZN(n7672) );
  AOI211_X1 U9392 ( .C1(n8314), .C2(n9957), .A(n7673), .B(n7672), .ZN(n7674)
         );
  OAI21_X1 U9393 ( .B1(n7675), .B2(n7709), .A(n7674), .ZN(P2_U3235) );
  OAI21_X1 U9394 ( .B1(n7678), .B2(n7677), .A(n7676), .ZN(n7679) );
  NAND2_X1 U9395 ( .A1(n7679), .A2(n9949), .ZN(n7684) );
  INV_X1 U9396 ( .A(n7680), .ZN(n8141) );
  INV_X1 U9397 ( .A(n7840), .ZN(n8112) );
  AOI22_X1 U9398 ( .A1(n8112), .A2(n9935), .B1(n9992), .B2(n7950), .ZN(n8146)
         );
  OAI22_X1 U9399 ( .A1(n7705), .A2(n8146), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7681), .ZN(n7682) );
  AOI21_X1 U9400 ( .B1(n8141), .B2(n7719), .A(n7682), .ZN(n7683) );
  OAI211_X1 U9401 ( .C1(n8143), .C2(n7723), .A(n7684), .B(n7683), .ZN(P2_U3237) );
  AOI22_X1 U9402 ( .A1(n9918), .A2(n7966), .B1(n9915), .B2(n9937), .ZN(n7693)
         );
  AOI22_X1 U9403 ( .A1(n9957), .A2(n7686), .B1(P2_REG3_REG_2__SCAN_IN), .B2(
        n7685), .ZN(n7692) );
  OAI21_X1 U9404 ( .B1(n7689), .B2(n7688), .A(n7687), .ZN(n7690) );
  NAND2_X1 U9405 ( .A1(n9949), .A2(n7690), .ZN(n7691) );
  NAND3_X1 U9406 ( .A1(n7693), .A2(n7692), .A3(n7691), .ZN(P2_U3239) );
  XNOR2_X1 U9407 ( .A(n7694), .B(n7695), .ZN(n7699) );
  NAND2_X1 U9408 ( .A1(P2_U3152), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8000) );
  OAI21_X1 U9409 ( .B1(n9966), .B2(n8206), .A(n8000), .ZN(n7697) );
  OAI22_X1 U9410 ( .A1(n8240), .A2(n9959), .B1(n9954), .B2(n8203), .ZN(n7696)
         );
  AOI211_X1 U9411 ( .C1(n8324), .C2(n9957), .A(n7697), .B(n7696), .ZN(n7698)
         );
  OAI21_X1 U9412 ( .B1(n7699), .B2(n7709), .A(n7698), .ZN(P2_U3240) );
  XNOR2_X1 U9413 ( .A(n7700), .B(n7701), .ZN(n7710) );
  NOR2_X1 U9414 ( .A1(n7702), .A2(n8241), .ZN(n7703) );
  AOI21_X1 U9415 ( .B1(n4696), .B2(n9935), .A(n7703), .ZN(n8280) );
  OAI22_X1 U9416 ( .A1(n8280), .A2(n7705), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7704), .ZN(n7706) );
  AOI21_X1 U9417 ( .B1(n8079), .B2(n7719), .A(n7706), .ZN(n7708) );
  NAND2_X1 U9418 ( .A1(n8282), .A2(n9957), .ZN(n7707) );
  OAI211_X1 U9419 ( .C1(n7710), .C2(n7709), .A(n7708), .B(n7707), .ZN(P2_U3242) );
  OAI21_X1 U9420 ( .B1(n7713), .B2(n7712), .A(n7711), .ZN(n7714) );
  NAND2_X1 U9421 ( .A1(n7714), .A2(n9949), .ZN(n7722) );
  INV_X1 U9422 ( .A(n7715), .ZN(n7720) );
  OAI22_X1 U9423 ( .A1(n8228), .A2(n9954), .B1(n9959), .B2(n7716), .ZN(n7717)
         );
  AOI211_X1 U9424 ( .C1(n7720), .C2(n7719), .A(n7718), .B(n7717), .ZN(n7721)
         );
  OAI211_X1 U9425 ( .C1(n9697), .C2(n7723), .A(n7722), .B(n7721), .ZN(P2_U3243) );
  NAND2_X1 U9426 ( .A1(n7725), .A2(n7724), .ZN(n7887) );
  INV_X1 U9427 ( .A(n7726), .ZN(n7729) );
  OAI21_X1 U9428 ( .B1(n8103), .B2(n8113), .A(n7851), .ZN(n7845) );
  NOR2_X1 U9429 ( .A1(n7845), .A2(n7727), .ZN(n7728) );
  MUX2_X1 U9430 ( .A(n7729), .B(n7728), .S(n7887), .Z(n7846) );
  NAND2_X1 U9431 ( .A1(n7741), .A2(n7730), .ZN(n7732) );
  INV_X1 U9432 ( .A(n7735), .ZN(n7731) );
  MUX2_X1 U9433 ( .A(n7732), .B(n7731), .S(n7887), .Z(n7740) );
  NAND2_X1 U9434 ( .A1(n7740), .A2(n7733), .ZN(n7739) );
  NAND2_X1 U9435 ( .A1(n7735), .A2(n7734), .ZN(n7738) );
  NOR2_X1 U9436 ( .A1(n7737), .A2(n7736), .ZN(n7761) );
  AOI21_X1 U9437 ( .B1(n7739), .B2(n7738), .A(n7761), .ZN(n7745) );
  INV_X1 U9438 ( .A(n7740), .ZN(n7759) );
  NAND2_X1 U9439 ( .A1(n7741), .A2(n7762), .ZN(n7742) );
  AOI21_X1 U9440 ( .B1(n7759), .B2(n7743), .A(n7742), .ZN(n7744) );
  MUX2_X1 U9441 ( .A(n7745), .B(n7744), .S(n7887), .Z(n7767) );
  NAND2_X1 U9442 ( .A1(n7750), .A2(n7921), .ZN(n7747) );
  NAND3_X1 U9443 ( .A1(n7747), .A2(n7752), .A3(n7746), .ZN(n7748) );
  NAND3_X1 U9444 ( .A1(n7748), .A2(n7755), .A3(n7751), .ZN(n7749) );
  NAND2_X1 U9445 ( .A1(n7749), .A2(n7753), .ZN(n7758) );
  NAND2_X1 U9446 ( .A1(n7751), .A2(n7750), .ZN(n7754) );
  NAND3_X1 U9447 ( .A1(n7754), .A2(n7753), .A3(n7752), .ZN(n7756) );
  NAND2_X1 U9448 ( .A1(n7756), .A2(n7755), .ZN(n7757) );
  MUX2_X1 U9449 ( .A(n7758), .B(n7757), .S(n7890), .Z(n7760) );
  NAND3_X1 U9450 ( .A1(n7760), .A2(n7759), .A3(n7894), .ZN(n7766) );
  INV_X1 U9451 ( .A(n7761), .ZN(n7763) );
  MUX2_X1 U9452 ( .A(n7763), .B(n7762), .S(n7890), .Z(n7764) );
  NAND2_X1 U9453 ( .A1(n7764), .A2(n7901), .ZN(n7765) );
  AOI21_X1 U9454 ( .B1(n7767), .B2(n7766), .A(n7765), .ZN(n7778) );
  MUX2_X1 U9455 ( .A(n7769), .B(n7768), .S(n7890), .Z(n7770) );
  NAND2_X1 U9456 ( .A1(n7770), .A2(n9990), .ZN(n7777) );
  NAND2_X1 U9457 ( .A1(n10082), .A2(n7961), .ZN(n7771) );
  NAND2_X1 U9458 ( .A1(n7781), .A2(n7771), .ZN(n7774) );
  INV_X1 U9459 ( .A(n7772), .ZN(n7773) );
  MUX2_X1 U9460 ( .A(n7774), .B(n7773), .S(n7890), .Z(n7775) );
  NOR2_X1 U9461 ( .A1(n7775), .A2(n4620), .ZN(n7776) );
  OAI21_X1 U9462 ( .B1(n7778), .B2(n7777), .A(n7776), .ZN(n7783) );
  AND2_X1 U9463 ( .A1(n7784), .A2(n7779), .ZN(n7780) );
  MUX2_X1 U9464 ( .A(n7781), .B(n7780), .S(n7887), .Z(n7782) );
  NAND3_X1 U9465 ( .A1(n7783), .A2(n7786), .A3(n7782), .ZN(n7790) );
  AND2_X1 U9466 ( .A1(n7785), .A2(n7784), .ZN(n7788) );
  AND2_X1 U9467 ( .A1(n7793), .A2(n7786), .ZN(n7787) );
  MUX2_X1 U9468 ( .A(n7788), .B(n7787), .S(n7887), .Z(n7789) );
  NAND2_X1 U9469 ( .A1(n7790), .A2(n7789), .ZN(n7795) );
  NAND2_X1 U9470 ( .A1(n7795), .A2(n7791), .ZN(n7792) );
  NAND3_X1 U9471 ( .A1(n7795), .A2(n7794), .A3(n7793), .ZN(n7797) );
  MUX2_X1 U9472 ( .A(n7801), .B(n7800), .S(n7890), .Z(n7806) );
  NAND4_X1 U9473 ( .A1(n7803), .A2(n7908), .A3(n7887), .A4(n7802), .ZN(n7804)
         );
  NAND3_X1 U9474 ( .A1(n7806), .A2(n7805), .A3(n7804), .ZN(n7810) );
  MUX2_X1 U9475 ( .A(n7808), .B(n7807), .S(n7887), .Z(n7809) );
  INV_X1 U9476 ( .A(n7811), .ZN(n7812) );
  MUX2_X1 U9477 ( .A(n7813), .B(n7812), .S(n7890), .Z(n7814) );
  OR2_X1 U9478 ( .A1(n8324), .A2(n8229), .ZN(n7823) );
  NAND2_X1 U9479 ( .A1(n7823), .A2(n7815), .ZN(n7818) );
  INV_X1 U9480 ( .A(n7816), .ZN(n7817) );
  MUX2_X1 U9481 ( .A(n7818), .B(n7817), .S(n7890), .Z(n7819) );
  NOR2_X1 U9482 ( .A1(n8318), .A2(n8203), .ZN(n7824) );
  AOI21_X1 U9483 ( .B1(n4420), .B2(n7826), .A(n7824), .ZN(n7821) );
  NAND2_X1 U9484 ( .A1(n7830), .A2(n4519), .ZN(n7820) );
  OAI211_X1 U9485 ( .C1(n7821), .C2(n7820), .A(n7827), .B(n7832), .ZN(n7822)
         );
  NAND3_X1 U9486 ( .A1(n7822), .A2(n7837), .A3(n7829), .ZN(n7835) );
  INV_X1 U9487 ( .A(n7823), .ZN(n7825) );
  NAND3_X1 U9488 ( .A1(n7831), .A2(n7830), .A3(n7829), .ZN(n7833) );
  NAND3_X1 U9489 ( .A1(n7833), .A2(n7836), .A3(n7832), .ZN(n7834) );
  MUX2_X1 U9490 ( .A(n7835), .B(n7834), .S(n7890), .Z(n7839) );
  MUX2_X1 U9491 ( .A(n7837), .B(n7836), .S(n7887), .Z(n7838) );
  NAND2_X1 U9492 ( .A1(n8112), .A2(n7890), .ZN(n7842) );
  NAND2_X1 U9493 ( .A1(n7840), .A2(n7887), .ZN(n7841) );
  MUX2_X1 U9494 ( .A(n7842), .B(n7841), .S(n8297), .Z(n7843) );
  INV_X1 U9495 ( .A(n7847), .ZN(n7849) );
  INV_X1 U9496 ( .A(n7851), .ZN(n8059) );
  INV_X1 U9497 ( .A(n7860), .ZN(n7856) );
  INV_X1 U9498 ( .A(n7852), .ZN(n7855) );
  OAI21_X1 U9499 ( .B1(n7859), .B2(n8062), .A(n7930), .ZN(n7858) );
  OAI21_X1 U9500 ( .B1(n7862), .B2(n7887), .A(n7858), .ZN(n7865) );
  INV_X1 U9501 ( .A(n7859), .ZN(n7861) );
  OAI211_X1 U9502 ( .C1(n7890), .C2(n8272), .A(n7861), .B(n7860), .ZN(n7864)
         );
  MUX2_X1 U9503 ( .A(n7862), .B(n7929), .S(n7890), .Z(n7863) );
  AOI21_X1 U9504 ( .B1(n7865), .B2(n7864), .A(n7863), .ZN(n7885) );
  NOR2_X1 U9505 ( .A1(n5091), .A2(n7866), .ZN(n7867) );
  NAND2_X1 U9506 ( .A1(n8264), .A2(n7948), .ZN(n7935) );
  INV_X1 U9507 ( .A(n8264), .ZN(n8030) );
  INV_X1 U9508 ( .A(n7948), .ZN(n7868) );
  NAND2_X1 U9509 ( .A1(n8030), .A2(n7868), .ZN(n7883) );
  NAND2_X1 U9510 ( .A1(n7935), .A2(n7883), .ZN(n7884) );
  INV_X1 U9511 ( .A(n7869), .ZN(n7870) );
  NAND2_X1 U9512 ( .A1(n7870), .A2(SI_30_), .ZN(n7874) );
  MUX2_X1 U9513 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n4478), .Z(n7876) );
  XNOR2_X1 U9514 ( .A(n7876), .B(SI_31_), .ZN(n7877) );
  NAND2_X1 U9515 ( .A1(n9623), .A2(n7879), .ZN(n7881) );
  OR2_X1 U9516 ( .A1(n5091), .A2(n6451), .ZN(n7880) );
  INV_X1 U9517 ( .A(n8025), .ZN(n7882) );
  OR2_X1 U9518 ( .A1(n8257), .A2(n7882), .ZN(n7891) );
  NAND2_X1 U9519 ( .A1(n7891), .A2(n7883), .ZN(n7934) );
  INV_X1 U9520 ( .A(n7934), .ZN(n7917) );
  INV_X1 U9521 ( .A(n8257), .ZN(n7886) );
  NOR2_X1 U9522 ( .A1(n7886), .A2(n8025), .ZN(n7937) );
  INV_X1 U9523 ( .A(n7937), .ZN(n7888) );
  NAND2_X1 U9524 ( .A1(n7888), .A2(n7935), .ZN(n7893) );
  AOI22_X1 U9525 ( .A1(n7889), .A2(n7888), .B1(n7893), .B2(n7887), .ZN(n7928)
         );
  INV_X1 U9526 ( .A(n7924), .ZN(n7892) );
  NOR2_X1 U9527 ( .A1(n7891), .A2(n7890), .ZN(n7927) );
  NOR3_X1 U9528 ( .A1(n7928), .A2(n7892), .A3(n7927), .ZN(n7922) );
  INV_X1 U9529 ( .A(n7893), .ZN(n7918) );
  INV_X1 U9530 ( .A(n8169), .ZN(n8172) );
  NAND4_X1 U9531 ( .A1(n7896), .A2(n7895), .A3(n7894), .A4(n7923), .ZN(n7898)
         );
  NOR4_X1 U9532 ( .A1(n7898), .A2(n7897), .A3(n10014), .A4(n10051), .ZN(n7902)
         );
  NAND4_X1 U9533 ( .A1(n7902), .A2(n7901), .A3(n7900), .A4(n7899), .ZN(n7904)
         );
  NOR4_X1 U9534 ( .A1(n7904), .A2(n7094), .A3(n4395), .A4(n7903), .ZN(n7905)
         );
  NAND4_X1 U9535 ( .A1(n7908), .A2(n7907), .A3(n7906), .A4(n7905), .ZN(n7909)
         );
  NOR4_X1 U9536 ( .A1(n8224), .A2(n8236), .A3(n7910), .A4(n7909), .ZN(n7912)
         );
  INV_X1 U9537 ( .A(n7911), .ZN(n8200) );
  NAND4_X1 U9538 ( .A1(n8172), .A2(n7912), .A3(n8193), .A4(n8200), .ZN(n7913)
         );
  NOR4_X1 U9539 ( .A1(n8107), .A2(n8144), .A3(n8160), .A4(n7913), .ZN(n7914)
         );
  NAND4_X1 U9540 ( .A1(n8072), .A2(n7914), .A3(n4928), .A4(n8092), .ZN(n7915)
         );
  NOR3_X1 U9541 ( .A1(n8035), .A2(n8060), .A3(n7915), .ZN(n7916) );
  NAND4_X1 U9542 ( .A1(n7918), .A2(n7930), .A3(n7917), .A4(n7916), .ZN(n7919)
         );
  XNOR2_X1 U9543 ( .A(n7919), .B(n8020), .ZN(n7920) );
  AOI21_X1 U9544 ( .B1(n7925), .B2(n7924), .A(n7923), .ZN(n7926) );
  OAI21_X1 U9545 ( .B1(n7928), .B2(n7927), .A(n7926), .ZN(n7940) );
  INV_X1 U9546 ( .A(n7933), .ZN(n7936) );
  NAND4_X1 U9547 ( .A1(n7943), .A2(n7942), .A3(n7941), .A4(n9992), .ZN(n7944)
         );
  OAI211_X1 U9548 ( .C1(n5048), .C2(n7946), .A(n7944), .B(P2_B_REG_SCAN_IN), 
        .ZN(n7945) );
  OAI21_X1 U9549 ( .B1(n7947), .B2(n7946), .A(n7945), .ZN(P2_U3244) );
  MUX2_X1 U9550 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n7948), .S(P2_U3966), .Z(
        P2_U3582) );
  MUX2_X1 U9551 ( .A(n7949), .B(P2_DATAO_REG_29__SCAN_IN), .S(n7967), .Z(
        P2_U3581) );
  MUX2_X1 U9552 ( .A(n8062), .B(P2_DATAO_REG_28__SCAN_IN), .S(n7967), .Z(
        P2_U3580) );
  MUX2_X1 U9553 ( .A(n4696), .B(P2_DATAO_REG_27__SCAN_IN), .S(n7967), .Z(
        P2_U3579) );
  MUX2_X1 U9554 ( .A(n8063), .B(P2_DATAO_REG_26__SCAN_IN), .S(n7967), .Z(
        P2_U3578) );
  MUX2_X1 U9555 ( .A(n8113), .B(P2_DATAO_REG_25__SCAN_IN), .S(n7967), .Z(
        P2_U3577) );
  MUX2_X1 U9556 ( .A(n8134), .B(P2_DATAO_REG_24__SCAN_IN), .S(n7967), .Z(
        P2_U3576) );
  MUX2_X1 U9557 ( .A(n8112), .B(P2_DATAO_REG_23__SCAN_IN), .S(n7967), .Z(
        P2_U3575) );
  MUX2_X1 U9558 ( .A(n8163), .B(P2_DATAO_REG_22__SCAN_IN), .S(n7967), .Z(
        P2_U3574) );
  MUX2_X1 U9559 ( .A(n7950), .B(P2_DATAO_REG_21__SCAN_IN), .S(n7967), .Z(
        P2_U3573) );
  INV_X1 U9560 ( .A(n7951), .ZN(n8162) );
  MUX2_X1 U9561 ( .A(n8162), .B(P2_DATAO_REG_20__SCAN_IN), .S(n7967), .Z(
        P2_U3572) );
  MUX2_X1 U9562 ( .A(n7952), .B(P2_DATAO_REG_19__SCAN_IN), .S(n7967), .Z(
        P2_U3571) );
  MUX2_X1 U9563 ( .A(n7953), .B(P2_DATAO_REG_18__SCAN_IN), .S(n7967), .Z(
        P2_U3570) );
  MUX2_X1 U9564 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n7954), .S(P2_U3966), .Z(
        P2_U3569) );
  MUX2_X1 U9565 ( .A(n7955), .B(P2_DATAO_REG_16__SCAN_IN), .S(n7967), .Z(
        P2_U3568) );
  MUX2_X1 U9566 ( .A(n7956), .B(P2_DATAO_REG_15__SCAN_IN), .S(n7967), .Z(
        P2_U3567) );
  MUX2_X1 U9567 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n7957), .S(P2_U3966), .Z(
        P2_U3566) );
  MUX2_X1 U9568 ( .A(n7958), .B(P2_DATAO_REG_13__SCAN_IN), .S(n7967), .Z(
        P2_U3565) );
  MUX2_X1 U9569 ( .A(n7959), .B(P2_DATAO_REG_12__SCAN_IN), .S(n7967), .Z(
        P2_U3564) );
  MUX2_X1 U9570 ( .A(n9914), .B(P2_DATAO_REG_11__SCAN_IN), .S(n7963), .Z(
        P2_U3563) );
  MUX2_X1 U9571 ( .A(n7960), .B(P2_DATAO_REG_10__SCAN_IN), .S(n7963), .Z(
        P2_U3562) );
  MUX2_X1 U9572 ( .A(n9917), .B(P2_DATAO_REG_9__SCAN_IN), .S(n7963), .Z(
        P2_U3561) );
  MUX2_X1 U9573 ( .A(n7961), .B(P2_DATAO_REG_8__SCAN_IN), .S(n7963), .Z(
        P2_U3560) );
  MUX2_X1 U9574 ( .A(n9993), .B(P2_DATAO_REG_7__SCAN_IN), .S(n7963), .Z(
        P2_U3559) );
  MUX2_X1 U9575 ( .A(n7962), .B(P2_DATAO_REG_6__SCAN_IN), .S(n7963), .Z(
        P2_U3558) );
  MUX2_X1 U9576 ( .A(n9936), .B(P2_DATAO_REG_5__SCAN_IN), .S(n7963), .Z(
        P2_U3557) );
  MUX2_X1 U9577 ( .A(n7964), .B(P2_DATAO_REG_4__SCAN_IN), .S(n7963), .Z(
        P2_U3556) );
  MUX2_X1 U9578 ( .A(n9937), .B(P2_DATAO_REG_3__SCAN_IN), .S(n7967), .Z(
        P2_U3555) );
  MUX2_X1 U9579 ( .A(n7965), .B(P2_DATAO_REG_2__SCAN_IN), .S(n7967), .Z(
        P2_U3554) );
  MUX2_X1 U9580 ( .A(n7966), .B(P2_DATAO_REG_1__SCAN_IN), .S(n7967), .Z(
        P2_U3553) );
  MUX2_X1 U9581 ( .A(n6764), .B(P2_DATAO_REG_0__SCAN_IN), .S(n7967), .Z(
        P2_U3552) );
  NAND2_X1 U9582 ( .A1(n9659), .A2(n7968), .ZN(n7979) );
  OAI211_X1 U9583 ( .C1(n7971), .C2(n7970), .A(n9968), .B(n7969), .ZN(n7978)
         );
  NOR2_X1 U9584 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8562), .ZN(n7972) );
  AOI21_X1 U9585 ( .B1(n9969), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n7972), .ZN(
        n7977) );
  OAI211_X1 U9586 ( .C1(n7975), .C2(n7974), .A(n9967), .B(n7973), .ZN(n7976)
         );
  NAND4_X1 U9587 ( .A1(n7979), .A2(n7978), .A3(n7977), .A4(n7976), .ZN(
        P2_U3255) );
  NAND2_X1 U9588 ( .A1(n7981), .A2(n7980), .ZN(n7983) );
  MUX2_X1 U9589 ( .A(P2_REG2_REG_17__SCAN_IN), .B(n8219), .S(n7996), .Z(n7982)
         );
  NAND2_X1 U9590 ( .A1(n7982), .A2(n7983), .ZN(n7992) );
  OAI211_X1 U9591 ( .C1(n7983), .C2(n7982), .A(n9968), .B(n7992), .ZN(n7991)
         );
  NOR2_X1 U9592 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8406), .ZN(n7989) );
  XNOR2_X1 U9593 ( .A(n7996), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n7986) );
  AOI211_X1 U9594 ( .C1(n7987), .C2(n7986), .A(n7995), .B(n9972), .ZN(n7988)
         );
  AOI211_X1 U9595 ( .C1(P2_ADDR_REG_17__SCAN_IN), .C2(n9969), .A(n7989), .B(
        n7988), .ZN(n7990) );
  OAI211_X1 U9596 ( .C1(n9971), .C2(n7993), .A(n7991), .B(n7990), .ZN(P2_U3262) );
  OAI21_X1 U9597 ( .B1(n7993), .B2(n8219), .A(n7992), .ZN(n8012) );
  XNOR2_X1 U9598 ( .A(n8012), .B(n8011), .ZN(n8010) );
  XOR2_X1 U9599 ( .A(P2_REG2_REG_18__SCAN_IN), .B(n8010), .Z(n8005) );
  INV_X1 U9600 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n8002) );
  XNOR2_X1 U9601 ( .A(n8011), .B(n7994), .ZN(n7998) );
  OAI21_X1 U9602 ( .B1(n7998), .B2(n7997), .A(n8007), .ZN(n7999) );
  NAND2_X1 U9603 ( .A1(n9967), .A2(n7999), .ZN(n8001) );
  OAI211_X1 U9604 ( .C1(n8022), .C2(n8002), .A(n8001), .B(n8000), .ZN(n8003)
         );
  AOI21_X1 U9605 ( .B1(n8011), .B2(n9659), .A(n8003), .ZN(n8004) );
  OAI21_X1 U9606 ( .B1(n8005), .B2(n9970), .A(n8004), .ZN(P2_U3263) );
  OR2_X1 U9607 ( .A1(n8011), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8006) );
  NAND2_X1 U9608 ( .A1(n8007), .A2(n8006), .ZN(n8008) );
  XNOR2_X1 U9609 ( .A(n8008), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8017) );
  OR2_X1 U9610 ( .A1(n8010), .A2(n8009), .ZN(n8014) );
  NAND2_X1 U9611 ( .A1(n8012), .A2(n8011), .ZN(n8013) );
  NAND2_X1 U9612 ( .A1(n8014), .A2(n8013), .ZN(n8015) );
  XNOR2_X1 U9613 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n8015), .ZN(n8019) );
  NAND2_X1 U9614 ( .A1(n8019), .A2(n9968), .ZN(n8016) );
  INV_X1 U9615 ( .A(n8017), .ZN(n8018) );
  NOR2_X1 U9616 ( .A1(n10035), .A2(n8023), .ZN(n8026) );
  NAND2_X1 U9617 ( .A1(n8025), .A2(n8024), .ZN(n8262) );
  NOR2_X1 U9618 ( .A1(n8208), .A2(n8262), .ZN(n8031) );
  AOI211_X1 U9619 ( .C1(n8257), .C2(n8071), .A(n8026), .B(n8031), .ZN(n8027)
         );
  OAI21_X1 U9620 ( .B1(n8259), .B2(n9986), .A(n8027), .ZN(P2_U3265) );
  INV_X1 U9621 ( .A(n8028), .ZN(n8029) );
  NAND2_X1 U9622 ( .A1(n8030), .A2(n8029), .ZN(n8261) );
  NAND3_X1 U9623 ( .A1(n8261), .A2(n8254), .A3(n8260), .ZN(n8033) );
  AOI21_X1 U9624 ( .B1(n8208), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8031), .ZN(
        n8032) );
  OAI211_X1 U9625 ( .C1(n8264), .C2(n10001), .A(n8033), .B(n8032), .ZN(
        P2_U3266) );
  OAI21_X1 U9626 ( .B1(n8036), .B2(n8035), .A(n8034), .ZN(n8037) );
  INV_X1 U9627 ( .A(n8037), .ZN(n8273) );
  XNOR2_X1 U9628 ( .A(n8039), .B(n8038), .ZN(n8040) );
  INV_X1 U9629 ( .A(n8055), .ZN(n8045) );
  INV_X1 U9630 ( .A(n8043), .ZN(n8044) );
  AOI211_X1 U9631 ( .C1(n8272), .C2(n8045), .A(n10102), .B(n8044), .ZN(n8271)
         );
  NAND2_X1 U9632 ( .A1(n8271), .A2(n8222), .ZN(n8048) );
  AOI22_X1 U9633 ( .A1(n8046), .A2(n8249), .B1(n8208), .B2(
        P2_REG2_REG_28__SCAN_IN), .ZN(n8047) );
  OAI211_X1 U9634 ( .C1(n8049), .C2(n10001), .A(n8048), .B(n8047), .ZN(n8050)
         );
  AOI21_X1 U9635 ( .B1(n8270), .B2(n10035), .A(n8050), .ZN(n8051) );
  OAI21_X1 U9636 ( .B1(n8273), .B2(n8232), .A(n8051), .ZN(P2_U3268) );
  OAI21_X1 U9637 ( .B1(n8053), .B2(n8060), .A(n8052), .ZN(n8054) );
  INV_X1 U9638 ( .A(n8054), .ZN(n8278) );
  AOI21_X1 U9639 ( .B1(n8274), .B2(n8077), .A(n8055), .ZN(n8275) );
  INV_X1 U9640 ( .A(n8056), .ZN(n8057) );
  AOI22_X1 U9641 ( .A1(n8208), .A2(P2_REG2_REG_27__SCAN_IN), .B1(n8057), .B2(
        n8249), .ZN(n8058) );
  OAI21_X1 U9642 ( .B1(n7576), .B2(n10001), .A(n8058), .ZN(n8066) );
  NOR2_X1 U9643 ( .A1(n8075), .A2(n8059), .ZN(n8061) );
  XNOR2_X1 U9644 ( .A(n8061), .B(n8060), .ZN(n8064) );
  NOR2_X1 U9645 ( .A1(n8277), .A2(n8208), .ZN(n8065) );
  AOI211_X1 U9646 ( .C1(n8275), .C2(n8254), .A(n8066), .B(n8065), .ZN(n8067)
         );
  OAI21_X1 U9647 ( .B1(n8278), .B2(n8232), .A(n8067), .ZN(P2_U3269) );
  OAI21_X1 U9648 ( .B1(n8070), .B2(n8069), .A(n8068), .ZN(n8279) );
  INV_X1 U9649 ( .A(n8279), .ZN(n8086) );
  AOI22_X1 U9650 ( .A1(n8282), .A2(n8071), .B1(n8208), .B2(
        P2_REG2_REG_26__SCAN_IN), .ZN(n8085) );
  NOR2_X1 U9651 ( .A1(n8073), .A2(n8072), .ZN(n8074) );
  NAND2_X1 U9652 ( .A1(n8076), .A2(n10012), .ZN(n8284) );
  INV_X1 U9653 ( .A(n8284), .ZN(n8083) );
  AOI21_X1 U9654 ( .B1(n8096), .B2(n8282), .A(n10102), .ZN(n8078) );
  NAND2_X1 U9655 ( .A1(n8078), .A2(n8077), .ZN(n8283) );
  NAND2_X1 U9656 ( .A1(n8079), .A2(n8249), .ZN(n8080) );
  OAI211_X1 U9657 ( .C1(n8283), .C2(n8081), .A(n8280), .B(n8080), .ZN(n8082)
         );
  OAI21_X1 U9658 ( .B1(n8083), .B2(n8082), .A(n10035), .ZN(n8084) );
  OAI211_X1 U9659 ( .C1(n8086), .C2(n8232), .A(n8085), .B(n8084), .ZN(P2_U3270) );
  OAI21_X1 U9660 ( .B1(n8089), .B2(n8088), .A(n8087), .ZN(n8090) );
  INV_X1 U9661 ( .A(n8090), .ZN(n8291) );
  XNOR2_X1 U9662 ( .A(n8092), .B(n8091), .ZN(n8093) );
  OAI222_X1 U9663 ( .A1(n9995), .A2(n8095), .B1(n8241), .B2(n8094), .C1(n8093), 
        .C2(n8226), .ZN(n8287) );
  INV_X1 U9664 ( .A(n8116), .ZN(n8098) );
  INV_X1 U9665 ( .A(n8096), .ZN(n8097) );
  AOI211_X1 U9666 ( .C1(n8289), .C2(n8098), .A(n10102), .B(n8097), .ZN(n8288)
         );
  NAND2_X1 U9667 ( .A1(n8288), .A2(n8222), .ZN(n8102) );
  INV_X1 U9668 ( .A(n8099), .ZN(n8100) );
  AOI22_X1 U9669 ( .A1(n8208), .A2(P2_REG2_REG_25__SCAN_IN), .B1(n8100), .B2(
        n8249), .ZN(n8101) );
  OAI211_X1 U9670 ( .C1(n8103), .C2(n10001), .A(n8102), .B(n8101), .ZN(n8104)
         );
  AOI21_X1 U9671 ( .B1(n8287), .B2(n10035), .A(n8104), .ZN(n8105) );
  OAI21_X1 U9672 ( .B1(n8291), .B2(n8232), .A(n8105), .ZN(P2_U3271) );
  XNOR2_X1 U9673 ( .A(n8106), .B(n8107), .ZN(n8296) );
  INV_X1 U9674 ( .A(n8133), .ZN(n8109) );
  OAI21_X1 U9675 ( .B1(n8109), .B2(n8108), .A(n8107), .ZN(n8111) );
  NAND3_X1 U9676 ( .A1(n8111), .A2(n10012), .A3(n8110), .ZN(n8115) );
  AOI22_X1 U9677 ( .A1(n8113), .A2(n9935), .B1(n9992), .B2(n8112), .ZN(n8114)
         );
  NAND2_X1 U9678 ( .A1(n8115), .A2(n8114), .ZN(n8292) );
  INV_X1 U9679 ( .A(n8128), .ZN(n8117) );
  AOI211_X1 U9680 ( .C1(n8294), .C2(n8117), .A(n10102), .B(n8116), .ZN(n8293)
         );
  NAND2_X1 U9681 ( .A1(n8293), .A2(n8222), .ZN(n8121) );
  INV_X1 U9682 ( .A(n8118), .ZN(n8119) );
  AOI22_X1 U9683 ( .A1(n8208), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n8119), .B2(
        n8249), .ZN(n8120) );
  OAI211_X1 U9684 ( .C1(n8122), .C2(n10001), .A(n8121), .B(n8120), .ZN(n8123)
         );
  AOI21_X1 U9685 ( .B1(n8292), .B2(n10035), .A(n8123), .ZN(n8124) );
  OAI21_X1 U9686 ( .B1(n8296), .B2(n8232), .A(n8124), .ZN(P2_U3272) );
  OAI21_X1 U9687 ( .B1(n8127), .B2(n8126), .A(n8125), .ZN(n8301) );
  INV_X1 U9688 ( .A(n8140), .ZN(n8129) );
  AOI21_X1 U9689 ( .B1(n8297), .B2(n8129), .A(n8128), .ZN(n8298) );
  AOI22_X1 U9690 ( .A1(n8208), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n8130), .B2(
        n8249), .ZN(n8131) );
  OAI21_X1 U9691 ( .B1(n8132), .B2(n10001), .A(n8131), .ZN(n8137) );
  OAI21_X1 U9692 ( .B1(n4417), .B2(n4928), .A(n8133), .ZN(n8135) );
  AOI222_X1 U9693 ( .A1(n10012), .A2(n8135), .B1(n8163), .B2(n9992), .C1(n8134), .C2(n9935), .ZN(n8300) );
  NOR2_X1 U9694 ( .A1(n8300), .A2(n8208), .ZN(n8136) );
  AOI211_X1 U9695 ( .C1(n8298), .C2(n8254), .A(n8137), .B(n8136), .ZN(n8138)
         );
  OAI21_X1 U9696 ( .B1(n8301), .B2(n8232), .A(n8138), .ZN(P2_U3273) );
  XOR2_X1 U9697 ( .A(n8139), .B(n8144), .Z(n8306) );
  AOI21_X1 U9698 ( .B1(n8302), .B2(n8154), .A(n8140), .ZN(n8303) );
  AOI22_X1 U9699 ( .A1(n8208), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8141), .B2(
        n8249), .ZN(n8142) );
  OAI21_X1 U9700 ( .B1(n8143), .B2(n10001), .A(n8142), .ZN(n8151) );
  AOI21_X1 U9701 ( .B1(n8145), .B2(n8144), .A(n8226), .ZN(n8149) );
  INV_X1 U9702 ( .A(n8146), .ZN(n8147) );
  AOI21_X1 U9703 ( .B1(n8149), .B2(n8148), .A(n8147), .ZN(n8305) );
  NOR2_X1 U9704 ( .A1(n8305), .A2(n8208), .ZN(n8150) );
  AOI211_X1 U9705 ( .C1(n8303), .C2(n8254), .A(n8151), .B(n8150), .ZN(n8152)
         );
  OAI21_X1 U9706 ( .B1(n8306), .B2(n8232), .A(n8152), .ZN(P2_U3274) );
  XNOR2_X1 U9707 ( .A(n4476), .B(n8160), .ZN(n8311) );
  INV_X1 U9708 ( .A(n8154), .ZN(n8155) );
  AOI21_X1 U9709 ( .B1(n8307), .B2(n8176), .A(n8155), .ZN(n8308) );
  INV_X1 U9710 ( .A(n8156), .ZN(n8157) );
  AOI22_X1 U9711 ( .A1(n8208), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8157), .B2(
        n8249), .ZN(n8158) );
  OAI21_X1 U9712 ( .B1(n8159), .B2(n10001), .A(n8158), .ZN(n8166) );
  XNOR2_X1 U9713 ( .A(n8161), .B(n8160), .ZN(n8164) );
  AOI222_X1 U9714 ( .A1(n10012), .A2(n8164), .B1(n8163), .B2(n9935), .C1(n8162), .C2(n9992), .ZN(n8310) );
  NOR2_X1 U9715 ( .A1(n8310), .A2(n8208), .ZN(n8165) );
  AOI211_X1 U9716 ( .C1(n8308), .C2(n8254), .A(n8166), .B(n8165), .ZN(n8167)
         );
  OAI21_X1 U9717 ( .B1(n8311), .B2(n8232), .A(n8167), .ZN(P2_U3275) );
  OAI21_X1 U9718 ( .B1(n8170), .B2(n8169), .A(n8168), .ZN(n8316) );
  NAND2_X1 U9719 ( .A1(n8171), .A2(n10012), .ZN(n8175) );
  AOI21_X1 U9720 ( .B1(n8191), .B2(n4519), .A(n8172), .ZN(n8174) );
  OAI21_X1 U9721 ( .B1(n8175), .B2(n8174), .A(n8173), .ZN(n8312) );
  AOI211_X1 U9722 ( .C1(n8314), .C2(n8185), .A(n10102), .B(n4545), .ZN(n8313)
         );
  NAND2_X1 U9723 ( .A1(n8313), .A2(n8222), .ZN(n8180) );
  INV_X1 U9724 ( .A(n8177), .ZN(n8178) );
  AOI22_X1 U9725 ( .A1(n8208), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8178), .B2(
        n8249), .ZN(n8179) );
  OAI211_X1 U9726 ( .C1(n8181), .C2(n10001), .A(n8180), .B(n8179), .ZN(n8182)
         );
  AOI21_X1 U9727 ( .B1(n8312), .B2(n10035), .A(n8182), .ZN(n8183) );
  OAI21_X1 U9728 ( .B1(n8316), .B2(n8232), .A(n8183), .ZN(P2_U3276) );
  XOR2_X1 U9729 ( .A(n8184), .B(n8193), .Z(n8321) );
  INV_X1 U9730 ( .A(n8204), .ZN(n8186) );
  AOI211_X1 U9731 ( .C1(n8318), .C2(n8186), .A(n10102), .B(n4546), .ZN(n8317)
         );
  INV_X1 U9732 ( .A(n8187), .ZN(n8188) );
  AOI22_X1 U9733 ( .A1(n8208), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n8188), .B2(
        n8249), .ZN(n8189) );
  OAI21_X1 U9734 ( .B1(n8190), .B2(n10001), .A(n8189), .ZN(n8197) );
  OAI21_X1 U9735 ( .B1(n8193), .B2(n8192), .A(n8191), .ZN(n8195) );
  AOI21_X1 U9736 ( .B1(n8195), .B2(n10012), .A(n8194), .ZN(n8320) );
  NOR2_X1 U9737 ( .A1(n8320), .A2(n8208), .ZN(n8196) );
  AOI211_X1 U9738 ( .C1(n8317), .C2(n8222), .A(n8197), .B(n8196), .ZN(n8198)
         );
  OAI21_X1 U9739 ( .B1(n8321), .B2(n8232), .A(n8198), .ZN(P2_U3277) );
  XNOR2_X1 U9740 ( .A(n8199), .B(n8200), .ZN(n8326) );
  XNOR2_X1 U9741 ( .A(n8201), .B(n8200), .ZN(n8202) );
  OAI222_X1 U9742 ( .A1(n9995), .A2(n8203), .B1(n8241), .B2(n8240), .C1(n8202), 
        .C2(n8226), .ZN(n8322) );
  INV_X1 U9743 ( .A(n8217), .ZN(n8205) );
  AOI211_X1 U9744 ( .C1(n8324), .C2(n8205), .A(n10102), .B(n8204), .ZN(n8323)
         );
  NAND2_X1 U9745 ( .A1(n8323), .A2(n8222), .ZN(n8210) );
  INV_X1 U9746 ( .A(n8206), .ZN(n8207) );
  AOI22_X1 U9747 ( .A1(n8208), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8207), .B2(
        n8249), .ZN(n8209) );
  OAI211_X1 U9748 ( .C1(n8211), .C2(n10001), .A(n8210), .B(n8209), .ZN(n8212)
         );
  AOI21_X1 U9749 ( .B1(n8322), .B2(n10035), .A(n8212), .ZN(n8213) );
  OAI21_X1 U9750 ( .B1(n8326), .B2(n8232), .A(n8213), .ZN(P2_U3278) );
  OAI21_X1 U9751 ( .B1(n8215), .B2(n8224), .A(n8214), .ZN(n8216) );
  INV_X1 U9752 ( .A(n8216), .ZN(n8332) );
  AOI211_X1 U9753 ( .C1(n8329), .C2(n8248), .A(n10102), .B(n8217), .ZN(n8328)
         );
  NOR2_X1 U9754 ( .A1(n4944), .A2(n10001), .ZN(n8221) );
  OAI22_X1 U9755 ( .A1(n10035), .A2(n8219), .B1(n8218), .B2(n10028), .ZN(n8220) );
  AOI211_X1 U9756 ( .C1(n8328), .C2(n8222), .A(n8221), .B(n8220), .ZN(n8231)
         );
  NAND2_X1 U9757 ( .A1(n8239), .A2(n8223), .ZN(n8225) );
  XNOR2_X1 U9758 ( .A(n8225), .B(n8224), .ZN(n8227) );
  OAI222_X1 U9759 ( .A1(n9995), .A2(n8229), .B1(n8241), .B2(n8228), .C1(n8227), 
        .C2(n8226), .ZN(n8327) );
  NAND2_X1 U9760 ( .A1(n8327), .A2(n10035), .ZN(n8230) );
  OAI211_X1 U9761 ( .C1(n8332), .C2(n8232), .A(n8231), .B(n8230), .ZN(P2_U3279) );
  NOR2_X1 U9762 ( .A1(n8233), .A2(n8236), .ZN(n8234) );
  NAND2_X1 U9763 ( .A1(n8237), .A2(n8236), .ZN(n8238) );
  NAND2_X1 U9764 ( .A1(n8239), .A2(n8238), .ZN(n8244) );
  OAI22_X1 U9765 ( .A1(n8242), .A2(n8241), .B1(n8240), .B2(n9995), .ZN(n8243)
         );
  AOI21_X1 U9766 ( .B1(n8244), .B2(n10012), .A(n8243), .ZN(n8245) );
  OAI21_X1 U9767 ( .B1(n8336), .B2(n9989), .A(n8245), .ZN(n8338) );
  NAND2_X1 U9768 ( .A1(n8338), .A2(n10035), .ZN(n8256) );
  NAND2_X1 U9769 ( .A1(n8246), .A2(n8333), .ZN(n8247) );
  AND2_X1 U9770 ( .A1(n8248), .A2(n8247), .ZN(n8334) );
  AOI22_X1 U9771 ( .A1(n8208), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n8250), .B2(
        n8249), .ZN(n8251) );
  OAI21_X1 U9772 ( .B1(n8252), .B2(n10001), .A(n8251), .ZN(n8253) );
  AOI21_X1 U9773 ( .B1(n8334), .B2(n8254), .A(n8253), .ZN(n8255) );
  OAI211_X1 U9774 ( .C1(n8336), .C2(n9987), .A(n8256), .B(n8255), .ZN(P2_U3280) );
  NAND2_X1 U9775 ( .A1(n8257), .A2(n10024), .ZN(n8258) );
  OAI211_X1 U9776 ( .C1(n8259), .C2(n10102), .A(n8258), .B(n8262), .ZN(n8339)
         );
  MUX2_X1 U9777 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n8339), .S(n10124), .Z(
        P2_U3551) );
  NAND3_X1 U9778 ( .A1(n8261), .A2(n10022), .A3(n8260), .ZN(n8263) );
  OAI211_X1 U9779 ( .C1(n8264), .C2(n10110), .A(n8263), .B(n8262), .ZN(n8610)
         );
  MUX2_X1 U9780 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n8610), .S(n10124), .Z(
        P2_U3550) );
  AOI22_X1 U9781 ( .A1(n8266), .A2(n10022), .B1(n10024), .B2(n8265), .ZN(n8267) );
  OAI211_X1 U9782 ( .C1(n8269), .C2(n8331), .A(n8268), .B(n8267), .ZN(n8611)
         );
  MUX2_X1 U9783 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n8611), .S(n10124), .Z(
        P2_U3549) );
  MUX2_X1 U9784 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n8612), .S(n10124), .Z(
        P2_U3548) );
  AOI22_X1 U9785 ( .A1(n8275), .A2(n10022), .B1(n10024), .B2(n8274), .ZN(n8276) );
  OAI211_X1 U9786 ( .C1(n8278), .C2(n8331), .A(n8277), .B(n8276), .ZN(n8613)
         );
  MUX2_X1 U9787 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n8613), .S(n10124), .Z(
        P2_U3547) );
  NAND2_X1 U9788 ( .A1(n8279), .A2(n10114), .ZN(n8286) );
  INV_X1 U9789 ( .A(n8280), .ZN(n8281) );
  AOI21_X1 U9790 ( .B1(n8282), .B2(n10024), .A(n8281), .ZN(n8285) );
  NAND4_X1 U9791 ( .A1(n8286), .A2(n8285), .A3(n8284), .A4(n8283), .ZN(n8614)
         );
  MUX2_X1 U9792 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n8614), .S(n10124), .Z(
        P2_U3546) );
  AOI211_X1 U9793 ( .C1(n10024), .C2(n8289), .A(n8288), .B(n8287), .ZN(n8290)
         );
  OAI21_X1 U9794 ( .B1(n8291), .B2(n8331), .A(n8290), .ZN(n8615) );
  MUX2_X1 U9795 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n8615), .S(n10124), .Z(
        P2_U3545) );
  AOI211_X1 U9796 ( .C1(n10024), .C2(n8294), .A(n8293), .B(n8292), .ZN(n8295)
         );
  OAI21_X1 U9797 ( .B1(n8296), .B2(n8331), .A(n8295), .ZN(n8616) );
  MUX2_X1 U9798 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8616), .S(n10124), .Z(
        P2_U3544) );
  AOI22_X1 U9799 ( .A1(n8298), .A2(n10022), .B1(n10024), .B2(n8297), .ZN(n8299) );
  OAI211_X1 U9800 ( .C1(n8301), .C2(n8331), .A(n8300), .B(n8299), .ZN(n8617)
         );
  MUX2_X1 U9801 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n8617), .S(n10124), .Z(
        P2_U3543) );
  AOI22_X1 U9802 ( .A1(n8303), .A2(n10022), .B1(n10024), .B2(n8302), .ZN(n8304) );
  OAI211_X1 U9803 ( .C1(n8306), .C2(n8331), .A(n8305), .B(n8304), .ZN(n8618)
         );
  MUX2_X1 U9804 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n8618), .S(n10124), .Z(
        P2_U3542) );
  AOI22_X1 U9805 ( .A1(n8308), .A2(n10022), .B1(n10024), .B2(n8307), .ZN(n8309) );
  OAI211_X1 U9806 ( .C1(n8311), .C2(n8331), .A(n8310), .B(n8309), .ZN(n8619)
         );
  MUX2_X1 U9807 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n8619), .S(n10124), .Z(
        P2_U3541) );
  AOI211_X1 U9808 ( .C1(n10024), .C2(n8314), .A(n8313), .B(n8312), .ZN(n8315)
         );
  OAI21_X1 U9809 ( .B1(n8316), .B2(n8331), .A(n8315), .ZN(n8620) );
  MUX2_X1 U9810 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n8620), .S(n10124), .Z(
        P2_U3540) );
  AOI21_X1 U9811 ( .B1(n10024), .B2(n8318), .A(n8317), .ZN(n8319) );
  OAI211_X1 U9812 ( .C1(n8321), .C2(n8331), .A(n8320), .B(n8319), .ZN(n8621)
         );
  MUX2_X1 U9813 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8621), .S(n10124), .Z(
        P2_U3539) );
  AOI211_X1 U9814 ( .C1(n10024), .C2(n8324), .A(n8323), .B(n8322), .ZN(n8325)
         );
  OAI21_X1 U9815 ( .B1(n8326), .B2(n8331), .A(n8325), .ZN(n8622) );
  MUX2_X1 U9816 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n8622), .S(n10124), .Z(
        P2_U3538) );
  AOI211_X1 U9817 ( .C1(n10024), .C2(n8329), .A(n8328), .B(n8327), .ZN(n8330)
         );
  OAI21_X1 U9818 ( .B1(n8332), .B2(n8331), .A(n8330), .ZN(n8623) );
  MUX2_X1 U9819 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n8623), .S(n10124), .Z(
        P2_U3537) );
  AOI22_X1 U9820 ( .A1(n8334), .A2(n10022), .B1(n10024), .B2(n8333), .ZN(n8335) );
  OAI21_X1 U9821 ( .B1(n8336), .B2(n10080), .A(n8335), .ZN(n8337) );
  OR2_X1 U9822 ( .A1(n8338), .A2(n8337), .ZN(n8624) );
  MUX2_X1 U9823 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n8624), .S(n10124), .Z(
        P2_U3536) );
  MUX2_X1 U9824 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n8339), .S(n10117), .Z(n8609) );
  NAND4_X1 U9825 ( .A1(P1_D_REG_24__SCAN_IN), .A2(P2_REG3_REG_0__SCAN_IN), 
        .A3(n8398), .A4(n8394), .ZN(n8347) );
  NAND4_X1 U9826 ( .A1(P1_REG1_REG_11__SCAN_IN), .A2(P2_REG1_REG_22__SCAN_IN), 
        .A3(n8501), .A4(n6356), .ZN(n8346) );
  NOR4_X1 U9827 ( .A1(SI_18_), .A2(P1_DATAO_REG_16__SCAN_IN), .A3(n8587), .A4(
        n8556), .ZN(n8344) );
  NOR4_X1 U9828 ( .A1(SI_22_), .A2(SI_20_), .A3(n8578), .A4(n8340), .ZN(n8343)
         );
  NOR4_X1 U9829 ( .A1(P2_IR_REG_28__SCAN_IN), .A2(P2_DATAO_REG_1__SCAN_IN), 
        .A3(P2_REG1_REG_31__SCAN_IN), .A4(n8590), .ZN(n8342) );
  NOR4_X1 U9830 ( .A1(P2_DATAO_REG_6__SCAN_IN), .A2(P2_DATAO_REG_10__SCAN_IN), 
        .A3(n8552), .A4(n8436), .ZN(n8341) );
  NAND4_X1 U9831 ( .A1(n8344), .A2(n8343), .A3(n8342), .A4(n8341), .ZN(n8345)
         );
  NOR3_X1 U9832 ( .A1(n8347), .A2(n8346), .A3(n8345), .ZN(n8390) );
  NOR4_X1 U9833 ( .A1(P1_IR_REG_30__SCAN_IN), .A2(P2_REG1_REG_15__SCAN_IN), 
        .A3(n8426), .A4(n8468), .ZN(n8348) );
  AND3_X1 U9834 ( .A1(P1_D_REG_19__SCAN_IN), .A2(P1_REG3_REG_5__SCAN_IN), .A3(
        n8348), .ZN(n8379) );
  AND4_X1 U9835 ( .A1(n8350), .A2(n4997), .A3(n8349), .A4(
        P1_REG0_REG_26__SCAN_IN), .ZN(n8359) );
  AND4_X1 U9836 ( .A1(n8409), .A2(n8351), .A3(P1_IR_REG_2__SCAN_IN), .A4(
        P2_DATAO_REG_27__SCAN_IN), .ZN(n8358) );
  INV_X1 U9837 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n8563) );
  NAND4_X1 U9838 ( .A1(P1_REG0_REG_21__SCAN_IN), .A2(P2_REG2_REG_17__SCAN_IN), 
        .A3(n8563), .A4(n6370), .ZN(n8353) );
  NAND4_X1 U9839 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(P2_REG1_REG_7__SCAN_IN), 
        .A3(P2_REG1_REG_6__SCAN_IN), .A4(n8516), .ZN(n8352) );
  NOR2_X1 U9840 ( .A1(n8353), .A2(n8352), .ZN(n8354) );
  INV_X1 U9841 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n8493) );
  AND4_X1 U9842 ( .A1(n8354), .A2(n5275), .A3(P2_IR_REG_4__SCAN_IN), .A4(
        P2_IR_REG_16__SCAN_IN), .ZN(n8355) );
  AND4_X1 U9843 ( .A1(n4712), .A2(P1_IR_REG_3__SCAN_IN), .A3(
        P1_IR_REG_4__SCAN_IN), .A4(n8355), .ZN(n8357) );
  NOR2_X1 U9844 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(P2_ADDR_REG_12__SCAN_IN), 
        .ZN(n8356) );
  NAND4_X1 U9845 ( .A1(n8359), .A2(n8358), .A3(n8357), .A4(n8356), .ZN(n8361)
         );
  INV_X1 U9846 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n9687) );
  NAND4_X1 U9847 ( .A1(P1_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_3__SCAN_IN), 
        .A3(P1_ADDR_REG_18__SCAN_IN), .A4(n9687), .ZN(n8360) );
  NOR2_X1 U9848 ( .A1(n8361), .A2(n8360), .ZN(n8373) );
  NAND2_X1 U9849 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n9673) );
  NAND4_X1 U9850 ( .A1(n8362), .A2(n9682), .A3(P2_REG3_REG_19__SCAN_IN), .A4(
        P2_REG1_REG_4__SCAN_IN), .ZN(n8365) );
  NAND4_X1 U9851 ( .A1(n8363), .A2(n8421), .A3(P2_IR_REG_19__SCAN_IN), .A4(
        P2_IR_REG_31__SCAN_IN), .ZN(n8364) );
  NOR3_X1 U9852 ( .A1(n9673), .A2(n8365), .A3(n8364), .ZN(n8372) );
  NAND4_X1 U9853 ( .A1(P1_REG1_REG_21__SCAN_IN), .A2(P1_REG2_REG_19__SCAN_IN), 
        .A3(n5990), .A4(n8576), .ZN(n8367) );
  INV_X1 U9854 ( .A(P1_WR_REG_SCAN_IN), .ZN(n8447) );
  NAND4_X1 U9855 ( .A1(P1_REG1_REG_7__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), 
        .A3(P2_REG2_REG_6__SCAN_IN), .A4(n8447), .ZN(n8366) );
  NOR2_X1 U9856 ( .A1(n8367), .A2(n8366), .ZN(n8371) );
  NAND4_X1 U9857 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_REG0_REG_24__SCAN_IN), 
        .A3(n5913), .A4(n8579), .ZN(n8369) );
  INV_X1 U9858 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10116) );
  NAND4_X1 U9859 ( .A1(P1_REG1_REG_16__SCAN_IN), .A2(P1_REG0_REG_19__SCAN_IN), 
        .A3(n8490), .A4(n10116), .ZN(n8368) );
  NOR2_X1 U9860 ( .A1(n8369), .A2(n8368), .ZN(n8370) );
  AND4_X1 U9861 ( .A1(n8373), .A2(n8372), .A3(n8371), .A4(n8370), .ZN(n8378)
         );
  NAND4_X1 U9862 ( .A1(P1_REG0_REG_28__SCAN_IN), .A2(P1_REG2_REG_11__SCAN_IN), 
        .A3(P1_REG2_REG_29__SCAN_IN), .A4(P2_REG2_REG_11__SCAN_IN), .ZN(n8374)
         );
  NOR3_X1 U9863 ( .A1(P1_REG3_REG_28__SCAN_IN), .A2(P2_REG1_REG_2__SCAN_IN), 
        .A3(n8374), .ZN(n8377) );
  NOR4_X1 U9864 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), 
        .A3(P2_STATE_REG_SCAN_IN), .A4(P2_D_REG_0__SCAN_IN), .ZN(n8375) );
  AND3_X1 U9865 ( .A1(SI_25_), .A2(n8375), .A3(n8411), .ZN(n8376) );
  NAND4_X1 U9866 ( .A1(n8379), .A2(n8378), .A3(n8377), .A4(n8376), .ZN(n8388)
         );
  NOR4_X1 U9867 ( .A1(P1_REG2_REG_24__SCAN_IN), .A2(P2_REG3_REG_17__SCAN_IN), 
        .A3(P2_REG3_REG_9__SCAN_IN), .A4(P2_REG1_REG_24__SCAN_IN), .ZN(n8386)
         );
  NOR4_X1 U9868 ( .A1(P1_REG2_REG_27__SCAN_IN), .A2(P2_REG3_REG_10__SCAN_IN), 
        .A3(P2_REG2_REG_29__SCAN_IN), .A4(n5848), .ZN(n8385) );
  INV_X1 U9869 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9879) );
  NAND4_X1 U9870 ( .A1(P2_REG2_REG_12__SCAN_IN), .A2(P2_REG1_REG_1__SCAN_IN), 
        .A3(n9136), .A4(n9879), .ZN(n8383) );
  NAND4_X1 U9871 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_REG3_REG_8__SCAN_IN), 
        .A3(P2_REG3_REG_8__SCAN_IN), .A4(P2_REG2_REG_13__SCAN_IN), .ZN(n8382)
         );
  NAND4_X1 U9872 ( .A1(P1_REG2_REG_20__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), 
        .A3(P2_REG3_REG_11__SCAN_IN), .A4(n8508), .ZN(n8381) );
  NAND4_X1 U9873 ( .A1(P1_REG1_REG_6__SCAN_IN), .A2(P2_REG0_REG_3__SCAN_IN), 
        .A3(n8506), .A4(n5793), .ZN(n8380) );
  NOR4_X1 U9874 ( .A1(n8383), .A2(n8382), .A3(n8381), .A4(n8380), .ZN(n8384)
         );
  NAND3_X1 U9875 ( .A1(n8386), .A2(n8385), .A3(n8384), .ZN(n8387) );
  NOR2_X1 U9876 ( .A1(n8388), .A2(n8387), .ZN(n8389) );
  NAND4_X1 U9877 ( .A1(n8392), .A2(n8391), .A3(n8390), .A4(n8389), .ZN(n8607)
         );
  AOI22_X1 U9878 ( .A1(n8394), .A2(keyinput101), .B1(keyinput3), .B2(P2_U3152), 
        .ZN(n8393) );
  OAI221_X1 U9879 ( .B1(n8394), .B2(keyinput101), .C1(P2_U3152), .C2(keyinput3), .A(n8393), .ZN(n8404) );
  INV_X1 U9880 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n9832) );
  AOI22_X1 U9881 ( .A1(n9832), .A2(keyinput98), .B1(keyinput113), .B2(n5049), 
        .ZN(n8395) );
  OAI221_X1 U9882 ( .B1(n9832), .B2(keyinput98), .C1(n5049), .C2(keyinput113), 
        .A(n8395), .ZN(n8403) );
  INV_X1 U9883 ( .A(SI_18_), .ZN(n8397) );
  AOI22_X1 U9884 ( .A1(n8398), .A2(keyinput119), .B1(n8397), .B2(keyinput0), 
        .ZN(n8396) );
  OAI221_X1 U9885 ( .B1(n8398), .B2(keyinput119), .C1(n8397), .C2(keyinput0), 
        .A(n8396), .ZN(n8402) );
  INV_X1 U9886 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n8400) );
  AOI22_X1 U9887 ( .A1(n8400), .A2(keyinput91), .B1(n6067), .B2(keyinput29), 
        .ZN(n8399) );
  OAI221_X1 U9888 ( .B1(n8400), .B2(keyinput91), .C1(n6067), .C2(keyinput29), 
        .A(n8399), .ZN(n8401) );
  NOR4_X1 U9889 ( .A1(n8404), .A2(n8403), .A3(n8402), .A4(n8401), .ZN(n8419)
         );
  AOI22_X1 U9890 ( .A1(n8407), .A2(keyinput83), .B1(n8406), .B2(keyinput7), 
        .ZN(n8405) );
  OAI221_X1 U9891 ( .B1(n8407), .B2(keyinput83), .C1(n8406), .C2(keyinput7), 
        .A(n8405), .ZN(n8417) );
  AOI22_X1 U9892 ( .A1(n9682), .A2(keyinput28), .B1(n8409), .B2(keyinput110), 
        .ZN(n8408) );
  OAI221_X1 U9893 ( .B1(n9682), .B2(keyinput28), .C1(n8409), .C2(keyinput110), 
        .A(n8408), .ZN(n8416) );
  AOI22_X1 U9894 ( .A1(n8412), .A2(keyinput64), .B1(n8411), .B2(keyinput13), 
        .ZN(n8410) );
  OAI221_X1 U9895 ( .B1(n8412), .B2(keyinput64), .C1(n8411), .C2(keyinput13), 
        .A(n8410), .ZN(n8415) );
  INV_X1 U9896 ( .A(P2_D_REG_19__SCAN_IN), .ZN(n10039) );
  AOI22_X1 U9897 ( .A1(n7424), .A2(keyinput81), .B1(n10039), .B2(keyinput80), 
        .ZN(n8413) );
  OAI221_X1 U9898 ( .B1(n7424), .B2(keyinput81), .C1(n10039), .C2(keyinput80), 
        .A(n8413), .ZN(n8414) );
  NOR4_X1 U9899 ( .A1(n8417), .A2(n8416), .A3(n8415), .A4(n8414), .ZN(n8418)
         );
  NAND2_X1 U9900 ( .A1(n8419), .A2(n8418), .ZN(n8605) );
  AOI22_X1 U9901 ( .A1(n5871), .A2(keyinput122), .B1(keyinput33), .B2(n8421), 
        .ZN(n8420) );
  OAI221_X1 U9902 ( .B1(n5871), .B2(keyinput122), .C1(n8421), .C2(keyinput33), 
        .A(n8420), .ZN(n8430) );
  AOI22_X1 U9903 ( .A1(n8423), .A2(keyinput105), .B1(n4712), .B2(keyinput46), 
        .ZN(n8422) );
  OAI221_X1 U9904 ( .B1(n8423), .B2(keyinput105), .C1(n4712), .C2(keyinput46), 
        .A(n8422), .ZN(n8429) );
  INV_X1 U9905 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n9833) );
  AOI22_X1 U9906 ( .A1(n9833), .A2(keyinput77), .B1(keyinput96), .B2(n5384), 
        .ZN(n8424) );
  OAI221_X1 U9907 ( .B1(n9833), .B2(keyinput77), .C1(n5384), .C2(keyinput96), 
        .A(n8424), .ZN(n8428) );
  AOI22_X1 U9908 ( .A1(n8426), .A2(keyinput120), .B1(keyinput94), .B2(n5911), 
        .ZN(n8425) );
  OAI221_X1 U9909 ( .B1(n8426), .B2(keyinput120), .C1(n5911), .C2(keyinput94), 
        .A(n8425), .ZN(n8427) );
  NOR4_X1 U9910 ( .A1(n8430), .A2(n8429), .A3(n8428), .A4(n8427), .ZN(n8549)
         );
  INV_X1 U9911 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n10041) );
  AOI22_X1 U9912 ( .A1(n10041), .A2(keyinput104), .B1(keyinput106), .B2(n6465), 
        .ZN(n8431) );
  OAI221_X1 U9913 ( .B1(n10041), .B2(keyinput104), .C1(n6465), .C2(keyinput106), .A(n8431), .ZN(n8434) );
  AOI22_X1 U9914 ( .A1(n10043), .A2(keyinput54), .B1(keyinput16), .B2(n7216), 
        .ZN(n8432) );
  OAI221_X1 U9915 ( .B1(n10043), .B2(keyinput54), .C1(n7216), .C2(keyinput16), 
        .A(n8432), .ZN(n8433) );
  NOR2_X1 U9916 ( .A1(n8434), .A2(n8433), .ZN(n8453) );
  AOI22_X1 U9917 ( .A1(n8436), .A2(keyinput17), .B1(keyinput44), .B2(n9136), 
        .ZN(n8435) );
  OAI221_X1 U9918 ( .B1(n8436), .B2(keyinput17), .C1(n9136), .C2(keyinput44), 
        .A(n8435), .ZN(n8440) );
  AOI22_X1 U9919 ( .A1(n8438), .A2(keyinput18), .B1(keyinput11), .B2(n6468), 
        .ZN(n8437) );
  OAI221_X1 U9920 ( .B1(n8438), .B2(keyinput18), .C1(n6468), .C2(keyinput11), 
        .A(n8437), .ZN(n8439) );
  NOR2_X1 U9921 ( .A1(n8440), .A2(n8439), .ZN(n8452) );
  AOI22_X1 U9922 ( .A1(n4966), .A2(keyinput20), .B1(keyinput66), .B2(n7365), 
        .ZN(n8441) );
  OAI221_X1 U9923 ( .B1(n4966), .B2(keyinput20), .C1(n7365), .C2(keyinput66), 
        .A(n8441), .ZN(n8444) );
  INV_X1 U9924 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n9642) );
  AOI22_X1 U9925 ( .A1(n6356), .A2(keyinput8), .B1(keyinput109), .B2(n9642), 
        .ZN(n8442) );
  OAI221_X1 U9926 ( .B1(n6356), .B2(keyinput8), .C1(n9642), .C2(keyinput109), 
        .A(n8442), .ZN(n8443) );
  NOR2_X1 U9927 ( .A1(n8444), .A2(n8443), .ZN(n8451) );
  AOI22_X1 U9928 ( .A1(n5793), .A2(keyinput79), .B1(keyinput121), .B2(n5083), 
        .ZN(n8445) );
  OAI221_X1 U9929 ( .B1(n5793), .B2(keyinput79), .C1(n5083), .C2(keyinput121), 
        .A(n8445), .ZN(n8449) );
  AOI22_X1 U9930 ( .A1(n6486), .A2(keyinput73), .B1(keyinput68), .B2(n8447), 
        .ZN(n8446) );
  OAI221_X1 U9931 ( .B1(n6486), .B2(keyinput73), .C1(n8447), .C2(keyinput68), 
        .A(n8446), .ZN(n8448) );
  NOR2_X1 U9932 ( .A1(n8449), .A2(n8448), .ZN(n8450) );
  NAND4_X1 U9933 ( .A1(n8453), .A2(n8452), .A3(n8451), .A4(n8450), .ZN(n8484)
         );
  INV_X1 U9934 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10177) );
  AOI22_X1 U9935 ( .A1(n10177), .A2(keyinput6), .B1(n7307), .B2(keyinput74), 
        .ZN(n8454) );
  OAI221_X1 U9936 ( .B1(n10177), .B2(keyinput6), .C1(n7307), .C2(keyinput74), 
        .A(n8454), .ZN(n8462) );
  AOI22_X1 U9937 ( .A1(n8457), .A2(keyinput116), .B1(n8456), .B2(keyinput1), 
        .ZN(n8455) );
  OAI221_X1 U9938 ( .B1(n8457), .B2(keyinput116), .C1(n8456), .C2(keyinput1), 
        .A(n8455), .ZN(n8461) );
  XNOR2_X1 U9939 ( .A(keyinput36), .B(P1_REG0_REG_7__SCAN_IN), .ZN(n8459) );
  XNOR2_X1 U9940 ( .A(keyinput27), .B(P2_REG1_REG_8__SCAN_IN), .ZN(n8458) );
  NAND2_X1 U9941 ( .A1(n8459), .A2(n8458), .ZN(n8460) );
  NOR3_X1 U9942 ( .A1(n8462), .A2(n8461), .A3(n8460), .ZN(n8482) );
  INV_X1 U9943 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n10038) );
  INV_X1 U9944 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n9836) );
  AOI22_X1 U9945 ( .A1(n10038), .A2(keyinput84), .B1(n9836), .B2(keyinput87), 
        .ZN(n8463) );
  OAI221_X1 U9946 ( .B1(n10038), .B2(keyinput84), .C1(n9836), .C2(keyinput87), 
        .A(n8463), .ZN(n8466) );
  AOI22_X1 U9947 ( .A1(n10171), .A2(keyinput30), .B1(n5764), .B2(keyinput89), 
        .ZN(n8464) );
  OAI221_X1 U9948 ( .B1(n10171), .B2(keyinput30), .C1(n5764), .C2(keyinput89), 
        .A(n8464), .ZN(n8465) );
  NOR2_X1 U9949 ( .A1(n8466), .A2(n8465), .ZN(n8481) );
  INV_X1 U9950 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n9617) );
  AOI22_X1 U9951 ( .A1(n8468), .A2(keyinput126), .B1(n9617), .B2(keyinput103), 
        .ZN(n8467) );
  OAI221_X1 U9952 ( .B1(n8468), .B2(keyinput126), .C1(n9617), .C2(keyinput103), 
        .A(n8467), .ZN(n8471) );
  INV_X1 U9953 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n9830) );
  AOI22_X1 U9954 ( .A1(n5275), .A2(keyinput21), .B1(n9830), .B2(keyinput49), 
        .ZN(n8469) );
  OAI221_X1 U9955 ( .B1(n5275), .B2(keyinput21), .C1(n9830), .C2(keyinput49), 
        .A(n8469), .ZN(n8470) );
  NOR2_X1 U9956 ( .A1(n8471), .A2(n8470), .ZN(n8480) );
  INV_X1 U9957 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n8473) );
  AOI22_X1 U9958 ( .A1(n8474), .A2(keyinput117), .B1(keyinput67), .B2(n8473), 
        .ZN(n8472) );
  OAI221_X1 U9959 ( .B1(n8474), .B2(keyinput117), .C1(n8473), .C2(keyinput67), 
        .A(n8472), .ZN(n8478) );
  INV_X1 U9960 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n9834) );
  AOI22_X1 U9961 ( .A1(n8476), .A2(keyinput107), .B1(n9834), .B2(keyinput58), 
        .ZN(n8475) );
  OAI221_X1 U9962 ( .B1(n8476), .B2(keyinput107), .C1(n9834), .C2(keyinput58), 
        .A(n8475), .ZN(n8477) );
  NOR2_X1 U9963 ( .A1(n8478), .A2(n8477), .ZN(n8479) );
  NAND4_X1 U9964 ( .A1(n8482), .A2(n8481), .A3(n8480), .A4(n8479), .ZN(n8483)
         );
  NOR2_X1 U9965 ( .A1(n8484), .A2(n8483), .ZN(n8548) );
  AOI22_X1 U9966 ( .A1(n6466), .A2(keyinput69), .B1(n6324), .B2(keyinput72), 
        .ZN(n8485) );
  OAI221_X1 U9967 ( .B1(n6466), .B2(keyinput69), .C1(n6324), .C2(keyinput72), 
        .A(n8485), .ZN(n8497) );
  AOI22_X1 U9968 ( .A1(n10116), .A2(keyinput37), .B1(n8487), .B2(keyinput90), 
        .ZN(n8486) );
  OAI221_X1 U9969 ( .B1(n10116), .B2(keyinput37), .C1(n8487), .C2(keyinput90), 
        .A(n8486), .ZN(n8496) );
  AOI22_X1 U9970 ( .A1(n8490), .A2(keyinput65), .B1(n8489), .B2(keyinput124), 
        .ZN(n8488) );
  OAI221_X1 U9971 ( .B1(n8490), .B2(keyinput65), .C1(n8489), .C2(keyinput124), 
        .A(n8488), .ZN(n8495) );
  AOI22_X1 U9972 ( .A1(n8493), .A2(keyinput92), .B1(n8492), .B2(keyinput48), 
        .ZN(n8491) );
  OAI221_X1 U9973 ( .B1(n8493), .B2(keyinput92), .C1(n8492), .C2(keyinput48), 
        .A(n8491), .ZN(n8494) );
  NOR4_X1 U9974 ( .A1(n8497), .A2(n8496), .A3(n8495), .A4(n8494), .ZN(n8547)
         );
  AOI22_X1 U9975 ( .A1(n9687), .A2(keyinput43), .B1(n8499), .B2(keyinput39), 
        .ZN(n8498) );
  OAI221_X1 U9976 ( .B1(n9687), .B2(keyinput43), .C1(n8499), .C2(keyinput39), 
        .A(n8498), .ZN(n8504) );
  AOI22_X1 U9977 ( .A1(n5988), .A2(keyinput50), .B1(keyinput9), .B2(n8501), 
        .ZN(n8500) );
  OAI221_X1 U9978 ( .B1(n5988), .B2(keyinput50), .C1(n8501), .C2(keyinput9), 
        .A(n8500), .ZN(n8503) );
  INV_X1 U9979 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n9835) );
  XNOR2_X1 U9980 ( .A(n9835), .B(keyinput42), .ZN(n8502) );
  NOR3_X1 U9981 ( .A1(n8504), .A2(n8503), .A3(n8502), .ZN(n8545) );
  AOI22_X1 U9982 ( .A1(n8506), .A2(keyinput86), .B1(keyinput15), .B2(n5890), 
        .ZN(n8505) );
  OAI221_X1 U9983 ( .B1(n8506), .B2(keyinput86), .C1(n5890), .C2(keyinput15), 
        .A(n8505), .ZN(n8514) );
  AOI22_X1 U9984 ( .A1(n9376), .A2(keyinput35), .B1(keyinput63), .B2(n8508), 
        .ZN(n8507) );
  OAI221_X1 U9985 ( .B1(n9376), .B2(keyinput35), .C1(n8508), .C2(keyinput63), 
        .A(n8507), .ZN(n8513) );
  INV_X1 U9986 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n8510) );
  AOI22_X1 U9987 ( .A1(n8511), .A2(keyinput45), .B1(keyinput75), .B2(n8510), 
        .ZN(n8509) );
  OAI221_X1 U9988 ( .B1(n8511), .B2(keyinput45), .C1(n8510), .C2(keyinput75), 
        .A(n8509), .ZN(n8512) );
  NOR3_X1 U9989 ( .A1(n8514), .A2(n8513), .A3(n8512), .ZN(n8544) );
  AOI22_X1 U9990 ( .A1(n8516), .A2(keyinput111), .B1(keyinput118), .B2(n6470), 
        .ZN(n8515) );
  OAI221_X1 U9991 ( .B1(n8516), .B2(keyinput111), .C1(n6470), .C2(keyinput118), 
        .A(n8515), .ZN(n8519) );
  INV_X1 U9992 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n8517) );
  XNOR2_X1 U9993 ( .A(n8517), .B(keyinput22), .ZN(n8518) );
  NOR2_X1 U9994 ( .A1(n8519), .A2(n8518), .ZN(n8543) );
  XNOR2_X1 U9995 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(keyinput25), .ZN(n8523) );
  XNOR2_X1 U9996 ( .A(P2_IR_REG_8__SCAN_IN), .B(keyinput56), .ZN(n8522) );
  XNOR2_X1 U9997 ( .A(P2_IR_REG_15__SCAN_IN), .B(keyinput88), .ZN(n8521) );
  XNOR2_X1 U9998 ( .A(P2_REG1_REG_22__SCAN_IN), .B(keyinput112), .ZN(n8520) );
  NAND4_X1 U9999 ( .A1(n8523), .A2(n8522), .A3(n8521), .A4(n8520), .ZN(n8529)
         );
  XNOR2_X1 U10000 ( .A(P1_REG2_REG_2__SCAN_IN), .B(keyinput102), .ZN(n8527) );
  XNOR2_X1 U10001 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput47), .ZN(n8526) );
  XNOR2_X1 U10002 ( .A(P2_IR_REG_28__SCAN_IN), .B(keyinput52), .ZN(n8525) );
  XNOR2_X1 U10003 ( .A(P2_IR_REG_19__SCAN_IN), .B(keyinput108), .ZN(n8524) );
  NAND4_X1 U10004 ( .A1(n8527), .A2(n8526), .A3(n8525), .A4(n8524), .ZN(n8528)
         );
  NOR2_X1 U10005 ( .A1(n8529), .A2(n8528), .ZN(n8541) );
  XNOR2_X1 U10006 ( .A(P1_IR_REG_8__SCAN_IN), .B(keyinput71), .ZN(n8533) );
  XNOR2_X1 U10007 ( .A(P2_IR_REG_31__SCAN_IN), .B(keyinput59), .ZN(n8532) );
  XNOR2_X1 U10008 ( .A(P2_REG3_REG_8__SCAN_IN), .B(keyinput34), .ZN(n8531) );
  XNOR2_X1 U10009 ( .A(P2_IR_REG_3__SCAN_IN), .B(keyinput62), .ZN(n8530) );
  NAND4_X1 U10010 ( .A1(n8533), .A2(n8532), .A3(n8531), .A4(n8530), .ZN(n8539)
         );
  XNOR2_X1 U10011 ( .A(P1_IR_REG_26__SCAN_IN), .B(keyinput51), .ZN(n8537) );
  XNOR2_X1 U10012 ( .A(P1_IR_REG_12__SCAN_IN), .B(keyinput53), .ZN(n8536) );
  XNOR2_X1 U10013 ( .A(P2_IR_REG_20__SCAN_IN), .B(keyinput70), .ZN(n8535) );
  XNOR2_X1 U10014 ( .A(keyinput40), .B(P2_REG3_REG_11__SCAN_IN), .ZN(n8534) );
  NAND4_X1 U10015 ( .A1(n8537), .A2(n8536), .A3(n8535), .A4(n8534), .ZN(n8538)
         );
  NOR2_X1 U10016 ( .A1(n8539), .A2(n8538), .ZN(n8540) );
  AND2_X1 U10017 ( .A1(n8541), .A2(n8540), .ZN(n8542) );
  AND4_X1 U10018 ( .A1(n8545), .A2(n8544), .A3(n8543), .A4(n8542), .ZN(n8546)
         );
  NAND4_X1 U10019 ( .A1(n8549), .A2(n8548), .A3(n8547), .A4(n8546), .ZN(n8604)
         );
  INV_X1 U10020 ( .A(P1_D_REG_25__SCAN_IN), .ZN(n9831) );
  AOI22_X1 U10021 ( .A1(n9831), .A2(keyinput93), .B1(keyinput57), .B2(n8219), 
        .ZN(n8550) );
  OAI221_X1 U10022 ( .B1(n9831), .B2(keyinput93), .C1(n8219), .C2(keyinput57), 
        .A(n8550), .ZN(n8560) );
  AOI22_X1 U10023 ( .A1(n6370), .A2(keyinput41), .B1(n8552), .B2(keyinput95), 
        .ZN(n8551) );
  OAI221_X1 U10024 ( .B1(n6370), .B2(keyinput41), .C1(n8552), .C2(keyinput95), 
        .A(n8551), .ZN(n8559) );
  INV_X1 U10025 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n10040) );
  AOI22_X1 U10026 ( .A1(n8554), .A2(keyinput115), .B1(keyinput55), .B2(n10040), 
        .ZN(n8553) );
  OAI221_X1 U10027 ( .B1(n8554), .B2(keyinput115), .C1(n10040), .C2(keyinput55), .A(n8553), .ZN(n8558) );
  AOI22_X1 U10028 ( .A1(n4551), .A2(keyinput97), .B1(n8556), .B2(keyinput10), 
        .ZN(n8555) );
  OAI221_X1 U10029 ( .B1(n4551), .B2(keyinput97), .C1(n8556), .C2(keyinput10), 
        .A(n8555), .ZN(n8557) );
  NOR4_X1 U10030 ( .A1(n8560), .A2(n8559), .A3(n8558), .A4(n8557), .ZN(n8602)
         );
  AOI22_X1 U10031 ( .A1(n8563), .A2(keyinput85), .B1(keyinput61), .B2(n8562), 
        .ZN(n8561) );
  OAI221_X1 U10032 ( .B1(n8563), .B2(keyinput85), .C1(n8562), .C2(keyinput61), 
        .A(n8561), .ZN(n8572) );
  AOI22_X1 U10033 ( .A1(n5848), .A2(keyinput32), .B1(n6274), .B2(keyinput19), 
        .ZN(n8564) );
  OAI221_X1 U10034 ( .B1(n5848), .B2(keyinput32), .C1(n6274), .C2(keyinput19), 
        .A(n8564), .ZN(n8571) );
  AOI22_X1 U10035 ( .A1(n8566), .A2(keyinput60), .B1(n4912), .B2(keyinput24), 
        .ZN(n8565) );
  OAI221_X1 U10036 ( .B1(n8566), .B2(keyinput60), .C1(n4912), .C2(keyinput24), 
        .A(n8565), .ZN(n8570) );
  INV_X1 U10037 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n9808) );
  AOI22_X1 U10038 ( .A1(n9808), .A2(keyinput26), .B1(n8568), .B2(keyinput100), 
        .ZN(n8567) );
  OAI221_X1 U10039 ( .B1(n9808), .B2(keyinput26), .C1(n8568), .C2(keyinput100), 
        .A(n8567), .ZN(n8569) );
  NOR4_X1 U10040 ( .A1(n8572), .A2(n8571), .A3(n8570), .A4(n8569), .ZN(n8601)
         );
  AOI22_X1 U10041 ( .A1(n8574), .A2(keyinput78), .B1(keyinput4), .B2(n6143), 
        .ZN(n8573) );
  OAI221_X1 U10042 ( .B1(n8574), .B2(keyinput78), .C1(n6143), .C2(keyinput4), 
        .A(n8573), .ZN(n8585) );
  AOI22_X1 U10043 ( .A1(n8576), .A2(keyinput5), .B1(n5990), .B2(keyinput31), 
        .ZN(n8575) );
  OAI221_X1 U10044 ( .B1(n8576), .B2(keyinput5), .C1(n5990), .C2(keyinput31), 
        .A(n8575), .ZN(n8584) );
  AOI22_X1 U10045 ( .A1(n8579), .A2(keyinput125), .B1(n8578), .B2(keyinput38), 
        .ZN(n8577) );
  OAI221_X1 U10046 ( .B1(n8579), .B2(keyinput125), .C1(n8578), .C2(keyinput38), 
        .A(n8577), .ZN(n8583) );
  AOI22_X1 U10047 ( .A1(n5913), .A2(keyinput114), .B1(keyinput23), .B2(n8581), 
        .ZN(n8580) );
  OAI221_X1 U10048 ( .B1(n5913), .B2(keyinput114), .C1(n8581), .C2(keyinput23), 
        .A(n8580), .ZN(n8582) );
  NOR4_X1 U10049 ( .A1(n8585), .A2(n8584), .A3(n8583), .A4(n8582), .ZN(n8600)
         );
  AOI22_X1 U10050 ( .A1(n8588), .A2(keyinput2), .B1(n8587), .B2(keyinput123), 
        .ZN(n8586) );
  OAI221_X1 U10051 ( .B1(n8588), .B2(keyinput2), .C1(n8587), .C2(keyinput123), 
        .A(n8586), .ZN(n8598) );
  AOI22_X1 U10052 ( .A1(n8590), .A2(keyinput14), .B1(keyinput127), .B2(n6506), 
        .ZN(n8589) );
  OAI221_X1 U10053 ( .B1(n8590), .B2(keyinput14), .C1(n6506), .C2(keyinput127), 
        .A(n8589), .ZN(n8597) );
  AOI22_X1 U10054 ( .A1(n8592), .A2(keyinput12), .B1(n5738), .B2(keyinput82), 
        .ZN(n8591) );
  OAI221_X1 U10055 ( .B1(n8592), .B2(keyinput12), .C1(n5738), .C2(keyinput82), 
        .A(n8591), .ZN(n8596) );
  AOI22_X1 U10056 ( .A1(n8594), .A2(keyinput99), .B1(keyinput76), .B2(n8681), 
        .ZN(n8593) );
  OAI221_X1 U10057 ( .B1(n8594), .B2(keyinput99), .C1(n8681), .C2(keyinput76), 
        .A(n8593), .ZN(n8595) );
  NOR4_X1 U10058 ( .A1(n8598), .A2(n8597), .A3(n8596), .A4(n8595), .ZN(n8599)
         );
  NAND4_X1 U10059 ( .A1(n8602), .A2(n8601), .A3(n8600), .A4(n8599), .ZN(n8603)
         );
  NOR3_X1 U10060 ( .A1(n8605), .A2(n8604), .A3(n8603), .ZN(n8606) );
  XOR2_X1 U10061 ( .A(n8607), .B(n8606), .Z(n8608) );
  XNOR2_X1 U10062 ( .A(n8609), .B(n8608), .ZN(P2_U3519) );
  MUX2_X1 U10063 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n8610), .S(n10117), .Z(
        P2_U3518) );
  MUX2_X1 U10064 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n8611), .S(n10117), .Z(
        P2_U3517) );
  MUX2_X1 U10065 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n8613), .S(n10117), .Z(
        P2_U3515) );
  MUX2_X1 U10066 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n8614), .S(n10117), .Z(
        P2_U3514) );
  MUX2_X1 U10067 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n8615), .S(n10117), .Z(
        P2_U3513) );
  MUX2_X1 U10068 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n8616), .S(n10117), .Z(
        P2_U3512) );
  MUX2_X1 U10069 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n8617), .S(n10117), .Z(
        P2_U3511) );
  MUX2_X1 U10070 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n8618), .S(n10117), .Z(
        P2_U3510) );
  MUX2_X1 U10071 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n8619), .S(n10117), .Z(
        P2_U3509) );
  MUX2_X1 U10072 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n8620), .S(n10117), .Z(
        P2_U3508) );
  MUX2_X1 U10073 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n8621), .S(n10117), .Z(
        P2_U3507) );
  MUX2_X1 U10074 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n8622), .S(n10117), .Z(
        P2_U3505) );
  MUX2_X1 U10075 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n8623), .S(n10117), .Z(
        P2_U3502) );
  MUX2_X1 U10076 ( .A(n8624), .B(P2_REG0_REG_16__SCAN_IN), .S(n10115), .Z(
        P2_U3499) );
  NAND3_X1 U10077 ( .A1(n8626), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .ZN(n8628) );
  OAI22_X1 U10078 ( .A1(n8625), .A2(n8628), .B1(n6451), .B2(n8627), .ZN(n8629)
         );
  AOI21_X1 U10079 ( .B1(n9623), .B2(n8630), .A(n8629), .ZN(n8631) );
  INV_X1 U10080 ( .A(n8631), .ZN(P2_U3327) );
  AOI21_X1 U10081 ( .B1(n8633), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n8632), .ZN(
        n8634) );
  OAI21_X1 U10082 ( .B1(n8636), .B2(n8635), .A(n8634), .ZN(P2_U3330) );
  MUX2_X1 U10083 ( .A(n8637), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  AND3_X1 U10084 ( .A1(n6990), .A2(n8639), .A3(n8638), .ZN(n8640) );
  OAI21_X1 U10085 ( .B1(n8641), .B2(n8640), .A(n8783), .ZN(n8650) );
  NOR2_X1 U10086 ( .A1(n8798), .A2(n8642), .ZN(n8643) );
  AOI211_X1 U10087 ( .C1(n8800), .C2(n9099), .A(n8644), .B(n8643), .ZN(n8649)
         );
  INV_X1 U10088 ( .A(n8645), .ZN(n8647) );
  AOI22_X1 U10089 ( .A1(n8789), .A2(n8647), .B1(n8804), .B2(n8646), .ZN(n8648)
         );
  NAND3_X1 U10090 ( .A1(n8650), .A2(n8649), .A3(n8648), .ZN(P1_U3211) );
  NAND2_X1 U10091 ( .A1(n8652), .A2(n8651), .ZN(n8653) );
  XOR2_X1 U10092 ( .A(n8654), .B(n8653), .Z(n8661) );
  NOR2_X1 U10093 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8655), .ZN(n9797) );
  NOR2_X1 U10094 ( .A1(n8798), .A2(n8842), .ZN(n8656) );
  AOI211_X1 U10095 ( .C1(n8800), .C2(n9452), .A(n9797), .B(n8656), .ZN(n8657)
         );
  OAI21_X1 U10096 ( .B1(n8658), .B2(n8802), .A(n8657), .ZN(n8659) );
  AOI21_X1 U10097 ( .B1(n8804), .B2(n9199), .A(n8659), .ZN(n8660) );
  OAI21_X1 U10098 ( .B1(n8661), .B2(n8806), .A(n8660), .ZN(P1_U3213) );
  NAND2_X1 U10099 ( .A1(n8663), .A2(n8662), .ZN(n8664) );
  XOR2_X1 U10100 ( .A(n8665), .B(n8664), .Z(n8670) );
  AOI22_X1 U10101 ( .A1(n8774), .A2(n9358), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3084), .ZN(n8667) );
  NAND2_X1 U10102 ( .A1(n9336), .A2(n8800), .ZN(n8666) );
  OAI211_X1 U10103 ( .C1(n8802), .C2(n9330), .A(n8667), .B(n8666), .ZN(n8668)
         );
  AOI21_X1 U10104 ( .B1(n9534), .B2(n8804), .A(n8668), .ZN(n8669) );
  OAI21_X1 U10105 ( .B1(n8670), .B2(n8806), .A(n8669), .ZN(P1_U3214) );
  XOR2_X1 U10106 ( .A(n8672), .B(n8671), .Z(n8673) );
  XNOR2_X1 U10107 ( .A(n8674), .B(n8673), .ZN(n8679) );
  NAND2_X1 U10108 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9183) );
  OAI21_X1 U10109 ( .B1(n8786), .B2(n9207), .A(n9183), .ZN(n8675) );
  AOI21_X1 U10110 ( .B1(n8774), .B2(n9436), .A(n8675), .ZN(n8676) );
  OAI21_X1 U10111 ( .B1(n9389), .B2(n8802), .A(n8676), .ZN(n8677) );
  AOI21_X1 U10112 ( .B1(n9554), .B2(n8804), .A(n8677), .ZN(n8678) );
  OAI21_X1 U10113 ( .B1(n8679), .B2(n8806), .A(n8678), .ZN(P1_U3217) );
  NAND2_X1 U10114 ( .A1(n8680), .A2(n8866), .ZN(n8683) );
  OR2_X1 U10115 ( .A1(n8869), .A2(n8681), .ZN(n8682) );
  NAND2_X1 U10116 ( .A1(n9512), .A2(n8684), .ZN(n8686) );
  NAND2_X1 U10117 ( .A1(n9279), .A2(n5845), .ZN(n8685) );
  NAND2_X1 U10118 ( .A1(n8686), .A2(n8685), .ZN(n8688) );
  XNOR2_X1 U10119 ( .A(n8688), .B(n5830), .ZN(n8691) );
  AOI22_X1 U10120 ( .A1(n9512), .A2(n5845), .B1(n8689), .B2(n9279), .ZN(n8690)
         );
  XNOR2_X1 U10121 ( .A(n8691), .B(n8690), .ZN(n8705) );
  NAND3_X1 U10122 ( .A1(n8692), .A2(n8783), .A3(n8705), .ZN(n8708) );
  OR2_X1 U10123 ( .A1(n9220), .A2(n4386), .ZN(n8699) );
  NAND2_X1 U10124 ( .A1(n8694), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n8696) );
  NAND2_X1 U10125 ( .A1(n5868), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n8695) );
  OAI211_X1 U10126 ( .C1(n6050), .C2(n8473), .A(n8696), .B(n8695), .ZN(n8697)
         );
  INV_X1 U10127 ( .A(n8697), .ZN(n8698) );
  INV_X1 U10128 ( .A(n9261), .ZN(n9094) );
  AOI22_X1 U10129 ( .A1(n9094), .A2(n8800), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n8702) );
  INV_X1 U10130 ( .A(n8700), .ZN(n9264) );
  NAND2_X1 U10131 ( .A1(n9264), .A2(n8789), .ZN(n8701) );
  OAI211_X1 U10132 ( .C1(n9289), .C2(n8798), .A(n8702), .B(n8701), .ZN(n8703)
         );
  AOI21_X1 U10133 ( .B1(n9512), .B2(n8804), .A(n8703), .ZN(n8707) );
  NAND3_X1 U10134 ( .A1(n8705), .A2(n8704), .A3(n8783), .ZN(n8706) );
  NAND4_X1 U10135 ( .A1(n8709), .A2(n8708), .A3(n8707), .A4(n8706), .ZN(
        P1_U3218) );
  NAND2_X1 U10136 ( .A1(n9368), .A2(n9892), .ZN(n9546) );
  INV_X1 U10137 ( .A(n8710), .ZN(n8711) );
  NAND2_X1 U10138 ( .A1(n8712), .A2(n8711), .ZN(n8721) );
  OAI21_X1 U10139 ( .B1(n8715), .B2(n8713), .A(n8714), .ZN(n8716) );
  NAND2_X1 U10140 ( .A1(n8716), .A2(n8783), .ZN(n8720) );
  AOI22_X1 U10141 ( .A1(n8774), .A2(n9396), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3084), .ZN(n8717) );
  OAI21_X1 U10142 ( .B1(n9210), .B2(n8786), .A(n8717), .ZN(n8718) );
  AOI21_X1 U10143 ( .B1(n9362), .B2(n8789), .A(n8718), .ZN(n8719) );
  OAI211_X1 U10144 ( .C1(n9546), .C2(n8721), .A(n8720), .B(n8719), .ZN(
        P1_U3221) );
  NOR2_X1 U10145 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8722), .ZN(n9116) );
  NOR2_X1 U10146 ( .A1(n8786), .A2(n8842), .ZN(n8723) );
  AOI211_X1 U10147 ( .C1(n8774), .C2(n9096), .A(n9116), .B(n8723), .ZN(n8724)
         );
  OAI21_X1 U10148 ( .B1(n8725), .B2(n8802), .A(n8724), .ZN(n8732) );
  OAI21_X1 U10149 ( .B1(n8728), .B2(n8727), .A(n8726), .ZN(n8730) );
  AOI21_X1 U10150 ( .B1(n8730), .B2(n8729), .A(n8806), .ZN(n8731) );
  AOI211_X1 U10151 ( .C1(n8804), .C2(n9586), .A(n8732), .B(n8731), .ZN(n8733)
         );
  INV_X1 U10152 ( .A(n8733), .ZN(P1_U3222) );
  OAI21_X1 U10153 ( .B1(n8736), .B2(n8734), .A(n8735), .ZN(n8737) );
  NAND2_X1 U10154 ( .A1(n8737), .A2(n8783), .ZN(n8742) );
  INV_X1 U10155 ( .A(n8738), .ZN(n9300) );
  AOI22_X1 U10156 ( .A1(n9336), .A2(n8774), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3084), .ZN(n8739) );
  OAI21_X1 U10157 ( .B1(n8859), .B2(n8786), .A(n8739), .ZN(n8740) );
  AOI21_X1 U10158 ( .B1(n9300), .B2(n8789), .A(n8740), .ZN(n8741) );
  OAI211_X1 U10159 ( .C1(n9302), .C2(n8792), .A(n8742), .B(n8741), .ZN(
        P1_U3223) );
  NAND2_X1 U10160 ( .A1(n8744), .A2(n8743), .ZN(n8745) );
  XOR2_X1 U10161 ( .A(n8746), .B(n8745), .Z(n8751) );
  NAND2_X1 U10162 ( .A1(P1_U3084), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9153) );
  OAI21_X1 U10163 ( .B1(n8786), .B2(n9204), .A(n9153), .ZN(n8747) );
  AOI21_X1 U10164 ( .B1(n8774), .B2(n9467), .A(n8747), .ZN(n8748) );
  OAI21_X1 U10165 ( .B1(n9430), .B2(n8802), .A(n8748), .ZN(n8749) );
  AOI21_X1 U10166 ( .B1(n9564), .B2(n8804), .A(n8749), .ZN(n8750) );
  OAI21_X1 U10167 ( .B1(n8751), .B2(n8806), .A(n8750), .ZN(P1_U3226) );
  INV_X1 U10168 ( .A(n8752), .ZN(n8753) );
  AOI21_X1 U10169 ( .B1(n8755), .B2(n8754), .A(n8753), .ZN(n8760) );
  AOI22_X1 U10170 ( .A1(n9316), .A2(n8800), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3084), .ZN(n8757) );
  NAND2_X1 U10171 ( .A1(n8789), .A2(n9320), .ZN(n8756) );
  OAI211_X1 U10172 ( .C1(n9212), .C2(n8798), .A(n8757), .B(n8756), .ZN(n8758)
         );
  AOI21_X1 U10173 ( .B1(n9530), .B2(n8804), .A(n8758), .ZN(n8759) );
  OAI21_X1 U10174 ( .B1(n8760), .B2(n8806), .A(n8759), .ZN(P1_U3227) );
  AOI21_X1 U10175 ( .B1(n8762), .B2(n8761), .A(n4418), .ZN(n8768) );
  INV_X1 U10176 ( .A(n9421), .ZN(n9205) );
  OAI22_X1 U10177 ( .A1(n8786), .A2(n9382), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8763), .ZN(n8764) );
  AOI21_X1 U10178 ( .B1(n8774), .B2(n9205), .A(n8764), .ZN(n8765) );
  OAI21_X1 U10179 ( .B1(n9375), .B2(n8802), .A(n8765), .ZN(n8766) );
  AOI21_X1 U10180 ( .B1(n9551), .B2(n8804), .A(n8766), .ZN(n8767) );
  OAI21_X1 U10181 ( .B1(n8768), .B2(n8806), .A(n8767), .ZN(P1_U3231) );
  NAND2_X1 U10182 ( .A1(n8770), .A2(n8769), .ZN(n8771) );
  XOR2_X1 U10183 ( .A(n8772), .B(n8771), .Z(n8779) );
  INV_X1 U10184 ( .A(n9382), .ZN(n9350) );
  AOI22_X1 U10185 ( .A1(n8774), .A2(n9350), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3084), .ZN(n8776) );
  NAND2_X1 U10186 ( .A1(n9349), .A2(n8800), .ZN(n8775) );
  OAI211_X1 U10187 ( .C1(n8802), .C2(n9343), .A(n8776), .B(n8775), .ZN(n8777)
         );
  AOI21_X1 U10188 ( .B1(n9539), .B2(n8804), .A(n8777), .ZN(n8778) );
  OAI21_X1 U10189 ( .B1(n8779), .B2(n8806), .A(n8778), .ZN(P1_U3233) );
  INV_X1 U10190 ( .A(n8735), .ZN(n8782) );
  OAI21_X1 U10191 ( .B1(n8782), .B2(n8781), .A(n8780), .ZN(n8784) );
  NAND3_X1 U10192 ( .A1(n8784), .A2(n8783), .A3(n6286), .ZN(n8791) );
  OAI22_X1 U10193 ( .A1(n9288), .A2(n8798), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8785), .ZN(n8788) );
  NOR2_X1 U10194 ( .A1(n9289), .A2(n8786), .ZN(n8787) );
  AOI211_X1 U10195 ( .C1(n8789), .C2(n9292), .A(n8788), .B(n8787), .ZN(n8790)
         );
  OAI211_X1 U10196 ( .C1(n9295), .C2(n8792), .A(n8791), .B(n8790), .ZN(
        P1_U3238) );
  NAND2_X1 U10197 ( .A1(n8794), .A2(n8793), .ZN(n8795) );
  XOR2_X1 U10198 ( .A(n8796), .B(n8795), .Z(n8807) );
  OAI21_X1 U10199 ( .B1(n8798), .B2(n9200), .A(n8797), .ZN(n8799) );
  AOI21_X1 U10200 ( .B1(n8800), .B2(n9467), .A(n8799), .ZN(n8801) );
  OAI21_X1 U10201 ( .B1(n9461), .B2(n8802), .A(n8801), .ZN(n8803) );
  AOI21_X1 U10202 ( .B1(n9574), .B2(n8804), .A(n8803), .ZN(n8805) );
  OAI21_X1 U10203 ( .B1(n8807), .B2(n8806), .A(n8805), .ZN(P1_U3239) );
  NOR2_X1 U10204 ( .A1(n8869), .A2(n6435), .ZN(n8808) );
  INV_X1 U10205 ( .A(n9498), .ZN(n8992) );
  INV_X1 U10206 ( .A(n9190), .ZN(n8809) );
  AND2_X1 U10207 ( .A1(n8992), .A2(n8809), .ZN(n8997) );
  NAND2_X1 U10208 ( .A1(n8810), .A2(n8866), .ZN(n8813) );
  OR2_X1 U10209 ( .A1(n8869), .A2(n8811), .ZN(n8812) );
  INV_X1 U10210 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n8817) );
  NAND2_X1 U10211 ( .A1(n8814), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n8816) );
  NAND2_X1 U10212 ( .A1(n5868), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n8815) );
  OAI211_X1 U10213 ( .C1(n6254), .C2(n8817), .A(n8816), .B(n8815), .ZN(n9246)
         );
  INV_X1 U10214 ( .A(n9246), .ZN(n8872) );
  NOR2_X1 U10215 ( .A1(n9193), .A2(n8872), .ZN(n8990) );
  NOR2_X1 U10216 ( .A1(n8997), .A2(n8990), .ZN(n9040) );
  OR2_X1 U10217 ( .A1(n9521), .A2(n8859), .ZN(n9242) );
  AND2_X1 U10218 ( .A1(n9242), .A2(n9238), .ZN(n8818) );
  NAND2_X1 U10219 ( .A1(n9257), .A2(n8818), .ZN(n8858) );
  NAND2_X1 U10220 ( .A1(n9312), .A2(n9336), .ZN(n8879) );
  NOR2_X1 U10221 ( .A1(n9534), .A2(n9212), .ZN(n9237) );
  INV_X1 U10222 ( .A(n9237), .ZN(n9005) );
  NAND2_X1 U10223 ( .A1(n8879), .A2(n9005), .ZN(n8966) );
  NOR2_X1 U10224 ( .A1(n8858), .A2(n8966), .ZN(n8857) );
  OR2_X1 U10225 ( .A1(n9539), .A2(n9210), .ZN(n9235) );
  OR2_X1 U10226 ( .A1(n9368), .A2(n9382), .ZN(n9007) );
  NAND2_X1 U10227 ( .A1(n9235), .A2(n9007), .ZN(n8958) );
  OR2_X1 U10228 ( .A1(n9561), .A2(n9204), .ZN(n9010) );
  OR2_X1 U10229 ( .A1(n9564), .A2(n9423), .ZN(n9415) );
  NAND2_X1 U10230 ( .A1(n9010), .A2(n9415), .ZN(n9227) );
  INV_X1 U10231 ( .A(n9227), .ZN(n8819) );
  NAND2_X1 U10232 ( .A1(n9554), .A2(n9421), .ZN(n9230) );
  NAND2_X1 U10233 ( .A1(n9561), .A2(n9204), .ZN(n9228) );
  NAND2_X1 U10234 ( .A1(n9230), .A2(n9228), .ZN(n8951) );
  OR2_X1 U10235 ( .A1(n9551), .A2(n9207), .ZN(n9231) );
  OR2_X1 U10236 ( .A1(n9554), .A2(n9421), .ZN(n9009) );
  AND2_X1 U10237 ( .A1(n9231), .A2(n9009), .ZN(n8952) );
  OAI21_X1 U10238 ( .B1(n8819), .B2(n8951), .A(n8952), .ZN(n8822) );
  AND2_X1 U10239 ( .A1(n9539), .A2(n9210), .ZN(n9234) );
  AND2_X1 U10240 ( .A1(n9551), .A2(n9207), .ZN(n9232) );
  NAND2_X1 U10241 ( .A1(n9007), .A2(n9232), .ZN(n8820) );
  NAND2_X1 U10242 ( .A1(n9368), .A2(n9382), .ZN(n9233) );
  NAND2_X1 U10243 ( .A1(n8820), .A2(n9233), .ZN(n8821) );
  OR2_X1 U10244 ( .A1(n9234), .A2(n8821), .ZN(n8824) );
  NAND2_X1 U10245 ( .A1(n8824), .A2(n9235), .ZN(n8963) );
  OAI21_X1 U10246 ( .B1(n8958), .B2(n8822), .A(n8963), .ZN(n8823) );
  NAND2_X1 U10247 ( .A1(n8857), .A2(n8823), .ZN(n9059) );
  INV_X1 U10248 ( .A(n9059), .ZN(n8865) );
  INV_X1 U10249 ( .A(n9230), .ZN(n8948) );
  NOR2_X1 U10250 ( .A1(n8824), .A2(n8948), .ZN(n9061) );
  NAND2_X1 U10251 ( .A1(n9564), .A2(n9423), .ZN(n9414) );
  NAND2_X1 U10252 ( .A1(n9228), .A2(n9414), .ZN(n8944) );
  NAND2_X1 U10253 ( .A1(n9570), .A2(n8852), .ZN(n9413) );
  INV_X1 U10254 ( .A(n9413), .ZN(n8825) );
  NOR2_X1 U10255 ( .A1(n8944), .A2(n8825), .ZN(n9229) );
  NAND2_X1 U10256 ( .A1(n8843), .A2(n8826), .ZN(n8928) );
  INV_X1 U10257 ( .A(n8827), .ZN(n8828) );
  NAND2_X1 U10258 ( .A1(n8922), .A2(n8828), .ZN(n8930) );
  NOR2_X1 U10259 ( .A1(n8930), .A2(n4709), .ZN(n8845) );
  NAND3_X1 U10260 ( .A1(n8845), .A2(n8913), .A3(n8900), .ZN(n8830) );
  NOR2_X1 U10261 ( .A1(n8928), .A2(n8830), .ZN(n8831) );
  NAND2_X1 U10262 ( .A1(n9574), .A2(n9201), .ZN(n9226) );
  AND2_X1 U10263 ( .A1(n8831), .A2(n9226), .ZN(n8832) );
  NAND2_X1 U10264 ( .A1(n9229), .A2(n8832), .ZN(n9058) );
  AND2_X1 U10265 ( .A1(n8833), .A2(n8887), .ZN(n9045) );
  INV_X1 U10266 ( .A(n9045), .ZN(n8839) );
  AOI21_X1 U10267 ( .B1(n9104), .B2(n9850), .A(n9069), .ZN(n8837) );
  INV_X1 U10268 ( .A(n8834), .ZN(n8835) );
  NAND4_X1 U10269 ( .A1(n8837), .A2(n9044), .A3(n8836), .A4(n8835), .ZN(n8838)
         );
  OR2_X1 U10270 ( .A1(n8839), .A2(n8838), .ZN(n8840) );
  INV_X1 U10271 ( .A(n8902), .ZN(n9053) );
  AOI21_X1 U10272 ( .B1(n8841), .B2(n8840), .A(n9053), .ZN(n8855) );
  AND2_X1 U10273 ( .A1(n9464), .A2(n9452), .ZN(n9225) );
  OR2_X1 U10274 ( .A1(n9579), .A2(n8842), .ZN(n8924) );
  OR2_X1 U10275 ( .A1(n9225), .A2(n8844), .ZN(n8883) );
  INV_X1 U10276 ( .A(n8928), .ZN(n8927) );
  INV_X1 U10277 ( .A(n8845), .ZN(n8849) );
  AND2_X1 U10278 ( .A1(n8909), .A2(n8917), .ZN(n8848) );
  INV_X1 U10279 ( .A(n8922), .ZN(n8846) );
  OAI21_X1 U10280 ( .B1(n8849), .B2(n8848), .A(n8925), .ZN(n8850) );
  AND2_X1 U10281 ( .A1(n8927), .A2(n8850), .ZN(n8851) );
  OAI21_X1 U10282 ( .B1(n8883), .B2(n8851), .A(n9226), .ZN(n8853) );
  OR2_X1 U10283 ( .A1(n9570), .A2(n8852), .ZN(n8941) );
  NAND2_X1 U10284 ( .A1(n8853), .A2(n8941), .ZN(n8854) );
  NAND2_X1 U10285 ( .A1(n9229), .A2(n8854), .ZN(n9056) );
  OAI21_X1 U10286 ( .B1(n9058), .B2(n8855), .A(n9056), .ZN(n8856) );
  NAND2_X1 U10287 ( .A1(n9061), .A2(n8856), .ZN(n8864) );
  INV_X1 U10288 ( .A(n8857), .ZN(n8863) );
  NAND2_X1 U10289 ( .A1(n9534), .A2(n9212), .ZN(n9236) );
  INV_X1 U10290 ( .A(n8858), .ZN(n8861) );
  NAND2_X1 U10291 ( .A1(n9524), .A2(n9288), .ZN(n9004) );
  NAND2_X1 U10292 ( .A1(n9530), .A2(n9214), .ZN(n9303) );
  AND2_X1 U10293 ( .A1(n9004), .A2(n9303), .ZN(n9240) );
  INV_X1 U10294 ( .A(n9240), .ZN(n8860) );
  AND2_X1 U10295 ( .A1(n9521), .A2(n8859), .ZN(n9241) );
  AOI22_X1 U10296 ( .A1(n8861), .A2(n8860), .B1(n9241), .B2(n9257), .ZN(n8862)
         );
  NAND2_X1 U10297 ( .A1(n9512), .A2(n9217), .ZN(n9243) );
  NAND2_X1 U10298 ( .A1(n9514), .A2(n9289), .ZN(n9003) );
  AND2_X1 U10299 ( .A1(n9243), .A2(n9003), .ZN(n8976) );
  OAI211_X1 U10300 ( .C1(n8863), .C2(n9236), .A(n8862), .B(n8976), .ZN(n9062)
         );
  AOI21_X1 U10301 ( .B1(n8865), .B2(n8864), .A(n9062), .ZN(n8874) );
  NAND2_X1 U10302 ( .A1(n8867), .A2(n8866), .ZN(n8871) );
  OR2_X1 U10303 ( .A1(n8869), .A2(n8868), .ZN(n8870) );
  NAND2_X1 U10304 ( .A1(n8978), .A2(n9002), .ZN(n9066) );
  AND2_X1 U10305 ( .A1(n9193), .A2(n8872), .ZN(n9039) );
  INV_X1 U10306 ( .A(n9039), .ZN(n8873) );
  NAND2_X1 U10307 ( .A1(n9507), .A2(n9261), .ZN(n9065) );
  OAI211_X1 U10308 ( .C1(n8874), .C2(n9066), .A(n8873), .B(n9065), .ZN(n8875)
         );
  AND2_X1 U10309 ( .A1(n9498), .A2(n9190), .ZN(n9068) );
  AOI21_X1 U10310 ( .B1(n9040), .B2(n8875), .A(n9068), .ZN(n9083) );
  NOR2_X1 U10311 ( .A1(n9083), .A2(n9321), .ZN(n9082) );
  INV_X1 U10312 ( .A(n9215), .ZN(n8876) );
  INV_X1 U10313 ( .A(n9285), .ZN(n9036) );
  NAND2_X1 U10314 ( .A1(n8966), .A2(n9303), .ZN(n8877) );
  NAND2_X1 U10315 ( .A1(n8877), .A2(n9238), .ZN(n8882) );
  INV_X1 U10316 ( .A(n9236), .ZN(n8878) );
  NAND2_X1 U10317 ( .A1(n8879), .A2(n8878), .ZN(n8880) );
  NAND2_X1 U10318 ( .A1(n9240), .A2(n8880), .ZN(n8881) );
  INV_X1 U10319 ( .A(n8995), .ZN(n8996) );
  MUX2_X1 U10320 ( .A(n8882), .B(n8881), .S(n8996), .Z(n8970) );
  INV_X1 U10321 ( .A(n8883), .ZN(n8938) );
  NAND2_X1 U10322 ( .A1(n8888), .A2(n9049), .ZN(n8886) );
  INV_X1 U10323 ( .A(n8884), .ZN(n8890) );
  NAND2_X1 U10324 ( .A1(n8891), .A2(n8887), .ZN(n9047) );
  INV_X1 U10325 ( .A(n9047), .ZN(n8885) );
  OAI22_X1 U10326 ( .A1(n8889), .A2(n8886), .B1(n8890), .B2(n8885), .ZN(n8896)
         );
  NAND3_X1 U10327 ( .A1(n8889), .A2(n8888), .A3(n8887), .ZN(n8894) );
  AOI21_X1 U10328 ( .B1(n8892), .B2(n8891), .A(n8890), .ZN(n8893) );
  NAND2_X1 U10329 ( .A1(n8894), .A2(n8893), .ZN(n8895) );
  INV_X1 U10330 ( .A(n8897), .ZN(n9019) );
  NAND3_X1 U10331 ( .A1(n8898), .A2(n9019), .A3(n9018), .ZN(n8907) );
  INV_X1 U10332 ( .A(n9050), .ZN(n8899) );
  AOI21_X1 U10333 ( .B1(n8899), .B2(n8900), .A(n9053), .ZN(n8905) );
  NAND2_X1 U10334 ( .A1(n8901), .A2(n8900), .ZN(n8903) );
  NAND2_X1 U10335 ( .A1(n8903), .A2(n8902), .ZN(n8904) );
  MUX2_X1 U10336 ( .A(n8905), .B(n8904), .S(n8995), .Z(n8906) );
  NAND2_X1 U10337 ( .A1(n8907), .A2(n8906), .ZN(n8912) );
  NAND2_X1 U10338 ( .A1(n8912), .A2(n8913), .ZN(n8910) );
  AOI21_X1 U10339 ( .B1(n8910), .B2(n8909), .A(n8908), .ZN(n8937) );
  NAND2_X1 U10340 ( .A1(n8912), .A2(n8911), .ZN(n8915) );
  NAND3_X1 U10341 ( .A1(n8915), .A2(n8914), .A3(n8913), .ZN(n8919) );
  AND4_X1 U10342 ( .A1(n8924), .A2(n8917), .A3(n8916), .A4(n8995), .ZN(n8918)
         );
  NAND4_X1 U10343 ( .A1(n8919), .A2(n8918), .A3(n8925), .A4(n9223), .ZN(n8935)
         );
  NAND4_X1 U10344 ( .A1(n8922), .A2(n8921), .A3(n8995), .A4(n8920), .ZN(n8923)
         );
  OAI211_X1 U10345 ( .C1(n8925), .C2(n8996), .A(n8924), .B(n8923), .ZN(n8926)
         );
  NAND2_X1 U10346 ( .A1(n8927), .A2(n8926), .ZN(n8933) );
  NAND2_X1 U10347 ( .A1(n8928), .A2(n8996), .ZN(n8932) );
  NAND3_X1 U10348 ( .A1(n8930), .A2(n8996), .A3(n8929), .ZN(n8931) );
  NAND4_X1 U10349 ( .A1(n8933), .A2(n9223), .A3(n8932), .A4(n8931), .ZN(n8934)
         );
  NAND2_X1 U10350 ( .A1(n8935), .A2(n8934), .ZN(n8936) );
  NAND2_X1 U10351 ( .A1(n8941), .A2(n9413), .ZN(n9441) );
  INV_X1 U10352 ( .A(n9441), .ZN(n9451) );
  MUX2_X1 U10353 ( .A(n9226), .B(n4729), .S(n8995), .Z(n8939) );
  NAND3_X1 U10354 ( .A1(n8940), .A2(n9451), .A3(n8939), .ZN(n8943) );
  NAND2_X1 U10355 ( .A1(n9415), .A2(n9414), .ZN(n9031) );
  MUX2_X1 U10356 ( .A(n8941), .B(n9413), .S(n8995), .Z(n8942) );
  NAND3_X1 U10357 ( .A1(n8943), .A2(n9434), .A3(n8942), .ZN(n8947) );
  MUX2_X1 U10358 ( .A(n8944), .B(n9227), .S(n8995), .Z(n8945) );
  INV_X1 U10359 ( .A(n8945), .ZN(n8946) );
  NAND2_X1 U10360 ( .A1(n8947), .A2(n8946), .ZN(n8955) );
  AND2_X1 U10361 ( .A1(n9009), .A2(n9010), .ZN(n8950) );
  OR2_X1 U10362 ( .A1(n9232), .A2(n8948), .ZN(n8949) );
  AOI21_X1 U10363 ( .B1(n8955), .B2(n8950), .A(n8949), .ZN(n8957) );
  INV_X1 U10364 ( .A(n8951), .ZN(n8954) );
  INV_X1 U10365 ( .A(n8952), .ZN(n8953) );
  AOI21_X1 U10366 ( .B1(n8955), .B2(n8954), .A(n8953), .ZN(n8956) );
  INV_X1 U10367 ( .A(n9231), .ZN(n9008) );
  OAI21_X1 U10368 ( .B1(n8961), .B2(n9008), .A(n9233), .ZN(n8959) );
  INV_X1 U10369 ( .A(n8958), .ZN(n8960) );
  NAND2_X1 U10370 ( .A1(n8961), .A2(n8960), .ZN(n8962) );
  NAND4_X1 U10371 ( .A1(n9303), .A2(n8963), .A3(n9236), .A4(n8962), .ZN(n8964)
         );
  MUX2_X1 U10372 ( .A(n9238), .B(n9004), .S(n8995), .Z(n8968) );
  OAI21_X1 U10373 ( .B1(n8970), .B2(n8969), .A(n8968), .ZN(n8971) );
  INV_X1 U10374 ( .A(n9241), .ZN(n8972) );
  MUX2_X1 U10375 ( .A(n9242), .B(n8972), .S(n8995), .Z(n8973) );
  NAND2_X1 U10376 ( .A1(n8974), .A2(n8973), .ZN(n8975) );
  NAND2_X1 U10377 ( .A1(n8975), .A2(n9257), .ZN(n8982) );
  NAND2_X1 U10378 ( .A1(n8982), .A2(n8976), .ZN(n8977) );
  NAND2_X1 U10379 ( .A1(n8977), .A2(n9002), .ZN(n8980) );
  INV_X1 U10380 ( .A(n8978), .ZN(n8979) );
  AOI21_X1 U10381 ( .B1(n8980), .B2(n9218), .A(n8979), .ZN(n8987) );
  INV_X1 U10382 ( .A(n9003), .ZN(n8981) );
  OAI211_X1 U10383 ( .C1(n8982), .C2(n8981), .A(n9257), .B(n9002), .ZN(n8983)
         );
  NAND2_X1 U10384 ( .A1(n8983), .A2(n9243), .ZN(n8985) );
  INV_X1 U10385 ( .A(n9065), .ZN(n8984) );
  AOI21_X1 U10386 ( .B1(n8985), .B2(n9218), .A(n8984), .ZN(n8986) );
  NAND2_X1 U10387 ( .A1(n9246), .A2(n9190), .ZN(n8988) );
  NAND2_X1 U10388 ( .A1(n9193), .A2(n8988), .ZN(n9064) );
  NAND2_X1 U10389 ( .A1(n8989), .A2(n9064), .ZN(n8994) );
  INV_X1 U10390 ( .A(n8990), .ZN(n8991) );
  NAND2_X1 U10391 ( .A1(n8991), .A2(n9190), .ZN(n8993) );
  NAND2_X1 U10392 ( .A1(n8993), .A2(n8992), .ZN(n9071) );
  INV_X1 U10393 ( .A(n9068), .ZN(n9076) );
  OAI21_X1 U10394 ( .B1(n8996), .B2(n9064), .A(n9076), .ZN(n8999) );
  INV_X1 U10395 ( .A(n8997), .ZN(n8998) );
  NAND2_X1 U10396 ( .A1(n8999), .A2(n8998), .ZN(n9000) );
  NAND2_X1 U10397 ( .A1(n9001), .A2(n9000), .ZN(n9077) );
  INV_X1 U10398 ( .A(n9218), .ZN(n9244) );
  NAND2_X1 U10399 ( .A1(n9002), .A2(n9243), .ZN(n9254) );
  INV_X1 U10400 ( .A(n9254), .ZN(n9256) );
  NAND2_X1 U10401 ( .A1(n9257), .A2(n9003), .ZN(n9277) );
  INV_X1 U10402 ( .A(n9277), .ZN(n9269) );
  XNOR2_X1 U10403 ( .A(n9530), .B(n9336), .ZN(n9314) );
  INV_X1 U10404 ( .A(n9314), .ZN(n9035) );
  NAND2_X1 U10405 ( .A1(n9005), .A2(n9236), .ZN(n9334) );
  INV_X1 U10406 ( .A(n9235), .ZN(n9006) );
  NOR2_X1 U10407 ( .A1(n9006), .A2(n9234), .ZN(n9347) );
  NAND2_X1 U10408 ( .A1(n9007), .A2(n9233), .ZN(n9363) );
  INV_X1 U10409 ( .A(n9363), .ZN(n9033) );
  NOR2_X1 U10410 ( .A1(n9008), .A2(n9232), .ZN(n9380) );
  INV_X1 U10411 ( .A(n9395), .ZN(n9385) );
  NAND2_X1 U10412 ( .A1(n9010), .A2(n9228), .ZN(n9418) );
  INV_X1 U10413 ( .A(n9226), .ZN(n9011) );
  NOR2_X1 U10414 ( .A1(n9225), .A2(n9011), .ZN(n9466) );
  NAND2_X1 U10415 ( .A1(n9013), .A2(n9012), .ZN(n9016) );
  NOR4_X1 U10416 ( .A1(n9016), .A2(n4599), .A3(n9015), .A4(n9014), .ZN(n9020)
         );
  NAND4_X1 U10417 ( .A1(n9020), .A2(n9019), .A3(n9018), .A4(n9017), .ZN(n9024)
         );
  OR4_X1 U10418 ( .A1(n9024), .A2(n9023), .A3(n9022), .A4(n9021), .ZN(n9028)
         );
  NOR4_X1 U10419 ( .A1(n9028), .A2(n9027), .A3(n9026), .A4(n9025), .ZN(n9029)
         );
  NAND4_X1 U10420 ( .A1(n9451), .A2(n9466), .A3(n9029), .A4(n9482), .ZN(n9030)
         );
  NOR4_X1 U10421 ( .A1(n9385), .A2(n9031), .A3(n9418), .A4(n9030), .ZN(n9032)
         );
  NAND4_X1 U10422 ( .A1(n9347), .A2(n9033), .A3(n9380), .A4(n9032), .ZN(n9034)
         );
  NOR4_X1 U10423 ( .A1(n9305), .A2(n9035), .A3(n9334), .A4(n9034), .ZN(n9037)
         );
  NAND4_X1 U10424 ( .A1(n9256), .A2(n9269), .A3(n9037), .A4(n9036), .ZN(n9038)
         );
  NOR4_X1 U10425 ( .A1(n9068), .A2(n9039), .A3(n9244), .A4(n9038), .ZN(n9041)
         );
  AOI21_X1 U10426 ( .B1(n9041), .B2(n9040), .A(n6309), .ZN(n9073) );
  INV_X1 U10427 ( .A(n9073), .ZN(n9042) );
  OAI21_X1 U10428 ( .B1(n9077), .B2(n9043), .A(n9042), .ZN(n9075) );
  NAND3_X1 U10429 ( .A1(n9046), .A2(n9045), .A3(n9044), .ZN(n9055) );
  AOI21_X1 U10430 ( .B1(n9049), .B2(n9048), .A(n9047), .ZN(n9052) );
  OAI21_X1 U10431 ( .B1(n9052), .B2(n9051), .A(n9050), .ZN(n9054) );
  AOI21_X1 U10432 ( .B1(n9055), .B2(n9054), .A(n9053), .ZN(n9057) );
  OAI21_X1 U10433 ( .B1(n9058), .B2(n9057), .A(n9056), .ZN(n9060) );
  AOI21_X1 U10434 ( .B1(n9061), .B2(n9060), .A(n9059), .ZN(n9063) );
  NOR2_X1 U10435 ( .A1(n9063), .A2(n9062), .ZN(n9067) );
  OAI211_X1 U10436 ( .C1(n9067), .C2(n9066), .A(n9065), .B(n9064), .ZN(n9070)
         );
  AOI211_X1 U10437 ( .C1(n9071), .C2(n9070), .A(n9069), .B(n9068), .ZN(n9072)
         );
  NOR2_X1 U10438 ( .A1(n9073), .A2(n9072), .ZN(n9074) );
  AND4_X1 U10439 ( .A1(n9077), .A2(n6309), .A3(n9076), .A4(n6308), .ZN(n9078)
         );
  NOR2_X1 U10440 ( .A1(n9079), .A2(n9078), .ZN(n9081) );
  INV_X1 U10441 ( .A(n9083), .ZN(n9086) );
  INV_X1 U10442 ( .A(n9090), .ZN(n9084) );
  OAI21_X1 U10443 ( .B1(n9086), .B2(n9085), .A(n9084), .ZN(n9092) );
  NAND4_X1 U10444 ( .A1(n9088), .A2(n9841), .A3(n9087), .A4(n9188), .ZN(n9089)
         );
  OAI211_X1 U10445 ( .C1(n6310), .C2(n9090), .A(n9089), .B(P1_B_REG_SCAN_IN), 
        .ZN(n9091) );
  OAI21_X1 U10446 ( .B1(n9093), .B2(n9092), .A(n9091), .ZN(P1_U3240) );
  MUX2_X1 U10447 ( .A(n9246), .B(P1_DATAO_REG_30__SCAN_IN), .S(n9105), .Z(
        P1_U3585) );
  MUX2_X1 U10448 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9094), .S(P1_U4006), .Z(
        P1_U3584) );
  MUX2_X1 U10449 ( .A(n9279), .B(P1_DATAO_REG_28__SCAN_IN), .S(n9105), .Z(
        P1_U3583) );
  MUX2_X1 U10450 ( .A(n9306), .B(P1_DATAO_REG_26__SCAN_IN), .S(n9105), .Z(
        P1_U3581) );
  MUX2_X1 U10451 ( .A(n9316), .B(P1_DATAO_REG_25__SCAN_IN), .S(n9105), .Z(
        P1_U3580) );
  MUX2_X1 U10452 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9336), .S(P1_U4006), .Z(
        P1_U3579) );
  MUX2_X1 U10453 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9349), .S(P1_U4006), .Z(
        P1_U3578) );
  MUX2_X1 U10454 ( .A(n9358), .B(P1_DATAO_REG_22__SCAN_IN), .S(n9105), .Z(
        P1_U3577) );
  MUX2_X1 U10455 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9350), .S(P1_U4006), .Z(
        P1_U3576) );
  MUX2_X1 U10456 ( .A(n9396), .B(P1_DATAO_REG_20__SCAN_IN), .S(n9105), .Z(
        P1_U3575) );
  MUX2_X1 U10457 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9205), .S(P1_U4006), .Z(
        P1_U3574) );
  MUX2_X1 U10458 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9436), .S(P1_U4006), .Z(
        P1_U3573) );
  MUX2_X1 U10459 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9453), .S(P1_U4006), .Z(
        P1_U3572) );
  MUX2_X1 U10460 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9467), .S(P1_U4006), .Z(
        P1_U3571) );
  MUX2_X1 U10461 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9452), .S(P1_U4006), .Z(
        P1_U3570) );
  MUX2_X1 U10462 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9485), .S(P1_U4006), .Z(
        P1_U3569) );
  MUX2_X1 U10463 ( .A(n9095), .B(P1_DATAO_REG_13__SCAN_IN), .S(n9105), .Z(
        P1_U3568) );
  MUX2_X1 U10464 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9487), .S(P1_U4006), .Z(
        P1_U3567) );
  MUX2_X1 U10465 ( .A(n9096), .B(P1_DATAO_REG_11__SCAN_IN), .S(n9105), .Z(
        P1_U3566) );
  MUX2_X1 U10466 ( .A(n9097), .B(P1_DATAO_REG_10__SCAN_IN), .S(n9105), .Z(
        P1_U3565) );
  MUX2_X1 U10467 ( .A(n9098), .B(P1_DATAO_REG_9__SCAN_IN), .S(n9105), .Z(
        P1_U3564) );
  MUX2_X1 U10468 ( .A(n9099), .B(P1_DATAO_REG_8__SCAN_IN), .S(n9105), .Z(
        P1_U3563) );
  MUX2_X1 U10469 ( .A(n9100), .B(P1_DATAO_REG_7__SCAN_IN), .S(n9105), .Z(
        P1_U3562) );
  MUX2_X1 U10470 ( .A(n9101), .B(P1_DATAO_REG_6__SCAN_IN), .S(n9105), .Z(
        P1_U3561) );
  MUX2_X1 U10471 ( .A(n9102), .B(P1_DATAO_REG_5__SCAN_IN), .S(n9105), .Z(
        P1_U3560) );
  MUX2_X1 U10472 ( .A(n9103), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9105), .Z(
        P1_U3559) );
  MUX2_X1 U10473 ( .A(n6677), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9105), .Z(
        P1_U3558) );
  MUX2_X1 U10474 ( .A(n9104), .B(P1_DATAO_REG_2__SCAN_IN), .S(n9105), .Z(
        P1_U3557) );
  MUX2_X1 U10475 ( .A(n9106), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9105), .Z(
        P1_U3556) );
  OAI21_X1 U10476 ( .B1(n9109), .B2(n9108), .A(n9107), .ZN(n9110) );
  NAND2_X1 U10477 ( .A1(n9110), .A2(n9824), .ZN(n9119) );
  AOI211_X1 U10478 ( .C1(n9113), .C2(n9112), .A(n9111), .B(n9819), .ZN(n9114)
         );
  AOI21_X1 U10479 ( .B1(n9815), .B2(n9115), .A(n9114), .ZN(n9118) );
  AOI21_X1 U10480 ( .B1(n9778), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n9116), .ZN(
        n9117) );
  NAND3_X1 U10481 ( .A1(n9119), .A2(n9118), .A3(n9117), .ZN(P1_U3253) );
  OAI21_X1 U10482 ( .B1(n9122), .B2(n9121), .A(n9120), .ZN(n9123) );
  NAND2_X1 U10483 ( .A1(n9123), .A2(n9824), .ZN(n9132) );
  AOI211_X1 U10484 ( .C1(n9126), .C2(n9125), .A(n9124), .B(n9819), .ZN(n9127)
         );
  AOI21_X1 U10485 ( .B1(n9815), .B2(n9128), .A(n9127), .ZN(n9130) );
  NAND2_X1 U10486 ( .A1(n9778), .A2(P1_ADDR_REG_13__SCAN_IN), .ZN(n9129) );
  NAND4_X1 U10487 ( .A1(n9132), .A2(n9131), .A3(n9130), .A4(n9129), .ZN(
        P1_U3254) );
  NOR2_X1 U10488 ( .A1(n9133), .A2(n9141), .ZN(n9135) );
  NOR2_X1 U10489 ( .A1(n9135), .A2(n9134), .ZN(n9139) );
  NOR2_X1 U10490 ( .A1(n9160), .A2(n9136), .ZN(n9137) );
  AOI21_X1 U10491 ( .B1(n9160), .B2(n9136), .A(n9137), .ZN(n9138) );
  NOR2_X1 U10492 ( .A1(n9139), .A2(n9138), .ZN(n9159) );
  AOI211_X1 U10493 ( .C1(n9139), .C2(n9138), .A(n9159), .B(n9819), .ZN(n9152)
         );
  NOR2_X1 U10494 ( .A1(n9141), .A2(n9140), .ZN(n9143) );
  NOR2_X1 U10495 ( .A1(n9143), .A2(n9142), .ZN(n9145) );
  XNOR2_X1 U10496 ( .A(n9160), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n9144) );
  NOR2_X1 U10497 ( .A1(n9145), .A2(n9144), .ZN(n9154) );
  AOI211_X1 U10498 ( .C1(n9145), .C2(n9144), .A(n9154), .B(n9769), .ZN(n9151)
         );
  NAND2_X1 U10499 ( .A1(P1_REG3_REG_16__SCAN_IN), .A2(P1_U3084), .ZN(n9147) );
  NAND2_X1 U10500 ( .A1(n9778), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n9146) );
  OAI211_X1 U10501 ( .C1(n9149), .C2(n9148), .A(n9147), .B(n9146), .ZN(n9150)
         );
  OR3_X1 U10502 ( .A1(n9152), .A2(n9151), .A3(n9150), .ZN(P1_U3257) );
  INV_X1 U10503 ( .A(n9153), .ZN(n9158) );
  AOI21_X1 U10504 ( .B1(n9160), .B2(P1_REG1_REG_16__SCAN_IN), .A(n9154), .ZN(
        n9156) );
  XNOR2_X1 U10505 ( .A(n9175), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n9155) );
  NOR2_X1 U10506 ( .A1(n9156), .A2(n9155), .ZN(n9174) );
  AOI211_X1 U10507 ( .C1(n9156), .C2(n9155), .A(n9174), .B(n9769), .ZN(n9157)
         );
  AOI211_X1 U10508 ( .C1(n9778), .C2(P1_ADDR_REG_17__SCAN_IN), .A(n9158), .B(
        n9157), .ZN(n9166) );
  NAND2_X1 U10509 ( .A1(n9175), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9161) );
  OAI21_X1 U10510 ( .B1(n9175), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9161), .ZN(
        n9162) );
  AOI211_X1 U10511 ( .C1(n9163), .C2(n9162), .A(n9167), .B(n9819), .ZN(n9164)
         );
  AOI21_X1 U10512 ( .B1(n9815), .B2(n9175), .A(n9164), .ZN(n9165) );
  NAND2_X1 U10513 ( .A1(n9166), .A2(n9165), .ZN(P1_U3258) );
  OR2_X1 U10514 ( .A1(n9814), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9169) );
  NAND2_X1 U10515 ( .A1(n9814), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9168) );
  NAND2_X1 U10516 ( .A1(n9169), .A2(n9168), .ZN(n9810) );
  AOI21_X1 U10517 ( .B1(n9814), .B2(P1_REG2_REG_18__SCAN_IN), .A(n9811), .ZN(
        n9170) );
  XNOR2_X1 U10518 ( .A(n9170), .B(n6143), .ZN(n9180) );
  NAND2_X1 U10519 ( .A1(n9180), .A2(n9171), .ZN(n9178) );
  AOI22_X1 U10520 ( .A1(n9814), .A2(P1_REG1_REG_18__SCAN_IN), .B1(n9173), .B2(
        n9172), .ZN(n9822) );
  AOI21_X1 U10521 ( .B1(P1_REG1_REG_17__SCAN_IN), .B2(n9175), .A(n9174), .ZN(
        n9823) );
  NAND2_X1 U10522 ( .A1(n9822), .A2(n9823), .ZN(n9821) );
  OAI21_X1 U10523 ( .B1(n9814), .B2(P1_REG1_REG_18__SCAN_IN), .A(n9821), .ZN(
        n9176) );
  XOR2_X1 U10524 ( .A(n9176), .B(P1_REG1_REG_19__SCAN_IN), .Z(n9179) );
  AOI21_X1 U10525 ( .B1(n9179), .B2(n9824), .A(n9815), .ZN(n9177) );
  NAND2_X1 U10526 ( .A1(n9178), .A2(n9177), .ZN(n9182) );
  OAI22_X1 U10527 ( .A1(n9180), .A2(n9819), .B1(n9179), .B2(n9769), .ZN(n9181)
         );
  MUX2_X1 U10528 ( .A(n9182), .B(n9181), .S(n9321), .Z(n9186) );
  OAI21_X1 U10529 ( .B1(n9828), .B2(n9184), .A(n9183), .ZN(n9185) );
  NAND2_X1 U10530 ( .A1(n9429), .A2(n9406), .ZN(n9403) );
  XNOR2_X1 U10531 ( .A(n9499), .B(n9498), .ZN(n9496) );
  NAND2_X1 U10532 ( .A1(n9496), .A2(n9493), .ZN(n9192) );
  INV_X1 U10533 ( .A(n9425), .ZN(n9447) );
  AND2_X1 U10534 ( .A1(n9188), .A2(P1_B_REG_SCAN_IN), .ZN(n9189) );
  NOR2_X1 U10535 ( .A1(n9422), .A2(n9189), .ZN(n9247) );
  NAND2_X1 U10536 ( .A1(n9247), .A2(n9190), .ZN(n9501) );
  NOR2_X1 U10537 ( .A1(n9447), .A2(n9501), .ZN(n9195) );
  AOI21_X1 U10538 ( .B1(n9490), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9195), .ZN(
        n9191) );
  OAI211_X1 U10539 ( .C1(n9498), .C2(n9480), .A(n9192), .B(n9191), .ZN(
        P1_U3261) );
  INV_X1 U10540 ( .A(n9219), .ZN(n9194) );
  NAND2_X1 U10541 ( .A1(n9194), .A2(n9193), .ZN(n9500) );
  NAND3_X1 U10542 ( .A1(n9500), .A2(n9499), .A3(n9493), .ZN(n9197) );
  AOI21_X1 U10543 ( .B1(n9490), .B2(P1_REG2_REG_30__SCAN_IN), .A(n9195), .ZN(
        n9196) );
  OAI211_X1 U10544 ( .C1(n9503), .C2(n9480), .A(n9197), .B(n9196), .ZN(
        P1_U3262) );
  NAND2_X1 U10545 ( .A1(n9392), .A2(n9421), .ZN(n9206) );
  NAND2_X1 U10546 ( .A1(n9551), .A2(n9396), .ZN(n9208) );
  AOI22_X1 U10547 ( .A1(n9372), .A2(n9208), .B1(n9207), .B2(n9374), .ZN(n9364)
         );
  NAND2_X1 U10548 ( .A1(n9333), .A2(n9212), .ZN(n9213) );
  INV_X1 U10549 ( .A(n9504), .ZN(n9252) );
  AOI211_X1 U10550 ( .C1(n9507), .C2(n9262), .A(n9883), .B(n9219), .ZN(n9506)
         );
  NOR2_X1 U10551 ( .A1(n4667), .A2(n9480), .ZN(n9222) );
  OAI22_X1 U10552 ( .A1(n9220), .A2(n9407), .B1(n9425), .B2(n8473), .ZN(n9221)
         );
  AOI211_X1 U10553 ( .C1(n9506), .C2(n9412), .A(n9222), .B(n9221), .ZN(n9251)
         );
  NAND2_X1 U10554 ( .A1(n9315), .A2(n9314), .ZN(n9313) );
  INV_X1 U10555 ( .A(n9238), .ZN(n9239) );
  NAND3_X1 U10556 ( .A1(n9258), .A2(n9256), .A3(n9257), .ZN(n9255) );
  NAND2_X1 U10557 ( .A1(n9255), .A2(n9243), .ZN(n9245) );
  XNOR2_X1 U10558 ( .A(n9245), .B(n9244), .ZN(n9249) );
  AOI22_X1 U10559 ( .A1(n9279), .A2(n9486), .B1(n9247), .B2(n9246), .ZN(n9248)
         );
  OAI21_X1 U10560 ( .B1(n9249), .B2(n9420), .A(n9248), .ZN(n9505) );
  NAND2_X1 U10561 ( .A1(n9505), .A2(n9425), .ZN(n9250) );
  OAI211_X1 U10562 ( .C1(n9252), .C2(n9495), .A(n9251), .B(n9250), .ZN(
        P1_U3355) );
  INV_X1 U10563 ( .A(n9255), .ZN(n9260) );
  AOI21_X1 U10564 ( .B1(n9258), .B2(n9257), .A(n9256), .ZN(n9259) );
  INV_X1 U10565 ( .A(n9262), .ZN(n9263) );
  AOI211_X1 U10566 ( .C1(n9512), .C2(n9271), .A(n9883), .B(n9263), .ZN(n9511)
         );
  NAND2_X1 U10567 ( .A1(n9511), .A2(n9412), .ZN(n9266) );
  AOI22_X1 U10568 ( .A1(n9264), .A2(n9477), .B1(P1_REG2_REG_28__SCAN_IN), .B2(
        n9490), .ZN(n9265) );
  OAI211_X1 U10569 ( .C1(n4666), .C2(n9480), .A(n9266), .B(n9265), .ZN(n9267)
         );
  AOI21_X1 U10570 ( .B1(n9510), .B2(n9425), .A(n9267), .ZN(n9268) );
  OAI21_X1 U10571 ( .B1(n9513), .B2(n9495), .A(n9268), .ZN(P1_U3263) );
  XNOR2_X1 U10572 ( .A(n9270), .B(n9269), .ZN(n9518) );
  INV_X1 U10573 ( .A(n9290), .ZN(n9273) );
  INV_X1 U10574 ( .A(n9271), .ZN(n9272) );
  AOI21_X1 U10575 ( .B1(n9514), .B2(n9273), .A(n9272), .ZN(n9515) );
  AOI22_X1 U10576 ( .A1(n9274), .A2(n9477), .B1(n9447), .B2(
        P1_REG2_REG_27__SCAN_IN), .ZN(n9275) );
  OAI21_X1 U10577 ( .B1(n9276), .B2(n9480), .A(n9275), .ZN(n9282) );
  XNOR2_X1 U10578 ( .A(n9278), .B(n9277), .ZN(n9280) );
  AOI222_X1 U10579 ( .A1(n9489), .A2(n9280), .B1(n9306), .B2(n9486), .C1(n9279), .C2(n9484), .ZN(n9517) );
  NOR2_X1 U10580 ( .A1(n9517), .A2(n9490), .ZN(n9281) );
  AOI211_X1 U10581 ( .C1(n9515), .C2(n9493), .A(n9282), .B(n9281), .ZN(n9283)
         );
  OAI21_X1 U10582 ( .B1(n9518), .B2(n9495), .A(n9283), .ZN(P1_U3264) );
  XNOR2_X1 U10583 ( .A(n9284), .B(n9285), .ZN(n9523) );
  XNOR2_X1 U10584 ( .A(n9286), .B(n9285), .ZN(n9287) );
  OAI222_X1 U10585 ( .A1(n9422), .A2(n9289), .B1(n9424), .B2(n9288), .C1(n9287), .C2(n9420), .ZN(n9519) );
  INV_X1 U10586 ( .A(n9299), .ZN(n9291) );
  AOI211_X1 U10587 ( .C1(n9521), .C2(n9291), .A(n9883), .B(n9290), .ZN(n9520)
         );
  NAND2_X1 U10588 ( .A1(n9520), .A2(n9412), .ZN(n9294) );
  AOI22_X1 U10589 ( .A1(P1_REG2_REG_26__SCAN_IN), .A2(n9447), .B1(n9292), .B2(
        n9477), .ZN(n9293) );
  OAI211_X1 U10590 ( .C1(n9295), .C2(n9480), .A(n9294), .B(n9293), .ZN(n9296)
         );
  AOI21_X1 U10591 ( .B1(n9519), .B2(n9425), .A(n9296), .ZN(n9297) );
  OAI21_X1 U10592 ( .B1(n9523), .B2(n9495), .A(n9297), .ZN(P1_U3265) );
  XOR2_X1 U10593 ( .A(n9298), .B(n9305), .Z(n9528) );
  AOI21_X1 U10594 ( .B1(n9524), .B2(n9318), .A(n9299), .ZN(n9525) );
  AOI22_X1 U10595 ( .A1(n9447), .A2(P1_REG2_REG_25__SCAN_IN), .B1(n9300), .B2(
        n9477), .ZN(n9301) );
  OAI21_X1 U10596 ( .B1(n9302), .B2(n9480), .A(n9301), .ZN(n9309) );
  NAND2_X1 U10597 ( .A1(n9313), .A2(n9303), .ZN(n9304) );
  XOR2_X1 U10598 ( .A(n9305), .B(n9304), .Z(n9307) );
  AOI222_X1 U10599 ( .A1(n9489), .A2(n9307), .B1(n9306), .B2(n9484), .C1(n9336), .C2(n9486), .ZN(n9527) );
  NOR2_X1 U10600 ( .A1(n9527), .A2(n9490), .ZN(n9308) );
  AOI211_X1 U10601 ( .C1(n9493), .C2(n9525), .A(n9309), .B(n9308), .ZN(n9310)
         );
  OAI21_X1 U10602 ( .B1(n9528), .B2(n9495), .A(n9310), .ZN(P1_U3266) );
  XNOR2_X1 U10603 ( .A(n9311), .B(n9314), .ZN(n9533) );
  NOR2_X1 U10604 ( .A1(n9312), .A2(n9480), .ZN(n9324) );
  OAI21_X1 U10605 ( .B1(n9315), .B2(n9314), .A(n9313), .ZN(n9317) );
  AOI222_X1 U10606 ( .A1(n9489), .A2(n9317), .B1(n9316), .B2(n9484), .C1(n9349), .C2(n9486), .ZN(n9532) );
  INV_X1 U10607 ( .A(n9318), .ZN(n9319) );
  AOI211_X1 U10608 ( .C1(n9530), .C2(n9327), .A(n9883), .B(n9319), .ZN(n9529)
         );
  AOI22_X1 U10609 ( .A1(n9529), .A2(n9321), .B1(n9477), .B2(n9320), .ZN(n9322)
         );
  AOI21_X1 U10610 ( .B1(n9532), .B2(n9322), .A(n9447), .ZN(n9323) );
  AOI211_X1 U10611 ( .C1(n9490), .C2(P1_REG2_REG_24__SCAN_IN), .A(n9324), .B(
        n9323), .ZN(n9325) );
  OAI21_X1 U10612 ( .B1(n9533), .B2(n9495), .A(n9325), .ZN(P1_U3267) );
  XNOR2_X1 U10613 ( .A(n9326), .B(n9334), .ZN(n9538) );
  INV_X1 U10614 ( .A(n9342), .ZN(n9329) );
  INV_X1 U10615 ( .A(n9327), .ZN(n9328) );
  AOI21_X1 U10616 ( .B1(n9534), .B2(n9329), .A(n9328), .ZN(n9535) );
  INV_X1 U10617 ( .A(n9330), .ZN(n9331) );
  AOI22_X1 U10618 ( .A1(n9447), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n9331), .B2(
        n9477), .ZN(n9332) );
  OAI21_X1 U10619 ( .B1(n9333), .B2(n9480), .A(n9332), .ZN(n9339) );
  XNOR2_X1 U10620 ( .A(n9335), .B(n9334), .ZN(n9337) );
  AOI222_X1 U10621 ( .A1(n9489), .A2(n9337), .B1(n9358), .B2(n9486), .C1(n9336), .C2(n9484), .ZN(n9537) );
  NOR2_X1 U10622 ( .A1(n9537), .A2(n9447), .ZN(n9338) );
  AOI211_X1 U10623 ( .C1(n9535), .C2(n9493), .A(n9339), .B(n9338), .ZN(n9340)
         );
  OAI21_X1 U10624 ( .B1(n9538), .B2(n9495), .A(n9340), .ZN(P1_U3268) );
  XOR2_X1 U10625 ( .A(n9341), .B(n9347), .Z(n9543) );
  AOI21_X1 U10626 ( .B1(n9539), .B2(n4453), .A(n9342), .ZN(n9540) );
  INV_X1 U10627 ( .A(n9343), .ZN(n9344) );
  AOI22_X1 U10628 ( .A1(n9447), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n9344), .B2(
        n9477), .ZN(n9345) );
  OAI21_X1 U10629 ( .B1(n9346), .B2(n9480), .A(n9345), .ZN(n9353) );
  XNOR2_X1 U10630 ( .A(n9348), .B(n9347), .ZN(n9351) );
  AOI222_X1 U10631 ( .A1(n9489), .A2(n9351), .B1(n9350), .B2(n9486), .C1(n9349), .C2(n9484), .ZN(n9542) );
  NOR2_X1 U10632 ( .A1(n9542), .A2(n9447), .ZN(n9352) );
  AOI211_X1 U10633 ( .C1(n9540), .C2(n9493), .A(n9353), .B(n9352), .ZN(n9354)
         );
  OAI21_X1 U10634 ( .B1(n9543), .B2(n9495), .A(n9354), .ZN(P1_U3269) );
  OAI211_X1 U10635 ( .C1(n9355), .C2(n9373), .A(n4453), .B(n9590), .ZN(n9545)
         );
  NOR2_X1 U10636 ( .A1(n9545), .A2(n9356), .ZN(n9361) );
  XNOR2_X1 U10637 ( .A(n9357), .B(n9363), .ZN(n9359) );
  AOI222_X1 U10638 ( .A1(n9489), .A2(n9359), .B1(n9358), .B2(n9484), .C1(n9396), .C2(n9486), .ZN(n9547) );
  INV_X1 U10639 ( .A(n9547), .ZN(n9360) );
  AOI211_X1 U10640 ( .C1(n9477), .C2(n9362), .A(n9361), .B(n9360), .ZN(n9371)
         );
  OR2_X1 U10641 ( .A1(n9364), .A2(n9363), .ZN(n9544) );
  NAND3_X1 U10642 ( .A1(n9544), .A2(n9365), .A3(n9366), .ZN(n9370) );
  AOI22_X1 U10643 ( .A1(n9368), .A2(n9367), .B1(n9447), .B2(
        P1_REG2_REG_21__SCAN_IN), .ZN(n9369) );
  OAI211_X1 U10644 ( .C1(n9490), .C2(n9371), .A(n9370), .B(n9369), .ZN(
        P1_U3270) );
  XNOR2_X1 U10645 ( .A(n9372), .B(n9380), .ZN(n9553) );
  AOI211_X1 U10646 ( .C1(n9551), .C2(n9387), .A(n9883), .B(n9373), .ZN(n9550)
         );
  NOR2_X1 U10647 ( .A1(n9374), .A2(n9480), .ZN(n9378) );
  OAI22_X1 U10648 ( .A1(n9425), .A2(n9376), .B1(n9375), .B2(n9407), .ZN(n9377)
         );
  AOI211_X1 U10649 ( .C1(n9550), .C2(n9412), .A(n9378), .B(n9377), .ZN(n9384)
         );
  XOR2_X1 U10650 ( .A(n9380), .B(n9379), .Z(n9381) );
  OAI222_X1 U10651 ( .A1(n9424), .A2(n9421), .B1(n9422), .B2(n9382), .C1(n9381), .C2(n9420), .ZN(n9549) );
  NAND2_X1 U10652 ( .A1(n9549), .A2(n9425), .ZN(n9383) );
  OAI211_X1 U10653 ( .C1(n9553), .C2(n9495), .A(n9384), .B(n9383), .ZN(
        P1_U3271) );
  XNOR2_X1 U10654 ( .A(n9386), .B(n9385), .ZN(n9558) );
  AOI21_X1 U10655 ( .B1(n9554), .B2(n9403), .A(n9388), .ZN(n9555) );
  INV_X1 U10656 ( .A(n9389), .ZN(n9390) );
  AOI22_X1 U10657 ( .A1(n9447), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9390), .B2(
        n9477), .ZN(n9391) );
  OAI21_X1 U10658 ( .B1(n9392), .B2(n9480), .A(n9391), .ZN(n9399) );
  OAI21_X1 U10659 ( .B1(n9395), .B2(n9394), .A(n9393), .ZN(n9397) );
  AOI222_X1 U10660 ( .A1(n9489), .A2(n9397), .B1(n9436), .B2(n9486), .C1(n9396), .C2(n9484), .ZN(n9557) );
  NOR2_X1 U10661 ( .A1(n9557), .A2(n9447), .ZN(n9398) );
  AOI211_X1 U10662 ( .C1(n9555), .C2(n9493), .A(n9399), .B(n9398), .ZN(n9400)
         );
  OAI21_X1 U10663 ( .B1(n9558), .B2(n9495), .A(n9400), .ZN(P1_U3272) );
  OAI21_X1 U10664 ( .B1(n9402), .B2(n9418), .A(n9401), .ZN(n9563) );
  INV_X1 U10665 ( .A(n9429), .ZN(n9405) );
  INV_X1 U10666 ( .A(n9403), .ZN(n9404) );
  AOI211_X1 U10667 ( .C1(n9561), .C2(n9405), .A(n9883), .B(n9404), .ZN(n9560)
         );
  NOR2_X1 U10668 ( .A1(n9406), .A2(n9480), .ZN(n9411) );
  OAI22_X1 U10669 ( .A1(n9425), .A2(n9409), .B1(n9408), .B2(n9407), .ZN(n9410)
         );
  AOI211_X1 U10670 ( .C1(n9560), .C2(n9412), .A(n9411), .B(n9410), .ZN(n9427)
         );
  NAND2_X1 U10671 ( .A1(n9449), .A2(n9413), .ZN(n9435) );
  INV_X1 U10672 ( .A(n9414), .ZN(n9416) );
  OAI21_X1 U10673 ( .B1(n9435), .B2(n9416), .A(n9415), .ZN(n9417) );
  XOR2_X1 U10674 ( .A(n9418), .B(n9417), .Z(n9419) );
  OAI222_X1 U10675 ( .A1(n9424), .A2(n9423), .B1(n9422), .B2(n9421), .C1(n9420), .C2(n9419), .ZN(n9559) );
  NAND2_X1 U10676 ( .A1(n9559), .A2(n9425), .ZN(n9426) );
  OAI211_X1 U10677 ( .C1(n9563), .C2(n9495), .A(n9427), .B(n9426), .ZN(
        P1_U3273) );
  XNOR2_X1 U10678 ( .A(n9428), .B(n9434), .ZN(n9568) );
  AOI21_X1 U10679 ( .B1(n9564), .B2(n9444), .A(n9429), .ZN(n9565) );
  INV_X1 U10680 ( .A(n9430), .ZN(n9431) );
  AOI22_X1 U10681 ( .A1(n9447), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9431), .B2(
        n9477), .ZN(n9432) );
  OAI21_X1 U10682 ( .B1(n9433), .B2(n9480), .A(n9432), .ZN(n9439) );
  XNOR2_X1 U10683 ( .A(n9435), .B(n9434), .ZN(n9437) );
  AOI222_X1 U10684 ( .A1(n9489), .A2(n9437), .B1(n9467), .B2(n9486), .C1(n9436), .C2(n9484), .ZN(n9567) );
  NOR2_X1 U10685 ( .A1(n9567), .A2(n9447), .ZN(n9438) );
  AOI211_X1 U10686 ( .C1(n9565), .C2(n9493), .A(n9439), .B(n9438), .ZN(n9440)
         );
  OAI21_X1 U10687 ( .B1(n9495), .B2(n9568), .A(n9440), .ZN(P1_U3274) );
  XNOR2_X1 U10688 ( .A(n9442), .B(n9441), .ZN(n9573) );
  INV_X1 U10689 ( .A(n9444), .ZN(n9445) );
  AOI211_X1 U10690 ( .C1(n9570), .C2(n4658), .A(n9883), .B(n9445), .ZN(n9569)
         );
  AOI22_X1 U10691 ( .A1(n9447), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9446), .B2(
        n9477), .ZN(n9448) );
  OAI21_X1 U10692 ( .B1(n9187), .B2(n9480), .A(n9448), .ZN(n9456) );
  OAI21_X1 U10693 ( .B1(n9451), .B2(n9450), .A(n9449), .ZN(n9454) );
  AOI222_X1 U10694 ( .A1(n9489), .A2(n9454), .B1(n9453), .B2(n9484), .C1(n9452), .C2(n9486), .ZN(n9572) );
  NOR2_X1 U10695 ( .A1(n9572), .A2(n9490), .ZN(n9455) );
  AOI211_X1 U10696 ( .C1(n9569), .C2(n9457), .A(n9456), .B(n9455), .ZN(n9458)
         );
  OAI21_X1 U10697 ( .B1(n9495), .B2(n9573), .A(n9458), .ZN(P1_U3275) );
  XOR2_X1 U10698 ( .A(n9459), .B(n9466), .Z(n9578) );
  AOI21_X1 U10699 ( .B1(n9574), .B2(n9460), .A(n9443), .ZN(n9575) );
  INV_X1 U10700 ( .A(n9461), .ZN(n9462) );
  AOI22_X1 U10701 ( .A1(n9447), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n9462), .B2(
        n9477), .ZN(n9463) );
  OAI21_X1 U10702 ( .B1(n9464), .B2(n9480), .A(n9463), .ZN(n9470) );
  XOR2_X1 U10703 ( .A(n9466), .B(n9465), .Z(n9468) );
  AOI222_X1 U10704 ( .A1(n9489), .A2(n9468), .B1(n9467), .B2(n9484), .C1(n9485), .C2(n9486), .ZN(n9577) );
  NOR2_X1 U10705 ( .A1(n9577), .A2(n9490), .ZN(n9469) );
  AOI211_X1 U10706 ( .C1(n9575), .C2(n9493), .A(n9470), .B(n9469), .ZN(n9471)
         );
  OAI21_X1 U10707 ( .B1(n9495), .B2(n9578), .A(n9471), .ZN(P1_U3276) );
  XNOR2_X1 U10708 ( .A(n9472), .B(n9482), .ZN(n9583) );
  INV_X1 U10709 ( .A(n9473), .ZN(n9475) );
  AOI21_X1 U10710 ( .B1(n9579), .B2(n9475), .A(n9474), .ZN(n9580) );
  INV_X1 U10711 ( .A(n9476), .ZN(n9478) );
  AOI22_X1 U10712 ( .A1(n9447), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n9478), .B2(
        n9477), .ZN(n9479) );
  OAI21_X1 U10713 ( .B1(n9481), .B2(n9480), .A(n9479), .ZN(n9492) );
  XNOR2_X1 U10714 ( .A(n9483), .B(n9482), .ZN(n9488) );
  AOI222_X1 U10715 ( .A1(n9489), .A2(n9488), .B1(n9487), .B2(n9486), .C1(n9485), .C2(n9484), .ZN(n9582) );
  NOR2_X1 U10716 ( .A1(n9582), .A2(n9490), .ZN(n9491) );
  AOI211_X1 U10717 ( .C1(n9580), .C2(n9493), .A(n9492), .B(n9491), .ZN(n9494)
         );
  OAI21_X1 U10718 ( .B1(n9583), .B2(n9495), .A(n9494), .ZN(P1_U3278) );
  NAND2_X1 U10719 ( .A1(n9496), .A2(n9590), .ZN(n9497) );
  OAI211_X1 U10720 ( .C1(n9498), .C2(n9881), .A(n9497), .B(n9501), .ZN(n9596)
         );
  MUX2_X1 U10721 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9596), .S(n9910), .Z(
        P1_U3554) );
  NAND3_X1 U10722 ( .A1(n9500), .A2(n9499), .A3(n9590), .ZN(n9502) );
  OAI211_X1 U10723 ( .C1(n9503), .C2(n9881), .A(n9502), .B(n9501), .ZN(n9597)
         );
  MUX2_X1 U10724 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n9597), .S(n9910), .Z(
        P1_U3553) );
  NAND2_X1 U10725 ( .A1(n9504), .A2(n9887), .ZN(n9509) );
  NAND2_X1 U10726 ( .A1(n9509), .A2(n9508), .ZN(n9598) );
  MUX2_X1 U10727 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9598), .S(n9910), .Z(
        P1_U3552) );
  AOI22_X1 U10728 ( .A1(n9515), .A2(n9590), .B1(n9892), .B2(n9514), .ZN(n9516)
         );
  OAI211_X1 U10729 ( .C1(n9518), .C2(n9894), .A(n9517), .B(n9516), .ZN(n9600)
         );
  MUX2_X1 U10730 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9600), .S(n9910), .Z(
        P1_U3550) );
  AOI211_X1 U10731 ( .C1(n9892), .C2(n9521), .A(n9520), .B(n9519), .ZN(n9522)
         );
  OAI21_X1 U10732 ( .B1(n9523), .B2(n9894), .A(n9522), .ZN(n9601) );
  MUX2_X1 U10733 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9601), .S(n9910), .Z(
        P1_U3549) );
  AOI22_X1 U10734 ( .A1(n9525), .A2(n9590), .B1(n9892), .B2(n9524), .ZN(n9526)
         );
  OAI211_X1 U10735 ( .C1(n9528), .C2(n9894), .A(n9527), .B(n9526), .ZN(n9602)
         );
  MUX2_X1 U10736 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9602), .S(n9910), .Z(
        P1_U3548) );
  AOI21_X1 U10737 ( .B1(n9892), .B2(n9530), .A(n9529), .ZN(n9531) );
  OAI211_X1 U10738 ( .C1(n9533), .C2(n9894), .A(n9532), .B(n9531), .ZN(n9603)
         );
  MUX2_X1 U10739 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9603), .S(n9910), .Z(
        P1_U3547) );
  AOI22_X1 U10740 ( .A1(n9535), .A2(n9590), .B1(n9892), .B2(n9534), .ZN(n9536)
         );
  OAI211_X1 U10741 ( .C1(n9538), .C2(n9894), .A(n9537), .B(n9536), .ZN(n9604)
         );
  MUX2_X1 U10742 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9604), .S(n9910), .Z(
        P1_U3546) );
  AOI22_X1 U10743 ( .A1(n9540), .A2(n9590), .B1(n9892), .B2(n9539), .ZN(n9541)
         );
  OAI211_X1 U10744 ( .C1(n9543), .C2(n9894), .A(n9542), .B(n9541), .ZN(n9605)
         );
  MUX2_X1 U10745 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9605), .S(n9910), .Z(
        P1_U3545) );
  NAND3_X1 U10746 ( .A1(n9544), .A2(n9365), .A3(n9887), .ZN(n9548) );
  NAND4_X1 U10747 ( .A1(n9548), .A2(n9547), .A3(n9546), .A4(n9545), .ZN(n9606)
         );
  MUX2_X1 U10748 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9606), .S(n9910), .Z(
        P1_U3544) );
  AOI211_X1 U10749 ( .C1(n9892), .C2(n9551), .A(n9550), .B(n9549), .ZN(n9552)
         );
  OAI21_X1 U10750 ( .B1(n9553), .B2(n9894), .A(n9552), .ZN(n9607) );
  MUX2_X1 U10751 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9607), .S(n9910), .Z(
        P1_U3543) );
  AOI22_X1 U10752 ( .A1(n9555), .A2(n9590), .B1(n9892), .B2(n9554), .ZN(n9556)
         );
  OAI211_X1 U10753 ( .C1(n9558), .C2(n9894), .A(n9557), .B(n9556), .ZN(n9608)
         );
  MUX2_X1 U10754 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9608), .S(n9910), .Z(
        P1_U3542) );
  AOI211_X1 U10755 ( .C1(n9892), .C2(n9561), .A(n9560), .B(n9559), .ZN(n9562)
         );
  OAI21_X1 U10756 ( .B1(n9563), .B2(n9894), .A(n9562), .ZN(n9609) );
  MUX2_X1 U10757 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9609), .S(n9910), .Z(
        P1_U3541) );
  AOI22_X1 U10758 ( .A1(n9565), .A2(n9590), .B1(n9892), .B2(n9564), .ZN(n9566)
         );
  OAI211_X1 U10759 ( .C1(n9568), .C2(n9894), .A(n9567), .B(n9566), .ZN(n9610)
         );
  MUX2_X1 U10760 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9610), .S(n9910), .Z(
        P1_U3540) );
  AOI21_X1 U10761 ( .B1(n9892), .B2(n9570), .A(n9569), .ZN(n9571) );
  OAI211_X1 U10762 ( .C1(n9573), .C2(n9894), .A(n9572), .B(n9571), .ZN(n9611)
         );
  MUX2_X1 U10763 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9611), .S(n9910), .Z(
        P1_U3539) );
  AOI22_X1 U10764 ( .A1(n9575), .A2(n9590), .B1(n9892), .B2(n9574), .ZN(n9576)
         );
  OAI211_X1 U10765 ( .C1(n9578), .C2(n9894), .A(n9577), .B(n9576), .ZN(n9612)
         );
  MUX2_X1 U10766 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n9612), .S(n9910), .Z(
        P1_U3538) );
  AOI22_X1 U10767 ( .A1(n9580), .A2(n9590), .B1(n9892), .B2(n9579), .ZN(n9581)
         );
  OAI211_X1 U10768 ( .C1(n9583), .C2(n9894), .A(n9582), .B(n9581), .ZN(n9613)
         );
  MUX2_X1 U10769 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n9613), .S(n9910), .Z(
        P1_U3536) );
  AOI211_X1 U10770 ( .C1(n9892), .C2(n9586), .A(n9585), .B(n9584), .ZN(n9587)
         );
  OAI21_X1 U10771 ( .B1(n9894), .B2(n9588), .A(n9587), .ZN(n9614) );
  MUX2_X1 U10772 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n9614), .S(n9910), .Z(
        P1_U3535) );
  AOI22_X1 U10773 ( .A1(n9591), .A2(n9590), .B1(n9892), .B2(n9589), .ZN(n9592)
         );
  OAI21_X1 U10774 ( .B1(n9593), .B2(n9843), .A(n9592), .ZN(n9594) );
  MUX2_X1 U10775 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n9615), .S(n9910), .Z(
        P1_U3534) );
  MUX2_X1 U10776 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9596), .S(n9900), .Z(
        P1_U3522) );
  MUX2_X1 U10777 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n9597), .S(n9900), .Z(
        P1_U3521) );
  MUX2_X1 U10778 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9598), .S(n9900), .Z(
        P1_U3520) );
  MUX2_X1 U10779 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9599), .S(n9900), .Z(
        P1_U3519) );
  MUX2_X1 U10780 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9600), .S(n9900), .Z(
        P1_U3518) );
  MUX2_X1 U10781 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9601), .S(n9900), .Z(
        P1_U3517) );
  MUX2_X1 U10782 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9602), .S(n9900), .Z(
        P1_U3516) );
  MUX2_X1 U10783 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9603), .S(n9900), .Z(
        P1_U3515) );
  MUX2_X1 U10784 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9604), .S(n9900), .Z(
        P1_U3514) );
  MUX2_X1 U10785 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9605), .S(n9900), .Z(
        P1_U3513) );
  MUX2_X1 U10786 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9606), .S(n9900), .Z(
        P1_U3512) );
  MUX2_X1 U10787 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9607), .S(n9900), .Z(
        P1_U3511) );
  MUX2_X1 U10788 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9608), .S(n9900), .Z(
        P1_U3510) );
  MUX2_X1 U10789 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9609), .S(n9900), .Z(
        P1_U3508) );
  MUX2_X1 U10790 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9610), .S(n9900), .Z(
        P1_U3505) );
  MUX2_X1 U10791 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9611), .S(n9900), .Z(
        P1_U3502) );
  MUX2_X1 U10792 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n9612), .S(n9900), .Z(
        P1_U3499) );
  MUX2_X1 U10793 ( .A(P1_REG0_REG_13__SCAN_IN), .B(n9613), .S(n9900), .Z(
        P1_U3493) );
  MUX2_X1 U10794 ( .A(P1_REG0_REG_12__SCAN_IN), .B(n9614), .S(n9900), .Z(
        P1_U3490) );
  MUX2_X1 U10795 ( .A(n9615), .B(P1_REG0_REG_11__SCAN_IN), .S(n9898), .Z(
        P1_U3487) );
  MUX2_X1 U10796 ( .A(P1_D_REG_0__SCAN_IN), .B(n9616), .S(n9841), .Z(P1_U3440)
         );
  NAND3_X1 U10797 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_STATE_REG_SCAN_IN), 
        .A3(n9617), .ZN(n9619) );
  OAI22_X1 U10798 ( .A1(n9620), .A2(n9619), .B1(n6435), .B2(n9618), .ZN(n9621)
         );
  AOI21_X1 U10799 ( .B1(n9623), .B2(n9622), .A(n9621), .ZN(n9624) );
  INV_X1 U10800 ( .A(n9624), .ZN(P1_U3322) );
  MUX2_X1 U10801 ( .A(n9625), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  OAI21_X1 U10802 ( .B1(n9627), .B2(n9626), .A(n4639), .ZN(n9639) );
  NAND2_X1 U10803 ( .A1(n9815), .A2(n9628), .ZN(n9638) );
  AND3_X1 U10804 ( .A1(n9631), .A2(n9630), .A3(n9629), .ZN(n9632) );
  OR3_X1 U10805 ( .A1(n9769), .A2(n9633), .A3(n9632), .ZN(n9636) );
  INV_X1 U10806 ( .A(n9634), .ZN(n9635) );
  AND2_X1 U10807 ( .A1(n9636), .A2(n9635), .ZN(n9637) );
  OAI211_X1 U10808 ( .C1(n9639), .C2(n9819), .A(n9638), .B(n9637), .ZN(n9640)
         );
  INV_X1 U10809 ( .A(n9640), .ZN(n9641) );
  OAI21_X1 U10810 ( .B1(n9642), .B2(n9828), .A(n9641), .ZN(P1_U3244) );
  AOI22_X1 U10811 ( .A1(n9969), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3152), .ZN(n9653) );
  AOI211_X1 U10812 ( .C1(n9645), .C2(n9644), .A(n9643), .B(n9972), .ZN(n9646)
         );
  AOI21_X1 U10813 ( .B1(n9659), .B2(n9647), .A(n9646), .ZN(n9652) );
  AND2_X1 U10814 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n9650) );
  OAI211_X1 U10815 ( .C1(n9650), .C2(n9649), .A(n9968), .B(n9648), .ZN(n9651)
         );
  NAND3_X1 U10816 ( .A1(n9653), .A2(n9652), .A3(n9651), .ZN(P2_U3246) );
  AOI22_X1 U10817 ( .A1(n9969), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n9665) );
  AOI211_X1 U10818 ( .C1(n9656), .C2(n9655), .A(n9654), .B(n9972), .ZN(n9657)
         );
  AOI21_X1 U10819 ( .B1(n9659), .B2(n9658), .A(n9657), .ZN(n9664) );
  OAI211_X1 U10820 ( .C1(n9662), .C2(n9661), .A(n9968), .B(n9660), .ZN(n9663)
         );
  NAND3_X1 U10821 ( .A1(n9665), .A2(n9664), .A3(n9663), .ZN(P2_U3247) );
  NOR2_X1 U10822 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n9666) );
  AOI21_X1 U10823 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n9666), .ZN(n10139) );
  NOR2_X1 U10824 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n9667) );
  AOI21_X1 U10825 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n9667), .ZN(n10142) );
  NOR2_X1 U10826 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n9668) );
  AOI21_X1 U10827 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n9668), .ZN(n10145) );
  NOR2_X1 U10828 ( .A1(P1_ADDR_REG_14__SCAN_IN), .A2(P2_ADDR_REG_14__SCAN_IN), 
        .ZN(n9669) );
  AOI21_X1 U10829 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n9669), .ZN(n10148) );
  NOR2_X1 U10830 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n9670) );
  AOI21_X1 U10831 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n9670), .ZN(n10151) );
  NOR2_X1 U10832 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n9671) );
  AOI21_X1 U10833 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(P1_ADDR_REG_4__SCAN_IN), 
        .A(n9671), .ZN(n10190) );
  INV_X1 U10834 ( .A(n9673), .ZN(n9674) );
  NAND2_X1 U10835 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n10135) );
  INV_X1 U10836 ( .A(n10135), .ZN(n9672) );
  NAND2_X1 U10837 ( .A1(n10135), .A2(n6608), .ZN(n10133) );
  AOI22_X1 U10838 ( .A1(n9672), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P2_ADDR_REG_1__SCAN_IN), .B2(n10133), .ZN(n10184) );
  OAI21_X1 U10839 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(P1_ADDR_REG_2__SCAN_IN), 
        .A(n9673), .ZN(n10183) );
  NOR2_X1 U10840 ( .A1(n10184), .A2(n10183), .ZN(n10182) );
  NOR2_X1 U10841 ( .A1(n9674), .A2(n10182), .ZN(n10187) );
  NAND2_X1 U10842 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n9675) );
  OAI21_X1 U10843 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(P2_ADDR_REG_3__SCAN_IN), 
        .A(n9675), .ZN(n10186) );
  NOR2_X1 U10844 ( .A1(n10187), .A2(n10186), .ZN(n10185) );
  AOI21_X1 U10845 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(P1_ADDR_REG_3__SCAN_IN), 
        .A(n10185), .ZN(n10189) );
  NAND2_X1 U10846 ( .A1(n10190), .A2(n10189), .ZN(n10188) );
  OAI21_X1 U10847 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(P2_ADDR_REG_4__SCAN_IN), 
        .A(n10188), .ZN(n9676) );
  INV_X1 U10848 ( .A(n9676), .ZN(n9677) );
  NOR2_X1 U10849 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n9677), .ZN(n10168) );
  INV_X1 U10850 ( .A(n10168), .ZN(n10169) );
  NAND2_X1 U10851 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n9677), .ZN(n10170) );
  NAND2_X1 U10852 ( .A1(n10171), .A2(n10170), .ZN(n10167) );
  NAND2_X1 U10853 ( .A1(n10169), .A2(n10167), .ZN(n9679) );
  NOR2_X1 U10854 ( .A1(n9679), .A2(n9678), .ZN(n9680) );
  XNOR2_X1 U10855 ( .A(n9679), .B(n9678), .ZN(n10166) );
  INV_X1 U10856 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n10165) );
  NOR2_X1 U10857 ( .A1(n9681), .A2(n9682), .ZN(n9683) );
  XNOR2_X1 U10858 ( .A(n9682), .B(n9681), .ZN(n10174) );
  INV_X1 U10859 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n10173) );
  INV_X1 U10860 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n9777) );
  NOR2_X1 U10861 ( .A1(n9684), .A2(n9777), .ZN(n9685) );
  XNOR2_X1 U10862 ( .A(n9777), .B(n9684), .ZN(n10163) );
  INV_X1 U10863 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n10162) );
  NOR2_X1 U10864 ( .A1(n9686), .A2(n9687), .ZN(n9688) );
  XNOR2_X1 U10865 ( .A(n9687), .B(n9686), .ZN(n10180) );
  NAND2_X1 U10866 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n9689) );
  OAI21_X1 U10867 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n9689), .ZN(n10159) );
  NAND2_X1 U10868 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n9690) );
  OAI21_X1 U10869 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n9690), .ZN(n10156) );
  NOR2_X1 U10870 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n9691) );
  AOI21_X1 U10871 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n9691), .ZN(n10153) );
  NAND2_X1 U10872 ( .A1(n10154), .A2(n10153), .ZN(n10152) );
  NAND2_X1 U10873 ( .A1(n10151), .A2(n10150), .ZN(n10149) );
  NAND2_X1 U10874 ( .A1(n10148), .A2(n10147), .ZN(n10146) );
  NAND2_X1 U10875 ( .A1(n10145), .A2(n10144), .ZN(n10143) );
  OAI21_X1 U10876 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10143), .ZN(n10141) );
  NAND2_X1 U10877 ( .A1(n10142), .A2(n10141), .ZN(n10140) );
  OAI21_X1 U10878 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10140), .ZN(n10138) );
  NAND2_X1 U10879 ( .A1(n10139), .A2(n10138), .ZN(n10137) );
  NOR2_X1 U10880 ( .A1(n10177), .A2(n10176), .ZN(n9692) );
  NAND2_X1 U10881 ( .A1(n10177), .A2(n10176), .ZN(n10175) );
  OAI21_X1 U10882 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n9692), .A(n10175), .ZN(
        n9694) );
  XOR2_X1 U10883 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .Z(n9693) );
  XNOR2_X1 U10884 ( .A(n9694), .B(n9693), .ZN(ADD_1071_U4) );
  OAI211_X1 U10885 ( .C1(n9697), .C2(n10110), .A(n9696), .B(n9695), .ZN(n9698)
         );
  AOI21_X1 U10886 ( .B1(n9699), .B2(n10114), .A(n9698), .ZN(n9711) );
  AOI22_X1 U10887 ( .A1(n10124), .A2(n9711), .B1(n5384), .B2(n10131), .ZN(
        P2_U3535) );
  OAI22_X1 U10888 ( .A1(n9701), .A2(n10102), .B1(n9700), .B2(n10110), .ZN(
        n9702) );
  AOI211_X1 U10889 ( .C1(n9704), .C2(n10114), .A(n9703), .B(n9702), .ZN(n9713)
         );
  AOI22_X1 U10890 ( .A1(n10124), .A2(n9713), .B1(n6867), .B2(n10131), .ZN(
        P2_U3534) );
  INV_X1 U10891 ( .A(n10080), .ZN(n10096) );
  INV_X1 U10892 ( .A(n9705), .ZN(n9710) );
  OAI22_X1 U10893 ( .A1(n9707), .A2(n10102), .B1(n4541), .B2(n10110), .ZN(
        n9709) );
  AOI211_X1 U10894 ( .C1(n10096), .C2(n9710), .A(n9709), .B(n9708), .ZN(n9715)
         );
  AOI22_X1 U10895 ( .A1(n10124), .A2(n9715), .B1(n5328), .B2(n10131), .ZN(
        P2_U3533) );
  AOI22_X1 U10896 ( .A1(n10117), .A2(n9711), .B1(n5388), .B2(n10115), .ZN(
        P2_U3496) );
  INV_X1 U10897 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n9712) );
  AOI22_X1 U10898 ( .A1(n10117), .A2(n9713), .B1(n9712), .B2(n10115), .ZN(
        P2_U3493) );
  INV_X1 U10899 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n9714) );
  AOI22_X1 U10900 ( .A1(n10117), .A2(n9715), .B1(n9714), .B2(n10115), .ZN(
        P2_U3490) );
  OAI21_X1 U10901 ( .B1(n4758), .B2(n9881), .A(n9716), .ZN(n9717) );
  AOI211_X1 U10902 ( .C1(n9719), .C2(n9887), .A(n9718), .B(n9717), .ZN(n9721)
         );
  AOI22_X1 U10903 ( .A1(n9910), .A2(n9721), .B1(n6046), .B2(n9908), .ZN(
        P1_U3537) );
  INV_X1 U10904 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n9720) );
  AOI22_X1 U10905 ( .A1(n9900), .A2(n9721), .B1(n9720), .B2(n9898), .ZN(
        P1_U3496) );
  XNOR2_X1 U10906 ( .A(P1_WR_REG_SCAN_IN), .B(P2_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U10907 ( .A(P2_RD_REG_SCAN_IN), .B(P1_RD_REG_SCAN_IN), .ZN(U126) );
  INV_X1 U10908 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n9729) );
  OAI22_X1 U10909 ( .A1(n9723), .A2(n9722), .B1(P1_IR_REG_0__SCAN_IN), .B2(
        n5826), .ZN(n9725) );
  OAI211_X1 U10910 ( .C1(n9726), .C2(n9725), .A(n9724), .B(n5838), .ZN(n9727)
         );
  OAI22_X1 U10911 ( .A1(n9828), .A2(n9729), .B1(n9728), .B2(n9727), .ZN(n9730)
         );
  INV_X1 U10912 ( .A(n9730), .ZN(n9732) );
  NAND3_X1 U10913 ( .A1(n9824), .A2(P1_IR_REG_0__SCAN_IN), .A3(n5826), .ZN(
        n9731) );
  OAI211_X1 U10914 ( .C1(P1_STATE_REG_SCAN_IN), .C2(n7027), .A(n9732), .B(
        n9731), .ZN(P1_U3241) );
  OAI21_X1 U10915 ( .B1(n4415), .B2(n9734), .A(n9733), .ZN(n9736) );
  AOI22_X1 U10916 ( .A1(n9765), .A2(n9736), .B1(n9815), .B2(n9735), .ZN(n9745)
         );
  AOI21_X1 U10917 ( .B1(n9739), .B2(n9738), .A(n9737), .ZN(n9740) );
  NOR2_X1 U10918 ( .A1(n9769), .A2(n9740), .ZN(n9741) );
  AOI211_X1 U10919 ( .C1(P1_ADDR_REG_4__SCAN_IN), .C2(n9778), .A(n9742), .B(
        n9741), .ZN(n9744) );
  NAND3_X1 U10920 ( .A1(n9745), .A2(n9744), .A3(n9743), .ZN(P1_U3245) );
  AOI22_X1 U10921 ( .A1(n9815), .A2(n9746), .B1(n9778), .B2(
        P1_ADDR_REG_5__SCAN_IN), .ZN(n9757) );
  INV_X1 U10922 ( .A(n9747), .ZN(n9756) );
  XNOR2_X1 U10923 ( .A(n9749), .B(n9748), .ZN(n9750) );
  NAND2_X1 U10924 ( .A1(n9765), .A2(n9750), .ZN(n9755) );
  OAI211_X1 U10925 ( .C1(n9753), .C2(n9752), .A(n9824), .B(n9751), .ZN(n9754)
         );
  NAND4_X1 U10926 ( .A1(n9757), .A2(n9756), .A3(n9755), .A4(n9754), .ZN(
        P1_U3246) );
  OAI21_X1 U10927 ( .B1(n9760), .B2(n9759), .A(n9758), .ZN(n9764) );
  AND3_X1 U10928 ( .A1(n9824), .A2(n9762), .A3(n9761), .ZN(n9763) );
  AOI21_X1 U10929 ( .B1(n9765), .B2(n9764), .A(n9763), .ZN(n9776) );
  INV_X1 U10930 ( .A(n9766), .ZN(n9771) );
  INV_X1 U10931 ( .A(n9767), .ZN(n9768) );
  AOI211_X1 U10932 ( .C1(n9771), .C2(n9770), .A(n9769), .B(n9768), .ZN(n9772)
         );
  AOI211_X1 U10933 ( .C1(n9815), .C2(n9774), .A(n9773), .B(n9772), .ZN(n9775)
         );
  OAI211_X1 U10934 ( .C1(n9828), .C2(n9777), .A(n9776), .B(n9775), .ZN(
        P1_U3249) );
  AOI22_X1 U10935 ( .A1(n9815), .A2(n9779), .B1(n9778), .B2(
        P1_ADDR_REG_10__SCAN_IN), .ZN(n9791) );
  OAI21_X1 U10936 ( .B1(n9782), .B2(n9781), .A(n9780), .ZN(n9789) );
  INV_X1 U10937 ( .A(n9783), .ZN(n9786) );
  AOI211_X1 U10938 ( .C1(n9786), .C2(n4649), .A(n9785), .B(n9819), .ZN(n9787)
         );
  AOI211_X1 U10939 ( .C1(n9824), .C2(n9789), .A(n9788), .B(n9787), .ZN(n9790)
         );
  NAND2_X1 U10940 ( .A1(n9791), .A2(n9790), .ZN(P1_U3251) );
  NAND2_X1 U10941 ( .A1(n9792), .A2(n7466), .ZN(n9795) );
  INV_X1 U10942 ( .A(n9793), .ZN(n9794) );
  NAND2_X1 U10943 ( .A1(n9795), .A2(n9794), .ZN(n9800) );
  NAND2_X1 U10944 ( .A1(n9815), .A2(n9796), .ZN(n9799) );
  INV_X1 U10945 ( .A(n9797), .ZN(n9798) );
  OAI211_X1 U10946 ( .C1(n9819), .C2(n9800), .A(n9799), .B(n9798), .ZN(n9801)
         );
  INV_X1 U10947 ( .A(n9801), .ZN(n9807) );
  OAI21_X1 U10948 ( .B1(n9804), .B2(n9803), .A(n9802), .ZN(n9805) );
  NAND2_X1 U10949 ( .A1(n9805), .A2(n9824), .ZN(n9806) );
  OAI211_X1 U10950 ( .C1(n9828), .C2(n9808), .A(n9807), .B(n9806), .ZN(
        P1_U3255) );
  NAND2_X1 U10951 ( .A1(n9810), .A2(n9809), .ZN(n9813) );
  INV_X1 U10952 ( .A(n9811), .ZN(n9812) );
  NAND2_X1 U10953 ( .A1(n9813), .A2(n9812), .ZN(n9818) );
  NAND2_X1 U10954 ( .A1(n9815), .A2(n9814), .ZN(n9817) );
  OAI211_X1 U10955 ( .C1(n9819), .C2(n9818), .A(n9817), .B(n9816), .ZN(n9820)
         );
  INV_X1 U10956 ( .A(n9820), .ZN(n9827) );
  OAI21_X1 U10957 ( .B1(n9823), .B2(n9822), .A(n9821), .ZN(n9825) );
  NAND2_X1 U10958 ( .A1(n9825), .A2(n9824), .ZN(n9826) );
  OAI211_X1 U10959 ( .C1(n9828), .C2(n10177), .A(n9827), .B(n9826), .ZN(
        P1_U3259) );
  AND2_X1 U10960 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9838), .ZN(P1_U3292) );
  AND2_X1 U10961 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9838), .ZN(P1_U3293) );
  AND2_X1 U10962 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9838), .ZN(P1_U3294) );
  AND2_X1 U10963 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9838), .ZN(P1_U3295) );
  NOR2_X1 U10964 ( .A1(n9837), .A2(n9830), .ZN(P1_U3296) );
  AND2_X1 U10965 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9838), .ZN(P1_U3297) );
  NOR2_X1 U10966 ( .A1(n9837), .A2(n9831), .ZN(P1_U3298) );
  NOR2_X1 U10967 ( .A1(n9837), .A2(n9832), .ZN(P1_U3299) );
  AND2_X1 U10968 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9838), .ZN(P1_U3300) );
  NOR2_X1 U10969 ( .A1(n9837), .A2(n9833), .ZN(P1_U3301) );
  AND2_X1 U10970 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9838), .ZN(P1_U3302) );
  AND2_X1 U10971 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9838), .ZN(P1_U3303) );
  NOR2_X1 U10972 ( .A1(n9837), .A2(n9834), .ZN(P1_U3304) );
  AND2_X1 U10973 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9838), .ZN(P1_U3305) );
  NOR2_X1 U10974 ( .A1(n9837), .A2(n9835), .ZN(P1_U3306) );
  AND2_X1 U10975 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9838), .ZN(P1_U3307) );
  AND2_X1 U10976 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9838), .ZN(P1_U3308) );
  AND2_X1 U10977 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9838), .ZN(P1_U3309) );
  AND2_X1 U10978 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9838), .ZN(P1_U3310) );
  AND2_X1 U10979 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9838), .ZN(P1_U3311) );
  AND2_X1 U10980 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9838), .ZN(P1_U3312) );
  AND2_X1 U10981 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9838), .ZN(P1_U3313) );
  NOR2_X1 U10982 ( .A1(n9837), .A2(n9836), .ZN(P1_U3314) );
  AND2_X1 U10983 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9838), .ZN(P1_U3315) );
  AND2_X1 U10984 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9838), .ZN(P1_U3316) );
  AND2_X1 U10985 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9838), .ZN(P1_U3317) );
  AND2_X1 U10986 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9838), .ZN(P1_U3318) );
  AND2_X1 U10987 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n9838), .ZN(P1_U3319) );
  AND2_X1 U10988 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9838), .ZN(P1_U3320) );
  AND2_X1 U10989 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9838), .ZN(P1_U3321) );
  INV_X1 U10990 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n9842) );
  NAND2_X1 U10991 ( .A1(n9839), .A2(n9841), .ZN(n9840) );
  OAI21_X1 U10992 ( .B1(n9842), .B2(n9841), .A(n9840), .ZN(P1_U3441) );
  INV_X1 U10993 ( .A(n9843), .ZN(n9860) );
  INV_X1 U10994 ( .A(n9844), .ZN(n9849) );
  OAI21_X1 U10995 ( .B1(n9881), .B2(n9846), .A(n9845), .ZN(n9848) );
  AOI211_X1 U10996 ( .C1(n9860), .C2(n9849), .A(n9848), .B(n9847), .ZN(n9901)
         );
  AOI22_X1 U10997 ( .A1(n9900), .A2(n9901), .B1(n5833), .B2(n9898), .ZN(
        P1_U3457) );
  OAI22_X1 U10998 ( .A1(n9851), .A2(n9883), .B1(n9850), .B2(n9881), .ZN(n9853)
         );
  AOI211_X1 U10999 ( .C1(n9887), .C2(n9854), .A(n9853), .B(n9852), .ZN(n9902)
         );
  AOI22_X1 U11000 ( .A1(n9900), .A2(n9902), .B1(n5793), .B2(n9898), .ZN(
        P1_U3460) );
  OAI22_X1 U11001 ( .A1(n9856), .A2(n9883), .B1(n9855), .B2(n9881), .ZN(n9858)
         );
  AOI211_X1 U11002 ( .C1(n9860), .C2(n9859), .A(n9858), .B(n9857), .ZN(n9903)
         );
  INV_X1 U11003 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n9861) );
  AOI22_X1 U11004 ( .A1(n9900), .A2(n9903), .B1(n9861), .B2(n9898), .ZN(
        P1_U3466) );
  OAI21_X1 U11005 ( .B1(n9863), .B2(n9881), .A(n9862), .ZN(n9865) );
  AOI211_X1 U11006 ( .C1(n9866), .C2(n9887), .A(n9865), .B(n9864), .ZN(n9904)
         );
  INV_X1 U11007 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n9867) );
  AOI22_X1 U11008 ( .A1(n9900), .A2(n9904), .B1(n9867), .B2(n9898), .ZN(
        P1_U3469) );
  OAI22_X1 U11009 ( .A1(n9869), .A2(n9883), .B1(n9868), .B2(n9881), .ZN(n9871)
         );
  AOI211_X1 U11010 ( .C1(n9887), .C2(n9872), .A(n9871), .B(n9870), .ZN(n9905)
         );
  INV_X1 U11011 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9873) );
  AOI22_X1 U11012 ( .A1(n9900), .A2(n9905), .B1(n9873), .B2(n9898), .ZN(
        P1_U3472) );
  OAI211_X1 U11013 ( .C1(n9876), .C2(n9881), .A(n9875), .B(n9874), .ZN(n9877)
         );
  AOI21_X1 U11014 ( .B1(n9887), .B2(n9878), .A(n9877), .ZN(n9906) );
  AOI22_X1 U11015 ( .A1(n9900), .A2(n9906), .B1(n9879), .B2(n9898), .ZN(
        P1_U3475) );
  INV_X1 U11016 ( .A(n9880), .ZN(n9888) );
  OAI22_X1 U11017 ( .A1(n9884), .A2(n9883), .B1(n9882), .B2(n9881), .ZN(n9886)
         );
  AOI211_X1 U11018 ( .C1(n9888), .C2(n9887), .A(n9886), .B(n9885), .ZN(n9907)
         );
  INV_X1 U11019 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n9889) );
  AOI22_X1 U11020 ( .A1(n9900), .A2(n9907), .B1(n9889), .B2(n9898), .ZN(
        P1_U3478) );
  AOI21_X1 U11021 ( .B1(n9892), .B2(n9891), .A(n9890), .ZN(n9893) );
  OAI21_X1 U11022 ( .B1(n9895), .B2(n9894), .A(n9893), .ZN(n9896) );
  NOR2_X1 U11023 ( .A1(n9897), .A2(n9896), .ZN(n9909) );
  INV_X1 U11024 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9899) );
  AOI22_X1 U11025 ( .A1(n9900), .A2(n9909), .B1(n9899), .B2(n9898), .ZN(
        P1_U3481) );
  AOI22_X1 U11026 ( .A1(n9910), .A2(n9901), .B1(n6361), .B2(n9908), .ZN(
        P1_U3524) );
  AOI22_X1 U11027 ( .A1(n9910), .A2(n9902), .B1(n6364), .B2(n9908), .ZN(
        P1_U3525) );
  AOI22_X1 U11028 ( .A1(n9910), .A2(n9903), .B1(n5848), .B2(n9908), .ZN(
        P1_U3527) );
  AOI22_X1 U11029 ( .A1(n9910), .A2(n9904), .B1(n5869), .B2(n9908), .ZN(
        P1_U3528) );
  AOI22_X1 U11030 ( .A1(n9910), .A2(n9905), .B1(n5890), .B2(n9908), .ZN(
        P1_U3529) );
  AOI22_X1 U11031 ( .A1(n9910), .A2(n9906), .B1(n5911), .B2(n9908), .ZN(
        P1_U3530) );
  AOI22_X1 U11032 ( .A1(n9910), .A2(n9907), .B1(n6369), .B2(n9908), .ZN(
        P1_U3531) );
  AOI22_X1 U11033 ( .A1(n9910), .A2(n9909), .B1(n6370), .B2(n9908), .ZN(
        P1_U3532) );
  OAI211_X1 U11034 ( .C1(n9913), .C2(n9912), .A(n9911), .B(n9949), .ZN(n9921)
         );
  AOI22_X1 U11035 ( .A1(n9915), .A2(n9914), .B1(P2_REG3_REG_10__SCAN_IN), .B2(
        P2_U3152), .ZN(n9920) );
  AOI22_X1 U11036 ( .A1(n9918), .A2(n9917), .B1(n9957), .B2(n9916), .ZN(n9919)
         );
  AND3_X1 U11037 ( .A1(n9921), .A2(n9920), .A3(n9919), .ZN(n9922) );
  OAI21_X1 U11038 ( .B1(n9966), .B2(n9923), .A(n9922), .ZN(P2_U3219) );
  OR2_X1 U11039 ( .A1(n9954), .A2(n9924), .ZN(n9933) );
  OR2_X1 U11040 ( .A1(n9959), .A2(n9925), .ZN(n9932) );
  AOI21_X1 U11041 ( .B1(n9957), .B2(n6754), .A(n9926), .ZN(n9931) );
  NAND2_X1 U11042 ( .A1(n9928), .A2(n9927), .ZN(n9929) );
  NAND3_X1 U11043 ( .A1(n9949), .A2(n9942), .A3(n9929), .ZN(n9930) );
  AND4_X1 U11044 ( .A1(n9933), .A2(n9932), .A3(n9931), .A4(n9930), .ZN(n9934)
         );
  OAI21_X1 U11045 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(n9966), .A(n9934), .ZN(
        P2_U3220) );
  NAND2_X1 U11046 ( .A1(n9936), .A2(n9935), .ZN(n9939) );
  NAND2_X1 U11047 ( .A1(n9937), .A2(n9992), .ZN(n9938) );
  NAND2_X1 U11048 ( .A1(n9939), .A2(n9938), .ZN(n10011) );
  AOI22_X1 U11049 ( .A1(n9940), .A2(n10011), .B1(P2_REG3_REG_4__SCAN_IN), .B2(
        P2_U3152), .ZN(n9948) );
  AND2_X1 U11050 ( .A1(n9942), .A2(n9941), .ZN(n9945) );
  OAI21_X1 U11051 ( .B1(n9945), .B2(n9944), .A(n9943), .ZN(n9946) );
  AOI22_X1 U11052 ( .A1(n9946), .A2(n9949), .B1(n9957), .B2(n10025), .ZN(n9947) );
  OAI211_X1 U11053 ( .C1(n9966), .C2(n10029), .A(n9948), .B(n9947), .ZN(
        P2_U3232) );
  OAI211_X1 U11054 ( .C1(n9952), .C2(n9951), .A(n9950), .B(n9949), .ZN(n9963)
         );
  OAI22_X1 U11055 ( .A1(n9954), .A2(n9953), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5302), .ZN(n9955) );
  INV_X1 U11056 ( .A(n9955), .ZN(n9962) );
  NAND2_X1 U11057 ( .A1(n9957), .A2(n9956), .ZN(n9961) );
  OR2_X1 U11058 ( .A1(n9959), .A2(n9958), .ZN(n9960) );
  OAI21_X1 U11059 ( .B1(n9966), .B2(n9965), .A(n9964), .ZN(P2_U3238) );
  AOI22_X1 U11060 ( .A1(P2_REG2_REG_0__SCAN_IN), .A2(n9968), .B1(n9967), .B2(
        P2_REG1_REG_0__SCAN_IN), .ZN(n9977) );
  AOI22_X1 U11061 ( .A1(n9969), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n9976) );
  NOR2_X1 U11062 ( .A1(n9970), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n9974) );
  OAI21_X1 U11063 ( .B1(n9972), .B2(P2_REG1_REG_0__SCAN_IN), .A(n9971), .ZN(
        n9973) );
  OAI21_X1 U11064 ( .B1(n9974), .B2(n9973), .A(P2_IR_REG_0__SCAN_IN), .ZN(
        n9975) );
  OAI211_X1 U11065 ( .C1(P2_IR_REG_0__SCAN_IN), .C2(n9977), .A(n9976), .B(
        n9975), .ZN(P2_U3245) );
  NAND2_X1 U11066 ( .A1(n9980), .A2(n9990), .ZN(n9981) );
  NAND2_X1 U11067 ( .A1(n9979), .A2(n9981), .ZN(n10081) );
  NAND2_X1 U11068 ( .A1(n9983), .A2(n9982), .ZN(n9984) );
  NAND2_X1 U11069 ( .A1(n9985), .A2(n9984), .ZN(n10083) );
  OAI22_X1 U11070 ( .A1(n10081), .A2(n9987), .B1(n9986), .B2(n10083), .ZN(
        n9988) );
  INV_X1 U11071 ( .A(n9988), .ZN(n10007) );
  OR2_X1 U11072 ( .A1(n10081), .A2(n9989), .ZN(n10000) );
  XNOR2_X1 U11073 ( .A(n9991), .B(n9990), .ZN(n9998) );
  NAND2_X1 U11074 ( .A1(n9993), .A2(n9992), .ZN(n9994) );
  OAI21_X1 U11075 ( .B1(n9996), .B2(n9995), .A(n9994), .ZN(n9997) );
  AOI21_X1 U11076 ( .B1(n9998), .B2(n10012), .A(n9997), .ZN(n9999) );
  NAND2_X1 U11077 ( .A1(n10000), .A2(n9999), .ZN(n10086) );
  NOR2_X1 U11078 ( .A1(n10001), .A2(n10082), .ZN(n10005) );
  OAI22_X1 U11079 ( .A1(n10035), .A2(n10003), .B1(n10002), .B2(n10028), .ZN(
        n10004) );
  AOI211_X1 U11080 ( .C1(n10086), .C2(n10035), .A(n10005), .B(n10004), .ZN(
        n10006) );
  NAND2_X1 U11081 ( .A1(n10007), .A2(n10006), .ZN(P2_U3288) );
  NAND2_X1 U11082 ( .A1(n6783), .A2(n10008), .ZN(n10010) );
  INV_X1 U11083 ( .A(n10014), .ZN(n10009) );
  XNOR2_X1 U11084 ( .A(n10010), .B(n10009), .ZN(n10013) );
  AOI21_X1 U11085 ( .B1(n10013), .B2(n10012), .A(n10011), .ZN(n10068) );
  OR2_X1 U11086 ( .A1(n10015), .A2(n10014), .ZN(n10016) );
  NAND2_X1 U11087 ( .A1(n10017), .A2(n10016), .ZN(n10066) );
  NAND2_X1 U11088 ( .A1(n10066), .A2(n10018), .ZN(n10019) );
  NAND2_X1 U11089 ( .A1(n10068), .A2(n10019), .ZN(n10033) );
  NAND2_X1 U11090 ( .A1(n10020), .A2(n10025), .ZN(n10021) );
  NAND3_X1 U11091 ( .A1(n10023), .A2(n10022), .A3(n10021), .ZN(n10027) );
  NAND2_X1 U11092 ( .A1(n10025), .A2(n10024), .ZN(n10026) );
  NAND2_X1 U11093 ( .A1(n10027), .A2(n10026), .ZN(n10065) );
  INV_X1 U11094 ( .A(n10065), .ZN(n10030) );
  OAI22_X1 U11095 ( .A1(n10031), .A2(n10030), .B1(n10029), .B2(n10028), .ZN(
        n10032) );
  AOI21_X1 U11096 ( .B1(n10033), .B2(n10035), .A(n10032), .ZN(n10034) );
  OAI21_X1 U11097 ( .B1(n10035), .B2(n6478), .A(n10034), .ZN(P2_U3292) );
  AND2_X1 U11098 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n10045), .ZN(P2_U3297) );
  AND2_X1 U11099 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n10045), .ZN(P2_U3298) );
  AND2_X1 U11100 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n10045), .ZN(P2_U3299) );
  AND2_X1 U11101 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n10045), .ZN(P2_U3300) );
  AND2_X1 U11102 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n10045), .ZN(P2_U3301) );
  NOR2_X1 U11103 ( .A1(n10042), .A2(n10038), .ZN(P2_U3302) );
  AND2_X1 U11104 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n10045), .ZN(P2_U3303) );
  AND2_X1 U11105 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n10045), .ZN(P2_U3304) );
  AND2_X1 U11106 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n10045), .ZN(P2_U3305) );
  AND2_X1 U11107 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n10045), .ZN(P2_U3306) );
  AND2_X1 U11108 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n10045), .ZN(P2_U3307) );
  AND2_X1 U11109 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n10045), .ZN(P2_U3308) );
  NOR2_X1 U11110 ( .A1(n10042), .A2(n10039), .ZN(P2_U3309) );
  AND2_X1 U11111 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n10045), .ZN(P2_U3310) );
  AND2_X1 U11112 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n10045), .ZN(P2_U3311) );
  AND2_X1 U11113 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n10045), .ZN(P2_U3312) );
  AND2_X1 U11114 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n10045), .ZN(P2_U3313) );
  AND2_X1 U11115 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n10045), .ZN(P2_U3314) );
  AND2_X1 U11116 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n10045), .ZN(P2_U3315) );
  AND2_X1 U11117 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n10045), .ZN(P2_U3316) );
  NOR2_X1 U11118 ( .A1(n10042), .A2(n10040), .ZN(P2_U3317) );
  NOR2_X1 U11119 ( .A1(n10042), .A2(n10041), .ZN(P2_U3318) );
  AND2_X1 U11120 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n10045), .ZN(P2_U3319) );
  AND2_X1 U11121 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n10045), .ZN(P2_U3320) );
  AND2_X1 U11122 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n10045), .ZN(P2_U3321) );
  AND2_X1 U11123 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n10045), .ZN(P2_U3322) );
  AND2_X1 U11124 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n10045), .ZN(P2_U3323) );
  AND2_X1 U11125 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n10045), .ZN(P2_U3324) );
  AND2_X1 U11126 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n10045), .ZN(P2_U3325) );
  AND2_X1 U11127 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n10045), .ZN(P2_U3326) );
  AOI22_X1 U11128 ( .A1(n10048), .A2(n10044), .B1(n10043), .B2(n10045), .ZN(
        P2_U3437) );
  AOI22_X1 U11129 ( .A1(n10048), .A2(n10047), .B1(n10046), .B2(n10045), .ZN(
        P2_U3438) );
  AOI22_X1 U11130 ( .A1(n10051), .A2(n10114), .B1(n10050), .B2(n10049), .ZN(
        n10052) );
  AND2_X1 U11131 ( .A1(n10053), .A2(n10052), .ZN(n10119) );
  AOI22_X1 U11132 ( .A1(n10117), .A2(n10119), .B1(n5050), .B2(n10115), .ZN(
        P2_U3451) );
  OAI21_X1 U11133 ( .B1(n10055), .B2(n10110), .A(n10054), .ZN(n10058) );
  INV_X1 U11134 ( .A(n10056), .ZN(n10057) );
  AOI211_X1 U11135 ( .C1(n10114), .C2(n10059), .A(n10058), .B(n10057), .ZN(
        n10120) );
  AOI22_X1 U11136 ( .A1(n10117), .A2(n10120), .B1(n5043), .B2(n10115), .ZN(
        P2_U3454) );
  NAND2_X1 U11137 ( .A1(n10061), .A2(n10060), .ZN(n10062) );
  AOI21_X1 U11138 ( .B1(n10114), .B2(n10063), .A(n10062), .ZN(n10121) );
  INV_X1 U11139 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10064) );
  AOI22_X1 U11140 ( .A1(n10117), .A2(n10121), .B1(n10064), .B2(n10115), .ZN(
        P2_U3457) );
  AOI21_X1 U11141 ( .B1(n10066), .B2(n10114), .A(n10065), .ZN(n10067) );
  AND2_X1 U11142 ( .A1(n10068), .A2(n10067), .ZN(n10122) );
  INV_X1 U11143 ( .A(n10122), .ZN(n10069) );
  MUX2_X1 U11144 ( .A(P2_REG0_REG_4__SCAN_IN), .B(n10069), .S(n10117), .Z(
        P2_U3463) );
  OAI22_X1 U11145 ( .A1(n10071), .A2(n10102), .B1(n10070), .B2(n10110), .ZN(
        n10073) );
  AOI211_X1 U11146 ( .C1(n10074), .C2(n10114), .A(n10073), .B(n10072), .ZN(
        n10123) );
  AOI22_X1 U11147 ( .A1(n10117), .A2(n10123), .B1(n5157), .B2(n10115), .ZN(
        P2_U3469) );
  OAI22_X1 U11148 ( .A1(n10076), .A2(n10102), .B1(n10075), .B2(n10110), .ZN(
        n10078) );
  AOI211_X1 U11149 ( .C1(n10114), .C2(n10079), .A(n10078), .B(n10077), .ZN(
        n10125) );
  AOI22_X1 U11150 ( .A1(n10117), .A2(n10125), .B1(n5175), .B2(n10115), .ZN(
        P2_U3472) );
  NOR2_X1 U11151 ( .A1(n10081), .A2(n10080), .ZN(n10085) );
  OAI22_X1 U11152 ( .A1(n10083), .A2(n10102), .B1(n10082), .B2(n10110), .ZN(
        n10084) );
  NOR3_X1 U11153 ( .A1(n10086), .A2(n10085), .A3(n10084), .ZN(n10126) );
  AOI22_X1 U11154 ( .A1(n10117), .A2(n10126), .B1(n5212), .B2(n10115), .ZN(
        P2_U3475) );
  OAI22_X1 U11155 ( .A1(n10088), .A2(n10102), .B1(n10087), .B2(n10110), .ZN(
        n10090) );
  AOI211_X1 U11156 ( .C1(n10114), .C2(n10091), .A(n10090), .B(n10089), .ZN(
        n10127) );
  INV_X1 U11157 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10092) );
  AOI22_X1 U11158 ( .A1(n10117), .A2(n10127), .B1(n10092), .B2(n10115), .ZN(
        P2_U3478) );
  OAI22_X1 U11159 ( .A1(n10094), .A2(n10102), .B1(n10093), .B2(n10110), .ZN(
        n10095) );
  AOI21_X1 U11160 ( .B1(n10097), .B2(n10096), .A(n10095), .ZN(n10098) );
  AND2_X1 U11161 ( .A1(n10099), .A2(n10098), .ZN(n10129) );
  AOI22_X1 U11162 ( .A1(n10117), .A2(n10129), .B1(n5258), .B2(n10115), .ZN(
        P2_U3481) );
  INV_X1 U11163 ( .A(n10100), .ZN(n10106) );
  OAI22_X1 U11164 ( .A1(n10103), .A2(n10102), .B1(n10101), .B2(n10110), .ZN(
        n10105) );
  AOI211_X1 U11165 ( .C1(n10106), .C2(n10114), .A(n10105), .B(n10104), .ZN(
        n10130) );
  INV_X1 U11166 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10107) );
  AOI22_X1 U11167 ( .A1(n10117), .A2(n10130), .B1(n10107), .B2(n10115), .ZN(
        P2_U3484) );
  OAI211_X1 U11168 ( .C1(n10111), .C2(n10110), .A(n10109), .B(n10108), .ZN(
        n10112) );
  AOI21_X1 U11169 ( .B1(n10114), .B2(n10113), .A(n10112), .ZN(n10132) );
  AOI22_X1 U11170 ( .A1(n10117), .A2(n10132), .B1(n10116), .B2(n10115), .ZN(
        P2_U3487) );
  INV_X1 U11171 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10118) );
  AOI22_X1 U11172 ( .A1(n10124), .A2(n10119), .B1(n10118), .B2(n10131), .ZN(
        P2_U3520) );
  AOI22_X1 U11173 ( .A1(n10124), .A2(n10120), .B1(n6465), .B2(n10131), .ZN(
        P2_U3521) );
  AOI22_X1 U11174 ( .A1(n10124), .A2(n10121), .B1(n6466), .B2(n10131), .ZN(
        P2_U3522) );
  AOI22_X1 U11175 ( .A1(n10124), .A2(n10122), .B1(n6468), .B2(n10131), .ZN(
        P2_U3524) );
  AOI22_X1 U11176 ( .A1(n10124), .A2(n10123), .B1(n6470), .B2(n10131), .ZN(
        P2_U3526) );
  AOI22_X1 U11177 ( .A1(n10124), .A2(n10125), .B1(n6506), .B2(n10131), .ZN(
        P2_U3527) );
  AOI22_X1 U11178 ( .A1(n10124), .A2(n10126), .B1(n8362), .B2(n10131), .ZN(
        P2_U3528) );
  AOI22_X1 U11179 ( .A1(n10124), .A2(n10127), .B1(n6523), .B2(n10131), .ZN(
        P2_U3529) );
  AOI22_X1 U11180 ( .A1(n10124), .A2(n10129), .B1(n10128), .B2(n10131), .ZN(
        P2_U3530) );
  AOI22_X1 U11181 ( .A1(n10124), .A2(n10130), .B1(n5275), .B2(n10131), .ZN(
        P2_U3531) );
  AOI22_X1 U11182 ( .A1(n10124), .A2(n10132), .B1(n6685), .B2(n10131), .ZN(
        P2_U3532) );
  OAI21_X1 U11183 ( .B1(n10135), .B2(n6608), .A(n10133), .ZN(n10134) );
  XNOR2_X1 U11184 ( .A(n10134), .B(P2_ADDR_REG_1__SCAN_IN), .ZN(ADD_1071_U5)
         );
  OAI21_X1 U11185 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(P2_ADDR_REG_0__SCAN_IN), 
        .A(n10135), .ZN(n10136) );
  INV_X1 U11186 ( .A(n10136), .ZN(ADD_1071_U46) );
  OAI21_X1 U11187 ( .B1(n10139), .B2(n10138), .A(n10137), .ZN(ADD_1071_U56) );
  OAI21_X1 U11188 ( .B1(n10142), .B2(n10141), .A(n10140), .ZN(ADD_1071_U57) );
  OAI21_X1 U11189 ( .B1(n10145), .B2(n10144), .A(n10143), .ZN(ADD_1071_U58) );
  OAI21_X1 U11190 ( .B1(n10148), .B2(n10147), .A(n10146), .ZN(ADD_1071_U59) );
  OAI21_X1 U11191 ( .B1(n10151), .B2(n10150), .A(n10149), .ZN(ADD_1071_U60) );
  OAI21_X1 U11192 ( .B1(n10154), .B2(n10153), .A(n10152), .ZN(ADD_1071_U61) );
  AOI21_X1 U11193 ( .B1(n10157), .B2(n10156), .A(n10155), .ZN(ADD_1071_U62) );
  AOI21_X1 U11194 ( .B1(n10160), .B2(n10159), .A(n10158), .ZN(ADD_1071_U63) );
  AOI21_X1 U11195 ( .B1(n10163), .B2(n10162), .A(n10161), .ZN(ADD_1071_U48) );
  AOI21_X1 U11196 ( .B1(n10166), .B2(n10165), .A(n10164), .ZN(ADD_1071_U50) );
  OAI222_X1 U11197 ( .A1(n10171), .A2(n10170), .B1(n10171), .B2(n10169), .C1(
        n10168), .C2(n10167), .ZN(ADD_1071_U51) );
  AOI21_X1 U11198 ( .B1(n10174), .B2(n10173), .A(n10172), .ZN(ADD_1071_U49) );
  OAI21_X1 U11199 ( .B1(n10177), .B2(n10176), .A(n10175), .ZN(n10178) );
  XNOR2_X1 U11200 ( .A(n10178), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  AOI21_X1 U11201 ( .B1(n10181), .B2(n10180), .A(n10179), .ZN(ADD_1071_U47) );
  AOI21_X1 U11202 ( .B1(n10184), .B2(n10183), .A(n10182), .ZN(ADD_1071_U54) );
  AOI21_X1 U11203 ( .B1(n10187), .B2(n10186), .A(n10185), .ZN(ADD_1071_U53) );
  OAI21_X1 U11204 ( .B1(n10190), .B2(n10189), .A(n10188), .ZN(ADD_1071_U52) );
  XNOR2_X1 U6563 ( .A(n5039), .B(n5036), .ZN(n7526) );
  INV_X1 U4897 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n6084) );
  NAND2_X2 U7334 ( .A1(n6828), .A2(n6321), .ZN(n5830) );
  CLKBUF_X1 U4893 ( .A(n5755), .Z(n5754) );
  CLKBUF_X1 U5056 ( .A(n5406), .Z(n6430) );
  CLKBUF_X1 U5223 ( .A(n8153), .Z(n4476) );
  CLKBUF_X1 U5986 ( .A(n6007), .Z(n6254) );
endmodule

