

module b20_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, P2_WR_REG_SCAN_IN, SI_31_, 
        SI_30_, SI_29_, SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, 
        SI_21_, SI_20_, SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, 
        SI_12_, SI_11_, SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, 
        SI_3_, SI_2_, SI_1_, SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, ADD_1068_U4, 
        ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, 
        ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, 
        ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, 
        ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, U126, U123, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, P1_U3468, 
        P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, 
        P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3509, 
        P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, 
        P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, 
        P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, 
        P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, 
        P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, 
        P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, 
        P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, P1_U3555, 
        P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, 
        P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, 
        P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, 
        P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, 
        P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U3973, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, P2_U3263, 
        P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, 
        P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, 
        P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, 
        P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, 
        P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, P2_U3405, 
        P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, P2_U3426, 
        P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, P2_U3446, 
        P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, P2_U3453, 
        P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, P2_U3460, 
        P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, P2_U3467, 
        P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, P2_U3474, 
        P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, P2_U3481, 
        P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, P2_U3488, 
        P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, 
        P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, 
        P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, 
        P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, P2_U3492, 
        P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, 
        P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, P2_U3178, 
        P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, 
        P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, 
        P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, 
        P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, P2_U3893
 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_,
         SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_,
         SI_20_, SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_,
         SI_12_, SI_11_, SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_,
         SI_3_, SI_2_, SI_1_, SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_REG3_REG_7__SCAN_IN, P2_REG3_REG_27__SCAN_IN,
         P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_23__SCAN_IN,
         P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_3__SCAN_IN,
         P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_28__SCAN_IN,
         P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_1__SCAN_IN,
         P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_12__SCAN_IN,
         P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_16__SCAN_IN,
         P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_17__SCAN_IN,
         P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_4__SCAN_IN,
         P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN,
         P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN,
         P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN,
         P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN,
         P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN,
         P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933,
         n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943,
         n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953,
         n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963,
         n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973,
         n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983,
         n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993,
         n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003,
         n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013,
         n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023,
         n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033,
         n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043,
         n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053,
         n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063,
         n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073,
         n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083,
         n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093,
         n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103,
         n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113,
         n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123,
         n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133,
         n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143,
         n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153,
         n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163,
         n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173,
         n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183,
         n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193,
         n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203,
         n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213,
         n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223,
         n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233,
         n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243,
         n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253,
         n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263,
         n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273,
         n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283,
         n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293,
         n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303,
         n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313,
         n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323,
         n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333,
         n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343,
         n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353,
         n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363,
         n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373,
         n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383,
         n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393,
         n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403,
         n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413,
         n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423,
         n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433,
         n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443,
         n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453,
         n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463,
         n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473,
         n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483,
         n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493,
         n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503,
         n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513,
         n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523,
         n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533,
         n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543,
         n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553,
         n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563,
         n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573,
         n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583,
         n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593,
         n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603,
         n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613,
         n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623,
         n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633,
         n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643,
         n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653,
         n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663,
         n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673,
         n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683,
         n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693,
         n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703,
         n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713,
         n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723,
         n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733,
         n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743,
         n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753,
         n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763,
         n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773,
         n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783,
         n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793,
         n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803,
         n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813,
         n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823,
         n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833,
         n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843,
         n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853,
         n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863,
         n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873,
         n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883,
         n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893,
         n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903,
         n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913,
         n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923,
         n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933,
         n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943,
         n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953,
         n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963,
         n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973,
         n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983,
         n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993,
         n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003,
         n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013,
         n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023,
         n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033,
         n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043,
         n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053,
         n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063,
         n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073,
         n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083,
         n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093,
         n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103,
         n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113,
         n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123,
         n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133,
         n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143,
         n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153,
         n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163,
         n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173,
         n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183,
         n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193,
         n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203,
         n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213,
         n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223,
         n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233,
         n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243,
         n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253,
         n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263,
         n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273,
         n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283,
         n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293,
         n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303,
         n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313,
         n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323,
         n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333,
         n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343,
         n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353,
         n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363,
         n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373,
         n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383,
         n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393,
         n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403,
         n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413,
         n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423,
         n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433,
         n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443,
         n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453,
         n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463,
         n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473,
         n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483,
         n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493,
         n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503,
         n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513,
         n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523,
         n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533,
         n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543,
         n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553,
         n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563,
         n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573,
         n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583,
         n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593,
         n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603,
         n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613,
         n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623,
         n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633,
         n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643,
         n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653,
         n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663,
         n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673,
         n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683,
         n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693,
         n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703,
         n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713,
         n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723,
         n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733,
         n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743,
         n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753,
         n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763,
         n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773,
         n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783,
         n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793,
         n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803,
         n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813,
         n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823,
         n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833,
         n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843,
         n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853,
         n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863,
         n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873,
         n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883,
         n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893,
         n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903,
         n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913,
         n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923,
         n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933,
         n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943,
         n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953,
         n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963,
         n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973,
         n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983,
         n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993,
         n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003,
         n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013,
         n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023,
         n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033,
         n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043,
         n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053,
         n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063,
         n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073,
         n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083,
         n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093,
         n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103,
         n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113,
         n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123,
         n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133,
         n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143,
         n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153,
         n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163,
         n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173,
         n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183,
         n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193,
         n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203,
         n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213,
         n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223,
         n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233,
         n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243,
         n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253,
         n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263,
         n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273,
         n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283,
         n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293,
         n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303,
         n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313,
         n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323,
         n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333,
         n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343,
         n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353,
         n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363,
         n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373,
         n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383,
         n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393,
         n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403,
         n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413,
         n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423,
         n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433,
         n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443,
         n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453,
         n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463,
         n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473,
         n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483,
         n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493,
         n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503,
         n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513,
         n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523,
         n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533,
         n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543,
         n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553,
         n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563,
         n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573,
         n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583,
         n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593,
         n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603,
         n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613,
         n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623,
         n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633,
         n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643,
         n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653,
         n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663,
         n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673,
         n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683,
         n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693,
         n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703,
         n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713,
         n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723,
         n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733,
         n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743,
         n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753,
         n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763,
         n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773,
         n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783,
         n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793,
         n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803,
         n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813,
         n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823,
         n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833,
         n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843,
         n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853,
         n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863,
         n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873,
         n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883,
         n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893,
         n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903,
         n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913,
         n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923,
         n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933,
         n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943,
         n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953,
         n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963,
         n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973,
         n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983,
         n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993,
         n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003,
         n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013,
         n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023,
         n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033,
         n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043,
         n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053,
         n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063,
         n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073,
         n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083,
         n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093,
         n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103,
         n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113,
         n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123,
         n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133,
         n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143,
         n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153,
         n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163,
         n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173,
         n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183,
         n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193,
         n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203,
         n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213,
         n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223,
         n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233,
         n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243,
         n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253,
         n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263,
         n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273,
         n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283,
         n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293,
         n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303,
         n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313,
         n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323,
         n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333,
         n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343,
         n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353,
         n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363,
         n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373,
         n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383,
         n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393,
         n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403,
         n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413,
         n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423,
         n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433,
         n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443,
         n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453,
         n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463,
         n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473,
         n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483,
         n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493,
         n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503,
         n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513,
         n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523,
         n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533,
         n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543,
         n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553,
         n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563,
         n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573,
         n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583,
         n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593,
         n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603,
         n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613,
         n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623,
         n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633,
         n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643,
         n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653,
         n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663,
         n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673,
         n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683,
         n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693,
         n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703,
         n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713,
         n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723,
         n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733,
         n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743,
         n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753,
         n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763,
         n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773,
         n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783,
         n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793,
         n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803,
         n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813,
         n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823,
         n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833,
         n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843,
         n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853,
         n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863,
         n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873,
         n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883,
         n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893,
         n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903,
         n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913,
         n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923,
         n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933,
         n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943,
         n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953,
         n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963,
         n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973,
         n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983,
         n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993,
         n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003,
         n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013,
         n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023,
         n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033,
         n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043,
         n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053,
         n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063,
         n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073,
         n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083,
         n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093,
         n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103,
         n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113,
         n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123,
         n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133,
         n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143,
         n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153,
         n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163,
         n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173,
         n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183,
         n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193,
         n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203,
         n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213,
         n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223,
         n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233,
         n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243,
         n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253,
         n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263,
         n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273,
         n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283,
         n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293,
         n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303,
         n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313,
         n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323,
         n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333,
         n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343,
         n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353,
         n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363,
         n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373,
         n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383,
         n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393,
         n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403,
         n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413,
         n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423,
         n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433,
         n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443,
         n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453,
         n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463,
         n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473,
         n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483,
         n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493,
         n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503,
         n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513,
         n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523,
         n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533,
         n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543,
         n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553,
         n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563,
         n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573,
         n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583,
         n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593,
         n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603,
         n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613,
         n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623,
         n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633,
         n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643,
         n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653,
         n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663,
         n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673,
         n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683,
         n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693,
         n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703,
         n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713,
         n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723,
         n9724, n9725, n9726, n9727, n9728, n9730, n9731, n9732, n9733, n9734,
         n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744,
         n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754,
         n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764,
         n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774,
         n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784,
         n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794,
         n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804,
         n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814,
         n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824,
         n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834,
         n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844,
         n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854,
         n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864,
         n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874,
         n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884,
         n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894,
         n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904,
         n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914,
         n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924,
         n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934,
         n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944,
         n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954,
         n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964,
         n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974,
         n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984,
         n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994,
         n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003,
         n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011,
         n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019,
         n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027,
         n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035,
         n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043,
         n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051,
         n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059,
         n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067,
         n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075,
         n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083,
         n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091,
         n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099,
         n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107,
         n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115,
         n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123,
         n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131,
         n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139,
         n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147,
         n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155,
         n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163,
         n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171,
         n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179,
         n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187,
         n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195,
         n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203,
         n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211,
         n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219,
         n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227,
         n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235,
         n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243,
         n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251,
         n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259,
         n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267,
         n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275,
         n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283,
         n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291,
         n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299,
         n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307,
         n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315,
         n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323,
         n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331,
         n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339,
         n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347,
         n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355,
         n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363,
         n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371,
         n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379,
         n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387,
         n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395,
         n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403,
         n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411,
         n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419,
         n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427,
         n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435,
         n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443,
         n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451,
         n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459,
         n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467,
         n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475,
         n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483,
         n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491,
         n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499,
         n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507,
         n10508, n10509, n10510, n10511, n10512, n10513, n10514, n10515,
         n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523,
         n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531,
         n10532, n10533, n10534, n10535, n10536, n10537, n10538, n10539,
         n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547,
         n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555,
         n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563,
         n10564, n10565, n10566, n10567, n10568, n10569, n10570, n10571,
         n10572, n10573, n10574, n10575, n10576, n10577, n10578, n10579,
         n10580, n10581, n10582, n10583, n10584, n10585, n10586, n10587,
         n10588, n10589, n10590, n10591, n10592, n10593, n10594, n10595,
         n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603,
         n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10611,
         n10612, n10613, n10614, n10615, n10616, n10617, n10618, n10619,
         n10620, n10621, n10622, n10623, n10624, n10625, n10626, n10627,
         n10628, n10629, n10630, n10631, n10632, n10633, n10634, n10635,
         n10636, n10637, n10638, n10639, n10640, n10641, n10642, n10643,
         n10644, n10645, n10646, n10647, n10648, n10649, n10650, n10651,
         n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659,
         n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667,
         n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675,
         n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10683,
         n10684, n10685, n10686, n10687, n10688, n10689, n10690, n10691,
         n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699,
         n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707,
         n10708, n10709, n10710, n10711, n10712, n10713, n10714, n10715,
         n10716, n10717, n10718, n10719, n10720, n10721, n10722, n10723,
         n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731,
         n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739,
         n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747,
         n10748, n10749, n10750, n10751, n10752, n10753, n10754, n10755,
         n10756, n10757, n10758, n10759, n10760, n10761, n10762, n10763,
         n10764;

  OAI21_X1 U4988 ( .B1(n5980), .B2(n5979), .A(n5978), .ZN(n5995) );
  CLKBUF_X2 U4989 ( .A(n8488), .Z(n4926) );
  CLKBUF_X3 U4990 ( .A(n5756), .Z(n4930) );
  XNOR2_X1 U4991 ( .A(n5569), .B(n5739), .ZN(n5648) );
  CLKBUF_X1 U4992 ( .A(n10558), .Z(n4924) );
  NOR2_X1 U4993 ( .A1(n6825), .A2(n4926), .ZN(n10558) );
  AND2_X1 U4994 ( .A1(n7810), .A2(n8286), .ZN(n8282) );
  INV_X2 U4995 ( .A(n8396), .ZN(n8387) );
  INV_X1 U4996 ( .A(n6936), .ZN(n7067) );
  INV_X1 U4997 ( .A(n8416), .ZN(n5046) );
  INV_X1 U4998 ( .A(n5765), .ZN(n6051) );
  INV_X2 U4999 ( .A(n6996), .ZN(n8745) );
  AOI21_X1 U5000 ( .B1(n7499), .B2(n7924), .A(n7415), .ZN(n7528) );
  NAND2_X1 U5001 ( .A1(n8820), .A2(n4997), .ZN(n8874) );
  XNOR2_X1 U5002 ( .A(n8439), .B(n4966), .ZN(n6294) );
  INV_X1 U5003 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5617) );
  XNOR2_X1 U5004 ( .A(n5478), .B(n5741), .ZN(n5744) );
  NAND2_X1 U5005 ( .A1(n6890), .A2(n6887), .ZN(n8743) );
  INV_X1 U5006 ( .A(n7122), .ZN(n6616) );
  NAND2_X1 U5007 ( .A1(n5561), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5563) );
  NAND2_X1 U5008 ( .A1(n5560), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6242) );
  INV_X1 U5009 ( .A(n6386), .ZN(n6579) );
  NAND4_X1 U5010 ( .A1(n5803), .A2(n5802), .A3(n5801), .A4(n5800), .ZN(n8939)
         );
  OAI211_X1 U5011 ( .C1(n5651), .C2(n5596), .A(n5595), .B(n5597), .ZN(n7289)
         );
  XNOR2_X1 U5012 ( .A(n6615), .B(P1_IR_REG_19__SCAN_IN), .ZN(n8488) );
  OR2_X1 U5013 ( .A1(n6249), .A2(n7499), .ZN(n8255) );
  NAND4_X2 U5014 ( .A1(n5760), .A2(n5759), .A3(n5758), .A4(n5757), .ZN(n6249)
         );
  BUF_X4 U5015 ( .A(n7289), .Z(n4925) );
  NOR2_X2 U5016 ( .A1(n10456), .A2(n10455), .ZN(n10454) );
  XNOR2_X2 U5017 ( .A(n5187), .B(n7145), .ZN(n10455) );
  AOI211_X2 U5018 ( .C1(n8376), .C2(n8375), .A(n8374), .B(n9080), .ZN(n8381)
         );
  XNOR2_X1 U5019 ( .A(n8941), .B(n8266), .ZN(n7760) );
  NAND4_X4 U5020 ( .A1(n5770), .A2(n5769), .A3(n5768), .A4(n5767), .ZN(n8941)
         );
  INV_X1 U5021 ( .A(n6889), .ZN(n8635) );
  NOR4_X2 U5022 ( .A1(n9117), .A2(n9080), .A3(n8467), .A4(n9050), .ZN(n8468)
         );
  NAND2_X2 U5023 ( .A1(n6891), .A2(n6890), .ZN(n8744) );
  OAI21_X2 U5024 ( .B1(n9172), .B2(n6277), .A(n6278), .ZN(n9160) );
  OAI22_X2 U5025 ( .A1(n7718), .A2(n7717), .B1(n7716), .B2(n8938), .ZN(n7719)
         );
  XNOR2_X2 U5026 ( .A(n5842), .B(n5841), .ZN(n5840) );
  NAND2_X2 U5027 ( .A1(n5826), .A2(n5825), .ZN(n5842) );
  INV_X1 U5028 ( .A(n8940), .ZN(n7438) );
  XNOR2_X2 U5029 ( .A(n5663), .B(n10418), .ZN(n10420) );
  NOR2_X2 U5030 ( .A1(n10395), .A2(n5662), .ZN(n5663) );
  NOR2_X1 U5031 ( .A1(n6848), .A2(n6847), .ZN(n6873) );
  NAND3_X1 U5032 ( .A1(n6293), .A2(n6292), .A3(n6291), .ZN(n6848) );
  NAND2_X1 U5033 ( .A1(n7854), .A2(n7856), .ZN(n7855) );
  INV_X2 U5034 ( .A(n7984), .ZN(n7924) );
  NAND2_X1 U5035 ( .A1(n5854), .A2(n5853), .ZN(n10619) );
  OR2_X1 U5036 ( .A1(n8937), .A2(n7715), .ZN(n8301) );
  NAND2_X1 U5037 ( .A1(n8263), .A2(n8256), .ZN(n6248) );
  NAND2_X1 U5038 ( .A1(n8295), .A2(n8276), .ZN(n8447) );
  NAND4_X1 U5039 ( .A1(n5784), .A2(n5783), .A3(n5782), .A4(n5781), .ZN(n8940)
         );
  AND4_X2 U5040 ( .A1(n5749), .A2(n5748), .A3(n5747), .A4(n5746), .ZN(n7628)
         );
  INV_X2 U5041 ( .A(n7366), .ZN(n6373) );
  NAND2_X2 U5042 ( .A1(n7409), .A2(n8479), .ZN(n7765) );
  INV_X2 U5043 ( .A(n8744), .ZN(n6919) );
  INV_X2 U5044 ( .A(n4931), .ZN(n4932) );
  INV_X2 U5045 ( .A(n4930), .ZN(n8424) );
  OR2_X1 U5046 ( .A1(n5744), .A2(n5745), .ZN(n6208) );
  AND2_X1 U5047 ( .A1(n9341), .A2(n5744), .ZN(n5756) );
  XNOR2_X1 U5048 ( .A(n5743), .B(n5742), .ZN(n5745) );
  NOR2_X1 U5049 ( .A1(n9039), .A2(n5006), .ZN(n5043) );
  OR2_X1 U5050 ( .A1(n8478), .A2(n7410), .ZN(n5287) );
  NAND2_X1 U5051 ( .A1(n5257), .A2(n5254), .ZN(n9255) );
  OAI21_X1 U5052 ( .B1(n6797), .B2(n10678), .A(n5177), .ZN(n6800) );
  OAI21_X1 U5053 ( .B1(n6797), .B2(n10676), .A(n5331), .ZN(n6795) );
  OAI21_X1 U5054 ( .B1(n9052), .B2(n4942), .A(n4979), .ZN(n5029) );
  NAND2_X1 U5055 ( .A1(n5259), .A2(n6286), .ZN(n9052) );
  OR2_X1 U5056 ( .A1(n6294), .A2(n10683), .ZN(n6293) );
  OR2_X1 U5057 ( .A1(n8386), .A2(n8385), .ZN(n5205) );
  NAND2_X1 U5058 ( .A1(n5225), .A2(n8592), .ZN(n8595) );
  OAI21_X1 U5059 ( .B1(n9105), .B2(n5038), .A(n5037), .ZN(n9081) );
  NAND2_X1 U5060 ( .A1(n9127), .A2(n8355), .ZN(n9112) );
  OR2_X1 U5061 ( .A1(n9669), .A2(n9667), .ZN(n9670) );
  NAND2_X1 U5062 ( .A1(n8822), .A2(n8821), .ZN(n8820) );
  NAND2_X1 U5063 ( .A1(n6276), .A2(n6275), .ZN(n9172) );
  AOI21_X1 U5064 ( .B1(n6958), .B2(n5079), .A(n5076), .ZN(n8138) );
  AND2_X1 U5065 ( .A1(n6957), .A2(n5077), .ZN(n5076) );
  NAND2_X1 U5066 ( .A1(n5291), .A2(n5290), .ZN(n5289) );
  NAND2_X1 U5067 ( .A1(n7976), .A2(n5476), .ZN(n8098) );
  NAND2_X1 U5068 ( .A1(n5099), .A2(n7821), .ZN(n5098) );
  NAND2_X1 U5069 ( .A1(n7926), .A2(n7925), .ZN(n7976) );
  NAND2_X1 U5070 ( .A1(n8163), .A2(n5673), .ZN(n8164) );
  OR2_X1 U5071 ( .A1(n6661), .A2(n9365), .ZN(n6670) );
  AND2_X1 U5072 ( .A1(n7801), .A2(n4998), .ZN(n9825) );
  AND2_X1 U5073 ( .A1(n5481), .A2(n4999), .ZN(n7718) );
  OR2_X1 U5074 ( .A1(n7576), .A2(n8695), .ZN(n7631) );
  OR2_X1 U5075 ( .A1(n7654), .A2(n7657), .ZN(n7599) );
  OAI21_X1 U5076 ( .B1(n5181), .B2(n5669), .A(n5182), .ZN(n5183) );
  AND2_X1 U5077 ( .A1(n6149), .A2(n8867), .ZN(n6167) );
  NAND2_X1 U5078 ( .A1(n5210), .A2(n5871), .ZN(n10642) );
  OAI21_X1 U5079 ( .B1(n5995), .B2(n5994), .A(n5993), .ZN(n6014) );
  AND2_X1 U5080 ( .A1(n5846), .A2(n5845), .ZN(n7715) );
  INV_X1 U5081 ( .A(n10571), .ZN(n7523) );
  OR2_X1 U5082 ( .A1(n7155), .A2(P2_D_REG_0__SCAN_IN), .ZN(n6304) );
  NAND4_X1 U5083 ( .A1(n6390), .A2(n6389), .A3(n6388), .A4(n6387), .ZN(n10544)
         );
  CLKBUF_X1 U5084 ( .A(n9821), .Z(n10541) );
  NAND4_X1 U5085 ( .A1(n6380), .A2(n6379), .A3(n6378), .A4(n6377), .ZN(n9512)
         );
  INV_X1 U5086 ( .A(n6896), .ZN(n6996) );
  AND3_X1 U5087 ( .A1(n5797), .A2(n5796), .A3(n5795), .ZN(n10577) );
  AND3_X1 U5088 ( .A1(n4989), .A2(n5317), .A3(n5316), .ZN(n8266) );
  INV_X2 U5089 ( .A(n8743), .ZN(n7069) );
  OR2_X1 U5090 ( .A1(n6517), .A2(n7358), .ZN(n6531) );
  NAND2_X1 U5091 ( .A1(n5808), .A2(n5807), .ZN(n5823) );
  NAND2_X1 U5092 ( .A1(n5765), .A2(n7103), .ZN(n5793) );
  NAND2_X1 U5093 ( .A1(n5765), .A2(n8416), .ZN(n5785) );
  NAND2_X2 U5094 ( .A1(n9339), .A2(n5745), .ZN(n5857) );
  INV_X1 U5095 ( .A(n5798), .ZN(n4931) );
  AND2_X2 U5096 ( .A1(n6342), .A2(n10009), .ZN(n8491) );
  XNOR2_X1 U5097 ( .A(n5546), .B(n5545), .ZN(n8240) );
  NAND2_X4 U5098 ( .A1(n7174), .A2(n9525), .ZN(n7122) );
  XNOR2_X1 U5099 ( .A(n5550), .B(n5549), .ZN(n6298) );
  NAND2_X1 U5100 ( .A1(n5790), .A2(n5789), .ZN(n5805) );
  MUX2_X1 U5101 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5571), .S(
        P2_IR_REG_27__SCAN_IN), .Z(n5572) );
  NAND2_X1 U5102 ( .A1(n9335), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5478) );
  MUX2_X1 U5103 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6361), .S(
        P1_IR_REG_28__SCAN_IN), .Z(n6362) );
  INV_X1 U5104 ( .A(n7900), .ZN(n5182) );
  NAND2_X1 U5105 ( .A1(n5556), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5575) );
  OR2_X1 U5106 ( .A1(n5740), .A2(n5617), .ZN(n5569) );
  AND2_X1 U5107 ( .A1(n7290), .A2(n7291), .ZN(n7293) );
  OR2_X1 U5108 ( .A1(n4995), .A2(n5617), .ZN(n5551) );
  AND2_X1 U5109 ( .A1(n6333), .A2(n6735), .ZN(n5475) );
  OAI21_X1 U5110 ( .B1(n8416), .B2(n5751), .A(n5750), .ZN(n5773) );
  NOR2_X1 U5111 ( .A1(n6332), .A2(P1_IR_REG_23__SCAN_IN), .ZN(n6333) );
  NAND2_X2 U5112 ( .A1(n7103), .A2(P1_U3086), .ZN(n7945) );
  AND2_X1 U5113 ( .A1(n5873), .A2(n5872), .ZN(n5889) );
  INV_X2 U5114 ( .A(n8416), .ZN(n7103) );
  AND4_X1 U5115 ( .A1(n5312), .A2(n5533), .A3(n5504), .A4(n5506), .ZN(n5311)
         );
  NAND2_X2 U5116 ( .A1(n8416), .A2(P2_U3151), .ZN(n8052) );
  OAI21_X1 U5117 ( .B1(n5696), .B2(n5652), .A(n5653), .ZN(n7270) );
  NAND2_X1 U5118 ( .A1(n5186), .A2(n5184), .ZN(n5696) );
  INV_X1 U5119 ( .A(n5597), .ZN(n5533) );
  AND3_X1 U5120 ( .A1(n6506), .A2(n6567), .A3(n5108), .ZN(n5176) );
  AND2_X1 U5121 ( .A1(n5537), .A2(n5538), .ZN(n5506) );
  NAND4_X1 U5122 ( .A1(n5539), .A2(n5579), .A3(n5629), .A4(n5576), .ZN(n5557)
         );
  AND2_X1 U5123 ( .A1(n5321), .A2(n6324), .ZN(n5175) );
  NAND3_X1 U5124 ( .A1(n5594), .A2(n5265), .A3(n5264), .ZN(n5597) );
  NAND3_X1 U5125 ( .A1(n5383), .A2(n5382), .A3(n5381), .ZN(n5380) );
  NAND3_X1 U5126 ( .A1(n5384), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n5379) );
  AND4_X1 U5127 ( .A1(n5313), .A2(n5534), .A3(n5536), .A4(n5535), .ZN(n5312)
         );
  NOR2_X1 U5128 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n6506) );
  INV_X2 U5129 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  NOR2_X1 U5130 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n6567) );
  INV_X1 U5131 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5629) );
  INV_X1 U5132 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5641) );
  INV_X1 U5133 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5555) );
  NOR2_X1 U5134 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n5108) );
  NOR2_X2 U5135 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n6381) );
  INV_X1 U5136 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5537) );
  NOR2_X1 U5137 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n5106) );
  INV_X1 U5138 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n6603) );
  NOR2_X1 U5139 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n5313) );
  NOR2_X1 U5140 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n5539) );
  NOR2_X2 U5141 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n5470) );
  INV_X1 U5142 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5579) );
  INV_X1 U5143 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5594) );
  INV_X1 U5144 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n6773) );
  INV_X1 U5145 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5384) );
  NOR2_X2 U5146 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n5651) );
  INV_X1 U5147 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5559) );
  NOR2_X1 U5148 ( .A1(n6248), .A2(n5244), .ZN(n5241) );
  OAI21_X1 U5149 ( .B1(n5049), .B2(n6248), .A(n8259), .ZN(n7785) );
  NAND2_X1 U5150 ( .A1(n5501), .A2(n5500), .ZN(n7923) );
  NAND2_X1 U5151 ( .A1(n5573), .A2(n5572), .ZN(n4927) );
  NAND2_X1 U5152 ( .A1(n5573), .A2(n5572), .ZN(n4928) );
  NAND2_X1 U5153 ( .A1(n5573), .A2(n5572), .ZN(n8480) );
  AND2_X4 U5154 ( .A1(n7122), .A2(n8416), .ZN(n6405) );
  BUF_X4 U5155 ( .A(n6208), .Z(n4929) );
  AND2_X1 U5156 ( .A1(n5744), .A2(n5745), .ZN(n5798) );
  NAND2_X1 U5157 ( .A1(n9339), .A2(n5745), .ZN(n4933) );
  NAND2_X1 U5158 ( .A1(n5197), .A2(n8387), .ZN(n5196) );
  NAND2_X1 U5159 ( .A1(n8260), .A2(n8387), .ZN(n8272) );
  INV_X1 U5160 ( .A(n8336), .ZN(n5338) );
  INV_X1 U5161 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5504) );
  AOI21_X1 U5162 ( .B1(n5843), .B2(n5839), .A(n5848), .ZN(n5061) );
  NOR2_X1 U5163 ( .A1(n4971), .A2(n5248), .ZN(n5247) );
  INV_X1 U5164 ( .A(n6282), .ZN(n5248) );
  AOI21_X1 U5165 ( .B1(n8355), .B2(n8356), .A(n8354), .ZN(n5351) );
  NAND2_X1 U5166 ( .A1(n5070), .A2(n4970), .ZN(n5069) );
  INV_X1 U5167 ( .A(n8904), .ZN(n5492) );
  NAND2_X1 U5168 ( .A1(n7289), .A2(n5656), .ZN(n5655) );
  AOI21_X1 U5169 ( .B1(P2_REG1_REG_4__SCAN_IN), .B2(n10406), .A(n10398), .ZN(
        n5604) );
  NOR2_X1 U5170 ( .A1(n10477), .A2(n10476), .ZN(n10475) );
  AOI21_X1 U5171 ( .B1(P2_REG1_REG_10__SCAN_IN), .B2(n7207), .A(n7903), .ZN(
        n5620) );
  NAND2_X1 U5172 ( .A1(n8177), .A2(n5625), .ZN(n5626) );
  OR2_X1 U5173 ( .A1(n9057), .A2(n9064), .ZN(n8388) );
  NAND2_X1 U5174 ( .A1(n9061), .A2(n4965), .ZN(n5259) );
  OR2_X1 U5175 ( .A1(n4929), .A2(n9065), .ZN(n6189) );
  NOR2_X1 U5176 ( .A1(n9154), .A2(n8351), .ZN(n5293) );
  AND2_X1 U5177 ( .A1(n5954), .A2(n5955), .ZN(n8325) );
  AOI21_X1 U5178 ( .B1(n8449), .B2(n7766), .A(n5780), .ZN(n8259) );
  AND2_X1 U5179 ( .A1(n5547), .A2(n5269), .ZN(n5268) );
  INV_X1 U5180 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5269) );
  NOR2_X1 U5181 ( .A1(n5542), .A2(n4952), .ZN(n5036) );
  NAND2_X1 U5182 ( .A1(n7469), .A2(n5448), .ZN(n5446) );
  OR2_X1 U5183 ( .A1(n6943), .A2(n7471), .ZN(n5448) );
  NAND2_X1 U5184 ( .A1(n6896), .A2(n6890), .ZN(n6898) );
  NAND3_X1 U5185 ( .A1(n6885), .A2(n6883), .A3(n6882), .ZN(n6896) );
  NOR2_X1 U5186 ( .A1(n9645), .A2(n9660), .ZN(n5365) );
  AOI21_X1 U5187 ( .B1(n9685), .B2(n6679), .A(n4941), .ZN(n5472) );
  AOI21_X1 U5188 ( .B1(n5147), .B2(n5145), .A(n4975), .ZN(n5144) );
  INV_X1 U5189 ( .A(n5465), .ZN(n5145) );
  NOR2_X1 U5190 ( .A1(n6752), .A2(n5326), .ZN(n5325) );
  INV_X1 U5191 ( .A(n8572), .ZN(n5326) );
  NAND2_X1 U5192 ( .A1(n5135), .A2(n5223), .ZN(n5133) );
  OR2_X1 U5193 ( .A1(n7018), .A2(n9763), .ZN(n8721) );
  OR2_X1 U5194 ( .A1(n9784), .A2(n9761), .ZN(n8563) );
  NOR2_X1 U5195 ( .A1(n9784), .A2(n5362), .ZN(n5361) );
  OR2_X1 U5196 ( .A1(n9925), .A2(n9463), .ZN(n8718) );
  NOR2_X1 U5197 ( .A1(n6410), .A2(n5461), .ZN(n5460) );
  AND2_X1 U5198 ( .A1(n8639), .A2(n8659), .ZN(n8632) );
  NAND2_X1 U5199 ( .A1(n8635), .A2(n8599), .ZN(n6882) );
  INV_X1 U5200 ( .A(n7146), .ZN(n6792) );
  NAND2_X1 U5201 ( .A1(n5475), .A2(n6734), .ZN(n6360) );
  NAND2_X1 U5202 ( .A1(n5392), .A2(n5390), .ZN(n6194) );
  AOI21_X1 U5203 ( .B1(n5393), .B2(n5395), .A(n5391), .ZN(n5390) );
  INV_X1 U5204 ( .A(n6176), .ZN(n5391) );
  AND2_X1 U5205 ( .A1(n6176), .A2(n6164), .ZN(n6174) );
  OAI21_X1 U5206 ( .B1(n6119), .B2(n6118), .A(n6117), .ZN(n6127) );
  AND2_X1 U5207 ( .A1(n6138), .A2(n6125), .ZN(n6126) );
  AND2_X1 U5208 ( .A1(n6602), .A2(n6603), .ZN(n6728) );
  INV_X1 U5209 ( .A(SI_18_), .ZN(n6034) );
  OAI211_X1 U5210 ( .C1(n5061), .C2(n5059), .A(n5058), .B(n5233), .ZN(n5910)
         );
  INV_X1 U5211 ( .A(n5234), .ZN(n5233) );
  INV_X1 U5212 ( .A(n5060), .ZN(n5059) );
  AOI21_X1 U5213 ( .B1(n5491), .B2(n5490), .A(n5489), .ZN(n5488) );
  INV_X1 U5214 ( .A(n8905), .ZN(n5489) );
  INV_X1 U5215 ( .A(n8792), .ZN(n5490) );
  NAND2_X1 U5216 ( .A1(n7611), .A2(n5479), .ZN(n5481) );
  NOR2_X1 U5217 ( .A1(n7422), .A2(n5480), .ZN(n5479) );
  INV_X1 U5218 ( .A(n5482), .ZN(n5480) );
  OR2_X1 U5219 ( .A1(n7977), .A2(n8042), .ZN(n5476) );
  NOR2_X1 U5220 ( .A1(n8231), .A2(n5497), .ZN(n5496) );
  INV_X1 U5221 ( .A(n5499), .ZN(n5497) );
  AND4_X1 U5222 ( .A1(n6173), .A2(n6172), .A3(n6171), .A4(n6170), .ZN(n8868)
         );
  AOI21_X1 U5223 ( .B1(P2_REG1_REG_16__SCAN_IN), .B2(n7610), .A(n9007), .ZN(
        n5639) );
  NAND2_X1 U5224 ( .A1(n5575), .A2(n5558), .ZN(n5642) );
  INV_X1 U5225 ( .A(n6874), .ZN(n8797) );
  INV_X1 U5226 ( .A(n4932), .ZN(n8426) );
  AND2_X1 U5227 ( .A1(n9096), .A2(n4958), .ZN(n5245) );
  OR2_X1 U5228 ( .A1(n8779), .A2(n9130), .ZN(n6282) );
  NAND2_X1 U5229 ( .A1(n9112), .A2(n5524), .ZN(n6283) );
  OR2_X1 U5230 ( .A1(n9323), .A2(n8833), .ZN(n5524) );
  NAND2_X1 U5231 ( .A1(n5048), .A2(n5047), .ZN(n6030) );
  NOR2_X1 U5232 ( .A1(n6025), .A2(n9188), .ZN(n5047) );
  AOI21_X1 U5233 ( .B1(n5251), .B2(n5253), .A(n4972), .ZN(n5249) );
  OR2_X1 U5234 ( .A1(n8072), .A2(n6270), .ZN(n5263) );
  OAI21_X1 U5235 ( .B1(n7387), .B2(n5244), .A(n7760), .ZN(n5243) );
  NAND2_X1 U5236 ( .A1(n6317), .A2(n6853), .ZN(n7620) );
  NAND2_X1 U5237 ( .A1(n6300), .A2(n8243), .ZN(n7155) );
  NAND2_X1 U5238 ( .A1(n5084), .A2(n5082), .ZN(n9389) );
  AOI21_X1 U5239 ( .B1(n5085), .B2(n5087), .A(n5083), .ZN(n5082) );
  INV_X1 U5240 ( .A(n7050), .ZN(n5083) );
  NAND2_X1 U5241 ( .A1(n6921), .A2(n6922), .ZN(n6923) );
  NOR2_X1 U5242 ( .A1(n6889), .A2(n8599), .ZN(n6891) );
  NAND2_X1 U5243 ( .A1(n6886), .A2(n6885), .ZN(n6887) );
  NAND2_X1 U5244 ( .A1(n10009), .A2(n10006), .ZN(n6386) );
  NAND2_X1 U5245 ( .A1(n9722), .A2(n8577), .ZN(n9704) );
  NAND2_X1 U5246 ( .A1(n9773), .A2(n8567), .ZN(n9758) );
  AOI21_X1 U5247 ( .B1(n4935), .B2(n6524), .A(n5011), .ZN(n5168) );
  NAND2_X1 U5248 ( .A1(n7793), .A2(n4935), .ZN(n5166) );
  NAND2_X1 U5249 ( .A1(n7797), .A2(n8704), .ZN(n7936) );
  NAND2_X1 U5250 ( .A1(n7141), .A2(n6490), .ZN(n5115) );
  NAND2_X1 U5251 ( .A1(n6397), .A2(n10571), .ZN(n6398) );
  NAND2_X1 U5252 ( .A1(n7122), .A2(n7103), .ZN(n6419) );
  AND2_X1 U5253 ( .A1(n6824), .A2(n4947), .ZN(n6836) );
  NAND2_X1 U5254 ( .A1(n5450), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6776) );
  INV_X1 U5255 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5451) );
  OAI21_X1 U5256 ( .B1(n6014), .B2(n5054), .A(n5052), .ZN(n5057) );
  AOI21_X1 U5257 ( .B1(n5055), .B2(n5053), .A(n5401), .ZN(n5052) );
  XNOR2_X1 U5258 ( .A(n5646), .B(P2_IR_REG_19__SCAN_IN), .ZN(n8479) );
  NAND2_X1 U5259 ( .A1(n5344), .A2(n8387), .ZN(n5343) );
  INV_X1 U5260 ( .A(n8550), .ZN(n5232) );
  NOR2_X1 U5261 ( .A1(n5231), .A2(n6551), .ZN(n5230) );
  NAND2_X1 U5262 ( .A1(n8546), .A2(n4961), .ZN(n5231) );
  OR2_X1 U5263 ( .A1(n5218), .A2(n5219), .ZN(n5214) );
  NAND2_X1 U5264 ( .A1(n5220), .A2(n5222), .ZN(n5215) );
  NOR2_X1 U5265 ( .A1(n5223), .A2(n8626), .ZN(n5219) );
  NAND2_X1 U5266 ( .A1(n6214), .A2(n5388), .ZN(n5387) );
  INV_X1 U5267 ( .A(n6195), .ZN(n5388) );
  INV_X1 U5268 ( .A(SI_9_), .ZN(n10146) );
  NOR2_X1 U5269 ( .A1(n5208), .A2(n9050), .ZN(n5200) );
  NAND2_X1 U5270 ( .A1(n5207), .A2(n5209), .ZN(n5206) );
  INV_X1 U5271 ( .A(n8392), .ZN(n5207) );
  NOR2_X1 U5272 ( .A1(n5844), .A2(n5665), .ZN(n5188) );
  OR4_X1 U5273 ( .A1(n8615), .A2(n8614), .A3(n8613), .A4(n8612), .ZN(n8616) );
  INV_X1 U5274 ( .A(n5394), .ZN(n5393) );
  OAI21_X1 U5275 ( .B1(n6144), .B2(n5395), .A(n6174), .ZN(n5394) );
  AND2_X1 U5276 ( .A1(n5107), .A2(n5106), .ZN(n6325) );
  NOR2_X1 U5277 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n5107) );
  OAI21_X1 U5278 ( .B1(n5945), .B2(n5408), .A(n5944), .ZN(n5407) );
  NAND2_X1 U5279 ( .A1(n5409), .A2(n5926), .ZN(n5408) );
  INV_X1 U5280 ( .A(SI_12_), .ZN(n10048) );
  INV_X1 U5281 ( .A(n8850), .ZN(n5508) );
  OR2_X1 U5282 ( .A1(n9030), .A2(n9033), .ZN(n8444) );
  NOR2_X1 U5283 ( .A1(n5302), .A2(n8383), .ZN(n5297) );
  NAND2_X1 U5284 ( .A1(n5301), .A2(n5300), .ZN(n5299) );
  INV_X1 U5285 ( .A(n5307), .ZN(n5300) );
  NOR2_X1 U5286 ( .A1(n5657), .A2(n5656), .ZN(n5658) );
  NAND2_X1 U5287 ( .A1(n5271), .A2(n5272), .ZN(n5274) );
  AOI21_X1 U5288 ( .B1(n5605), .B2(n5273), .A(n5608), .ZN(n5272) );
  NOR2_X1 U5289 ( .A1(n10469), .A2(n5614), .ZN(n5615) );
  NOR2_X1 U5290 ( .A1(n10473), .A2(n5613), .ZN(n5614) );
  OR2_X1 U5291 ( .A1(n10752), .A2(n10739), .ZN(n8342) );
  OR2_X1 U5292 ( .A1(n10725), .A2(n9237), .ZN(n8330) );
  INV_X1 U5293 ( .A(n5305), .ZN(n5304) );
  OAI22_X1 U5294 ( .A1(n6874), .A2(n5306), .B1(n9045), .B2(n9053), .ZN(n5305)
         );
  NAND2_X1 U5295 ( .A1(n6213), .A2(n8389), .ZN(n5306) );
  NOR2_X1 U5296 ( .A1(n6874), .A2(n5308), .ZN(n5307) );
  INV_X1 U5297 ( .A(n8389), .ZN(n5308) );
  INV_X1 U5298 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5538) );
  INV_X1 U5299 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5534) );
  OR2_X1 U5300 ( .A1(n5606), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n5586) );
  NAND2_X1 U5301 ( .A1(n7040), .A2(n5436), .ZN(n5435) );
  OR2_X1 U5302 ( .A1(n4953), .A2(n5434), .ZN(n5433) );
  INV_X1 U5303 ( .A(n7028), .ZN(n5436) );
  AOI21_X1 U5304 ( .B1(n5431), .B2(n4937), .A(n5089), .ZN(n5088) );
  NAND2_X1 U5305 ( .A1(n5423), .A2(n6981), .ZN(n5422) );
  INV_X1 U5306 ( .A(n5421), .ZN(n5420) );
  OAI21_X1 U5307 ( .B1(n9440), .B2(n5422), .A(n9350), .ZN(n5421) );
  INV_X1 U5308 ( .A(n5418), .ZN(n5417) );
  OAI21_X1 U5309 ( .B1(n9440), .B2(n5419), .A(n9351), .ZN(n5418) );
  NOR2_X1 U5310 ( .A1(n8667), .A2(n8597), .ZN(n5074) );
  AND2_X1 U5311 ( .A1(n9621), .A2(n9498), .ZN(n5224) );
  NAND2_X1 U5312 ( .A1(n5069), .A2(n5226), .ZN(n5225) );
  NOR2_X1 U5313 ( .A1(n8604), .A2(n5227), .ZN(n5226) );
  AND2_X1 U5314 ( .A1(n9621), .A2(n8597), .ZN(n5399) );
  NAND2_X1 U5315 ( .A1(n9616), .A2(n9498), .ZN(n5397) );
  NAND2_X1 U5316 ( .A1(n5125), .A2(n8638), .ZN(n5124) );
  NAND2_X1 U5317 ( .A1(n6625), .A2(n5172), .ZN(n5171) );
  NOR2_X1 U5318 ( .A1(n8605), .A2(n5464), .ZN(n5463) );
  INV_X1 U5319 ( .A(n6613), .ZN(n5172) );
  NAND2_X1 U5320 ( .A1(n6750), .A2(n5131), .ZN(n5130) );
  NOR2_X1 U5321 ( .A1(n6751), .A2(n5132), .ZN(n5131) );
  INV_X1 U5322 ( .A(n8705), .ZN(n5132) );
  NAND2_X1 U5323 ( .A1(n6558), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n6577) );
  OR2_X1 U5324 ( .A1(n9858), .A2(n8203), .ZN(n8700) );
  INV_X1 U5325 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n6482) );
  INV_X1 U5326 ( .A(n6450), .ZN(n5157) );
  OR2_X1 U5327 ( .A1(n7657), .A2(n7959), .ZN(n8525) );
  NAND2_X1 U5328 ( .A1(n7638), .A2(n7678), .ZN(n8510) );
  NAND2_X1 U5329 ( .A1(n7574), .A2(n8612), .ZN(n7573) );
  NAND2_X1 U5330 ( .A1(n8501), .A2(n8514), .ZN(n5149) );
  NAND2_X1 U5331 ( .A1(n5159), .A2(n5158), .ZN(n6725) );
  AOI21_X1 U5332 ( .B1(n5160), .B2(n5163), .A(n4976), .ZN(n5158) );
  AND3_X1 U5333 ( .A1(n4967), .A2(n5475), .A3(n5319), .ZN(n6359) );
  INV_X1 U5334 ( .A(n6360), .ZN(n6356) );
  NOR2_X1 U5335 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n6355) );
  INV_X1 U5336 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n6326) );
  AOI21_X1 U5337 ( .B1(n5402), .B2(n5056), .A(n5016), .ZN(n5400) );
  AND2_X1 U5338 ( .A1(n6086), .A2(n6071), .ZN(n6084) );
  OAI21_X1 U5339 ( .B1(n6014), .B2(n6013), .A(n6000), .ZN(n6032) );
  NOR2_X1 U5340 ( .A1(n5927), .A2(n5411), .ZN(n5410) );
  INV_X1 U5341 ( .A(n5912), .ZN(n5411) );
  OR2_X1 U5342 ( .A1(n6462), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n6508) );
  INV_X1 U5343 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n6324) );
  AND2_X1 U5344 ( .A1(n8441), .A2(n8484), .ZN(n8396) );
  NAND2_X1 U5345 ( .A1(n5889), .A2(n10195), .ZN(n5901) );
  OR2_X1 U5346 ( .A1(n8764), .A2(n8917), .ZN(n8765) );
  NOR2_X1 U5347 ( .A1(n8857), .A2(n5511), .ZN(n5510) );
  INV_X1 U5348 ( .A(n8765), .ZN(n5511) );
  NAND2_X1 U5349 ( .A1(n7420), .A2(n8940), .ZN(n5482) );
  OR2_X1 U5350 ( .A1(n7719), .A2(n7720), .ZN(n5502) );
  NOR2_X1 U5351 ( .A1(n6861), .A2(n6860), .ZN(n7442) );
  INV_X1 U5352 ( .A(n5557), .ZN(n5541) );
  AND4_X1 U5353 ( .A1(n6112), .A2(n6111), .A3(n6110), .A4(n6109), .ZN(n8833)
         );
  NAND2_X1 U5354 ( .A1(n6038), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5782) );
  OAI21_X1 U5355 ( .B1(n5696), .B2(n5598), .A(n5600), .ZN(n7277) );
  NAND2_X1 U5356 ( .A1(n4925), .A2(n5766), .ZN(n5601) );
  NOR2_X1 U5357 ( .A1(n10473), .A2(n10646), .ZN(n5373) );
  XNOR2_X1 U5358 ( .A(n5615), .B(n7881), .ZN(n7877) );
  NAND2_X1 U5359 ( .A1(n5275), .A2(n5623), .ZN(n8177) );
  OAI21_X1 U5360 ( .B1(n8065), .B2(n10701), .A(n5276), .ZN(n5275) );
  XNOR2_X1 U5361 ( .A(n5626), .B(n7314), .ZN(n8954) );
  NOR2_X1 U5362 ( .A1(n8954), .A2(n10715), .ZN(n8953) );
  OR2_X1 U5363 ( .A1(n6219), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n6319) );
  XNOR2_X1 U5364 ( .A(n9052), .B(n9050), .ZN(n5258) );
  NOR2_X1 U5365 ( .A1(n9053), .A2(n10754), .ZN(n5255) );
  OR2_X1 U5366 ( .A1(n9078), .A2(n9090), .ZN(n6284) );
  OR2_X1 U5367 ( .A1(n9314), .A2(n8868), .ZN(n5515) );
  AND4_X1 U5368 ( .A1(n6156), .A2(n6155), .A3(n6154), .A4(n6153), .ZN(n9076)
         );
  AND4_X1 U5369 ( .A1(n6191), .A2(n6190), .A3(n6189), .A4(n6188), .ZN(n9077)
         );
  OR2_X1 U5370 ( .A1(n9096), .A2(n8368), .ZN(n5039) );
  NOR2_X1 U5371 ( .A1(n9105), .A2(n9104), .ZN(n5040) );
  AND4_X1 U5372 ( .A1(n6137), .A2(n6136), .A3(n6135), .A4(n6134), .ZN(n9114)
         );
  AND2_X1 U5373 ( .A1(n6279), .A2(n6083), .ZN(n9154) );
  NAND2_X1 U5374 ( .A1(n9180), .A2(n8342), .ZN(n9164) );
  NAND2_X1 U5375 ( .A1(n6016), .A2(n6015), .ZN(n8848) );
  AND4_X1 U5376 ( .A1(n5953), .A2(n5952), .A3(n5951), .A4(n5950), .ZN(n9235)
         );
  INV_X1 U5377 ( .A(n8325), .ZN(n6271) );
  AND2_X1 U5378 ( .A1(n6271), .A2(n8150), .ZN(n5262) );
  NAND2_X1 U5379 ( .A1(n5263), .A2(n8150), .ZN(n7991) );
  INV_X1 U5380 ( .A(n10686), .ZN(n8073) );
  NAND2_X1 U5381 ( .A1(n5033), .A2(n5035), .ZN(n5030) );
  INV_X1 U5382 ( .A(n5309), .ZN(n5035) );
  NAND2_X1 U5383 ( .A1(n8150), .A2(n7983), .ZN(n8459) );
  AOI21_X1 U5384 ( .B1(n5907), .B2(n8454), .A(n5310), .ZN(n5309) );
  INV_X1 U5385 ( .A(n8314), .ZN(n5310) );
  AND2_X1 U5386 ( .A1(n8316), .A2(n8318), .ZN(n8458) );
  OR2_X1 U5387 ( .A1(n5895), .A2(n8042), .ZN(n8284) );
  INV_X1 U5388 ( .A(n9216), .ZN(n9236) );
  AND2_X1 U5389 ( .A1(n7435), .A2(n8396), .ZN(n9216) );
  OR2_X1 U5390 ( .A1(n5785), .A2(n7108), .ZN(n5317) );
  NAND2_X1 U5391 ( .A1(n6105), .A2(n6104), .ZN(n8779) );
  AND2_X1 U5392 ( .A1(n8396), .A2(n6247), .ZN(n10658) );
  OR3_X1 U5393 ( .A1(n7619), .A2(n8479), .A3(n6243), .ZN(n10683) );
  NOR2_X1 U5394 ( .A1(n10740), .A2(n7432), .ZN(n7430) );
  NAND2_X1 U5395 ( .A1(n8254), .A2(n7948), .ZN(n10740) );
  NAND2_X1 U5396 ( .A1(n7444), .A2(n7228), .ZN(n7432) );
  INV_X1 U5397 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n5741) );
  NAND2_X1 U5398 ( .A1(n5270), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5743) );
  AND2_X1 U5399 ( .A1(n5268), .A2(n5739), .ZN(n5267) );
  NAND2_X1 U5400 ( .A1(n5543), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5550) );
  INV_X1 U5401 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5549) );
  INV_X1 U5402 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n6241) );
  NAND2_X1 U5403 ( .A1(n6946), .A2(n6945), .ZN(n5099) );
  NAND2_X1 U5404 ( .A1(n5446), .A2(n5444), .ZN(n6947) );
  NOR2_X1 U5405 ( .A1(n6945), .A2(n5445), .ZN(n5444) );
  INV_X1 U5406 ( .A(n5447), .ZN(n5445) );
  NAND2_X1 U5407 ( .A1(n6933), .A2(n5518), .ZN(n5427) );
  AOI21_X1 U5408 ( .B1(n5088), .B2(n5432), .A(n5086), .ZN(n5085) );
  INV_X1 U5409 ( .A(n9419), .ZN(n5086) );
  INV_X1 U5410 ( .A(n5088), .ZN(n5087) );
  NAND2_X1 U5411 ( .A1(n6465), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n6483) );
  INV_X1 U5412 ( .A(n6467), .ZN(n6465) );
  INV_X1 U5413 ( .A(n9431), .ZN(n5091) );
  NAND2_X1 U5414 ( .A1(n9381), .A2(n4953), .ZN(n9448) );
  NAND2_X1 U5415 ( .A1(n5430), .A2(n7040), .ZN(n9447) );
  NAND2_X1 U5416 ( .A1(n9381), .A2(n7028), .ZN(n5430) );
  NOR2_X1 U5417 ( .A1(n5080), .A2(n7954), .ZN(n5079) );
  NOR2_X1 U5418 ( .A1(n5080), .A2(n5078), .ZN(n5077) );
  XNOR2_X1 U5419 ( .A(n6907), .B(n6996), .ZN(n6911) );
  INV_X1 U5420 ( .A(n6975), .ZN(n5105) );
  NAND2_X1 U5421 ( .A1(n5420), .A2(n5422), .ZN(n5413) );
  NAND2_X1 U5422 ( .A1(n5417), .A2(n5419), .ZN(n5414) );
  AND2_X1 U5423 ( .A1(n5415), .A2(n5104), .ZN(n5103) );
  OR2_X1 U5424 ( .A1(n8198), .A2(n5105), .ZN(n5104) );
  OR2_X1 U5425 ( .A1(n5417), .A2(n5420), .ZN(n5415) );
  AND2_X1 U5426 ( .A1(n8596), .A2(n8668), .ZN(n8603) );
  INV_X1 U5427 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n6727) );
  NOR4_X1 U5428 ( .A1(n8634), .A2(n8728), .A3(n8664), .A4(n8633), .ZN(n8675)
         );
  OR2_X1 U5429 ( .A1(n6386), .A2(n6343), .ZN(n6344) );
  OR2_X1 U5430 ( .A1(n9684), .A2(n9685), .ZN(n9682) );
  NOR2_X1 U5431 ( .A1(n6678), .A2(n5330), .ZN(n5329) );
  INV_X1 U5432 ( .A(n8648), .ZN(n5330) );
  AOI21_X1 U5433 ( .B1(n5466), .B2(n9747), .A(n4977), .ZN(n5465) );
  NAND2_X1 U5434 ( .A1(n9758), .A2(n5325), .ZN(n8663) );
  OAI21_X1 U5435 ( .B1(n9804), .B2(n5134), .A(n4981), .ZN(n9722) );
  INV_X1 U5436 ( .A(n5135), .ZN(n5134) );
  INV_X1 U5437 ( .A(n5323), .ZN(n5322) );
  NAND2_X1 U5438 ( .A1(n6646), .A2(n6645), .ZN(n9744) );
  NAND2_X1 U5439 ( .A1(n9804), .A2(n8566), .ZN(n9773) );
  NAND2_X1 U5440 ( .A1(n5454), .A2(n5457), .ZN(n8183) );
  INV_X1 U5441 ( .A(n5458), .ZN(n5457) );
  OAI21_X1 U5442 ( .B1(n9834), .B2(n5459), .A(n8626), .ZN(n5458) );
  NAND2_X1 U5443 ( .A1(n8087), .A2(n6566), .ZN(n9835) );
  NAND2_X1 U5444 ( .A1(n9835), .A2(n9834), .ZN(n9833) );
  INV_X1 U5445 ( .A(n9998), .ZN(n5354) );
  NOR2_X1 U5446 ( .A1(n5165), .A2(n8623), .ZN(n5164) );
  INV_X1 U5447 ( .A(n5168), .ZN(n5165) );
  AND2_X1 U5448 ( .A1(n8707), .A2(n8705), .ZN(n8622) );
  NAND2_X1 U5449 ( .A1(n6504), .A2(n6503), .ZN(n7793) );
  NAND2_X1 U5450 ( .A1(n5112), .A2(n5114), .ZN(n5110) );
  NAND2_X1 U5451 ( .A1(n7594), .A2(n7595), .ZN(n7593) );
  OR2_X1 U5452 ( .A1(n7638), .A2(n7678), .ZN(n7645) );
  NAND2_X1 U5453 ( .A1(n7680), .A2(n8613), .ZN(n7679) );
  NAND2_X1 U5454 ( .A1(n5150), .A2(n5460), .ZN(n5152) );
  AOI21_X1 U5455 ( .B1(n5460), .B2(n8608), .A(n4954), .ZN(n5153) );
  INV_X1 U5456 ( .A(n5149), .ZN(n8610) );
  INV_X1 U5457 ( .A(n10543), .ZN(n9764) );
  OR2_X1 U5458 ( .A1(n7122), .A2(n5367), .ZN(n6371) );
  INV_X1 U5459 ( .A(n9515), .ZN(n5367) );
  NAND2_X1 U5460 ( .A1(n6695), .A2(n6694), .ZN(n9660) );
  NAND2_X1 U5461 ( .A1(n6669), .A2(n6668), .ZN(n9695) );
  AND3_X1 U5462 ( .A1(n6395), .A2(n6396), .A3(n5180), .ZN(n10571) );
  OR2_X1 U5463 ( .A1(n7113), .A2(n6419), .ZN(n5180) );
  NAND2_X1 U5464 ( .A1(n6882), .A2(n6755), .ZN(n10546) );
  NAND2_X1 U5465 ( .A1(n6786), .A2(n6780), .ZN(n7146) );
  XNOR2_X1 U5466 ( .A(n6336), .B(n6335), .ZN(n6342) );
  INV_X1 U5467 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n6335) );
  NAND2_X1 U5468 ( .A1(n10001), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6336) );
  XNOR2_X1 U5469 ( .A(n8415), .B(n8414), .ZN(n9338) );
  XNOR2_X1 U5470 ( .A(n6215), .B(n6214), .ZN(n8246) );
  NAND2_X1 U5471 ( .A1(n6160), .A2(n6159), .ZN(n6175) );
  INV_X1 U5472 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n6735) );
  NAND2_X1 U5473 ( .A1(n5403), .A2(n6033), .ZN(n6044) );
  NAND2_X1 U5474 ( .A1(n5051), .A2(n5055), .ZN(n5403) );
  NAND2_X1 U5475 ( .A1(n6014), .A2(n6000), .ZN(n5051) );
  XNOR2_X1 U5476 ( .A(n5995), .B(n5991), .ZN(n7402) );
  XNOR2_X1 U5477 ( .A(n5928), .B(n5927), .ZN(n7219) );
  NAND2_X1 U5478 ( .A1(n5412), .A2(n5912), .ZN(n5928) );
  NAND2_X1 U5479 ( .A1(n5238), .A2(n5334), .ZN(n5896) );
  NAND2_X1 U5480 ( .A1(n5852), .A2(n5236), .ZN(n5238) );
  XNOR2_X1 U5481 ( .A(n5883), .B(n5882), .ZN(n7141) );
  NAND2_X1 U5482 ( .A1(n5333), .A2(n5866), .ZN(n5883) );
  NAND2_X1 U5483 ( .A1(n6129), .A2(n6128), .ZN(n9273) );
  AND2_X1 U5484 ( .A1(n7418), .A2(n7614), .ZN(n7419) );
  AOI21_X1 U5485 ( .B1(n5486), .B2(n5485), .A(n5014), .ZN(n5484) );
  INV_X1 U5486 ( .A(n10741), .ZN(n8862) );
  AND2_X1 U5487 ( .A1(n7920), .A2(n8031), .ZN(n7921) );
  INV_X1 U5488 ( .A(n8031), .ZN(n10620) );
  AOI21_X1 U5489 ( .B1(n8830), .B2(n8831), .A(n5527), .ZN(n8885) );
  INV_X1 U5490 ( .A(n8868), .ZN(n9090) );
  INV_X1 U5491 ( .A(n9076), .ZN(n9102) );
  INV_X1 U5492 ( .A(n9114), .ZN(n9089) );
  INV_X1 U5493 ( .A(n10755), .ZN(n8931) );
  INV_X1 U5494 ( .A(n8035), .ZN(n10657) );
  INV_X1 U5495 ( .A(n7628), .ZN(n8942) );
  OR2_X1 U5496 ( .A1(n10502), .A2(n10501), .ZN(n10513) );
  NOR2_X1 U5497 ( .A1(n10505), .A2(n10504), .ZN(n10503) );
  AND2_X1 U5498 ( .A1(n5686), .A2(n5370), .ZN(n5369) );
  NAND2_X1 U5499 ( .A1(n5726), .A2(n5683), .ZN(n5370) );
  NOR2_X1 U5500 ( .A1(n10499), .A2(n5645), .ZN(n5647) );
  OAI21_X1 U5501 ( .B1(n4950), .B2(n7872), .A(n5734), .ZN(n5735) );
  OAI21_X1 U5502 ( .B1(n9049), .B2(n6213), .A(n8389), .ZN(n6877) );
  INV_X1 U5503 ( .A(n9328), .ZN(n9138) );
  INV_X1 U5504 ( .A(n9230), .ZN(n10639) );
  INV_X1 U5505 ( .A(n9222), .ZN(n10638) );
  NOR2_X1 U5506 ( .A1(n6294), .A2(n10684), .ZN(n6847) );
  NAND2_X1 U5507 ( .A1(n5765), .A2(n5045), .ZN(n5044) );
  OAI21_X1 U5508 ( .B1(n7106), .B2(n5046), .A(n4943), .ZN(n5045) );
  NAND2_X1 U5509 ( .A1(n6302), .A2(n6301), .ZN(n7135) );
  OR2_X1 U5510 ( .A1(n7155), .A2(P2_D_REG_1__SCAN_IN), .ZN(n6302) );
  AND2_X1 U5511 ( .A1(n8226), .A2(n8112), .ZN(n6785) );
  OAI21_X1 U5512 ( .B1(n7073), .B2(n7074), .A(n7075), .ZN(n7081) );
  XNOR2_X1 U5513 ( .A(n6921), .B(n6920), .ZN(n7249) );
  NAND2_X1 U5514 ( .A1(n6618), .A2(n6617), .ZN(n9784) );
  INV_X1 U5515 ( .A(n9706), .ZN(n9743) );
  NAND2_X1 U5516 ( .A1(n6576), .A2(n6575), .ZN(n9830) );
  INV_X1 U5517 ( .A(n9491), .ZN(n9451) );
  INV_X1 U5518 ( .A(n9494), .ZN(n9480) );
  AND2_X1 U5519 ( .A1(n5067), .A2(n4926), .ZN(n5064) );
  INV_X1 U5520 ( .A(n9640), .ZN(n9499) );
  AND2_X1 U5521 ( .A1(n6831), .A2(n6830), .ZN(n6832) );
  AOI21_X1 U5522 ( .B1(n6822), .B2(n10546), .A(n6821), .ZN(n6838) );
  INV_X1 U5523 ( .A(n6820), .ZN(n6821) );
  XNOR2_X1 U5524 ( .A(n6815), .B(n6814), .ZN(n6822) );
  AOI22_X1 U5525 ( .A1(n9499), .A2(n9821), .B1(n9615), .B2(n9498), .ZN(n6820)
         );
  NAND2_X1 U5526 ( .A1(n6481), .A2(n6480), .ZN(n7961) );
  INV_X1 U5527 ( .A(n5140), .ZN(n6839) );
  NAND2_X1 U5528 ( .A1(n6529), .A2(n6528), .ZN(n9846) );
  OR2_X1 U5529 ( .A1(n5332), .A2(n5179), .ZN(n6797) );
  OAI21_X1 U5530 ( .B1(n9629), .B2(n9937), .A(n9625), .ZN(n5332) );
  INV_X1 U5531 ( .A(n9634), .ZN(n5179) );
  INV_X1 U5532 ( .A(n8290), .ZN(n8311) );
  NOR2_X1 U5533 ( .A1(n8681), .A2(n8686), .ZN(n8500) );
  AOI21_X1 U5534 ( .B1(n8334), .B2(n8333), .A(n9203), .ZN(n5340) );
  INV_X1 U5535 ( .A(n8553), .ZN(n5228) );
  OAI211_X1 U5536 ( .C1(n5232), .C2(n4983), .A(n8547), .B(n5230), .ZN(n5229)
         );
  NAND2_X1 U5537 ( .A1(n4984), .A2(n9738), .ZN(n5222) );
  AOI21_X1 U5538 ( .B1(n4973), .B2(n9738), .A(n5221), .ZN(n5220) );
  OAI21_X1 U5539 ( .B1(n5003), .B2(n8568), .A(n8597), .ZN(n5221) );
  NOR2_X1 U5540 ( .A1(n5217), .A2(n5220), .ZN(n5216) );
  INV_X1 U5541 ( .A(n5218), .ZN(n5217) );
  NOR2_X1 U5542 ( .A1(n8497), .A2(n8496), .ZN(n8681) );
  NAND2_X1 U5543 ( .A1(n8394), .A2(n8393), .ZN(n5350) );
  NAND2_X1 U5544 ( .A1(n8390), .A2(n8391), .ZN(n5209) );
  INV_X1 U5545 ( .A(SI_22_), .ZN(n10121) );
  INV_X1 U5546 ( .A(SI_14_), .ZN(n10139) );
  INV_X1 U5547 ( .A(n5410), .ZN(n5409) );
  INV_X1 U5548 ( .A(n8435), .ZN(n5202) );
  INV_X1 U5549 ( .A(n5209), .ZN(n5208) );
  INV_X1 U5550 ( .A(n10443), .ZN(n5273) );
  INV_X1 U5551 ( .A(n9450), .ZN(n5434) );
  INV_X1 U5552 ( .A(n8590), .ZN(n5227) );
  AOI21_X1 U5553 ( .B1(n5144), .B2(n5146), .A(n5142), .ZN(n5141) );
  INV_X1 U5554 ( .A(n6679), .ZN(n5142) );
  INV_X1 U5555 ( .A(n8642), .ZN(n5324) );
  INV_X1 U5556 ( .A(n6626), .ZN(n5464) );
  NAND2_X1 U5557 ( .A1(n7494), .A2(n9510), .ZN(n8514) );
  AND2_X1 U5558 ( .A1(n5468), .A2(n5161), .ZN(n5160) );
  NAND2_X1 U5559 ( .A1(n8630), .A2(n5162), .ZN(n5161) );
  AND2_X1 U5560 ( .A1(n5125), .A2(n6705), .ZN(n5468) );
  INV_X1 U5561 ( .A(n6692), .ZN(n5162) );
  OAI21_X1 U5562 ( .B1(n6196), .B2(n5386), .A(n5385), .ZN(n8399) );
  NAND2_X1 U5563 ( .A1(n6214), .A2(n4945), .ZN(n5386) );
  NAND2_X1 U5564 ( .A1(n5021), .A2(n4945), .ZN(n5385) );
  INV_X1 U5565 ( .A(n6159), .ZN(n5395) );
  INV_X1 U5566 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n6068) );
  INV_X1 U5567 ( .A(SI_17_), .ZN(n10133) );
  INV_X1 U5568 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n5996) );
  INV_X1 U5569 ( .A(SI_15_), .ZN(n10042) );
  INV_X1 U5570 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n5963) );
  AND2_X1 U5571 ( .A1(n5236), .A2(n5517), .ZN(n5060) );
  OAI21_X1 U5572 ( .B1(n5334), .B2(n5235), .A(n5897), .ZN(n5234) );
  NAND2_X1 U5573 ( .A1(n5337), .A2(n5866), .ZN(n5336) );
  INV_X1 U5574 ( .A(n5882), .ZN(n5337) );
  OR3_X1 U5575 ( .A1(n10751), .A2(n8396), .A3(n5522), .ZN(n7423) );
  AOI21_X1 U5576 ( .B1(n5205), .B2(n5203), .A(n5201), .ZN(n5348) );
  NOR2_X1 U5577 ( .A1(n5208), .A2(n5204), .ZN(n5203) );
  NOR2_X1 U5578 ( .A1(n4936), .A2(n5202), .ZN(n5201) );
  NAND2_X1 U5579 ( .A1(n9051), .A2(n8435), .ZN(n5204) );
  NOR2_X1 U5580 ( .A1(n8438), .A2(n8387), .ZN(n5346) );
  OR2_X1 U5581 ( .A1(n7269), .A2(n5654), .ZN(n7290) );
  NOR2_X1 U5582 ( .A1(n5810), .A2(n5661), .ZN(n5662) );
  INV_X1 U5583 ( .A(n5187), .ZN(n5666) );
  NOR2_X1 U5584 ( .A1(n8970), .A2(n5632), .ZN(n5633) );
  NOR2_X1 U5585 ( .A1(n8997), .A2(n5371), .ZN(n5680) );
  NOR2_X1 U5586 ( .A1(n9012), .A2(n6017), .ZN(n5371) );
  NAND2_X1 U5587 ( .A1(n6114), .A2(n5294), .ZN(n5291) );
  INV_X1 U5588 ( .A(n5526), .ZN(n5290) );
  INV_X1 U5589 ( .A(n5293), .ZN(n5292) );
  OR2_X1 U5590 ( .A1(n9138), .A2(n8930), .ZN(n8355) );
  INV_X1 U5591 ( .A(n8252), .ZN(n5294) );
  INV_X1 U5592 ( .A(n5252), .ZN(n5251) );
  OAI21_X1 U5593 ( .B1(n9213), .B2(n5253), .A(n9203), .ZN(n5252) );
  INV_X1 U5594 ( .A(n5984), .ZN(n5985) );
  AND2_X1 U5595 ( .A1(n5034), .A2(n8458), .ZN(n5033) );
  NAND2_X1 U5596 ( .A1(n5309), .A2(n8309), .ZN(n5034) );
  INV_X1 U5597 ( .A(n5542), .ZN(n5314) );
  INV_X1 U5598 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5552) );
  INV_X1 U5599 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5584) );
  INV_X1 U5600 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5532) );
  NAND2_X1 U5601 ( .A1(n7471), .A2(n6943), .ZN(n5447) );
  NAND2_X1 U5602 ( .A1(n5443), .A2(n5442), .ZN(n5441) );
  INV_X1 U5603 ( .A(n9460), .ZN(n5442) );
  INV_X1 U5604 ( .A(n9459), .ZN(n5443) );
  INV_X1 U5605 ( .A(n8141), .ZN(n5080) );
  OR4_X1 U5606 ( .A1(n8626), .A2(n9834), .A3(n8625), .A4(n8624), .ZN(n8627) );
  OR2_X1 U5607 ( .A1(n9628), .A2(n9499), .ZN(n8639) );
  NOR2_X1 U5608 ( .A1(n5120), .A2(n8630), .ZN(n5117) );
  INV_X1 U5609 ( .A(n5121), .ZN(n5120) );
  NOR2_X1 U5610 ( .A1(n6812), .A2(n5122), .ZN(n5121) );
  INV_X1 U5611 ( .A(n5124), .ZN(n5122) );
  NAND2_X1 U5612 ( .A1(n9628), .A2(n5365), .ZN(n5364) );
  INV_X1 U5613 ( .A(n5147), .ZN(n5146) );
  NOR2_X1 U5614 ( .A1(n5324), .A2(n5136), .ZN(n5135) );
  OAI21_X1 U5615 ( .B1(n5325), .B2(n5324), .A(n9724), .ZN(n5323) );
  INV_X1 U5616 ( .A(n9780), .ZN(n5072) );
  INV_X1 U5617 ( .A(n6585), .ZN(n5459) );
  NOR2_X1 U5618 ( .A1(n5459), .A2(n5456), .ZN(n5455) );
  INV_X1 U5619 ( .A(n6566), .ZN(n5456) );
  INV_X1 U5620 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n8120) );
  OR2_X1 U5621 ( .A1(n9830), .A2(n6584), .ZN(n8716) );
  NAND2_X1 U5622 ( .A1(n6543), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n6560) );
  INV_X1 U5623 ( .A(n9943), .ZN(n5355) );
  INV_X1 U5624 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n6530) );
  OR2_X1 U5625 ( .A1(n6531), .A2(n6530), .ZN(n6545) );
  NOR2_X1 U5626 ( .A1(n8542), .A2(n9846), .ZN(n5356) );
  INV_X1 U5627 ( .A(n5113), .ZN(n5112) );
  OAI21_X1 U5628 ( .B1(n7595), .B2(n5114), .A(n8700), .ZN(n5113) );
  OR2_X1 U5629 ( .A1(n8520), .A2(n6746), .ZN(n8698) );
  INV_X1 U5630 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n6454) );
  AND2_X1 U5631 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n6411) );
  AND2_X1 U5632 ( .A1(n6742), .A2(n8684), .ZN(n7369) );
  NAND2_X1 U5633 ( .A1(n7369), .A2(n8607), .ZN(n7368) );
  NAND2_X1 U5634 ( .A1(n8635), .A2(n8739), .ZN(n8671) );
  INV_X1 U5635 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n10195) );
  NAND2_X1 U5636 ( .A1(n5176), .A2(n6325), .ZN(n6599) );
  INV_X1 U5637 ( .A(n10001), .ZN(n6338) );
  XNOR2_X1 U5638 ( .A(n8399), .B(n8400), .ZN(n8397) );
  AND2_X1 U5639 ( .A1(n6195), .A2(n6182), .ZN(n6193) );
  AND2_X1 U5640 ( .A1(n6159), .A2(n6143), .ZN(n6144) );
  AND4_X1 U5641 ( .A1(n5175), .A2(n6735), .A3(n5470), .A4(n6381), .ZN(n5174)
         );
  INV_X1 U5642 ( .A(n6000), .ZN(n5053) );
  INV_X1 U5643 ( .A(n5055), .ZN(n5054) );
  AOI21_X1 U5644 ( .B1(n6013), .B2(n6000), .A(n5056), .ZN(n5055) );
  NAND2_X1 U5645 ( .A1(n4980), .A2(n5908), .ZN(n5404) );
  INV_X1 U5646 ( .A(n5407), .ZN(n5406) );
  NAND2_X1 U5647 ( .A1(n5062), .A2(n5061), .ZN(n5852) );
  NAND2_X1 U5648 ( .A1(n5840), .A2(n5843), .ZN(n5062) );
  NOR2_X1 U5649 ( .A1(n5336), .A2(n5237), .ZN(n5236) );
  INV_X1 U5650 ( .A(n5851), .ZN(n5237) );
  INV_X1 U5651 ( .A(n5335), .ZN(n5334) );
  OAI21_X1 U5652 ( .B1(n5336), .B2(n5863), .A(n5881), .ZN(n5335) );
  NAND2_X1 U5653 ( .A1(n5852), .A2(n5851), .ZN(n5864) );
  OAI21_X1 U5654 ( .B1(n7103), .B2(n5792), .A(n5791), .ZN(n5806) );
  NAND2_X1 U5655 ( .A1(n7103), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n5791) );
  INV_X1 U5656 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n5751) );
  OR2_X1 U5657 ( .A1(n8229), .A2(n9235), .ZN(n5499) );
  INV_X1 U5658 ( .A(n8806), .ZN(n5487) );
  NOR2_X1 U5659 ( .A1(n5985), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6019) );
  INV_X1 U5660 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n10090) );
  NAND2_X1 U5661 ( .A1(n10090), .A2(n6019), .ZN(n6018) );
  INV_X1 U5662 ( .A(n8266), .ZN(n7481) );
  AOI21_X1 U5663 ( .B1(n5510), .B2(n5508), .A(n4969), .ZN(n5507) );
  INV_X1 U5664 ( .A(n5510), .ZN(n5509) );
  NOR2_X1 U5665 ( .A1(n6018), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n6037) );
  NAND2_X1 U5666 ( .A1(n8894), .A2(n6037), .ZN(n6054) );
  OR2_X1 U5667 ( .A1(n5833), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5855) );
  AND3_X1 U5668 ( .A1(n7406), .A2(n7135), .A3(n6864), .ZN(n7450) );
  OR2_X1 U5669 ( .A1(n8387), .A2(n6297), .ZN(n7433) );
  AND2_X1 U5670 ( .A1(n8437), .A2(n5299), .ZN(n5298) );
  AND2_X1 U5671 ( .A1(n8444), .A2(n5530), .ZN(n8437) );
  AND4_X1 U5672 ( .A1(n8431), .A2(n8430), .A3(n8429), .A4(n8428), .ZN(n9033)
         );
  OR2_X1 U5673 ( .A1(n7277), .A2(n5599), .ZN(n7278) );
  AND2_X1 U5674 ( .A1(n7294), .A2(n7295), .ZN(n7297) );
  OAI21_X1 U5675 ( .B1(n10420), .B2(n5374), .A(n5189), .ZN(n10433) );
  NAND2_X1 U5676 ( .A1(n5375), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5374) );
  NAND2_X1 U5677 ( .A1(n5664), .A2(n5375), .ZN(n5189) );
  INV_X1 U5678 ( .A(n10434), .ZN(n5375) );
  NOR2_X1 U5679 ( .A1(n10420), .A2(n10421), .ZN(n10419) );
  NOR2_X1 U5680 ( .A1(n5610), .A2(n10450), .ZN(n10471) );
  OR2_X1 U5681 ( .A1(n5586), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n5611) );
  OAI21_X1 U5682 ( .B1(n7877), .B2(n5281), .A(n5280), .ZN(n7903) );
  NAND2_X1 U5683 ( .A1(n5282), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5281) );
  NAND2_X1 U5684 ( .A1(n5616), .A2(n5282), .ZN(n5280) );
  NOR2_X1 U5685 ( .A1(n7877), .A2(n10665), .ZN(n7876) );
  INV_X1 U5686 ( .A(n5372), .ZN(n5668) );
  NAND2_X1 U5687 ( .A1(n8164), .A2(n5674), .ZN(n5675) );
  NOR2_X1 U5688 ( .A1(n8953), .A2(n5628), .ZN(n8972) );
  NOR2_X1 U5689 ( .A1(n8972), .A2(n8971), .ZN(n8970) );
  OAI21_X1 U5690 ( .B1(n8990), .B2(n5284), .A(n5283), .ZN(n9007) );
  NAND2_X1 U5691 ( .A1(n5285), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n5284) );
  NAND2_X1 U5692 ( .A1(n5634), .A2(n5285), .ZN(n5283) );
  INV_X1 U5693 ( .A(n9008), .ZN(n5285) );
  NOR2_X1 U5694 ( .A1(n8990), .A2(n10729), .ZN(n8989) );
  NOR2_X1 U5695 ( .A1(n9018), .A2(n9192), .ZN(n9017) );
  INV_X1 U5696 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n8894) );
  OAI21_X1 U5697 ( .B1(n9016), .B2(n5278), .A(n5277), .ZN(n10499) );
  NAND2_X1 U5698 ( .A1(n5279), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n5278) );
  NAND2_X1 U5699 ( .A1(n5640), .A2(n5279), .ZN(n5277) );
  NAND2_X1 U5700 ( .A1(n8465), .A2(n6158), .ZN(n5038) );
  NAND2_X1 U5701 ( .A1(n5039), .A2(n6158), .ZN(n5037) );
  NAND2_X1 U5702 ( .A1(n9126), .A2(n6281), .ZN(n9127) );
  NOR2_X1 U5703 ( .A1(n6090), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n6106) );
  NAND2_X1 U5704 ( .A1(n10203), .A2(n6076), .ZN(n6090) );
  NAND2_X1 U5705 ( .A1(n8350), .A2(n8349), .ZN(n9159) );
  INV_X1 U5706 ( .A(n9181), .ZN(n9173) );
  NAND2_X1 U5707 ( .A1(n9242), .A2(n5977), .ZN(n9210) );
  INV_X1 U5708 ( .A(n5971), .ZN(n5972) );
  NOR2_X1 U5709 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(n5972), .ZN(n5984) );
  AND2_X1 U5710 ( .A1(n6272), .A2(n8326), .ZN(n9232) );
  AOI21_X1 U5711 ( .B1(n5262), .B2(n6270), .A(n4964), .ZN(n5261) );
  INV_X1 U5712 ( .A(n9232), .ZN(n9243) );
  NAND2_X1 U5713 ( .A1(n5933), .A2(n5932), .ZN(n5949) );
  NOR2_X1 U5714 ( .A1(n5855), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5873) );
  AND2_X1 U5715 ( .A1(n8282), .A2(n8301), .ZN(n5315) );
  AND3_X1 U5716 ( .A1(n5813), .A2(n5812), .A3(n5811), .ZN(n7413) );
  INV_X1 U5717 ( .A(n8255), .ZN(n5050) );
  NAND2_X1 U5718 ( .A1(n6248), .A2(n7387), .ZN(n5242) );
  CLKBUF_X1 U5719 ( .A(n7760), .Z(n7768) );
  OR2_X1 U5720 ( .A1(n8396), .A2(n6296), .ZN(n6850) );
  NAND2_X1 U5721 ( .A1(n8422), .A2(n8421), .ZN(n9030) );
  NAND2_X1 U5722 ( .A1(n5303), .A2(n5304), .ZN(n8439) );
  NAND2_X1 U5723 ( .A1(n9049), .A2(n5307), .ZN(n5303) );
  INV_X1 U5724 ( .A(n9135), .ZN(n9284) );
  AND4_X1 U5725 ( .A1(n6042), .A2(n6041), .A3(n6040), .A4(n6039), .ZN(n10739)
         );
  NAND2_X1 U5726 ( .A1(n5983), .A2(n5982), .ZN(n10725) );
  AND3_X1 U5727 ( .A1(n5829), .A2(n5828), .A3(n5827), .ZN(n10600) );
  INV_X1 U5728 ( .A(n10658), .ZN(n10754) );
  XNOR2_X1 U5729 ( .A(n5551), .B(n5552), .ZN(n7443) );
  XNOR2_X1 U5730 ( .A(n5548), .B(n5547), .ZN(n6303) );
  NOR2_X1 U5731 ( .A1(n9371), .A2(n5438), .ZN(n5437) );
  INV_X1 U5732 ( .A(n5440), .ZN(n5438) );
  NAND2_X1 U5733 ( .A1(n9459), .A2(n9460), .ZN(n5440) );
  NAND2_X1 U5734 ( .A1(n9458), .A2(n5441), .ZN(n5439) );
  OR2_X1 U5735 ( .A1(n6577), .A2(n8120), .ZN(n6592) );
  AND2_X1 U5736 ( .A1(n7050), .A2(n7049), .ZN(n9419) );
  OR2_X1 U5737 ( .A1(n6455), .A2(n6454), .ZN(n6467) );
  NAND2_X1 U5738 ( .A1(n6619), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n6630) );
  OR2_X1 U5739 ( .A1(n6630), .A2(n9433), .ZN(n6638) );
  AOI21_X1 U5740 ( .B1(n5437), .B2(n5095), .A(n5094), .ZN(n5093) );
  INV_X1 U5741 ( .A(n7010), .ZN(n5094) );
  INV_X1 U5742 ( .A(n5441), .ZN(n5095) );
  INV_X1 U5743 ( .A(n5437), .ZN(n5096) );
  INV_X1 U5744 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n9433) );
  NAND2_X1 U5745 ( .A1(n6650), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n6661) );
  NAND2_X1 U5746 ( .A1(n6494), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n6517) );
  NAND2_X1 U5747 ( .A1(n6590), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n6609) );
  INV_X1 U5748 ( .A(n6592), .ZN(n6590) );
  NAND2_X1 U5749 ( .A1(n5427), .A2(n5424), .ZN(n5425) );
  NAND2_X1 U5750 ( .A1(n5398), .A2(n5397), .ZN(n5396) );
  AOI21_X1 U5751 ( .B1(n8595), .B2(n9955), .A(n4986), .ZN(n5075) );
  AOI21_X1 U5752 ( .B1(n8595), .B2(n5224), .A(n5074), .ZN(n5073) );
  NAND2_X1 U5753 ( .A1(n5116), .A2(n5118), .ZN(n6815) );
  AOI21_X1 U5754 ( .B1(n5121), .B2(n5127), .A(n5119), .ZN(n5118) );
  NAND2_X1 U5755 ( .A1(n9654), .A2(n5117), .ZN(n5116) );
  INV_X1 U5756 ( .A(n8639), .ZN(n5119) );
  NAND2_X1 U5757 ( .A1(n5123), .A2(n5124), .ZN(n6813) );
  NAND2_X1 U5758 ( .A1(n9653), .A2(n5126), .ZN(n5123) );
  INV_X1 U5759 ( .A(n8632), .ZN(n6812) );
  NOR2_X1 U5760 ( .A1(n9675), .A2(n5363), .ZN(n9644) );
  INV_X1 U5761 ( .A(n5365), .ZN(n5363) );
  AND2_X1 U5762 ( .A1(n6720), .A2(n6828), .ZN(n9626) );
  NAND2_X1 U5763 ( .A1(n9654), .A2(n5163), .ZN(n9653) );
  NAND2_X1 U5764 ( .A1(n9688), .A2(n8645), .ZN(n9669) );
  OR2_X1 U5765 ( .A1(n6670), .A2(n9424), .ZN(n6684) );
  NAND2_X1 U5766 ( .A1(n6754), .A2(n8648), .ZN(n9686) );
  AND2_X1 U5767 ( .A1(n8578), .A2(n8648), .ZN(n9703) );
  NOR2_X1 U5768 ( .A1(n5359), .A2(n7018), .ZN(n5357) );
  NAND2_X1 U5769 ( .A1(n5170), .A2(n5169), .ZN(n9746) );
  AOI21_X1 U5770 ( .B1(n4938), .B2(n5173), .A(n5012), .ZN(n5169) );
  NAND2_X1 U5771 ( .A1(n8563), .A2(n8567), .ZN(n9780) );
  NAND2_X1 U5772 ( .A1(n9794), .A2(n5361), .ZN(n9782) );
  NAND2_X1 U5773 ( .A1(n9794), .A2(n9989), .ZN(n9795) );
  AND2_X1 U5774 ( .A1(n6612), .A2(n6611), .ZN(n9412) );
  NAND2_X1 U5775 ( .A1(n5130), .A2(n8708), .ZN(n8080) );
  NOR2_X1 U5776 ( .A1(n8625), .A2(n5129), .ZN(n5128) );
  INV_X1 U5777 ( .A(n8708), .ZN(n5129) );
  NAND2_X1 U5778 ( .A1(n7801), .A2(n4939), .ZN(n8088) );
  NAND2_X1 U5779 ( .A1(n7801), .A2(n7838), .ZN(n7934) );
  AND2_X1 U5780 ( .A1(n8701), .A2(n8704), .ZN(n8621) );
  AND2_X1 U5781 ( .A1(n7739), .A2(n8149), .ZN(n7801) );
  NOR2_X1 U5782 ( .A1(n7599), .A2(n7961), .ZN(n7739) );
  AOI21_X1 U5783 ( .B1(n8614), .B2(n5157), .A(n4974), .ZN(n5156) );
  AND2_X1 U5784 ( .A1(n7681), .A2(n7734), .ZN(n7682) );
  NAND2_X1 U5785 ( .A1(n7682), .A2(n10630), .ZN(n7654) );
  NOR2_X1 U5786 ( .A1(n7581), .A2(n10609), .ZN(n7681) );
  OR2_X1 U5787 ( .A1(n7544), .A2(n7491), .ZN(n7581) );
  NAND2_X1 U5788 ( .A1(n7545), .A2(n10593), .ZN(n7544) );
  OAI211_X1 U5789 ( .C1(n8608), .C2(n8496), .A(n5328), .B(n8609), .ZN(n7540)
         );
  AND2_X1 U5790 ( .A1(n6743), .A2(n8495), .ZN(n5327) );
  NOR2_X1 U5791 ( .A1(n10536), .A2(n7523), .ZN(n7545) );
  NAND2_X1 U5792 ( .A1(n8497), .A2(n8608), .ZN(n7538) );
  NAND2_X1 U5793 ( .A1(n5025), .A2(n10538), .ZN(n10536) );
  NAND2_X1 U5794 ( .A1(n8683), .A2(n6743), .ZN(n10540) );
  INV_X1 U5795 ( .A(n7369), .ZN(n6741) );
  NAND2_X1 U5796 ( .A1(n6707), .A2(n6706), .ZN(n9645) );
  NAND2_X1 U5797 ( .A1(n6660), .A2(n6659), .ZN(n9711) );
  NAND2_X1 U5798 ( .A1(n5167), .A2(n6523), .ZN(n7933) );
  OR2_X1 U5799 ( .A1(n7793), .A2(n6524), .ZN(n5167) );
  NAND2_X1 U5800 ( .A1(n7593), .A2(n8529), .ZN(n7741) );
  OR2_X1 U5801 ( .A1(n6883), .A2(n6793), .ZN(n10669) );
  AOI21_X1 U5802 ( .B1(n6792), .B2(n10278), .A(n6784), .ZN(n7078) );
  NOR2_X1 U5803 ( .A1(n6420), .A2(n5320), .ZN(n5318) );
  NAND2_X1 U5804 ( .A1(n5474), .A2(n5321), .ZN(n5320) );
  INV_X1 U5805 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5474) );
  NAND2_X1 U5806 ( .A1(n6340), .A2(n6339), .ZN(n6341) );
  OR3_X1 U5807 ( .A1(n6359), .A2(n6334), .A3(n6509), .ZN(n6340) );
  NOR2_X1 U5808 ( .A1(n6338), .A2(n6337), .ZN(n6339) );
  NOR2_X1 U5809 ( .A1(P1_IR_REG_29__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n6337) );
  XNOR2_X1 U5810 ( .A(n8397), .B(SI_29_), .ZN(n6802) );
  XNOR2_X1 U5811 ( .A(n6216), .B(n6230), .ZN(n9343) );
  NAND2_X1 U5812 ( .A1(n6215), .A2(n6214), .ZN(n6233) );
  NAND2_X1 U5813 ( .A1(n6354), .A2(n6353), .ZN(n6358) );
  NOR2_X1 U5814 ( .A1(n6331), .A2(n6509), .ZN(n6353) );
  XNOR2_X1 U5815 ( .A(n6736), .B(n6735), .ZN(n8598) );
  INV_X1 U5816 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n6732) );
  NAND2_X1 U5817 ( .A1(n6731), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6733) );
  NAND2_X1 U5818 ( .A1(n5405), .A2(n5926), .ZN(n5946) );
  NAND2_X1 U5819 ( .A1(n5412), .A2(n5410), .ZN(n5405) );
  INV_X1 U5820 ( .A(n6729), .ZN(n6462) );
  OAI21_X1 U5821 ( .B1(n5840), .B2(n5839), .A(n5843), .ZN(n5849) );
  NAND2_X1 U5822 ( .A1(n5502), .A2(n4934), .ZN(n7848) );
  INV_X1 U5823 ( .A(n5494), .ZN(n8761) );
  NAND2_X1 U5824 ( .A1(n8228), .A2(n5499), .ZN(n8230) );
  AND2_X1 U5825 ( .A1(n6319), .A2(n6220), .ZN(n9041) );
  AOI21_X1 U5826 ( .B1(n4934), .B2(n7720), .A(n4982), .ZN(n5500) );
  AND4_X1 U5827 ( .A1(n5989), .A2(n5988), .A3(n5987), .A4(n5986), .ZN(n9237)
         );
  NAND2_X1 U5828 ( .A1(n8851), .A2(n8850), .ZN(n8849) );
  NAND2_X1 U5829 ( .A1(n8849), .A2(n8765), .ZN(n8856) );
  NAND2_X1 U5830 ( .A1(n6148), .A2(n6147), .ZN(n9093) );
  NAND2_X1 U5831 ( .A1(n8820), .A2(n8773), .ZN(n8876) );
  AOI21_X1 U5832 ( .B1(n8154), .B2(n8153), .A(n8152), .ZN(n8156) );
  AND4_X1 U5833 ( .A1(n6094), .A2(n6093), .A3(n6092), .A4(n6091), .ZN(n9148)
         );
  INV_X1 U5834 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n10205) );
  AND2_X1 U5835 ( .A1(n6206), .A2(n6187), .ZN(n9065) );
  NAND2_X1 U5836 ( .A1(n7431), .A2(n10638), .ZN(n8910) );
  AND4_X1 U5837 ( .A1(n6024), .A2(n6023), .A3(n6022), .A4(n6021), .ZN(n8917)
         );
  OR2_X1 U5838 ( .A1(n7436), .A2(n7435), .ZN(n8918) );
  NAND2_X1 U5839 ( .A1(n5494), .A2(n5493), .ZN(n8915) );
  NOR2_X1 U5840 ( .A1(n5498), .A2(n8760), .ZN(n5493) );
  INV_X1 U5841 ( .A(n8916), .ZN(n5498) );
  INV_X1 U5842 ( .A(n8912), .ZN(n8914) );
  AND2_X1 U5843 ( .A1(n7434), .A2(n7435), .ZN(n8922) );
  XNOR2_X1 U5844 ( .A(n5564), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8484) );
  NOR2_X1 U5845 ( .A1(n5542), .A2(n5505), .ZN(n5503) );
  INV_X1 U5846 ( .A(n8917), .ZN(n9217) );
  INV_X1 U5847 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n7223) );
  INV_X1 U5848 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n7210) );
  AND4_X1 U5849 ( .A1(n5894), .A2(n5893), .A3(n5892), .A4(n5891), .ZN(n8042)
         );
  INV_X1 U5850 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n7208) );
  AND4_X1 U5851 ( .A1(n5878), .A2(n5877), .A3(n5876), .A4(n5875), .ZN(n8031)
         );
  NAND2_X1 U5852 ( .A1(n6038), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5800) );
  NAND2_X1 U5853 ( .A1(n4930), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5781) );
  INV_X1 U5854 ( .A(P2_U3893), .ZN(n10508) );
  NOR2_X1 U5855 ( .A1(n10444), .A2(n10443), .ZN(n10442) );
  NOR2_X1 U5856 ( .A1(n10415), .A2(n5605), .ZN(n10444) );
  XNOR2_X1 U5857 ( .A(n5675), .B(n7314), .ZN(n8945) );
  AND2_X1 U5858 ( .A1(n5675), .A2(n7314), .ZN(n5676) );
  NOR2_X1 U5859 ( .A1(n8945), .A2(n8944), .ZN(n8943) );
  OAI21_X1 U5860 ( .B1(n8945), .B2(n5377), .A(n5376), .ZN(n8961) );
  NAND2_X1 U5861 ( .A1(n5378), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n5377) );
  NAND2_X1 U5862 ( .A1(n5676), .A2(n5378), .ZN(n5376) );
  INV_X1 U5863 ( .A(n8962), .ZN(n5378) );
  NOR2_X1 U5864 ( .A1(n8981), .A2(n8980), .ZN(n8979) );
  OAI21_X1 U5865 ( .B1(n8981), .B2(n5191), .A(n5190), .ZN(n8997) );
  NAND2_X1 U5866 ( .A1(n5192), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n5191) );
  NAND2_X1 U5867 ( .A1(n5679), .A2(n5192), .ZN(n5190) );
  INV_X1 U5868 ( .A(n8998), .ZN(n5192) );
  INV_X1 U5869 ( .A(n10507), .ZN(n10474) );
  OAI22_X1 U5870 ( .A1(n6876), .A2(n9234), .B1(n9064), .B2(n9236), .ZN(n9039)
         );
  NOR2_X1 U5871 ( .A1(n5256), .A2(n5255), .ZN(n5254) );
  NAND2_X1 U5872 ( .A1(n5258), .A2(n9211), .ZN(n5257) );
  NOR2_X1 U5873 ( .A1(n9077), .A2(n9236), .ZN(n5256) );
  NAND2_X1 U5874 ( .A1(n6204), .A2(n6203), .ZN(n9057) );
  NAND2_X1 U5875 ( .A1(n6184), .A2(n6183), .ZN(n9260) );
  NAND2_X1 U5876 ( .A1(n6166), .A2(n6165), .ZN(n9078) );
  AND2_X1 U5877 ( .A1(n6168), .A2(n6151), .ZN(n9094) );
  NOR2_X1 U5878 ( .A1(n5040), .A2(n5039), .ZN(n9098) );
  AND2_X1 U5879 ( .A1(n5246), .A2(n4958), .ZN(n9088) );
  NAND2_X1 U5880 ( .A1(n6283), .A2(n6282), .ZN(n9101) );
  AND2_X1 U5881 ( .A1(n9115), .A2(n9134), .ZN(n9135) );
  NAND2_X1 U5882 ( .A1(n9162), .A2(n8350), .ZN(n9155) );
  NAND2_X1 U5883 ( .A1(n6053), .A2(n6052), .ZN(n9296) );
  AND3_X1 U5884 ( .A1(n6062), .A2(n6061), .A3(n6060), .ZN(n10755) );
  NAND2_X1 U5885 ( .A1(n6030), .A2(n6029), .ZN(n9182) );
  NAND2_X1 U5886 ( .A1(n6036), .A2(n6035), .ZN(n10752) );
  INV_X1 U5887 ( .A(n10739), .ZN(n9194) );
  AND2_X1 U5888 ( .A1(n6007), .A2(n6006), .ZN(n10741) );
  OR2_X1 U5889 ( .A1(n10740), .A2(n6318), .ZN(n9240) );
  NAND2_X1 U5890 ( .A1(n5263), .A2(n5262), .ZN(n7993) );
  NAND2_X1 U5891 ( .A1(n8029), .A2(n5907), .ZN(n5032) );
  AND4_X1 U5892 ( .A1(n5925), .A2(n5924), .A3(n5923), .A4(n5922), .ZN(n10686)
         );
  AND4_X1 U5893 ( .A1(n5906), .A2(n5905), .A3(n5904), .A4(n5903), .ZN(n8035)
         );
  NAND2_X1 U5894 ( .A1(n5888), .A2(n5887), .ZN(n5895) );
  INV_X1 U5895 ( .A(n10641), .ZN(n9225) );
  NAND2_X1 U5896 ( .A1(n5756), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5767) );
  NAND2_X1 U5897 ( .A1(n10643), .A2(n7695), .ZN(n9230) );
  NAND2_X1 U5898 ( .A1(n5756), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5746) );
  NAND2_X1 U5899 ( .A1(n10761), .A2(n10751), .ZN(n9288) );
  INV_X1 U5900 ( .A(n9030), .ZN(n9302) );
  AND2_X1 U5901 ( .A1(n8412), .A2(n8411), .ZN(n9305) );
  INV_X1 U5902 ( .A(n8779), .ZN(n9323) );
  AND2_X1 U5903 ( .A1(n6089), .A2(n6088), .ZN(n9328) );
  NAND2_X1 U5904 ( .A1(n6074), .A2(n6073), .ZN(n9331) );
  NAND2_X1 U5905 ( .A1(n7141), .A2(n5981), .ZN(n5210) );
  INV_X1 U5906 ( .A(n7432), .ZN(n7428) );
  AND2_X1 U5907 ( .A1(n7443), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7228) );
  AND2_X1 U5908 ( .A1(n5739), .A2(n5742), .ZN(n5477) );
  INV_X1 U5909 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5545) );
  NAND2_X1 U5910 ( .A1(n5544), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5546) );
  INV_X1 U5911 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7946) );
  INV_X1 U5912 ( .A(n8484), .ZN(n7948) );
  INV_X1 U5913 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5562) );
  INV_X1 U5914 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7865) );
  INV_X1 U5915 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7831) );
  INV_X1 U5916 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n7335) );
  AND2_X1 U5917 ( .A1(n4946), .A2(n5537), .ZN(n5618) );
  INV_X1 U5918 ( .A(n7908), .ZN(n7207) );
  INV_X1 U5919 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n7200) );
  NAND2_X1 U5920 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n5596) );
  NAND2_X1 U5921 ( .A1(n5617), .A2(n5594), .ZN(n5595) );
  NAND3_X1 U5922 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_IR_REG_0__SCAN_IN), .ZN(n5186) );
  NAND2_X1 U5923 ( .A1(n5264), .A2(n5185), .ZN(n5184) );
  AND2_X1 U5924 ( .A1(n7124), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7101) );
  NAND2_X1 U5925 ( .A1(n9448), .A2(n9450), .ZN(n9363) );
  NAND2_X1 U5926 ( .A1(n6958), .A2(n6960), .ZN(n7953) );
  NAND2_X1 U5927 ( .A1(n5439), .A2(n5440), .ZN(n9370) );
  INV_X1 U5928 ( .A(n9508), .ZN(n7826) );
  INV_X1 U5929 ( .A(n5098), .ZN(n5097) );
  NOR2_X1 U5930 ( .A1(n6996), .A2(n8606), .ZN(n6897) );
  NOR2_X1 U5931 ( .A1(n5428), .A2(n5426), .ZN(n7378) );
  INV_X1 U5932 ( .A(n6930), .ZN(n5428) );
  INV_X1 U5933 ( .A(n5427), .ZN(n5426) );
  NAND2_X1 U5934 ( .A1(n6589), .A2(n6588), .ZN(n9925) );
  OAI21_X1 U5935 ( .B1(n9381), .B2(n5087), .A(n5085), .ZN(n9421) );
  NAND2_X1 U5936 ( .A1(n8197), .A2(n8198), .ZN(n5102) );
  NAND2_X1 U5937 ( .A1(n6649), .A2(n6648), .ZN(n9721) );
  OR2_X1 U5938 ( .A1(n7092), .A2(n7087), .ZN(n9434) );
  NAND2_X1 U5939 ( .A1(n7951), .A2(n6960), .ZN(n8139) );
  NAND2_X1 U5940 ( .A1(n9388), .A2(n7062), .ZN(n9471) );
  INV_X1 U5941 ( .A(n9496), .ZN(n9472) );
  OR2_X1 U5942 ( .A1(n7092), .A2(n7088), .ZN(n9491) );
  AOI21_X1 U5943 ( .B1(n5103), .B2(n5105), .A(n4985), .ZN(n5101) );
  NAND2_X1 U5944 ( .A1(n7086), .A2(n9854), .ZN(n9494) );
  AND2_X1 U5945 ( .A1(n8602), .A2(n5240), .ZN(n8601) );
  NAND2_X1 U5946 ( .A1(n8603), .A2(n8597), .ZN(n5240) );
  OR2_X1 U5947 ( .A1(n8733), .A2(n5068), .ZN(n5067) );
  INV_X1 U5948 ( .A(n8740), .ZN(n5068) );
  NAND2_X1 U5949 ( .A1(n8679), .A2(n8740), .ZN(n5063) );
  NAND2_X1 U5950 ( .A1(n6712), .A2(n6711), .ZN(n9656) );
  NAND2_X1 U5951 ( .A1(n6691), .A2(n6690), .ZN(n9689) );
  NAND4_X1 U5952 ( .A1(n6404), .A2(n6403), .A3(n6402), .A4(n6401), .ZN(n9511)
         );
  CLKBUF_X1 U5953 ( .A(n6902), .Z(n10542) );
  NOR2_X1 U5954 ( .A1(n9614), .A2(n9797), .ZN(n9865) );
  NAND2_X1 U5955 ( .A1(n5469), .A2(n6705), .ZN(n9635) );
  NAND2_X1 U5956 ( .A1(n9652), .A2(n8630), .ZN(n5469) );
  NAND2_X1 U5957 ( .A1(n6681), .A2(n6680), .ZN(n9883) );
  NAND2_X1 U5958 ( .A1(n9682), .A2(n6679), .ZN(n9668) );
  NAND2_X1 U5959 ( .A1(n8663), .A2(n8642), .ZN(n9723) );
  NAND2_X1 U5961 ( .A1(n9744), .A2(n5466), .ZN(n9730) );
  NAND2_X1 U5962 ( .A1(n9758), .A2(n8572), .ZN(n9739) );
  NAND2_X1 U5963 ( .A1(n6627), .A2(n6626), .ZN(n9756) );
  NAND2_X1 U5964 ( .A1(n9781), .A2(n6625), .ZN(n6627) );
  NAND2_X1 U5965 ( .A1(n9833), .A2(n6585), .ZN(n8184) );
  NAND2_X1 U5966 ( .A1(n5166), .A2(n5168), .ZN(n7968) );
  NAND2_X1 U5967 ( .A1(n6750), .A2(n8705), .ZN(n7964) );
  NAND2_X1 U5968 ( .A1(n6464), .A2(n6463), .ZN(n7657) );
  NAND2_X1 U5969 ( .A1(n7633), .A2(n8614), .ZN(n7632) );
  NAND2_X1 U5970 ( .A1(n7679), .A2(n6450), .ZN(n7633) );
  NAND2_X1 U5971 ( .A1(n5153), .A2(n5152), .ZN(n7392) );
  AND2_X1 U5972 ( .A1(n7588), .A2(n6811), .ZN(n9836) );
  NAND2_X1 U5973 ( .A1(n5462), .A2(n6398), .ZN(n7536) );
  AND2_X1 U5974 ( .A1(n10524), .A2(n6826), .ZN(n10552) );
  INV_X1 U5975 ( .A(n9836), .ZN(n10559) );
  INV_X1 U5976 ( .A(n10552), .ZN(n9802) );
  INV_X1 U5977 ( .A(n9854), .ZN(n10554) );
  NAND2_X1 U5978 ( .A1(n5239), .A2(n6493), .ZN(n9858) );
  NAND2_X1 U5979 ( .A1(n7219), .A2(n6490), .ZN(n5239) );
  NAND2_X1 U5980 ( .A1(n10681), .A2(n10675), .ZN(n5473) );
  NOR2_X1 U5981 ( .A1(n6801), .A2(n5516), .ZN(n6805) );
  NAND2_X1 U5982 ( .A1(n6838), .A2(n6837), .ZN(n5140) );
  INV_X1 U5983 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n5178) );
  INV_X1 U5984 ( .A(n9660), .ZN(n9963) );
  INV_X1 U5985 ( .A(n9695), .ZN(n9968) );
  INV_X1 U5986 ( .A(n9711), .ZN(n9972) );
  INV_X1 U5987 ( .A(n9721), .ZN(n9976) );
  INV_X1 U5988 ( .A(n9830), .ZN(n9994) );
  NAND2_X1 U5989 ( .A1(n6557), .A2(n6556), .ZN(n9998) );
  INV_X1 U5990 ( .A(n6341), .ZN(n10009) );
  NAND2_X1 U5991 ( .A1(n6774), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6775) );
  XNOR2_X1 U5992 ( .A(n6778), .B(P1_IR_REG_24__SCAN_IN), .ZN(n8112) );
  AND2_X1 U5993 ( .A1(n6735), .A2(n5452), .ZN(n5449) );
  INV_X1 U5994 ( .A(n8598), .ZN(n8739) );
  NAND2_X1 U5995 ( .A1(n6614), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6615) );
  AND2_X1 U5996 ( .A1(n6540), .A2(n6553), .ZN(n10324) );
  AND2_X1 U5997 ( .A1(n6527), .A2(n6537), .ZN(n10375) );
  AND2_X1 U5998 ( .A1(n6514), .A2(n6526), .ZN(n8124) );
  AND2_X1 U5999 ( .A1(n6479), .A2(n6491), .ZN(n10389) );
  NOR2_X1 U6000 ( .A1(n7103), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10003) );
  OAI21_X1 U6001 ( .B1(n10503), .B2(n4940), .A(n5686), .ZN(n5193) );
  OAI211_X1 U6002 ( .C1(n10503), .C2(n5027), .A(n5369), .B(n5368), .ZN(n5737)
         );
  NOR2_X1 U6003 ( .A1(n6870), .A2(n5531), .ZN(n6871) );
  NAND2_X1 U6004 ( .A1(n5041), .A2(n4944), .ZN(P2_U3455) );
  NAND2_X1 U6005 ( .A1(n5042), .A2(n10764), .ZN(n5041) );
  NAND2_X1 U6006 ( .A1(n10676), .A2(n6723), .ZN(n5331) );
  NAND2_X1 U6007 ( .A1(n5139), .A2(n5137), .ZN(P1_U3519) );
  INV_X1 U6008 ( .A(n5138), .ZN(n5137) );
  NAND2_X1 U6009 ( .A1(n5140), .A2(n10681), .ZN(n5139) );
  OAI21_X1 U6010 ( .B1(n6840), .B2(n5473), .A(n6842), .ZN(n5138) );
  NAND2_X1 U6011 ( .A1(n10678), .A2(n5178), .ZN(n5177) );
  NAND2_X1 U6012 ( .A1(n6786), .A2(n6785), .ZN(n6890) );
  NAND2_X2 U6013 ( .A1(n5648), .A2(n4927), .ZN(n5765) );
  AND2_X1 U6014 ( .A1(n4948), .A2(n7751), .ZN(n4934) );
  AND2_X1 U6015 ( .A1(n5295), .A2(n5294), .ZN(n9115) );
  INV_X1 U6016 ( .A(n5491), .ZN(n5485) );
  OAI211_X1 U6017 ( .C1(n6419), .C2(n7108), .A(n6383), .B(n6382), .ZN(n10553)
         );
  INV_X1 U6018 ( .A(n10553), .ZN(n10538) );
  AND2_X1 U6019 ( .A1(n6523), .A2(n4968), .ZN(n4935) );
  AND2_X1 U6020 ( .A1(n8576), .A2(n8577), .ZN(n9724) );
  AND2_X1 U6021 ( .A1(n4987), .A2(n5206), .ZN(n4936) );
  NOR2_X1 U6022 ( .A1(n7040), .A2(n9450), .ZN(n4937) );
  AND2_X1 U6023 ( .A1(n5463), .A2(n5171), .ZN(n4938) );
  AND2_X1 U6024 ( .A1(n5356), .A2(n5355), .ZN(n4939) );
  INV_X1 U6025 ( .A(n6599), .ZN(n5319) );
  NAND2_X1 U6026 ( .A1(n8594), .A2(n8593), .ZN(n9621) );
  INV_X1 U6027 ( .A(n9621), .ZN(n9955) );
  AND2_X1 U6028 ( .A1(n10505), .A2(n10504), .ZN(n4940) );
  INV_X1 U6029 ( .A(n9747), .ZN(n6645) );
  AND2_X1 U6030 ( .A1(n8721), .A2(n8573), .ZN(n9747) );
  INV_X1 U6031 ( .A(n5467), .ZN(n5466) );
  NAND2_X1 U6032 ( .A1(n9731), .A2(n6647), .ZN(n5467) );
  INV_X1 U6033 ( .A(n7018), .ZN(n9980) );
  NAND2_X1 U6034 ( .A1(n6635), .A2(n6634), .ZN(n7018) );
  NOR2_X1 U6035 ( .A1(n9883), .A2(n9689), .ZN(n4941) );
  AND2_X1 U6036 ( .A1(n9309), .A2(n9064), .ZN(n4942) );
  INV_X1 U6037 ( .A(n5302), .ZN(n5301) );
  NAND2_X1 U6038 ( .A1(n5304), .A2(n8395), .ZN(n5302) );
  NAND2_X1 U6039 ( .A1(n7103), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n4943) );
  INV_X1 U6040 ( .A(n5506), .ZN(n5505) );
  NAND2_X1 U6041 ( .A1(n5097), .A2(n6947), .ZN(n7820) );
  AND2_X1 U6042 ( .A1(n6881), .A2(n5019), .ZN(n4944) );
  INV_X1 U6043 ( .A(n6031), .ZN(n5056) );
  INV_X1 U6044 ( .A(n8599), .ZN(n6888) );
  XNOR2_X1 U6045 ( .A(n6737), .B(P1_IR_REG_20__SCAN_IN), .ZN(n8599) );
  OR2_X1 U6046 ( .A1(n6231), .A2(n6230), .ZN(n4945) );
  INV_X1 U6047 ( .A(n5857), .ZN(n6038) );
  AND2_X1 U6048 ( .A1(n5312), .A2(n5533), .ZN(n4946) );
  OR3_X1 U6049 ( .A1(n9675), .A2(n5364), .A3(n6823), .ZN(n4947) );
  AND2_X1 U6050 ( .A1(n5754), .A2(n5044), .ZN(n7414) );
  NAND2_X1 U6051 ( .A1(n7748), .A2(n8937), .ZN(n4948) );
  INV_X1 U6052 ( .A(n5398), .ZN(n8634) );
  OR2_X1 U6053 ( .A1(n8596), .A2(n8668), .ZN(n5398) );
  NAND2_X1 U6054 ( .A1(n5533), .A2(n5532), .ZN(n5583) );
  AND4_X1 U6055 ( .A1(n6347), .A2(n6346), .A3(n6345), .A4(n6344), .ZN(n6895)
         );
  XOR2_X1 U6056 ( .A(n6927), .B(n8745), .Z(n4949) );
  INV_X1 U6057 ( .A(n5810), .ZN(n10406) );
  INV_X1 U6058 ( .A(n8529), .ZN(n5114) );
  XNOR2_X1 U6059 ( .A(n5896), .B(n5517), .ZN(n6461) );
  OAI21_X1 U6060 ( .B1(n9381), .B2(n4937), .A(n5431), .ZN(n9361) );
  NOR2_X1 U6061 ( .A1(n5521), .A2(n5492), .ZN(n5491) );
  INV_X1 U6062 ( .A(n9351), .ZN(n5423) );
  XOR2_X1 U6063 ( .A(n5728), .B(n5727), .Z(n4950) );
  AND4_X1 U6064 ( .A1(n6328), .A2(n6327), .A3(n6603), .A4(n6326), .ZN(n4951)
         );
  OR3_X1 U6065 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .A3(
        P2_IR_REG_23__SCAN_IN), .ZN(n4952) );
  AND2_X1 U6066 ( .A1(n7039), .A2(n7028), .ZN(n4953) );
  XNOR2_X1 U6067 ( .A(n5773), .B(n10066), .ZN(n5772) );
  NAND2_X1 U6068 ( .A1(n5389), .A2(n6086), .ZN(n6095) );
  NOR2_X1 U6069 ( .A1(n6451), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n6729) );
  NAND2_X1 U6070 ( .A1(n5109), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6737) );
  AND2_X1 U6071 ( .A1(n9511), .A2(n7547), .ZN(n4954) );
  NAND2_X1 U6072 ( .A1(n6898), .A2(n8743), .ZN(n6915) );
  INV_X1 U6073 ( .A(n8596), .ZN(n9951) );
  NAND2_X1 U6074 ( .A1(n6516), .A2(n6515), .ZN(n8542) );
  OR2_X1 U6075 ( .A1(n10708), .A2(n10696), .ZN(n4955) );
  AND2_X1 U6076 ( .A1(n5439), .A2(n5437), .ZN(n4956) );
  AND2_X1 U6077 ( .A1(n9744), .A2(n6647), .ZN(n4957) );
  NAND2_X1 U6078 ( .A1(n9273), .A2(n9089), .ZN(n4958) );
  OR2_X1 U6079 ( .A1(n9675), .A2(n5364), .ZN(n4959) );
  AND2_X1 U6080 ( .A1(n9173), .A2(n6029), .ZN(n4960) );
  AND4_X1 U6081 ( .A1(n5861), .A2(n5860), .A3(n5859), .A4(n5858), .ZN(n7750)
         );
  NAND2_X1 U6082 ( .A1(n6381), .A2(n5470), .ZN(n6406) );
  AND2_X1 U6083 ( .A1(n5311), .A2(n5036), .ZN(n5568) );
  INV_X1 U6084 ( .A(n5568), .ZN(n5567) );
  OR2_X1 U6085 ( .A1(n8548), .A2(n8549), .ZN(n4961) );
  NOR2_X1 U6086 ( .A1(n8979), .A2(n5679), .ZN(n4962) );
  NOR2_X1 U6087 ( .A1(n8989), .A2(n5634), .ZN(n4963) );
  AND2_X1 U6088 ( .A1(n10714), .A2(n8934), .ZN(n4964) );
  INV_X1 U6089 ( .A(n5432), .ZN(n5431) );
  OR2_X1 U6090 ( .A1(n8382), .A2(n9077), .ZN(n4965) );
  AND2_X1 U6091 ( .A1(n8395), .A2(n8435), .ZN(n4966) );
  AND2_X1 U6092 ( .A1(n5318), .A2(n4951), .ZN(n4967) );
  NAND2_X1 U6093 ( .A1(n9846), .A2(n9502), .ZN(n4968) );
  AND2_X1 U6094 ( .A1(n8767), .A2(n9201), .ZN(n4969) );
  AND2_X1 U6095 ( .A1(n8632), .A2(n8589), .ZN(n4970) );
  INV_X1 U6096 ( .A(n5127), .ZN(n5126) );
  NAND2_X1 U6097 ( .A1(n8638), .A2(n8654), .ZN(n5127) );
  INV_X1 U6098 ( .A(n5366), .ZN(n9659) );
  NOR2_X1 U6099 ( .A1(n9675), .A2(n9660), .ZN(n5366) );
  AND2_X1 U6100 ( .A1(n8388), .A2(n8389), .ZN(n9051) );
  INV_X1 U6101 ( .A(n9051), .ZN(n9050) );
  AND2_X1 U6102 ( .A1(n9106), .A2(n9114), .ZN(n4971) );
  INV_X1 U6103 ( .A(n5223), .ZN(n8566) );
  NAND2_X1 U6104 ( .A1(n5072), .A2(n9771), .ZN(n5223) );
  AND2_X1 U6105 ( .A1(n8848), .A2(n9217), .ZN(n4972) );
  NOR2_X1 U6106 ( .A1(n8562), .A2(n5514), .ZN(n4973) );
  NOR2_X1 U6107 ( .A1(n7638), .A2(n9507), .ZN(n4974) );
  NOR2_X1 U6108 ( .A1(n9711), .A2(n9726), .ZN(n4975) );
  NOR2_X1 U6109 ( .A1(n9645), .A2(n9656), .ZN(n4976) );
  NOR2_X1 U6110 ( .A1(n9721), .A2(n9706), .ZN(n4977) );
  AND2_X1 U6111 ( .A1(n8708), .A2(n8711), .ZN(n8623) );
  INV_X1 U6112 ( .A(n9685), .ZN(n6678) );
  AND2_X1 U6113 ( .A1(n8645), .A2(n8649), .ZN(n9685) );
  INV_X1 U6114 ( .A(n5359), .ZN(n5358) );
  NAND2_X1 U6115 ( .A1(n5361), .A2(n5360), .ZN(n5359) );
  AND2_X1 U6116 ( .A1(n8572), .A2(n9738), .ZN(n8605) );
  NAND2_X1 U6117 ( .A1(n6542), .A2(n6541), .ZN(n9943) );
  AND3_X1 U6118 ( .A1(n5175), .A2(n5470), .A3(n6381), .ZN(n6424) );
  AND2_X1 U6119 ( .A1(n8638), .A2(n8658), .ZN(n9636) );
  INV_X1 U6120 ( .A(n9636), .ZN(n5125) );
  AND2_X1 U6121 ( .A1(n5215), .A2(n5214), .ZN(n4978) );
  NAND2_X1 U6122 ( .A1(n9057), .A2(n9259), .ZN(n4979) );
  XNOR2_X1 U6123 ( .A(n6918), .B(n8745), .ZN(n6921) );
  AND2_X1 U6124 ( .A1(n5942), .A2(n5926), .ZN(n4980) );
  AND2_X1 U6125 ( .A1(n5322), .A2(n5133), .ZN(n4981) );
  INV_X1 U6126 ( .A(n8465), .ZN(n9104) );
  AND2_X1 U6127 ( .A1(n7847), .A2(n7750), .ZN(n4982) );
  NAND4_X1 U6128 ( .A1(n8705), .A2(n8597), .A3(n8704), .A4(n8530), .ZN(n4983)
         );
  NOR2_X1 U6129 ( .A1(n8562), .A2(n8626), .ZN(n4984) );
  NAND2_X1 U6130 ( .A1(n5092), .A2(n5090), .ZN(n9377) );
  NAND2_X1 U6131 ( .A1(n5414), .A2(n5413), .ZN(n4985) );
  NAND2_X1 U6132 ( .A1(n8942), .A2(n7414), .ZN(n8256) );
  OR2_X1 U6133 ( .A1(n8603), .A2(n5399), .ZN(n4986) );
  AND2_X1 U6134 ( .A1(n4966), .A2(n5350), .ZN(n4987) );
  INV_X1 U6135 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n5264) );
  OR2_X1 U6136 ( .A1(n9296), .A2(n10755), .ZN(n8350) );
  AND3_X1 U6137 ( .A1(n6735), .A2(n5452), .A3(n5451), .ZN(n4988) );
  INV_X1 U6138 ( .A(n10453), .ZN(n7145) );
  AND2_X1 U6139 ( .A1(n5588), .A2(n5611), .ZN(n10453) );
  OR2_X1 U6140 ( .A1(n5765), .A2(n4925), .ZN(n4989) );
  AND2_X1 U6141 ( .A1(n9711), .A2(n9726), .ZN(n4990) );
  NOR2_X1 U6142 ( .A1(n9140), .A2(n6280), .ZN(n4991) );
  OR2_X1 U6143 ( .A1(n5040), .A2(n8368), .ZN(n4992) );
  NOR2_X1 U6144 ( .A1(n9015), .A2(n5640), .ZN(n4993) );
  NOR2_X1 U6145 ( .A1(n5526), .A2(n5292), .ZN(n4994) );
  INV_X1 U6146 ( .A(n5517), .ZN(n5235) );
  NAND2_X1 U6147 ( .A1(n9162), .A2(n5293), .ZN(n5295) );
  AND2_X1 U6148 ( .A1(n5311), .A2(n5314), .ZN(n4995) );
  AND2_X1 U6149 ( .A1(n8360), .A2(n8359), .ZN(n4996) );
  AND2_X1 U6150 ( .A1(n8774), .A2(n8773), .ZN(n4997) );
  AND2_X1 U6151 ( .A1(n4939), .A2(n5354), .ZN(n4998) );
  NAND2_X1 U6152 ( .A1(n8002), .A2(n7503), .ZN(n4999) );
  OR2_X1 U6153 ( .A1(n8346), .A2(n9159), .ZN(n5000) );
  OR2_X1 U6154 ( .A1(n8353), .A2(n9154), .ZN(n5001) );
  INV_X1 U6155 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5321) );
  AND2_X1 U6156 ( .A1(n5488), .A2(n5487), .ZN(n5486) );
  NAND2_X1 U6157 ( .A1(n6957), .A2(n6956), .ZN(n6960) );
  NAND2_X1 U6158 ( .A1(n8228), .A2(n5496), .ZN(n5494) );
  INV_X1 U6159 ( .A(n6956), .ZN(n5078) );
  XNOR2_X1 U6160 ( .A(n6733), .B(n6732), .ZN(n6889) );
  INV_X1 U6161 ( .A(n10473), .ZN(n7154) );
  OR2_X1 U6162 ( .A1(n8029), .A2(n8454), .ZN(n8027) );
  NAND2_X1 U6163 ( .A1(n6030), .A2(n4960), .ZN(n9180) );
  OAI21_X1 U6164 ( .B1(n9210), .B2(n5990), .A(n8330), .ZN(n9187) );
  INV_X1 U6165 ( .A(n9187), .ZN(n5048) );
  NAND2_X1 U6166 ( .A1(n9784), .A2(n9761), .ZN(n8567) );
  INV_X1 U6167 ( .A(n8567), .ZN(n5136) );
  INV_X1 U6168 ( .A(n7881), .ZN(n7202) );
  AND2_X1 U6169 ( .A1(n9794), .A2(n5358), .ZN(n5002) );
  OAI21_X1 U6170 ( .B1(n8098), .B2(n7982), .A(n7981), .ZN(n8154) );
  NAND2_X1 U6171 ( .A1(n9212), .A2(n6274), .ZN(n9199) );
  NAND2_X1 U6172 ( .A1(n7002), .A2(n7001), .ZN(n9458) );
  NAND2_X1 U6173 ( .A1(n5416), .A2(n6981), .ZN(n9349) );
  NAND2_X1 U6174 ( .A1(n5102), .A2(n6975), .ZN(n9439) );
  NAND2_X1 U6175 ( .A1(n6304), .A2(n7226), .ZN(n7406) );
  INV_X1 U6176 ( .A(n9418), .ZN(n5089) );
  AND2_X1 U6177 ( .A1(n8572), .A2(n8563), .ZN(n5003) );
  AND2_X1 U6178 ( .A1(n8565), .A2(n8564), .ZN(n5004) );
  NOR2_X1 U6179 ( .A1(n8943), .A2(n5676), .ZN(n5005) );
  NOR2_X1 U6180 ( .A1(n9040), .A2(n10754), .ZN(n5006) );
  AND2_X1 U6181 ( .A1(n6960), .A2(n6959), .ZN(n5007) );
  AND2_X1 U6182 ( .A1(n8849), .A2(n5510), .ZN(n5008) );
  NOR2_X1 U6183 ( .A1(n8064), .A2(n5621), .ZN(n5009) );
  NAND2_X1 U6184 ( .A1(n6218), .A2(n6217), .ZN(n9045) );
  NAND2_X1 U6185 ( .A1(n6958), .A2(n5007), .ZN(n7951) );
  AND2_X1 U6186 ( .A1(n5494), .A2(n5495), .ZN(n5010) );
  NOR2_X1 U6187 ( .A1(n9846), .A2(n9502), .ZN(n5011) );
  NOR2_X1 U6188 ( .A1(n9909), .A2(n9777), .ZN(n5012) );
  NAND2_X1 U6189 ( .A1(n5166), .A2(n5164), .ZN(n7966) );
  NAND2_X1 U6190 ( .A1(n6729), .A2(n6602), .ZN(n5013) );
  NOR2_X1 U6191 ( .A1(n8795), .A2(n9064), .ZN(n5014) );
  INV_X1 U6192 ( .A(n8760), .ZN(n5495) );
  NAND2_X1 U6193 ( .A1(n4946), .A2(n5503), .ZN(n5015) );
  NAND2_X1 U6194 ( .A1(n6065), .A2(n6064), .ZN(n5016) );
  AND2_X1 U6195 ( .A1(n6096), .A2(n6086), .ZN(n5017) );
  AND2_X1 U6196 ( .A1(n6715), .A2(n6714), .ZN(n9628) );
  AND2_X1 U6197 ( .A1(n6043), .A2(n6033), .ZN(n5402) );
  INV_X1 U6198 ( .A(n5402), .ZN(n5401) );
  NAND2_X1 U6199 ( .A1(n6629), .A2(n6628), .ZN(n9909) );
  INV_X1 U6200 ( .A(n9909), .ZN(n5360) );
  NAND2_X1 U6201 ( .A1(n6889), .A2(n8598), .ZN(n6883) );
  NAND2_X1 U6202 ( .A1(n7801), .A2(n5356), .ZN(n5018) );
  OR2_X1 U6203 ( .A1(n10764), .A2(n6879), .ZN(n5019) );
  XNOR2_X1 U6204 ( .A(n6775), .B(P1_IR_REG_26__SCAN_IN), .ZN(n6786) );
  NAND2_X1 U6205 ( .A1(n5032), .A2(n5309), .ZN(n8020) );
  AND2_X1 U6206 ( .A1(n6607), .A2(n6606), .ZN(n9989) );
  INV_X1 U6207 ( .A(n9989), .ZN(n5362) );
  NAND2_X1 U6208 ( .A1(n5098), .A2(n6947), .ZN(n7854) );
  NAND2_X1 U6209 ( .A1(n5847), .A2(n8301), .ZN(n7891) );
  NOR2_X1 U6210 ( .A1(n7876), .A2(n5616), .ZN(n5020) );
  AND2_X1 U6211 ( .A1(n6228), .A2(n6202), .ZN(n6214) );
  NAND2_X1 U6212 ( .A1(n5387), .A2(n6232), .ZN(n5021) );
  NAND2_X1 U6213 ( .A1(n7306), .A2(n6935), .ZN(n5429) );
  AND2_X1 U6214 ( .A1(n5502), .A2(n4948), .ZN(n5022) );
  AND2_X1 U6215 ( .A1(n5099), .A2(n6947), .ZN(n5023) );
  XOR2_X1 U6216 ( .A(n8479), .B(P2_REG1_REG_19__SCAN_IN), .Z(n5024) );
  AND2_X2 U6217 ( .A1(n6796), .A2(n7079), .ZN(n10677) );
  AND2_X1 U6218 ( .A1(n6373), .A2(n10518), .ZN(n5025) );
  INV_X1 U6219 ( .A(n8254), .ZN(n8441) );
  INV_X1 U6220 ( .A(n9211), .ZN(n9234) );
  NAND2_X1 U6221 ( .A1(n6289), .A2(n6862), .ZN(n9211) );
  NAND2_X1 U6222 ( .A1(n5242), .A2(n6250), .ZN(n7759) );
  NAND2_X1 U6223 ( .A1(n6933), .A2(n6932), .ZN(n7306) );
  AND2_X2 U6224 ( .A1(n6796), .A2(n6808), .ZN(n10681) );
  AND2_X1 U6225 ( .A1(n7517), .A2(n10613), .ZN(n9937) );
  NOR2_X1 U6226 ( .A1(n10419), .A2(n5664), .ZN(n5026) );
  OR2_X1 U6227 ( .A1(n5726), .A2(n5683), .ZN(n5027) );
  INV_X1 U6228 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5452) );
  XNOR2_X1 U6229 ( .A(n5620), .B(n8069), .ZN(n8065) );
  XNOR2_X1 U6230 ( .A(n5633), .B(n8994), .ZN(n8990) );
  MUX2_X1 U6231 ( .A(n8559), .B(n8558), .S(n8591), .Z(n8561) );
  OAI21_X1 U6232 ( .B1(n5223), .B2(n5004), .A(n8591), .ZN(n5218) );
  MUX2_X1 U6233 ( .A(n8524), .B(n8523), .S(n8591), .Z(n8535) );
  MUX2_X1 U6234 ( .A(n8504), .B(n8503), .S(n8591), .Z(n8513) );
  AOI211_X1 U6235 ( .C1(n10474), .C2(n9023), .A(n9022), .B(n9021), .ZN(n9028)
         );
  XNOR2_X1 U6236 ( .A(n5680), .B(n9023), .ZN(n9018) );
  AOI211_X1 U6237 ( .C1(n9632), .C2(n4924), .A(n9631), .B(n9630), .ZN(n9633)
         );
  NOR3_X1 U6238 ( .A1(n8341), .A2(n8340), .A3(n9181), .ZN(n8348) );
  AND2_X1 U6239 ( .A1(n8433), .A2(n8444), .ZN(n8478) );
  NAND2_X1 U6240 ( .A1(n8320), .A2(n8319), .ZN(n5198) );
  AOI21_X1 U6241 ( .B1(n5196), .B2(n5194), .A(n8324), .ZN(n8334) );
  OAI21_X1 U6242 ( .B1(n8477), .B2(n7409), .A(n5287), .ZN(n5286) );
  NAND2_X1 U6243 ( .A1(n5199), .A2(n4936), .ZN(n5349) );
  OAI21_X1 U6244 ( .B1(n8332), .B2(n8331), .A(n8330), .ZN(n5344) );
  NAND2_X1 U6245 ( .A1(n5028), .A2(n8304), .ZN(n8313) );
  NAND2_X1 U6246 ( .A1(n8292), .A2(n8293), .ZN(n5028) );
  OAI211_X1 U6247 ( .C1(n8283), .C2(n8387), .A(n8284), .B(n5352), .ZN(n8290)
         );
  NAND2_X1 U6248 ( .A1(n5349), .A2(n5346), .ZN(n5345) );
  INV_X1 U6249 ( .A(n5195), .ZN(n5194) );
  NOR2_X1 U6250 ( .A1(n8334), .A2(n9232), .ZN(n8332) );
  NAND2_X1 U6251 ( .A1(n8678), .A2(n6738), .ZN(n8679) );
  AOI22_X1 U6252 ( .A1(n8637), .A2(n5064), .B1(n5067), .B2(n5063), .ZN(n5065)
         );
  OAI211_X1 U6253 ( .C1(n8432), .C2(n8434), .A(n8470), .B(n8443), .ZN(n8433)
         );
  NAND2_X1 U6254 ( .A1(n5342), .A2(n8396), .ZN(n5341) );
  AOI21_X1 U6255 ( .B1(n8288), .B2(n8287), .A(n8396), .ZN(n5353) );
  OAI21_X1 U6256 ( .B1(n5213), .B2(n5001), .A(n5351), .ZN(n5212) );
  NAND2_X1 U6257 ( .A1(n5266), .A2(n4991), .ZN(n9126) );
  INV_X1 U6258 ( .A(n5029), .ZN(n6875) );
  INV_X1 U6259 ( .A(n5042), .ZN(n9250) );
  OAI21_X2 U6260 ( .B1(n8021), .B2(n6269), .A(n6268), .ZN(n8072) );
  NAND2_X1 U6261 ( .A1(n6878), .A2(n5043), .ZN(n5042) );
  OR2_X2 U6262 ( .A1(n10619), .A2(n7750), .ZN(n7810) );
  NAND2_X1 U6263 ( .A1(n5246), .A2(n5245), .ZN(n9087) );
  NAND2_X1 U6264 ( .A1(n5250), .A2(n5249), .ZN(n9185) );
  INV_X1 U6265 ( .A(n9160), .ZN(n5266) );
  NAND2_X1 U6266 ( .A1(n5198), .A2(n4955), .ZN(n5197) );
  XNOR2_X1 U6267 ( .A(n5286), .B(n8479), .ZN(n8487) );
  INV_X1 U6268 ( .A(n5353), .ZN(n5352) );
  OAI21_X1 U6269 ( .B1(n8332), .B2(n8327), .A(n8329), .ZN(n5342) );
  NAND2_X1 U6270 ( .A1(n5348), .A2(n8387), .ZN(n5347) );
  NAND2_X1 U6271 ( .A1(n5347), .A2(n5345), .ZN(n8432) );
  NAND2_X1 U6272 ( .A1(n5212), .A2(n4996), .ZN(n5211) );
  NAND2_X1 U6273 ( .A1(n5211), .A2(n8364), .ZN(n8365) );
  OAI21_X1 U6274 ( .B1(n8321), .B2(n8387), .A(n8325), .ZN(n5195) );
  NOR3_X1 U6275 ( .A1(n8347), .A2(n8348), .A3(n5000), .ZN(n5213) );
  NAND2_X1 U6276 ( .A1(n8029), .A2(n5033), .ZN(n5031) );
  NAND3_X1 U6277 ( .A1(n5031), .A2(n8318), .A3(n5030), .ZN(n8076) );
  AND2_X1 U6278 ( .A1(n5568), .A2(n5268), .ZN(n5740) );
  AOI21_X1 U6279 ( .B1(n9081), .B2(n8377), .A(n8378), .ZN(n9070) );
  NAND2_X1 U6280 ( .A1(n5050), .A2(n8449), .ZN(n5049) );
  NOR2_X1 U6281 ( .A1(n6248), .A2(n8255), .ZN(n7767) );
  NAND2_X1 U6282 ( .A1(n5057), .A2(n6064), .ZN(n6050) );
  NAND3_X1 U6283 ( .A1(n5840), .A2(n5843), .A3(n5060), .ZN(n5058) );
  NAND2_X1 U6284 ( .A1(n8734), .A2(n5067), .ZN(n5066) );
  NAND2_X1 U6285 ( .A1(n5066), .A2(n5065), .ZN(P1_U3242) );
  NAND3_X1 U6286 ( .A1(n5071), .A2(n8588), .A3(n9636), .ZN(n5070) );
  NAND4_X1 U6287 ( .A1(n8587), .A2(n8586), .A3(n8656), .A4(n8585), .ZN(n5071)
         );
  OAI22_X2 U6288 ( .A1(n5075), .A2(n5396), .B1(n5073), .B2(n9951), .ZN(n8602)
         );
  NAND2_X1 U6289 ( .A1(n5081), .A2(n7460), .ZN(n7469) );
  NAND3_X1 U6290 ( .A1(n5425), .A2(n5429), .A3(n7459), .ZN(n5081) );
  NAND2_X1 U6291 ( .A1(n9381), .A2(n5085), .ZN(n5084) );
  NAND2_X1 U6292 ( .A1(n9458), .A2(n5093), .ZN(n5092) );
  OAI21_X1 U6293 ( .B1(n9458), .B2(n5096), .A(n5093), .ZN(n9430) );
  AOI21_X1 U6294 ( .B1(n5093), .B2(n5096), .A(n5091), .ZN(n5090) );
  NAND2_X1 U6295 ( .A1(n8197), .A2(n5103), .ZN(n5100) );
  NAND2_X1 U6296 ( .A1(n5100), .A2(n5101), .ZN(n9481) );
  NAND3_X1 U6297 ( .A1(n6729), .A2(n6728), .A3(n6727), .ZN(n5109) );
  OAI21_X1 U6298 ( .B1(n7594), .B2(n5114), .A(n5112), .ZN(n7795) );
  NAND3_X1 U6299 ( .A1(n5111), .A2(n8530), .A3(n5110), .ZN(n6749) );
  NAND2_X1 U6300 ( .A1(n7594), .A2(n5112), .ZN(n5111) );
  NAND2_X2 U6301 ( .A1(n5115), .A2(n6453), .ZN(n7638) );
  NAND2_X1 U6302 ( .A1(n9653), .A2(n8654), .ZN(n9637) );
  NAND2_X1 U6303 ( .A1(n5130), .A2(n5128), .ZN(n9812) );
  OAI21_X1 U6304 ( .B1(n6646), .B2(n5146), .A(n5144), .ZN(n9684) );
  NAND2_X1 U6305 ( .A1(n5143), .A2(n5141), .ZN(n5471) );
  NAND2_X1 U6306 ( .A1(n6646), .A2(n5144), .ZN(n5143) );
  OAI21_X1 U6307 ( .B1(n6646), .B2(n5467), .A(n5465), .ZN(n9702) );
  AOI21_X1 U6308 ( .B1(n5465), .B2(n5467), .A(n4990), .ZN(n5147) );
  NAND2_X1 U6309 ( .A1(n5148), .A2(n5151), .ZN(n7574) );
  NAND3_X1 U6310 ( .A1(n5153), .A2(n5152), .A3(n5149), .ZN(n5148) );
  INV_X1 U6311 ( .A(n7511), .ZN(n5150) );
  OR2_X1 U6312 ( .A1(n7491), .A2(n9510), .ZN(n5151) );
  NAND2_X1 U6313 ( .A1(n5154), .A2(n5156), .ZN(n7651) );
  NAND2_X1 U6314 ( .A1(n7680), .A2(n5155), .ZN(n5154) );
  AND2_X1 U6315 ( .A1(n8613), .A2(n8614), .ZN(n5155) );
  NAND2_X1 U6316 ( .A1(n6693), .A2(n5160), .ZN(n5159) );
  INV_X1 U6317 ( .A(n8630), .ZN(n5163) );
  NAND2_X1 U6318 ( .A1(n6693), .A2(n6692), .ZN(n9652) );
  NAND2_X1 U6319 ( .A1(n9791), .A2(n4938), .ZN(n5170) );
  INV_X1 U6320 ( .A(n6625), .ZN(n5173) );
  NAND2_X1 U6321 ( .A1(n9791), .A2(n6613), .ZN(n9781) );
  NAND4_X1 U6322 ( .A1(n4951), .A2(n5176), .A3(n6325), .A4(n5174), .ZN(n6787)
         );
  NAND3_X1 U6323 ( .A1(n6381), .A2(n5470), .A3(n6324), .ZN(n6420) );
  AND3_X2 U6324 ( .A1(n5319), .A2(n6424), .A3(n4951), .ZN(n6734) );
  NOR2_X1 U6325 ( .A1(n7868), .A2(n8034), .ZN(n5181) );
  XNOR2_X2 U6326 ( .A(n5372), .B(n7202), .ZN(n7868) );
  NOR2_X1 U6327 ( .A1(n7867), .A2(n5669), .ZN(n7901) );
  NOR2_X1 U6328 ( .A1(n7868), .A2(n8034), .ZN(n7867) );
  INV_X1 U6329 ( .A(n5183), .ZN(n7899) );
  NAND2_X1 U6330 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n5185) );
  OR2_X2 U6331 ( .A1(n10433), .A2(n5188), .ZN(n5187) );
  XNOR2_X1 U6332 ( .A(n5678), .B(n8994), .ZN(n8981) );
  NAND4_X1 U6333 ( .A1(n5193), .A2(n10513), .A3(n10512), .A4(n10514), .ZN(
        P2_U3200) );
  NAND2_X1 U6334 ( .A1(n5205), .A2(n5200), .ZN(n5199) );
  NAND3_X1 U6335 ( .A1(n8311), .A2(n8285), .A3(n8282), .ZN(n8293) );
  OAI21_X1 U6336 ( .B1(n5216), .B2(n8561), .A(n4978), .ZN(n8570) );
  OAI21_X1 U6337 ( .B1(n8556), .B2(n8713), .A(n8714), .ZN(n8555) );
  AND2_X1 U6338 ( .A1(n5229), .A2(n5228), .ZN(n8556) );
  OAI21_X2 U6339 ( .B1(n5241), .B2(n5243), .A(n6251), .ZN(n7786) );
  INV_X1 U6340 ( .A(n6250), .ZN(n5244) );
  NAND2_X1 U6341 ( .A1(n6283), .A2(n5247), .ZN(n5246) );
  NAND2_X1 U6342 ( .A1(n9214), .A2(n5251), .ZN(n5250) );
  INV_X1 U6343 ( .A(n6274), .ZN(n5253) );
  NAND2_X1 U6344 ( .A1(n9214), .A2(n9213), .ZN(n9212) );
  NAND2_X1 U6345 ( .A1(n5260), .A2(n5261), .ZN(n9231) );
  NAND2_X1 U6346 ( .A1(n8072), .A2(n5262), .ZN(n5260) );
  INV_X2 U6347 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n5265) );
  NAND2_X1 U6348 ( .A1(n5568), .A2(n5547), .ZN(n5570) );
  NAND2_X1 U6349 ( .A1(n5568), .A2(n5267), .ZN(n5270) );
  NAND2_X1 U6350 ( .A1(n10415), .A2(n5273), .ZN(n5271) );
  XNOR2_X1 U6351 ( .A(n5274), .B(n7145), .ZN(n10451) );
  INV_X1 U6352 ( .A(n5274), .ZN(n5609) );
  INV_X1 U6353 ( .A(n5621), .ZN(n5276) );
  NOR2_X1 U6354 ( .A1(n8065), .A2(n10701), .ZN(n8064) );
  NOR2_X1 U6355 ( .A1(n9016), .A2(n10746), .ZN(n9015) );
  INV_X1 U6356 ( .A(n10500), .ZN(n5279) );
  INV_X1 U6357 ( .A(n7904), .ZN(n5282) );
  NOR2_X1 U6358 ( .A1(n10626), .A2(n10451), .ZN(n10450) );
  NOR2_X1 U6359 ( .A1(n10471), .A2(n10470), .ZN(n10469) );
  NAND2_X1 U6360 ( .A1(n9252), .A2(n9251), .ZN(n9253) );
  NAND2_X1 U6361 ( .A1(n6257), .A2(n6256), .ZN(n7665) );
  AOI211_X1 U6362 ( .C1(n8515), .C2(n8514), .A(n8695), .B(n8513), .ZN(n8519)
         );
  NAND2_X1 U6363 ( .A1(n6744), .A2(n6743), .ZN(n8497) );
  NAND2_X1 U6364 ( .A1(n5650), .A2(n5649), .ZN(n5738) );
  NAND2_X1 U6365 ( .A1(n5288), .A2(n5289), .ZN(n6116) );
  NAND2_X1 U6366 ( .A1(n9162), .A2(n4994), .ZN(n5288) );
  NAND2_X1 U6367 ( .A1(n9071), .A2(n5297), .ZN(n5296) );
  NAND2_X1 U6368 ( .A1(n9071), .A2(n6192), .ZN(n9049) );
  NAND2_X1 U6369 ( .A1(n5296), .A2(n5298), .ZN(n8476) );
  NAND2_X1 U6370 ( .A1(n5541), .A2(n5512), .ZN(n5542) );
  NAND2_X1 U6371 ( .A1(n5847), .A2(n5315), .ZN(n7809) );
  NAND2_X1 U6372 ( .A1(n7809), .A2(n5879), .ZN(n5880) );
  OR2_X1 U6373 ( .A1(n5793), .A2(n5777), .ZN(n5316) );
  INV_X1 U6374 ( .A(n5740), .ZN(n5573) );
  NAND4_X1 U6375 ( .A1(n5475), .A2(n4967), .A3(n6334), .A4(n5319), .ZN(n10001)
         );
  NAND2_X1 U6376 ( .A1(n6744), .A2(n5327), .ZN(n5328) );
  NAND2_X1 U6377 ( .A1(n7368), .A2(n6742), .ZN(n10539) );
  NAND2_X1 U6378 ( .A1(n6754), .A2(n5329), .ZN(n9688) );
  NAND2_X1 U6379 ( .A1(n5864), .A2(n5863), .ZN(n5333) );
  AND2_X1 U6380 ( .A1(n5339), .A2(n5338), .ZN(n8341) );
  NAND3_X1 U6381 ( .A1(n5343), .A2(n5341), .A3(n5340), .ZN(n5339) );
  NAND2_X1 U6382 ( .A1(n9794), .A2(n5357), .ZN(n9749) );
  NAND2_X2 U6383 ( .A1(n6362), .A2(n6363), .ZN(n7174) );
  OR2_X2 U6384 ( .A1(n8055), .A2(n5672), .ZN(n8163) );
  NOR2_X1 U6385 ( .A1(n8057), .A2(n8056), .ZN(n8055) );
  XNOR2_X1 U6386 ( .A(n5671), .B(n8069), .ZN(n8057) );
  NAND2_X1 U6387 ( .A1(n10503), .A2(n5726), .ZN(n5368) );
  OR2_X2 U6388 ( .A1(n10475), .A2(n5373), .ZN(n5372) );
  INV_X1 U6389 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n5382) );
  INV_X1 U6390 ( .A(P1_RD_REG_SCAN_IN), .ZN(n5381) );
  AND2_X4 U6391 ( .A1(n5380), .A2(n5379), .ZN(n8416) );
  INV_X1 U6392 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n5383) );
  NAND2_X1 U6393 ( .A1(n6196), .A2(n6195), .ZN(n6215) );
  NAND2_X1 U6394 ( .A1(n6085), .A2(n6084), .ZN(n5389) );
  NAND2_X1 U6395 ( .A1(n5389), .A2(n5017), .ZN(n6099) );
  NAND2_X1 U6396 ( .A1(n6145), .A2(n5393), .ZN(n5392) );
  NAND2_X1 U6397 ( .A1(n6145), .A2(n6144), .ZN(n6160) );
  OAI21_X1 U6398 ( .B1(n6032), .B2(n5401), .A(n5400), .ZN(n6067) );
  OAI21_X1 U6399 ( .B1(n5910), .B2(n5404), .A(n5406), .ZN(n5959) );
  OR2_X1 U6400 ( .A1(n5910), .A2(n5909), .ZN(n5412) );
  NAND2_X1 U6401 ( .A1(n9439), .A2(n9440), .ZN(n5416) );
  INV_X1 U6402 ( .A(n6981), .ZN(n5419) );
  AND2_X1 U6403 ( .A1(n6930), .A2(n7379), .ZN(n5424) );
  AND2_X1 U6404 ( .A1(n5429), .A2(n5425), .ZN(n7461) );
  NAND3_X1 U6405 ( .A1(n9362), .A2(n5435), .A3(n5433), .ZN(n5432) );
  NAND2_X1 U6406 ( .A1(n5446), .A2(n5447), .ZN(n6946) );
  NAND2_X1 U6407 ( .A1(n6734), .A2(n5449), .ZN(n6777) );
  NAND2_X1 U6408 ( .A1(n6734), .A2(n4988), .ZN(n5450) );
  NAND2_X1 U6409 ( .A1(n5453), .A2(n10540), .ZN(n6385) );
  XNOR2_X1 U6410 ( .A(n5453), .B(n10540), .ZN(n10560) );
  NAND2_X1 U6411 ( .A1(n6375), .A2(n6374), .ZN(n5453) );
  NAND2_X1 U6412 ( .A1(n8087), .A2(n5455), .ZN(n5454) );
  INV_X1 U6413 ( .A(n6398), .ZN(n5461) );
  NAND2_X1 U6414 ( .A1(n7511), .A2(n6745), .ZN(n5462) );
  NAND2_X1 U6415 ( .A1(n5471), .A2(n5472), .ZN(n6693) );
  XNOR2_X1 U6416 ( .A(n6805), .B(n6814), .ZN(n6840) );
  OAI21_X1 U6417 ( .B1(n6840), .B2(n9937), .A(n6839), .ZN(n6843) );
  NAND2_X1 U6418 ( .A1(n5740), .A2(n5477), .ZN(n9335) );
  NAND2_X1 U6419 ( .A1(n7613), .A2(n7612), .ZN(n7611) );
  NAND2_X1 U6420 ( .A1(n7611), .A2(n5482), .ZN(n7421) );
  INV_X1 U6421 ( .A(n5481), .ZN(n7504) );
  NAND2_X1 U6422 ( .A1(n8839), .A2(n5486), .ZN(n5483) );
  NAND2_X1 U6423 ( .A1(n5483), .A2(n5484), .ZN(n8799) );
  OAI21_X1 U6424 ( .B1(n8839), .B2(n5485), .A(n5488), .ZN(n8805) );
  AOI21_X1 U6425 ( .B1(n8839), .B2(n8792), .A(n5521), .ZN(n8903) );
  NAND2_X1 U6426 ( .A1(n7719), .A2(n4934), .ZN(n5501) );
  INV_X1 U6427 ( .A(n5502), .ZN(n7749) );
  NAND2_X1 U6428 ( .A1(n4946), .A2(n5506), .ZN(n5554) );
  OAI21_X1 U6429 ( .B1(n8851), .B2(n5509), .A(n5507), .ZN(n8891) );
  OAI21_X1 U6430 ( .B1(n6848), .B2(n5520), .A(n10643), .ZN(n6323) );
  NAND2_X1 U6431 ( .A1(n9250), .A2(n10761), .ZN(n9252) );
  NAND2_X1 U6432 ( .A1(n9038), .A2(n10749), .ZN(n6878) );
  OR2_X1 U6433 ( .A1(n6823), .A2(n8753), .ZN(n8660) );
  NAND2_X1 U6434 ( .A1(n9471), .A2(n7076), .ZN(n8742) );
  AOI21_X1 U6435 ( .B1(n8476), .B2(n5529), .A(n5513), .ZN(n8477) );
  OR2_X1 U6436 ( .A1(n6386), .A2(n6364), .ZN(n6366) );
  NAND2_X1 U6437 ( .A1(n6902), .A2(n6919), .ZN(n6899) );
  NOR2_X1 U6438 ( .A1(n8671), .A2(n7174), .ZN(n9821) );
  NAND2_X1 U6439 ( .A1(n7628), .A2(n5755), .ZN(n8263) );
  INV_X1 U6440 ( .A(n6342), .ZN(n10006) );
  INV_X1 U6441 ( .A(n8488), .ZN(n6738) );
  OR2_X1 U6442 ( .A1(n6840), .A2(n9836), .ZN(n6835) );
  NAND2_X1 U6443 ( .A1(n6915), .A2(n7366), .ZN(n6900) );
  AND4_X1 U6444 ( .A1(n5540), .A2(n5559), .A3(n5641), .A4(n5555), .ZN(n5512)
         );
  AND2_X1 U6445 ( .A1(n8475), .A2(n8254), .ZN(n5513) );
  AND2_X1 U6446 ( .A1(n9771), .A2(n8718), .ZN(n5514) );
  AND2_X1 U6447 ( .A1(n8755), .A2(n9499), .ZN(n5516) );
  INV_X1 U6448 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n5656) );
  AND2_X1 U6449 ( .A1(P2_U3893), .A2(n5648), .ZN(n10495) );
  INV_X1 U6450 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n8223) );
  INV_X1 U6451 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n5613) );
  AND2_X1 U6452 ( .A1(n5897), .A2(n5886), .ZN(n5517) );
  NOR2_X1 U6453 ( .A1(n6931), .A2(n4949), .ZN(n5518) );
  OR2_X1 U6454 ( .A1(n9959), .A2(n9480), .ZN(n5519) );
  AND2_X1 U6455 ( .A1(n6846), .A2(n7693), .ZN(n5520) );
  NOR2_X1 U6456 ( .A1(n8791), .A2(n8842), .ZN(n5521) );
  NOR2_X1 U6457 ( .A1(n7409), .A2(n6862), .ZN(n5522) );
  AND2_X1 U6458 ( .A1(n7758), .A2(n7750), .ZN(n5523) );
  INV_X1 U6459 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5816) );
  INV_X1 U6460 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n5777) );
  INV_X1 U6461 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n6002) );
  INV_X1 U6462 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n5872) );
  INV_X1 U6463 ( .A(n10764), .ZN(n6872) );
  NAND2_X1 U6464 ( .A1(n7620), .A2(n10638), .ZN(n10643) );
  INV_X1 U6465 ( .A(n9201), .ZN(n8932) );
  NOR2_X1 U6466 ( .A1(n5889), .A2(n5874), .ZN(n5525) );
  NOR2_X1 U6467 ( .A1(n8361), .A2(n9116), .ZN(n5526) );
  NAND2_X1 U6468 ( .A1(n10681), .A2(n10610), .ZN(n9995) );
  INV_X1 U6469 ( .A(n9995), .ZN(n6798) );
  NAND2_X2 U6470 ( .A1(n6825), .A2(n9854), .ZN(n10524) );
  INV_X1 U6471 ( .A(n8604), .ZN(n6814) );
  AND2_X1 U6472 ( .A1(n8778), .A2(n9148), .ZN(n5527) );
  INV_X1 U6473 ( .A(n5844), .ZN(n10435) );
  INV_X1 U6474 ( .A(n10510), .ZN(n10494) );
  OR2_X1 U6475 ( .A1(n7765), .A2(n8484), .ZN(n10684) );
  AND2_X2 U6476 ( .A1(n6854), .A2(n6853), .ZN(n10761) );
  NOR2_X1 U6477 ( .A1(n8282), .A2(n7885), .ZN(n5528) );
  AND2_X1 U6478 ( .A1(n8442), .A2(n8441), .ZN(n5529) );
  AND3_X1 U6479 ( .A1(n8469), .A2(n8436), .A3(n8435), .ZN(n5530) );
  INV_X1 U6480 ( .A(n6922), .ZN(n6920) );
  INV_X1 U6481 ( .A(n7414), .ZN(n5755) );
  INV_X1 U6482 ( .A(n8448), .ZN(n5830) );
  NOR2_X1 U6483 ( .A1(n6869), .A2(n9327), .ZN(n5531) );
  INV_X1 U6484 ( .A(n9327), .ZN(n6880) );
  INV_X1 U6485 ( .A(n8623), .ZN(n6551) );
  NAND2_X1 U6486 ( .A1(n8941), .A2(n8266), .ZN(n8267) );
  AND2_X1 U6487 ( .A1(n8294), .A2(n8267), .ZN(n8268) );
  NAND2_X1 U6488 ( .A1(n8269), .A2(n8268), .ZN(n8270) );
  NAND2_X1 U6489 ( .A1(n8270), .A2(n8396), .ZN(n8271) );
  NAND2_X1 U6490 ( .A1(n8272), .A2(n8271), .ZN(n8274) );
  NAND2_X1 U6491 ( .A1(n8567), .A2(n8565), .ZN(n8562) );
  INV_X1 U6492 ( .A(n9117), .ZN(n8359) );
  INV_X1 U6493 ( .A(n8363), .ZN(n8364) );
  OR2_X1 U6494 ( .A1(n9030), .A2(n9305), .ZN(n8436) );
  MUX2_X1 U6495 ( .A(n8665), .B(n8660), .S(n8591), .Z(n8592) );
  INV_X1 U6496 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n6331) );
  NAND2_X1 U6497 ( .A1(n8440), .A2(n9030), .ZN(n8442) );
  INV_X1 U6498 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n5661) );
  INV_X1 U6499 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n6329) );
  INV_X1 U6500 ( .A(n4925), .ZN(n5657) );
  NOR2_X1 U6501 ( .A1(n5528), .A2(n5523), .ZN(n6259) );
  INV_X1 U6502 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n6730) );
  AND2_X1 U6503 ( .A1(n7765), .A2(n8254), .ZN(n7407) );
  NOR2_X1 U6504 ( .A1(n5844), .A2(n5832), .ZN(n5608) );
  INV_X1 U6505 ( .A(n5631), .ZN(n5632) );
  OR2_X1 U6506 ( .A1(n9407), .A2(n9408), .ZN(n7000) );
  INV_X1 U6507 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n6001) );
  OAI21_X1 U6508 ( .B1(n4925), .B2(n5656), .A(n5655), .ZN(n7291) );
  NOR2_X1 U6509 ( .A1(n5603), .A2(n7318), .ZN(n10400) );
  OR2_X1 U6510 ( .A1(n9260), .A2(n8929), .ZN(n6286) );
  INV_X1 U6511 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n5932) );
  INV_X1 U6512 ( .A(n7760), .ZN(n8449) );
  INV_X1 U6513 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5739) );
  INV_X1 U6514 ( .A(n6638), .ZN(n6636) );
  INV_X1 U6515 ( .A(n6545), .ZN(n6543) );
  OAI22_X1 U6516 ( .A1(n6895), .A2(n8744), .B1(n6892), .B2(n6890), .ZN(n6893)
         );
  INV_X1 U6517 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n7358) );
  INV_X1 U6518 ( .A(n6621), .ZN(n6619) );
  INV_X1 U6519 ( .A(SI_25_), .ZN(n10123) );
  INV_X1 U6520 ( .A(SI_19_), .ZN(n10129) );
  INV_X1 U6521 ( .A(SI_16_), .ZN(n10140) );
  INV_X1 U6522 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n6446) );
  NOR2_X1 U6523 ( .A1(n6054), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6076) );
  NAND2_X1 U6524 ( .A1(n4930), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5759) );
  NOR2_X1 U6525 ( .A1(n5660), .A2(n7326), .ZN(n10397) );
  NOR2_X1 U6526 ( .A1(n10510), .A2(n5643), .ZN(n5645) );
  NAND2_X1 U6527 ( .A1(n6167), .A2(n10184), .ZN(n6186) );
  AND2_X1 U6528 ( .A1(n8366), .A2(n8367), .ZN(n8465) );
  NOR2_X1 U6529 ( .A1(n5949), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5971) );
  OR2_X1 U6530 ( .A1(n7155), .A2(n6315), .ZN(n6864) );
  INV_X1 U6531 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5742) );
  INV_X1 U6532 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5576) );
  NAND2_X1 U6533 ( .A1(n9481), .A2(n9483), .ZN(n6984) );
  INV_X1 U6534 ( .A(n6931), .ZN(n6932) );
  INV_X1 U6535 ( .A(n6496), .ZN(n6494) );
  NAND2_X1 U6536 ( .A1(n6696), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n6719) );
  NAND2_X1 U6537 ( .A1(n6636), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n6652) );
  OR2_X1 U6538 ( .A1(n6483), .A2(n6482), .ZN(n6496) );
  AND2_X1 U6539 ( .A1(n6898), .A2(n8743), .ZN(n6936) );
  NAND2_X1 U6540 ( .A1(n9805), .A2(n9806), .ZN(n9804) );
  NAND2_X1 U6541 ( .A1(n10571), .A2(n10544), .ZN(n8498) );
  INV_X1 U6542 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n10203) );
  INV_X1 U6543 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n6334) );
  NOR2_X1 U6544 ( .A1(n6356), .A2(n6355), .ZN(n6357) );
  INV_X1 U6545 ( .A(SI_21_), .ZN(n6087) );
  AND2_X1 U6546 ( .A1(n6570), .A2(n6569), .ZN(n6573) );
  NOR2_X1 U6547 ( .A1(n6508), .A2(n6507), .ZN(n6513) );
  INV_X1 U6548 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n5792) );
  INV_X1 U6549 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5547) );
  OR2_X1 U6550 ( .A1(n8770), .A2(n10739), .ZN(n8771) );
  XNOR2_X1 U6551 ( .A(n7416), .B(n7628), .ZN(n7527) );
  OR2_X1 U6552 ( .A1(n8762), .A2(n9237), .ZN(n8763) );
  INV_X1 U6553 ( .A(n8922), .ZN(n8897) );
  AOI21_X1 U6554 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n7337), .A(n8961), .ZN(
        n5678) );
  INV_X1 U6555 ( .A(n8928), .ZN(n9053) );
  NAND2_X1 U6556 ( .A1(n7430), .A2(n6318), .ZN(n9238) );
  OR2_X1 U6557 ( .A1(n7406), .A2(n7135), .ZN(n6861) );
  INV_X1 U6558 ( .A(n9512), .ZN(n7513) );
  INV_X1 U6559 ( .A(n6902), .ZN(n7215) );
  OR2_X1 U6560 ( .A1(n6609), .A2(n6608), .ZN(n6621) );
  INV_X1 U6561 ( .A(n9689), .ZN(n9476) );
  OR2_X1 U6562 ( .A1(n6719), .A2(n6718), .ZN(n6828) );
  AND2_X1 U6563 ( .A1(n10519), .A2(n6888), .ZN(n10537) );
  INV_X1 U6564 ( .A(n9505), .ZN(n7860) );
  INV_X1 U6565 ( .A(n10546), .ZN(n9759) );
  INV_X1 U6566 ( .A(n10537), .ZN(n9797) );
  AND2_X1 U6567 ( .A1(n8512), .A2(n8499), .ZN(n8609) );
  AND2_X1 U6568 ( .A1(n6033), .A2(n6005), .ZN(n6031) );
  OR2_X1 U6569 ( .A1(n6526), .A2(P1_IR_REG_13__SCAN_IN), .ZN(n6537) );
  OAI21_X1 U6570 ( .B1(n5778), .B2(n5777), .A(n5776), .ZN(n5788) );
  AOI21_X1 U6571 ( .B1(n7923), .B2(n7922), .A(n7921), .ZN(n7926) );
  INV_X1 U6572 ( .A(n8918), .ZN(n8895) );
  OR2_X1 U6573 ( .A1(n4929), .A2(n9041), .ZN(n6222) );
  AND2_X1 U6574 ( .A1(n6012), .A2(n6011), .ZN(n9201) );
  INV_X1 U6575 ( .A(n8163), .ZN(n8167) );
  AND2_X1 U6576 ( .A1(n5729), .A2(n9344), .ZN(n7259) );
  AND2_X1 U6577 ( .A1(n8305), .A2(n8314), .ZN(n8457) );
  INV_X1 U6578 ( .A(n9238), .ZN(n9222) );
  OAI21_X1 U6579 ( .B1(n6869), .B2(n9288), .A(n6857), .ZN(n6858) );
  AND2_X1 U6580 ( .A1(n6861), .A2(n6316), .ZN(n6853) );
  NOR2_X1 U6581 ( .A1(n10764), .A2(n6867), .ZN(n6870) );
  INV_X1 U6582 ( .A(n10749), .ZN(n10710) );
  INV_X1 U6583 ( .A(n10740), .ZN(n10751) );
  NAND2_X1 U6584 ( .A1(n10683), .A2(n10684), .ZN(n10749) );
  NAND2_X1 U6585 ( .A1(n6866), .A2(n6865), .ZN(n6868) );
  INV_X1 U6586 ( .A(n6303), .ZN(n8243) );
  AND2_X1 U6587 ( .A1(n7214), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9486) );
  INV_X1 U6588 ( .A(n9434), .ZN(n9488) );
  NAND2_X1 U6589 ( .A1(n6676), .A2(n6675), .ZN(n9707) );
  INV_X1 U6590 ( .A(n8491), .ZN(n6759) );
  OR2_X1 U6591 ( .A1(n6386), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n6389) );
  OR2_X1 U6592 ( .A1(n6386), .A2(n6376), .ZN(n6379) );
  INV_X1 U6593 ( .A(n10383), .ZN(n10329) );
  INV_X1 U6594 ( .A(n10338), .ZN(n10390) );
  INV_X1 U6595 ( .A(n8605), .ZN(n9757) );
  NAND2_X1 U6596 ( .A1(n10537), .A2(n6809), .ZN(n9854) );
  AOI21_X1 U6597 ( .B1(n6792), .B2(n7148), .A(n7150), .ZN(n7079) );
  INV_X1 U6598 ( .A(n10669), .ZN(n10610) );
  INV_X1 U6599 ( .A(n9937), .ZN(n10675) );
  AND2_X1 U6600 ( .A1(n6789), .A2(n10277), .ZN(n6796) );
  XNOR2_X1 U6601 ( .A(n6788), .B(n5452), .ZN(n7124) );
  AND2_X1 U6602 ( .A1(n6574), .A2(n6586), .ZN(n8214) );
  CLKBUF_X1 U6603 ( .A(n10003), .Z(n10012) );
  OR3_X1 U6604 ( .A1(n8240), .A2(n6303), .A3(n6298), .ZN(n7444) );
  AND2_X1 U6605 ( .A1(n7453), .A2(n7452), .ZN(n8919) );
  NAND2_X1 U6606 ( .A1(n7429), .A2(n7428), .ZN(n8912) );
  AND4_X1 U6607 ( .A1(n8431), .A2(n6240), .A3(n6239), .A4(n6238), .ZN(n9040)
         );
  INV_X1 U6608 ( .A(n8833), .ZN(n9130) );
  INV_X1 U6609 ( .A(n9235), .ZN(n8934) );
  OR2_X1 U6610 ( .A1(P2_U3150), .A2(n5731), .ZN(n10489) );
  NAND2_X1 U6611 ( .A1(n7259), .A2(n5685), .ZN(n10506) );
  INV_X1 U6612 ( .A(n5735), .ZN(n5736) );
  INV_X1 U6613 ( .A(n9223), .ZN(n10647) );
  INV_X1 U6614 ( .A(n10643), .ZN(n9223) );
  INV_X1 U6615 ( .A(n6858), .ZN(n6859) );
  INV_X1 U6616 ( .A(n10761), .ZN(n10760) );
  AND3_X1 U6617 ( .A1(n10588), .A2(n10587), .A3(n10586), .ZN(n10591) );
  AND2_X2 U6618 ( .A1(n6868), .A2(n7428), .ZN(n10764) );
  NAND2_X1 U6619 ( .A1(n7428), .A2(n7155), .ZN(n7225) );
  INV_X1 U6620 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n8238) );
  INV_X1 U6621 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7608) );
  INV_X1 U6622 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n7152) );
  INV_X1 U6623 ( .A(n9345), .ZN(n8237) );
  INV_X1 U6624 ( .A(n9486), .ZN(n9454) );
  INV_X1 U6625 ( .A(n9858), .ZN(n8149) );
  OR2_X1 U6626 ( .A1(n7092), .A2(n7080), .ZN(n9496) );
  NAND2_X1 U6627 ( .A1(n6704), .A2(n6703), .ZN(n9673) );
  INV_X1 U6628 ( .A(n9412), .ZN(n9776) );
  NAND2_X1 U6629 ( .A1(n7126), .A2(n7127), .ZN(n10394) );
  INV_X1 U6630 ( .A(n10524), .ZN(n10555) );
  INV_X1 U6631 ( .A(n10524), .ZN(n9800) );
  NAND2_X1 U6632 ( .A1(n8755), .A2(n9940), .ZN(n6794) );
  NAND2_X1 U6633 ( .A1(n10677), .A2(n10610), .ZN(n9934) );
  INV_X1 U6634 ( .A(n10677), .ZN(n10676) );
  INV_X1 U6635 ( .A(n9645), .ZN(n9959) );
  NAND2_X1 U6636 ( .A1(n7149), .A2(n7146), .ZN(n10018) );
  NAND2_X1 U6637 ( .A1(n6890), .A2(n7101), .ZN(n10279) );
  OAI21_X1 U6638 ( .B1(n6873), .B2(n10760), .A(n6859), .ZN(P2_U3488) );
  OAI21_X1 U6639 ( .B1(n6873), .B2(n6872), .A(n6871), .ZN(P2_U3456) );
  NAND2_X1 U6640 ( .A1(n6835), .A2(n6834), .ZN(P1_U3356) );
  NOR2_X1 U6641 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n5536) );
  NOR2_X1 U6642 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n5535) );
  NOR2_X1 U6643 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n5540) );
  NAND2_X1 U6644 ( .A1(n5551), .A2(n5552), .ZN(n5543) );
  NAND2_X1 U6645 ( .A1(n5550), .A2(n5549), .ZN(n5544) );
  NAND2_X1 U6646 ( .A1(n5567), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5548) );
  INV_X1 U6647 ( .A(n7228), .ZN(n5553) );
  NOR2_X4 U6648 ( .A1(n7444), .A2(n5553), .ZN(P2_U3893) );
  INV_X1 U6649 ( .A(n7444), .ZN(n5565) );
  NAND2_X1 U6650 ( .A1(n5554), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5622) );
  NAND2_X1 U6651 ( .A1(n5622), .A2(n5555), .ZN(n5556) );
  NAND2_X1 U6652 ( .A1(n5557), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5558) );
  OAI21_X2 U6653 ( .B1(n5642), .B2(P2_IR_REG_18__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5646) );
  NAND2_X1 U6654 ( .A1(n5646), .A2(n5559), .ZN(n5560) );
  NAND2_X1 U6655 ( .A1(n6242), .A2(n6241), .ZN(n5561) );
  XNOR2_X2 U6656 ( .A(n5563), .B(n5562), .ZN(n8254) );
  NAND2_X1 U6657 ( .A1(n5015), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5564) );
  OR2_X1 U6658 ( .A1(n5565), .A2(n8396), .ZN(n5566) );
  NAND2_X1 U6659 ( .A1(n5566), .A2(n7443), .ZN(n5729) );
  NAND2_X1 U6660 ( .A1(n5570), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5571) );
  NAND2_X1 U6661 ( .A1(n5729), .A2(n5765), .ZN(n5574) );
  NAND2_X1 U6662 ( .A1(n5574), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  NAND2_X1 U6663 ( .A1(n5575), .A2(n5576), .ZN(n5577) );
  NAND2_X1 U6664 ( .A1(n5577), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5630) );
  NAND2_X1 U6665 ( .A1(n5630), .A2(n5629), .ZN(n5578) );
  NAND2_X1 U6666 ( .A1(n5578), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5581) );
  NAND2_X1 U6667 ( .A1(n5581), .A2(n5579), .ZN(n5580) );
  NAND2_X1 U6668 ( .A1(n5580), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5636) );
  XNOR2_X1 U6669 ( .A(n5636), .B(P2_IR_REG_16__SCAN_IN), .ZN(n9012) );
  INV_X1 U6670 ( .A(n9012), .ZN(n7610) );
  XNOR2_X1 U6671 ( .A(n5581), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8994) );
  OR2_X1 U6672 ( .A1(n4946), .A2(n5617), .ZN(n5582) );
  XNOR2_X1 U6673 ( .A(n5582), .B(P2_IR_REG_10__SCAN_IN), .ZN(n7908) );
  NOR2_X1 U6674 ( .A1(n5583), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n5589) );
  NAND2_X1 U6675 ( .A1(n5589), .A2(n5584), .ZN(n5606) );
  OAI21_X1 U6676 ( .B1(n5611), .B2(P2_IR_REG_8__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5585) );
  XNOR2_X1 U6677 ( .A(n5585), .B(P2_IR_REG_9__SCAN_IN), .ZN(n7881) );
  NAND2_X1 U6678 ( .A1(n5586), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5587) );
  MUX2_X1 U6679 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5587), .S(
        P2_IR_REG_7__SCAN_IN), .Z(n5588) );
  OR2_X1 U6680 ( .A1(n5589), .A2(n5617), .ZN(n5590) );
  XNOR2_X1 U6681 ( .A(n5590), .B(P2_IR_REG_5__SCAN_IN), .ZN(n10418) );
  NAND2_X1 U6682 ( .A1(n5583), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5591) );
  XNOR2_X1 U6683 ( .A(n5591), .B(P2_IR_REG_4__SCAN_IN), .ZN(n5810) );
  NAND2_X1 U6684 ( .A1(n5597), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5592) );
  MUX2_X1 U6685 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5592), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n5593) );
  AND2_X1 U6686 ( .A1(n5593), .A2(n5583), .ZN(n5794) );
  AND2_X1 U6687 ( .A1(n5265), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5598) );
  NAND2_X1 U6688 ( .A1(n5651), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5600) );
  INV_X1 U6689 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n5599) );
  NAND2_X1 U6690 ( .A1(n7278), .A2(n5600), .ZN(n7294) );
  OAI21_X1 U6691 ( .B1(n4925), .B2(n5766), .A(n5601), .ZN(n7295) );
  AOI21_X1 U6692 ( .B1(P2_REG1_REG_2__SCAN_IN), .B2(n4925), .A(n7297), .ZN(
        n5602) );
  NOR2_X1 U6693 ( .A1(n5794), .A2(n5602), .ZN(n5603) );
  INV_X1 U6694 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10581) );
  XNOR2_X1 U6695 ( .A(n5794), .B(n5602), .ZN(n7319) );
  NOR2_X1 U6696 ( .A1(n10581), .A2(n7319), .ZN(n7318) );
  INV_X1 U6697 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10589) );
  AOI22_X1 U6698 ( .A1(n5810), .A2(P2_REG1_REG_4__SCAN_IN), .B1(n10589), .B2(
        n10406), .ZN(n10399) );
  NOR2_X1 U6699 ( .A1(n10400), .A2(n10399), .ZN(n10398) );
  NOR2_X1 U6700 ( .A1(n10418), .A2(n5604), .ZN(n5605) );
  INV_X1 U6701 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n10605) );
  INV_X1 U6702 ( .A(n10418), .ZN(n7118) );
  XOR2_X1 U6703 ( .A(n7118), .B(n5604), .Z(n10416) );
  NOR2_X1 U6704 ( .A1(n10605), .A2(n10416), .ZN(n10415) );
  INV_X1 U6705 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n5832) );
  NAND2_X1 U6706 ( .A1(n5606), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5607) );
  XNOR2_X1 U6707 ( .A(n5607), .B(P2_IR_REG_6__SCAN_IN), .ZN(n5844) );
  MUX2_X1 U6708 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n5832), .S(n5844), .Z(n10443)
         );
  NOR2_X1 U6709 ( .A1(n10453), .A2(n5609), .ZN(n5610) );
  INV_X1 U6710 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n10626) );
  NAND2_X1 U6711 ( .A1(n5611), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5612) );
  XNOR2_X1 U6712 ( .A(n5612), .B(P2_IR_REG_8__SCAN_IN), .ZN(n10473) );
  AOI22_X1 U6713 ( .A1(n10473), .A2(P2_REG1_REG_8__SCAN_IN), .B1(n5613), .B2(
        n7154), .ZN(n10470) );
  NOR2_X1 U6714 ( .A1(n7881), .A2(n5615), .ZN(n5616) );
  INV_X1 U6715 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n10665) );
  INV_X1 U6716 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n10691) );
  AOI22_X1 U6717 ( .A1(n7908), .A2(P2_REG1_REG_10__SCAN_IN), .B1(n10691), .B2(
        n7207), .ZN(n7904) );
  OR2_X1 U6718 ( .A1(n5618), .A2(n5617), .ZN(n5619) );
  XNOR2_X1 U6719 ( .A(n5619), .B(P2_IR_REG_11__SCAN_IN), .ZN(n8069) );
  INV_X1 U6720 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n10701) );
  NOR2_X1 U6721 ( .A1(n8069), .A2(n5620), .ZN(n5621) );
  INV_X1 U6722 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n5624) );
  XNOR2_X1 U6723 ( .A(n5622), .B(P2_IR_REG_12__SCAN_IN), .ZN(n8180) );
  MUX2_X1 U6724 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n5624), .S(n8180), .Z(n8175)
         );
  INV_X1 U6725 ( .A(n8175), .ZN(n5623) );
  OR2_X1 U6726 ( .A1(n8180), .A2(n5624), .ZN(n5625) );
  XNOR2_X1 U6727 ( .A(n5575), .B(P2_IR_REG_13__SCAN_IN), .ZN(n8958) );
  INV_X1 U6728 ( .A(n8958), .ZN(n7314) );
  INV_X1 U6729 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n10715) );
  INV_X1 U6730 ( .A(n5626), .ZN(n5627) );
  NOR2_X1 U6731 ( .A1(n8958), .A2(n5627), .ZN(n5628) );
  XNOR2_X1 U6732 ( .A(n5630), .B(n5629), .ZN(n7337) );
  NAND2_X1 U6733 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n7337), .ZN(n5631) );
  OAI21_X1 U6734 ( .B1(P2_REG1_REG_14__SCAN_IN), .B2(n7337), .A(n5631), .ZN(
        n8971) );
  NOR2_X1 U6735 ( .A1(n8994), .A2(n5633), .ZN(n5634) );
  INV_X1 U6736 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n10729) );
  INV_X1 U6737 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n10736) );
  AOI22_X1 U6738 ( .A1(n9012), .A2(P2_REG1_REG_16__SCAN_IN), .B1(n10736), .B2(
        n7610), .ZN(n9008) );
  INV_X1 U6739 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5635) );
  NAND2_X1 U6740 ( .A1(n5636), .A2(n5635), .ZN(n5637) );
  NAND2_X1 U6741 ( .A1(n5637), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5638) );
  XNOR2_X1 U6742 ( .A(n5638), .B(P2_IR_REG_17__SCAN_IN), .ZN(n9023) );
  XNOR2_X1 U6743 ( .A(n5639), .B(n9023), .ZN(n9016) );
  INV_X1 U6744 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n10746) );
  NOR2_X1 U6745 ( .A1(n9023), .A2(n5639), .ZN(n5640) );
  XNOR2_X1 U6746 ( .A(n5642), .B(n5641), .ZN(n10510) );
  INV_X1 U6747 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n5643) );
  NOR2_X1 U6748 ( .A1(n10494), .A2(n5643), .ZN(n5644) );
  AOI21_X1 U6749 ( .B1(n10494), .B2(n5643), .A(n5644), .ZN(n10500) );
  XNOR2_X1 U6750 ( .A(n5647), .B(n5024), .ZN(n5650) );
  NOR2_X1 U6751 ( .A1(n5648), .A2(P2_U3151), .ZN(n9344) );
  NAND2_X1 U6752 ( .A1(n7259), .A2(n4928), .ZN(n10501) );
  INV_X1 U6753 ( .A(n10501), .ZN(n5649) );
  INV_X1 U6754 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n8056) );
  AND2_X1 U6755 ( .A1(n5265), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5652) );
  NAND2_X1 U6756 ( .A1(n5651), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5653) );
  INV_X1 U6757 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n7271) );
  NOR2_X1 U6758 ( .A1(n7270), .A2(n7271), .ZN(n7269) );
  INV_X1 U6759 ( .A(n5653), .ZN(n5654) );
  NOR2_X2 U6760 ( .A1(n7293), .A2(n5658), .ZN(n5659) );
  NOR2_X1 U6761 ( .A1(n5794), .A2(n5659), .ZN(n5660) );
  INV_X1 U6762 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n7328) );
  INV_X1 U6763 ( .A(n5794), .ZN(n7334) );
  XNOR2_X1 U6764 ( .A(n5659), .B(n5794), .ZN(n7327) );
  NOR2_X1 U6765 ( .A1(n7328), .A2(n7327), .ZN(n7326) );
  AOI22_X1 U6766 ( .A1(n5810), .A2(P2_REG2_REG_4__SCAN_IN), .B1(n5661), .B2(
        n10406), .ZN(n10396) );
  NOR2_X1 U6767 ( .A1(n10397), .A2(n10396), .ZN(n10395) );
  NOR2_X1 U6768 ( .A1(n10418), .A2(n5663), .ZN(n5664) );
  INV_X1 U6769 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n10421) );
  INV_X1 U6770 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n5665) );
  AOI22_X1 U6771 ( .A1(P2_REG2_REG_6__SCAN_IN), .A2(n5844), .B1(n10435), .B2(
        n5665), .ZN(n10434) );
  NOR2_X1 U6772 ( .A1(n10453), .A2(n5666), .ZN(n5667) );
  INV_X1 U6773 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n10456) );
  NOR2_X1 U6774 ( .A1(n5667), .A2(n10454), .ZN(n10477) );
  INV_X1 U6775 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n10646) );
  AOI22_X1 U6776 ( .A1(n10473), .A2(P2_REG2_REG_8__SCAN_IN), .B1(n10646), .B2(
        n7154), .ZN(n10476) );
  NOR2_X1 U6777 ( .A1(n7881), .A2(n5668), .ZN(n5669) );
  INV_X1 U6778 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n8034) );
  INV_X1 U6779 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n5670) );
  AOI22_X1 U6780 ( .A1(n7908), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n5670), .B2(
        n7207), .ZN(n7900) );
  AOI21_X2 U6781 ( .B1(P2_REG2_REG_10__SCAN_IN), .B2(n7207), .A(n7899), .ZN(
        n5671) );
  NOR2_X1 U6782 ( .A1(n8069), .A2(n5671), .ZN(n5672) );
  INV_X1 U6783 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n5935) );
  MUX2_X1 U6784 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n5935), .S(n8180), .Z(n8166)
         );
  INV_X1 U6785 ( .A(n8166), .ZN(n5673) );
  OR2_X1 U6786 ( .A1(n8180), .A2(n5935), .ZN(n5674) );
  INV_X1 U6787 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n8944) );
  NAND2_X1 U6788 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n7337), .ZN(n5677) );
  OAI21_X1 U6789 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n7337), .A(n5677), .ZN(
        n8962) );
  NOR2_X1 U6790 ( .A1(n8994), .A2(n5678), .ZN(n5679) );
  INV_X1 U6791 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8980) );
  INV_X1 U6792 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n6017) );
  MUX2_X1 U6793 ( .A(P2_REG2_REG_16__SCAN_IN), .B(n6017), .S(n9012), .Z(n8998)
         );
  NOR2_X1 U6794 ( .A1(n9023), .A2(n5680), .ZN(n5681) );
  INV_X1 U6795 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n9192) );
  NOR2_X1 U6796 ( .A1(n5681), .A2(n9017), .ZN(n10505) );
  NAND2_X1 U6797 ( .A1(n10494), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n5682) );
  OAI21_X1 U6798 ( .B1(n10494), .B2(P2_REG2_REG_18__SCAN_IN), .A(n5682), .ZN(
        n10504) );
  INV_X1 U6799 ( .A(n5682), .ZN(n5683) );
  INV_X1 U6800 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n5684) );
  MUX2_X1 U6801 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n5684), .S(n8479), .Z(n5726)
         );
  INV_X1 U6802 ( .A(n8480), .ZN(n5685) );
  INV_X1 U6803 ( .A(n10506), .ZN(n5686) );
  MUX2_X1 U6804 ( .A(P2_REG2_REG_17__SCAN_IN), .B(P2_REG1_REG_17__SCAN_IN), 
        .S(n8480), .Z(n5722) );
  XNOR2_X1 U6805 ( .A(n5722), .B(n9023), .ZN(n9025) );
  MUX2_X1 U6806 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n4928), .Z(n5721) );
  XNOR2_X1 U6807 ( .A(n5721), .B(n9012), .ZN(n9002) );
  MUX2_X1 U6808 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n8480), .Z(n5688) );
  INV_X1 U6809 ( .A(n5688), .ZN(n5687) );
  NAND2_X1 U6810 ( .A1(n8994), .A2(n5687), .ZN(n5720) );
  XNOR2_X1 U6811 ( .A(n5688), .B(n8994), .ZN(n8984) );
  MUX2_X1 U6812 ( .A(P2_REG2_REG_14__SCAN_IN), .B(P2_REG1_REG_14__SCAN_IN), 
        .S(n4928), .Z(n5689) );
  OR2_X1 U6813 ( .A1(n5689), .A2(n7337), .ZN(n5719) );
  INV_X1 U6814 ( .A(n7337), .ZN(n8976) );
  XNOR2_X1 U6815 ( .A(n5689), .B(n8976), .ZN(n8965) );
  MUX2_X1 U6816 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n8480), .Z(n5690) );
  OR2_X1 U6817 ( .A1(n5690), .A2(n7314), .ZN(n5718) );
  XNOR2_X1 U6818 ( .A(n5690), .B(n8958), .ZN(n8948) );
  MUX2_X1 U6819 ( .A(P2_REG2_REG_12__SCAN_IN), .B(P2_REG1_REG_12__SCAN_IN), 
        .S(n8480), .Z(n5692) );
  INV_X1 U6820 ( .A(n5692), .ZN(n5691) );
  NAND2_X1 U6821 ( .A1(n8180), .A2(n5691), .ZN(n5717) );
  XNOR2_X1 U6822 ( .A(n5692), .B(n8180), .ZN(n8170) );
  MUX2_X1 U6823 ( .A(P2_REG2_REG_11__SCAN_IN), .B(P2_REG1_REG_11__SCAN_IN), 
        .S(n4928), .Z(n5715) );
  INV_X1 U6824 ( .A(n5715), .ZN(n5693) );
  NAND2_X1 U6825 ( .A1(n8069), .A2(n5693), .ZN(n5716) );
  MUX2_X1 U6826 ( .A(P2_REG2_REG_9__SCAN_IN), .B(P2_REG1_REG_9__SCAN_IN), .S(
        n4928), .Z(n5710) );
  NOR2_X1 U6827 ( .A1(n5710), .A2(n7202), .ZN(n5713) );
  MUX2_X1 U6828 ( .A(P2_REG2_REG_8__SCAN_IN), .B(P2_REG1_REG_8__SCAN_IN), .S(
        n8480), .Z(n5708) );
  NOR2_X1 U6829 ( .A1(n5708), .A2(n7154), .ZN(n5709) );
  MUX2_X1 U6830 ( .A(P2_REG2_REG_7__SCAN_IN), .B(P2_REG1_REG_7__SCAN_IN), .S(
        n4928), .Z(n5707) );
  MUX2_X1 U6831 ( .A(P2_REG2_REG_6__SCAN_IN), .B(P2_REG1_REG_6__SCAN_IN), .S(
        n8480), .Z(n5706) );
  MUX2_X1 U6832 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n8480), .Z(n5694) );
  INV_X1 U6833 ( .A(n5694), .ZN(n5704) );
  XNOR2_X1 U6834 ( .A(n5694), .B(n5810), .ZN(n10411) );
  MUX2_X1 U6835 ( .A(n7328), .B(n10581), .S(n4928), .Z(n5703) );
  XNOR2_X1 U6836 ( .A(n5703), .B(n5794), .ZN(n7323) );
  INV_X1 U6837 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n5766) );
  MUX2_X1 U6838 ( .A(n5656), .B(n5766), .S(n8480), .Z(n5700) );
  INV_X1 U6839 ( .A(n5700), .ZN(n5695) );
  NAND2_X1 U6840 ( .A1(n5695), .A2(n4925), .ZN(n5702) );
  MUX2_X1 U6841 ( .A(P2_REG2_REG_1__SCAN_IN), .B(P2_REG1_REG_1__SCAN_IN), .S(
        n8480), .Z(n5698) );
  INV_X1 U6842 ( .A(n5696), .ZN(n7285) );
  XNOR2_X1 U6843 ( .A(n5698), .B(n5696), .ZN(n7275) );
  MUX2_X1 U6844 ( .A(P2_REG2_REG_0__SCAN_IN), .B(P2_REG1_REG_0__SCAN_IN), .S(
        n4928), .Z(n5697) );
  NOR2_X1 U6845 ( .A1(n5697), .A2(n5265), .ZN(n7274) );
  INV_X1 U6846 ( .A(n5698), .ZN(n5699) );
  OAI22_X1 U6847 ( .A1(n7275), .A2(n7274), .B1(n7285), .B2(n5699), .ZN(n7288)
         );
  XNOR2_X1 U6848 ( .A(n5700), .B(n4925), .ZN(n7287) );
  NAND2_X1 U6849 ( .A1(n7288), .A2(n7287), .ZN(n5701) );
  NAND2_X1 U6850 ( .A1(n5702), .A2(n5701), .ZN(n7322) );
  NOR2_X1 U6851 ( .A1(n7323), .A2(n7322), .ZN(n7321) );
  AOI21_X1 U6852 ( .B1(n5703), .B2(n5794), .A(n7321), .ZN(n10410) );
  NAND2_X1 U6853 ( .A1(n10411), .A2(n10410), .ZN(n10409) );
  OAI21_X1 U6854 ( .B1(n5810), .B2(n5704), .A(n10409), .ZN(n10428) );
  MUX2_X1 U6855 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n4928), .Z(n5705) );
  XNOR2_X1 U6856 ( .A(n5705), .B(n10418), .ZN(n10427) );
  AOI22_X1 U6857 ( .A1(n10428), .A2(n10427), .B1(n5705), .B2(n7118), .ZN(
        n10440) );
  XNOR2_X1 U6858 ( .A(n5706), .B(n5844), .ZN(n10439) );
  NAND2_X1 U6859 ( .A1(n10440), .A2(n10439), .ZN(n10438) );
  OAI21_X1 U6860 ( .B1(n5706), .B2(n10435), .A(n10438), .ZN(n10464) );
  XNOR2_X1 U6861 ( .A(n5707), .B(n10453), .ZN(n10463) );
  NAND2_X1 U6862 ( .A1(n10464), .A2(n10463), .ZN(n10462) );
  OAI21_X1 U6863 ( .B1(n5707), .B2(n7145), .A(n10462), .ZN(n10484) );
  AOI21_X1 U6864 ( .B1(n5708), .B2(n7154), .A(n5709), .ZN(n10483) );
  AND2_X1 U6865 ( .A1(n10484), .A2(n10483), .ZN(n10486) );
  NOR2_X1 U6866 ( .A1(n5709), .A2(n10486), .ZN(n7870) );
  INV_X1 U6867 ( .A(n5710), .ZN(n5712) );
  INV_X1 U6868 ( .A(n5713), .ZN(n5711) );
  OAI21_X1 U6869 ( .B1(n7881), .B2(n5712), .A(n5711), .ZN(n7871) );
  NOR2_X1 U6870 ( .A1(n7870), .A2(n7871), .ZN(n7869) );
  NOR2_X1 U6871 ( .A1(n5713), .A2(n7869), .ZN(n7912) );
  MUX2_X1 U6872 ( .A(n5670), .B(n10691), .S(n8480), .Z(n5714) );
  NAND2_X1 U6873 ( .A1(n5714), .A2(n7908), .ZN(n7909) );
  NOR2_X1 U6874 ( .A1(n5714), .A2(n7908), .ZN(n7911) );
  AOI21_X1 U6875 ( .B1(n7912), .B2(n7909), .A(n7911), .ZN(n8060) );
  XNOR2_X1 U6876 ( .A(n5715), .B(n8069), .ZN(n8059) );
  NAND2_X1 U6877 ( .A1(n8060), .A2(n8059), .ZN(n8058) );
  NAND2_X1 U6878 ( .A1(n5716), .A2(n8058), .ZN(n8169) );
  NAND2_X1 U6879 ( .A1(n8170), .A2(n8169), .ZN(n8168) );
  NAND2_X1 U6880 ( .A1(n5717), .A2(n8168), .ZN(n8947) );
  NAND2_X1 U6881 ( .A1(n8948), .A2(n8947), .ZN(n8946) );
  NAND2_X1 U6882 ( .A1(n5718), .A2(n8946), .ZN(n8964) );
  NAND2_X1 U6883 ( .A1(n8965), .A2(n8964), .ZN(n8963) );
  NAND2_X1 U6884 ( .A1(n5719), .A2(n8963), .ZN(n8983) );
  NAND2_X1 U6885 ( .A1(n8984), .A2(n8983), .ZN(n8982) );
  NAND2_X1 U6886 ( .A1(n5720), .A2(n8982), .ZN(n9001) );
  NAND2_X1 U6887 ( .A1(n9002), .A2(n9001), .ZN(n9000) );
  OAI21_X1 U6888 ( .B1(n5721), .B2(n7610), .A(n9000), .ZN(n9024) );
  INV_X1 U6889 ( .A(n5722), .ZN(n5723) );
  AOI22_X1 U6890 ( .A1(n9025), .A2(n9024), .B1(n9023), .B2(n5723), .ZN(n5725)
         );
  MUX2_X1 U6891 ( .A(P2_REG2_REG_18__SCAN_IN), .B(P2_REG1_REG_18__SCAN_IN), 
        .S(n4928), .Z(n5724) );
  NOR2_X1 U6892 ( .A1(n5725), .A2(n5724), .ZN(n10491) );
  NAND2_X1 U6893 ( .A1(n5725), .A2(n5724), .ZN(n10492) );
  OAI21_X1 U6894 ( .B1(n10491), .B2(n10510), .A(n10492), .ZN(n5728) );
  MUX2_X1 U6895 ( .A(n5726), .B(n5024), .S(n4928), .Z(n5727) );
  NOR2_X1 U6896 ( .A1(n4928), .A2(P2_U3151), .ZN(n8249) );
  NAND2_X1 U6897 ( .A1(n5729), .A2(n8249), .ZN(n5730) );
  INV_X1 U6898 ( .A(n5648), .ZN(n8481) );
  MUX2_X1 U6899 ( .A(n5730), .B(n10508), .S(n8481), .Z(n10507) );
  INV_X1 U6900 ( .A(n8479), .ZN(n7833) );
  INV_X1 U6901 ( .A(n7443), .ZN(n8050) );
  NOR2_X1 U6902 ( .A1(n7444), .A2(n8050), .ZN(n5731) );
  INV_X1 U6903 ( .A(n10489), .ZN(n10498) );
  NAND2_X1 U6904 ( .A1(n10498), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n5732) );
  NAND2_X1 U6905 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8823) );
  OAI211_X1 U6906 ( .C1(n10507), .C2(n7833), .A(n5732), .B(n8823), .ZN(n5733)
         );
  INV_X1 U6907 ( .A(n5733), .ZN(n5734) );
  NAND3_X1 U6908 ( .A1(n5738), .A2(n5737), .A3(n5736), .ZN(P2_U3201) );
  INV_X1 U6909 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n7698) );
  OR2_X1 U6910 ( .A1(n6208), .A2(n7698), .ZN(n5749) );
  INV_X1 U6911 ( .A(n5744), .ZN(n9339) );
  OR2_X1 U6912 ( .A1(n4933), .A2(n7271), .ZN(n5748) );
  NAND2_X1 U6913 ( .A1(n5798), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5747) );
  INV_X1 U6914 ( .A(n5745), .ZN(n9341) );
  NAND2_X1 U6915 ( .A1(n8416), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5750) );
  INV_X1 U6916 ( .A(SI_1_), .ZN(n10066) );
  INV_X1 U6917 ( .A(n8416), .ZN(n5778) );
  AND2_X1 U6918 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5752) );
  NAND2_X1 U6919 ( .A1(n5778), .A2(n5752), .ZN(n6349) );
  AND2_X1 U6920 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n5753) );
  NAND2_X1 U6921 ( .A1(n8416), .A2(n5753), .ZN(n5763) );
  NAND2_X1 U6922 ( .A1(n6349), .A2(n5763), .ZN(n5771) );
  XNOR2_X1 U6923 ( .A(n5772), .B(n5771), .ZN(n7106) );
  INV_X1 U6924 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n7105) );
  OR2_X1 U6925 ( .A1(n5765), .A2(n5696), .ZN(n5754) );
  INV_X1 U6926 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n10198) );
  OR2_X1 U6927 ( .A1(n4929), .A2(n10198), .ZN(n5760) );
  INV_X1 U6928 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n7256) );
  OR2_X1 U6929 ( .A1(n5857), .A2(n7256), .ZN(n5758) );
  NAND2_X1 U6930 ( .A1(n4932), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5757) );
  NAND2_X1 U6931 ( .A1(n8416), .A2(SI_0_), .ZN(n5762) );
  INV_X1 U6932 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5761) );
  NAND2_X1 U6933 ( .A1(n5762), .A2(n5761), .ZN(n5764) );
  NAND2_X1 U6934 ( .A1(n5764), .A2(n5763), .ZN(n9347) );
  MUX2_X1 U6935 ( .A(n5265), .B(n9347), .S(n5765), .Z(n7499) );
  INV_X1 U6936 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n7300) );
  OR2_X1 U6937 ( .A1(n4929), .A2(n7300), .ZN(n5770) );
  NAND2_X1 U6938 ( .A1(n5798), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5769) );
  OR2_X1 U6939 ( .A1(n4933), .A2(n5656), .ZN(n5768) );
  NAND2_X1 U6940 ( .A1(n5772), .A2(n5771), .ZN(n5775) );
  NAND2_X1 U6941 ( .A1(n5773), .A2(SI_1_), .ZN(n5774) );
  NAND2_X1 U6942 ( .A1(n5775), .A2(n5774), .ZN(n5787) );
  NAND2_X1 U6943 ( .A1(n5778), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5776) );
  INV_X1 U6944 ( .A(SI_2_), .ZN(n5779) );
  XNOR2_X1 U6945 ( .A(n5788), .B(n5779), .ZN(n5786) );
  XNOR2_X1 U6946 ( .A(n5787), .B(n5786), .ZN(n7108) );
  INV_X1 U6947 ( .A(n8263), .ZN(n7766) );
  INV_X1 U6948 ( .A(n8941), .ZN(n7614) );
  NOR2_X1 U6949 ( .A1(n8941), .A2(n8266), .ZN(n5780) );
  NAND2_X1 U6950 ( .A1(n4932), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5784) );
  OR2_X1 U6951 ( .A1(n4929), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5783) );
  NAND2_X1 U6952 ( .A1(n5787), .A2(n5786), .ZN(n5790) );
  NAND2_X1 U6953 ( .A1(n5788), .A2(SI_2_), .ZN(n5789) );
  INV_X1 U6954 ( .A(SI_3_), .ZN(n10062) );
  XNOR2_X1 U6955 ( .A(n5806), .B(n10062), .ZN(n5804) );
  XNOR2_X1 U6956 ( .A(n5805), .B(n5804), .ZN(n7113) );
  OR2_X1 U6957 ( .A1(n5785), .A2(n7113), .ZN(n5797) );
  OR2_X1 U6958 ( .A1(n5793), .A2(n5792), .ZN(n5796) );
  NAND2_X1 U6959 ( .A1(n6051), .A2(n5794), .ZN(n5795) );
  OR2_X1 U6960 ( .A1(n8940), .A2(n10577), .ZN(n8275) );
  NAND2_X1 U6961 ( .A1(n8940), .A2(n10577), .ZN(n8294) );
  NAND2_X1 U6962 ( .A1(n8275), .A2(n8294), .ZN(n8446) );
  INV_X1 U6963 ( .A(n8446), .ZN(n7784) );
  NAND2_X1 U6964 ( .A1(n7785), .A2(n7784), .ZN(n7783) );
  NAND2_X1 U6965 ( .A1(n7783), .A2(n8275), .ZN(n7774) );
  NAND2_X1 U6966 ( .A1(n4932), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5803) );
  OR2_X1 U6967 ( .A1(n8424), .A2(n10589), .ZN(n5802) );
  NOR2_X1 U6968 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5815) );
  AND2_X1 U6969 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5799) );
  NOR2_X1 U6970 ( .A1(n5815), .A2(n5799), .ZN(n7454) );
  OR2_X1 U6971 ( .A1(n4929), .A2(n7454), .ZN(n5801) );
  NAND2_X1 U6972 ( .A1(n5805), .A2(n5804), .ZN(n5808) );
  NAND2_X1 U6973 ( .A1(n5806), .A2(SI_3_), .ZN(n5807) );
  MUX2_X1 U6974 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n7103), .Z(n5824) );
  INV_X1 U6975 ( .A(SI_4_), .ZN(n5809) );
  XNOR2_X1 U6976 ( .A(n5824), .B(n5809), .ZN(n5822) );
  XNOR2_X1 U6977 ( .A(n5823), .B(n5822), .ZN(n7111) );
  OR2_X1 U6978 ( .A1(n5785), .A2(n7111), .ZN(n5813) );
  INV_X1 U6979 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n7110) );
  OR2_X1 U6980 ( .A1(n5793), .A2(n7110), .ZN(n5812) );
  NAND2_X1 U6981 ( .A1(n6051), .A2(n5810), .ZN(n5811) );
  NAND2_X1 U6982 ( .A1(n8939), .A2(n7413), .ZN(n8276) );
  NAND2_X1 U6983 ( .A1(n7774), .A2(n8276), .ZN(n5814) );
  OR2_X1 U6984 ( .A1(n8939), .A2(n7413), .ZN(n8295) );
  NAND2_X1 U6985 ( .A1(n5814), .A2(n8295), .ZN(n8008) );
  INV_X1 U6986 ( .A(n8008), .ZN(n5831) );
  NAND2_X1 U6987 ( .A1(n4932), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5821) );
  OR2_X1 U6988 ( .A1(n8424), .A2(n10605), .ZN(n5820) );
  NAND2_X1 U6989 ( .A1(n5815), .A2(n5816), .ZN(n5833) );
  OR2_X1 U6990 ( .A1(n5816), .A2(n5815), .ZN(n5817) );
  AND2_X1 U6991 ( .A1(n5833), .A2(n5817), .ZN(n8004) );
  OR2_X1 U6992 ( .A1(n4929), .A2(n8004), .ZN(n5819) );
  OR2_X1 U6993 ( .A1(n5857), .A2(n10421), .ZN(n5818) );
  NAND4_X1 U6994 ( .A1(n5821), .A2(n5820), .A3(n5819), .A4(n5818), .ZN(n8938)
         );
  NAND2_X1 U6995 ( .A1(n5823), .A2(n5822), .ZN(n5826) );
  NAND2_X1 U6996 ( .A1(n5824), .A2(SI_4_), .ZN(n5825) );
  MUX2_X1 U6997 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n7103), .Z(n5841) );
  XNOR2_X1 U6998 ( .A(n5840), .B(SI_5_), .ZN(n7114) );
  INV_X2 U6999 ( .A(n5785), .ZN(n5981) );
  NAND2_X1 U7000 ( .A1(n7114), .A2(n5981), .ZN(n5829) );
  INV_X2 U7001 ( .A(n5793), .ZN(n6072) );
  NAND2_X1 U7002 ( .A1(n6072), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n5828) );
  NAND2_X1 U7003 ( .A1(n6051), .A2(n10418), .ZN(n5827) );
  OR2_X1 U7004 ( .A1(n8938), .A2(n10600), .ZN(n8296) );
  NAND2_X1 U7005 ( .A1(n8938), .A2(n10600), .ZN(n7663) );
  NAND2_X1 U7006 ( .A1(n8296), .A2(n7663), .ZN(n8448) );
  NAND2_X1 U7007 ( .A1(n5831), .A2(n5830), .ZN(n7662) );
  NAND2_X1 U7008 ( .A1(n4932), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5838) );
  OR2_X1 U7009 ( .A1(n8424), .A2(n5832), .ZN(n5837) );
  NAND2_X1 U7010 ( .A1(n5833), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5834) );
  AND2_X1 U7011 ( .A1(n5855), .A2(n5834), .ZN(n7714) );
  OR2_X1 U7012 ( .A1(n4929), .A2(n7714), .ZN(n5836) );
  OR2_X1 U7013 ( .A1(n5857), .A2(n5665), .ZN(n5835) );
  NAND4_X1 U7014 ( .A1(n5838), .A2(n5837), .A3(n5836), .A4(n5835), .ZN(n8937)
         );
  INV_X1 U7015 ( .A(SI_5_), .ZN(n5839) );
  NAND2_X1 U7016 ( .A1(n5842), .A2(n5841), .ZN(n5843) );
  MUX2_X1 U7017 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n7103), .Z(n5850) );
  XNOR2_X1 U7018 ( .A(n5850), .B(SI_6_), .ZN(n5848) );
  XNOR2_X1 U7019 ( .A(n5849), .B(n5848), .ZN(n7119) );
  NAND2_X1 U7020 ( .A1(n7119), .A2(n5981), .ZN(n5846) );
  AOI22_X1 U7021 ( .A1(n6072), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n6051), .B2(
        n5844), .ZN(n5845) );
  NAND2_X1 U7022 ( .A1(n8937), .A2(n7715), .ZN(n8278) );
  AND2_X1 U7023 ( .A1(n8278), .A2(n7663), .ZN(n8299) );
  NAND2_X1 U7024 ( .A1(n7662), .A2(n8299), .ZN(n5847) );
  NAND2_X1 U7025 ( .A1(n5850), .A2(SI_6_), .ZN(n5851) );
  MUX2_X1 U7026 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n7103), .Z(n5865) );
  XNOR2_X1 U7027 ( .A(n5865), .B(SI_7_), .ZN(n5862) );
  XNOR2_X1 U7028 ( .A(n5864), .B(n5862), .ZN(n7139) );
  NAND2_X1 U7029 ( .A1(n7139), .A2(n5981), .ZN(n5854) );
  AOI22_X1 U7030 ( .A1(n6072), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n6051), .B2(
        n10453), .ZN(n5853) );
  NAND2_X1 U7031 ( .A1(n4932), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5861) );
  OR2_X1 U7032 ( .A1(n8424), .A2(n10626), .ZN(n5860) );
  AND2_X1 U7033 ( .A1(n5855), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5856) );
  NOR2_X1 U7034 ( .A1(n5873), .A2(n5856), .ZN(n7893) );
  OR2_X1 U7035 ( .A1(n4929), .A2(n7893), .ZN(n5859) );
  OR2_X1 U7036 ( .A1(n5857), .A2(n10456), .ZN(n5858) );
  NAND2_X1 U7037 ( .A1(n10619), .A2(n7750), .ZN(n8286) );
  INV_X1 U7038 ( .A(n8282), .ZN(n8453) );
  INV_X1 U7039 ( .A(n5862), .ZN(n5863) );
  NAND2_X1 U7040 ( .A1(n5865), .A2(SI_7_), .ZN(n5866) );
  MUX2_X1 U7041 ( .A(n7152), .B(n7208), .S(n7103), .Z(n5868) );
  INV_X1 U7042 ( .A(SI_8_), .ZN(n5867) );
  NAND2_X1 U7043 ( .A1(n5868), .A2(n5867), .ZN(n5881) );
  INV_X1 U7044 ( .A(n5868), .ZN(n5869) );
  NAND2_X1 U7045 ( .A1(n5869), .A2(SI_8_), .ZN(n5870) );
  NAND2_X1 U7046 ( .A1(n5881), .A2(n5870), .ZN(n5882) );
  AOI22_X1 U7047 ( .A1(n6072), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6051), .B2(
        n10473), .ZN(n5871) );
  NAND2_X1 U7048 ( .A1(n4932), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5878) );
  OR2_X1 U7049 ( .A1(n8424), .A2(n5613), .ZN(n5877) );
  NOR2_X1 U7050 ( .A1(n5873), .A2(n5872), .ZN(n5874) );
  OR2_X1 U7051 ( .A1(n4929), .A2(n5525), .ZN(n5876) );
  OR2_X1 U7052 ( .A1(n5857), .A2(n10646), .ZN(n5875) );
  OR2_X1 U7053 ( .A1(n10642), .A2(n8031), .ZN(n8283) );
  NAND2_X1 U7054 ( .A1(n8283), .A2(n7810), .ZN(n8310) );
  INV_X1 U7055 ( .A(n8310), .ZN(n5879) );
  NAND2_X1 U7056 ( .A1(n10642), .A2(n8031), .ZN(n8287) );
  NAND2_X1 U7057 ( .A1(n5880), .A2(n8287), .ZN(n8029) );
  MUX2_X1 U7058 ( .A(n7200), .B(n7210), .S(n7103), .Z(n5884) );
  NAND2_X1 U7059 ( .A1(n5884), .A2(n10146), .ZN(n5897) );
  INV_X1 U7060 ( .A(n5884), .ZN(n5885) );
  NAND2_X1 U7061 ( .A1(n5885), .A2(SI_9_), .ZN(n5886) );
  NAND2_X1 U7062 ( .A1(n6461), .A2(n5981), .ZN(n5888) );
  AOI22_X1 U7063 ( .A1(n6072), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6051), .B2(
        n7881), .ZN(n5887) );
  NAND2_X1 U7064 ( .A1(n4932), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5894) );
  OR2_X1 U7065 ( .A1(n8424), .A2(n10665), .ZN(n5893) );
  OR2_X1 U7066 ( .A1(n5889), .A2(n10195), .ZN(n5890) );
  AND2_X1 U7067 ( .A1(n5901), .A2(n5890), .ZN(n8033) );
  OR2_X1 U7068 ( .A1(n4929), .A2(n8033), .ZN(n5892) );
  OR2_X1 U7069 ( .A1(n5857), .A2(n8034), .ZN(n5891) );
  NAND2_X1 U7070 ( .A1(n5895), .A2(n8042), .ZN(n8288) );
  NAND2_X1 U7071 ( .A1(n8284), .A2(n8288), .ZN(n8454) );
  MUX2_X1 U7072 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .S(n7103), .Z(n5911) );
  INV_X1 U7073 ( .A(SI_10_), .ZN(n5898) );
  XNOR2_X1 U7074 ( .A(n5911), .B(n5898), .ZN(n5908) );
  XNOR2_X1 U7075 ( .A(n5910), .B(n5908), .ZN(n7203) );
  NAND2_X1 U7076 ( .A1(n7203), .A2(n5981), .ZN(n5900) );
  AOI22_X1 U7077 ( .A1(n6072), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6051), .B2(
        n7908), .ZN(n5899) );
  NAND2_X1 U7078 ( .A1(n5900), .A2(n5899), .ZN(n10685) );
  NAND2_X1 U7079 ( .A1(n4932), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5906) );
  OR2_X1 U7080 ( .A1(n8424), .A2(n10691), .ZN(n5905) );
  OR2_X2 U7081 ( .A1(n5901), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5920) );
  NAND2_X1 U7082 ( .A1(n5901), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5902) );
  AND2_X1 U7083 ( .A1(n5920), .A2(n5902), .ZN(n8044) );
  OR2_X1 U7084 ( .A1(n4929), .A2(n8044), .ZN(n5904) );
  OR2_X1 U7085 ( .A1(n5857), .A2(n5670), .ZN(n5903) );
  OR2_X1 U7086 ( .A1(n10685), .A2(n8035), .ZN(n8305) );
  NAND2_X1 U7087 ( .A1(n8305), .A2(n8284), .ZN(n8309) );
  INV_X1 U7088 ( .A(n8309), .ZN(n5907) );
  NAND2_X1 U7089 ( .A1(n10685), .A2(n8035), .ZN(n8314) );
  INV_X1 U7090 ( .A(n5908), .ZN(n5909) );
  NAND2_X1 U7091 ( .A1(n5911), .A2(SI_10_), .ZN(n5912) );
  INV_X1 U7092 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n5913) );
  MUX2_X1 U7093 ( .A(n5913), .B(n7223), .S(n7103), .Z(n5915) );
  INV_X1 U7094 ( .A(SI_11_), .ZN(n5914) );
  NAND2_X1 U7095 ( .A1(n5915), .A2(n5914), .ZN(n5926) );
  INV_X1 U7096 ( .A(n5915), .ZN(n5916) );
  NAND2_X1 U7097 ( .A1(n5916), .A2(SI_11_), .ZN(n5917) );
  NAND2_X1 U7098 ( .A1(n5926), .A2(n5917), .ZN(n5927) );
  NAND2_X1 U7099 ( .A1(n7219), .A2(n5981), .ZN(n5919) );
  AOI22_X1 U7100 ( .A1(n6072), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6051), .B2(
        n8069), .ZN(n5918) );
  NAND2_X1 U7101 ( .A1(n5919), .A2(n5918), .ZN(n10695) );
  NAND2_X1 U7102 ( .A1(n4932), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5925) );
  OR2_X1 U7103 ( .A1(n5857), .A2(n8056), .ZN(n5924) );
  NOR2_X2 U7104 ( .A1(n5920), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5933) );
  AND2_X1 U7105 ( .A1(n5920), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5921) );
  NOR2_X1 U7106 ( .A1(n5933), .A2(n5921), .ZN(n8107) );
  OR2_X1 U7107 ( .A1(n4929), .A2(n8107), .ZN(n5923) );
  OR2_X1 U7108 ( .A1(n8424), .A2(n10701), .ZN(n5922) );
  OR2_X1 U7109 ( .A1(n10695), .A2(n10686), .ZN(n8316) );
  NAND2_X1 U7110 ( .A1(n10695), .A2(n10686), .ZN(n8318) );
  MUX2_X1 U7111 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .S(n5046), .Z(n5943) );
  XNOR2_X1 U7112 ( .A(n5943), .B(n10048), .ZN(n5942) );
  XNOR2_X1 U7113 ( .A(n5946), .B(n5942), .ZN(n7263) );
  NAND2_X1 U7114 ( .A1(n7263), .A2(n5981), .ZN(n5930) );
  AOI22_X1 U7115 ( .A1(n6072), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6051), .B2(
        n8180), .ZN(n5929) );
  NAND2_X1 U7116 ( .A1(n5930), .A2(n5929), .ZN(n10708) );
  NAND2_X1 U7117 ( .A1(n4930), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5939) );
  INV_X1 U7118 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n5931) );
  OR2_X1 U7119 ( .A1(n8426), .A2(n5931), .ZN(n5938) );
  OR2_X1 U7120 ( .A1(n5933), .A2(n5932), .ZN(n5934) );
  AND2_X1 U7121 ( .A1(n5949), .A2(n5934), .ZN(n8075) );
  OR2_X1 U7122 ( .A1(n4929), .A2(n8075), .ZN(n5937) );
  OR2_X1 U7123 ( .A1(n5857), .A2(n5935), .ZN(n5936) );
  NAND4_X1 U7124 ( .A1(n5939), .A2(n5938), .A3(n5937), .A4(n5936), .ZN(n8935)
         );
  INV_X1 U7125 ( .A(n8935), .ZN(n10696) );
  NAND2_X1 U7126 ( .A1(n8076), .A2(n4955), .ZN(n5941) );
  AND2_X1 U7127 ( .A1(n10708), .A2(n10696), .ZN(n8307) );
  INV_X1 U7128 ( .A(n8307), .ZN(n5940) );
  NAND2_X1 U7129 ( .A1(n5941), .A2(n5940), .ZN(n7990) );
  INV_X1 U7130 ( .A(n5942), .ZN(n5945) );
  NAND2_X1 U7131 ( .A1(n5943), .A2(SI_12_), .ZN(n5944) );
  MUX2_X1 U7132 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n5046), .Z(n5960) );
  XNOR2_X1 U7133 ( .A(n5960), .B(SI_13_), .ZN(n5957) );
  XNOR2_X1 U7134 ( .A(n5959), .B(n5957), .ZN(n7267) );
  NAND2_X1 U7135 ( .A1(n7267), .A2(n5981), .ZN(n5948) );
  AOI22_X1 U7136 ( .A1(n6072), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6051), .B2(
        n8958), .ZN(n5947) );
  NAND2_X1 U7137 ( .A1(n5948), .A2(n5947), .ZN(n10714) );
  NAND2_X1 U7138 ( .A1(n4932), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5953) );
  OR2_X1 U7139 ( .A1(n8424), .A2(n10715), .ZN(n5952) );
  AOI21_X1 U7140 ( .B1(n5949), .B2(P2_REG3_REG_13__SCAN_IN), .A(n5971), .ZN(
        n8157) );
  OR2_X1 U7141 ( .A1(n4929), .A2(n8157), .ZN(n5951) );
  OR2_X1 U7142 ( .A1(n5857), .A2(n8944), .ZN(n5950) );
  NOR2_X1 U7143 ( .A1(n10714), .A2(n9235), .ZN(n8322) );
  INV_X1 U7144 ( .A(n8322), .ZN(n5954) );
  AND2_X1 U7145 ( .A1(n10714), .A2(n9235), .ZN(n8323) );
  INV_X1 U7146 ( .A(n8323), .ZN(n5955) );
  NAND2_X1 U7147 ( .A1(n7990), .A2(n8325), .ZN(n5956) );
  NAND2_X1 U7148 ( .A1(n5956), .A2(n5955), .ZN(n9244) );
  INV_X1 U7149 ( .A(n5957), .ZN(n5958) );
  NAND2_X1 U7150 ( .A1(n5959), .A2(n5958), .ZN(n5962) );
  NAND2_X1 U7151 ( .A1(n5960), .A2(SI_13_), .ZN(n5961) );
  NAND2_X1 U7152 ( .A1(n5962), .A2(n5961), .ZN(n5980) );
  MUX2_X1 U7153 ( .A(n7335), .B(n5963), .S(n5046), .Z(n5964) );
  NAND2_X1 U7154 ( .A1(n5964), .A2(n10139), .ZN(n5978) );
  INV_X1 U7155 ( .A(n5964), .ZN(n5965) );
  NAND2_X1 U7156 ( .A1(n5965), .A2(SI_14_), .ZN(n5966) );
  NAND2_X1 U7157 ( .A1(n5978), .A2(n5966), .ZN(n5979) );
  XNOR2_X1 U7158 ( .A(n5980), .B(n5979), .ZN(n7316) );
  NAND2_X1 U7159 ( .A1(n7316), .A2(n5981), .ZN(n5968) );
  AOI22_X1 U7160 ( .A1(n6072), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6051), .B2(
        n8976), .ZN(n5967) );
  NAND2_X1 U7161 ( .A1(n5968), .A2(n5967), .ZN(n8328) );
  NAND2_X1 U7162 ( .A1(n4932), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5976) );
  INV_X1 U7163 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n5969) );
  OR2_X1 U7164 ( .A1(n8424), .A2(n5969), .ZN(n5975) );
  INV_X1 U7165 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n5970) );
  OR2_X1 U7166 ( .A1(n5857), .A2(n5970), .ZN(n5974) );
  AOI21_X1 U7167 ( .B1(P2_REG3_REG_14__SCAN_IN), .B2(n5972), .A(n5984), .ZN(
        n9239) );
  OR2_X1 U7168 ( .A1(n4929), .A2(n9239), .ZN(n5973) );
  NAND4_X1 U7169 ( .A1(n5976), .A2(n5975), .A3(n5974), .A4(n5973), .ZN(n9215)
         );
  OR2_X1 U7170 ( .A1(n8328), .A2(n9215), .ZN(n6272) );
  NAND2_X1 U7171 ( .A1(n8328), .A2(n9215), .ZN(n8326) );
  NAND2_X1 U7172 ( .A1(n9244), .A2(n9243), .ZN(n9242) );
  INV_X1 U7173 ( .A(n9215), .ZN(n8758) );
  NAND2_X1 U7174 ( .A1(n8328), .A2(n8758), .ZN(n5977) );
  MUX2_X1 U7175 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n5046), .Z(n5992) );
  XNOR2_X1 U7176 ( .A(n5992), .B(n10042), .ZN(n5991) );
  NAND2_X1 U7177 ( .A1(n7402), .A2(n5981), .ZN(n5983) );
  AOI22_X1 U7178 ( .A1(n6072), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n6051), .B2(
        n8994), .ZN(n5982) );
  NAND2_X1 U7179 ( .A1(n4932), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5989) );
  AOI21_X1 U7180 ( .B1(P2_REG3_REG_15__SCAN_IN), .B2(n5985), .A(n6019), .ZN(
        n9220) );
  OR2_X1 U7181 ( .A1(n4929), .A2(n9220), .ZN(n5988) );
  OR2_X1 U7182 ( .A1(n8424), .A2(n10729), .ZN(n5987) );
  OR2_X1 U7183 ( .A1(n5857), .A2(n8980), .ZN(n5986) );
  NAND2_X1 U7184 ( .A1(n10725), .A2(n9237), .ZN(n8329) );
  INV_X1 U7185 ( .A(n8329), .ZN(n5990) );
  INV_X1 U7186 ( .A(n5991), .ZN(n5994) );
  NAND2_X1 U7187 ( .A1(n5992), .A2(SI_15_), .ZN(n5993) );
  MUX2_X1 U7188 ( .A(n7608), .B(n5996), .S(n5046), .Z(n5997) );
  NAND2_X1 U7189 ( .A1(n5997), .A2(n10140), .ZN(n6000) );
  INV_X1 U7190 ( .A(n5997), .ZN(n5998) );
  NAND2_X1 U7191 ( .A1(n5998), .A2(SI_16_), .ZN(n5999) );
  NAND2_X1 U7192 ( .A1(n6000), .A2(n5999), .ZN(n6013) );
  MUX2_X1 U7193 ( .A(n6002), .B(n6001), .S(n5046), .Z(n6003) );
  NAND2_X1 U7194 ( .A1(n6003), .A2(n10133), .ZN(n6033) );
  INV_X1 U7195 ( .A(n6003), .ZN(n6004) );
  NAND2_X1 U7196 ( .A1(n6004), .A2(SI_17_), .ZN(n6005) );
  XNOR2_X1 U7197 ( .A(n6032), .B(n6031), .ZN(n7629) );
  NAND2_X1 U7198 ( .A1(n7629), .A2(n5981), .ZN(n6007) );
  AOI22_X1 U7199 ( .A1(n6072), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n9023), .B2(
        n6051), .ZN(n6006) );
  NAND2_X1 U7200 ( .A1(n4932), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n6009) );
  NAND2_X1 U7201 ( .A1(n6038), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n6008) );
  OAI211_X1 U7202 ( .C1(n10746), .C2(n8424), .A(n6009), .B(n6008), .ZN(n6010)
         );
  INV_X1 U7203 ( .A(n6010), .ZN(n6012) );
  AOI21_X1 U7204 ( .B1(P2_REG3_REG_17__SCAN_IN), .B2(n6018), .A(n6037), .ZN(
        n9191) );
  OR2_X1 U7205 ( .A1(n9191), .A2(n4929), .ZN(n6011) );
  NOR2_X1 U7206 ( .A1(n8862), .A2(n9201), .ZN(n6025) );
  XNOR2_X1 U7207 ( .A(n6014), .B(n6013), .ZN(n7534) );
  NAND2_X1 U7208 ( .A1(n7534), .A2(n5981), .ZN(n6016) );
  AOI22_X1 U7209 ( .A1(n6072), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6051), .B2(
        n9012), .ZN(n6015) );
  NAND2_X1 U7210 ( .A1(n4932), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n6024) );
  OR2_X1 U7211 ( .A1(n5857), .A2(n6017), .ZN(n6023) );
  OR2_X1 U7212 ( .A1(n8424), .A2(n10736), .ZN(n6022) );
  OAI21_X1 U7213 ( .B1(n10090), .B2(n6019), .A(n6018), .ZN(n9204) );
  INV_X1 U7214 ( .A(n9204), .ZN(n6020) );
  OR2_X1 U7215 ( .A1(n4929), .A2(n6020), .ZN(n6021) );
  NOR2_X1 U7216 ( .A1(n8848), .A2(n8917), .ZN(n9188) );
  NAND2_X1 U7217 ( .A1(n8848), .A2(n8917), .ZN(n6026) );
  NAND2_X1 U7218 ( .A1(n6026), .A2(n8932), .ZN(n6028) );
  NOR2_X1 U7219 ( .A1(n8932), .A2(n9217), .ZN(n6027) );
  AOI22_X1 U7220 ( .A1(n8862), .A2(n6028), .B1(n6027), .B2(n8848), .ZN(n6029)
         );
  MUX2_X1 U7221 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n5046), .Z(n6045) );
  XNOR2_X1 U7222 ( .A(n6045), .B(n6034), .ZN(n6043) );
  XNOR2_X1 U7223 ( .A(n6044), .B(n6043), .ZN(n7703) );
  NAND2_X1 U7224 ( .A1(n7703), .A2(n5981), .ZN(n6036) );
  AOI22_X1 U7225 ( .A1(n6072), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6051), .B2(
        n10510), .ZN(n6035) );
  OAI21_X1 U7226 ( .B1(n8894), .B2(n6037), .A(n6054), .ZN(n9176) );
  INV_X1 U7227 ( .A(n4929), .ZN(n6056) );
  NAND2_X1 U7228 ( .A1(n9176), .A2(n6056), .ZN(n6042) );
  NAND2_X1 U7229 ( .A1(n4930), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n6041) );
  NAND2_X1 U7230 ( .A1(n4932), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n6040) );
  NAND2_X1 U7231 ( .A1(n6038), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n6039) );
  NAND2_X1 U7232 ( .A1(n10752), .A2(n10739), .ZN(n8343) );
  NAND2_X1 U7233 ( .A1(n8342), .A2(n8343), .ZN(n9181) );
  NAND2_X1 U7234 ( .A1(n6045), .A2(SI_18_), .ZN(n6064) );
  INV_X1 U7235 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n6046) );
  MUX2_X1 U7236 ( .A(n7831), .B(n6046), .S(n5046), .Z(n6047) );
  NAND2_X1 U7237 ( .A1(n6047), .A2(n10129), .ZN(n6066) );
  INV_X1 U7238 ( .A(n6047), .ZN(n6048) );
  NAND2_X1 U7239 ( .A1(n6048), .A2(SI_19_), .ZN(n6049) );
  NAND2_X1 U7240 ( .A1(n6066), .A2(n6049), .ZN(n6063) );
  XNOR2_X1 U7241 ( .A(n6050), .B(n6063), .ZN(n7772) );
  NAND2_X1 U7242 ( .A1(n7772), .A2(n5981), .ZN(n6053) );
  AOI22_X1 U7243 ( .A1(n6072), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n8479), .B2(
        n6051), .ZN(n6052) );
  NAND2_X1 U7244 ( .A1(n6054), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6055) );
  INV_X1 U7245 ( .A(n6076), .ZN(n6078) );
  NAND2_X1 U7246 ( .A1(n6055), .A2(n6078), .ZN(n9165) );
  NAND2_X1 U7247 ( .A1(n9165), .A2(n6056), .ZN(n6062) );
  INV_X1 U7248 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n6057) );
  OR2_X1 U7249 ( .A1(n8426), .A2(n6057), .ZN(n6059) );
  OR2_X1 U7250 ( .A1(n5857), .A2(n5684), .ZN(n6058) );
  AND2_X1 U7251 ( .A1(n6059), .A2(n6058), .ZN(n6061) );
  NAND2_X1 U7252 ( .A1(n4930), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n6060) );
  NAND2_X1 U7253 ( .A1(n9296), .A2(n10755), .ZN(n8349) );
  INV_X1 U7254 ( .A(n9159), .ZN(n9163) );
  NAND2_X1 U7255 ( .A1(n9164), .A2(n9163), .ZN(n9162) );
  INV_X1 U7256 ( .A(n6063), .ZN(n6065) );
  NAND2_X1 U7257 ( .A1(n6067), .A2(n6066), .ZN(n6085) );
  MUX2_X1 U7258 ( .A(n7865), .B(n6068), .S(n5046), .Z(n6069) );
  INV_X1 U7259 ( .A(SI_20_), .ZN(n10131) );
  NAND2_X1 U7260 ( .A1(n6069), .A2(n10131), .ZN(n6086) );
  INV_X1 U7261 ( .A(n6069), .ZN(n6070) );
  NAND2_X1 U7262 ( .A1(n6070), .A2(SI_20_), .ZN(n6071) );
  XNOR2_X1 U7263 ( .A(n6085), .B(n6084), .ZN(n7843) );
  NAND2_X1 U7264 ( .A1(n7843), .A2(n5981), .ZN(n6074) );
  NAND2_X1 U7265 ( .A1(n6072), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n6073) );
  NAND2_X1 U7266 ( .A1(n4930), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n6082) );
  INV_X1 U7267 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n6075) );
  OR2_X1 U7268 ( .A1(n8426), .A2(n6075), .ZN(n6081) );
  INV_X1 U7269 ( .A(n6090), .ZN(n6077) );
  AOI21_X1 U7270 ( .B1(P2_REG3_REG_20__SCAN_IN), .B2(n6078), .A(n6077), .ZN(
        n9151) );
  OR2_X1 U7271 ( .A1(n4929), .A2(n9151), .ZN(n6080) );
  INV_X1 U7272 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n9152) );
  OR2_X1 U7273 ( .A1(n5857), .A2(n9152), .ZN(n6079) );
  NAND4_X1 U7274 ( .A1(n6082), .A2(n6081), .A3(n6080), .A4(n6079), .ZN(n9295)
         );
  OR2_X1 U7275 ( .A1(n9331), .A2(n9295), .ZN(n6279) );
  NAND2_X1 U7276 ( .A1(n9331), .A2(n9295), .ZN(n6083) );
  INV_X1 U7277 ( .A(n9295), .ZN(n8825) );
  AND2_X1 U7278 ( .A1(n9331), .A2(n8825), .ZN(n8252) );
  MUX2_X1 U7279 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n5046), .Z(n6097) );
  XNOR2_X1 U7280 ( .A(n6097), .B(n6087), .ZN(n6096) );
  XNOR2_X1 U7281 ( .A(n6095), .B(n6096), .ZN(n7918) );
  NAND2_X1 U7282 ( .A1(n7918), .A2(n5981), .ZN(n6089) );
  NAND2_X1 U7283 ( .A1(n6072), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n6088) );
  NAND2_X1 U7284 ( .A1(n4930), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n6094) );
  INV_X1 U7285 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n9325) );
  OR2_X1 U7286 ( .A1(n8426), .A2(n9325), .ZN(n6093) );
  AOI21_X1 U7287 ( .B1(P2_REG3_REG_21__SCAN_IN), .B2(n6090), .A(n6106), .ZN(
        n9132) );
  OR2_X1 U7288 ( .A1(n4929), .A2(n9132), .ZN(n6092) );
  INV_X1 U7289 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n9133) );
  OR2_X1 U7290 ( .A1(n5857), .A2(n9133), .ZN(n6091) );
  INV_X1 U7291 ( .A(n9148), .ZN(n8930) );
  NAND2_X1 U7292 ( .A1(n9138), .A2(n8930), .ZN(n8357) );
  NAND2_X1 U7293 ( .A1(n8355), .A2(n8357), .ZN(n9134) );
  NAND2_X1 U7294 ( .A1(n6097), .A2(SI_21_), .ZN(n6098) );
  NAND2_X1 U7295 ( .A1(n6099), .A2(n6098), .ZN(n6119) );
  INV_X1 U7296 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n6100) );
  MUX2_X1 U7297 ( .A(n7946), .B(n6100), .S(n5046), .Z(n6101) );
  NAND2_X1 U7298 ( .A1(n6101), .A2(n10121), .ZN(n6117) );
  INV_X1 U7299 ( .A(n6101), .ZN(n6102) );
  NAND2_X1 U7300 ( .A1(n6102), .A2(SI_22_), .ZN(n6103) );
  NAND2_X1 U7301 ( .A1(n6117), .A2(n6103), .ZN(n6118) );
  XNOR2_X1 U7302 ( .A(n6119), .B(n6118), .ZN(n7943) );
  NAND2_X1 U7303 ( .A1(n7943), .A2(n5981), .ZN(n6105) );
  NAND2_X1 U7304 ( .A1(n6072), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n6104) );
  NAND2_X1 U7305 ( .A1(n4930), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n6112) );
  INV_X1 U7306 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n9321) );
  OR2_X1 U7307 ( .A1(n8426), .A2(n9321), .ZN(n6111) );
  NAND2_X1 U7308 ( .A1(n10205), .A2(n6106), .ZN(n6132) );
  INV_X1 U7309 ( .A(n6106), .ZN(n6107) );
  NAND2_X1 U7310 ( .A1(P2_REG3_REG_22__SCAN_IN), .A2(n6107), .ZN(n6108) );
  AND2_X1 U7311 ( .A1(n6132), .A2(n6108), .ZN(n9119) );
  OR2_X1 U7312 ( .A1(n4929), .A2(n9119), .ZN(n6110) );
  INV_X1 U7313 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n9120) );
  OR2_X1 U7314 ( .A1(n5857), .A2(n9120), .ZN(n6109) );
  AND2_X1 U7315 ( .A1(n8779), .A2(n8833), .ZN(n8361) );
  INV_X1 U7316 ( .A(n8361), .ZN(n6113) );
  AND2_X1 U7317 ( .A1(n9134), .A2(n6113), .ZN(n6114) );
  OR2_X1 U7318 ( .A1(n9138), .A2(n9148), .ZN(n9116) );
  NOR2_X1 U7319 ( .A1(n8779), .A2(n8833), .ZN(n8362) );
  INV_X1 U7320 ( .A(n8362), .ZN(n6115) );
  NAND2_X1 U7321 ( .A1(n6116), .A2(n6115), .ZN(n9105) );
  INV_X1 U7322 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n6121) );
  INV_X1 U7323 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n6120) );
  MUX2_X1 U7324 ( .A(n6121), .B(n6120), .S(n5046), .Z(n6123) );
  INV_X1 U7325 ( .A(SI_23_), .ZN(n6122) );
  NAND2_X1 U7326 ( .A1(n6123), .A2(n6122), .ZN(n6138) );
  INV_X1 U7327 ( .A(n6123), .ZN(n6124) );
  NAND2_X1 U7328 ( .A1(n6124), .A2(SI_23_), .ZN(n6125) );
  NAND2_X1 U7329 ( .A1(n6127), .A2(n6126), .ZN(n6139) );
  OAI21_X1 U7330 ( .B1(n6127), .B2(n6126), .A(n6139), .ZN(n8049) );
  NAND2_X1 U7331 ( .A1(n8049), .A2(n5981), .ZN(n6129) );
  NAND2_X1 U7332 ( .A1(n6072), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n6128) );
  NAND2_X1 U7333 ( .A1(n4930), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n6137) );
  INV_X1 U7334 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n6130) );
  OR2_X1 U7335 ( .A1(n8426), .A2(n6130), .ZN(n6136) );
  INV_X1 U7336 ( .A(n6132), .ZN(n6131) );
  INV_X1 U7337 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8814) );
  NAND2_X1 U7338 ( .A1(n6131), .A2(n8814), .ZN(n6150) );
  NAND2_X1 U7339 ( .A1(n6132), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6133) );
  AND2_X1 U7340 ( .A1(n6150), .A2(n6133), .ZN(n9107) );
  OR2_X1 U7341 ( .A1(n4929), .A2(n9107), .ZN(n6135) );
  INV_X1 U7342 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n9108) );
  OR2_X1 U7343 ( .A1(n5857), .A2(n9108), .ZN(n6134) );
  OR2_X1 U7344 ( .A1(n9273), .A2(n9114), .ZN(n8366) );
  NAND2_X1 U7345 ( .A1(n9273), .A2(n9114), .ZN(n8367) );
  NAND2_X1 U7346 ( .A1(n6139), .A2(n6138), .ZN(n6145) );
  INV_X1 U7347 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n6140) );
  MUX2_X1 U7348 ( .A(n8223), .B(n6140), .S(n5046), .Z(n6141) );
  INV_X1 U7349 ( .A(SI_24_), .ZN(n10120) );
  NAND2_X1 U7350 ( .A1(n6141), .A2(n10120), .ZN(n6159) );
  INV_X1 U7351 ( .A(n6141), .ZN(n6142) );
  NAND2_X1 U7352 ( .A1(n6142), .A2(SI_24_), .ZN(n6143) );
  OR2_X1 U7353 ( .A1(n6145), .A2(n6144), .ZN(n6146) );
  NAND2_X1 U7354 ( .A1(n6160), .A2(n6146), .ZN(n8111) );
  NAND2_X1 U7355 ( .A1(n8111), .A2(n5981), .ZN(n6148) );
  NAND2_X1 U7356 ( .A1(n6072), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n6147) );
  NAND2_X1 U7357 ( .A1(n4930), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n6156) );
  INV_X1 U7358 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n9316) );
  OR2_X1 U7359 ( .A1(n8426), .A2(n9316), .ZN(n6155) );
  INV_X1 U7360 ( .A(n6150), .ZN(n6149) );
  INV_X1 U7361 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n8867) );
  INV_X1 U7362 ( .A(n6167), .ZN(n6168) );
  NAND2_X1 U7363 ( .A1(n6150), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6151) );
  OR2_X1 U7364 ( .A1(n4929), .A2(n9094), .ZN(n6154) );
  INV_X1 U7365 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n6152) );
  OR2_X1 U7366 ( .A1(n5857), .A2(n6152), .ZN(n6153) );
  NOR2_X1 U7367 ( .A1(n9093), .A2(n9076), .ZN(n8371) );
  INV_X1 U7368 ( .A(n8371), .ZN(n6158) );
  AND2_X1 U7369 ( .A1(n9093), .A2(n9076), .ZN(n8372) );
  INV_X1 U7370 ( .A(n8372), .ZN(n6157) );
  NAND2_X1 U7371 ( .A1(n6158), .A2(n6157), .ZN(n9096) );
  INV_X1 U7372 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n6161) );
  MUX2_X1 U7373 ( .A(n8238), .B(n6161), .S(n5046), .Z(n6162) );
  NAND2_X1 U7374 ( .A1(n6162), .A2(n10123), .ZN(n6176) );
  INV_X1 U7375 ( .A(n6162), .ZN(n6163) );
  NAND2_X1 U7376 ( .A1(n6163), .A2(SI_25_), .ZN(n6164) );
  XNOR2_X1 U7377 ( .A(n6175), .B(n6174), .ZN(n8225) );
  NAND2_X1 U7378 ( .A1(n8225), .A2(n5981), .ZN(n6166) );
  NAND2_X1 U7379 ( .A1(n6072), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n6165) );
  NAND2_X1 U7380 ( .A1(n4930), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n6173) );
  INV_X1 U7381 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n9312) );
  OR2_X1 U7382 ( .A1(n8426), .A2(n9312), .ZN(n6172) );
  INV_X1 U7383 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n10184) );
  NAND2_X1 U7384 ( .A1(n6168), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6169) );
  AND2_X1 U7385 ( .A1(n6186), .A2(n6169), .ZN(n9082) );
  OR2_X1 U7386 ( .A1(n4929), .A2(n9082), .ZN(n6171) );
  INV_X1 U7387 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n9083) );
  OR2_X1 U7388 ( .A1(n5857), .A2(n9083), .ZN(n6170) );
  OR2_X1 U7389 ( .A1(n9078), .A2(n8868), .ZN(n8377) );
  NAND2_X1 U7390 ( .A1(n9078), .A2(n8868), .ZN(n8373) );
  INV_X1 U7391 ( .A(n8373), .ZN(n8378) );
  INV_X1 U7392 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n6178) );
  INV_X1 U7393 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n6177) );
  MUX2_X1 U7394 ( .A(n6178), .B(n6177), .S(n5046), .Z(n6180) );
  INV_X1 U7395 ( .A(SI_26_), .ZN(n6179) );
  NAND2_X1 U7396 ( .A1(n6180), .A2(n6179), .ZN(n6195) );
  INV_X1 U7397 ( .A(n6180), .ZN(n6181) );
  NAND2_X1 U7398 ( .A1(n6181), .A2(SI_26_), .ZN(n6182) );
  XNOR2_X1 U7399 ( .A(n6194), .B(n6193), .ZN(n8241) );
  NAND2_X1 U7400 ( .A1(n8241), .A2(n5981), .ZN(n6184) );
  NAND2_X1 U7401 ( .A1(n6072), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n6183) );
  NAND2_X1 U7402 ( .A1(n4930), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n6191) );
  INV_X1 U7403 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n6185) );
  OR2_X1 U7404 ( .A1(n8426), .A2(n6185), .ZN(n6190) );
  OR2_X2 U7405 ( .A1(n6186), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6206) );
  NAND2_X1 U7406 ( .A1(n6186), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6187) );
  INV_X1 U7407 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n9066) );
  OR2_X1 U7408 ( .A1(n5857), .A2(n9066), .ZN(n6188) );
  XNOR2_X1 U7409 ( .A(n9260), .B(n9077), .ZN(n9062) );
  INV_X1 U7410 ( .A(n9062), .ZN(n9069) );
  NAND2_X1 U7411 ( .A1(n9070), .A2(n9069), .ZN(n9071) );
  NOR2_X1 U7412 ( .A1(n9260), .A2(n9077), .ZN(n8383) );
  INV_X1 U7413 ( .A(n8383), .ZN(n6192) );
  NAND2_X1 U7414 ( .A1(n6194), .A2(n6193), .ZN(n6196) );
  INV_X1 U7415 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n6198) );
  INV_X1 U7416 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n6197) );
  MUX2_X1 U7417 ( .A(n6198), .B(n6197), .S(n5046), .Z(n6200) );
  INV_X1 U7418 ( .A(SI_27_), .ZN(n6199) );
  NAND2_X1 U7419 ( .A1(n6200), .A2(n6199), .ZN(n6228) );
  INV_X1 U7420 ( .A(n6200), .ZN(n6201) );
  NAND2_X1 U7421 ( .A1(n6201), .A2(SI_27_), .ZN(n6202) );
  NAND2_X1 U7422 ( .A1(n8246), .A2(n5981), .ZN(n6204) );
  NAND2_X1 U7423 ( .A1(n6072), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n6203) );
  NAND2_X1 U7424 ( .A1(n4930), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n6212) );
  INV_X1 U7425 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n9307) );
  OR2_X1 U7426 ( .A1(n8426), .A2(n9307), .ZN(n6211) );
  INV_X1 U7427 ( .A(n6206), .ZN(n6205) );
  INV_X1 U7428 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n8807) );
  NAND2_X1 U7429 ( .A1(n6205), .A2(n8807), .ZN(n6219) );
  NAND2_X1 U7430 ( .A1(n6206), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6207) );
  AND2_X1 U7431 ( .A1(n6219), .A2(n6207), .ZN(n9054) );
  OR2_X1 U7432 ( .A1(n4929), .A2(n9054), .ZN(n6210) );
  INV_X1 U7433 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n9055) );
  OR2_X1 U7434 ( .A1(n5857), .A2(n9055), .ZN(n6209) );
  AND4_X2 U7435 ( .A1(n6212), .A2(n6211), .A3(n6210), .A4(n6209), .ZN(n9064)
         );
  INV_X1 U7436 ( .A(n8388), .ZN(n6213) );
  NAND2_X1 U7437 ( .A1(n9057), .A2(n9064), .ZN(n8389) );
  NAND2_X1 U7438 ( .A1(n6233), .A2(n6228), .ZN(n6216) );
  MUX2_X1 U7439 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n7103), .Z(n6225) );
  INV_X1 U7440 ( .A(SI_28_), .ZN(n6226) );
  XNOR2_X1 U7441 ( .A(n6225), .B(n6226), .ZN(n6230) );
  NAND2_X1 U7442 ( .A1(n9343), .A2(n5981), .ZN(n6218) );
  NAND2_X1 U7443 ( .A1(n6072), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n6217) );
  NAND2_X1 U7444 ( .A1(n4930), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6224) );
  INV_X1 U7445 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n6879) );
  OR2_X1 U7446 ( .A1(n8426), .A2(n6879), .ZN(n6223) );
  NAND2_X1 U7447 ( .A1(n6219), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n6220) );
  INV_X1 U7448 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n9042) );
  OR2_X1 U7449 ( .A1(n5857), .A2(n9042), .ZN(n6221) );
  NAND4_X1 U7450 ( .A1(n6224), .A2(n6223), .A3(n6222), .A4(n6221), .ZN(n8928)
         );
  XNOR2_X1 U7451 ( .A(n9045), .B(n9053), .ZN(n6874) );
  INV_X1 U7452 ( .A(n6225), .ZN(n6227) );
  NAND2_X1 U7453 ( .A1(n6227), .A2(n6226), .ZN(n6229) );
  AND2_X1 U7454 ( .A1(n6228), .A2(n6229), .ZN(n6232) );
  INV_X1 U7455 ( .A(n6229), .ZN(n6231) );
  INV_X1 U7456 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n6235) );
  INV_X1 U7457 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n6234) );
  MUX2_X1 U7458 ( .A(n6235), .B(n6234), .S(n8416), .Z(n8400) );
  NAND2_X1 U7459 ( .A1(n6802), .A2(n5981), .ZN(n6237) );
  NAND2_X1 U7460 ( .A1(n6072), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n6236) );
  NAND2_X1 U7461 ( .A1(n6237), .A2(n6236), .ZN(n6855) );
  OR2_X1 U7462 ( .A1(n4929), .A2(n6319), .ZN(n8431) );
  INV_X1 U7463 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n6867) );
  OR2_X1 U7464 ( .A1(n8426), .A2(n6867), .ZN(n6240) );
  INV_X1 U7465 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n6320) );
  OR2_X1 U7466 ( .A1(n5857), .A2(n6320), .ZN(n6239) );
  INV_X1 U7467 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n6856) );
  OR2_X1 U7468 ( .A1(n8424), .A2(n6856), .ZN(n6238) );
  OR2_X1 U7469 ( .A1(n6855), .A2(n9040), .ZN(n8395) );
  NAND2_X1 U7470 ( .A1(n6855), .A2(n9040), .ZN(n8435) );
  XNOR2_X2 U7471 ( .A(n6242), .B(n6241), .ZN(n7409) );
  NAND2_X1 U7472 ( .A1(n7409), .A2(n7833), .ZN(n6297) );
  NAND2_X1 U7473 ( .A1(n7433), .A2(n10740), .ZN(n7619) );
  NOR2_X1 U7474 ( .A1(n7409), .A2(n8484), .ZN(n6243) );
  INV_X1 U7475 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n6245) );
  AOI22_X1 U7476 ( .A1(n4930), .A2(P2_REG1_REG_30__SCAN_IN), .B1(n4932), .B2(
        P2_REG0_REG_30__SCAN_IN), .ZN(n6244) );
  OAI211_X1 U7477 ( .C1(n5857), .C2(n6245), .A(n8431), .B(n6244), .ZN(n8927)
         );
  OAI21_X1 U7478 ( .B1(n5648), .B2(n8480), .A(n5765), .ZN(n6247) );
  NAND2_X1 U7479 ( .A1(n5765), .A2(P2_B_REG_SCAN_IN), .ZN(n6246) );
  AND2_X1 U7480 ( .A1(n10658), .A2(n6246), .ZN(n9031) );
  INV_X1 U7481 ( .A(n6247), .ZN(n7435) );
  AOI22_X1 U7482 ( .A1(n8927), .A2(n9031), .B1(n9216), .B2(n8928), .ZN(n6292)
         );
  INV_X1 U7483 ( .A(n7499), .ZN(n7626) );
  NAND2_X1 U7484 ( .A1(n6249), .A2(n7626), .ZN(n7387) );
  NAND2_X1 U7485 ( .A1(n7628), .A2(n7414), .ZN(n6250) );
  OR2_X1 U7486 ( .A1(n8941), .A2(n7481), .ZN(n6251) );
  INV_X1 U7487 ( .A(n10577), .ZN(n6252) );
  NOR2_X1 U7488 ( .A1(n8940), .A2(n6252), .ZN(n6253) );
  OAI22_X1 U7489 ( .A1(n7786), .A2(n6253), .B1(n7438), .B2(n10577), .ZN(n7776)
         );
  NAND2_X1 U7490 ( .A1(n7776), .A2(n8447), .ZN(n8000) );
  INV_X1 U7491 ( .A(n7413), .ZN(n10585) );
  NAND2_X1 U7492 ( .A1(n8939), .A2(n10585), .ZN(n7999) );
  INV_X1 U7493 ( .A(n10600), .ZN(n8007) );
  NAND2_X1 U7494 ( .A1(n8007), .A2(n8938), .ZN(n6254) );
  AND2_X1 U7495 ( .A1(n7999), .A2(n6254), .ZN(n6255) );
  NAND2_X1 U7496 ( .A1(n8000), .A2(n6255), .ZN(n6257) );
  OR2_X1 U7497 ( .A1(n8938), .A2(n8007), .ZN(n6256) );
  AND2_X1 U7498 ( .A1(n8301), .A2(n8278), .ZN(n8451) );
  INV_X1 U7499 ( .A(n8451), .ZN(n7884) );
  AND2_X1 U7500 ( .A1(n7884), .A2(n8453), .ZN(n6258) );
  NAND2_X1 U7501 ( .A1(n7665), .A2(n6258), .ZN(n6260) );
  INV_X1 U7502 ( .A(n8937), .ZN(n10601) );
  NAND2_X1 U7503 ( .A1(n10601), .A2(n7715), .ZN(n7885) );
  INV_X1 U7504 ( .A(n10619), .ZN(n7758) );
  NAND2_X1 U7505 ( .A1(n6260), .A2(n6259), .ZN(n7812) );
  NAND2_X1 U7506 ( .A1(n8283), .A2(n8287), .ZN(n8452) );
  NAND2_X1 U7507 ( .A1(n7812), .A2(n8452), .ZN(n6262) );
  OR2_X1 U7508 ( .A1(n10642), .A2(n10620), .ZN(n6261) );
  NAND2_X1 U7509 ( .A1(n6262), .A2(n6261), .ZN(n8030) );
  NAND2_X1 U7510 ( .A1(n8030), .A2(n8454), .ZN(n6264) );
  INV_X1 U7511 ( .A(n8042), .ZN(n8015) );
  OR2_X1 U7512 ( .A1(n5895), .A2(n8015), .ZN(n6263) );
  NAND2_X1 U7513 ( .A1(n6264), .A2(n6263), .ZN(n8041) );
  INV_X1 U7514 ( .A(n8457), .ZN(n6265) );
  NAND2_X1 U7515 ( .A1(n8041), .A2(n6265), .ZN(n6267) );
  OR2_X1 U7516 ( .A1(n10685), .A2(n10657), .ZN(n6266) );
  NAND2_X1 U7517 ( .A1(n6267), .A2(n6266), .ZN(n8021) );
  NOR2_X1 U7518 ( .A1(n10695), .A2(n8073), .ZN(n6269) );
  NAND2_X1 U7519 ( .A1(n10695), .A2(n8073), .ZN(n6268) );
  NAND2_X1 U7520 ( .A1(n10708), .A2(n8935), .ZN(n7983) );
  INV_X1 U7521 ( .A(n7983), .ZN(n6270) );
  OR2_X1 U7522 ( .A1(n10708), .A2(n8935), .ZN(n8150) );
  NAND2_X1 U7523 ( .A1(n9231), .A2(n6272), .ZN(n6273) );
  NAND2_X1 U7524 ( .A1(n6273), .A2(n8326), .ZN(n9214) );
  NAND2_X1 U7525 ( .A1(n8330), .A2(n8329), .ZN(n9213) );
  INV_X1 U7526 ( .A(n9237), .ZN(n8933) );
  NAND2_X1 U7527 ( .A1(n10725), .A2(n8933), .ZN(n6274) );
  XNOR2_X1 U7528 ( .A(n8848), .B(n8917), .ZN(n9203) );
  XNOR2_X1 U7529 ( .A(n8862), .B(n9201), .ZN(n9190) );
  NAND2_X1 U7530 ( .A1(n9185), .A2(n9190), .ZN(n6276) );
  OR2_X1 U7531 ( .A1(n10741), .A2(n9201), .ZN(n6275) );
  AND2_X1 U7532 ( .A1(n10752), .A2(n9194), .ZN(n6277) );
  OR2_X1 U7533 ( .A1(n10752), .A2(n9194), .ZN(n6278) );
  NOR2_X1 U7534 ( .A1(n9296), .A2(n8931), .ZN(n9140) );
  INV_X1 U7535 ( .A(n6279), .ZN(n6280) );
  INV_X1 U7536 ( .A(n9134), .ZN(n9129) );
  NAND2_X1 U7537 ( .A1(n9296), .A2(n8931), .ZN(n9142) );
  AND2_X1 U7538 ( .A1(n9154), .A2(n9142), .ZN(n9141) );
  OR2_X1 U7539 ( .A1(n6280), .A2(n9141), .ZN(n9125) );
  AND2_X1 U7540 ( .A1(n9129), .A2(n9125), .ZN(n6281) );
  INV_X1 U7541 ( .A(n9273), .ZN(n9106) );
  OAI21_X1 U7542 ( .B1(n9093), .B2(n9102), .A(n9087), .ZN(n9074) );
  INV_X1 U7543 ( .A(n9078), .ZN(n9314) );
  NAND2_X1 U7544 ( .A1(n9074), .A2(n5515), .ZN(n6285) );
  NAND2_X1 U7545 ( .A1(n6285), .A2(n6284), .ZN(n9061) );
  INV_X1 U7546 ( .A(n9260), .ZN(n8382) );
  INV_X1 U7547 ( .A(n9077), .ZN(n8929) );
  INV_X1 U7548 ( .A(n9057), .ZN(n9309) );
  INV_X1 U7549 ( .A(n9064), .ZN(n9259) );
  OR2_X1 U7550 ( .A1(n9045), .A2(n8928), .ZN(n8393) );
  INV_X1 U7551 ( .A(n8393), .ZN(n6287) );
  NAND2_X1 U7552 ( .A1(n9045), .A2(n8928), .ZN(n8391) );
  OAI21_X1 U7553 ( .B1(n6875), .B2(n6287), .A(n8391), .ZN(n6288) );
  XNOR2_X1 U7554 ( .A(n6288), .B(n4966), .ZN(n6290) );
  OR2_X1 U7555 ( .A1(n8254), .A2(n7409), .ZN(n6289) );
  NAND2_X1 U7556 ( .A1(n8479), .A2(n8484), .ZN(n6862) );
  NAND2_X1 U7557 ( .A1(n6290), .A2(n9211), .ZN(n6291) );
  INV_X1 U7558 ( .A(n6294), .ZN(n6846) );
  NOR2_X1 U7559 ( .A1(n8254), .A2(n7765), .ZN(n7693) );
  OR2_X1 U7560 ( .A1(n8479), .A2(n7948), .ZN(n6295) );
  NOR2_X1 U7561 ( .A1(n7409), .A2(n6295), .ZN(n6296) );
  NAND2_X1 U7562 ( .A1(n8396), .A2(n6297), .ZN(n7445) );
  NAND2_X1 U7563 ( .A1(n6850), .A2(n7445), .ZN(n6852) );
  XNOR2_X1 U7564 ( .A(n6298), .B(P2_B_REG_SCAN_IN), .ZN(n6299) );
  NAND2_X1 U7565 ( .A1(n6299), .A2(n8240), .ZN(n6300) );
  NAND2_X1 U7566 ( .A1(n8240), .A2(n6303), .ZN(n6301) );
  NAND2_X1 U7567 ( .A1(n6298), .A2(n6303), .ZN(n7226) );
  AOI22_X1 U7568 ( .A1(n6852), .A2(n7135), .B1(n7406), .B2(n6850), .ZN(n6317)
         );
  NOR2_X1 U7569 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .ZN(
        n6308) );
  NOR4_X1 U7570 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n6307) );
  NOR4_X1 U7571 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n6306) );
  NOR4_X1 U7572 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n6305) );
  NAND4_X1 U7573 ( .A1(n6308), .A2(n6307), .A3(n6306), .A4(n6305), .ZN(n6314)
         );
  NOR4_X1 U7574 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n6312) );
  NOR4_X1 U7575 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n6311) );
  NOR4_X1 U7576 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6310) );
  NOR4_X1 U7577 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n6309) );
  NAND4_X1 U7578 ( .A1(n6312), .A2(n6311), .A3(n6310), .A4(n6309), .ZN(n6313)
         );
  NOR2_X1 U7579 ( .A1(n6314), .A2(n6313), .ZN(n6315) );
  AND2_X1 U7580 ( .A1(n6864), .A2(n7428), .ZN(n6316) );
  INV_X1 U7581 ( .A(n7765), .ZN(n6318) );
  NOR2_X2 U7582 ( .A1(n7620), .A2(n9240), .ZN(n10641) );
  NOR2_X1 U7583 ( .A1(n9238), .A2(n6319), .ZN(n9034) );
  NOR2_X1 U7584 ( .A1(n10643), .A2(n6320), .ZN(n6321) );
  AOI211_X1 U7585 ( .C1(n6855), .C2(n10641), .A(n9034), .B(n6321), .ZN(n6322)
         );
  NAND2_X1 U7586 ( .A1(n6323), .A2(n6322), .ZN(P2_U3204) );
  NOR2_X1 U7587 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n6328) );
  NOR2_X1 U7588 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), .ZN(
        n6327) );
  NAND2_X1 U7589 ( .A1(n6773), .A2(n6329), .ZN(n6330) );
  NOR2_X2 U7590 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(n6330), .ZN(n6351) );
  NAND2_X1 U7591 ( .A1(n6331), .A2(n6351), .ZN(n6332) );
  NAND2_X1 U7592 ( .A1(n8491), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6347) );
  AND2_X2 U7593 ( .A1(n10006), .A2(n6341), .ZN(n6400) );
  NAND2_X1 U7594 ( .A1(n6400), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6346) );
  AND2_X2 U7595 ( .A1(n6342), .A2(n6341), .ZN(n6441) );
  NAND2_X1 U7596 ( .A1(n6441), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n6345) );
  INV_X1 U7597 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n6343) );
  INV_X1 U7598 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n9526) );
  INV_X1 U7599 ( .A(SI_0_), .ZN(n10162) );
  INV_X1 U7600 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n6348) );
  OAI21_X1 U7601 ( .B1(n8416), .B2(n10162), .A(n6348), .ZN(n6350) );
  NAND2_X1 U7602 ( .A1(n6350), .A2(n6349), .ZN(n10016) );
  NOR2_X1 U7603 ( .A1(n6787), .A2(P1_IR_REG_23__SCAN_IN), .ZN(n6352) );
  NAND2_X1 U7604 ( .A1(n6352), .A2(n6351), .ZN(n6354) );
  NAND2_X2 U7605 ( .A1(n6358), .A2(n6357), .ZN(n9525) );
  INV_X1 U7606 ( .A(n6359), .ZN(n6363) );
  NAND2_X1 U7607 ( .A1(n6360), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6361) );
  MUX2_X1 U7608 ( .A(n9526), .B(n10016), .S(n7122), .Z(n10518) );
  OR2_X1 U7609 ( .A1(n6895), .A2(n10518), .ZN(n7365) );
  INV_X1 U7610 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n6364) );
  NAND2_X1 U7611 ( .A1(n6400), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6365) );
  AND2_X1 U7612 ( .A1(n6366), .A2(n6365), .ZN(n6369) );
  NAND2_X1 U7613 ( .A1(n6441), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n6368) );
  NAND2_X1 U7614 ( .A1(n8491), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6367) );
  NAND3_X2 U7615 ( .A1(n6369), .A2(n6368), .A3(n6367), .ZN(n6902) );
  NAND2_X1 U7616 ( .A1(n6405), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n6372) );
  NAND2_X1 U7617 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n6370) );
  XNOR2_X1 U7618 ( .A(n6370), .B(P1_IR_REG_1__SCAN_IN), .ZN(n9515) );
  OAI211_X2 U7619 ( .C1(n6419), .C2(n7106), .A(n6372), .B(n6371), .ZN(n7366)
         );
  NAND2_X1 U7620 ( .A1(n7215), .A2(n7366), .ZN(n6742) );
  NAND2_X1 U7621 ( .A1(n6902), .A2(n6373), .ZN(n8684) );
  NAND2_X1 U7622 ( .A1(n7365), .A2(n6741), .ZN(n6375) );
  NAND2_X1 U7623 ( .A1(n7215), .A2(n6373), .ZN(n6374) );
  NAND2_X1 U7624 ( .A1(n8491), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6380) );
  INV_X1 U7625 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n6376) );
  NAND2_X1 U7626 ( .A1(n6400), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6378) );
  NAND2_X1 U7627 ( .A1(n6441), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n6377) );
  NAND2_X1 U7628 ( .A1(n6405), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n6383) );
  OR2_X1 U7629 ( .A1(n6381), .A2(n6509), .ZN(n6392) );
  XNOR2_X1 U7630 ( .A(n6392), .B(P1_IR_REG_2__SCAN_IN), .ZN(n9535) );
  NAND2_X1 U7631 ( .A1(n6616), .A2(n9535), .ZN(n6382) );
  NAND2_X1 U7632 ( .A1(n9512), .A2(n10538), .ZN(n8683) );
  NAND2_X1 U7633 ( .A1(n7513), .A2(n10553), .ZN(n6743) );
  NAND2_X1 U7634 ( .A1(n7513), .A2(n10538), .ZN(n6384) );
  NAND2_X1 U7635 ( .A1(n6385), .A2(n6384), .ZN(n7511) );
  NAND2_X1 U7636 ( .A1(n8491), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6390) );
  NAND2_X1 U7637 ( .A1(n6400), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6388) );
  NAND2_X1 U7638 ( .A1(n6441), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n6387) );
  INV_X1 U7639 ( .A(n10544), .ZN(n6397) );
  NAND2_X1 U7640 ( .A1(n6405), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n6396) );
  INV_X1 U7641 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n6391) );
  NAND2_X1 U7642 ( .A1(n6392), .A2(n6391), .ZN(n6393) );
  NAND2_X1 U7643 ( .A1(n6393), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6394) );
  XNOR2_X1 U7644 ( .A(n6394), .B(P1_IR_REG_3__SCAN_IN), .ZN(n9548) );
  NAND2_X1 U7645 ( .A1(n6616), .A2(n9548), .ZN(n6395) );
  NAND2_X1 U7646 ( .A1(n6397), .A2(n7523), .ZN(n8495) );
  NAND2_X1 U7647 ( .A1(n8495), .A2(n8498), .ZN(n6745) );
  NAND2_X1 U7648 ( .A1(n8491), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6404) );
  INV_X1 U7649 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n6399) );
  XNOR2_X1 U7650 ( .A(n6399), .B(P1_REG3_REG_3__SCAN_IN), .ZN(n7546) );
  NAND2_X1 U7651 ( .A1(n6579), .A2(n7546), .ZN(n6403) );
  NAND2_X1 U7652 ( .A1(n6400), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6402) );
  NAND2_X1 U7653 ( .A1(n6441), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n6401) );
  NAND2_X1 U7654 ( .A1(n6405), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n6409) );
  NAND2_X1 U7655 ( .A1(n6406), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6407) );
  XNOR2_X1 U7656 ( .A(n6407), .B(P1_IR_REG_4__SCAN_IN), .ZN(n9558) );
  NAND2_X1 U7657 ( .A1(n6616), .A2(n9558), .ZN(n6408) );
  OAI211_X1 U7658 ( .C1(n6419), .C2(n7111), .A(n6409), .B(n6408), .ZN(n7547)
         );
  NOR2_X1 U7659 ( .A1(n9511), .A2(n7547), .ZN(n6410) );
  NAND2_X1 U7660 ( .A1(n8491), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6418) );
  NAND2_X1 U7661 ( .A1(n6411), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n6430) );
  INV_X1 U7662 ( .A(n6411), .ZN(n6413) );
  INV_X1 U7663 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n6412) );
  NAND2_X1 U7664 ( .A1(n6413), .A2(n6412), .ZN(n6414) );
  AND2_X1 U7665 ( .A1(n6430), .A2(n6414), .ZN(n7397) );
  NAND2_X1 U7666 ( .A1(n6579), .A2(n7397), .ZN(n6417) );
  NAND2_X1 U7667 ( .A1(n6400), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6416) );
  NAND2_X1 U7668 ( .A1(n6441), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n6415) );
  NAND4_X1 U7669 ( .A1(n6418), .A2(n6417), .A3(n6416), .A4(n6415), .ZN(n9510)
         );
  INV_X1 U7670 ( .A(n9510), .ZN(n7575) );
  INV_X2 U7671 ( .A(n6419), .ZN(n6490) );
  NAND2_X1 U7672 ( .A1(n7114), .A2(n6490), .ZN(n6423) );
  NAND2_X1 U7673 ( .A1(n6420), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6421) );
  XNOR2_X1 U7674 ( .A(n6421), .B(P1_IR_REG_5__SCAN_IN), .ZN(n9575) );
  AOI22_X1 U7675 ( .A1(n6405), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n6616), .B2(
        n9575), .ZN(n6422) );
  NAND2_X1 U7676 ( .A1(n6423), .A2(n6422), .ZN(n7491) );
  NAND2_X1 U7677 ( .A1(n7575), .A2(n7491), .ZN(n8501) );
  INV_X1 U7678 ( .A(n7491), .ZN(n7494) );
  NAND2_X1 U7679 ( .A1(n7119), .A2(n6490), .ZN(n6427) );
  OR2_X1 U7680 ( .A1(n6424), .A2(n6509), .ZN(n6425) );
  XNOR2_X1 U7681 ( .A(n6425), .B(P1_IR_REG_6__SCAN_IN), .ZN(n9588) );
  AOI22_X1 U7682 ( .A1(n6405), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n6616), .B2(
        n9588), .ZN(n6426) );
  NAND2_X1 U7683 ( .A1(n6427), .A2(n6426), .ZN(n10609) );
  INV_X1 U7684 ( .A(n10609), .ZN(n7584) );
  NAND2_X1 U7685 ( .A1(n8491), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6435) );
  INV_X1 U7686 ( .A(n6430), .ZN(n6428) );
  NAND2_X1 U7687 ( .A1(n6428), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n6439) );
  INV_X1 U7688 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6429) );
  NAND2_X1 U7689 ( .A1(n6430), .A2(n6429), .ZN(n6431) );
  AND2_X1 U7690 ( .A1(n6439), .A2(n6431), .ZN(n7582) );
  NAND2_X1 U7691 ( .A1(n6579), .A2(n7582), .ZN(n6434) );
  NAND2_X1 U7692 ( .A1(n6400), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6433) );
  NAND2_X1 U7693 ( .A1(n6441), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n6432) );
  NAND4_X1 U7694 ( .A1(n6435), .A2(n6434), .A3(n6433), .A4(n6432), .ZN(n9509)
         );
  NAND2_X1 U7695 ( .A1(n7584), .A2(n9509), .ZN(n8505) );
  INV_X1 U7696 ( .A(n9509), .ZN(n7677) );
  NAND2_X1 U7697 ( .A1(n7677), .A2(n10609), .ZN(n8506) );
  NAND2_X1 U7698 ( .A1(n8505), .A2(n8506), .ZN(n8612) );
  NAND2_X1 U7699 ( .A1(n7584), .A2(n7677), .ZN(n6436) );
  NAND2_X1 U7700 ( .A1(n7573), .A2(n6436), .ZN(n7680) );
  NAND2_X1 U7701 ( .A1(n8491), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6445) );
  INV_X1 U7702 ( .A(n6439), .ZN(n6437) );
  NAND2_X1 U7703 ( .A1(n6437), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n6455) );
  INV_X1 U7704 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n6438) );
  NAND2_X1 U7705 ( .A1(n6439), .A2(n6438), .ZN(n6440) );
  AND2_X1 U7706 ( .A1(n6455), .A2(n6440), .ZN(n7685) );
  NAND2_X1 U7707 ( .A1(n6579), .A2(n7685), .ZN(n6444) );
  NAND2_X1 U7708 ( .A1(n6400), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6443) );
  NAND2_X1 U7709 ( .A1(n6441), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n6442) );
  NAND4_X1 U7710 ( .A1(n6445), .A2(n6444), .A3(n6443), .A4(n6442), .ZN(n9508)
         );
  NAND2_X1 U7711 ( .A1(n7139), .A2(n6490), .ZN(n6449) );
  NAND2_X1 U7712 ( .A1(n6424), .A2(n6446), .ZN(n6451) );
  NAND2_X1 U7713 ( .A1(n6451), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6447) );
  XNOR2_X1 U7714 ( .A(n6447), .B(P1_IR_REG_7__SCAN_IN), .ZN(n10291) );
  AOI22_X1 U7715 ( .A1(n6405), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n6616), .B2(
        n10291), .ZN(n6448) );
  NAND2_X1 U7716 ( .A1(n6449), .A2(n6448), .ZN(n7684) );
  OR2_X1 U7717 ( .A1(n7826), .A2(n7684), .ZN(n8508) );
  NAND2_X1 U7718 ( .A1(n7684), .A2(n7826), .ZN(n8516) );
  NAND2_X1 U7719 ( .A1(n8508), .A2(n8516), .ZN(n8613) );
  OR2_X1 U7720 ( .A1(n7684), .A2(n9508), .ZN(n6450) );
  NAND2_X1 U7721 ( .A1(n6462), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6452) );
  XNOR2_X1 U7722 ( .A(n6452), .B(P1_IR_REG_8__SCAN_IN), .ZN(n10295) );
  AOI22_X1 U7723 ( .A1(n6405), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n6616), .B2(
        n10295), .ZN(n6453) );
  NAND2_X1 U7724 ( .A1(n6455), .A2(n6454), .ZN(n6456) );
  AND2_X1 U7725 ( .A1(n6467), .A2(n6456), .ZN(n7822) );
  NAND2_X1 U7726 ( .A1(n6579), .A2(n7822), .ZN(n6460) );
  NAND2_X1 U7727 ( .A1(n8491), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6459) );
  NAND2_X1 U7728 ( .A1(n6400), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6458) );
  NAND2_X1 U7729 ( .A1(n6441), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n6457) );
  NAND4_X1 U7730 ( .A1(n6460), .A2(n6459), .A3(n6458), .A4(n6457), .ZN(n9507)
         );
  INV_X1 U7731 ( .A(n9507), .ZN(n7678) );
  NAND2_X1 U7732 ( .A1(n7645), .A2(n8510), .ZN(n8614) );
  NAND2_X1 U7733 ( .A1(n6461), .A2(n6490), .ZN(n6464) );
  NAND2_X1 U7734 ( .A1(n6508), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6475) );
  XNOR2_X1 U7735 ( .A(n6475), .B(P1_IR_REG_9__SCAN_IN), .ZN(n7354) );
  AOI22_X1 U7736 ( .A1(n6405), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n6616), .B2(
        n7354), .ZN(n6463) );
  INV_X1 U7737 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n6466) );
  NAND2_X1 U7738 ( .A1(n6467), .A2(n6466), .ZN(n6468) );
  AND2_X1 U7739 ( .A1(n6483), .A2(n6468), .ZN(n7862) );
  NAND2_X1 U7740 ( .A1(n6579), .A2(n7862), .ZN(n6472) );
  NAND2_X1 U7741 ( .A1(n8491), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6471) );
  NAND2_X1 U7742 ( .A1(n6400), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6470) );
  NAND2_X1 U7743 ( .A1(n6441), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n6469) );
  NAND4_X1 U7744 ( .A1(n6472), .A2(n6471), .A3(n6470), .A4(n6469), .ZN(n9506)
         );
  INV_X1 U7745 ( .A(n9506), .ZN(n7959) );
  NAND2_X1 U7746 ( .A1(n7657), .A2(n7959), .ZN(n8526) );
  NAND2_X1 U7747 ( .A1(n8525), .A2(n8526), .ZN(n8617) );
  NAND2_X1 U7748 ( .A1(n7651), .A2(n8617), .ZN(n7653) );
  OR2_X1 U7749 ( .A1(n7657), .A2(n9506), .ZN(n6473) );
  NAND2_X1 U7750 ( .A1(n7653), .A2(n6473), .ZN(n7598) );
  NAND2_X1 U7751 ( .A1(n7203), .A2(n6490), .ZN(n6481) );
  INV_X1 U7752 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n6474) );
  INV_X1 U7753 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n6509) );
  AOI21_X1 U7754 ( .B1(n6475), .B2(n6474), .A(n6509), .ZN(n6476) );
  NAND2_X1 U7755 ( .A1(n6476), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n6479) );
  INV_X1 U7756 ( .A(n6476), .ZN(n6478) );
  INV_X1 U7757 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n6477) );
  NAND2_X1 U7758 ( .A1(n6478), .A2(n6477), .ZN(n6491) );
  AOI22_X1 U7759 ( .A1(n6405), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6616), .B2(
        n10389), .ZN(n6480) );
  NAND2_X1 U7760 ( .A1(n8491), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6488) );
  NAND2_X1 U7761 ( .A1(n6483), .A2(n6482), .ZN(n6484) );
  AND2_X1 U7762 ( .A1(n6496), .A2(n6484), .ZN(n7955) );
  NAND2_X1 U7763 ( .A1(n6579), .A2(n7955), .ZN(n6487) );
  NAND2_X1 U7764 ( .A1(n6400), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6486) );
  NAND2_X1 U7765 ( .A1(n6441), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n6485) );
  NAND4_X1 U7766 ( .A1(n6488), .A2(n6487), .A3(n6486), .A4(n6485), .ZN(n9505)
         );
  OR2_X1 U7767 ( .A1(n7961), .A2(n7860), .ZN(n8534) );
  NAND2_X1 U7768 ( .A1(n7961), .A2(n7860), .ZN(n8529) );
  NAND2_X1 U7769 ( .A1(n8534), .A2(n8529), .ZN(n8618) );
  NAND2_X1 U7770 ( .A1(n7598), .A2(n8618), .ZN(n7597) );
  OR2_X1 U7771 ( .A1(n7961), .A2(n9505), .ZN(n6489) );
  NAND2_X1 U7772 ( .A1(n7597), .A2(n6489), .ZN(n7738) );
  NAND2_X1 U7773 ( .A1(n6491), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6492) );
  XNOR2_X1 U7774 ( .A(n6492), .B(P1_IR_REG_11__SCAN_IN), .ZN(n10320) );
  AOI22_X1 U7775 ( .A1(n6405), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n6616), .B2(
        n10320), .ZN(n6493) );
  NAND2_X1 U7776 ( .A1(n8491), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n6501) );
  INV_X1 U7777 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n6495) );
  NAND2_X1 U7778 ( .A1(n6496), .A2(n6495), .ZN(n6497) );
  AND2_X1 U7779 ( .A1(n6517), .A2(n6497), .ZN(n9853) );
  NAND2_X1 U7780 ( .A1(n6579), .A2(n9853), .ZN(n6500) );
  NAND2_X1 U7781 ( .A1(n6400), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6499) );
  NAND2_X1 U7782 ( .A1(n6441), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n6498) );
  NAND4_X1 U7783 ( .A1(n6501), .A2(n6500), .A3(n6499), .A4(n6498), .ZN(n9504)
         );
  NAND2_X1 U7784 ( .A1(n9858), .A2(n9504), .ZN(n6502) );
  NAND2_X1 U7785 ( .A1(n7738), .A2(n6502), .ZN(n6504) );
  OR2_X1 U7786 ( .A1(n9858), .A2(n9504), .ZN(n6503) );
  NAND2_X1 U7787 ( .A1(n7263), .A2(n6490), .ZN(n6516) );
  INV_X1 U7788 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n6505) );
  NAND2_X1 U7789 ( .A1(n6506), .A2(n6505), .ZN(n6507) );
  NOR2_X1 U7790 ( .A1(n6513), .A2(n6509), .ZN(n6510) );
  MUX2_X1 U7791 ( .A(n6509), .B(n6510), .S(P1_IR_REG_12__SCAN_IN), .Z(n6511)
         );
  INV_X1 U7792 ( .A(n6511), .ZN(n6514) );
  INV_X1 U7793 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n6512) );
  NAND2_X1 U7794 ( .A1(n6513), .A2(n6512), .ZN(n6526) );
  AOI22_X1 U7795 ( .A1(n6405), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n6616), .B2(
        n8124), .ZN(n6515) );
  NAND2_X1 U7796 ( .A1(n8491), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n6522) );
  NAND2_X1 U7797 ( .A1(n6517), .A2(n7358), .ZN(n6518) );
  AND2_X1 U7798 ( .A1(n6531), .A2(n6518), .ZN(n8199) );
  NAND2_X1 U7799 ( .A1(n6579), .A2(n8199), .ZN(n6521) );
  NAND2_X1 U7800 ( .A1(n6400), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n6520) );
  NAND2_X1 U7801 ( .A1(n6441), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n6519) );
  NAND4_X1 U7802 ( .A1(n6522), .A2(n6521), .A3(n6520), .A4(n6519), .ZN(n9503)
         );
  NOR2_X1 U7803 ( .A1(n8542), .A2(n9503), .ZN(n6524) );
  NAND2_X1 U7804 ( .A1(n8542), .A2(n9503), .ZN(n6523) );
  NAND2_X1 U7805 ( .A1(n7267), .A2(n6490), .ZN(n6529) );
  NAND2_X1 U7806 ( .A1(n6526), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6525) );
  MUX2_X1 U7807 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6525), .S(
        P1_IR_REG_13__SCAN_IN), .Z(n6527) );
  AOI22_X1 U7808 ( .A1(n6405), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n6616), .B2(
        n10375), .ZN(n6528) );
  NAND2_X1 U7809 ( .A1(n8491), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n6536) );
  NAND2_X1 U7810 ( .A1(n6531), .A2(n6530), .ZN(n6532) );
  AND2_X1 U7811 ( .A1(n6545), .A2(n6532), .ZN(n9842) );
  NAND2_X1 U7812 ( .A1(n6579), .A2(n9842), .ZN(n6535) );
  NAND2_X1 U7813 ( .A1(n6400), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n6534) );
  NAND2_X1 U7814 ( .A1(n6441), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n6533) );
  NAND4_X1 U7815 ( .A1(n6536), .A2(n6535), .A3(n6534), .A4(n6533), .ZN(n9502)
         );
  NAND2_X1 U7816 ( .A1(n7316), .A2(n6490), .ZN(n6542) );
  NAND2_X1 U7817 ( .A1(n6537), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6570) );
  INV_X1 U7818 ( .A(n6570), .ZN(n6538) );
  NAND2_X1 U7819 ( .A1(n6538), .A2(P1_IR_REG_14__SCAN_IN), .ZN(n6540) );
  INV_X1 U7820 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n6539) );
  NAND2_X1 U7821 ( .A1(n6570), .A2(n6539), .ZN(n6553) );
  AOI22_X1 U7822 ( .A1(n6405), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n6616), .B2(
        n10324), .ZN(n6541) );
  INV_X1 U7823 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n6544) );
  NAND2_X1 U7824 ( .A1(n6545), .A2(n6544), .ZN(n6546) );
  AND2_X1 U7825 ( .A1(n6560), .A2(n6546), .ZN(n9353) );
  NAND2_X1 U7826 ( .A1(n6579), .A2(n9353), .ZN(n6550) );
  NAND2_X1 U7827 ( .A1(n8491), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n6549) );
  NAND2_X1 U7828 ( .A1(n6400), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n6548) );
  NAND2_X1 U7829 ( .A1(n6441), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n6547) );
  NAND4_X1 U7830 ( .A1(n6550), .A2(n6549), .A3(n6548), .A4(n6547), .ZN(n9501)
         );
  INV_X1 U7831 ( .A(n9501), .ZN(n9492) );
  OR2_X1 U7832 ( .A1(n9943), .A2(n9492), .ZN(n8708) );
  NAND2_X1 U7833 ( .A1(n9943), .A2(n9492), .ZN(n8711) );
  NAND2_X1 U7834 ( .A1(n9943), .A2(n9501), .ZN(n6552) );
  NAND2_X1 U7835 ( .A1(n7966), .A2(n6552), .ZN(n8085) );
  NAND2_X1 U7836 ( .A1(n7402), .A2(n6490), .ZN(n6557) );
  NAND2_X1 U7837 ( .A1(n6553), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6555) );
  INV_X1 U7838 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n6554) );
  XNOR2_X1 U7839 ( .A(n6555), .B(n6554), .ZN(n8128) );
  INV_X1 U7840 ( .A(n8128), .ZN(n10350) );
  AOI22_X1 U7841 ( .A1(n6616), .A2(n10350), .B1(n6405), .B2(
        P2_DATAO_REG_15__SCAN_IN), .ZN(n6556) );
  NAND2_X1 U7842 ( .A1(n8491), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n6565) );
  INV_X1 U7843 ( .A(n6560), .ZN(n6558) );
  INV_X1 U7844 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n6559) );
  NAND2_X1 U7845 ( .A1(n6560), .A2(n6559), .ZN(n6561) );
  AND2_X1 U7846 ( .A1(n6577), .A2(n6561), .ZN(n9485) );
  NAND2_X1 U7847 ( .A1(n6579), .A2(n9485), .ZN(n6564) );
  NAND2_X1 U7848 ( .A1(n6400), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n6563) );
  NAND2_X1 U7849 ( .A1(n6441), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n6562) );
  NAND4_X1 U7850 ( .A1(n6565), .A2(n6564), .A3(n6563), .A4(n6562), .ZN(n9820)
         );
  INV_X1 U7851 ( .A(n9820), .ZN(n9402) );
  OR2_X1 U7852 ( .A1(n9998), .A2(n9402), .ZN(n8554) );
  NAND2_X1 U7853 ( .A1(n9998), .A2(n9402), .ZN(n9813) );
  NAND2_X1 U7854 ( .A1(n8554), .A2(n9813), .ZN(n8625) );
  NAND2_X1 U7855 ( .A1(n8085), .A2(n8625), .ZN(n8087) );
  NAND2_X1 U7856 ( .A1(n9998), .A2(n9820), .ZN(n6566) );
  NAND2_X1 U7857 ( .A1(n7534), .A2(n6490), .ZN(n6576) );
  INV_X1 U7858 ( .A(n6567), .ZN(n6568) );
  NAND2_X1 U7859 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n6568), .ZN(n6569) );
  INV_X1 U7860 ( .A(n6573), .ZN(n6571) );
  NAND2_X1 U7861 ( .A1(n6571), .A2(P1_IR_REG_16__SCAN_IN), .ZN(n6574) );
  INV_X1 U7862 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n6572) );
  NAND2_X1 U7863 ( .A1(n6573), .A2(n6572), .ZN(n6586) );
  AOI22_X1 U7864 ( .A1(n6405), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n8214), .B2(
        n6616), .ZN(n6575) );
  NAND2_X1 U7865 ( .A1(n8491), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n6583) );
  NAND2_X1 U7866 ( .A1(n6577), .A2(n8120), .ZN(n6578) );
  AND2_X1 U7867 ( .A1(n6592), .A2(n6578), .ZN(n9826) );
  NAND2_X1 U7868 ( .A1(n6579), .A2(n9826), .ZN(n6582) );
  NAND2_X1 U7869 ( .A1(n6400), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n6581) );
  NAND2_X1 U7870 ( .A1(n6441), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n6580) );
  NAND4_X1 U7871 ( .A1(n6583), .A2(n6582), .A3(n6581), .A4(n6580), .ZN(n9500)
         );
  INV_X1 U7872 ( .A(n9500), .ZN(n6584) );
  NAND2_X1 U7873 ( .A1(n9830), .A2(n6584), .ZN(n8714) );
  NAND2_X1 U7874 ( .A1(n8716), .A2(n8714), .ZN(n9834) );
  NAND2_X1 U7875 ( .A1(n9830), .A2(n9500), .ZN(n6585) );
  NAND2_X1 U7876 ( .A1(n7629), .A2(n6490), .ZN(n6589) );
  NAND2_X1 U7877 ( .A1(n6586), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6587) );
  XNOR2_X1 U7878 ( .A(n6587), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9604) );
  AOI22_X1 U7879 ( .A1(n9604), .A2(n6616), .B1(n6405), .B2(
        P2_DATAO_REG_17__SCAN_IN), .ZN(n6588) );
  NAND2_X1 U7880 ( .A1(n8491), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n6597) );
  INV_X1 U7881 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n6591) );
  NAND2_X1 U7882 ( .A1(n6592), .A2(n6591), .ZN(n6593) );
  AND2_X1 U7883 ( .A1(n6609), .A2(n6593), .ZN(n9414) );
  NAND2_X1 U7884 ( .A1(n6579), .A2(n9414), .ZN(n6596) );
  NAND2_X1 U7885 ( .A1(n6400), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n6595) );
  NAND2_X1 U7886 ( .A1(n6441), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n6594) );
  NAND4_X1 U7887 ( .A1(n6597), .A2(n6596), .A3(n6595), .A4(n6594), .ZN(n9819)
         );
  INV_X1 U7888 ( .A(n9819), .ZN(n9463) );
  NAND2_X1 U7889 ( .A1(n9925), .A2(n9463), .ZN(n8564) );
  NAND2_X1 U7890 ( .A1(n8718), .A2(n8564), .ZN(n8626) );
  NAND2_X1 U7891 ( .A1(n9925), .A2(n9819), .ZN(n6598) );
  NAND2_X1 U7892 ( .A1(n8183), .A2(n6598), .ZN(n9793) );
  NAND2_X1 U7893 ( .A1(n7703), .A2(n6490), .ZN(n6607) );
  INV_X1 U7894 ( .A(n6599), .ZN(n6602) );
  NAND2_X1 U7895 ( .A1(n5013), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6600) );
  MUX2_X1 U7896 ( .A(n6600), .B(P1_IR_REG_31__SCAN_IN), .S(n6603), .Z(n6601)
         );
  INV_X1 U7897 ( .A(n6601), .ZN(n6605) );
  NAND2_X1 U7898 ( .A1(n6728), .A2(n6729), .ZN(n6614) );
  INV_X1 U7899 ( .A(n6614), .ZN(n6604) );
  NOR2_X1 U7900 ( .A1(n6605), .A2(n6604), .ZN(n10363) );
  AOI22_X1 U7901 ( .A1(n6405), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n6616), .B2(
        n10363), .ZN(n6606) );
  INV_X1 U7902 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n6608) );
  NAND2_X1 U7903 ( .A1(n6609), .A2(n6608), .ZN(n6610) );
  AND2_X1 U7904 ( .A1(n6621), .A2(n6610), .ZN(n9799) );
  AOI22_X1 U7905 ( .A1(n9799), .A2(n6579), .B1(n6441), .B2(
        P1_REG0_REG_18__SCAN_IN), .ZN(n6612) );
  AOI22_X1 U7906 ( .A1(n8491), .A2(P1_REG1_REG_18__SCAN_IN), .B1(n6400), .B2(
        P1_REG2_REG_18__SCAN_IN), .ZN(n6611) );
  OR2_X1 U7907 ( .A1(n9989), .A2(n9776), .ZN(n8565) );
  NAND2_X1 U7908 ( .A1(n9989), .A2(n9776), .ZN(n9771) );
  NAND2_X1 U7909 ( .A1(n8565), .A2(n9771), .ZN(n9792) );
  NAND2_X1 U7910 ( .A1(n9793), .A2(n9792), .ZN(n9791) );
  OR2_X1 U7911 ( .A1(n9989), .A2(n9412), .ZN(n6613) );
  NAND2_X1 U7912 ( .A1(n7772), .A2(n6490), .ZN(n6618) );
  AOI22_X1 U7913 ( .A1(n6405), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n4926), .B2(
        n6616), .ZN(n6617) );
  INV_X1 U7914 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9915) );
  INV_X1 U7915 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n6620) );
  NAND2_X1 U7916 ( .A1(n6621), .A2(n6620), .ZN(n6622) );
  NAND2_X1 U7917 ( .A1(n6630), .A2(n6622), .ZN(n9785) );
  OR2_X1 U7918 ( .A1(n9785), .A2(n6386), .ZN(n6624) );
  AOI22_X1 U7919 ( .A1(n6400), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n6441), .B2(
        P1_REG0_REG_19__SCAN_IN), .ZN(n6623) );
  OAI211_X1 U7920 ( .C1(n6759), .C2(n9915), .A(n6624), .B(n6623), .ZN(n9807)
         );
  OR2_X1 U7921 ( .A1(n9784), .A2(n9807), .ZN(n6625) );
  NAND2_X1 U7922 ( .A1(n9784), .A2(n9807), .ZN(n6626) );
  NAND2_X1 U7923 ( .A1(n7843), .A2(n6490), .ZN(n6629) );
  NAND2_X1 U7924 ( .A1(n6405), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n6628) );
  NAND2_X1 U7925 ( .A1(n6630), .A2(n9433), .ZN(n6631) );
  NAND2_X1 U7926 ( .A1(n6638), .A2(n6631), .ZN(n9765) );
  AOI22_X1 U7927 ( .A1(n6400), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n6441), .B2(
        P1_REG0_REG_20__SCAN_IN), .ZN(n6633) );
  NAND2_X1 U7928 ( .A1(n8491), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n6632) );
  OAI211_X1 U7929 ( .C1(n9765), .C2(n6386), .A(n6633), .B(n6632), .ZN(n9777)
         );
  INV_X1 U7930 ( .A(n9777), .ZN(n9742) );
  OR2_X1 U7931 ( .A1(n9909), .A2(n9742), .ZN(n8572) );
  NAND2_X1 U7932 ( .A1(n9909), .A2(n9742), .ZN(n9738) );
  INV_X1 U7933 ( .A(n9746), .ZN(n6646) );
  NAND2_X1 U7934 ( .A1(n7918), .A2(n6490), .ZN(n6635) );
  NAND2_X1 U7935 ( .A1(n6405), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n6634) );
  INV_X1 U7936 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n6637) );
  NAND2_X1 U7937 ( .A1(n6638), .A2(n6637), .ZN(n6639) );
  NAND2_X1 U7938 ( .A1(n6652), .A2(n6639), .ZN(n9383) );
  OR2_X1 U7939 ( .A1(n9383), .A2(n6386), .ZN(n6644) );
  INV_X1 U7940 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n9905) );
  NAND2_X1 U7941 ( .A1(n6400), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n6641) );
  NAND2_X1 U7942 ( .A1(n6441), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n6640) );
  OAI211_X1 U7943 ( .C1(n6759), .C2(n9905), .A(n6641), .B(n6640), .ZN(n6642)
         );
  INV_X1 U7944 ( .A(n6642), .ZN(n6643) );
  NAND2_X1 U7945 ( .A1(n6644), .A2(n6643), .ZN(n9725) );
  INV_X1 U7946 ( .A(n9725), .ZN(n9763) );
  NAND2_X1 U7947 ( .A1(n7018), .A2(n9763), .ZN(n8573) );
  NAND2_X1 U7948 ( .A1(n7018), .A2(n9725), .ZN(n6647) );
  NAND2_X1 U7949 ( .A1(n7943), .A2(n6490), .ZN(n6649) );
  NAND2_X1 U7950 ( .A1(n6405), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n6648) );
  INV_X1 U7951 ( .A(n6652), .ZN(n6650) );
  INV_X1 U7952 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n6651) );
  NAND2_X1 U7953 ( .A1(n6652), .A2(n6651), .ZN(n6653) );
  NAND2_X1 U7954 ( .A1(n6661), .A2(n6653), .ZN(n9732) );
  OR2_X1 U7955 ( .A1(n9732), .A2(n6386), .ZN(n6658) );
  INV_X1 U7956 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n9900) );
  NAND2_X1 U7957 ( .A1(n6400), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n6655) );
  NAND2_X1 U7958 ( .A1(n6441), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n6654) );
  OAI211_X1 U7959 ( .C1(n9900), .C2(n6759), .A(n6655), .B(n6654), .ZN(n6656)
         );
  INV_X1 U7960 ( .A(n6656), .ZN(n6657) );
  NAND2_X1 U7961 ( .A1(n6658), .A2(n6657), .ZN(n9706) );
  OR2_X1 U7962 ( .A1(n9721), .A2(n9743), .ZN(n8576) );
  NAND2_X1 U7963 ( .A1(n9721), .A2(n9743), .ZN(n8577) );
  NAND2_X1 U7964 ( .A1(n8049), .A2(n6490), .ZN(n6660) );
  NAND2_X1 U7965 ( .A1(n6405), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n6659) );
  INV_X1 U7966 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n9365) );
  NAND2_X1 U7967 ( .A1(n6661), .A2(n9365), .ZN(n6662) );
  NAND2_X1 U7968 ( .A1(n6670), .A2(n6662), .ZN(n9712) );
  OR2_X1 U7969 ( .A1(n9712), .A2(n6386), .ZN(n6667) );
  INV_X1 U7970 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n9895) );
  NAND2_X1 U7971 ( .A1(n6400), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n6664) );
  NAND2_X1 U7972 ( .A1(n6441), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n6663) );
  OAI211_X1 U7973 ( .C1(n9895), .C2(n6759), .A(n6664), .B(n6663), .ZN(n6665)
         );
  INV_X1 U7974 ( .A(n6665), .ZN(n6666) );
  NAND2_X1 U7975 ( .A1(n6667), .A2(n6666), .ZN(n9726) );
  NAND2_X1 U7976 ( .A1(n8111), .A2(n6490), .ZN(n6669) );
  NAND2_X1 U7977 ( .A1(n6405), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n6668) );
  INV_X1 U7978 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9424) );
  NAND2_X1 U7979 ( .A1(n6670), .A2(n9424), .ZN(n6671) );
  AND2_X1 U7980 ( .A1(n6684), .A2(n6671), .ZN(n9696) );
  NAND2_X1 U7981 ( .A1(n9696), .A2(n6579), .ZN(n6676) );
  INV_X1 U7982 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n9890) );
  NAND2_X1 U7983 ( .A1(n6400), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n6673) );
  NAND2_X1 U7984 ( .A1(n6441), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n6672) );
  OAI211_X1 U7985 ( .C1(n9890), .C2(n6759), .A(n6673), .B(n6672), .ZN(n6674)
         );
  INV_X1 U7986 ( .A(n6674), .ZN(n6675) );
  INV_X1 U7987 ( .A(n9707), .ZN(n6677) );
  OR2_X1 U7988 ( .A1(n9695), .A2(n6677), .ZN(n8645) );
  NAND2_X1 U7989 ( .A1(n9695), .A2(n6677), .ZN(n8649) );
  NAND2_X1 U7990 ( .A1(n9695), .A2(n9707), .ZN(n6679) );
  NAND2_X1 U7991 ( .A1(n8225), .A2(n6490), .ZN(n6681) );
  NAND2_X1 U7992 ( .A1(n6405), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n6680) );
  INV_X1 U7993 ( .A(n6684), .ZN(n6682) );
  NAND2_X1 U7994 ( .A1(n6682), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n6698) );
  INV_X1 U7995 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n6683) );
  NAND2_X1 U7996 ( .A1(n6684), .A2(n6683), .ZN(n6685) );
  NAND2_X1 U7997 ( .A1(n6698), .A2(n6685), .ZN(n9678) );
  OR2_X1 U7998 ( .A1(n9678), .A2(n6386), .ZN(n6691) );
  INV_X1 U7999 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n6688) );
  NAND2_X1 U8000 ( .A1(n6400), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n6687) );
  NAND2_X1 U8001 ( .A1(n6441), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n6686) );
  OAI211_X1 U8002 ( .C1(n6759), .C2(n6688), .A(n6687), .B(n6686), .ZN(n6689)
         );
  INV_X1 U8003 ( .A(n6689), .ZN(n6690) );
  NAND2_X1 U8004 ( .A1(n9883), .A2(n9689), .ZN(n6692) );
  NAND2_X1 U8005 ( .A1(n8241), .A2(n6490), .ZN(n6695) );
  NAND2_X1 U8006 ( .A1(n6405), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n6694) );
  INV_X1 U8007 ( .A(n6698), .ZN(n6696) );
  INV_X1 U8008 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n6697) );
  NAND2_X1 U8009 ( .A1(n6698), .A2(n6697), .ZN(n6699) );
  NAND2_X1 U8010 ( .A1(n6719), .A2(n6699), .ZN(n9474) );
  OR2_X1 U8011 ( .A1(n9474), .A2(n6386), .ZN(n6704) );
  INV_X1 U8012 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n9880) );
  NAND2_X1 U8013 ( .A1(n6400), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n6701) );
  NAND2_X1 U8014 ( .A1(n6441), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n6700) );
  OAI211_X1 U8015 ( .C1(n9880), .C2(n6759), .A(n6701), .B(n6700), .ZN(n6702)
         );
  INV_X1 U8016 ( .A(n6702), .ZN(n6703) );
  INV_X1 U8017 ( .A(n9673), .ZN(n9639) );
  OR2_X1 U8018 ( .A1(n9660), .A2(n9639), .ZN(n8656) );
  NAND2_X1 U8019 ( .A1(n9660), .A2(n9639), .ZN(n8654) );
  NAND2_X1 U8020 ( .A1(n8656), .A2(n8654), .ZN(n8630) );
  NAND2_X1 U8021 ( .A1(n9660), .A2(n9673), .ZN(n6705) );
  NAND2_X1 U8022 ( .A1(n8246), .A2(n6490), .ZN(n6707) );
  NAND2_X1 U8023 ( .A1(n6405), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n6706) );
  XNOR2_X1 U8024 ( .A(n6719), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n9646) );
  NAND2_X1 U8025 ( .A1(n9646), .A2(n6579), .ZN(n6712) );
  INV_X1 U8026 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n9875) );
  NAND2_X1 U8027 ( .A1(n6400), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n6709) );
  NAND2_X1 U8028 ( .A1(n6441), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n6708) );
  OAI211_X1 U8029 ( .C1(n9875), .C2(n6759), .A(n6709), .B(n6708), .ZN(n6710)
         );
  INV_X1 U8030 ( .A(n6710), .ZN(n6711) );
  INV_X1 U8031 ( .A(n9656), .ZN(n6713) );
  NAND2_X1 U8032 ( .A1(n9645), .A2(n6713), .ZN(n8638) );
  OR2_X1 U8033 ( .A1(n9645), .A2(n6713), .ZN(n8658) );
  NAND2_X1 U8034 ( .A1(n9343), .A2(n6490), .ZN(n6715) );
  NAND2_X1 U8035 ( .A1(n6405), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n6714) );
  INV_X1 U8036 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n6717) );
  INV_X1 U8037 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n6716) );
  OAI21_X1 U8038 ( .B1(n6719), .B2(n6717), .A(n6716), .ZN(n6720) );
  NAND2_X1 U8039 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n6718) );
  INV_X1 U8040 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n6723) );
  NAND2_X1 U8041 ( .A1(n6400), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n6722) );
  NAND2_X1 U8042 ( .A1(n6441), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n6721) );
  OAI211_X1 U8043 ( .C1(n6723), .C2(n6759), .A(n6722), .B(n6721), .ZN(n6724)
         );
  AOI21_X1 U8044 ( .B1(n9626), .B2(n6579), .A(n6724), .ZN(n9640) );
  NAND2_X1 U8045 ( .A1(n9628), .A2(n9499), .ZN(n8659) );
  NOR2_X1 U8046 ( .A1(n6725), .A2(n8632), .ZN(n6801) );
  AND2_X1 U8047 ( .A1(n6725), .A2(n8632), .ZN(n6726) );
  OR2_X1 U8048 ( .A1(n6801), .A2(n6726), .ZN(n9629) );
  NAND2_X1 U8049 ( .A1(n6737), .A2(n6730), .ZN(n6731) );
  OR2_X1 U8050 ( .A1(n6734), .A2(n6509), .ZN(n6736) );
  NAND2_X1 U8051 ( .A1(n6888), .A2(n6738), .ZN(n8730) );
  NAND2_X1 U8052 ( .A1(n6738), .A2(n8739), .ZN(n6884) );
  NAND2_X1 U8053 ( .A1(n8730), .A2(n6884), .ZN(n6739) );
  AND2_X1 U8054 ( .A1(n6883), .A2(n6739), .ZN(n6740) );
  OR2_X1 U8055 ( .A1(n8671), .A2(n8730), .ZN(n10515) );
  NAND2_X1 U8056 ( .A1(n6740), .A2(n10515), .ZN(n7517) );
  OR2_X1 U8057 ( .A1(n8599), .A2(n6738), .ZN(n8680) );
  OR2_X1 U8058 ( .A1(n8680), .A2(n8739), .ZN(n10613) );
  INV_X1 U8059 ( .A(n10518), .ZN(n8606) );
  AND2_X1 U8060 ( .A1(n6895), .A2(n8606), .ZN(n8607) );
  NAND2_X1 U8061 ( .A1(n10539), .A2(n8683), .ZN(n6744) );
  INV_X1 U8062 ( .A(n6745), .ZN(n8608) );
  INV_X1 U8063 ( .A(n9511), .ZN(n7512) );
  NAND2_X1 U8064 ( .A1(n7512), .A2(n7547), .ZN(n8512) );
  INV_X1 U8065 ( .A(n7547), .ZN(n10593) );
  NAND2_X1 U8066 ( .A1(n9511), .A2(n10593), .ZN(n8499) );
  NAND2_X1 U8067 ( .A1(n7540), .A2(n8512), .ZN(n7394) );
  NAND2_X1 U8068 ( .A1(n7394), .A2(n8610), .ZN(n7393) );
  NAND2_X1 U8069 ( .A1(n7393), .A2(n8501), .ZN(n7576) );
  INV_X1 U8070 ( .A(n8506), .ZN(n8695) );
  NAND2_X1 U8071 ( .A1(n8525), .A2(n7645), .ZN(n8520) );
  NAND2_X1 U8072 ( .A1(n8508), .A2(n8505), .ZN(n8518) );
  NOR2_X1 U8073 ( .A1(n8520), .A2(n8518), .ZN(n8694) );
  NAND2_X1 U8074 ( .A1(n7631), .A2(n8694), .ZN(n6748) );
  AND2_X1 U8075 ( .A1(n8510), .A2(n8516), .ZN(n6746) );
  AND2_X1 U8076 ( .A1(n8698), .A2(n8526), .ZN(n6747) );
  NAND2_X1 U8077 ( .A1(n6748), .A2(n6747), .ZN(n7594) );
  INV_X1 U8078 ( .A(n8618), .ZN(n7595) );
  INV_X1 U8079 ( .A(n9504), .ZN(n8203) );
  NAND2_X1 U8080 ( .A1(n9858), .A2(n8203), .ZN(n8530) );
  INV_X1 U8081 ( .A(n9503), .ZN(n9443) );
  OR2_X1 U8082 ( .A1(n8542), .A2(n9443), .ZN(n8701) );
  NAND2_X1 U8083 ( .A1(n8542), .A2(n9443), .ZN(n8704) );
  NAND2_X1 U8084 ( .A1(n6749), .A2(n8621), .ZN(n7797) );
  INV_X1 U8085 ( .A(n9502), .ZN(n9357) );
  OR2_X1 U8086 ( .A1(n9846), .A2(n9357), .ZN(n8707) );
  NAND2_X1 U8087 ( .A1(n9846), .A2(n9357), .ZN(n8705) );
  NAND2_X1 U8088 ( .A1(n7936), .A2(n8622), .ZN(n6750) );
  INV_X1 U8089 ( .A(n8711), .ZN(n6751) );
  AND2_X1 U8090 ( .A1(n8714), .A2(n9813), .ZN(n8712) );
  NAND2_X1 U8091 ( .A1(n9812), .A2(n8712), .ZN(n9817) );
  NAND2_X1 U8092 ( .A1(n9817), .A2(n8716), .ZN(n8192) );
  INV_X1 U8093 ( .A(n8626), .ZN(n8560) );
  NAND2_X1 U8094 ( .A1(n8192), .A2(n8560), .ZN(n8191) );
  NAND2_X1 U8095 ( .A1(n8191), .A2(n8718), .ZN(n9805) );
  INV_X1 U8096 ( .A(n9792), .ZN(n9806) );
  INV_X1 U8097 ( .A(n9807), .ZN(n9761) );
  INV_X1 U8098 ( .A(n9771), .ZN(n8719) );
  INV_X1 U8099 ( .A(n8721), .ZN(n6752) );
  INV_X1 U8100 ( .A(n9738), .ZN(n8568) );
  NAND2_X1 U8101 ( .A1(n8721), .A2(n8568), .ZN(n6753) );
  AND2_X1 U8102 ( .A1(n6753), .A2(n8573), .ZN(n8642) );
  INV_X1 U8103 ( .A(n9726), .ZN(n9425) );
  OR2_X1 U8104 ( .A1(n9711), .A2(n9425), .ZN(n8578) );
  NAND2_X1 U8105 ( .A1(n9711), .A2(n9425), .ZN(n8648) );
  NAND2_X1 U8106 ( .A1(n9704), .A2(n9703), .ZN(n6754) );
  OR2_X1 U8107 ( .A1(n9883), .A2(n9476), .ZN(n8650) );
  NAND2_X1 U8108 ( .A1(n9883), .A2(n9476), .ZN(n8653) );
  NAND2_X1 U8109 ( .A1(n8650), .A2(n8653), .ZN(n9667) );
  NAND2_X1 U8110 ( .A1(n9670), .A2(n8653), .ZN(n9654) );
  XNOR2_X1 U8111 ( .A(n6813), .B(n6812), .ZN(n6764) );
  NAND2_X1 U8112 ( .A1(n4926), .A2(n8739), .ZN(n6755) );
  INV_X1 U8113 ( .A(n6828), .ZN(n6761) );
  INV_X1 U8114 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n6758) );
  NAND2_X1 U8115 ( .A1(n6441), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6757) );
  NAND2_X1 U8116 ( .A1(n6400), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n6756) );
  OAI211_X1 U8117 ( .C1(n6759), .C2(n6758), .A(n6757), .B(n6756), .ZN(n6760)
         );
  AOI21_X1 U8118 ( .B1(n6761), .B2(n6579), .A(n6760), .ZN(n8753) );
  INV_X1 U8119 ( .A(n7174), .ZN(n10013) );
  NOR2_X2 U8120 ( .A1(n10013), .A2(n8671), .ZN(n10543) );
  NAND2_X1 U8121 ( .A1(n9656), .A2(n10541), .ZN(n6762) );
  OAI21_X1 U8122 ( .B1(n8753), .B2(n9764), .A(n6762), .ZN(n6763) );
  AOI21_X1 U8123 ( .B1(n6764), .B2(n10546), .A(n6763), .ZN(n9634) );
  INV_X1 U8124 ( .A(n7684), .ZN(n7734) );
  INV_X1 U8125 ( .A(n7638), .ZN(n10630) );
  INV_X1 U8126 ( .A(n8542), .ZN(n7838) );
  NAND2_X1 U8127 ( .A1(n9825), .A2(n9994), .ZN(n9824) );
  NOR2_X2 U8128 ( .A1(n9925), .A2(n9824), .ZN(n9794) );
  OR2_X2 U8129 ( .A1(n9721), .A2(n9749), .ZN(n9719) );
  NOR2_X2 U8130 ( .A1(n9711), .A2(n9719), .ZN(n9710) );
  NAND2_X1 U8131 ( .A1(n9968), .A2(n9710), .ZN(n9692) );
  OR2_X2 U8132 ( .A1(n9883), .A2(n9692), .ZN(n9675) );
  INV_X1 U8133 ( .A(n6883), .ZN(n10519) );
  OAI211_X1 U8134 ( .C1(n9628), .C2(n9644), .A(n10537), .B(n4959), .ZN(n9625)
         );
  NOR2_X1 U8135 ( .A1(P1_D_REG_31__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .ZN(
        n6768) );
  NOR4_X1 U8136 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_29__SCAN_IN), .A4(P1_D_REG_28__SCAN_IN), .ZN(n6767) );
  NOR4_X1 U8137 ( .A1(P1_D_REG_23__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_21__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n6766) );
  NOR4_X1 U8138 ( .A1(P1_D_REG_27__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_25__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n6765) );
  NAND4_X1 U8139 ( .A1(n6768), .A2(n6767), .A3(n6766), .A4(n6765), .ZN(n6782)
         );
  NOR4_X1 U8140 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n6772) );
  NOR4_X1 U8141 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n6771) );
  NOR4_X1 U8142 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n6770) );
  NOR4_X1 U8143 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n6769) );
  NAND4_X1 U8144 ( .A1(n6772), .A2(n6771), .A3(n6770), .A4(n6769), .ZN(n6781)
         );
  NAND2_X1 U8145 ( .A1(n6776), .A2(n6773), .ZN(n6774) );
  XNOR2_X1 U8146 ( .A(n6776), .B(P1_IR_REG_25__SCAN_IN), .ZN(n8226) );
  INV_X1 U8147 ( .A(n8226), .ZN(n6783) );
  NAND2_X1 U8148 ( .A1(n6783), .A2(P1_B_REG_SCAN_IN), .ZN(n6779) );
  NAND2_X1 U8149 ( .A1(n6777), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6778) );
  MUX2_X1 U8150 ( .A(n6779), .B(P1_B_REG_SCAN_IN), .S(n8112), .Z(n6780) );
  OAI21_X1 U8151 ( .B1(n6782), .B2(n6781), .A(n6792), .ZN(n7077) );
  INV_X1 U8152 ( .A(n8730), .ZN(n6793) );
  OR2_X1 U8153 ( .A1(n8671), .A2(n6793), .ZN(n7093) );
  NAND2_X1 U8154 ( .A1(n7077), .A2(n7093), .ZN(n6806) );
  AOI21_X1 U8155 ( .B1(n4926), .B2(n10537), .A(n6806), .ZN(n6789) );
  INV_X1 U8156 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n10278) );
  INV_X1 U8157 ( .A(n6786), .ZN(n6791) );
  AND2_X1 U8158 ( .A1(n6791), .A2(n6783), .ZN(n6784) );
  NAND2_X1 U8159 ( .A1(n6787), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6788) );
  NOR2_X1 U8160 ( .A1(n7078), .A2(n10279), .ZN(n10277) );
  INV_X1 U8161 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n7148) );
  INV_X1 U8162 ( .A(n8112), .ZN(n6790) );
  AND2_X1 U8163 ( .A1(n6791), .A2(n6790), .ZN(n7150) );
  NAND2_X1 U8164 ( .A1(n6795), .A2(n6794), .ZN(P1_U3550) );
  INV_X1 U8165 ( .A(n7079), .ZN(n6808) );
  NAND2_X1 U8166 ( .A1(n8755), .A2(n6798), .ZN(n6799) );
  NAND2_X1 U8167 ( .A1(n6800), .A2(n6799), .ZN(P1_U3518) );
  INV_X1 U8168 ( .A(n9628), .ZN(n8755) );
  NAND2_X1 U8169 ( .A1(n6802), .A2(n6490), .ZN(n6804) );
  NAND2_X1 U8170 ( .A1(n6405), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n6803) );
  NAND2_X1 U8171 ( .A1(n6804), .A2(n6803), .ZN(n6823) );
  NAND2_X1 U8172 ( .A1(n6823), .A2(n8753), .ZN(n8665) );
  NAND2_X1 U8173 ( .A1(n8660), .A2(n8665), .ZN(n8604) );
  INV_X1 U8174 ( .A(n6806), .ZN(n6807) );
  INV_X1 U8175 ( .A(n10279), .ZN(n7149) );
  NAND4_X1 U8176 ( .A1(n6808), .A2(n6807), .A3(n7149), .A4(n7078), .ZN(n6825)
         );
  NOR2_X1 U8177 ( .A1(n10279), .A2(n6738), .ZN(n6809) );
  NOR2_X1 U8178 ( .A1(n6889), .A2(n8680), .ZN(n6810) );
  NAND2_X1 U8179 ( .A1(n10524), .A2(n6810), .ZN(n7588) );
  INV_X1 U8180 ( .A(n7517), .ZN(n7635) );
  NAND2_X1 U8181 ( .A1(n10524), .A2(n7635), .ZN(n6811) );
  INV_X1 U8182 ( .A(n9525), .ZN(n8247) );
  NAND2_X1 U8183 ( .A1(n8247), .A2(P1_B_REG_SCAN_IN), .ZN(n6816) );
  AND2_X1 U8184 ( .A1(n10543), .A2(n6816), .ZN(n9615) );
  NAND2_X1 U8185 ( .A1(n8491), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n6819) );
  NAND2_X1 U8186 ( .A1(n6400), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n6818) );
  NAND2_X1 U8187 ( .A1(n6441), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n6817) );
  NAND3_X1 U8188 ( .A1(n6819), .A2(n6818), .A3(n6817), .ZN(n9498) );
  AOI21_X1 U8189 ( .B1(n6823), .B2(n4959), .A(n9797), .ZN(n6824) );
  NAND2_X1 U8190 ( .A1(n6836), .A2(n4924), .ZN(n6831) );
  OR2_X1 U8191 ( .A1(n6883), .A2(n6888), .ZN(n7083) );
  INV_X1 U8192 ( .A(n7083), .ZN(n6826) );
  INV_X1 U8193 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n6827) );
  OAI22_X1 U8194 ( .A1(n6828), .A2(n9854), .B1(n6827), .B2(n10524), .ZN(n6829)
         );
  AOI21_X1 U8195 ( .B1(n6823), .B2(n10552), .A(n6829), .ZN(n6830) );
  OAI21_X1 U8196 ( .B1(n6838), .B2(n9800), .A(n6832), .ZN(n6833) );
  INV_X1 U8197 ( .A(n6833), .ZN(n6834) );
  AOI21_X1 U8198 ( .B1(n10610), .B2(n6823), .A(n6836), .ZN(n6837) );
  INV_X1 U8199 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n6841) );
  OR2_X1 U8200 ( .A1(n10681), .A2(n6841), .ZN(n6842) );
  NAND2_X1 U8201 ( .A1(n6843), .A2(n10677), .ZN(n6845) );
  OR2_X1 U8202 ( .A1(n10677), .A2(n6758), .ZN(n6844) );
  NAND2_X1 U8203 ( .A1(n6845), .A2(n6844), .ZN(P1_U3551) );
  NOR2_X1 U8204 ( .A1(n8441), .A2(n10684), .ZN(n6849) );
  OR2_X1 U8205 ( .A1(n7406), .A2(n6849), .ZN(n6851) );
  AOI22_X1 U8206 ( .A1(n6852), .A2(n6851), .B1(n7135), .B2(n6850), .ZN(n6854)
         );
  INV_X1 U8207 ( .A(n6855), .ZN(n6869) );
  OR2_X1 U8208 ( .A1(n10761), .A2(n6856), .ZN(n6857) );
  INV_X1 U8209 ( .A(n6864), .ZN(n6860) );
  NAND2_X1 U8210 ( .A1(n5522), .A2(n8254), .ZN(n7448) );
  NAND2_X1 U8211 ( .A1(n7433), .A2(n7448), .ZN(n6863) );
  NAND2_X1 U8212 ( .A1(n7442), .A2(n6863), .ZN(n6866) );
  NAND2_X1 U8213 ( .A1(n7423), .A2(n9240), .ZN(n7440) );
  NAND2_X1 U8214 ( .A1(n7450), .A2(n7440), .ZN(n6865) );
  NAND2_X1 U8215 ( .A1(n6868), .A2(n7430), .ZN(n9327) );
  XNOR2_X1 U8216 ( .A(n6875), .B(n8797), .ZN(n6876) );
  XNOR2_X1 U8217 ( .A(n6877), .B(n8797), .ZN(n9038) );
  INV_X1 U8218 ( .A(n9045), .ZN(n9254) );
  NAND2_X1 U8219 ( .A1(n9045), .A2(n6880), .ZN(n6881) );
  INV_X2 U8220 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  NAND2_X1 U8221 ( .A1(n6889), .A2(n4926), .ZN(n6885) );
  AND2_X1 U8222 ( .A1(n6888), .A2(n6884), .ZN(n6886) );
  INV_X1 U8223 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n6892) );
  INV_X1 U8224 ( .A(n6893), .ZN(n6894) );
  OAI21_X1 U8225 ( .B1(n6936), .B2(n10518), .A(n6894), .ZN(n7213) );
  OAI222_X1 U8226 ( .A1(n8744), .A2(n10518), .B1(n8743), .B2(n6895), .C1(n6890), .C2(n9526), .ZN(n7212) );
  AOI21_X1 U8227 ( .B1(n7213), .B2(n7212), .A(n6897), .ZN(n7231) );
  AND2_X1 U8228 ( .A1(n6900), .A2(n6899), .ZN(n6901) );
  XNOR2_X1 U8229 ( .A(n6901), .B(n6996), .ZN(n7232) );
  AOI22_X1 U8230 ( .A1(n10542), .A2(n7069), .B1(n6919), .B2(n7366), .ZN(n7230)
         );
  AOI21_X1 U8231 ( .B1(n7231), .B2(n7232), .A(n7230), .ZN(n6904) );
  NOR2_X1 U8232 ( .A1(n7232), .A2(n7231), .ZN(n6903) );
  NOR2_X1 U8233 ( .A1(n6904), .A2(n6903), .ZN(n7239) );
  NAND2_X1 U8234 ( .A1(n10553), .A2(n6915), .ZN(n6906) );
  NAND2_X1 U8235 ( .A1(n9512), .A2(n6919), .ZN(n6905) );
  NAND2_X1 U8236 ( .A1(n6906), .A2(n6905), .ZN(n6907) );
  NAND2_X1 U8237 ( .A1(n9512), .A2(n7069), .ZN(n6909) );
  NAND2_X1 U8238 ( .A1(n10553), .A2(n6919), .ZN(n6908) );
  NAND2_X1 U8239 ( .A1(n6909), .A2(n6908), .ZN(n6910) );
  AND2_X1 U8240 ( .A1(n6911), .A2(n6910), .ZN(n6912) );
  NOR2_X1 U8241 ( .A1(n6911), .A2(n6910), .ZN(n6913) );
  NOR2_X1 U8242 ( .A1(n6912), .A2(n6913), .ZN(n7240) );
  NAND2_X1 U8243 ( .A1(n7239), .A2(n7240), .ZN(n7238) );
  INV_X1 U8244 ( .A(n6913), .ZN(n6914) );
  NAND2_X1 U8245 ( .A1(n7238), .A2(n6914), .ZN(n7248) );
  BUF_X4 U8246 ( .A(n6919), .Z(n7070) );
  NAND2_X1 U8247 ( .A1(n10544), .A2(n7070), .ZN(n6917) );
  NAND2_X1 U8248 ( .A1(n7523), .A2(n6915), .ZN(n6916) );
  NAND2_X1 U8249 ( .A1(n6917), .A2(n6916), .ZN(n6918) );
  AOI22_X1 U8250 ( .A1(n10544), .A2(n7069), .B1(n6919), .B2(n7523), .ZN(n6922)
         );
  NAND2_X1 U8251 ( .A1(n7248), .A2(n7249), .ZN(n7247) );
  NAND2_X1 U8252 ( .A1(n7247), .A2(n6923), .ZN(n7305) );
  INV_X1 U8253 ( .A(n7305), .ZN(n6933) );
  NAND2_X1 U8254 ( .A1(n9511), .A2(n7070), .ZN(n6925) );
  NAND2_X1 U8255 ( .A1(n7547), .A2(n6915), .ZN(n6924) );
  NAND2_X1 U8256 ( .A1(n6925), .A2(n6924), .ZN(n6926) );
  XNOR2_X1 U8257 ( .A(n6926), .B(n8745), .ZN(n6928) );
  AOI22_X1 U8258 ( .A1(n9511), .A2(n7069), .B1(n7070), .B2(n7547), .ZN(n6929)
         );
  XNOR2_X1 U8259 ( .A(n6928), .B(n6929), .ZN(n6931) );
  AOI22_X1 U8260 ( .A1(n9510), .A2(n7070), .B1(n7491), .B2(n6915), .ZN(n6927)
         );
  OR2_X1 U8261 ( .A1(n6929), .A2(n6928), .ZN(n6934) );
  OR2_X1 U8262 ( .A1(n4949), .A2(n6934), .ZN(n6930) );
  AOI22_X1 U8263 ( .A1(n9510), .A2(n7069), .B1(n7070), .B2(n7491), .ZN(n7379)
         );
  AND2_X1 U8264 ( .A1(n4949), .A2(n6934), .ZN(n6935) );
  NAND2_X1 U8265 ( .A1(n10609), .A2(n7067), .ZN(n6938) );
  NAND2_X1 U8266 ( .A1(n9509), .A2(n7070), .ZN(n6937) );
  NAND2_X1 U8267 ( .A1(n6938), .A2(n6937), .ZN(n6939) );
  XNOR2_X1 U8268 ( .A(n6939), .B(n8745), .ZN(n6941) );
  AOI22_X1 U8269 ( .A1(n10609), .A2(n7070), .B1(n9509), .B2(n7069), .ZN(n6940)
         );
  NAND2_X1 U8270 ( .A1(n6941), .A2(n6940), .ZN(n7459) );
  OR2_X1 U8271 ( .A1(n6941), .A2(n6940), .ZN(n7460) );
  OAI22_X1 U8272 ( .A1(n7734), .A2(n8744), .B1(n7826), .B2(n8743), .ZN(n6943)
         );
  INV_X1 U8273 ( .A(n6943), .ZN(n7470) );
  AOI22_X1 U8274 ( .A1(n7684), .A2(n7067), .B1(n7070), .B2(n9508), .ZN(n6942)
         );
  XNOR2_X1 U8275 ( .A(n6942), .B(n8745), .ZN(n7471) );
  AOI22_X1 U8276 ( .A1(n7638), .A2(n7067), .B1(n6919), .B2(n9507), .ZN(n6944)
         );
  XNOR2_X1 U8277 ( .A(n6944), .B(n8745), .ZN(n6945) );
  AOI22_X1 U8278 ( .A1(n7638), .A2(n7070), .B1(n7069), .B2(n9507), .ZN(n7821)
         );
  AOI22_X1 U8279 ( .A1(n7657), .A2(n7070), .B1(n7069), .B2(n9506), .ZN(n6951)
         );
  NAND2_X1 U8280 ( .A1(n7657), .A2(n7067), .ZN(n6949) );
  NAND2_X1 U8281 ( .A1(n9506), .A2(n7070), .ZN(n6948) );
  NAND2_X1 U8282 ( .A1(n6949), .A2(n6948), .ZN(n6950) );
  XNOR2_X1 U8283 ( .A(n6950), .B(n8745), .ZN(n6952) );
  XOR2_X1 U8284 ( .A(n6951), .B(n6952), .Z(n7856) );
  NAND2_X1 U8285 ( .A1(n6952), .A2(n6951), .ZN(n6953) );
  NAND2_X1 U8286 ( .A1(n7855), .A2(n6953), .ZN(n6957) );
  INV_X1 U8287 ( .A(n6957), .ZN(n6955) );
  AOI22_X1 U8288 ( .A1(n7961), .A2(n7067), .B1(n6919), .B2(n9505), .ZN(n6954)
         );
  XOR2_X1 U8289 ( .A(n8745), .B(n6954), .Z(n6956) );
  NAND2_X1 U8290 ( .A1(n6955), .A2(n5078), .ZN(n6958) );
  INV_X1 U8291 ( .A(n7961), .ZN(n10670) );
  OAI22_X1 U8292 ( .A1(n10670), .A2(n8744), .B1(n7860), .B2(n8743), .ZN(n7954)
         );
  INV_X1 U8293 ( .A(n7954), .ZN(n6959) );
  NAND2_X1 U8294 ( .A1(n9858), .A2(n7067), .ZN(n6962) );
  NAND2_X1 U8295 ( .A1(n9504), .A2(n7070), .ZN(n6961) );
  NAND2_X1 U8296 ( .A1(n6962), .A2(n6961), .ZN(n6963) );
  XNOR2_X1 U8297 ( .A(n6963), .B(n6996), .ZN(n6966) );
  NAND2_X1 U8298 ( .A1(n9858), .A2(n7070), .ZN(n6965) );
  NAND2_X1 U8299 ( .A1(n9504), .A2(n7069), .ZN(n6964) );
  NAND2_X1 U8300 ( .A1(n6965), .A2(n6964), .ZN(n6967) );
  NAND2_X1 U8301 ( .A1(n6966), .A2(n6967), .ZN(n8141) );
  INV_X1 U8302 ( .A(n6966), .ZN(n6969) );
  INV_X1 U8303 ( .A(n6967), .ZN(n6968) );
  NAND2_X1 U8304 ( .A1(n6969), .A2(n6968), .ZN(n8140) );
  NAND2_X1 U8305 ( .A1(n8138), .A2(n8140), .ZN(n8197) );
  AOI22_X1 U8306 ( .A1(n8542), .A2(n7070), .B1(n7069), .B2(n9503), .ZN(n6974)
         );
  NAND2_X1 U8307 ( .A1(n8542), .A2(n7067), .ZN(n6971) );
  NAND2_X1 U8308 ( .A1(n9503), .A2(n7070), .ZN(n6970) );
  NAND2_X1 U8309 ( .A1(n6971), .A2(n6970), .ZN(n6972) );
  XNOR2_X1 U8310 ( .A(n6972), .B(n8745), .ZN(n6973) );
  XOR2_X1 U8311 ( .A(n6974), .B(n6973), .Z(n8198) );
  NAND2_X1 U8312 ( .A1(n6973), .A2(n6974), .ZN(n6975) );
  AOI22_X1 U8313 ( .A1(n9846), .A2(n7070), .B1(n7069), .B2(n9502), .ZN(n6979)
         );
  NAND2_X1 U8314 ( .A1(n9846), .A2(n7067), .ZN(n6977) );
  NAND2_X1 U8315 ( .A1(n9502), .A2(n7070), .ZN(n6976) );
  NAND2_X1 U8316 ( .A1(n6977), .A2(n6976), .ZN(n6978) );
  XNOR2_X1 U8317 ( .A(n6978), .B(n8745), .ZN(n6980) );
  XOR2_X1 U8318 ( .A(n6979), .B(n6980), .Z(n9440) );
  NAND2_X1 U8319 ( .A1(n6980), .A2(n6979), .ZN(n6981) );
  AOI22_X1 U8320 ( .A1(n9943), .A2(n7067), .B1(n6919), .B2(n9501), .ZN(n6982)
         );
  XOR2_X1 U8321 ( .A(n8745), .B(n6982), .Z(n9351) );
  AOI22_X1 U8322 ( .A1(n9943), .A2(n7070), .B1(n7069), .B2(n9501), .ZN(n9350)
         );
  AOI22_X1 U8323 ( .A1(n9998), .A2(n7067), .B1(n6919), .B2(n9820), .ZN(n6983)
         );
  XOR2_X1 U8324 ( .A(n8745), .B(n6983), .Z(n9483) );
  AOI22_X1 U8325 ( .A1(n9998), .A2(n7070), .B1(n7069), .B2(n9820), .ZN(n9482)
         );
  OAI21_X1 U8326 ( .B1(n9481), .B2(n9483), .A(n9482), .ZN(n6985) );
  NAND2_X1 U8327 ( .A1(n6985), .A2(n6984), .ZN(n9397) );
  AOI22_X1 U8328 ( .A1(n9830), .A2(n7070), .B1(n7069), .B2(n9500), .ZN(n6990)
         );
  NAND2_X1 U8329 ( .A1(n9830), .A2(n7067), .ZN(n6987) );
  NAND2_X1 U8330 ( .A1(n9500), .A2(n7070), .ZN(n6986) );
  NAND2_X1 U8331 ( .A1(n6987), .A2(n6986), .ZN(n6988) );
  XNOR2_X1 U8332 ( .A(n6988), .B(n8745), .ZN(n6989) );
  XOR2_X1 U8333 ( .A(n6990), .B(n6989), .Z(n9398) );
  INV_X1 U8334 ( .A(n6989), .ZN(n6992) );
  INV_X1 U8335 ( .A(n6990), .ZN(n6991) );
  NOR2_X1 U8336 ( .A1(n6992), .A2(n6991), .ZN(n6993) );
  AOI21_X1 U8337 ( .B1(n9397), .B2(n9398), .A(n6993), .ZN(n9406) );
  NAND2_X1 U8338 ( .A1(n9925), .A2(n7067), .ZN(n6995) );
  NAND2_X1 U8339 ( .A1(n9819), .A2(n7070), .ZN(n6994) );
  NAND2_X1 U8340 ( .A1(n6995), .A2(n6994), .ZN(n6997) );
  XNOR2_X1 U8341 ( .A(n6997), .B(n6996), .ZN(n9407) );
  NAND2_X1 U8342 ( .A1(n9925), .A2(n6919), .ZN(n6999) );
  NAND2_X1 U8343 ( .A1(n9819), .A2(n7069), .ZN(n6998) );
  NAND2_X1 U8344 ( .A1(n6999), .A2(n6998), .ZN(n9408) );
  NAND2_X1 U8345 ( .A1(n9406), .A2(n7000), .ZN(n7002) );
  NAND2_X1 U8346 ( .A1(n9407), .A2(n9408), .ZN(n7001) );
  OAI22_X1 U8347 ( .A1(n9989), .A2(n6936), .B1(n9412), .B2(n8744), .ZN(n7003)
         );
  XOR2_X1 U8348 ( .A(n8745), .B(n7003), .Z(n9459) );
  OAI22_X1 U8349 ( .A1(n9989), .A2(n8744), .B1(n9412), .B2(n8743), .ZN(n9460)
         );
  NAND2_X1 U8350 ( .A1(n9784), .A2(n7067), .ZN(n7005) );
  NAND2_X1 U8351 ( .A1(n9807), .A2(n7070), .ZN(n7004) );
  NAND2_X1 U8352 ( .A1(n7005), .A2(n7004), .ZN(n7006) );
  XNOR2_X1 U8353 ( .A(n7006), .B(n8745), .ZN(n7009) );
  AND2_X1 U8354 ( .A1(n9807), .A2(n7069), .ZN(n7007) );
  AOI21_X1 U8355 ( .B1(n9784), .B2(n7070), .A(n7007), .ZN(n7008) );
  NAND2_X1 U8356 ( .A1(n7009), .A2(n7008), .ZN(n7010) );
  OAI21_X1 U8357 ( .B1(n7009), .B2(n7008), .A(n7010), .ZN(n9371) );
  AOI22_X1 U8358 ( .A1(n9909), .A2(n7070), .B1(n7069), .B2(n9777), .ZN(n7020)
         );
  NAND2_X1 U8359 ( .A1(n9909), .A2(n7067), .ZN(n7012) );
  NAND2_X1 U8360 ( .A1(n9777), .A2(n6919), .ZN(n7011) );
  NAND2_X1 U8361 ( .A1(n7012), .A2(n7011), .ZN(n7013) );
  XNOR2_X1 U8362 ( .A(n7013), .B(n8745), .ZN(n7019) );
  XOR2_X1 U8363 ( .A(n7020), .B(n7019), .Z(n9431) );
  NAND2_X1 U8364 ( .A1(n7018), .A2(n7067), .ZN(n7015) );
  NAND2_X1 U8365 ( .A1(n9725), .A2(n7070), .ZN(n7014) );
  NAND2_X1 U8366 ( .A1(n7015), .A2(n7014), .ZN(n7016) );
  XNOR2_X1 U8367 ( .A(n7016), .B(n8745), .ZN(n7024) );
  AND2_X1 U8368 ( .A1(n9725), .A2(n7069), .ZN(n7017) );
  AOI21_X1 U8369 ( .B1(n7018), .B2(n7070), .A(n7017), .ZN(n7025) );
  XNOR2_X1 U8370 ( .A(n7024), .B(n7025), .ZN(n9378) );
  INV_X1 U8371 ( .A(n7019), .ZN(n7022) );
  INV_X1 U8372 ( .A(n7020), .ZN(n7021) );
  NOR2_X1 U8373 ( .A1(n7022), .A2(n7021), .ZN(n9379) );
  NOR2_X1 U8374 ( .A1(n9378), .A2(n9379), .ZN(n7023) );
  NAND2_X1 U8375 ( .A1(n9377), .A2(n7023), .ZN(n9381) );
  INV_X1 U8376 ( .A(n7024), .ZN(n7027) );
  INV_X1 U8377 ( .A(n7025), .ZN(n7026) );
  NAND2_X1 U8378 ( .A1(n7027), .A2(n7026), .ZN(n7028) );
  AOI22_X1 U8379 ( .A1(n9721), .A2(n7067), .B1(n6919), .B2(n9706), .ZN(n7029)
         );
  XOR2_X1 U8380 ( .A(n8745), .B(n7029), .Z(n7039) );
  OAI22_X1 U8381 ( .A1(n9976), .A2(n8744), .B1(n9743), .B2(n8743), .ZN(n9450)
         );
  NAND2_X1 U8382 ( .A1(n9711), .A2(n7067), .ZN(n7031) );
  NAND2_X1 U8383 ( .A1(n9726), .A2(n6919), .ZN(n7030) );
  NAND2_X1 U8384 ( .A1(n7031), .A2(n7030), .ZN(n7032) );
  XNOR2_X1 U8385 ( .A(n7032), .B(n8745), .ZN(n7034) );
  AND2_X1 U8386 ( .A1(n9726), .A2(n7069), .ZN(n7033) );
  AOI21_X1 U8387 ( .B1(n9711), .B2(n7070), .A(n7033), .ZN(n7035) );
  NAND2_X1 U8388 ( .A1(n7034), .A2(n7035), .ZN(n9418) );
  INV_X1 U8389 ( .A(n7034), .ZN(n7037) );
  INV_X1 U8390 ( .A(n7035), .ZN(n7036) );
  NAND2_X1 U8391 ( .A1(n7037), .A2(n7036), .ZN(n7038) );
  AND2_X1 U8392 ( .A1(n9418), .A2(n7038), .ZN(n9362) );
  INV_X1 U8393 ( .A(n7039), .ZN(n7040) );
  NAND2_X1 U8394 ( .A1(n9695), .A2(n7067), .ZN(n7042) );
  NAND2_X1 U8395 ( .A1(n9707), .A2(n7070), .ZN(n7041) );
  NAND2_X1 U8396 ( .A1(n7042), .A2(n7041), .ZN(n7043) );
  XNOR2_X1 U8397 ( .A(n7043), .B(n8745), .ZN(n7045) );
  AND2_X1 U8398 ( .A1(n9707), .A2(n7069), .ZN(n7044) );
  AOI21_X1 U8399 ( .B1(n9695), .B2(n6919), .A(n7044), .ZN(n7046) );
  NAND2_X1 U8400 ( .A1(n7045), .A2(n7046), .ZN(n7050) );
  INV_X1 U8401 ( .A(n7045), .ZN(n7048) );
  INV_X1 U8402 ( .A(n7046), .ZN(n7047) );
  NAND2_X1 U8403 ( .A1(n7048), .A2(n7047), .ZN(n7049) );
  AOI22_X1 U8404 ( .A1(n9883), .A2(n7070), .B1(n7069), .B2(n9689), .ZN(n7059)
         );
  NAND2_X1 U8405 ( .A1(n9883), .A2(n7067), .ZN(n7052) );
  NAND2_X1 U8406 ( .A1(n9689), .A2(n6919), .ZN(n7051) );
  NAND2_X1 U8407 ( .A1(n7052), .A2(n7051), .ZN(n7053) );
  XNOR2_X1 U8408 ( .A(n7053), .B(n8745), .ZN(n7058) );
  XOR2_X1 U8409 ( .A(n7059), .B(n7058), .Z(n9390) );
  NAND2_X1 U8410 ( .A1(n9389), .A2(n9390), .ZN(n9388) );
  NAND2_X1 U8411 ( .A1(n9660), .A2(n7067), .ZN(n7055) );
  NAND2_X1 U8412 ( .A1(n9673), .A2(n7070), .ZN(n7054) );
  NAND2_X1 U8413 ( .A1(n7055), .A2(n7054), .ZN(n7056) );
  XNOR2_X1 U8414 ( .A(n7056), .B(n8745), .ZN(n7063) );
  AND2_X1 U8415 ( .A1(n9673), .A2(n7069), .ZN(n7057) );
  AOI21_X1 U8416 ( .B1(n9660), .B2(n6919), .A(n7057), .ZN(n7064) );
  XNOR2_X1 U8417 ( .A(n7063), .B(n7064), .ZN(n9468) );
  INV_X1 U8418 ( .A(n7058), .ZN(n7061) );
  INV_X1 U8419 ( .A(n7059), .ZN(n7060) );
  NOR2_X1 U8420 ( .A1(n7061), .A2(n7060), .ZN(n9469) );
  NOR2_X1 U8421 ( .A1(n9468), .A2(n9469), .ZN(n7062) );
  INV_X1 U8422 ( .A(n9471), .ZN(n7073) );
  INV_X1 U8423 ( .A(n7063), .ZN(n7066) );
  INV_X1 U8424 ( .A(n7064), .ZN(n7065) );
  AND2_X1 U8425 ( .A1(n7066), .A2(n7065), .ZN(n7074) );
  AOI22_X1 U8426 ( .A1(n9645), .A2(n7067), .B1(n6919), .B2(n9656), .ZN(n7068)
         );
  XOR2_X1 U8427 ( .A(n8745), .B(n7068), .Z(n7072) );
  AOI22_X1 U8428 ( .A1(n9645), .A2(n7070), .B1(n7069), .B2(n9656), .ZN(n7071)
         );
  NAND2_X1 U8429 ( .A1(n7072), .A2(n7071), .ZN(n8741) );
  OAI21_X1 U8430 ( .B1(n7072), .B2(n7071), .A(n8741), .ZN(n7075) );
  NOR2_X1 U8431 ( .A1(n7075), .A2(n7074), .ZN(n7076) );
  NAND3_X1 U8432 ( .A1(n7079), .A2(n7078), .A3(n7077), .ZN(n7092) );
  NAND2_X1 U8433 ( .A1(n10669), .A2(n8671), .ZN(n7089) );
  OR2_X1 U8434 ( .A1(n7089), .A2(n10279), .ZN(n7080) );
  AOI21_X1 U8435 ( .B1(n7081), .B2(n8742), .A(n9496), .ZN(n7082) );
  INV_X1 U8436 ( .A(n7082), .ZN(n7100) );
  INV_X1 U8437 ( .A(n7092), .ZN(n7085) );
  NOR2_X1 U8438 ( .A1(n7083), .A2(n10279), .ZN(n7084) );
  NAND2_X1 U8439 ( .A1(n7085), .A2(n7084), .ZN(n7086) );
  OR2_X1 U8440 ( .A1(n10515), .A2(n10279), .ZN(n7090) );
  INV_X1 U8441 ( .A(n7090), .ZN(n8736) );
  NAND2_X1 U8442 ( .A1(n8736), .A2(n7174), .ZN(n7087) );
  NAND2_X1 U8443 ( .A1(n8736), .A2(n10013), .ZN(n7088) );
  AOI22_X1 U8444 ( .A1(n9673), .A2(n9451), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3086), .ZN(n7097) );
  NAND2_X1 U8445 ( .A1(n8599), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7845) );
  NAND3_X1 U8446 ( .A1(n7090), .A2(n7089), .A3(n7845), .ZN(n7091) );
  NAND2_X1 U8447 ( .A1(n7092), .A2(n7091), .ZN(n7095) );
  AND3_X1 U8448 ( .A1(n7093), .A2(n6890), .A3(n7124), .ZN(n7094) );
  NAND2_X1 U8449 ( .A1(n7095), .A2(n7094), .ZN(n7214) );
  NAND2_X1 U8450 ( .A1(n9646), .A2(n9486), .ZN(n7096) );
  OAI211_X1 U8451 ( .C1(n9640), .C2(n9434), .A(n7097), .B(n7096), .ZN(n7098)
         );
  INV_X1 U8452 ( .A(n7098), .ZN(n7099) );
  NAND3_X1 U8453 ( .A1(n7100), .A2(n5519), .A3(n7099), .ZN(P1_U3214) );
  INV_X1 U8454 ( .A(n7101), .ZN(n7102) );
  NOR2_X2 U8455 ( .A1(n6890), .A2(n7102), .ZN(P1_U3973) );
  AOI22_X1 U8456 ( .A1(n10003), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        P1_STATE_REG_SCAN_IN), .B2(n9515), .ZN(n7104) );
  OAI21_X1 U8457 ( .B1(n7106), .B2(n7945), .A(n7104), .ZN(P1_U3354) );
  NOR2_X1 U8458 ( .A1(n8416), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9345) );
  OAI222_X1 U8459 ( .A1(n5696), .A2(P2_U3151), .B1(n8052), .B2(n7106), .C1(
        n7105), .C2(n8237), .ZN(P2_U3294) );
  OAI222_X1 U8460 ( .A1(n4925), .A2(P2_U3151), .B1(n8052), .B2(n7108), .C1(
        n5777), .C2(n8237), .ZN(P2_U3293) );
  AOI22_X1 U8461 ( .A1(n10003), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(
        P1_STATE_REG_SCAN_IN), .B2(n9535), .ZN(n7107) );
  OAI21_X1 U8462 ( .B1(n7108), .B2(n7945), .A(n7107), .ZN(P1_U3353) );
  AOI22_X1 U8463 ( .A1(n10003), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n9558), .B2(
        P1_STATE_REG_SCAN_IN), .ZN(n7109) );
  OAI21_X1 U8464 ( .B1(n7111), .B2(n7945), .A(n7109), .ZN(P1_U3351) );
  OAI222_X1 U8465 ( .A1(n10406), .A2(P2_U3151), .B1(n8052), .B2(n7111), .C1(
        n7110), .C2(n8237), .ZN(P2_U3291) );
  OAI222_X1 U8466 ( .A1(n7334), .A2(P2_U3151), .B1(n8052), .B2(n7113), .C1(
        n5792), .C2(n8237), .ZN(P2_U3292) );
  AOI22_X1 U8467 ( .A1(P2_DATAO_REG_3__SCAN_IN), .A2(n10012), .B1(n9548), .B2(
        P1_STATE_REG_SCAN_IN), .ZN(n7112) );
  OAI21_X1 U8468 ( .B1(n7113), .B2(n7945), .A(n7112), .ZN(P1_U3352) );
  INV_X1 U8469 ( .A(n7114), .ZN(n7117) );
  AOI22_X1 U8470 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9575), .B1(n10012), .B2(
        P2_DATAO_REG_5__SCAN_IN), .ZN(n7115) );
  OAI21_X1 U8471 ( .B1(n7117), .B2(n7945), .A(n7115), .ZN(P1_U3350) );
  INV_X1 U8472 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n7116) );
  OAI222_X1 U8473 ( .A1(n7118), .A2(P2_U3151), .B1(n8052), .B2(n7117), .C1(
        n7116), .C2(n8237), .ZN(P2_U3290) );
  INV_X1 U8474 ( .A(n7119), .ZN(n7134) );
  AOI22_X1 U8475 ( .A1(n9588), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n10012), .ZN(n7120) );
  OAI21_X1 U8476 ( .B1(n7134), .B2(n7945), .A(n7120), .ZN(P1_U3349) );
  INV_X1 U8477 ( .A(n7124), .ZN(n7121) );
  OR2_X1 U8478 ( .A1(n8671), .A2(n7121), .ZN(n7123) );
  NAND2_X1 U8479 ( .A1(n7123), .A2(n7122), .ZN(n7126) );
  OR2_X1 U8480 ( .A1(n7124), .A2(P1_U3086), .ZN(n8738) );
  NAND2_X1 U8481 ( .A1(n10279), .A2(n8738), .ZN(n7127) );
  INV_X1 U8482 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n7132) );
  NOR2_X1 U8483 ( .A1(n7174), .A2(n9525), .ZN(n8735) );
  AOI22_X1 U8484 ( .A1(n8735), .A2(P1_REG2_REG_0__SCAN_IN), .B1(
        P1_REG1_REG_0__SCAN_IN), .B2(n9525), .ZN(n7125) );
  XNOR2_X1 U8485 ( .A(n7125), .B(P1_IR_REG_0__SCAN_IN), .ZN(n7129) );
  INV_X1 U8486 ( .A(n7126), .ZN(n7128) );
  AND2_X1 U8487 ( .A1(n7128), .A2(n7127), .ZN(n7190) );
  NAND2_X1 U8488 ( .A1(n7129), .A2(n7190), .ZN(n7131) );
  NAND2_X1 U8489 ( .A1(P1_U3086), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n7130) );
  OAI211_X1 U8490 ( .C1(n10394), .C2(n7132), .A(n7131), .B(n7130), .ZN(
        P1_U3243) );
  INV_X1 U8491 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n7133) );
  OAI222_X1 U8492 ( .A1(n10435), .A2(P2_U3151), .B1(n8052), .B2(n7134), .C1(
        n7133), .C2(n8237), .ZN(P2_U3289) );
  INV_X1 U8493 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n7138) );
  INV_X1 U8494 ( .A(n7135), .ZN(n7136) );
  NAND2_X1 U8495 ( .A1(n7136), .A2(n7428), .ZN(n7137) );
  OAI21_X1 U8496 ( .B1(n7428), .B2(n7138), .A(n7137), .ZN(P2_U3377) );
  INV_X1 U8497 ( .A(n7139), .ZN(n7144) );
  AOI22_X1 U8498 ( .A1(n10291), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n10012), .ZN(n7140) );
  OAI21_X1 U8499 ( .B1(n7144), .B2(n7945), .A(n7140), .ZN(P1_U3348) );
  INV_X1 U8500 ( .A(n7141), .ZN(n7153) );
  AOI22_X1 U8501 ( .A1(n10295), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n10012), .ZN(n7142) );
  OAI21_X1 U8502 ( .B1(n7153), .B2(n7945), .A(n7142), .ZN(P1_U3347) );
  INV_X1 U8503 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n7143) );
  OAI222_X1 U8504 ( .A1(n7145), .A2(P2_U3151), .B1(n8052), .B2(n7144), .C1(
        n7143), .C2(n8237), .ZN(P2_U3288) );
  INV_X1 U8505 ( .A(n10018), .ZN(n7147) );
  NOR2_X1 U8506 ( .A1(n7147), .A2(P1_D_REG_0__SCAN_IN), .ZN(n7151) );
  OAI22_X1 U8507 ( .A1(n7151), .A2(n7150), .B1(n7149), .B2(n7148), .ZN(
        P1_U3439) );
  OAI222_X1 U8508 ( .A1(n7154), .A2(P2_U3151), .B1(n8052), .B2(n7153), .C1(
        n7152), .C2(n8237), .ZN(P2_U3287) );
  AND2_X1 U8509 ( .A1(n7225), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U8510 ( .A1(n7225), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  AND2_X1 U8511 ( .A1(n7225), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3262) );
  AND2_X1 U8512 ( .A1(n7225), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  AND2_X1 U8513 ( .A1(n7225), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  AND2_X1 U8514 ( .A1(n7225), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U8515 ( .A1(n7225), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U8516 ( .A1(n7225), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U8517 ( .A1(n7225), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  AND2_X1 U8518 ( .A1(n7225), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  INV_X1 U8519 ( .A(n10394), .ZN(n9607) );
  NOR2_X1 U8520 ( .A1(n9607), .A2(P1_U3973), .ZN(P1_U3085) );
  INV_X1 U8521 ( .A(n6461), .ZN(n7201) );
  AOI22_X1 U8522 ( .A1(n7354), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n10012), .ZN(n7156) );
  OAI21_X1 U8523 ( .B1(n7201), .B2(n7945), .A(n7156), .ZN(P1_U3346) );
  NAND2_X1 U8524 ( .A1(n7190), .A2(n8735), .ZN(n10383) );
  NOR2_X1 U8525 ( .A1(n7354), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n7157) );
  AOI21_X1 U8526 ( .B1(P1_REG2_REG_9__SCAN_IN), .B2(n7354), .A(n7157), .ZN(
        n7173) );
  INV_X1 U8527 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n7158) );
  MUX2_X1 U8528 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n7158), .S(n9535), .Z(n9541)
         );
  INV_X1 U8529 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n7159) );
  MUX2_X1 U8530 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n7159), .S(n9515), .Z(n9518)
         );
  AND2_X1 U8531 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n9517) );
  NAND2_X1 U8532 ( .A1(n9518), .A2(n9517), .ZN(n9516) );
  NAND2_X1 U8533 ( .A1(n9515), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n7160) );
  NAND2_X1 U8534 ( .A1(n9516), .A2(n7160), .ZN(n9540) );
  NAND2_X1 U8535 ( .A1(n9541), .A2(n9540), .ZN(n9539) );
  NAND2_X1 U8536 ( .A1(n9535), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n7161) );
  NAND2_X1 U8537 ( .A1(n9539), .A2(n7161), .ZN(n9553) );
  INV_X1 U8538 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n7518) );
  XNOR2_X1 U8539 ( .A(n9548), .B(n7518), .ZN(n9554) );
  NAND2_X1 U8540 ( .A1(n9553), .A2(n9554), .ZN(n9552) );
  NAND2_X1 U8541 ( .A1(n9548), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n7162) );
  NAND2_X1 U8542 ( .A1(n9552), .A2(n7162), .ZN(n9563) );
  INV_X1 U8543 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n7163) );
  XNOR2_X1 U8544 ( .A(n9558), .B(n7163), .ZN(n9564) );
  NAND2_X1 U8545 ( .A1(n9563), .A2(n9564), .ZN(n9562) );
  NAND2_X1 U8546 ( .A1(n9558), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n7164) );
  NAND2_X1 U8547 ( .A1(n9562), .A2(n7164), .ZN(n9580) );
  INV_X1 U8548 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n7165) );
  MUX2_X1 U8549 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n7165), .S(n9575), .Z(n9581)
         );
  NAND2_X1 U8550 ( .A1(n9580), .A2(n9581), .ZN(n9579) );
  NAND2_X1 U8551 ( .A1(n9575), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n7166) );
  NAND2_X1 U8552 ( .A1(n9579), .A2(n7166), .ZN(n9593) );
  INV_X1 U8553 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n7167) );
  MUX2_X1 U8554 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n7167), .S(n9588), .Z(n9594)
         );
  NAND2_X1 U8555 ( .A1(n9593), .A2(n9594), .ZN(n9592) );
  NAND2_X1 U8556 ( .A1(n9588), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n7168) );
  NAND2_X1 U8557 ( .A1(n9592), .A2(n7168), .ZN(n10280) );
  OR2_X1 U8558 ( .A1(n10291), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n7170) );
  NAND2_X1 U8559 ( .A1(P1_REG2_REG_7__SCAN_IN), .A2(n10291), .ZN(n7169) );
  AND2_X1 U8560 ( .A1(n7170), .A2(n7169), .ZN(n10281) );
  AND2_X1 U8561 ( .A1(n10280), .A2(n10281), .ZN(n10282) );
  AOI21_X1 U8562 ( .B1(n10291), .B2(P1_REG2_REG_7__SCAN_IN), .A(n10282), .ZN(
        n10297) );
  NAND2_X1 U8563 ( .A1(n10295), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n7171) );
  OAI21_X1 U8564 ( .B1(n10295), .B2(P1_REG2_REG_8__SCAN_IN), .A(n7171), .ZN(
        n10298) );
  NOR2_X1 U8565 ( .A1(n10297), .A2(n10298), .ZN(n10296) );
  AOI21_X1 U8566 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n10295), .A(n10296), .ZN(
        n7172) );
  NAND2_X1 U8567 ( .A1(n7173), .A2(n7172), .ZN(n7345) );
  OAI21_X1 U8568 ( .B1(n7173), .B2(n7172), .A(n7345), .ZN(n7197) );
  NAND2_X1 U8569 ( .A1(n7190), .A2(n7174), .ZN(n10338) );
  INV_X1 U8570 ( .A(n7354), .ZN(n7195) );
  INV_X1 U8571 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10654) );
  AOI22_X1 U8572 ( .A1(n7354), .A2(P1_REG1_REG_9__SCAN_IN), .B1(n10654), .B2(
        n7195), .ZN(n7189) );
  INV_X1 U8573 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10549) );
  MUX2_X1 U8574 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n10549), .S(n9535), .Z(n9538)
         );
  INV_X1 U8575 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10533) );
  MUX2_X1 U8576 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n10533), .S(n9515), .Z(n9521)
         );
  AND2_X1 U8577 ( .A1(P1_REG1_REG_0__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n9520) );
  NAND2_X1 U8578 ( .A1(n9521), .A2(n9520), .ZN(n9519) );
  NAND2_X1 U8579 ( .A1(n9515), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n7175) );
  NAND2_X1 U8580 ( .A1(n9519), .A2(n7175), .ZN(n9537) );
  NAND2_X1 U8581 ( .A1(n9538), .A2(n9537), .ZN(n9536) );
  NAND2_X1 U8582 ( .A1(n9535), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n7176) );
  NAND2_X1 U8583 ( .A1(n9536), .A2(n7176), .ZN(n9550) );
  INV_X1 U8584 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n7177) );
  XNOR2_X1 U8585 ( .A(n9548), .B(n7177), .ZN(n9551) );
  NAND2_X1 U8586 ( .A1(n9550), .A2(n9551), .ZN(n9549) );
  NAND2_X1 U8587 ( .A1(n9548), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n7178) );
  NAND2_X1 U8588 ( .A1(n9549), .A2(n7178), .ZN(n9566) );
  INV_X1 U8589 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n7179) );
  XNOR2_X1 U8590 ( .A(n9558), .B(n7179), .ZN(n9567) );
  NAND2_X1 U8591 ( .A1(n9566), .A2(n9567), .ZN(n9565) );
  NAND2_X1 U8592 ( .A1(n9558), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n7180) );
  NAND2_X1 U8593 ( .A1(n9565), .A2(n7180), .ZN(n9577) );
  INV_X1 U8594 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n7181) );
  MUX2_X1 U8595 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n7181), .S(n9575), .Z(n9578)
         );
  NAND2_X1 U8596 ( .A1(n9577), .A2(n9578), .ZN(n9576) );
  NAND2_X1 U8597 ( .A1(n9575), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n7182) );
  NAND2_X1 U8598 ( .A1(n9576), .A2(n7182), .ZN(n9590) );
  INV_X1 U8599 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n10616) );
  MUX2_X1 U8600 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n10616), .S(n9588), .Z(n9591)
         );
  NAND2_X1 U8601 ( .A1(n9590), .A2(n9591), .ZN(n9589) );
  NAND2_X1 U8602 ( .A1(n9588), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n7183) );
  NAND2_X1 U8603 ( .A1(n9589), .A2(n7183), .ZN(n10284) );
  OR2_X1 U8604 ( .A1(n10291), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n7185) );
  NAND2_X1 U8605 ( .A1(P1_REG1_REG_7__SCAN_IN), .A2(n10291), .ZN(n7184) );
  AND2_X1 U8606 ( .A1(n7185), .A2(n7184), .ZN(n10285) );
  AND2_X1 U8607 ( .A1(n10284), .A2(n10285), .ZN(n10286) );
  AND2_X1 U8608 ( .A1(n10291), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n7186) );
  NOR2_X1 U8609 ( .A1(n10286), .A2(n7186), .ZN(n10301) );
  INV_X1 U8610 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n7187) );
  MUX2_X1 U8611 ( .A(n7187), .B(P1_REG1_REG_8__SCAN_IN), .S(n10295), .Z(n10300) );
  NOR2_X1 U8612 ( .A1(n10301), .A2(n10300), .ZN(n10302) );
  AOI21_X1 U8613 ( .B1(P1_REG1_REG_8__SCAN_IN), .B2(n10295), .A(n10302), .ZN(
        n7188) );
  NAND2_X1 U8614 ( .A1(n7189), .A2(n7188), .ZN(n7353) );
  OAI21_X1 U8615 ( .B1(n7189), .B2(n7188), .A(n7353), .ZN(n7192) );
  INV_X1 U8616 ( .A(n7190), .ZN(n7191) );
  NOR2_X2 U8617 ( .A1(n7191), .A2(n8247), .ZN(n10334) );
  NAND2_X1 U8618 ( .A1(n7192), .A2(n10334), .ZN(n7194) );
  AND2_X1 U8619 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7858) );
  AOI21_X1 U8620 ( .B1(n9607), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n7858), .ZN(
        n7193) );
  OAI211_X1 U8621 ( .C1(n10338), .C2(n7195), .A(n7194), .B(n7193), .ZN(n7196)
         );
  AOI21_X1 U8622 ( .B1(n10329), .B2(n7197), .A(n7196), .ZN(n7198) );
  INV_X1 U8623 ( .A(n7198), .ZN(P1_U3252) );
  NAND2_X1 U8624 ( .A1(n9819), .A2(P1_U3973), .ZN(n7199) );
  OAI21_X1 U8625 ( .B1(n6002), .B2(P1_U3973), .A(n7199), .ZN(P1_U3571) );
  OAI222_X1 U8626 ( .A1(P2_U3151), .A2(n7202), .B1(n8052), .B2(n7201), .C1(
        n7200), .C2(n8237), .ZN(P2_U3286) );
  INV_X1 U8627 ( .A(n7203), .ZN(n7206) );
  AOI22_X1 U8628 ( .A1(n10389), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n10012), .ZN(n7204) );
  OAI21_X1 U8629 ( .B1(n7206), .B2(n7945), .A(n7204), .ZN(P1_U3345) );
  INV_X1 U8630 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n7205) );
  OAI222_X1 U8631 ( .A1(P2_U3151), .A2(n7207), .B1(n8052), .B2(n7206), .C1(
        n7205), .C2(n8237), .ZN(P2_U3285) );
  MUX2_X1 U8632 ( .A(n7208), .B(n8031), .S(P2_U3893), .Z(n7209) );
  INV_X1 U8633 ( .A(n7209), .ZN(P2_U3499) );
  MUX2_X1 U8634 ( .A(n7210), .B(n8042), .S(P2_U3893), .Z(n7211) );
  INV_X1 U8635 ( .A(n7211), .ZN(P2_U3500) );
  XOR2_X1 U8636 ( .A(n7213), .B(n7212), .Z(n9532) );
  INV_X1 U8637 ( .A(n9532), .ZN(n7218) );
  OR2_X1 U8638 ( .A1(n7214), .A2(P1_U3086), .ZN(n7241) );
  OAI22_X1 U8639 ( .A1(n9480), .A2(n10518), .B1(n7215), .B2(n9434), .ZN(n7216)
         );
  AOI21_X1 U8640 ( .B1(P1_REG3_REG_0__SCAN_IN), .B2(n7241), .A(n7216), .ZN(
        n7217) );
  OAI21_X1 U8641 ( .B1(n7218), .B2(n9496), .A(n7217), .ZN(P1_U3232) );
  INV_X1 U8642 ( .A(n7219), .ZN(n7222) );
  AOI22_X1 U8643 ( .A1(n8069), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n9345), .ZN(n7220) );
  OAI21_X1 U8644 ( .B1(n7222), .B2(n8052), .A(n7220), .ZN(P2_U3284) );
  AOI22_X1 U8645 ( .A1(n10320), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n10012), .ZN(n7221) );
  OAI21_X1 U8646 ( .B1(n7222), .B2(n7945), .A(n7221), .ZN(P1_U3344) );
  MUX2_X1 U8647 ( .A(n7223), .B(n10686), .S(P2_U3893), .Z(n7224) );
  INV_X1 U8648 ( .A(n7224), .ZN(P2_U3502) );
  INV_X1 U8649 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n7229) );
  INV_X1 U8650 ( .A(n7226), .ZN(n7227) );
  AOI22_X1 U8651 ( .A1(n7225), .A2(n7229), .B1(n7228), .B2(n7227), .ZN(
        P2_U3376) );
  XNOR2_X1 U8652 ( .A(n7231), .B(n7230), .ZN(n7233) );
  XNOR2_X1 U8653 ( .A(n7233), .B(n7232), .ZN(n7237) );
  NOR2_X1 U8654 ( .A1(n9480), .A2(n6373), .ZN(n7235) );
  OAI22_X1 U8655 ( .A1(n7513), .A2(n9434), .B1(n6895), .B2(n9491), .ZN(n7234)
         );
  AOI211_X1 U8656 ( .C1(P1_REG3_REG_1__SCAN_IN), .C2(n7241), .A(n7235), .B(
        n7234), .ZN(n7236) );
  OAI21_X1 U8657 ( .B1(n7237), .B2(n9496), .A(n7236), .ZN(P1_U3222) );
  OAI21_X1 U8658 ( .B1(n7240), .B2(n7239), .A(n7238), .ZN(n7245) );
  AOI22_X1 U8659 ( .A1(n9451), .A2(n10542), .B1(n9488), .B2(n10544), .ZN(n7243) );
  NAND2_X1 U8660 ( .A1(n7241), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n7242) );
  OAI211_X1 U8661 ( .C1(n10538), .C2(n9480), .A(n7243), .B(n7242), .ZN(n7244)
         );
  AOI21_X1 U8662 ( .B1(n7245), .B2(n9472), .A(n7244), .ZN(n7246) );
  INV_X1 U8663 ( .A(n7246), .ZN(P1_U3237) );
  AND2_X1 U8664 ( .A1(n7225), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  AND2_X1 U8665 ( .A1(n7225), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  AND2_X1 U8666 ( .A1(n7225), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U8667 ( .A1(n7225), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U8668 ( .A1(n7225), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  AND2_X1 U8669 ( .A1(n7225), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U8670 ( .A1(n7225), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3255) );
  AND2_X1 U8671 ( .A1(n7225), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U8672 ( .A1(n7225), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U8673 ( .A1(n7225), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U8674 ( .A1(n7225), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U8675 ( .A1(n7225), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U8676 ( .A1(n7225), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U8677 ( .A1(n7225), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  AND2_X1 U8678 ( .A1(n7225), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U8679 ( .A1(n7225), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U8680 ( .A1(n7225), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U8681 ( .A1(n7225), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U8682 ( .A1(n7225), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U8683 ( .A1(n7225), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  OAI21_X1 U8684 ( .B1(n7249), .B2(n7248), .A(n7247), .ZN(n7250) );
  NAND2_X1 U8685 ( .A1(n7250), .A2(n9472), .ZN(n7254) );
  NAND2_X1 U8686 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9545) );
  INV_X1 U8687 ( .A(n9545), .ZN(n7252) );
  OAI22_X1 U8688 ( .A1(n9480), .A2(n10571), .B1(n7513), .B2(n9491), .ZN(n7251)
         );
  AOI211_X1 U8689 ( .C1(n9488), .C2(n9511), .A(n7252), .B(n7251), .ZN(n7253)
         );
  OAI211_X1 U8690 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n9454), .A(n7254), .B(
        n7253), .ZN(P1_U3218) );
  INV_X1 U8691 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n7255) );
  MUX2_X1 U8692 ( .A(n7256), .B(n7255), .S(n8480), .Z(n7257) );
  NOR2_X1 U8693 ( .A1(n7257), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n7258) );
  OAI22_X1 U8694 ( .A1(n7259), .A2(n10495), .B1(n7274), .B2(n7258), .ZN(n7260)
         );
  OAI21_X1 U8695 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n10198), .A(n7260), .ZN(
        n7261) );
  AOI21_X1 U8696 ( .B1(n10498), .B2(P2_ADDR_REG_0__SCAN_IN), .A(n7261), .ZN(
        n7262) );
  OAI21_X1 U8697 ( .B1(n5265), .B2(n10507), .A(n7262), .ZN(P2_U3182) );
  INV_X1 U8698 ( .A(n7263), .ZN(n7266) );
  AOI22_X1 U8699 ( .A1(n8180), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_12__SCAN_IN), .B2(n9345), .ZN(n7264) );
  OAI21_X1 U8700 ( .B1(n7266), .B2(n8052), .A(n7264), .ZN(P2_U3283) );
  AOI22_X1 U8701 ( .A1(n8124), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n10012), .ZN(n7265) );
  OAI21_X1 U8702 ( .B1(n7266), .B2(n7945), .A(n7265), .ZN(P1_U3343) );
  INV_X1 U8703 ( .A(n7267), .ZN(n7313) );
  AOI22_X1 U8704 ( .A1(n10375), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n10003), .ZN(n7268) );
  OAI21_X1 U8705 ( .B1(n7313), .B2(n7945), .A(n7268), .ZN(P1_U3342) );
  INV_X1 U8706 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n7273) );
  AOI21_X1 U8707 ( .B1(n7271), .B2(n7270), .A(n7269), .ZN(n7272) );
  OAI22_X1 U8708 ( .A1(n10489), .A2(n7273), .B1(n10506), .B2(n7272), .ZN(n7284) );
  XOR2_X1 U8709 ( .A(n7275), .B(n7274), .Z(n7276) );
  NAND2_X1 U8710 ( .A1(n7276), .A2(n10495), .ZN(n7282) );
  INV_X1 U8711 ( .A(n7277), .ZN(n7279) );
  OAI21_X1 U8712 ( .B1(n7279), .B2(P2_REG1_REG_1__SCAN_IN), .A(n7278), .ZN(
        n7280) );
  NAND2_X1 U8713 ( .A1(n5649), .A2(n7280), .ZN(n7281) );
  OAI211_X1 U8714 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n7698), .A(n7282), .B(n7281), .ZN(n7283) );
  AOI211_X1 U8715 ( .C1(n10474), .C2(n7285), .A(n7284), .B(n7283), .ZN(n7286)
         );
  INV_X1 U8716 ( .A(n7286), .ZN(P2_U3183) );
  INV_X1 U8717 ( .A(n10495), .ZN(n7872) );
  XNOR2_X1 U8718 ( .A(n7288), .B(n7287), .ZN(n7304) );
  NOR2_X1 U8719 ( .A1(n10507), .A2(n4925), .ZN(n7302) );
  NOR2_X1 U8720 ( .A1(n7291), .A2(n7290), .ZN(n7292) );
  OAI21_X1 U8721 ( .B1(n7293), .B2(n7292), .A(n5686), .ZN(n7299) );
  NOR2_X1 U8722 ( .A1(n7295), .A2(n7294), .ZN(n7296) );
  OAI21_X1 U8723 ( .B1(n7297), .B2(n7296), .A(n5649), .ZN(n7298) );
  OAI211_X1 U8724 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n7300), .A(n7299), .B(n7298), .ZN(n7301) );
  AOI211_X1 U8725 ( .C1(n10498), .C2(P2_ADDR_REG_2__SCAN_IN), .A(n7302), .B(
        n7301), .ZN(n7303) );
  OAI21_X1 U8726 ( .B1(n7872), .B2(n7304), .A(n7303), .ZN(P2_U3184) );
  INV_X1 U8727 ( .A(n7546), .ZN(n7311) );
  AOI21_X1 U8728 ( .B1(n7305), .B2(n6931), .A(n9496), .ZN(n7307) );
  NAND2_X1 U8729 ( .A1(n7307), .A2(n7306), .ZN(n7310) );
  AND2_X1 U8730 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n9561) );
  OAI22_X1 U8731 ( .A1(n9480), .A2(n10593), .B1(n7575), .B2(n9434), .ZN(n7308)
         );
  AOI211_X1 U8732 ( .C1(n9451), .C2(n10544), .A(n9561), .B(n7308), .ZN(n7309)
         );
  OAI211_X1 U8733 ( .C1(n9454), .C2(n7311), .A(n7310), .B(n7309), .ZN(P1_U3230) );
  INV_X1 U8734 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n7312) );
  OAI222_X1 U8735 ( .A1(n7314), .A2(P2_U3151), .B1(n8052), .B2(n7313), .C1(
        n7312), .C2(n8237), .ZN(P2_U3282) );
  NAND2_X1 U8736 ( .A1(n9707), .A2(P1_U3973), .ZN(n7315) );
  OAI21_X1 U8737 ( .B1(P1_U3973), .B2(n8223), .A(n7315), .ZN(P1_U3578) );
  INV_X1 U8738 ( .A(n7316), .ZN(n7336) );
  AOI22_X1 U8739 ( .A1(n10324), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n10003), .ZN(n7317) );
  OAI21_X1 U8740 ( .B1(n7336), .B2(n7945), .A(n7317), .ZN(P1_U3341) );
  AOI21_X1 U8741 ( .B1(n7319), .B2(n10581), .A(n7318), .ZN(n7320) );
  NOR2_X1 U8742 ( .A1(n10501), .A2(n7320), .ZN(n7332) );
  INV_X1 U8743 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n7325) );
  AOI21_X1 U8744 ( .B1(n7323), .B2(n7322), .A(n7321), .ZN(n7324) );
  OAI22_X1 U8745 ( .A1(n10489), .A2(n7325), .B1(n7324), .B2(n7872), .ZN(n7331)
         );
  AOI21_X1 U8746 ( .B1(n7328), .B2(n7327), .A(n7326), .ZN(n7329) );
  NOR2_X1 U8747 ( .A1(n10506), .A2(n7329), .ZN(n7330) );
  INV_X1 U8748 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n10080) );
  NOR2_X1 U8749 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10080), .ZN(n7616) );
  NOR4_X1 U8750 ( .A1(n7332), .A2(n7331), .A3(n7330), .A4(n7616), .ZN(n7333)
         );
  OAI21_X1 U8751 ( .B1(n7334), .B2(n10507), .A(n7333), .ZN(P2_U3185) );
  OAI222_X1 U8752 ( .A1(n7337), .A2(P2_U3151), .B1(n8052), .B2(n7336), .C1(
        n7335), .C2(n8237), .ZN(P2_U3281) );
  NAND2_X1 U8753 ( .A1(n6249), .A2(n7499), .ZN(n8261) );
  NAND2_X1 U8754 ( .A1(n8255), .A2(n8261), .ZN(n8445) );
  INV_X1 U8755 ( .A(n8445), .ZN(n7339) );
  NOR2_X1 U8756 ( .A1(n10749), .A2(n9211), .ZN(n7338) );
  OAI222_X1 U8757 ( .A1(n7499), .A2(n10740), .B1(n7339), .B2(n7338), .C1(
        n10754), .C2(n7628), .ZN(n7341) );
  NAND2_X1 U8758 ( .A1(n7341), .A2(n10761), .ZN(n7340) );
  OAI21_X1 U8759 ( .B1(n10761), .B2(n7255), .A(n7340), .ZN(P2_U3459) );
  INV_X1 U8760 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n7343) );
  NAND2_X1 U8761 ( .A1(n7341), .A2(n10764), .ZN(n7342) );
  OAI21_X1 U8762 ( .B1(n10764), .B2(n7343), .A(n7342), .ZN(P2_U3390) );
  NOR2_X1 U8763 ( .A1(n8124), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n7344) );
  AOI21_X1 U8764 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n8124), .A(n7344), .ZN(
        n7349) );
  OAI21_X1 U8765 ( .B1(n7354), .B2(P1_REG2_REG_9__SCAN_IN), .A(n7345), .ZN(
        n10386) );
  NAND2_X1 U8766 ( .A1(P1_REG2_REG_10__SCAN_IN), .A2(n10389), .ZN(n7346) );
  OAI21_X1 U8767 ( .B1(P1_REG2_REG_10__SCAN_IN), .B2(n10389), .A(n7346), .ZN(
        n10385) );
  NOR2_X1 U8768 ( .A1(n10386), .A2(n10385), .ZN(n10384) );
  AOI21_X1 U8769 ( .B1(n10389), .B2(P1_REG2_REG_10__SCAN_IN), .A(n10384), .ZN(
        n10314) );
  NAND2_X1 U8770 ( .A1(n10320), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n7347) );
  OAI21_X1 U8771 ( .B1(n10320), .B2(P1_REG2_REG_11__SCAN_IN), .A(n7347), .ZN(
        n10313) );
  NOR2_X1 U8772 ( .A1(n10314), .A2(n10313), .ZN(n10312) );
  AOI21_X1 U8773 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n10320), .A(n10312), .ZN(
        n7348) );
  NAND2_X1 U8774 ( .A1(n7349), .A2(n7348), .ZN(n8123) );
  OAI21_X1 U8775 ( .B1(n7349), .B2(n7348), .A(n8123), .ZN(n7350) );
  INV_X1 U8776 ( .A(n7350), .ZN(n7364) );
  INV_X1 U8777 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n7351) );
  INV_X1 U8778 ( .A(n8124), .ZN(n7360) );
  AOI22_X1 U8779 ( .A1(n8124), .A2(P1_REG1_REG_12__SCAN_IN), .B1(n7351), .B2(
        n7360), .ZN(n7357) );
  INV_X1 U8780 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n7352) );
  MUX2_X1 U8781 ( .A(n7352), .B(P1_REG1_REG_10__SCAN_IN), .S(n10389), .Z(
        n10381) );
  OAI21_X1 U8782 ( .B1(n7354), .B2(P1_REG1_REG_9__SCAN_IN), .A(n7353), .ZN(
        n10382) );
  NOR2_X1 U8783 ( .A1(n10381), .A2(n10382), .ZN(n10380) );
  AOI21_X1 U8784 ( .B1(n10389), .B2(P1_REG1_REG_10__SCAN_IN), .A(n10380), .ZN(
        n10317) );
  INV_X1 U8785 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n7355) );
  MUX2_X1 U8786 ( .A(n7355), .B(P1_REG1_REG_11__SCAN_IN), .S(n10320), .Z(
        n10316) );
  NOR2_X1 U8787 ( .A1(n10317), .A2(n10316), .ZN(n10315) );
  AOI21_X1 U8788 ( .B1(P1_REG1_REG_11__SCAN_IN), .B2(n10320), .A(n10315), .ZN(
        n7356) );
  NAND2_X1 U8789 ( .A1(n7357), .A2(n7356), .ZN(n8115) );
  OAI21_X1 U8790 ( .B1(n7357), .B2(n7356), .A(n8115), .ZN(n7362) );
  NOR2_X1 U8791 ( .A1(n7358), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8200) );
  AOI21_X1 U8792 ( .B1(n9607), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n8200), .ZN(
        n7359) );
  OAI21_X1 U8793 ( .B1(n10338), .B2(n7360), .A(n7359), .ZN(n7361) );
  AOI21_X1 U8794 ( .B1(n7362), .B2(n10334), .A(n7361), .ZN(n7363) );
  OAI21_X1 U8795 ( .B1(n7364), .B2(n10383), .A(n7363), .ZN(P1_U3255) );
  INV_X1 U8796 ( .A(n7588), .ZN(n7642) );
  XNOR2_X1 U8797 ( .A(n6741), .B(n7365), .ZN(n10532) );
  AOI211_X1 U8798 ( .C1(n8606), .C2(n7366), .A(n9797), .B(n5025), .ZN(n10528)
         );
  AOI22_X1 U8799 ( .A1(n10528), .A2(n4924), .B1(P1_REG3_REG_1__SCAN_IN), .B2(
        n10554), .ZN(n7367) );
  OAI21_X1 U8800 ( .B1(n6373), .B2(n9802), .A(n7367), .ZN(n7375) );
  OAI21_X1 U8801 ( .B1(n7369), .B2(n8607), .A(n7368), .ZN(n7370) );
  NAND2_X1 U8802 ( .A1(n7370), .A2(n10546), .ZN(n7373) );
  NAND2_X1 U8803 ( .A1(n10532), .A2(n7635), .ZN(n7372) );
  INV_X1 U8804 ( .A(n6895), .ZN(n9513) );
  AOI22_X1 U8805 ( .A1(n9513), .A2(n10541), .B1(n10543), .B2(n9512), .ZN(n7371) );
  NAND3_X1 U8806 ( .A1(n7373), .A2(n7372), .A3(n7371), .ZN(n10531) );
  MUX2_X1 U8807 ( .A(n10531), .B(P1_REG2_REG_1__SCAN_IN), .S(n10555), .Z(n7374) );
  AOI211_X1 U8808 ( .C1(n7642), .C2(n10532), .A(n7375), .B(n7374), .ZN(n7376)
         );
  INV_X1 U8809 ( .A(n7376), .ZN(P1_U3292) );
  INV_X2 U8810 ( .A(P1_U3973), .ZN(n9528) );
  NAND2_X1 U8811 ( .A1(n9528), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n7377) );
  OAI21_X1 U8812 ( .B1(n8753), .B2(n9528), .A(n7377), .ZN(P1_U3583) );
  NAND2_X1 U8813 ( .A1(n5429), .A2(n7378), .ZN(n7380) );
  XNOR2_X1 U8814 ( .A(n7380), .B(n7379), .ZN(n7386) );
  NAND2_X1 U8815 ( .A1(n9486), .A2(n7397), .ZN(n7383) );
  NAND2_X1 U8816 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n9572) );
  INV_X1 U8817 ( .A(n9572), .ZN(n7381) );
  AOI21_X1 U8818 ( .B1(n9488), .B2(n9509), .A(n7381), .ZN(n7382) );
  OAI211_X1 U8819 ( .C1(n7512), .C2(n9491), .A(n7383), .B(n7382), .ZN(n7384)
         );
  AOI21_X1 U8820 ( .B1(n7491), .B2(n9494), .A(n7384), .ZN(n7385) );
  OAI21_X1 U8821 ( .B1(n7386), .B2(n9496), .A(n7385), .ZN(P1_U3227) );
  AOI21_X1 U8822 ( .B1(n8255), .B2(n6248), .A(n7767), .ZN(n7702) );
  OAI22_X1 U8823 ( .A1(n7702), .A2(n10710), .B1(n7614), .B2(n10754), .ZN(n7390) );
  INV_X1 U8824 ( .A(n7387), .ZN(n7415) );
  XNOR2_X1 U8825 ( .A(n6248), .B(n7415), .ZN(n7389) );
  INV_X1 U8826 ( .A(n6249), .ZN(n7388) );
  OAI22_X1 U8827 ( .A1(n7389), .A2(n9234), .B1(n7388), .B2(n9236), .ZN(n7696)
         );
  NOR2_X1 U8828 ( .A1(n7390), .A2(n7696), .ZN(n7592) );
  INV_X1 U8829 ( .A(n9288), .ZN(n9293) );
  AOI22_X1 U8830 ( .A1(n9293), .A2(n5755), .B1(n10760), .B2(
        P2_REG1_REG_1__SCAN_IN), .ZN(n7391) );
  OAI21_X1 U8831 ( .B1(n7592), .B2(n10760), .A(n7391), .ZN(P2_U3460) );
  XOR2_X1 U8832 ( .A(n8610), .B(n7392), .Z(n7486) );
  OAI21_X1 U8833 ( .B1(n8610), .B2(n7394), .A(n7393), .ZN(n7395) );
  AOI222_X1 U8834 ( .A1(n10546), .A2(n7395), .B1(n9509), .B2(n10543), .C1(
        n9511), .C2(n10541), .ZN(n7487) );
  MUX2_X1 U8835 ( .A(n7165), .B(n7487), .S(n10524), .Z(n7401) );
  INV_X1 U8836 ( .A(n7581), .ZN(n7396) );
  AOI211_X1 U8837 ( .C1(n7491), .C2(n7544), .A(n9797), .B(n7396), .ZN(n7489)
         );
  INV_X1 U8838 ( .A(n7397), .ZN(n7398) );
  OAI22_X1 U8839 ( .A1(n9802), .A2(n7494), .B1(n9854), .B2(n7398), .ZN(n7399)
         );
  AOI21_X1 U8840 ( .B1(n7489), .B2(n4924), .A(n7399), .ZN(n7400) );
  OAI211_X1 U8841 ( .C1(n9836), .C2(n7486), .A(n7401), .B(n7400), .ZN(P1_U3288) );
  INV_X1 U8842 ( .A(n7402), .ZN(n7405) );
  AOI22_X1 U8843 ( .A1(n8994), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_15__SCAN_IN), .B2(n9345), .ZN(n7403) );
  OAI21_X1 U8844 ( .B1(n7405), .B2(n8052), .A(n7403), .ZN(P2_U3280) );
  AOI22_X1 U8845 ( .A1(n10350), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n10003), .ZN(n7404) );
  OAI21_X1 U8846 ( .B1(n7405), .B2(n7945), .A(n7404), .ZN(P1_U3340) );
  INV_X1 U8847 ( .A(n7406), .ZN(n7408) );
  NAND2_X1 U8848 ( .A1(n7408), .A2(n7407), .ZN(n7412) );
  INV_X1 U8849 ( .A(n7409), .ZN(n7410) );
  OR2_X1 U8850 ( .A1(n8254), .A2(n7410), .ZN(n7411) );
  NAND2_X2 U8851 ( .A1(n7412), .A2(n7411), .ZN(n7417) );
  INV_X2 U8852 ( .A(n7417), .ZN(n7984) );
  XNOR2_X1 U8853 ( .A(n7924), .B(n7413), .ZN(n7502) );
  XNOR2_X1 U8854 ( .A(n7502), .B(n8939), .ZN(n7422) );
  XNOR2_X1 U8855 ( .A(n7924), .B(n10577), .ZN(n7420) );
  XNOR2_X1 U8856 ( .A(n7417), .B(n7414), .ZN(n7416) );
  NAND2_X1 U8857 ( .A1(n7527), .A2(n7528), .ZN(n7526) );
  OAI21_X1 U8858 ( .B1(n7416), .B2(n8942), .A(n7526), .ZN(n7479) );
  XNOR2_X1 U8859 ( .A(n7417), .B(n7481), .ZN(n7418) );
  XNOR2_X1 U8860 ( .A(n7418), .B(n8941), .ZN(n7480) );
  AOI21_X1 U8861 ( .B1(n7479), .B2(n7480), .A(n7419), .ZN(n7613) );
  XNOR2_X1 U8862 ( .A(n7420), .B(n7438), .ZN(n7612) );
  AOI21_X1 U8863 ( .B1(n7422), .B2(n7421), .A(n7504), .ZN(n7457) );
  INV_X1 U8864 ( .A(n7423), .ZN(n7424) );
  NAND2_X1 U8865 ( .A1(n7442), .A2(n7424), .ZN(n7427) );
  INV_X1 U8866 ( .A(n7448), .ZN(n7425) );
  NAND2_X1 U8867 ( .A1(n7450), .A2(n7425), .ZN(n7426) );
  NAND2_X1 U8868 ( .A1(n7427), .A2(n7426), .ZN(n7429) );
  NAND2_X1 U8869 ( .A1(n7442), .A2(n7430), .ZN(n7431) );
  INV_X1 U8870 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n10193) );
  NOR2_X1 U8871 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10193), .ZN(n10402) );
  NOR2_X1 U8872 ( .A1(n7433), .A2(n7432), .ZN(n8482) );
  AND2_X1 U8873 ( .A1(n7450), .A2(n8482), .ZN(n7434) );
  INV_X1 U8874 ( .A(n8938), .ZN(n7437) );
  INV_X1 U8875 ( .A(n7434), .ZN(n7436) );
  OAI22_X1 U8876 ( .A1(n8897), .A2(n7438), .B1(n7437), .B2(n8918), .ZN(n7439)
         );
  AOI211_X1 U8877 ( .C1(n10585), .C2(n8910), .A(n10402), .B(n7439), .ZN(n7456)
         );
  INV_X1 U8878 ( .A(n7440), .ZN(n7441) );
  OR2_X1 U8879 ( .A1(n7442), .A2(n7441), .ZN(n7447) );
  AND3_X1 U8880 ( .A1(n7445), .A2(n7444), .A3(n7443), .ZN(n7446) );
  OAI211_X1 U8881 ( .C1(n7450), .C2(n7448), .A(n7447), .B(n7446), .ZN(n7449)
         );
  NAND2_X1 U8882 ( .A1(n7449), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7453) );
  INV_X1 U8883 ( .A(n8482), .ZN(n7451) );
  OR2_X1 U8884 ( .A1(n7451), .A2(n7450), .ZN(n7452) );
  INV_X1 U8885 ( .A(n8919), .ZN(n8899) );
  INV_X1 U8886 ( .A(n7454), .ZN(n7780) );
  NAND2_X1 U8887 ( .A1(n8899), .A2(n7780), .ZN(n7455) );
  OAI211_X1 U8888 ( .C1(n7457), .C2(n8912), .A(n7456), .B(n7455), .ZN(P2_U3170) );
  NAND2_X1 U8889 ( .A1(n9090), .A2(P2_U3893), .ZN(n7458) );
  OAI21_X1 U8890 ( .B1(P2_U3893), .B2(n6161), .A(n7458), .ZN(P2_U3516) );
  NAND2_X1 U8891 ( .A1(n7460), .A2(n7459), .ZN(n7462) );
  XOR2_X1 U8892 ( .A(n7462), .B(n7461), .Z(n7468) );
  NAND2_X1 U8893 ( .A1(n9486), .A2(n7582), .ZN(n7465) );
  NAND2_X1 U8894 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9585) );
  INV_X1 U8895 ( .A(n9585), .ZN(n7463) );
  AOI21_X1 U8896 ( .B1(n9488), .B2(n9508), .A(n7463), .ZN(n7464) );
  OAI211_X1 U8897 ( .C1(n7575), .C2(n9491), .A(n7465), .B(n7464), .ZN(n7466)
         );
  AOI21_X1 U8898 ( .B1(n10609), .B2(n9494), .A(n7466), .ZN(n7467) );
  OAI21_X1 U8899 ( .B1(n7468), .B2(n9496), .A(n7467), .ZN(P1_U3239) );
  XNOR2_X1 U8900 ( .A(n7471), .B(n7470), .ZN(n7472) );
  XNOR2_X1 U8901 ( .A(n7469), .B(n7472), .ZN(n7478) );
  NAND2_X1 U8902 ( .A1(n9486), .A2(n7685), .ZN(n7475) );
  NAND2_X1 U8903 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n10292) );
  INV_X1 U8904 ( .A(n10292), .ZN(n7473) );
  AOI21_X1 U8905 ( .B1(n9488), .B2(n9507), .A(n7473), .ZN(n7474) );
  OAI211_X1 U8906 ( .C1(n7677), .C2(n9491), .A(n7475), .B(n7474), .ZN(n7476)
         );
  AOI21_X1 U8907 ( .B1(n7684), .B2(n9494), .A(n7476), .ZN(n7477) );
  OAI21_X1 U8908 ( .B1(n7478), .B2(n9496), .A(n7477), .ZN(P1_U3213) );
  XOR2_X1 U8909 ( .A(n7480), .B(n7479), .Z(n7485) );
  NAND2_X1 U8910 ( .A1(n8919), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7498) );
  AOI22_X1 U8911 ( .A1(n8895), .A2(n8940), .B1(n8910), .B2(n7481), .ZN(n7482)
         );
  OAI21_X1 U8912 ( .B1(n7628), .B2(n8897), .A(n7482), .ZN(n7483) );
  AOI21_X1 U8913 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(n7498), .A(n7483), .ZN(
        n7484) );
  OAI21_X1 U8914 ( .B1(n7485), .B2(n8912), .A(n7484), .ZN(P2_U3177) );
  INV_X1 U8915 ( .A(n7486), .ZN(n7490) );
  INV_X1 U8916 ( .A(n7487), .ZN(n7488) );
  AOI211_X1 U8917 ( .C1(n7490), .C2(n10675), .A(n7489), .B(n7488), .ZN(n7497)
         );
  INV_X1 U8918 ( .A(n9934), .ZN(n9940) );
  AOI22_X1 U8919 ( .A1(n9940), .A2(n7491), .B1(n10676), .B2(
        P1_REG1_REG_5__SCAN_IN), .ZN(n7492) );
  OAI21_X1 U8920 ( .B1(n7497), .B2(n10676), .A(n7492), .ZN(P1_U3527) );
  INV_X1 U8921 ( .A(n10681), .ZN(n10678) );
  INV_X1 U8922 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n7493) );
  OAI22_X1 U8923 ( .A1(n9995), .A2(n7494), .B1(n10681), .B2(n7493), .ZN(n7495)
         );
  INV_X1 U8924 ( .A(n7495), .ZN(n7496) );
  OAI21_X1 U8925 ( .B1(n7497), .B2(n10678), .A(n7496), .ZN(P1_U3468) );
  INV_X1 U8926 ( .A(n7498), .ZN(n7533) );
  INV_X1 U8927 ( .A(n8910), .ZN(n8925) );
  OAI22_X1 U8928 ( .A1(n8925), .A2(n7499), .B1(n7628), .B2(n8918), .ZN(n7500)
         );
  AOI21_X1 U8929 ( .B1(n8914), .B2(n8445), .A(n7500), .ZN(n7501) );
  OAI21_X1 U8930 ( .B1(n7533), .B2(n10198), .A(n7501), .ZN(P2_U3172) );
  INV_X1 U8931 ( .A(n8939), .ZN(n8002) );
  INV_X1 U8932 ( .A(n7502), .ZN(n7503) );
  XNOR2_X1 U8933 ( .A(n10600), .B(n8796), .ZN(n7716) );
  XNOR2_X1 U8934 ( .A(n7716), .B(n8938), .ZN(n7717) );
  XOR2_X1 U8935 ( .A(n7718), .B(n7717), .Z(n7509) );
  NOR2_X1 U8936 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5816), .ZN(n10417) );
  AOI21_X1 U8937 ( .B1(n8895), .B2(n8937), .A(n10417), .ZN(n7506) );
  NAND2_X1 U8938 ( .A1(n8922), .A2(n8939), .ZN(n7505) );
  OAI211_X1 U8939 ( .C1(n8919), .C2(n8004), .A(n7506), .B(n7505), .ZN(n7507)
         );
  AOI21_X1 U8940 ( .B1(n8007), .B2(n8910), .A(n7507), .ZN(n7508) );
  OAI21_X1 U8941 ( .B1(n7509), .B2(n8912), .A(n7508), .ZN(P2_U3167) );
  NAND2_X1 U8942 ( .A1(n10508), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n7510) );
  OAI21_X1 U8943 ( .B1(n9040), .B2(n10508), .A(n7510), .ZN(P2_U3520) );
  XNOR2_X1 U8944 ( .A(n7511), .B(n8608), .ZN(n10569) );
  OAI21_X1 U8945 ( .B1(n8608), .B2(n8497), .A(n7538), .ZN(n7515) );
  INV_X1 U8946 ( .A(n9821), .ZN(n9762) );
  OAI22_X1 U8947 ( .A1(n7513), .A2(n9762), .B1(n7512), .B2(n9764), .ZN(n7514)
         );
  AOI21_X1 U8948 ( .B1(n7515), .B2(n10546), .A(n7514), .ZN(n7516) );
  OAI21_X1 U8949 ( .B1(n10569), .B2(n7517), .A(n7516), .ZN(n10572) );
  NAND2_X1 U8950 ( .A1(n10572), .A2(n10524), .ZN(n7525) );
  OAI22_X1 U8951 ( .A1(n10524), .A2(n7518), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n9854), .ZN(n7522) );
  INV_X1 U8952 ( .A(n10536), .ZN(n7520) );
  INV_X1 U8953 ( .A(n7545), .ZN(n7519) );
  OAI211_X1 U8954 ( .C1(n10571), .C2(n7520), .A(n7519), .B(n10537), .ZN(n10570) );
  INV_X1 U8955 ( .A(n4924), .ZN(n9832) );
  NOR2_X1 U8956 ( .A1(n10570), .A2(n9832), .ZN(n7521) );
  AOI211_X1 U8957 ( .C1(n10552), .C2(n7523), .A(n7522), .B(n7521), .ZN(n7524)
         );
  OAI211_X1 U8958 ( .C1(n10569), .C2(n7588), .A(n7525), .B(n7524), .ZN(
        P1_U3290) );
  OAI21_X1 U8959 ( .B1(n7528), .B2(n7527), .A(n7526), .ZN(n7529) );
  NAND2_X1 U8960 ( .A1(n7529), .A2(n8914), .ZN(n7532) );
  OAI22_X1 U8961 ( .A1(n8925), .A2(n7414), .B1(n7614), .B2(n8918), .ZN(n7530)
         );
  AOI21_X1 U8962 ( .B1(n8922), .B2(n6249), .A(n7530), .ZN(n7531) );
  OAI211_X1 U8963 ( .C1(n7533), .C2(n7698), .A(n7532), .B(n7531), .ZN(P2_U3162) );
  INV_X1 U8964 ( .A(n7534), .ZN(n7609) );
  AOI22_X1 U8965 ( .A1(n8214), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n10003), .ZN(n7535) );
  OAI21_X1 U8966 ( .B1(n7609), .B2(n7945), .A(n7535), .ZN(P1_U3339) );
  XOR2_X1 U8967 ( .A(n7536), .B(n8609), .Z(n10596) );
  INV_X1 U8968 ( .A(n10596), .ZN(n7552) );
  INV_X1 U8969 ( .A(n8609), .ZN(n7537) );
  NAND3_X1 U8970 ( .A1(n7538), .A2(n7537), .A3(n8495), .ZN(n7539) );
  NAND2_X1 U8971 ( .A1(n7540), .A2(n7539), .ZN(n7541) );
  NAND2_X1 U8972 ( .A1(n7541), .A2(n10546), .ZN(n7543) );
  AOI22_X1 U8973 ( .A1(n10541), .A2(n10544), .B1(n9510), .B2(n10543), .ZN(
        n7542) );
  NAND2_X1 U8974 ( .A1(n7543), .A2(n7542), .ZN(n10594) );
  OAI211_X1 U8975 ( .C1(n7545), .C2(n10593), .A(n7544), .B(n10537), .ZN(n10592) );
  AOI22_X1 U8976 ( .A1(n10555), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n7546), .B2(
        n10554), .ZN(n7549) );
  NAND2_X1 U8977 ( .A1(n10552), .A2(n7547), .ZN(n7548) );
  OAI211_X1 U8978 ( .C1(n10592), .C2(n9832), .A(n7549), .B(n7548), .ZN(n7550)
         );
  AOI21_X1 U8979 ( .B1(n10594), .B2(n10524), .A(n7550), .ZN(n7551) );
  OAI21_X1 U8980 ( .B1(n7552), .B2(n9836), .A(n7551), .ZN(P1_U3289) );
  NOR2_X1 U8981 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(P1_ADDR_REG_18__SCAN_IN), 
        .ZN(n7553) );
  AOI21_X1 U8982 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(P2_ADDR_REG_18__SCAN_IN), 
        .A(n7553), .ZN(n10276) );
  NOR2_X1 U8983 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7554) );
  AOI21_X1 U8984 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n7554), .ZN(n10273) );
  NOR2_X1 U8985 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7555) );
  AOI21_X1 U8986 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n7555), .ZN(n10270) );
  NOR2_X1 U8987 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7556) );
  AOI21_X1 U8988 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n7556), .ZN(n10267) );
  NOR2_X1 U8989 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7557) );
  AOI21_X1 U8990 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n7557), .ZN(n10264) );
  NOR2_X1 U8991 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7558) );
  AOI21_X1 U8992 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n7558), .ZN(n10261) );
  NOR2_X1 U8993 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7559) );
  AOI21_X1 U8994 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n7559), .ZN(n10258) );
  NOR2_X1 U8995 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n7560) );
  AOI21_X1 U8996 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n7560), .ZN(n10255) );
  NOR2_X1 U8997 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n7561) );
  AOI21_X1 U8998 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n7561), .ZN(n10252) );
  NOR2_X1 U8999 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n7562) );
  AOI21_X1 U9000 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(P2_ADDR_REG_9__SCAN_IN), 
        .A(n7562), .ZN(n10249) );
  NOR2_X1 U9001 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n7563) );
  AOI21_X1 U9002 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(P2_ADDR_REG_8__SCAN_IN), 
        .A(n7563), .ZN(n10246) );
  NOR2_X1 U9003 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n7564) );
  AOI21_X1 U9004 ( .B1(P1_ADDR_REG_7__SCAN_IN), .B2(P2_ADDR_REG_7__SCAN_IN), 
        .A(n7564), .ZN(n10243) );
  NOR2_X1 U9005 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n7565) );
  AOI21_X1 U9006 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(P2_ADDR_REG_6__SCAN_IN), 
        .A(n7565), .ZN(n10240) );
  NOR2_X1 U9007 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n7566) );
  AOI21_X1 U9008 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(P2_ADDR_REG_5__SCAN_IN), 
        .A(n7566), .ZN(n10237) );
  NAND2_X1 U9009 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .ZN(n10223) );
  INV_X1 U9010 ( .A(n10223), .ZN(n7567) );
  INV_X1 U9011 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10224) );
  NAND2_X1 U9012 ( .A1(n10224), .A2(n10223), .ZN(n10222) );
  AOI22_X1 U9013 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n7567), .B1(
        P2_ADDR_REG_1__SCAN_IN), .B2(n10222), .ZN(n10228) );
  NAND2_X1 U9014 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n7568) );
  OAI21_X1 U9015 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(P2_ADDR_REG_2__SCAN_IN), 
        .A(n7568), .ZN(n10227) );
  NOR2_X1 U9016 ( .A1(n10228), .A2(n10227), .ZN(n10226) );
  AOI21_X1 U9017 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(P1_ADDR_REG_2__SCAN_IN), 
        .A(n10226), .ZN(n10231) );
  NAND2_X1 U9018 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(P1_ADDR_REG_3__SCAN_IN), 
        .ZN(n7569) );
  OAI21_X1 U9019 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(P1_ADDR_REG_3__SCAN_IN), 
        .A(n7569), .ZN(n10230) );
  NOR2_X1 U9020 ( .A1(n10231), .A2(n10230), .ZN(n10229) );
  AOI21_X1 U9021 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(P2_ADDR_REG_3__SCAN_IN), 
        .A(n10229), .ZN(n10234) );
  NOR2_X1 U9022 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7570) );
  AOI21_X1 U9023 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(P1_ADDR_REG_4__SCAN_IN), 
        .A(n7570), .ZN(n10233) );
  NAND2_X1 U9024 ( .A1(n10234), .A2(n10233), .ZN(n10232) );
  OAI21_X1 U9025 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(P2_ADDR_REG_4__SCAN_IN), 
        .A(n10232), .ZN(n10236) );
  NAND2_X1 U9026 ( .A1(n10237), .A2(n10236), .ZN(n10235) );
  OAI21_X1 U9027 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(P1_ADDR_REG_5__SCAN_IN), 
        .A(n10235), .ZN(n10239) );
  NAND2_X1 U9028 ( .A1(n10240), .A2(n10239), .ZN(n10238) );
  OAI21_X1 U9029 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(P1_ADDR_REG_6__SCAN_IN), 
        .A(n10238), .ZN(n10242) );
  NAND2_X1 U9030 ( .A1(n10243), .A2(n10242), .ZN(n10241) );
  OAI21_X1 U9031 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(P1_ADDR_REG_7__SCAN_IN), 
        .A(n10241), .ZN(n10245) );
  NAND2_X1 U9032 ( .A1(n10246), .A2(n10245), .ZN(n10244) );
  OAI21_X1 U9033 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(P1_ADDR_REG_8__SCAN_IN), 
        .A(n10244), .ZN(n10248) );
  NAND2_X1 U9034 ( .A1(n10249), .A2(n10248), .ZN(n10247) );
  OAI21_X1 U9035 ( .B1(P2_ADDR_REG_9__SCAN_IN), .B2(P1_ADDR_REG_9__SCAN_IN), 
        .A(n10247), .ZN(n10251) );
  NAND2_X1 U9036 ( .A1(n10252), .A2(n10251), .ZN(n10250) );
  OAI21_X1 U9037 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10250), .ZN(n10254) );
  NAND2_X1 U9038 ( .A1(n10255), .A2(n10254), .ZN(n10253) );
  OAI21_X1 U9039 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10253), .ZN(n10257) );
  NAND2_X1 U9040 ( .A1(n10258), .A2(n10257), .ZN(n10256) );
  OAI21_X1 U9041 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10256), .ZN(n10260) );
  NAND2_X1 U9042 ( .A1(n10261), .A2(n10260), .ZN(n10259) );
  OAI21_X1 U9043 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10259), .ZN(n10263) );
  NAND2_X1 U9044 ( .A1(n10264), .A2(n10263), .ZN(n10262) );
  OAI21_X1 U9045 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10262), .ZN(n10266) );
  NAND2_X1 U9046 ( .A1(n10267), .A2(n10266), .ZN(n10265) );
  OAI21_X1 U9047 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10265), .ZN(n10269) );
  NAND2_X1 U9048 ( .A1(n10270), .A2(n10269), .ZN(n10268) );
  OAI21_X1 U9049 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10268), .ZN(n10272) );
  NAND2_X1 U9050 ( .A1(n10273), .A2(n10272), .ZN(n10271) );
  OAI21_X1 U9051 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10271), .ZN(n10275) );
  NAND2_X1 U9052 ( .A1(n10276), .A2(n10275), .ZN(n10274) );
  OAI21_X1 U9053 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(P1_ADDR_REG_18__SCAN_IN), 
        .A(n10274), .ZN(n7572) );
  XNOR2_X1 U9054 ( .A(n5382), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n7571) );
  XNOR2_X1 U9055 ( .A(n7572), .B(n7571), .ZN(ADD_1068_U4) );
  OAI21_X1 U9056 ( .B1(n7574), .B2(n8612), .A(n7573), .ZN(n7580) );
  INV_X1 U9057 ( .A(n7580), .ZN(n10614) );
  OAI22_X1 U9058 ( .A1(n7575), .A2(n9762), .B1(n7826), .B2(n9764), .ZN(n7579)
         );
  XNOR2_X1 U9059 ( .A(n7576), .B(n8612), .ZN(n7577) );
  NOR2_X1 U9060 ( .A1(n7577), .A2(n9759), .ZN(n7578) );
  AOI211_X1 U9061 ( .C1(n7635), .C2(n7580), .A(n7579), .B(n7578), .ZN(n10612)
         );
  MUX2_X1 U9062 ( .A(n7167), .B(n10612), .S(n10524), .Z(n7587) );
  AOI211_X1 U9063 ( .C1(n10609), .C2(n7581), .A(n9797), .B(n7681), .ZN(n10608)
         );
  INV_X1 U9064 ( .A(n7582), .ZN(n7583) );
  OAI22_X1 U9065 ( .A1(n9802), .A2(n7584), .B1(n9854), .B2(n7583), .ZN(n7585)
         );
  AOI21_X1 U9066 ( .B1(n10608), .B2(n4924), .A(n7585), .ZN(n7586) );
  OAI211_X1 U9067 ( .C1(n10614), .C2(n7588), .A(n7587), .B(n7586), .ZN(
        P1_U3287) );
  INV_X1 U9068 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n7589) );
  OAI22_X1 U9069 ( .A1(n9327), .A2(n7414), .B1(n10764), .B2(n7589), .ZN(n7590)
         );
  INV_X1 U9070 ( .A(n7590), .ZN(n7591) );
  OAI21_X1 U9071 ( .B1(n7592), .B2(n6872), .A(n7591), .ZN(P2_U3393) );
  OAI21_X1 U9072 ( .B1(n7595), .B2(n7594), .A(n7593), .ZN(n7596) );
  AOI222_X1 U9073 ( .A1(n10546), .A2(n7596), .B1(n9504), .B2(n10543), .C1(
        n9506), .C2(n10541), .ZN(n10671) );
  OAI21_X1 U9074 ( .B1(n7598), .B2(n8618), .A(n7597), .ZN(n10674) );
  NAND2_X1 U9075 ( .A1(n7599), .A2(n7961), .ZN(n7600) );
  NAND2_X1 U9076 ( .A1(n7600), .A2(n10537), .ZN(n7601) );
  OR2_X1 U9077 ( .A1(n7739), .A2(n7601), .ZN(n10668) );
  INV_X1 U9078 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7603) );
  INV_X1 U9079 ( .A(n7955), .ZN(n7602) );
  OAI22_X1 U9080 ( .A1(n10524), .A2(n7603), .B1(n7602), .B2(n9854), .ZN(n7604)
         );
  AOI21_X1 U9081 ( .B1(n7961), .B2(n10552), .A(n7604), .ZN(n7605) );
  OAI21_X1 U9082 ( .B1(n10668), .B2(n9832), .A(n7605), .ZN(n7606) );
  AOI21_X1 U9083 ( .B1(n10674), .B2(n10559), .A(n7606), .ZN(n7607) );
  OAI21_X1 U9084 ( .B1(n10555), .B2(n10671), .A(n7607), .ZN(P1_U3283) );
  OAI222_X1 U9085 ( .A1(n7610), .A2(P2_U3151), .B1(n8052), .B2(n7609), .C1(
        n7608), .C2(n8237), .ZN(P2_U3279) );
  OAI211_X1 U9086 ( .C1(n7613), .C2(n7612), .A(n7611), .B(n8914), .ZN(n7618)
         );
  OAI22_X1 U9087 ( .A1(n7614), .A2(n8897), .B1(n8925), .B2(n10577), .ZN(n7615)
         );
  AOI211_X1 U9088 ( .C1(n8895), .C2(n8939), .A(n7616), .B(n7615), .ZN(n7617)
         );
  OAI211_X1 U9089 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n8919), .A(n7618), .B(
        n7617), .ZN(P2_U3158) );
  NAND2_X1 U9090 ( .A1(n10643), .A2(n10658), .ZN(n9178) );
  NOR2_X1 U9091 ( .A1(n10643), .A2(n7256), .ZN(n7625) );
  INV_X1 U9092 ( .A(n7619), .ZN(n7622) );
  INV_X1 U9093 ( .A(n7620), .ZN(n7621) );
  NAND3_X1 U9094 ( .A1(n8445), .A2(n7622), .A3(n7621), .ZN(n7623) );
  OAI21_X1 U9095 ( .B1(n9238), .B2(n10198), .A(n7623), .ZN(n7624) );
  AOI211_X1 U9096 ( .C1(n10641), .C2(n7626), .A(n7625), .B(n7624), .ZN(n7627)
         );
  OAI21_X1 U9097 ( .B1(n7628), .B2(n9178), .A(n7627), .ZN(P2_U3233) );
  INV_X1 U9098 ( .A(n7629), .ZN(n7691) );
  AOI22_X1 U9099 ( .A1(n9604), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n10012), .ZN(n7630) );
  OAI21_X1 U9100 ( .B1(n7691), .B2(n7945), .A(n7630), .ZN(P1_U3338) );
  NAND2_X1 U9101 ( .A1(n7631), .A2(n8505), .ZN(n7675) );
  OR2_X1 U9102 ( .A1(n7675), .A2(n8613), .ZN(n7673) );
  NAND2_X1 U9103 ( .A1(n7673), .A2(n8516), .ZN(n7647) );
  XNOR2_X1 U9104 ( .A(n7647), .B(n8614), .ZN(n7637) );
  OAI21_X1 U9105 ( .B1(n7633), .B2(n8614), .A(n7632), .ZN(n10633) );
  OAI22_X1 U9106 ( .A1(n7826), .A2(n9762), .B1(n7959), .B2(n9764), .ZN(n7634)
         );
  AOI21_X1 U9107 ( .B1(n10633), .B2(n7635), .A(n7634), .ZN(n7636) );
  OAI21_X1 U9108 ( .B1(n7637), .B2(n9759), .A(n7636), .ZN(n10631) );
  INV_X1 U9109 ( .A(n10631), .ZN(n7644) );
  OAI211_X1 U9110 ( .C1(n7682), .C2(n10630), .A(n10537), .B(n7654), .ZN(n10629) );
  AOI22_X1 U9111 ( .A1(n9800), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n7822), .B2(
        n10554), .ZN(n7640) );
  NAND2_X1 U9112 ( .A1(n7638), .A2(n10552), .ZN(n7639) );
  OAI211_X1 U9113 ( .C1(n10629), .C2(n9832), .A(n7640), .B(n7639), .ZN(n7641)
         );
  AOI21_X1 U9114 ( .B1(n10633), .B2(n7642), .A(n7641), .ZN(n7643) );
  OAI21_X1 U9115 ( .B1(n7644), .B2(n9800), .A(n7643), .ZN(P1_U3285) );
  INV_X1 U9116 ( .A(n8510), .ZN(n7646) );
  OAI21_X1 U9117 ( .B1(n7647), .B2(n7646), .A(n7645), .ZN(n7648) );
  XNOR2_X1 U9118 ( .A(n7648), .B(n8617), .ZN(n7650) );
  AND2_X1 U9119 ( .A1(n9507), .A2(n9821), .ZN(n7649) );
  AOI21_X1 U9120 ( .B1(n7650), .B2(n10546), .A(n7649), .ZN(n10653) );
  OR2_X1 U9121 ( .A1(n7651), .A2(n8617), .ZN(n7652) );
  NAND2_X1 U9122 ( .A1(n7653), .A2(n7652), .ZN(n10651) );
  INV_X1 U9123 ( .A(n7657), .ZN(n10649) );
  XNOR2_X1 U9124 ( .A(n7654), .B(n10649), .ZN(n7656) );
  AND2_X1 U9125 ( .A1(n9505), .A2(n10543), .ZN(n7655) );
  AOI21_X1 U9126 ( .B1(n7656), .B2(n10537), .A(n7655), .ZN(n10648) );
  AOI22_X1 U9127 ( .A1(n9800), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n7862), .B2(
        n10554), .ZN(n7659) );
  NAND2_X1 U9128 ( .A1(n7657), .A2(n10552), .ZN(n7658) );
  OAI211_X1 U9129 ( .C1(n10648), .C2(n9832), .A(n7659), .B(n7658), .ZN(n7660)
         );
  AOI21_X1 U9130 ( .B1(n10651), .B2(n10559), .A(n7660), .ZN(n7661) );
  OAI21_X1 U9131 ( .B1(n10653), .B2(n9800), .A(n7661), .ZN(P1_U3284) );
  NAND2_X1 U9132 ( .A1(n7662), .A2(n7663), .ZN(n7664) );
  XNOR2_X1 U9133 ( .A(n7664), .B(n7884), .ZN(n7705) );
  XNOR2_X1 U9134 ( .A(n7665), .B(n7884), .ZN(n7666) );
  AOI22_X1 U9135 ( .A1(n7666), .A2(n9211), .B1(n9216), .B2(n8938), .ZN(n7706)
         );
  OAI21_X1 U9136 ( .B1(n7750), .B2(n10754), .A(n7706), .ZN(n7667) );
  AOI21_X1 U9137 ( .B1(n10749), .B2(n7705), .A(n7667), .ZN(n7672) );
  INV_X1 U9138 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n7668) );
  OAI22_X1 U9139 ( .A1(n9327), .A2(n7715), .B1(n10764), .B2(n7668), .ZN(n7669)
         );
  INV_X1 U9140 ( .A(n7669), .ZN(n7670) );
  OAI21_X1 U9141 ( .B1(n7672), .B2(n6872), .A(n7670), .ZN(P2_U3408) );
  INV_X1 U9142 ( .A(n7715), .ZN(n7723) );
  AOI22_X1 U9143 ( .A1(n9293), .A2(n7723), .B1(n10760), .B2(
        P2_REG1_REG_6__SCAN_IN), .ZN(n7671) );
  OAI21_X1 U9144 ( .B1(n7672), .B2(n10760), .A(n7671), .ZN(P2_U3465) );
  INV_X1 U9145 ( .A(n7673), .ZN(n7674) );
  AOI21_X1 U9146 ( .B1(n8613), .B2(n7675), .A(n7674), .ZN(n7676) );
  OAI222_X1 U9147 ( .A1(n9764), .A2(n7678), .B1(n9762), .B2(n7677), .C1(n9759), 
        .C2(n7676), .ZN(n7727) );
  INV_X1 U9148 ( .A(n7727), .ZN(n7690) );
  OAI21_X1 U9149 ( .B1(n7680), .B2(n8613), .A(n7679), .ZN(n7729) );
  INV_X1 U9150 ( .A(n7681), .ZN(n7683) );
  AOI211_X1 U9151 ( .C1(n7684), .C2(n7683), .A(n9797), .B(n7682), .ZN(n7728)
         );
  NAND2_X1 U9152 ( .A1(n7728), .A2(n4924), .ZN(n7687) );
  AOI22_X1 U9153 ( .A1(n9800), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n7685), .B2(
        n10554), .ZN(n7686) );
  OAI211_X1 U9154 ( .C1(n7734), .C2(n9802), .A(n7687), .B(n7686), .ZN(n7688)
         );
  AOI21_X1 U9155 ( .B1(n7729), .B2(n10559), .A(n7688), .ZN(n7689) );
  OAI21_X1 U9156 ( .B1(n7690), .B2(n10555), .A(n7689), .ZN(P1_U3286) );
  INV_X1 U9157 ( .A(n9023), .ZN(n7692) );
  OAI222_X1 U9158 ( .A1(n7692), .A2(P2_U3151), .B1(n8237), .B2(n6002), .C1(
        n7691), .C2(n8052), .ZN(P2_U3278) );
  INV_X1 U9159 ( .A(n7693), .ZN(n7694) );
  NAND2_X1 U9160 ( .A1(n10683), .A2(n7694), .ZN(n7695) );
  INV_X1 U9161 ( .A(n7696), .ZN(n7697) );
  MUX2_X1 U9162 ( .A(n7697), .B(n7271), .S(n9223), .Z(n7701) );
  INV_X1 U9163 ( .A(n9178), .ZN(n9195) );
  OAI22_X1 U9164 ( .A1(n9225), .A2(n7414), .B1(n7698), .B2(n10638), .ZN(n7699)
         );
  AOI21_X1 U9165 ( .B1(n9195), .B2(n8941), .A(n7699), .ZN(n7700) );
  OAI211_X1 U9166 ( .C1(n7702), .C2(n9230), .A(n7701), .B(n7700), .ZN(P2_U3232) );
  INV_X1 U9167 ( .A(n7703), .ZN(n7725) );
  AOI22_X1 U9168 ( .A1(n10363), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n10012), .ZN(n7704) );
  OAI21_X1 U9169 ( .B1(n7725), .B2(n7945), .A(n7704), .ZN(P1_U3337) );
  INV_X1 U9170 ( .A(n7705), .ZN(n7710) );
  MUX2_X1 U9171 ( .A(n5665), .B(n7706), .S(n10643), .Z(n7709) );
  OAI22_X1 U9172 ( .A1(n9178), .A2(n7750), .B1(n7714), .B2(n10638), .ZN(n7707)
         );
  AOI21_X1 U9173 ( .B1(n10641), .B2(n7723), .A(n7707), .ZN(n7708) );
  OAI211_X1 U9174 ( .C1(n7710), .C2(n9230), .A(n7709), .B(n7708), .ZN(P2_U3227) );
  INV_X1 U9175 ( .A(n7750), .ZN(n8936) );
  NAND2_X1 U9176 ( .A1(P2_U3151), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n10448) );
  INV_X1 U9177 ( .A(n10448), .ZN(n7711) );
  AOI21_X1 U9178 ( .B1(n8895), .B2(n8936), .A(n7711), .ZN(n7713) );
  NAND2_X1 U9179 ( .A1(n8922), .A2(n8938), .ZN(n7712) );
  OAI211_X1 U9180 ( .C1(n8919), .C2(n7714), .A(n7713), .B(n7712), .ZN(n7722)
         );
  XNOR2_X1 U9181 ( .A(n7715), .B(n7924), .ZN(n7748) );
  XNOR2_X1 U9182 ( .A(n7748), .B(n8937), .ZN(n7720) );
  AOI211_X1 U9183 ( .C1(n7720), .C2(n7719), .A(n8912), .B(n7749), .ZN(n7721)
         );
  AOI211_X1 U9184 ( .C1(n7723), .C2(n8910), .A(n7722), .B(n7721), .ZN(n7724)
         );
  INV_X1 U9185 ( .A(n7724), .ZN(P2_U3179) );
  INV_X1 U9186 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7726) );
  OAI222_X1 U9187 ( .A1(n8237), .A2(n7726), .B1(P2_U3151), .B2(n10494), .C1(
        n7725), .C2(n8052), .ZN(P2_U3277) );
  AOI211_X1 U9188 ( .C1(n10675), .C2(n7729), .A(n7728), .B(n7727), .ZN(n7737)
         );
  INV_X1 U9189 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n7730) );
  OAI22_X1 U9190 ( .A1(n9934), .A2(n7734), .B1(n10677), .B2(n7730), .ZN(n7731)
         );
  INV_X1 U9191 ( .A(n7731), .ZN(n7732) );
  OAI21_X1 U9192 ( .B1(n7737), .B2(n10676), .A(n7732), .ZN(P1_U3529) );
  INV_X1 U9193 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n7733) );
  OAI22_X1 U9194 ( .A1(n9995), .A2(n7734), .B1(n10681), .B2(n7733), .ZN(n7735)
         );
  INV_X1 U9195 ( .A(n7735), .ZN(n7736) );
  OAI21_X1 U9196 ( .B1(n7737), .B2(n10678), .A(n7736), .ZN(P1_U3474) );
  NAND2_X1 U9197 ( .A1(n8700), .A2(n8530), .ZN(n8619) );
  XNOR2_X1 U9198 ( .A(n7738), .B(n8619), .ZN(n9852) );
  OAI21_X1 U9199 ( .B1(n7739), .B2(n8149), .A(n10537), .ZN(n7740) );
  NOR2_X1 U9200 ( .A1(n7740), .A2(n7801), .ZN(n9860) );
  XNOR2_X1 U9201 ( .A(n7741), .B(n8619), .ZN(n7742) );
  OAI222_X1 U9202 ( .A1(n9764), .A2(n9443), .B1(n9762), .B2(n7860), .C1(n7742), 
        .C2(n9759), .ZN(n9859) );
  AOI211_X1 U9203 ( .C1(n10675), .C2(n9852), .A(n9860), .B(n9859), .ZN(n7747)
         );
  AOI22_X1 U9204 ( .A1(n9858), .A2(n9940), .B1(n10676), .B2(
        P1_REG1_REG_11__SCAN_IN), .ZN(n7743) );
  OAI21_X1 U9205 ( .B1(n7747), .B2(n10676), .A(n7743), .ZN(P1_U3533) );
  INV_X1 U9206 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n7744) );
  OAI22_X1 U9207 ( .A1(n8149), .A2(n9995), .B1(n10681), .B2(n7744), .ZN(n7745)
         );
  INV_X1 U9208 ( .A(n7745), .ZN(n7746) );
  OAI21_X1 U9209 ( .B1(n7747), .B2(n10678), .A(n7746), .ZN(P1_U3486) );
  XNOR2_X1 U9210 ( .A(n7758), .B(n8796), .ZN(n7846) );
  XNOR2_X1 U9211 ( .A(n7846), .B(n7750), .ZN(n7751) );
  OAI21_X1 U9212 ( .B1(n5022), .B2(n7751), .A(n7848), .ZN(n7752) );
  NAND2_X1 U9213 ( .A1(n7752), .A2(n8914), .ZN(n7757) );
  INV_X1 U9214 ( .A(n7893), .ZN(n7755) );
  AND2_X1 U9215 ( .A1(P2_U3151), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n10452) );
  AOI21_X1 U9216 ( .B1(n8895), .B2(n10620), .A(n10452), .ZN(n7753) );
  OAI21_X1 U9217 ( .B1(n8897), .B2(n10601), .A(n7753), .ZN(n7754) );
  AOI21_X1 U9218 ( .B1(n8899), .B2(n7755), .A(n7754), .ZN(n7756) );
  OAI211_X1 U9219 ( .C1(n7758), .C2(n8925), .A(n7757), .B(n7756), .ZN(P2_U3153) );
  NOR2_X1 U9220 ( .A1(n8266), .A2(n10740), .ZN(n10565) );
  NOR2_X1 U9221 ( .A1(n9238), .A2(n7300), .ZN(n7764) );
  XNOR2_X1 U9222 ( .A(n7759), .B(n7768), .ZN(n7761) );
  NAND2_X1 U9223 ( .A1(n7761), .A2(n9211), .ZN(n7763) );
  AOI22_X1 U9224 ( .A1(n9216), .A2(n8942), .B1(n8940), .B2(n10658), .ZN(n7762)
         );
  NAND2_X1 U9225 ( .A1(n7763), .A2(n7762), .ZN(n10564) );
  AOI211_X1 U9226 ( .C1(n10565), .C2(n7765), .A(n7764), .B(n10564), .ZN(n7771)
         );
  NOR2_X1 U9227 ( .A1(n7767), .A2(n7766), .ZN(n7769) );
  XNOR2_X1 U9228 ( .A(n7769), .B(n7768), .ZN(n10566) );
  AOI22_X1 U9229 ( .A1(n10566), .A2(n10639), .B1(n9223), .B2(
        P2_REG2_REG_2__SCAN_IN), .ZN(n7770) );
  OAI21_X1 U9230 ( .B1(n7771), .B2(n9223), .A(n7770), .ZN(P2_U3231) );
  INV_X1 U9231 ( .A(n7772), .ZN(n7832) );
  AOI22_X1 U9232 ( .A1(n4926), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n10012), .ZN(n7773) );
  OAI21_X1 U9233 ( .B1(n7832), .B2(n7945), .A(n7773), .ZN(P1_U3336) );
  XNOR2_X1 U9234 ( .A(n7774), .B(n8447), .ZN(n10584) );
  INV_X1 U9235 ( .A(n8447), .ZN(n7775) );
  XNOR2_X1 U9236 ( .A(n7776), .B(n7775), .ZN(n7777) );
  NAND2_X1 U9237 ( .A1(n7777), .A2(n9211), .ZN(n7779) );
  AOI22_X1 U9238 ( .A1(n10658), .A2(n8938), .B1(n8940), .B2(n9216), .ZN(n7778)
         );
  AND2_X1 U9239 ( .A1(n7779), .A2(n7778), .ZN(n10588) );
  MUX2_X1 U9240 ( .A(n10588), .B(n5661), .S(n9223), .Z(n7782) );
  AOI22_X1 U9241 ( .A1(n10641), .A2(n10585), .B1(n9222), .B2(n7780), .ZN(n7781) );
  OAI211_X1 U9242 ( .C1(n9230), .C2(n10584), .A(n7782), .B(n7781), .ZN(
        P2_U3229) );
  OAI21_X1 U9243 ( .B1(n7785), .B2(n7784), .A(n7783), .ZN(n10580) );
  OAI22_X1 U9244 ( .A1(n9225), .A2(n10577), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n10638), .ZN(n7791) );
  XNOR2_X1 U9245 ( .A(n7786), .B(n8446), .ZN(n7787) );
  NAND2_X1 U9246 ( .A1(n7787), .A2(n9211), .ZN(n7789) );
  AOI22_X1 U9247 ( .A1(n9216), .A2(n8941), .B1(n8939), .B2(n10658), .ZN(n7788)
         );
  NAND2_X1 U9248 ( .A1(n7789), .A2(n7788), .ZN(n10578) );
  MUX2_X1 U9249 ( .A(n10578), .B(P2_REG2_REG_3__SCAN_IN), .S(n9223), .Z(n7790)
         );
  AOI211_X1 U9250 ( .C1(n10639), .C2(n10580), .A(n7791), .B(n7790), .ZN(n7792)
         );
  INV_X1 U9251 ( .A(n7792), .ZN(P2_U3230) );
  XOR2_X1 U9252 ( .A(n7793), .B(n8621), .Z(n7836) );
  INV_X1 U9253 ( .A(n7836), .ZN(n7808) );
  INV_X1 U9254 ( .A(n8621), .ZN(n7794) );
  NAND3_X1 U9255 ( .A1(n7795), .A2(n7794), .A3(n8530), .ZN(n7796) );
  NAND2_X1 U9256 ( .A1(n7797), .A2(n7796), .ZN(n7798) );
  NAND2_X1 U9257 ( .A1(n7798), .A2(n10546), .ZN(n7800) );
  AOI22_X1 U9258 ( .A1(n10541), .A2(n9504), .B1(n9502), .B2(n10543), .ZN(n7799) );
  NAND2_X1 U9259 ( .A1(n7800), .A2(n7799), .ZN(n7834) );
  INV_X1 U9260 ( .A(n7801), .ZN(n7803) );
  INV_X1 U9261 ( .A(n7934), .ZN(n7802) );
  AOI211_X1 U9262 ( .C1(n8542), .C2(n7803), .A(n9797), .B(n7802), .ZN(n7835)
         );
  NAND2_X1 U9263 ( .A1(n7835), .A2(n4924), .ZN(n7805) );
  AOI22_X1 U9264 ( .A1(n9800), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n8199), .B2(
        n10554), .ZN(n7804) );
  OAI211_X1 U9265 ( .C1(n7838), .C2(n9802), .A(n7805), .B(n7804), .ZN(n7806)
         );
  AOI21_X1 U9266 ( .B1(n10524), .B2(n7834), .A(n7806), .ZN(n7807) );
  OAI21_X1 U9267 ( .B1(n7808), .B2(n9836), .A(n7807), .ZN(P1_U3281) );
  NAND2_X1 U9268 ( .A1(n7809), .A2(n7810), .ZN(n7811) );
  XNOR2_X1 U9269 ( .A(n7811), .B(n8452), .ZN(n10640) );
  XNOR2_X1 U9270 ( .A(n7812), .B(n8452), .ZN(n7813) );
  AOI222_X1 U9271 ( .A1(n9211), .A2(n7813), .B1(n8936), .B2(n9216), .C1(n8015), 
        .C2(n10658), .ZN(n10637) );
  INV_X1 U9272 ( .A(n10637), .ZN(n7814) );
  AOI21_X1 U9273 ( .B1(n10749), .B2(n10640), .A(n7814), .ZN(n7819) );
  INV_X1 U9274 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n7815) );
  NOR2_X1 U9275 ( .A1(n10764), .A2(n7815), .ZN(n7816) );
  AOI21_X1 U9276 ( .B1(n6880), .B2(n10642), .A(n7816), .ZN(n7817) );
  OAI21_X1 U9277 ( .B1(n7819), .B2(n6872), .A(n7817), .ZN(P2_U3414) );
  AOI22_X1 U9278 ( .A1(n9293), .A2(n10642), .B1(n10760), .B2(
        P2_REG1_REG_8__SCAN_IN), .ZN(n7818) );
  OAI21_X1 U9279 ( .B1(n7819), .B2(n10760), .A(n7818), .ZN(P2_U3467) );
  OAI21_X1 U9280 ( .B1(n7821), .B2(n5023), .A(n7820), .ZN(n7829) );
  NOR2_X1 U9281 ( .A1(n10630), .A2(n9480), .ZN(n7828) );
  NAND2_X1 U9282 ( .A1(n9486), .A2(n7822), .ZN(n7825) );
  NAND2_X1 U9283 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n10309) );
  INV_X1 U9284 ( .A(n10309), .ZN(n7823) );
  AOI21_X1 U9285 ( .B1(n9488), .B2(n9506), .A(n7823), .ZN(n7824) );
  OAI211_X1 U9286 ( .C1(n7826), .C2(n9491), .A(n7825), .B(n7824), .ZN(n7827)
         );
  AOI211_X1 U9287 ( .C1(n7829), .C2(n9472), .A(n7828), .B(n7827), .ZN(n7830)
         );
  INV_X1 U9288 ( .A(n7830), .ZN(P1_U3221) );
  OAI222_X1 U9289 ( .A1(n7833), .A2(P2_U3151), .B1(n8052), .B2(n7832), .C1(
        n7831), .C2(n8237), .ZN(P2_U3276) );
  AOI211_X1 U9290 ( .C1(n7836), .C2(n10675), .A(n7835), .B(n7834), .ZN(n7842)
         );
  INV_X1 U9291 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n7837) );
  OAI22_X1 U9292 ( .A1(n7838), .A2(n9995), .B1(n10681), .B2(n7837), .ZN(n7839)
         );
  INV_X1 U9293 ( .A(n7839), .ZN(n7840) );
  OAI21_X1 U9294 ( .B1(n7842), .B2(n10678), .A(n7840), .ZN(P1_U3489) );
  AOI22_X1 U9295 ( .A1(n8542), .A2(n9940), .B1(n10676), .B2(
        P1_REG1_REG_12__SCAN_IN), .ZN(n7841) );
  OAI21_X1 U9296 ( .B1(n7842), .B2(n10676), .A(n7841), .ZN(P1_U3534) );
  INV_X1 U9297 ( .A(n7843), .ZN(n7866) );
  NAND2_X1 U9298 ( .A1(n10003), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n7844) );
  OAI211_X1 U9299 ( .C1(n7866), .C2(n7945), .A(n7845), .B(n7844), .ZN(P1_U3335) );
  XNOR2_X1 U9300 ( .A(n10642), .B(n8796), .ZN(n7920) );
  XNOR2_X1 U9301 ( .A(n7920), .B(n10620), .ZN(n7922) );
  INV_X1 U9302 ( .A(n7846), .ZN(n7847) );
  XOR2_X1 U9303 ( .A(n7922), .B(n7923), .Z(n7853) );
  NOR2_X1 U9304 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5872), .ZN(n10472) );
  AOI21_X1 U9305 ( .B1(n8895), .B2(n8015), .A(n10472), .ZN(n7850) );
  NAND2_X1 U9306 ( .A1(n8922), .A2(n8936), .ZN(n7849) );
  OAI211_X1 U9307 ( .C1(n8919), .C2(n5525), .A(n7850), .B(n7849), .ZN(n7851)
         );
  AOI21_X1 U9308 ( .B1(n10642), .B2(n8910), .A(n7851), .ZN(n7852) );
  OAI21_X1 U9309 ( .B1(n7853), .B2(n8912), .A(n7852), .ZN(P2_U3161) );
  OAI21_X1 U9310 ( .B1(n7856), .B2(n7854), .A(n7855), .ZN(n7857) );
  NAND2_X1 U9311 ( .A1(n7857), .A2(n9472), .ZN(n7864) );
  AOI21_X1 U9312 ( .B1(n9451), .B2(n9507), .A(n7858), .ZN(n7859) );
  OAI21_X1 U9313 ( .B1(n7860), .B2(n9434), .A(n7859), .ZN(n7861) );
  AOI21_X1 U9314 ( .B1(n7862), .B2(n9486), .A(n7861), .ZN(n7863) );
  OAI211_X1 U9315 ( .C1(n10649), .C2(n9480), .A(n7864), .B(n7863), .ZN(
        P1_U3231) );
  OAI222_X1 U9316 ( .A1(P2_U3151), .A2(n7409), .B1(n8052), .B2(n7866), .C1(
        n7865), .C2(n8237), .ZN(P2_U3275) );
  AOI21_X1 U9317 ( .B1(n8034), .B2(n7868), .A(n7867), .ZN(n7883) );
  INV_X1 U9318 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n7875) );
  AOI21_X1 U9319 ( .B1(n7871), .B2(n7870), .A(n7869), .ZN(n7873) );
  OR2_X1 U9320 ( .A1(n7873), .A2(n7872), .ZN(n7874) );
  OR2_X1 U9321 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10195), .ZN(n7927) );
  OAI211_X1 U9322 ( .C1(n10489), .C2(n7875), .A(n7874), .B(n7927), .ZN(n7880)
         );
  AOI21_X1 U9323 ( .B1(n10665), .B2(n7877), .A(n7876), .ZN(n7878) );
  NOR2_X1 U9324 ( .A1(n7878), .A2(n10501), .ZN(n7879) );
  AOI211_X1 U9325 ( .C1(n10474), .C2(n7881), .A(n7880), .B(n7879), .ZN(n7882)
         );
  OAI21_X1 U9326 ( .B1(n7883), .B2(n10506), .A(n7882), .ZN(P2_U3191) );
  NAND2_X1 U9327 ( .A1(n7665), .A2(n7884), .ZN(n7886) );
  NAND2_X1 U9328 ( .A1(n7886), .A2(n7885), .ZN(n7887) );
  XNOR2_X1 U9329 ( .A(n7887), .B(n8453), .ZN(n7888) );
  NAND2_X1 U9330 ( .A1(n7888), .A2(n9211), .ZN(n7890) );
  NAND2_X1 U9331 ( .A1(n8937), .A2(n9216), .ZN(n7889) );
  NAND2_X1 U9332 ( .A1(n7890), .A2(n7889), .ZN(n10623) );
  NAND2_X1 U9333 ( .A1(n7891), .A2(n8453), .ZN(n7892) );
  NAND2_X1 U9334 ( .A1(n7809), .A2(n7892), .ZN(n10622) );
  OAI22_X1 U9335 ( .A1(n10643), .A2(n10456), .B1(n7893), .B2(n10638), .ZN(
        n7894) );
  AOI21_X1 U9336 ( .B1(n9195), .B2(n10620), .A(n7894), .ZN(n7896) );
  NAND2_X1 U9337 ( .A1(n10641), .A2(n10619), .ZN(n7895) );
  OAI211_X1 U9338 ( .C1(n10622), .C2(n9230), .A(n7896), .B(n7895), .ZN(n7897)
         );
  AOI21_X1 U9339 ( .B1(n10647), .B2(n10623), .A(n7897), .ZN(n7898) );
  INV_X1 U9340 ( .A(n7898), .ZN(P2_U3226) );
  AOI21_X1 U9341 ( .B1(n7901), .B2(n7900), .A(n7899), .ZN(n7917) );
  INV_X1 U9342 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n7902) );
  NAND2_X1 U9343 ( .A1(P2_U3151), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n8013) );
  OAI21_X1 U9344 ( .B1(n10489), .B2(n7902), .A(n8013), .ZN(n7907) );
  AOI21_X1 U9345 ( .B1(n5020), .B2(n7904), .A(n7903), .ZN(n7905) );
  NOR2_X1 U9346 ( .A1(n7905), .A2(n10501), .ZN(n7906) );
  AOI211_X1 U9347 ( .C1(n10474), .C2(n7908), .A(n7907), .B(n7906), .ZN(n7916)
         );
  INV_X1 U9348 ( .A(n7909), .ZN(n7910) );
  NOR2_X1 U9349 ( .A1(n7911), .A2(n7910), .ZN(n7913) );
  XOR2_X1 U9350 ( .A(n7913), .B(n7912), .Z(n7914) );
  NAND2_X1 U9351 ( .A1(n7914), .A2(n10495), .ZN(n7915) );
  OAI211_X1 U9352 ( .C1(n7917), .C2(n10506), .A(n7916), .B(n7915), .ZN(
        P2_U3192) );
  INV_X1 U9353 ( .A(n7918), .ZN(n7950) );
  AOI22_X1 U9354 ( .A1(n8635), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n10012), .ZN(n7919) );
  OAI21_X1 U9355 ( .B1(n7950), .B2(n7945), .A(n7919), .ZN(P1_U3334) );
  INV_X1 U9356 ( .A(n5895), .ZN(n7932) );
  XNOR2_X1 U9357 ( .A(n5895), .B(n8796), .ZN(n7977) );
  XNOR2_X1 U9358 ( .A(n7977), .B(n8015), .ZN(n7925) );
  OAI211_X1 U9359 ( .C1(n7926), .C2(n7925), .A(n7976), .B(n8914), .ZN(n7931)
         );
  OAI21_X1 U9360 ( .B1(n8918), .B2(n8035), .A(n7927), .ZN(n7929) );
  NOR2_X1 U9361 ( .A1(n8919), .A2(n8033), .ZN(n7928) );
  AOI211_X1 U9362 ( .C1(n8922), .C2(n10620), .A(n7929), .B(n7928), .ZN(n7930)
         );
  OAI211_X1 U9363 ( .C1(n7932), .C2(n8925), .A(n7931), .B(n7930), .ZN(P2_U3171) );
  XNOR2_X1 U9364 ( .A(n7933), .B(n8622), .ZN(n9841) );
  AOI21_X1 U9365 ( .B1(n7934), .B2(n9846), .A(n9797), .ZN(n7935) );
  AND2_X1 U9366 ( .A1(n7935), .A2(n5018), .ZN(n9847) );
  XOR2_X1 U9367 ( .A(n8622), .B(n7936), .Z(n7937) );
  OAI222_X1 U9368 ( .A1(n9764), .A2(n9492), .B1(n9762), .B2(n9443), .C1(n7937), 
        .C2(n9759), .ZN(n9840) );
  AOI211_X1 U9369 ( .C1(n9841), .C2(n10675), .A(n9847), .B(n9840), .ZN(n7942)
         );
  INV_X1 U9370 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n8114) );
  AOI22_X1 U9371 ( .A1(n9846), .A2(n9940), .B1(n10676), .B2(
        P1_REG1_REG_13__SCAN_IN), .ZN(n7938) );
  OAI21_X1 U9372 ( .B1(n7942), .B2(n10676), .A(n7938), .ZN(P1_U3535) );
  INV_X1 U9373 ( .A(n9846), .ZN(n8549) );
  INV_X1 U9374 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n7939) );
  OAI22_X1 U9375 ( .A1(n8549), .A2(n9995), .B1(n10681), .B2(n7939), .ZN(n7940)
         );
  INV_X1 U9376 ( .A(n7940), .ZN(n7941) );
  OAI21_X1 U9377 ( .B1(n7942), .B2(n10678), .A(n7941), .ZN(P1_U3492) );
  INV_X1 U9378 ( .A(n7943), .ZN(n7947) );
  AOI22_X1 U9379 ( .A1(n8739), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n10012), .ZN(n7944) );
  OAI21_X1 U9380 ( .B1(n7947), .B2(n7945), .A(n7944), .ZN(P1_U3333) );
  OAI222_X1 U9381 ( .A1(n7948), .A2(P2_U3151), .B1(n8052), .B2(n7947), .C1(
        n7946), .C2(n8237), .ZN(P2_U3273) );
  INV_X1 U9382 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7949) );
  OAI222_X1 U9383 ( .A1(P2_U3151), .A2(n8254), .B1(n8052), .B2(n7950), .C1(
        n7949), .C2(n8237), .ZN(P2_U3274) );
  INV_X1 U9384 ( .A(n7951), .ZN(n7952) );
  AOI21_X1 U9385 ( .B1(n7954), .B2(n7953), .A(n7952), .ZN(n7963) );
  NAND2_X1 U9386 ( .A1(n9486), .A2(n7955), .ZN(n7958) );
  NAND2_X1 U9387 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n10391) );
  INV_X1 U9388 ( .A(n10391), .ZN(n7956) );
  AOI21_X1 U9389 ( .B1(n9488), .B2(n9504), .A(n7956), .ZN(n7957) );
  OAI211_X1 U9390 ( .C1(n7959), .C2(n9491), .A(n7958), .B(n7957), .ZN(n7960)
         );
  AOI21_X1 U9391 ( .B1(n7961), .B2(n9494), .A(n7960), .ZN(n7962) );
  OAI21_X1 U9392 ( .B1(n7963), .B2(n9496), .A(n7962), .ZN(P1_U3217) );
  XNOR2_X1 U9393 ( .A(n7964), .B(n8623), .ZN(n7965) );
  AOI222_X1 U9394 ( .A1(n10546), .A2(n7965), .B1(n9820), .B2(n10543), .C1(
        n9502), .C2(n10541), .ZN(n9946) );
  INV_X1 U9395 ( .A(n7966), .ZN(n7967) );
  AOI21_X1 U9396 ( .B1(n8623), .B2(n7968), .A(n7967), .ZN(n9942) );
  AOI21_X1 U9397 ( .B1(n5018), .B2(n9943), .A(n9797), .ZN(n7969) );
  NAND2_X1 U9398 ( .A1(n7969), .A2(n8088), .ZN(n9945) );
  INV_X1 U9399 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7971) );
  INV_X1 U9400 ( .A(n9353), .ZN(n7970) );
  OAI22_X1 U9401 ( .A1(n10524), .A2(n7971), .B1(n7970), .B2(n9854), .ZN(n7972)
         );
  AOI21_X1 U9402 ( .B1(n9943), .B2(n10552), .A(n7972), .ZN(n7973) );
  OAI21_X1 U9403 ( .B1(n9945), .B2(n9832), .A(n7973), .ZN(n7974) );
  AOI21_X1 U9404 ( .B1(n9942), .B2(n10559), .A(n7974), .ZN(n7975) );
  OAI21_X1 U9405 ( .B1(n10555), .B2(n9946), .A(n7975), .ZN(P1_U3279) );
  XNOR2_X1 U9406 ( .A(n10695), .B(n8796), .ZN(n8101) );
  XNOR2_X1 U9407 ( .A(n10685), .B(n7984), .ZN(n8099) );
  INV_X1 U9408 ( .A(n8099), .ZN(n7978) );
  OAI22_X1 U9409 ( .A1(n8101), .A2(n10686), .B1(n8035), .B2(n7978), .ZN(n7982)
         );
  OAI21_X1 U9410 ( .B1(n8099), .B2(n10657), .A(n8073), .ZN(n7980) );
  NOR2_X1 U9411 ( .A1(n8073), .A2(n10657), .ZN(n7979) );
  AOI22_X1 U9412 ( .A1(n8101), .A2(n7980), .B1(n7979), .B2(n7978), .ZN(n7981)
         );
  INV_X2 U9413 ( .A(n7984), .ZN(n8796) );
  XNOR2_X1 U9414 ( .A(n8459), .B(n8796), .ZN(n8153) );
  XOR2_X1 U9415 ( .A(n8154), .B(n8153), .Z(n7989) );
  NAND2_X1 U9416 ( .A1(P2_U3151), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n8172) );
  OAI21_X1 U9417 ( .B1(n8918), .B2(n9235), .A(n8172), .ZN(n7985) );
  AOI21_X1 U9418 ( .B1(n8922), .B2(n8073), .A(n7985), .ZN(n7986) );
  OAI21_X1 U9419 ( .B1(n8919), .B2(n8075), .A(n7986), .ZN(n7987) );
  AOI21_X1 U9420 ( .B1(n10708), .B2(n8910), .A(n7987), .ZN(n7988) );
  OAI21_X1 U9421 ( .B1(n7989), .B2(n8912), .A(n7988), .ZN(P2_U3164) );
  XNOR2_X1 U9422 ( .A(n7990), .B(n6271), .ZN(n10711) );
  NAND2_X1 U9423 ( .A1(n7991), .A2(n8325), .ZN(n7992) );
  NAND3_X1 U9424 ( .A1(n7993), .A2(n9211), .A3(n7992), .ZN(n7995) );
  AOI22_X1 U9425 ( .A1(n10658), .A2(n9215), .B1(n8935), .B2(n9216), .ZN(n7994)
         );
  NAND2_X1 U9426 ( .A1(n7995), .A2(n7994), .ZN(n10712) );
  INV_X1 U9427 ( .A(n10714), .ZN(n8162) );
  OAI22_X1 U9428 ( .A1(n8162), .A2(n9240), .B1(n8157), .B2(n10638), .ZN(n7996)
         );
  OAI21_X1 U9429 ( .B1(n10712), .B2(n7996), .A(n10647), .ZN(n7998) );
  NAND2_X1 U9430 ( .A1(n9223), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n7997) );
  OAI211_X1 U9431 ( .C1(n9230), .C2(n10711), .A(n7998), .B(n7997), .ZN(
        P2_U3220) );
  NAND2_X1 U9432 ( .A1(n8000), .A2(n7999), .ZN(n8001) );
  XNOR2_X1 U9433 ( .A(n8001), .B(n8448), .ZN(n8003) );
  OAI22_X1 U9434 ( .A1(n8003), .A2(n9234), .B1(n8002), .B2(n9236), .ZN(n10602)
         );
  INV_X1 U9435 ( .A(n10602), .ZN(n8012) );
  OAI22_X1 U9436 ( .A1(n10647), .A2(n10421), .B1(n8004), .B2(n10638), .ZN(
        n8006) );
  NOR2_X1 U9437 ( .A1(n9178), .A2(n10601), .ZN(n8005) );
  AOI211_X1 U9438 ( .C1(n10641), .C2(n8007), .A(n8006), .B(n8005), .ZN(n8011)
         );
  AND2_X1 U9439 ( .A1(n8008), .A2(n8448), .ZN(n10599) );
  INV_X1 U9440 ( .A(n10599), .ZN(n8009) );
  NAND3_X1 U9441 ( .A1(n8009), .A2(n10639), .A3(n7662), .ZN(n8010) );
  OAI211_X1 U9442 ( .C1(n8012), .C2(n9223), .A(n8011), .B(n8010), .ZN(P2_U3228) );
  XNOR2_X1 U9443 ( .A(n8098), .B(n8099), .ZN(n8100) );
  XNOR2_X1 U9444 ( .A(n8100), .B(n8035), .ZN(n8019) );
  OAI21_X1 U9445 ( .B1(n8918), .B2(n10686), .A(n8013), .ZN(n8014) );
  AOI21_X1 U9446 ( .B1(n8922), .B2(n8015), .A(n8014), .ZN(n8016) );
  OAI21_X1 U9447 ( .B1(n8919), .B2(n8044), .A(n8016), .ZN(n8017) );
  AOI21_X1 U9448 ( .B1(n10685), .B2(n8910), .A(n8017), .ZN(n8018) );
  OAI21_X1 U9449 ( .B1(n8019), .B2(n8912), .A(n8018), .ZN(P2_U3157) );
  XOR2_X1 U9450 ( .A(n8020), .B(n8458), .Z(n10694) );
  XNOR2_X1 U9451 ( .A(n8021), .B(n8458), .ZN(n8022) );
  OAI22_X1 U9452 ( .A1(n8022), .A2(n9234), .B1(n8035), .B2(n9236), .ZN(n10698)
         );
  NAND2_X1 U9453 ( .A1(n10698), .A2(n10643), .ZN(n8026) );
  NOR2_X1 U9454 ( .A1(n9178), .A2(n10696), .ZN(n8024) );
  OAI22_X1 U9455 ( .A1(n10647), .A2(n8056), .B1(n8107), .B2(n10638), .ZN(n8023) );
  AOI211_X1 U9456 ( .C1(n10695), .C2(n10641), .A(n8024), .B(n8023), .ZN(n8025)
         );
  OAI211_X1 U9457 ( .C1(n10694), .C2(n9230), .A(n8026), .B(n8025), .ZN(
        P2_U3222) );
  INV_X1 U9458 ( .A(n8027), .ZN(n8028) );
  AOI21_X1 U9459 ( .B1(n8454), .B2(n8029), .A(n8028), .ZN(n10663) );
  INV_X1 U9460 ( .A(n10663), .ZN(n10660) );
  XOR2_X1 U9461 ( .A(n8030), .B(n8454), .Z(n8032) );
  OAI22_X1 U9462 ( .A1(n8032), .A2(n9234), .B1(n8031), .B2(n9236), .ZN(n10661)
         );
  NAND2_X1 U9463 ( .A1(n10661), .A2(n10643), .ZN(n8039) );
  OAI22_X1 U9464 ( .A1(n10647), .A2(n8034), .B1(n8033), .B2(n10638), .ZN(n8037) );
  NOR2_X1 U9465 ( .A1(n9178), .A2(n8035), .ZN(n8036) );
  AOI211_X1 U9466 ( .C1(n10641), .C2(n5895), .A(n8037), .B(n8036), .ZN(n8038)
         );
  OAI211_X1 U9467 ( .C1(n10660), .C2(n9230), .A(n8039), .B(n8038), .ZN(
        P2_U3224) );
  NAND2_X1 U9468 ( .A1(n8027), .A2(n8284), .ZN(n8040) );
  XNOR2_X1 U9469 ( .A(n8040), .B(n8457), .ZN(n10682) );
  XNOR2_X1 U9470 ( .A(n8041), .B(n8457), .ZN(n8043) );
  OAI22_X1 U9471 ( .A1(n8043), .A2(n9234), .B1(n8042), .B2(n9236), .ZN(n10690)
         );
  NAND2_X1 U9472 ( .A1(n10690), .A2(n10643), .ZN(n8048) );
  OAI22_X1 U9473 ( .A1(n10647), .A2(n5670), .B1(n8044), .B2(n10638), .ZN(n8046) );
  NOR2_X1 U9474 ( .A1(n9178), .A2(n10686), .ZN(n8045) );
  AOI211_X1 U9475 ( .C1(n10685), .C2(n10641), .A(n8046), .B(n8045), .ZN(n8047)
         );
  OAI211_X1 U9476 ( .C1(n10682), .C2(n9230), .A(n8048), .B(n8047), .ZN(
        P2_U3223) );
  INV_X1 U9477 ( .A(n8049), .ZN(n8054) );
  NAND2_X1 U9478 ( .A1(n9345), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n8051) );
  NAND2_X1 U9479 ( .A1(n8050), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8486) );
  OAI211_X1 U9480 ( .C1(n8054), .C2(n8052), .A(n8051), .B(n8486), .ZN(P2_U3272) );
  NAND2_X1 U9481 ( .A1(n10003), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n8053) );
  OAI211_X1 U9482 ( .C1(n8054), .C2(n7945), .A(n8738), .B(n8053), .ZN(P1_U3332) );
  AOI21_X1 U9483 ( .B1(n8057), .B2(n8056), .A(n8055), .ZN(n8071) );
  INV_X1 U9484 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n8063) );
  OAI21_X1 U9485 ( .B1(n8060), .B2(n8059), .A(n8058), .ZN(n8061) );
  NAND2_X1 U9486 ( .A1(n8061), .A2(n10495), .ZN(n8062) );
  NAND2_X1 U9487 ( .A1(P2_U3151), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n8104) );
  OAI211_X1 U9488 ( .C1(n10489), .C2(n8063), .A(n8062), .B(n8104), .ZN(n8068)
         );
  AOI21_X1 U9489 ( .B1(n10701), .B2(n8065), .A(n8064), .ZN(n8066) );
  NOR2_X1 U9490 ( .A1(n8066), .A2(n10501), .ZN(n8067) );
  AOI211_X1 U9491 ( .C1(n10474), .C2(n8069), .A(n8068), .B(n8067), .ZN(n8070)
         );
  OAI21_X1 U9492 ( .B1(n8071), .B2(n10506), .A(n8070), .ZN(P2_U3193) );
  XNOR2_X1 U9493 ( .A(n8072), .B(n8459), .ZN(n8074) );
  AOI222_X1 U9494 ( .A1(n9211), .A2(n8074), .B1(n8073), .B2(n9216), .C1(n8934), 
        .C2(n10658), .ZN(n10705) );
  OAI22_X1 U9495 ( .A1(n10647), .A2(n5935), .B1(n8075), .B2(n10638), .ZN(n8078) );
  XOR2_X1 U9496 ( .A(n8076), .B(n8459), .Z(n10704) );
  NOR2_X1 U9497 ( .A1(n10704), .A2(n9230), .ZN(n8077) );
  AOI211_X1 U9498 ( .C1(n10641), .C2(n10708), .A(n8078), .B(n8077), .ZN(n8079)
         );
  OAI21_X1 U9499 ( .B1(n9223), .B2(n10705), .A(n8079), .ZN(P2_U3221) );
  NAND2_X1 U9500 ( .A1(n8080), .A2(n8625), .ZN(n8081) );
  NAND2_X1 U9501 ( .A1(n9812), .A2(n8081), .ZN(n8082) );
  NAND2_X1 U9502 ( .A1(n8082), .A2(n10546), .ZN(n8084) );
  AOI22_X1 U9503 ( .A1(n10541), .A2(n9501), .B1(n9500), .B2(n10543), .ZN(n8083) );
  AND2_X1 U9504 ( .A1(n8084), .A2(n8083), .ZN(n9936) );
  OR2_X1 U9505 ( .A1(n8085), .A2(n8625), .ZN(n8086) );
  NAND2_X1 U9506 ( .A1(n8087), .A2(n8086), .ZN(n9938) );
  INV_X1 U9507 ( .A(n9938), .ZN(n8096) );
  INV_X1 U9508 ( .A(n9825), .ZN(n8090) );
  AOI21_X1 U9509 ( .B1(n8088), .B2(n9998), .A(n9797), .ZN(n8089) );
  NAND2_X1 U9510 ( .A1(n8090), .A2(n8089), .ZN(n9935) );
  INV_X1 U9511 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n8092) );
  INV_X1 U9512 ( .A(n9485), .ZN(n8091) );
  OAI22_X1 U9513 ( .A1(n10524), .A2(n8092), .B1(n8091), .B2(n9854), .ZN(n8093)
         );
  AOI21_X1 U9514 ( .B1(n9998), .B2(n10552), .A(n8093), .ZN(n8094) );
  OAI21_X1 U9515 ( .B1(n9935), .B2(n9832), .A(n8094), .ZN(n8095) );
  AOI21_X1 U9516 ( .B1(n8096), .B2(n10559), .A(n8095), .ZN(n8097) );
  OAI21_X1 U9517 ( .B1(n10555), .B2(n9936), .A(n8097), .ZN(P1_U3278) );
  OAI22_X1 U9518 ( .A1(n8100), .A2(n10657), .B1(n8099), .B2(n8098), .ZN(n8103)
         );
  XNOR2_X1 U9519 ( .A(n8101), .B(n10686), .ZN(n8102) );
  XNOR2_X1 U9520 ( .A(n8103), .B(n8102), .ZN(n8110) );
  OAI21_X1 U9521 ( .B1(n8918), .B2(n10696), .A(n8104), .ZN(n8105) );
  AOI21_X1 U9522 ( .B1(n8922), .B2(n10657), .A(n8105), .ZN(n8106) );
  OAI21_X1 U9523 ( .B1(n8919), .B2(n8107), .A(n8106), .ZN(n8108) );
  AOI21_X1 U9524 ( .B1(n10695), .B2(n8910), .A(n8108), .ZN(n8109) );
  OAI21_X1 U9525 ( .B1(n8110), .B2(n8912), .A(n8109), .ZN(P2_U3176) );
  INV_X1 U9526 ( .A(n8111), .ZN(n8224) );
  AOI22_X1 U9527 ( .A1(n8112), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n10012), .ZN(n8113) );
  OAI21_X1 U9528 ( .B1(n8224), .B2(n7945), .A(n8113), .ZN(P1_U3331) );
  INV_X1 U9529 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9932) );
  INV_X1 U9530 ( .A(n8214), .ZN(n8122) );
  AOI22_X1 U9531 ( .A1(n8214), .A2(P1_REG1_REG_16__SCAN_IN), .B1(n9932), .B2(
        n8122), .ZN(n8119) );
  MUX2_X1 U9532 ( .A(n8114), .B(P1_REG1_REG_13__SCAN_IN), .S(n10375), .Z(
        n10368) );
  OAI21_X1 U9533 ( .B1(n8124), .B2(P1_REG1_REG_12__SCAN_IN), .A(n8115), .ZN(
        n10369) );
  NOR2_X1 U9534 ( .A1(n10368), .A2(n10369), .ZN(n10367) );
  AOI21_X1 U9535 ( .B1(n10375), .B2(P1_REG1_REG_13__SCAN_IN), .A(n10367), .ZN(
        n10331) );
  XNOR2_X1 U9536 ( .A(n10324), .B(P1_REG1_REG_14__SCAN_IN), .ZN(n10332) );
  NOR2_X1 U9537 ( .A1(n10331), .A2(n10332), .ZN(n10330) );
  AOI21_X1 U9538 ( .B1(P1_REG1_REG_14__SCAN_IN), .B2(n10324), .A(n10330), .ZN(
        n8116) );
  NOR2_X1 U9539 ( .A1(n8116), .A2(n8128), .ZN(n8117) );
  INV_X1 U9540 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n10344) );
  XNOR2_X1 U9541 ( .A(n8128), .B(n8116), .ZN(n10345) );
  NOR2_X1 U9542 ( .A1(n10344), .A2(n10345), .ZN(n10343) );
  NOR2_X1 U9543 ( .A1(n8117), .A2(n10343), .ZN(n8118) );
  NAND2_X1 U9544 ( .A1(n8119), .A2(n8118), .ZN(n8213) );
  OAI21_X1 U9545 ( .B1(n8119), .B2(n8118), .A(n8213), .ZN(n8135) );
  NOR2_X1 U9546 ( .A1(n8120), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9399) );
  AOI21_X1 U9547 ( .B1(n9607), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n9399), .ZN(
        n8121) );
  OAI21_X1 U9548 ( .B1(n10338), .B2(n8122), .A(n8121), .ZN(n8134) );
  OAI21_X1 U9549 ( .B1(n8124), .B2(P1_REG2_REG_12__SCAN_IN), .A(n8123), .ZN(
        n10372) );
  NAND2_X1 U9550 ( .A1(n10375), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n8125) );
  OAI21_X1 U9551 ( .B1(n10375), .B2(P1_REG2_REG_13__SCAN_IN), .A(n8125), .ZN(
        n10371) );
  NOR2_X1 U9552 ( .A1(n10372), .A2(n10371), .ZN(n10370) );
  AOI21_X1 U9553 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(n10375), .A(n10370), .ZN(
        n10326) );
  NAND2_X1 U9554 ( .A1(n10324), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n8126) );
  OAI21_X1 U9555 ( .B1(n10324), .B2(P1_REG2_REG_14__SCAN_IN), .A(n8126), .ZN(
        n10327) );
  NOR2_X1 U9556 ( .A1(n10326), .A2(n10327), .ZN(n10325) );
  AOI21_X1 U9557 ( .B1(P1_REG2_REG_14__SCAN_IN), .B2(n10324), .A(n10325), .ZN(
        n8127) );
  NOR2_X1 U9558 ( .A1(n8127), .A2(n8128), .ZN(n8129) );
  XNOR2_X1 U9559 ( .A(n8128), .B(n8127), .ZN(n10347) );
  NOR2_X1 U9560 ( .A1(n8092), .A2(n10347), .ZN(n10346) );
  NOR2_X1 U9561 ( .A1(n8129), .A2(n10346), .ZN(n8132) );
  NAND2_X1 U9562 ( .A1(n8214), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n8130) );
  OAI21_X1 U9563 ( .B1(n8214), .B2(P1_REG2_REG_16__SCAN_IN), .A(n8130), .ZN(
        n8131) );
  NOR2_X1 U9564 ( .A1(n8132), .A2(n8131), .ZN(n8208) );
  AOI211_X1 U9565 ( .C1(n8132), .C2(n8131), .A(n8208), .B(n10383), .ZN(n8133)
         );
  AOI211_X1 U9566 ( .C1(n10334), .C2(n8135), .A(n8134), .B(n8133), .ZN(n8136)
         );
  INV_X1 U9567 ( .A(n8136), .ZN(P1_U3259) );
  INV_X1 U9568 ( .A(n8140), .ZN(n8137) );
  NOR2_X1 U9569 ( .A1(n8138), .A2(n8137), .ZN(n8143) );
  AOI21_X1 U9570 ( .B1(n8141), .B2(n8140), .A(n8139), .ZN(n8142) );
  OAI21_X1 U9571 ( .B1(n8143), .B2(n8142), .A(n9472), .ZN(n8148) );
  NAND2_X1 U9572 ( .A1(P1_U3086), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n10321) );
  INV_X1 U9573 ( .A(n10321), .ZN(n8144) );
  AOI21_X1 U9574 ( .B1(n9451), .B2(n9505), .A(n8144), .ZN(n8145) );
  OAI21_X1 U9575 ( .B1(n9443), .B2(n9434), .A(n8145), .ZN(n8146) );
  AOI21_X1 U9576 ( .B1(n9853), .B2(n9486), .A(n8146), .ZN(n8147) );
  OAI211_X1 U9577 ( .C1(n8149), .C2(n9480), .A(n8148), .B(n8147), .ZN(P1_U3236) );
  INV_X1 U9578 ( .A(n8150), .ZN(n8151) );
  MUX2_X1 U9579 ( .A(n8151), .B(n8307), .S(n8796), .Z(n8152) );
  XNOR2_X1 U9580 ( .A(n10714), .B(n8796), .ZN(n8229) );
  XNOR2_X1 U9581 ( .A(n8229), .B(n8934), .ZN(n8155) );
  NAND2_X1 U9582 ( .A1(n8156), .A2(n8155), .ZN(n8228) );
  OAI211_X1 U9583 ( .C1(n8156), .C2(n8155), .A(n8228), .B(n8914), .ZN(n8161)
         );
  NAND2_X1 U9584 ( .A1(P2_U3151), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n8951) );
  OAI21_X1 U9585 ( .B1(n8918), .B2(n8758), .A(n8951), .ZN(n8159) );
  NOR2_X1 U9586 ( .A1(n8919), .A2(n8157), .ZN(n8158) );
  AOI211_X1 U9587 ( .C1(n8922), .C2(n8935), .A(n8159), .B(n8158), .ZN(n8160)
         );
  OAI211_X1 U9588 ( .C1(n8162), .C2(n8925), .A(n8161), .B(n8160), .ZN(P2_U3174) );
  INV_X1 U9589 ( .A(n8164), .ZN(n8165) );
  AOI21_X1 U9590 ( .B1(n8167), .B2(n8166), .A(n8165), .ZN(n8182) );
  INV_X1 U9591 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n8174) );
  OAI21_X1 U9592 ( .B1(n8170), .B2(n8169), .A(n8168), .ZN(n8171) );
  NAND2_X1 U9593 ( .A1(n8171), .A2(n10495), .ZN(n8173) );
  OAI211_X1 U9594 ( .C1(n10489), .C2(n8174), .A(n8173), .B(n8172), .ZN(n8179)
         );
  NAND2_X1 U9595 ( .A1(n5009), .A2(n8175), .ZN(n8176) );
  AOI21_X1 U9596 ( .B1(n8177), .B2(n8176), .A(n10501), .ZN(n8178) );
  AOI211_X1 U9597 ( .C1(n10474), .C2(n8180), .A(n8179), .B(n8178), .ZN(n8181)
         );
  OAI21_X1 U9598 ( .B1(n8182), .B2(n10506), .A(n8181), .ZN(P2_U3194) );
  OAI21_X1 U9599 ( .B1(n8184), .B2(n8626), .A(n8183), .ZN(n9927) );
  NAND2_X1 U9600 ( .A1(n9925), .A2(n9824), .ZN(n8185) );
  NAND2_X1 U9601 ( .A1(n8185), .A2(n10537), .ZN(n8186) );
  NOR2_X1 U9602 ( .A1(n9794), .A2(n8186), .ZN(n9924) );
  INV_X1 U9603 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n8189) );
  NAND2_X1 U9604 ( .A1(n9925), .A2(n10552), .ZN(n8188) );
  NAND2_X1 U9605 ( .A1(n10554), .A2(n9414), .ZN(n8187) );
  OAI211_X1 U9606 ( .C1(n10524), .C2(n8189), .A(n8188), .B(n8187), .ZN(n8190)
         );
  AOI21_X1 U9607 ( .B1(n9924), .B2(n4924), .A(n8190), .ZN(n8196) );
  OAI211_X1 U9608 ( .C1(n8192), .C2(n8560), .A(n8191), .B(n10546), .ZN(n8194)
         );
  NAND2_X1 U9609 ( .A1(n9500), .A2(n9821), .ZN(n8193) );
  OAI211_X1 U9610 ( .C1(n9412), .C2(n9764), .A(n8194), .B(n8193), .ZN(n9923)
         );
  NAND2_X1 U9611 ( .A1(n9923), .A2(n10524), .ZN(n8195) );
  OAI211_X1 U9612 ( .C1(n9927), .C2(n9836), .A(n8196), .B(n8195), .ZN(P1_U3276) );
  XOR2_X1 U9613 ( .A(n8197), .B(n8198), .Z(n8206) );
  NAND2_X1 U9614 ( .A1(n9486), .A2(n8199), .ZN(n8202) );
  AOI21_X1 U9615 ( .B1(n9488), .B2(n9502), .A(n8200), .ZN(n8201) );
  OAI211_X1 U9616 ( .C1(n8203), .C2(n9491), .A(n8202), .B(n8201), .ZN(n8204)
         );
  AOI21_X1 U9617 ( .B1(n8542), .B2(n9494), .A(n8204), .ZN(n8205) );
  OAI21_X1 U9618 ( .B1(n8206), .B2(n9496), .A(n8205), .ZN(P1_U3224) );
  NOR2_X1 U9619 ( .A1(n9604), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n8207) );
  AOI21_X1 U9620 ( .B1(P1_REG2_REG_17__SCAN_IN), .B2(n9604), .A(n8207), .ZN(
        n8210) );
  AOI21_X1 U9621 ( .B1(P1_REG2_REG_16__SCAN_IN), .B2(n8214), .A(n8208), .ZN(
        n8209) );
  NAND2_X1 U9622 ( .A1(n8210), .A2(n8209), .ZN(n9598) );
  OAI21_X1 U9623 ( .B1(n8210), .B2(n8209), .A(n9598), .ZN(n8211) );
  INV_X1 U9624 ( .A(n8211), .ZN(n8222) );
  INV_X1 U9625 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n8212) );
  INV_X1 U9626 ( .A(n9604), .ZN(n8218) );
  AOI22_X1 U9627 ( .A1(n9604), .A2(P1_REG1_REG_17__SCAN_IN), .B1(n8212), .B2(
        n8218), .ZN(n8216) );
  OAI21_X1 U9628 ( .B1(n8214), .B2(P1_REG1_REG_16__SCAN_IN), .A(n8213), .ZN(
        n8215) );
  NAND2_X1 U9629 ( .A1(n8216), .A2(n8215), .ZN(n9603) );
  OAI21_X1 U9630 ( .B1(n8216), .B2(n8215), .A(n9603), .ZN(n8220) );
  NAND2_X1 U9631 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9410) );
  NAND2_X1 U9632 ( .A1(n9607), .A2(P1_ADDR_REG_17__SCAN_IN), .ZN(n8217) );
  OAI211_X1 U9633 ( .C1(n10338), .C2(n8218), .A(n9410), .B(n8217), .ZN(n8219)
         );
  AOI21_X1 U9634 ( .B1(n8220), .B2(n10334), .A(n8219), .ZN(n8221) );
  OAI21_X1 U9635 ( .B1(n8222), .B2(n10383), .A(n8221), .ZN(P1_U3260) );
  OAI222_X1 U9636 ( .A1(P2_U3151), .A2(n6298), .B1(n8052), .B2(n8224), .C1(
        n8223), .C2(n8237), .ZN(P2_U3271) );
  INV_X1 U9637 ( .A(n8225), .ZN(n8239) );
  AOI22_X1 U9638 ( .A1(n8226), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n10012), .ZN(n8227) );
  OAI21_X1 U9639 ( .B1(n8239), .B2(n7945), .A(n8227), .ZN(P1_U3330) );
  XNOR2_X1 U9640 ( .A(n8328), .B(n8796), .ZN(n8759) );
  XNOR2_X1 U9641 ( .A(n8759), .B(n8758), .ZN(n8231) );
  AOI21_X1 U9642 ( .B1(n8231), .B2(n8230), .A(n8761), .ZN(n8236) );
  NAND2_X1 U9643 ( .A1(P2_U3151), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n8968) );
  OAI21_X1 U9644 ( .B1(n8918), .B2(n9237), .A(n8968), .ZN(n8232) );
  AOI21_X1 U9645 ( .B1(n8922), .B2(n8934), .A(n8232), .ZN(n8233) );
  OAI21_X1 U9646 ( .B1(n8919), .B2(n9239), .A(n8233), .ZN(n8234) );
  AOI21_X1 U9647 ( .B1(n8328), .B2(n8910), .A(n8234), .ZN(n8235) );
  OAI21_X1 U9648 ( .B1(n8236), .B2(n8912), .A(n8235), .ZN(P2_U3155) );
  OAI222_X1 U9649 ( .A1(n8240), .A2(P2_U3151), .B1(n8052), .B2(n8239), .C1(
        n8238), .C2(n8237), .ZN(P2_U3270) );
  INV_X1 U9650 ( .A(n8241), .ZN(n8245) );
  AOI22_X1 U9651 ( .A1(n6786), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n10012), .ZN(n8242) );
  OAI21_X1 U9652 ( .B1(n8245), .B2(n7945), .A(n8242), .ZN(P1_U3329) );
  AOI22_X1 U9653 ( .A1(n8243), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n9345), .ZN(n8244) );
  OAI21_X1 U9654 ( .B1(n8245), .B2(n8052), .A(n8244), .ZN(P2_U3269) );
  INV_X1 U9655 ( .A(n8246), .ZN(n8251) );
  AOI22_X1 U9656 ( .A1(n8247), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n10012), .ZN(n8248) );
  OAI21_X1 U9657 ( .B1(n8251), .B2(n7945), .A(n8248), .ZN(P1_U3328) );
  AOI21_X1 U9658 ( .B1(P1_DATAO_REG_27__SCAN_IN), .B2(n9345), .A(n8249), .ZN(
        n8250) );
  OAI21_X1 U9659 ( .B1(n8251), .B2(n8052), .A(n8250), .ZN(P2_U3268) );
  MUX2_X1 U9660 ( .A(n8928), .B(n9045), .S(n8387), .Z(n8390) );
  INV_X1 U9661 ( .A(n8390), .ZN(n8394) );
  MUX2_X1 U9662 ( .A(n9328), .B(n9148), .S(n8387), .Z(n8356) );
  NOR2_X1 U9663 ( .A1(n9331), .A2(n8825), .ZN(n8253) );
  MUX2_X1 U9664 ( .A(n8253), .B(n8252), .S(n8387), .Z(n8354) );
  NAND2_X1 U9665 ( .A1(n8255), .A2(n8254), .ZN(n8257) );
  NAND4_X1 U9666 ( .A1(n8449), .A2(n8257), .A3(n8261), .A4(n8256), .ZN(n8258)
         );
  NAND3_X1 U9667 ( .A1(n8259), .A2(n8258), .A3(n8275), .ZN(n8260) );
  INV_X1 U9668 ( .A(n8261), .ZN(n8262) );
  NAND2_X1 U9669 ( .A1(n8263), .A2(n8262), .ZN(n8264) );
  NAND2_X1 U9670 ( .A1(n8264), .A2(n8256), .ZN(n8265) );
  NAND2_X1 U9671 ( .A1(n8265), .A2(n8449), .ZN(n8269) );
  MUX2_X1 U9672 ( .A(n8295), .B(n8276), .S(n8387), .Z(n8273) );
  NAND2_X1 U9673 ( .A1(n8274), .A2(n8273), .ZN(n8298) );
  INV_X1 U9674 ( .A(n8275), .ZN(n8277) );
  OAI211_X1 U9675 ( .C1(n8298), .C2(n8277), .A(n8299), .B(n8276), .ZN(n8281)
         );
  NAND2_X1 U9676 ( .A1(n8301), .A2(n8296), .ZN(n8279) );
  AOI21_X1 U9677 ( .B1(n8279), .B2(n8278), .A(n8387), .ZN(n8280) );
  NAND2_X1 U9678 ( .A1(n8281), .A2(n8280), .ZN(n8285) );
  AND2_X1 U9679 ( .A1(n8287), .A2(n8286), .ZN(n8289) );
  OAI211_X1 U9680 ( .C1(n8290), .C2(n8289), .A(n8314), .B(n8288), .ZN(n8291)
         );
  NAND2_X1 U9681 ( .A1(n8291), .A2(n8396), .ZN(n8292) );
  INV_X1 U9682 ( .A(n8294), .ZN(n8297) );
  OAI211_X1 U9683 ( .C1(n8298), .C2(n8297), .A(n8296), .B(n8295), .ZN(n8300)
         );
  NAND2_X1 U9684 ( .A1(n8300), .A2(n8299), .ZN(n8302) );
  NAND2_X1 U9685 ( .A1(n8302), .A2(n8301), .ZN(n8303) );
  NAND2_X1 U9686 ( .A1(n8303), .A2(n8387), .ZN(n8304) );
  NAND2_X1 U9687 ( .A1(n8316), .A2(n8305), .ZN(n8306) );
  OAI21_X1 U9688 ( .B1(n8313), .B2(n8306), .A(n8318), .ZN(n8308) );
  AOI21_X1 U9689 ( .B1(n8308), .B2(n8459), .A(n8307), .ZN(n8321) );
  AOI21_X1 U9690 ( .B1(n8311), .B2(n8310), .A(n8309), .ZN(n8312) );
  NAND2_X1 U9691 ( .A1(n8313), .A2(n8312), .ZN(n8315) );
  NAND2_X1 U9692 ( .A1(n8315), .A2(n8314), .ZN(n8317) );
  NAND2_X1 U9693 ( .A1(n8317), .A2(n8316), .ZN(n8320) );
  AND2_X1 U9694 ( .A1(n8459), .A2(n8318), .ZN(n8319) );
  MUX2_X1 U9695 ( .A(n8323), .B(n8322), .S(n8396), .Z(n8324) );
  NOR2_X1 U9696 ( .A1(n9213), .A2(n8326), .ZN(n8333) );
  NAND2_X1 U9697 ( .A1(n8330), .A2(n8758), .ZN(n8327) );
  INV_X1 U9698 ( .A(n8328), .ZN(n10718) );
  NAND2_X1 U9699 ( .A1(n8329), .A2(n10718), .ZN(n8331) );
  MUX2_X1 U9700 ( .A(n8387), .B(n9217), .S(n8848), .Z(n8335) );
  AOI21_X1 U9701 ( .B1(n8917), .B2(n8396), .A(n8335), .ZN(n8336) );
  MUX2_X1 U9702 ( .A(n9201), .B(n10741), .S(n8387), .Z(n8340) );
  NAND2_X1 U9703 ( .A1(n8343), .A2(n10741), .ZN(n8338) );
  NAND2_X1 U9704 ( .A1(n8342), .A2(n9201), .ZN(n8337) );
  MUX2_X1 U9705 ( .A(n8338), .B(n8337), .S(n8387), .Z(n8339) );
  AOI21_X1 U9706 ( .B1(n8341), .B2(n8340), .A(n8339), .ZN(n8347) );
  INV_X1 U9707 ( .A(n8342), .ZN(n8345) );
  INV_X1 U9708 ( .A(n8343), .ZN(n8344) );
  MUX2_X1 U9709 ( .A(n8345), .B(n8344), .S(n8387), .Z(n8346) );
  INV_X1 U9710 ( .A(n8349), .ZN(n8352) );
  INV_X1 U9711 ( .A(n8350), .ZN(n8351) );
  MUX2_X1 U9712 ( .A(n8352), .B(n8351), .S(n8387), .Z(n8353) );
  INV_X1 U9713 ( .A(n8356), .ZN(n8358) );
  NAND2_X1 U9714 ( .A1(n8358), .A2(n8357), .ZN(n8360) );
  XNOR2_X1 U9715 ( .A(n8779), .B(n8833), .ZN(n9117) );
  MUX2_X1 U9716 ( .A(n8362), .B(n8361), .S(n8387), .Z(n8363) );
  NAND2_X1 U9717 ( .A1(n8365), .A2(n8465), .ZN(n8376) );
  INV_X1 U9718 ( .A(n8366), .ZN(n8369) );
  INV_X1 U9719 ( .A(n8367), .ZN(n8368) );
  MUX2_X1 U9720 ( .A(n8369), .B(n8368), .S(n8387), .Z(n8370) );
  NOR2_X1 U9721 ( .A1(n9096), .A2(n8370), .ZN(n8375) );
  MUX2_X1 U9722 ( .A(n8372), .B(n8371), .S(n8387), .Z(n8374) );
  NAND2_X1 U9723 ( .A1(n8377), .A2(n8373), .ZN(n9080) );
  INV_X1 U9724 ( .A(n8377), .ZN(n8379) );
  MUX2_X1 U9725 ( .A(n8379), .B(n8378), .S(n8387), .Z(n8380) );
  NOR3_X1 U9726 ( .A1(n8381), .A2(n9062), .A3(n8380), .ZN(n8386) );
  NOR2_X1 U9727 ( .A1(n8382), .A2(n8929), .ZN(n8384) );
  MUX2_X1 U9728 ( .A(n8384), .B(n8383), .S(n8387), .Z(n8385) );
  MUX2_X1 U9729 ( .A(n8389), .B(n8388), .S(n8387), .Z(n8392) );
  INV_X1 U9730 ( .A(n8395), .ZN(n8438) );
  INV_X1 U9731 ( .A(n8397), .ZN(n8398) );
  NAND2_X1 U9732 ( .A1(n8398), .A2(SI_29_), .ZN(n8404) );
  INV_X1 U9733 ( .A(n8399), .ZN(n8402) );
  INV_X1 U9734 ( .A(n8400), .ZN(n8401) );
  NAND2_X1 U9735 ( .A1(n8402), .A2(n8401), .ZN(n8403) );
  NAND2_X1 U9736 ( .A1(n8404), .A2(n8403), .ZN(n8415) );
  INV_X1 U9737 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8406) );
  INV_X1 U9738 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8405) );
  MUX2_X1 U9739 ( .A(n8406), .B(n8405), .S(n8416), .Z(n8408) );
  INV_X1 U9740 ( .A(SI_30_), .ZN(n8407) );
  NAND2_X1 U9741 ( .A1(n8408), .A2(n8407), .ZN(n8413) );
  INV_X1 U9742 ( .A(n8408), .ZN(n8409) );
  NAND2_X1 U9743 ( .A1(n8409), .A2(SI_30_), .ZN(n8410) );
  NAND2_X1 U9744 ( .A1(n8413), .A2(n8410), .ZN(n8414) );
  NAND2_X1 U9745 ( .A1(n9338), .A2(n5981), .ZN(n8412) );
  NAND2_X1 U9746 ( .A1(n6072), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n8411) );
  NOR2_X1 U9747 ( .A1(n9305), .A2(n8927), .ZN(n8434) );
  NAND2_X1 U9748 ( .A1(n9305), .A2(n8927), .ZN(n8470) );
  OAI21_X1 U9749 ( .B1(n8415), .B2(n8414), .A(n8413), .ZN(n8420) );
  MUX2_X1 U9750 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n8416), .Z(n8418) );
  INV_X1 U9751 ( .A(SI_31_), .ZN(n8417) );
  XNOR2_X1 U9752 ( .A(n8418), .B(n8417), .ZN(n8419) );
  XNOR2_X1 U9753 ( .A(n8420), .B(n8419), .ZN(n9334) );
  NAND2_X1 U9754 ( .A1(n9334), .A2(n5981), .ZN(n8422) );
  NAND2_X1 U9755 ( .A1(n6072), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n8421) );
  INV_X1 U9756 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n8423) );
  OR2_X1 U9757 ( .A1(n8424), .A2(n8423), .ZN(n8430) );
  INV_X1 U9758 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n8425) );
  OR2_X1 U9759 ( .A1(n8426), .A2(n8425), .ZN(n8429) );
  INV_X1 U9760 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n8427) );
  OR2_X1 U9761 ( .A1(n5857), .A2(n8427), .ZN(n8428) );
  NAND2_X1 U9762 ( .A1(n9030), .A2(n9033), .ZN(n8443) );
  INV_X1 U9763 ( .A(n8434), .ZN(n8469) );
  INV_X1 U9764 ( .A(n9033), .ZN(n8926) );
  NAND2_X1 U9765 ( .A1(n8470), .A2(n8926), .ZN(n8440) );
  INV_X1 U9766 ( .A(n8443), .ZN(n8474) );
  INV_X1 U9767 ( .A(n8444), .ZN(n8473) );
  INV_X1 U9768 ( .A(n9096), .ZN(n8466) );
  NOR4_X1 U9769 ( .A1(n8447), .A2(n8446), .A3(n6248), .A4(n8445), .ZN(n8450)
         );
  NAND4_X1 U9770 ( .A1(n8451), .A2(n8450), .A3(n5830), .A4(n8449), .ZN(n8455)
         );
  NOR4_X1 U9771 ( .A1(n8455), .A2(n8454), .A3(n8453), .A4(n8452), .ZN(n8456)
         );
  NAND4_X1 U9772 ( .A1(n8459), .A2(n8458), .A3(n8457), .A4(n8456), .ZN(n8460)
         );
  NOR4_X1 U9773 ( .A1(n9213), .A2(n9232), .A3(n6271), .A4(n8460), .ZN(n8462)
         );
  INV_X1 U9774 ( .A(n9203), .ZN(n8461) );
  NAND3_X1 U9775 ( .A1(n9173), .A2(n8462), .A3(n8461), .ZN(n8463) );
  NOR4_X1 U9776 ( .A1(n9154), .A2(n9190), .A3(n9159), .A4(n8463), .ZN(n8464)
         );
  NAND4_X1 U9777 ( .A1(n8466), .A2(n8465), .A3(n8464), .A4(n9134), .ZN(n8467)
         );
  NAND4_X1 U9778 ( .A1(n4966), .A2(n8468), .A3(n8797), .A4(n9069), .ZN(n8472)
         );
  NAND2_X1 U9779 ( .A1(n8470), .A2(n8469), .ZN(n8471) );
  NOR4_X1 U9780 ( .A1(n8474), .A2(n8473), .A3(n8472), .A4(n8471), .ZN(n8475)
         );
  NAND3_X1 U9781 ( .A1(n8482), .A2(n8481), .A3(n8480), .ZN(n8483) );
  OAI211_X1 U9782 ( .C1(n8484), .C2(n8486), .A(n8483), .B(P2_B_REG_SCAN_IN), 
        .ZN(n8485) );
  OAI21_X1 U9783 ( .B1(n8487), .B2(n8486), .A(n8485), .ZN(P2_U3296) );
  NAND2_X1 U9784 ( .A1(n4926), .A2(n8598), .ZN(n8591) );
  INV_X1 U9785 ( .A(n8591), .ZN(n8597) );
  NAND2_X1 U9786 ( .A1(n9334), .A2(n6490), .ZN(n8490) );
  NAND2_X1 U9787 ( .A1(n6405), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n8489) );
  NAND2_X1 U9788 ( .A1(n8490), .A2(n8489), .ZN(n8596) );
  NAND2_X1 U9789 ( .A1(n8491), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n8494) );
  NAND2_X1 U9790 ( .A1(n6400), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n8493) );
  NAND2_X1 U9791 ( .A1(n6441), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n8492) );
  AND3_X1 U9792 ( .A1(n8494), .A2(n8493), .A3(n8492), .ZN(n8668) );
  INV_X1 U9793 ( .A(n8668), .ZN(n9616) );
  MUX2_X1 U9794 ( .A(n8659), .B(n8639), .S(n8591), .Z(n8590) );
  INV_X1 U9795 ( .A(n8495), .ZN(n8496) );
  NAND2_X1 U9796 ( .A1(n8499), .A2(n8498), .ZN(n8686) );
  NAND2_X1 U9797 ( .A1(n8501), .A2(n8512), .ZN(n8690) );
  OAI21_X1 U9798 ( .B1(n8500), .B2(n8690), .A(n8514), .ZN(n8504) );
  INV_X1 U9799 ( .A(n8500), .ZN(n8502) );
  INV_X1 U9800 ( .A(n8514), .ZN(n8691) );
  OAI21_X1 U9801 ( .B1(n8502), .B2(n8691), .A(n8501), .ZN(n8503) );
  INV_X1 U9802 ( .A(n8505), .ZN(n8507) );
  OAI211_X1 U9803 ( .C1(n8513), .C2(n8507), .A(n8516), .B(n8506), .ZN(n8509)
         );
  INV_X1 U9804 ( .A(n8614), .ZN(n8517) );
  NAND3_X1 U9805 ( .A1(n8509), .A2(n8517), .A3(n8508), .ZN(n8511) );
  NAND3_X1 U9806 ( .A1(n8511), .A2(n8526), .A3(n8510), .ZN(n8524) );
  INV_X1 U9807 ( .A(n8512), .ZN(n8515) );
  OAI211_X1 U9808 ( .C1(n8519), .C2(n8518), .A(n8517), .B(n8516), .ZN(n8522)
         );
  INV_X1 U9809 ( .A(n8520), .ZN(n8521) );
  NAND2_X1 U9810 ( .A1(n8522), .A2(n8521), .ZN(n8523) );
  OAI211_X1 U9811 ( .C1(n5114), .C2(n8525), .A(n8700), .B(n8534), .ZN(n8531)
         );
  INV_X1 U9812 ( .A(n8526), .ZN(n8527) );
  NAND2_X1 U9813 ( .A1(n8534), .A2(n8527), .ZN(n8528) );
  NAND3_X1 U9814 ( .A1(n8530), .A2(n8529), .A3(n8528), .ZN(n8702) );
  MUX2_X1 U9815 ( .A(n8531), .B(n8702), .S(n8591), .Z(n8537) );
  INV_X1 U9816 ( .A(n8537), .ZN(n8532) );
  OAI21_X1 U9817 ( .B1(n8535), .B2(n5114), .A(n8532), .ZN(n8550) );
  NAND2_X1 U9818 ( .A1(n9443), .A2(n8591), .ZN(n8539) );
  INV_X1 U9819 ( .A(n8539), .ZN(n8533) );
  AOI22_X1 U9820 ( .A1(n8542), .A2(n8533), .B1(n9357), .B2(n8591), .ZN(n8548)
         );
  INV_X1 U9821 ( .A(n8534), .ZN(n8697) );
  NOR2_X1 U9822 ( .A1(n8535), .A2(n8697), .ZN(n8538) );
  AND4_X1 U9823 ( .A1(n8707), .A2(n8701), .A3(n8700), .A4(n8591), .ZN(n8536)
         );
  OAI21_X1 U9824 ( .B1(n8538), .B2(n8537), .A(n8536), .ZN(n8547) );
  NAND2_X1 U9825 ( .A1(n9503), .A2(n8597), .ZN(n8540) );
  OAI22_X1 U9826 ( .A1(n8542), .A2(n8540), .B1(n9357), .B2(n8591), .ZN(n8545)
         );
  OAI21_X1 U9827 ( .B1(n9502), .B2(n8539), .A(n8542), .ZN(n8544) );
  NOR2_X1 U9828 ( .A1(n8540), .A2(n9357), .ZN(n8541) );
  OR2_X1 U9829 ( .A1(n8542), .A2(n8541), .ZN(n8543) );
  AOI22_X1 U9830 ( .A1(n8549), .A2(n8545), .B1(n8544), .B2(n8543), .ZN(n8546)
         );
  NAND2_X1 U9831 ( .A1(n8554), .A2(n8708), .ZN(n8552) );
  NAND2_X1 U9832 ( .A1(n9813), .A2(n8711), .ZN(n8551) );
  MUX2_X1 U9833 ( .A(n8552), .B(n8551), .S(n8597), .Z(n8553) );
  INV_X1 U9834 ( .A(n8554), .ZN(n8713) );
  NAND2_X1 U9835 ( .A1(n8555), .A2(n8716), .ZN(n8559) );
  INV_X1 U9836 ( .A(n8556), .ZN(n8557) );
  INV_X1 U9837 ( .A(n8716), .ZN(n9818) );
  AOI21_X1 U9838 ( .B1(n8557), .B2(n8712), .A(n9818), .ZN(n8558) );
  OAI21_X1 U9839 ( .B1(n8568), .B2(n5136), .A(n8591), .ZN(n8569) );
  NAND2_X1 U9840 ( .A1(n8570), .A2(n8569), .ZN(n8571) );
  OAI211_X1 U9841 ( .C1(n8597), .C2(n8572), .A(n8571), .B(n9747), .ZN(n8575)
         );
  MUX2_X1 U9842 ( .A(n8721), .B(n8573), .S(n8591), .Z(n8574) );
  INV_X1 U9843 ( .A(n9724), .ZN(n9731) );
  AOI21_X1 U9844 ( .B1(n8575), .B2(n8574), .A(n9731), .ZN(n8581) );
  NAND2_X1 U9845 ( .A1(n8578), .A2(n8576), .ZN(n8647) );
  NAND2_X1 U9846 ( .A1(n8648), .A2(n8577), .ZN(n8640) );
  MUX2_X1 U9847 ( .A(n8647), .B(n8640), .S(n8591), .Z(n8580) );
  MUX2_X1 U9848 ( .A(n8648), .B(n8578), .S(n8591), .Z(n8579) );
  OAI211_X1 U9849 ( .C1(n8581), .C2(n8580), .A(n9685), .B(n8579), .ZN(n8582)
         );
  NAND4_X1 U9850 ( .A1(n8582), .A2(n8653), .A3(n8649), .A4(n8591), .ZN(n8587)
         );
  INV_X1 U9851 ( .A(n9667), .ZN(n9671) );
  NAND4_X1 U9852 ( .A1(n8582), .A2(n9671), .A3(n8597), .A4(n8645), .ZN(n8586)
         );
  OAI21_X1 U9853 ( .B1(n9689), .B2(n8591), .A(n9883), .ZN(n8584) );
  INV_X1 U9854 ( .A(n9883), .ZN(n9396) );
  OAI21_X1 U9855 ( .B1(n9476), .B2(n8597), .A(n9396), .ZN(n8583) );
  INV_X1 U9856 ( .A(n8654), .ZN(n8644) );
  AOI21_X1 U9857 ( .B1(n8584), .B2(n8583), .A(n8644), .ZN(n8585) );
  MUX2_X1 U9858 ( .A(n8656), .B(n8654), .S(n8591), .Z(n8588) );
  MUX2_X1 U9859 ( .A(n8638), .B(n8658), .S(n8591), .Z(n8589) );
  NAND2_X1 U9860 ( .A1(n9338), .A2(n6490), .ZN(n8594) );
  NAND2_X1 U9861 ( .A1(n6405), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n8593) );
  NAND2_X1 U9862 ( .A1(n9955), .A2(n9498), .ZN(n8667) );
  OAI211_X1 U9863 ( .C1(n5398), .C2(n6738), .A(n8635), .B(n8598), .ZN(n8600)
         );
  OAI21_X1 U9864 ( .B1(n8601), .B2(n8600), .A(n8599), .ZN(n8734) );
  NAND2_X1 U9865 ( .A1(n8602), .A2(n8739), .ZN(n8636) );
  INV_X1 U9866 ( .A(n8603), .ZN(n8672) );
  NAND2_X1 U9867 ( .A1(n8672), .A2(n8667), .ZN(n8728) );
  NOR2_X1 U9868 ( .A1(n9955), .A2(n9498), .ZN(n8664) );
  NOR2_X1 U9869 ( .A1(n6895), .A2(n8606), .ZN(n8682) );
  OR2_X1 U9870 ( .A1(n8607), .A2(n8682), .ZN(n10516) );
  NOR4_X1 U9871 ( .A1(n10516), .A2(n6741), .A3(n10540), .A4(n8635), .ZN(n8611)
         );
  NAND4_X1 U9872 ( .A1(n8611), .A2(n8610), .A3(n8609), .A4(n8608), .ZN(n8615)
         );
  NOR4_X1 U9873 ( .A1(n8619), .A2(n8618), .A3(n8617), .A4(n8616), .ZN(n8620)
         );
  NAND4_X1 U9874 ( .A1(n8623), .A2(n8622), .A3(n8621), .A4(n8620), .ZN(n8624)
         );
  NOR4_X1 U9875 ( .A1(n9757), .A2(n9780), .A3(n9792), .A4(n8627), .ZN(n8628)
         );
  NAND4_X1 U9876 ( .A1(n9703), .A2(n9724), .A3(n9747), .A4(n8628), .ZN(n8629)
         );
  NOR4_X1 U9877 ( .A1(n6678), .A2(n8630), .A3(n9667), .A4(n8629), .ZN(n8631)
         );
  NAND4_X1 U9878 ( .A1(n6814), .A2(n8632), .A3(n9636), .A4(n8631), .ZN(n8633)
         );
  AOI21_X1 U9879 ( .B1(n8636), .B2(n8635), .A(n8675), .ZN(n8637) );
  NAND2_X1 U9880 ( .A1(n8639), .A2(n8638), .ZN(n8661) );
  INV_X1 U9881 ( .A(n8640), .ZN(n8641) );
  NAND4_X1 U9882 ( .A1(n8653), .A2(n8642), .A3(n8641), .A4(n8649), .ZN(n8643)
         );
  NOR3_X1 U9883 ( .A1(n8661), .A2(n8644), .A3(n8643), .ZN(n8725) );
  INV_X1 U9884 ( .A(n8645), .ZN(n8646) );
  AOI21_X1 U9885 ( .B1(n8648), .B2(n8647), .A(n8646), .ZN(n8652) );
  INV_X1 U9886 ( .A(n8649), .ZN(n8651) );
  OAI21_X1 U9887 ( .B1(n8652), .B2(n8651), .A(n8650), .ZN(n8655) );
  NAND3_X1 U9888 ( .A1(n8655), .A2(n8654), .A3(n8653), .ZN(n8657) );
  AND3_X1 U9889 ( .A1(n8658), .A2(n8657), .A3(n8656), .ZN(n8662) );
  OAI211_X1 U9890 ( .C1(n8662), .C2(n8661), .A(n8660), .B(n8659), .ZN(n8723)
         );
  AOI21_X1 U9891 ( .B1(n8725), .B2(n8663), .A(n8723), .ZN(n8669) );
  INV_X1 U9892 ( .A(n8664), .ZN(n8666) );
  NAND2_X1 U9893 ( .A1(n8666), .A2(n8665), .ZN(n8726) );
  OAI22_X1 U9894 ( .A1(n8669), .A2(n8726), .B1(n8668), .B2(n8667), .ZN(n8670)
         );
  OAI211_X1 U9895 ( .C1(n9955), .C2(n9616), .A(n8670), .B(n5398), .ZN(n8674)
         );
  INV_X1 U9896 ( .A(n8671), .ZN(n8673) );
  NAND3_X1 U9897 ( .A1(n8674), .A2(n8673), .A3(n8672), .ZN(n8677) );
  INV_X1 U9898 ( .A(n8675), .ZN(n8676) );
  NAND2_X1 U9899 ( .A1(n8677), .A2(n8676), .ZN(n8678) );
  INV_X1 U9900 ( .A(n8680), .ZN(n10517) );
  INV_X1 U9901 ( .A(n8681), .ZN(n8689) );
  INV_X1 U9902 ( .A(n8682), .ZN(n8685) );
  AND4_X1 U9903 ( .A1(n8685), .A2(n8635), .A3(n8684), .A4(n8683), .ZN(n8688)
         );
  INV_X1 U9904 ( .A(n8686), .ZN(n8687) );
  OAI21_X1 U9905 ( .B1(n8689), .B2(n8688), .A(n8687), .ZN(n8693) );
  INV_X1 U9906 ( .A(n8690), .ZN(n8692) );
  AOI21_X1 U9907 ( .B1(n8693), .B2(n8692), .A(n8691), .ZN(n8696) );
  OAI21_X1 U9908 ( .B1(n8696), .B2(n8695), .A(n8694), .ZN(n8699) );
  AOI21_X1 U9909 ( .B1(n8699), .B2(n8698), .A(n8697), .ZN(n8703) );
  OAI211_X1 U9910 ( .C1(n8703), .C2(n8702), .A(n8701), .B(n8700), .ZN(n8706)
         );
  NAND3_X1 U9911 ( .A1(n8706), .A2(n8705), .A3(n8704), .ZN(n8709) );
  NAND3_X1 U9912 ( .A1(n8709), .A2(n8708), .A3(n8707), .ZN(n8710) );
  NAND3_X1 U9913 ( .A1(n8712), .A2(n8711), .A3(n8710), .ZN(n8717) );
  NAND2_X1 U9914 ( .A1(n8714), .A2(n8713), .ZN(n8715) );
  NAND4_X1 U9915 ( .A1(n8718), .A2(n8717), .A3(n8716), .A4(n8715), .ZN(n8720)
         );
  AOI21_X1 U9916 ( .B1(n5004), .B2(n8720), .A(n8719), .ZN(n8722) );
  OAI211_X1 U9917 ( .C1(n5136), .C2(n8722), .A(n8721), .B(n5003), .ZN(n8724)
         );
  AOI21_X1 U9918 ( .B1(n8725), .B2(n8724), .A(n8723), .ZN(n8727) );
  NOR2_X1 U9919 ( .A1(n8727), .A2(n8726), .ZN(n8729) );
  OAI21_X1 U9920 ( .B1(n8729), .B2(n8728), .A(n5398), .ZN(n8732) );
  NOR2_X1 U9921 ( .A1(n8732), .A2(n8730), .ZN(n8731) );
  AOI211_X1 U9922 ( .C1(n10517), .C2(n8732), .A(n8738), .B(n8731), .ZN(n8733)
         );
  NAND2_X1 U9923 ( .A1(n8736), .A2(n8735), .ZN(n8737) );
  OAI211_X1 U9924 ( .C1(n8739), .C2(n8738), .A(n8737), .B(P1_B_REG_SCAN_IN), 
        .ZN(n8740) );
  NAND2_X1 U9925 ( .A1(n8742), .A2(n8741), .ZN(n8750) );
  OAI22_X1 U9926 ( .A1(n9628), .A2(n6936), .B1(n9640), .B2(n8744), .ZN(n8748)
         );
  OAI22_X1 U9927 ( .A1(n9628), .A2(n8744), .B1(n9640), .B2(n8743), .ZN(n8746)
         );
  XNOR2_X1 U9928 ( .A(n8746), .B(n8745), .ZN(n8747) );
  XOR2_X1 U9929 ( .A(n8748), .B(n8747), .Z(n8749) );
  XNOR2_X1 U9930 ( .A(n8750), .B(n8749), .ZN(n8757) );
  AOI22_X1 U9931 ( .A1(n9626), .A2(n9486), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n8752) );
  NAND2_X1 U9932 ( .A1(n9656), .A2(n9451), .ZN(n8751) );
  OAI211_X1 U9933 ( .C1(n8753), .C2(n9434), .A(n8752), .B(n8751), .ZN(n8754)
         );
  AOI21_X1 U9934 ( .B1(n8755), .B2(n9494), .A(n8754), .ZN(n8756) );
  OAI21_X1 U9935 ( .B1(n8757), .B2(n9496), .A(n8756), .ZN(P1_U3220) );
  AND2_X1 U9936 ( .A1(n8759), .A2(n8758), .ZN(n8760) );
  XNOR2_X1 U9937 ( .A(n10725), .B(n8796), .ZN(n8762) );
  XNOR2_X1 U9938 ( .A(n8762), .B(n8933), .ZN(n8916) );
  NAND2_X1 U9939 ( .A1(n8915), .A2(n8763), .ZN(n8851) );
  XNOR2_X1 U9940 ( .A(n8848), .B(n8796), .ZN(n8764) );
  XNOR2_X1 U9941 ( .A(n8764), .B(n9217), .ZN(n8850) );
  XNOR2_X1 U9942 ( .A(n10741), .B(n8796), .ZN(n8766) );
  XNOR2_X1 U9943 ( .A(n8766), .B(n8932), .ZN(n8857) );
  INV_X1 U9944 ( .A(n8766), .ZN(n8767) );
  INV_X1 U9945 ( .A(n8891), .ZN(n8769) );
  XNOR2_X1 U9946 ( .A(n10752), .B(n8796), .ZN(n8770) );
  XNOR2_X1 U9947 ( .A(n8770), .B(n10739), .ZN(n8890) );
  INV_X1 U9948 ( .A(n8890), .ZN(n8768) );
  NAND2_X1 U9949 ( .A1(n8769), .A2(n8768), .ZN(n8892) );
  NAND2_X1 U9950 ( .A1(n8892), .A2(n8771), .ZN(n8822) );
  XNOR2_X1 U9951 ( .A(n9159), .B(n7984), .ZN(n8821) );
  INV_X1 U9952 ( .A(n8821), .ZN(n8772) );
  NAND2_X1 U9953 ( .A1(n8772), .A2(n8931), .ZN(n8773) );
  XNOR2_X1 U9954 ( .A(n9331), .B(n8796), .ZN(n8775) );
  XNOR2_X1 U9955 ( .A(n8775), .B(n8825), .ZN(n8877) );
  INV_X1 U9956 ( .A(n8877), .ZN(n8774) );
  NAND2_X1 U9957 ( .A1(n8775), .A2(n8825), .ZN(n8776) );
  NAND2_X1 U9958 ( .A1(n8874), .A2(n8776), .ZN(n8830) );
  XNOR2_X1 U9959 ( .A(n9328), .B(n8796), .ZN(n8777) );
  XNOR2_X1 U9960 ( .A(n8777), .B(n9148), .ZN(n8831) );
  INV_X1 U9961 ( .A(n8777), .ZN(n8778) );
  XNOR2_X1 U9962 ( .A(n8779), .B(n8796), .ZN(n8780) );
  XNOR2_X1 U9963 ( .A(n8780), .B(n9130), .ZN(n8884) );
  NAND2_X1 U9964 ( .A1(n8885), .A2(n8884), .ZN(n8883) );
  INV_X1 U9965 ( .A(n8780), .ZN(n8781) );
  NAND2_X1 U9966 ( .A1(n8781), .A2(n9130), .ZN(n8782) );
  NAND2_X1 U9967 ( .A1(n8883), .A2(n8782), .ZN(n8783) );
  XNOR2_X1 U9968 ( .A(n9273), .B(n8796), .ZN(n8784) );
  XNOR2_X1 U9969 ( .A(n8783), .B(n8784), .ZN(n8813) );
  NAND2_X1 U9970 ( .A1(n8813), .A2(n9114), .ZN(n8787) );
  INV_X1 U9971 ( .A(n8783), .ZN(n8785) );
  NAND2_X1 U9972 ( .A1(n8785), .A2(n8784), .ZN(n8786) );
  NAND2_X1 U9973 ( .A1(n8787), .A2(n8786), .ZN(n8865) );
  XNOR2_X1 U9974 ( .A(n9093), .B(n8796), .ZN(n8788) );
  XNOR2_X1 U9975 ( .A(n8788), .B(n9102), .ZN(n8866) );
  NAND2_X1 U9976 ( .A1(n8865), .A2(n8866), .ZN(n8839) );
  NAND2_X1 U9977 ( .A1(n8788), .A2(n9076), .ZN(n8840) );
  XNOR2_X1 U9978 ( .A(n9078), .B(n8796), .ZN(n8790) );
  NAND2_X1 U9979 ( .A1(n8790), .A2(n8868), .ZN(n8789) );
  AND2_X1 U9980 ( .A1(n8840), .A2(n8789), .ZN(n8792) );
  INV_X1 U9981 ( .A(n8789), .ZN(n8791) );
  XNOR2_X1 U9982 ( .A(n8790), .B(n9090), .ZN(n8842) );
  XNOR2_X1 U9983 ( .A(n9260), .B(n7984), .ZN(n8793) );
  NAND2_X1 U9984 ( .A1(n8793), .A2(n8929), .ZN(n8904) );
  INV_X1 U9985 ( .A(n8793), .ZN(n8794) );
  NAND2_X1 U9986 ( .A1(n8794), .A2(n9077), .ZN(n8905) );
  XNOR2_X1 U9987 ( .A(n9057), .B(n8796), .ZN(n8795) );
  XNOR2_X1 U9988 ( .A(n8795), .B(n9064), .ZN(n8806) );
  XNOR2_X1 U9989 ( .A(n8797), .B(n8796), .ZN(n8798) );
  XNOR2_X1 U9990 ( .A(n8799), .B(n8798), .ZN(n8804) );
  NOR2_X1 U9991 ( .A1(n8919), .A2(n9041), .ZN(n8802) );
  AOI22_X1 U9992 ( .A1(n8922), .A2(n9259), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n8800) );
  OAI21_X1 U9993 ( .B1(n9040), .B2(n8918), .A(n8800), .ZN(n8801) );
  AOI211_X1 U9994 ( .C1(n9045), .C2(n8910), .A(n8802), .B(n8801), .ZN(n8803)
         );
  OAI21_X1 U9995 ( .B1(n8804), .B2(n8912), .A(n8803), .ZN(P2_U3160) );
  XNOR2_X1 U9996 ( .A(n8805), .B(n8806), .ZN(n8812) );
  OAI22_X1 U9997 ( .A1(n8918), .A2(n9053), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8807), .ZN(n8808) );
  AOI21_X1 U9998 ( .B1(n8922), .B2(n8929), .A(n8808), .ZN(n8809) );
  OAI21_X1 U9999 ( .B1(n9054), .B2(n8919), .A(n8809), .ZN(n8810) );
  AOI21_X1 U10000 ( .B1(n9057), .B2(n8910), .A(n8810), .ZN(n8811) );
  OAI21_X1 U10001 ( .B1(n8812), .B2(n8912), .A(n8811), .ZN(P2_U3154) );
  XNOR2_X1 U10002 ( .A(n8813), .B(n9089), .ZN(n8819) );
  OAI22_X1 U10003 ( .A1(n8918), .A2(n9076), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8814), .ZN(n8815) );
  AOI21_X1 U10004 ( .B1(n8922), .B2(n9130), .A(n8815), .ZN(n8816) );
  OAI21_X1 U10005 ( .B1(n9107), .B2(n8919), .A(n8816), .ZN(n8817) );
  AOI21_X1 U10006 ( .B1(n9273), .B2(n8910), .A(n8817), .ZN(n8818) );
  OAI21_X1 U10007 ( .B1(n8819), .B2(n8912), .A(n8818), .ZN(P2_U3156) );
  INV_X1 U10008 ( .A(n9296), .ZN(n8829) );
  OAI211_X1 U10009 ( .C1(n8822), .C2(n8821), .A(n8820), .B(n8914), .ZN(n8828)
         );
  NAND2_X1 U10010 ( .A1(n9194), .A2(n8922), .ZN(n8824) );
  OAI211_X1 U10011 ( .C1(n8825), .C2(n8918), .A(n8824), .B(n8823), .ZN(n8826)
         );
  AOI21_X1 U10012 ( .B1(n8899), .B2(n9165), .A(n8826), .ZN(n8827) );
  OAI211_X1 U10013 ( .C1(n8829), .C2(n8925), .A(n8828), .B(n8827), .ZN(
        P2_U3159) );
  XOR2_X1 U10014 ( .A(n8831), .B(n8830), .Z(n8838) );
  INV_X1 U10015 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n8832) );
  OAI22_X1 U10016 ( .A1(n8918), .A2(n8833), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8832), .ZN(n8834) );
  AOI21_X1 U10017 ( .B1(n8922), .B2(n9295), .A(n8834), .ZN(n8835) );
  OAI21_X1 U10018 ( .B1(n9132), .B2(n8919), .A(n8835), .ZN(n8836) );
  AOI21_X1 U10019 ( .B1(n9138), .B2(n8910), .A(n8836), .ZN(n8837) );
  OAI21_X1 U10020 ( .B1(n8838), .B2(n8912), .A(n8837), .ZN(P2_U3163) );
  NAND2_X1 U10021 ( .A1(n8839), .A2(n8840), .ZN(n8841) );
  XOR2_X1 U10022 ( .A(n8842), .B(n8841), .Z(n8847) );
  OAI22_X1 U10023 ( .A1(n8918), .A2(n9077), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10184), .ZN(n8843) );
  AOI21_X1 U10024 ( .B1(n8922), .B2(n9102), .A(n8843), .ZN(n8844) );
  OAI21_X1 U10025 ( .B1(n9082), .B2(n8919), .A(n8844), .ZN(n8845) );
  AOI21_X1 U10026 ( .B1(n9078), .B2(n8910), .A(n8845), .ZN(n8846) );
  OAI21_X1 U10027 ( .B1(n8847), .B2(n8912), .A(n8846), .ZN(P2_U3165) );
  INV_X1 U10028 ( .A(n8848), .ZN(n10732) );
  OAI211_X1 U10029 ( .C1(n8851), .C2(n8850), .A(n8849), .B(n8914), .ZN(n8855)
         );
  NOR2_X1 U10030 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10090), .ZN(n8999) );
  AOI21_X1 U10031 ( .B1(n8932), .B2(n8895), .A(n8999), .ZN(n8852) );
  OAI21_X1 U10032 ( .B1(n9237), .B2(n8897), .A(n8852), .ZN(n8853) );
  AOI21_X1 U10033 ( .B1(n9204), .B2(n8899), .A(n8853), .ZN(n8854) );
  OAI211_X1 U10034 ( .C1(n10732), .C2(n8925), .A(n8855), .B(n8854), .ZN(
        P2_U3166) );
  AOI21_X1 U10035 ( .B1(n8857), .B2(n8856), .A(n5008), .ZN(n8864) );
  INV_X1 U10036 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8858) );
  OAI22_X1 U10037 ( .A1(n10739), .A2(n8918), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8858), .ZN(n8859) );
  AOI21_X1 U10038 ( .B1(n8922), .B2(n9217), .A(n8859), .ZN(n8860) );
  OAI21_X1 U10039 ( .B1(n9191), .B2(n8919), .A(n8860), .ZN(n8861) );
  AOI21_X1 U10040 ( .B1(n8862), .B2(n8910), .A(n8861), .ZN(n8863) );
  OAI21_X1 U10041 ( .B1(n8864), .B2(n8912), .A(n8863), .ZN(P2_U3168) );
  XOR2_X1 U10042 ( .A(n8866), .B(n8865), .Z(n8873) );
  OAI22_X1 U10043 ( .A1(n8918), .A2(n8868), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8867), .ZN(n8869) );
  AOI21_X1 U10044 ( .B1(n8922), .B2(n9089), .A(n8869), .ZN(n8870) );
  OAI21_X1 U10045 ( .B1(n9094), .B2(n8919), .A(n8870), .ZN(n8871) );
  AOI21_X1 U10046 ( .B1(n9093), .B2(n8910), .A(n8871), .ZN(n8872) );
  OAI21_X1 U10047 ( .B1(n8873), .B2(n8912), .A(n8872), .ZN(P2_U3169) );
  INV_X1 U10048 ( .A(n8874), .ZN(n8875) );
  AOI21_X1 U10049 ( .B1(n8877), .B2(n8876), .A(n8875), .ZN(n8882) );
  OAI22_X1 U10050 ( .A1(n8918), .A2(n9148), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10203), .ZN(n8878) );
  AOI21_X1 U10051 ( .B1(n8922), .B2(n8931), .A(n8878), .ZN(n8879) );
  OAI21_X1 U10052 ( .B1(n9151), .B2(n8919), .A(n8879), .ZN(n8880) );
  AOI21_X1 U10053 ( .B1(n9331), .B2(n8910), .A(n8880), .ZN(n8881) );
  OAI21_X1 U10054 ( .B1(n8882), .B2(n8912), .A(n8881), .ZN(P2_U3173) );
  OAI211_X1 U10055 ( .C1(n8885), .C2(n8884), .A(n8883), .B(n8914), .ZN(n8889)
         );
  OAI22_X1 U10056 ( .A1(n8897), .A2(n9148), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10205), .ZN(n8887) );
  NOR2_X1 U10057 ( .A1(n8919), .A2(n9119), .ZN(n8886) );
  AOI211_X1 U10058 ( .C1(n8895), .C2(n9089), .A(n8887), .B(n8886), .ZN(n8888)
         );
  OAI211_X1 U10059 ( .C1(n9323), .C2(n8925), .A(n8889), .B(n8888), .ZN(
        P2_U3175) );
  INV_X1 U10060 ( .A(n10752), .ZN(n8902) );
  AOI21_X1 U10061 ( .B1(n8891), .B2(n8890), .A(n8912), .ZN(n8893) );
  NAND2_X1 U10062 ( .A1(n8893), .A2(n8892), .ZN(n8901) );
  NOR2_X1 U10063 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8894), .ZN(n10497) );
  AOI21_X1 U10064 ( .B1(n8931), .B2(n8895), .A(n10497), .ZN(n8896) );
  OAI21_X1 U10065 ( .B1(n9201), .B2(n8897), .A(n8896), .ZN(n8898) );
  AOI21_X1 U10066 ( .B1(n9176), .B2(n8899), .A(n8898), .ZN(n8900) );
  OAI211_X1 U10067 ( .C1(n8902), .C2(n8925), .A(n8901), .B(n8900), .ZN(
        P2_U3178) );
  NAND2_X1 U10068 ( .A1(n8905), .A2(n8904), .ZN(n8906) );
  XNOR2_X1 U10069 ( .A(n8903), .B(n8906), .ZN(n8913) );
  NOR2_X1 U10070 ( .A1(n8919), .A2(n9065), .ZN(n8909) );
  AOI22_X1 U10071 ( .A1(n8922), .A2(n9090), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n8907) );
  OAI21_X1 U10072 ( .B1(n9064), .B2(n8918), .A(n8907), .ZN(n8908) );
  AOI211_X1 U10073 ( .C1(n9260), .C2(n8910), .A(n8909), .B(n8908), .ZN(n8911)
         );
  OAI21_X1 U10074 ( .B1(n8913), .B2(n8912), .A(n8911), .ZN(P2_U3180) );
  INV_X1 U10075 ( .A(n10725), .ZN(n9226) );
  OAI211_X1 U10076 ( .C1(n5010), .C2(n8916), .A(n8915), .B(n8914), .ZN(n8924)
         );
  INV_X1 U10077 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n10212) );
  OR2_X1 U10078 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10212), .ZN(n8987) );
  OAI21_X1 U10079 ( .B1(n8918), .B2(n8917), .A(n8987), .ZN(n8921) );
  NOR2_X1 U10080 ( .A1(n8919), .A2(n9220), .ZN(n8920) );
  AOI211_X1 U10081 ( .C1(n8922), .C2(n9215), .A(n8921), .B(n8920), .ZN(n8923)
         );
  OAI211_X1 U10082 ( .C1(n9226), .C2(n8925), .A(n8924), .B(n8923), .ZN(
        P2_U3181) );
  MUX2_X1 U10083 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n8926), .S(P2_U3893), .Z(
        P2_U3522) );
  MUX2_X1 U10084 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8927), .S(P2_U3893), .Z(
        P2_U3521) );
  MUX2_X1 U10085 ( .A(n8928), .B(P2_DATAO_REG_28__SCAN_IN), .S(n10508), .Z(
        P2_U3519) );
  MUX2_X1 U10086 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n9259), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U10087 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n8929), .S(P2_U3893), .Z(
        P2_U3517) );
  MUX2_X1 U10088 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n9102), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U10089 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n9089), .S(P2_U3893), .Z(
        P2_U3514) );
  MUX2_X1 U10090 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n9130), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U10091 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8930), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U10092 ( .A(n9295), .B(P2_DATAO_REG_20__SCAN_IN), .S(n10508), .Z(
        P2_U3511) );
  MUX2_X1 U10093 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8931), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U10094 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n9194), .S(P2_U3893), .Z(
        P2_U3509) );
  MUX2_X1 U10095 ( .A(n8932), .B(P2_DATAO_REG_17__SCAN_IN), .S(n10508), .Z(
        P2_U3508) );
  MUX2_X1 U10096 ( .A(n9217), .B(P2_DATAO_REG_16__SCAN_IN), .S(n10508), .Z(
        P2_U3507) );
  MUX2_X1 U10097 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8933), .S(P2_U3893), .Z(
        P2_U3506) );
  MUX2_X1 U10098 ( .A(n9215), .B(P2_DATAO_REG_14__SCAN_IN), .S(n10508), .Z(
        P2_U3505) );
  MUX2_X1 U10099 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n8934), .S(P2_U3893), .Z(
        P2_U3504) );
  MUX2_X1 U10100 ( .A(n8935), .B(P2_DATAO_REG_12__SCAN_IN), .S(n10508), .Z(
        P2_U3503) );
  MUX2_X1 U10101 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n10657), .S(P2_U3893), .Z(
        P2_U3501) );
  MUX2_X1 U10102 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n8936), .S(P2_U3893), .Z(
        P2_U3498) );
  MUX2_X1 U10103 ( .A(n8937), .B(P2_DATAO_REG_6__SCAN_IN), .S(n10508), .Z(
        P2_U3497) );
  MUX2_X1 U10104 ( .A(n8938), .B(P2_DATAO_REG_5__SCAN_IN), .S(n10508), .Z(
        P2_U3496) );
  MUX2_X1 U10105 ( .A(n8939), .B(P2_DATAO_REG_4__SCAN_IN), .S(n10508), .Z(
        P2_U3495) );
  MUX2_X1 U10106 ( .A(n8940), .B(P2_DATAO_REG_3__SCAN_IN), .S(n10508), .Z(
        P2_U3494) );
  MUX2_X1 U10107 ( .A(n8941), .B(P2_DATAO_REG_2__SCAN_IN), .S(n10508), .Z(
        P2_U3493) );
  MUX2_X1 U10108 ( .A(n8942), .B(P2_DATAO_REG_1__SCAN_IN), .S(n10508), .Z(
        P2_U3492) );
  MUX2_X1 U10109 ( .A(n6249), .B(P2_DATAO_REG_0__SCAN_IN), .S(n10508), .Z(
        P2_U3491) );
  AOI21_X1 U10110 ( .B1(n8945), .B2(n8944), .A(n8943), .ZN(n8960) );
  INV_X1 U10111 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n8952) );
  OAI21_X1 U10112 ( .B1(n8948), .B2(n8947), .A(n8946), .ZN(n8949) );
  NAND2_X1 U10113 ( .A1(n8949), .A2(n10495), .ZN(n8950) );
  OAI211_X1 U10114 ( .C1(n10489), .C2(n8952), .A(n8951), .B(n8950), .ZN(n8957)
         );
  AOI21_X1 U10115 ( .B1(n10715), .B2(n8954), .A(n8953), .ZN(n8955) );
  NOR2_X1 U10116 ( .A1(n8955), .A2(n10501), .ZN(n8956) );
  AOI211_X1 U10117 ( .C1(n10474), .C2(n8958), .A(n8957), .B(n8956), .ZN(n8959)
         );
  OAI21_X1 U10118 ( .B1(n8960), .B2(n10506), .A(n8959), .ZN(P2_U3195) );
  AOI21_X1 U10119 ( .B1(n5005), .B2(n8962), .A(n8961), .ZN(n8978) );
  INV_X1 U10120 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n8969) );
  OAI21_X1 U10121 ( .B1(n8965), .B2(n8964), .A(n8963), .ZN(n8966) );
  NAND2_X1 U10122 ( .A1(n8966), .A2(n10495), .ZN(n8967) );
  OAI211_X1 U10123 ( .C1(n10489), .C2(n8969), .A(n8968), .B(n8967), .ZN(n8975)
         );
  AOI21_X1 U10124 ( .B1(n8972), .B2(n8971), .A(n8970), .ZN(n8973) );
  NOR2_X1 U10125 ( .A1(n8973), .A2(n10501), .ZN(n8974) );
  AOI211_X1 U10126 ( .C1(n10474), .C2(n8976), .A(n8975), .B(n8974), .ZN(n8977)
         );
  OAI21_X1 U10127 ( .B1(n8978), .B2(n10506), .A(n8977), .ZN(P2_U3196) );
  AOI21_X1 U10128 ( .B1(n8981), .B2(n8980), .A(n8979), .ZN(n8996) );
  INV_X1 U10129 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n8988) );
  OAI21_X1 U10130 ( .B1(n8984), .B2(n8983), .A(n8982), .ZN(n8985) );
  NAND2_X1 U10131 ( .A1(n8985), .A2(n10495), .ZN(n8986) );
  OAI211_X1 U10132 ( .C1(n10489), .C2(n8988), .A(n8987), .B(n8986), .ZN(n8993)
         );
  AOI21_X1 U10133 ( .B1(n10729), .B2(n8990), .A(n8989), .ZN(n8991) );
  NOR2_X1 U10134 ( .A1(n8991), .A2(n10501), .ZN(n8992) );
  AOI211_X1 U10135 ( .C1(n10474), .C2(n8994), .A(n8993), .B(n8992), .ZN(n8995)
         );
  OAI21_X1 U10136 ( .B1(n8996), .B2(n10506), .A(n8995), .ZN(P2_U3197) );
  AOI21_X1 U10137 ( .B1(n4962), .B2(n8998), .A(n8997), .ZN(n9014) );
  INV_X1 U10138 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n9006) );
  INV_X1 U10139 ( .A(n8999), .ZN(n9005) );
  OAI21_X1 U10140 ( .B1(n9002), .B2(n9001), .A(n9000), .ZN(n9003) );
  NAND2_X1 U10141 ( .A1(n9003), .A2(n10495), .ZN(n9004) );
  OAI211_X1 U10142 ( .C1(n10489), .C2(n9006), .A(n9005), .B(n9004), .ZN(n9011)
         );
  AOI21_X1 U10143 ( .B1(n4963), .B2(n9008), .A(n9007), .ZN(n9009) );
  NOR2_X1 U10144 ( .A1(n9009), .A2(n10501), .ZN(n9010) );
  AOI211_X1 U10145 ( .C1(n10474), .C2(n9012), .A(n9011), .B(n9010), .ZN(n9013)
         );
  OAI21_X1 U10146 ( .B1(n9014), .B2(n10506), .A(n9013), .ZN(P2_U3198) );
  AOI21_X1 U10147 ( .B1(n10746), .B2(n9016), .A(n9015), .ZN(n9029) );
  AOI21_X1 U10148 ( .B1(n9018), .B2(n9192), .A(n9017), .ZN(n9019) );
  NOR2_X1 U10149 ( .A1(n10506), .A2(n9019), .ZN(n9022) );
  INV_X1 U10150 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n9020) );
  OAI22_X1 U10151 ( .A1(n10489), .A2(n9020), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8858), .ZN(n9021) );
  XNOR2_X1 U10152 ( .A(n9025), .B(n9024), .ZN(n9026) );
  NAND2_X1 U10153 ( .A1(n9026), .A2(n10495), .ZN(n9027) );
  OAI211_X1 U10154 ( .C1(n9029), .C2(n10501), .A(n9028), .B(n9027), .ZN(
        P2_U3199) );
  INV_X1 U10155 ( .A(n9031), .ZN(n9032) );
  NOR2_X1 U10156 ( .A1(n9033), .A2(n9032), .ZN(n9300) );
  NOR3_X1 U10157 ( .A1(n9300), .A2(n9223), .A3(n9034), .ZN(n9037) );
  NOR2_X1 U10158 ( .A1(n10643), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n9035) );
  OAI22_X1 U10159 ( .A1(n9302), .A2(n9225), .B1(n9037), .B2(n9035), .ZN(
        P2_U3202) );
  NOR2_X1 U10160 ( .A1(n10643), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n9036) );
  OAI22_X1 U10161 ( .A1(n9305), .A2(n9225), .B1(n9037), .B2(n9036), .ZN(
        P2_U3203) );
  INV_X1 U10162 ( .A(n9038), .ZN(n9048) );
  NAND2_X1 U10163 ( .A1(n9039), .A2(n10647), .ZN(n9047) );
  NOR2_X1 U10164 ( .A1(n9178), .A2(n9040), .ZN(n9044) );
  OAI22_X1 U10165 ( .A1(n10643), .A2(n9042), .B1(n9041), .B2(n9238), .ZN(n9043) );
  AOI211_X1 U10166 ( .C1(n9045), .C2(n10641), .A(n9044), .B(n9043), .ZN(n9046)
         );
  OAI211_X1 U10167 ( .C1(n9048), .C2(n9230), .A(n9047), .B(n9046), .ZN(
        P2_U3205) );
  XNOR2_X1 U10168 ( .A(n9049), .B(n9050), .ZN(n9256) );
  INV_X1 U10169 ( .A(n9256), .ZN(n9060) );
  NAND2_X1 U10170 ( .A1(n9255), .A2(n10647), .ZN(n9059) );
  OAI22_X1 U10171 ( .A1(n10643), .A2(n9055), .B1(n9054), .B2(n9238), .ZN(n9056) );
  AOI21_X1 U10172 ( .B1(n9057), .B2(n10641), .A(n9056), .ZN(n9058) );
  OAI211_X1 U10173 ( .C1(n9060), .C2(n9230), .A(n9059), .B(n9058), .ZN(
        P2_U3206) );
  XNOR2_X1 U10174 ( .A(n9061), .B(n9062), .ZN(n9063) );
  AOI22_X1 U10175 ( .A1(n9063), .A2(n9211), .B1(n9216), .B2(n9090), .ZN(n9264)
         );
  NOR2_X1 U10176 ( .A1(n9178), .A2(n9064), .ZN(n9068) );
  OAI22_X1 U10177 ( .A1(n10647), .A2(n9066), .B1(n9065), .B2(n9238), .ZN(n9067) );
  AOI211_X1 U10178 ( .C1(n9260), .C2(n10641), .A(n9068), .B(n9067), .ZN(n9073)
         );
  OR2_X1 U10179 ( .A1(n9070), .A2(n9069), .ZN(n9261) );
  NAND3_X1 U10180 ( .A1(n9261), .A2(n9071), .A3(n10639), .ZN(n9072) );
  OAI211_X1 U10181 ( .C1(n9264), .C2(n9223), .A(n9073), .B(n9072), .ZN(
        P2_U3207) );
  INV_X1 U10182 ( .A(n9240), .ZN(n9079) );
  XOR2_X1 U10183 ( .A(n9074), .B(n9080), .Z(n9075) );
  OAI222_X1 U10184 ( .A1(n10754), .A2(n9077), .B1(n9236), .B2(n9076), .C1(
        n9234), .C2(n9075), .ZN(n9265) );
  AOI21_X1 U10185 ( .B1(n9079), .B2(n9078), .A(n9265), .ZN(n9086) );
  XOR2_X1 U10186 ( .A(n9081), .B(n9080), .Z(n9266) );
  OAI22_X1 U10187 ( .A1(n10643), .A2(n9083), .B1(n9082), .B2(n9238), .ZN(n9084) );
  AOI21_X1 U10188 ( .B1(n9266), .B2(n10639), .A(n9084), .ZN(n9085) );
  OAI21_X1 U10189 ( .B1(n9086), .B2(n9223), .A(n9085), .ZN(P2_U3208) );
  OAI21_X1 U10190 ( .B1(n9088), .B2(n9096), .A(n9087), .ZN(n9091) );
  AOI222_X1 U10191 ( .A1(n9211), .A2(n9091), .B1(n9090), .B2(n10658), .C1(
        n9089), .C2(n9216), .ZN(n9092) );
  INV_X1 U10192 ( .A(n9092), .ZN(n9269) );
  INV_X1 U10193 ( .A(n9093), .ZN(n9318) );
  OAI22_X1 U10194 ( .A1(n9318), .A2(n9240), .B1(n9094), .B2(n9238), .ZN(n9095)
         );
  OAI21_X1 U10195 ( .B1(n9269), .B2(n9095), .A(n10647), .ZN(n9100) );
  AND2_X1 U10196 ( .A1(n4992), .A2(n9096), .ZN(n9097) );
  NOR2_X1 U10197 ( .A1(n9098), .A2(n9097), .ZN(n9270) );
  AOI22_X1 U10198 ( .A1(n9270), .A2(n10639), .B1(P2_REG2_REG_24__SCAN_IN), 
        .B2(n9223), .ZN(n9099) );
  NAND2_X1 U10199 ( .A1(n9100), .A2(n9099), .ZN(P2_U3209) );
  XNOR2_X1 U10200 ( .A(n9101), .B(n9104), .ZN(n9103) );
  AOI222_X1 U10201 ( .A1(n9211), .A2(n9103), .B1(n9130), .B2(n9216), .C1(n9102), .C2(n10658), .ZN(n9276) );
  XNOR2_X1 U10202 ( .A(n9105), .B(n9104), .ZN(n9274) );
  NOR2_X1 U10203 ( .A1(n9106), .A2(n9225), .ZN(n9110) );
  OAI22_X1 U10204 ( .A1(n10643), .A2(n9108), .B1(n9107), .B2(n9238), .ZN(n9109) );
  AOI211_X1 U10205 ( .C1(n9274), .C2(n10639), .A(n9110), .B(n9109), .ZN(n9111)
         );
  OAI21_X1 U10206 ( .B1(n9276), .B2(n9223), .A(n9111), .ZN(P2_U3210) );
  XOR2_X1 U10207 ( .A(n9112), .B(n9117), .Z(n9113) );
  OAI222_X1 U10208 ( .A1(n9236), .A2(n9148), .B1(n10754), .B2(n9114), .C1(
        n9113), .C2(n9234), .ZN(n9277) );
  INV_X1 U10209 ( .A(n9277), .ZN(n9124) );
  NAND2_X1 U10210 ( .A1(n9284), .A2(n9116), .ZN(n9118) );
  XNOR2_X1 U10211 ( .A(n9118), .B(n9117), .ZN(n9278) );
  NOR2_X1 U10212 ( .A1(n9323), .A2(n9225), .ZN(n9122) );
  OAI22_X1 U10213 ( .A1(n10647), .A2(n9120), .B1(n9119), .B2(n9238), .ZN(n9121) );
  AOI211_X1 U10214 ( .C1(n9278), .C2(n10639), .A(n9122), .B(n9121), .ZN(n9123)
         );
  OAI21_X1 U10215 ( .B1(n9124), .B2(n9223), .A(n9123), .ZN(P2_U3211) );
  AND2_X1 U10216 ( .A1(n9126), .A2(n9125), .ZN(n9128) );
  OAI21_X1 U10217 ( .B1(n9129), .B2(n9128), .A(n9127), .ZN(n9131) );
  AOI222_X1 U10218 ( .A1(n9211), .A2(n9131), .B1(n9295), .B2(n9216), .C1(n9130), .C2(n10658), .ZN(n9282) );
  OAI22_X1 U10219 ( .A1(n10647), .A2(n9133), .B1(n9132), .B2(n10638), .ZN(
        n9137) );
  NOR2_X1 U10220 ( .A1(n9115), .A2(n9134), .ZN(n9281) );
  NOR3_X1 U10221 ( .A1(n9281), .A2(n9135), .A3(n9230), .ZN(n9136) );
  AOI211_X1 U10222 ( .C1(n10641), .C2(n9138), .A(n9137), .B(n9136), .ZN(n9139)
         );
  OAI21_X1 U10223 ( .B1(n9282), .B2(n9223), .A(n9139), .ZN(P2_U3212) );
  OR2_X1 U10224 ( .A1(n9160), .A2(n9140), .ZN(n9143) );
  NAND2_X1 U10225 ( .A1(n9143), .A2(n9141), .ZN(n9147) );
  NAND2_X1 U10226 ( .A1(n9143), .A2(n9142), .ZN(n9145) );
  INV_X1 U10227 ( .A(n9154), .ZN(n9144) );
  NAND2_X1 U10228 ( .A1(n9145), .A2(n9144), .ZN(n9146) );
  NAND2_X1 U10229 ( .A1(n9147), .A2(n9146), .ZN(n9150) );
  OAI22_X1 U10230 ( .A1(n10755), .A2(n9236), .B1(n9148), .B2(n10754), .ZN(
        n9149) );
  AOI21_X1 U10231 ( .B1(n9150), .B2(n9211), .A(n9149), .ZN(n9291) );
  OAI22_X1 U10232 ( .A1(n10647), .A2(n9152), .B1(n9151), .B2(n9238), .ZN(n9153) );
  AOI21_X1 U10233 ( .B1(n9331), .B2(n10641), .A(n9153), .ZN(n9158) );
  NAND2_X1 U10234 ( .A1(n9155), .A2(n9154), .ZN(n9156) );
  NAND2_X1 U10235 ( .A1(n5295), .A2(n9156), .ZN(n9289) );
  NAND2_X1 U10236 ( .A1(n9289), .A2(n10639), .ZN(n9157) );
  OAI211_X1 U10237 ( .C1(n9291), .C2(n9223), .A(n9158), .B(n9157), .ZN(
        P2_U3213) );
  XNOR2_X1 U10238 ( .A(n9160), .B(n9159), .ZN(n9161) );
  AOI22_X1 U10239 ( .A1(n9161), .A2(n9211), .B1(n9216), .B2(n9194), .ZN(n9298)
         );
  OAI21_X1 U10240 ( .B1(n9164), .B2(n9163), .A(n9162), .ZN(n9299) );
  INV_X1 U10241 ( .A(n9165), .ZN(n9166) );
  OAI22_X1 U10242 ( .A1(n10647), .A2(n5684), .B1(n9166), .B2(n10638), .ZN(
        n9167) );
  AOI21_X1 U10243 ( .B1(n9195), .B2(n9295), .A(n9167), .ZN(n9169) );
  NAND2_X1 U10244 ( .A1(n9296), .A2(n10641), .ZN(n9168) );
  OAI211_X1 U10245 ( .C1(n9299), .C2(n9230), .A(n9169), .B(n9168), .ZN(n9170)
         );
  INV_X1 U10246 ( .A(n9170), .ZN(n9171) );
  OAI21_X1 U10247 ( .B1(n9298), .B2(n9223), .A(n9171), .ZN(P2_U3214) );
  XNOR2_X1 U10248 ( .A(n9172), .B(n9173), .ZN(n9175) );
  NOR2_X1 U10249 ( .A1(n9201), .A2(n9236), .ZN(n9174) );
  AOI21_X1 U10250 ( .B1(n9175), .B2(n9211), .A(n9174), .ZN(n10759) );
  AOI22_X1 U10251 ( .A1(n9223), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n9176), .B2(
        n9222), .ZN(n9177) );
  OAI21_X1 U10252 ( .B1(n10755), .B2(n9178), .A(n9177), .ZN(n9179) );
  AOI21_X1 U10253 ( .B1(n10752), .B2(n10641), .A(n9179), .ZN(n9184) );
  NAND2_X1 U10254 ( .A1(n9182), .A2(n9181), .ZN(n10750) );
  NAND3_X1 U10255 ( .A1(n9180), .A2(n10639), .A3(n10750), .ZN(n9183) );
  OAI211_X1 U10256 ( .C1(n10759), .C2(n9223), .A(n9184), .B(n9183), .ZN(
        P2_U3215) );
  XOR2_X1 U10257 ( .A(n9185), .B(n9190), .Z(n9186) );
  AOI22_X1 U10258 ( .A1(n9186), .A2(n9211), .B1(n9216), .B2(n9217), .ZN(n10742) );
  NOR2_X1 U10259 ( .A1(n5048), .A2(n9203), .ZN(n9202) );
  NOR2_X1 U10260 ( .A1(n9202), .A2(n9188), .ZN(n9189) );
  XOR2_X1 U10261 ( .A(n9190), .B(n9189), .Z(n10745) );
  OAI22_X1 U10262 ( .A1(n10647), .A2(n9192), .B1(n9191), .B2(n10638), .ZN(
        n9193) );
  AOI21_X1 U10263 ( .B1(n9195), .B2(n9194), .A(n9193), .ZN(n9196) );
  OAI21_X1 U10264 ( .B1(n10741), .B2(n9225), .A(n9196), .ZN(n9197) );
  AOI21_X1 U10265 ( .B1(n10745), .B2(n10639), .A(n9197), .ZN(n9198) );
  OAI21_X1 U10266 ( .B1(n10742), .B2(n9223), .A(n9198), .ZN(P2_U3216) );
  XNOR2_X1 U10267 ( .A(n9199), .B(n9203), .ZN(n9200) );
  OAI222_X1 U10268 ( .A1(n10754), .A2(n9201), .B1(n9236), .B2(n9237), .C1(
        n9234), .C2(n9200), .ZN(n10733) );
  INV_X1 U10269 ( .A(n10733), .ZN(n9208) );
  AOI21_X1 U10270 ( .B1(n5048), .B2(n9203), .A(n9202), .ZN(n10735) );
  AOI22_X1 U10271 ( .A1(n9223), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n9204), .B2(
        n9222), .ZN(n9205) );
  OAI21_X1 U10272 ( .B1(n10732), .B2(n9225), .A(n9205), .ZN(n9206) );
  AOI21_X1 U10273 ( .B1(n10735), .B2(n10639), .A(n9206), .ZN(n9207) );
  OAI21_X1 U10274 ( .B1(n9208), .B2(n9223), .A(n9207), .ZN(P2_U3217) );
  INV_X1 U10275 ( .A(n9213), .ZN(n9209) );
  XNOR2_X1 U10276 ( .A(n9210), .B(n9209), .ZN(n10724) );
  INV_X1 U10277 ( .A(n10724), .ZN(n9229) );
  OAI211_X1 U10278 ( .C1(n9214), .C2(n9213), .A(n9212), .B(n9211), .ZN(n9219)
         );
  AOI22_X1 U10279 ( .A1(n9217), .A2(n10658), .B1(n9216), .B2(n9215), .ZN(n9218) );
  NAND2_X1 U10280 ( .A1(n9219), .A2(n9218), .ZN(n10728) );
  INV_X1 U10281 ( .A(n9220), .ZN(n9221) );
  AOI22_X1 U10282 ( .A1(n9223), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n9222), .B2(
        n9221), .ZN(n9224) );
  OAI21_X1 U10283 ( .B1(n9226), .B2(n9225), .A(n9224), .ZN(n9227) );
  AOI21_X1 U10284 ( .B1(n10728), .B2(n10643), .A(n9227), .ZN(n9228) );
  OAI21_X1 U10285 ( .B1(n9230), .B2(n9229), .A(n9228), .ZN(P2_U3218) );
  XNOR2_X1 U10286 ( .A(n9231), .B(n9232), .ZN(n9233) );
  OAI222_X1 U10287 ( .A1(n10754), .A2(n9237), .B1(n9236), .B2(n9235), .C1(
        n9234), .C2(n9233), .ZN(n10719) );
  OAI22_X1 U10288 ( .A1(n10718), .A2(n9240), .B1(n9239), .B2(n9238), .ZN(n9241) );
  OAI21_X1 U10289 ( .B1(n10719), .B2(n9241), .A(n10643), .ZN(n9246) );
  OAI21_X1 U10290 ( .B1(n9244), .B2(n9243), .A(n9242), .ZN(n10721) );
  NAND2_X1 U10291 ( .A1(n10721), .A2(n10639), .ZN(n9245) );
  OAI211_X1 U10292 ( .C1(n5970), .C2(n10647), .A(n9246), .B(n9245), .ZN(
        P2_U3219) );
  NAND2_X1 U10293 ( .A1(n9300), .A2(n10761), .ZN(n9248) );
  NAND2_X1 U10294 ( .A1(n10760), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n9247) );
  OAI211_X1 U10295 ( .C1(n9302), .C2(n9288), .A(n9248), .B(n9247), .ZN(
        P2_U3490) );
  NAND2_X1 U10296 ( .A1(n10760), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n9249) );
  OAI211_X1 U10297 ( .C1(n9305), .C2(n9288), .A(n9249), .B(n9248), .ZN(
        P2_U3489) );
  OR2_X1 U10298 ( .A1(n10761), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n9251) );
  OAI21_X1 U10299 ( .B1(n9254), .B2(n9288), .A(n9253), .ZN(P2_U3487) );
  INV_X1 U10300 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n9257) );
  AOI21_X1 U10301 ( .B1(n10749), .B2(n9256), .A(n9255), .ZN(n9306) );
  MUX2_X1 U10302 ( .A(n9257), .B(n9306), .S(n10761), .Z(n9258) );
  OAI21_X1 U10303 ( .B1(n9309), .B2(n9288), .A(n9258), .ZN(P2_U3486) );
  AOI22_X1 U10304 ( .A1(n9260), .A2(n10751), .B1(n10658), .B2(n9259), .ZN(
        n9263) );
  NAND3_X1 U10305 ( .A1(n9261), .A2(n9071), .A3(n10749), .ZN(n9262) );
  NAND3_X1 U10306 ( .A1(n9264), .A2(n9263), .A3(n9262), .ZN(n9310) );
  MUX2_X1 U10307 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n9310), .S(n10761), .Z(
        P2_U3485) );
  INV_X1 U10308 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n9267) );
  AOI21_X1 U10309 ( .B1(n10749), .B2(n9266), .A(n9265), .ZN(n9311) );
  MUX2_X1 U10310 ( .A(n9267), .B(n9311), .S(n10761), .Z(n9268) );
  OAI21_X1 U10311 ( .B1(n9314), .B2(n9288), .A(n9268), .ZN(P2_U3484) );
  INV_X1 U10312 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n9271) );
  AOI21_X1 U10313 ( .B1(n9270), .B2(n10749), .A(n9269), .ZN(n9315) );
  MUX2_X1 U10314 ( .A(n9271), .B(n9315), .S(n10761), .Z(n9272) );
  OAI21_X1 U10315 ( .B1(n9318), .B2(n9288), .A(n9272), .ZN(P2_U3483) );
  AOI22_X1 U10316 ( .A1(n9274), .A2(n10749), .B1(n10751), .B2(n9273), .ZN(
        n9275) );
  NAND2_X1 U10317 ( .A1(n9276), .A2(n9275), .ZN(n9319) );
  MUX2_X1 U10318 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n9319), .S(n10761), .Z(
        P2_U3482) );
  INV_X1 U10319 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n9279) );
  AOI21_X1 U10320 ( .B1(n9278), .B2(n10749), .A(n9277), .ZN(n9320) );
  MUX2_X1 U10321 ( .A(n9279), .B(n9320), .S(n10761), .Z(n9280) );
  OAI21_X1 U10322 ( .B1(n9323), .B2(n9288), .A(n9280), .ZN(P2_U3481) );
  INV_X1 U10323 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n9286) );
  NOR2_X1 U10324 ( .A1(n9281), .A2(n10710), .ZN(n9285) );
  INV_X1 U10325 ( .A(n9282), .ZN(n9283) );
  AOI21_X1 U10326 ( .B1(n9285), .B2(n9284), .A(n9283), .ZN(n9324) );
  MUX2_X1 U10327 ( .A(n9286), .B(n9324), .S(n10761), .Z(n9287) );
  OAI21_X1 U10328 ( .B1(n9328), .B2(n9288), .A(n9287), .ZN(P2_U3480) );
  NAND2_X1 U10329 ( .A1(n9289), .A2(n10749), .ZN(n9290) );
  NAND2_X1 U10330 ( .A1(n9291), .A2(n9290), .ZN(n9329) );
  MUX2_X1 U10331 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n9329), .S(n10761), .Z(
        n9292) );
  AOI21_X1 U10332 ( .B1(n9293), .B2(n9331), .A(n9292), .ZN(n9294) );
  INV_X1 U10333 ( .A(n9294), .ZN(P2_U3479) );
  AOI22_X1 U10334 ( .A1(n9296), .A2(n10751), .B1(n10658), .B2(n9295), .ZN(
        n9297) );
  OAI211_X1 U10335 ( .C1(n10710), .C2(n9299), .A(n9298), .B(n9297), .ZN(n9333)
         );
  MUX2_X1 U10336 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n9333), .S(n10761), .Z(
        P2_U3478) );
  NAND2_X1 U10337 ( .A1(n10764), .A2(n9300), .ZN(n9303) );
  NAND2_X1 U10338 ( .A1(n6872), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n9301) );
  OAI211_X1 U10339 ( .C1(n9302), .C2(n9327), .A(n9303), .B(n9301), .ZN(
        P2_U3458) );
  NAND2_X1 U10340 ( .A1(n6872), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n9304) );
  OAI211_X1 U10341 ( .C1(n9305), .C2(n9327), .A(n9304), .B(n9303), .ZN(
        P2_U3457) );
  MUX2_X1 U10342 ( .A(n9307), .B(n9306), .S(n10764), .Z(n9308) );
  OAI21_X1 U10343 ( .B1(n9309), .B2(n9327), .A(n9308), .ZN(P2_U3454) );
  MUX2_X1 U10344 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n9310), .S(n10764), .Z(
        P2_U3453) );
  MUX2_X1 U10345 ( .A(n9312), .B(n9311), .S(n10764), .Z(n9313) );
  OAI21_X1 U10346 ( .B1(n9314), .B2(n9327), .A(n9313), .ZN(P2_U3452) );
  MUX2_X1 U10347 ( .A(n9316), .B(n9315), .S(n10764), .Z(n9317) );
  OAI21_X1 U10348 ( .B1(n9318), .B2(n9327), .A(n9317), .ZN(P2_U3451) );
  MUX2_X1 U10349 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n9319), .S(n10764), .Z(
        P2_U3450) );
  MUX2_X1 U10350 ( .A(n9321), .B(n9320), .S(n10764), .Z(n9322) );
  OAI21_X1 U10351 ( .B1(n9323), .B2(n9327), .A(n9322), .ZN(P2_U3449) );
  MUX2_X1 U10352 ( .A(n9325), .B(n9324), .S(n10764), .Z(n9326) );
  OAI21_X1 U10353 ( .B1(n9328), .B2(n9327), .A(n9326), .ZN(P2_U3448) );
  MUX2_X1 U10354 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n9329), .S(n10764), .Z(
        n9330) );
  AOI21_X1 U10355 ( .B1(n6880), .B2(n9331), .A(n9330), .ZN(n9332) );
  INV_X1 U10356 ( .A(n9332), .ZN(P2_U3447) );
  MUX2_X1 U10357 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n9333), .S(n10764), .Z(
        P2_U3446) );
  INV_X1 U10358 ( .A(n9334), .ZN(n10005) );
  NOR4_X1 U10359 ( .A1(n9335), .A2(P2_IR_REG_30__SCAN_IN), .A3(P2_U3151), .A4(
        n5617), .ZN(n9336) );
  AOI21_X1 U10360 ( .B1(n9345), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n9336), .ZN(
        n9337) );
  OAI21_X1 U10361 ( .B1(n10005), .B2(n8052), .A(n9337), .ZN(P2_U3264) );
  INV_X1 U10362 ( .A(n9338), .ZN(n10008) );
  AOI22_X1 U10363 ( .A1(n9339), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n9345), .ZN(n9340) );
  OAI21_X1 U10364 ( .B1(n10008), .B2(n8052), .A(n9340), .ZN(P2_U3265) );
  INV_X1 U10365 ( .A(n6802), .ZN(n10011) );
  AOI22_X1 U10366 ( .A1(n9341), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n9345), .ZN(n9342) );
  OAI21_X1 U10367 ( .B1(n10011), .B2(n8052), .A(n9342), .ZN(P2_U3266) );
  INV_X1 U10368 ( .A(n9343), .ZN(n10015) );
  AOI21_X1 U10369 ( .B1(P1_DATAO_REG_28__SCAN_IN), .B2(n9345), .A(n9344), .ZN(
        n9346) );
  OAI21_X1 U10370 ( .B1(n10015), .B2(n8052), .A(n9346), .ZN(P2_U3267) );
  INV_X1 U10371 ( .A(n9347), .ZN(n9348) );
  MUX2_X1 U10372 ( .A(n9348), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  XNOR2_X1 U10373 ( .A(n9351), .B(n9350), .ZN(n9352) );
  XNOR2_X1 U10374 ( .A(n9349), .B(n9352), .ZN(n9360) );
  NAND2_X1 U10375 ( .A1(n9486), .A2(n9353), .ZN(n9356) );
  NAND2_X1 U10376 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n10340)
         );
  INV_X1 U10377 ( .A(n10340), .ZN(n9354) );
  AOI21_X1 U10378 ( .B1(n9488), .B2(n9820), .A(n9354), .ZN(n9355) );
  OAI211_X1 U10379 ( .C1(n9357), .C2(n9491), .A(n9356), .B(n9355), .ZN(n9358)
         );
  AOI21_X1 U10380 ( .B1(n9943), .B2(n9494), .A(n9358), .ZN(n9359) );
  OAI21_X1 U10381 ( .B1(n9360), .B2(n9496), .A(n9359), .ZN(P1_U3215) );
  INV_X1 U10382 ( .A(n9361), .ZN(n9420) );
  AOI21_X1 U10383 ( .B1(n9363), .B2(n9447), .A(n9362), .ZN(n9364) );
  OAI21_X1 U10384 ( .B1(n9420), .B2(n9364), .A(n9472), .ZN(n9369) );
  NOR2_X1 U10385 ( .A1(n9712), .A2(n9454), .ZN(n9367) );
  OAI22_X1 U10386 ( .A1(n9743), .A2(n9491), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9365), .ZN(n9366) );
  AOI211_X1 U10387 ( .C1(n9488), .C2(n9707), .A(n9367), .B(n9366), .ZN(n9368)
         );
  OAI211_X1 U10388 ( .C1(n9972), .C2(n9480), .A(n9369), .B(n9368), .ZN(
        P1_U3216) );
  AOI21_X1 U10389 ( .B1(n9371), .B2(n9370), .A(n4956), .ZN(n9376) );
  NOR2_X1 U10390 ( .A1(n9454), .A2(n9785), .ZN(n9374) );
  NAND2_X1 U10391 ( .A1(n9777), .A2(n9488), .ZN(n9372) );
  NAND2_X1 U10392 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9609) );
  OAI211_X1 U10393 ( .C1(n9412), .C2(n9491), .A(n9372), .B(n9609), .ZN(n9373)
         );
  AOI211_X1 U10394 ( .C1(n9784), .C2(n9494), .A(n9374), .B(n9373), .ZN(n9375)
         );
  OAI21_X1 U10395 ( .B1(n9376), .B2(n9496), .A(n9375), .ZN(P1_U3219) );
  INV_X1 U10396 ( .A(n9377), .ZN(n9380) );
  OAI21_X1 U10397 ( .B1(n9380), .B2(n9379), .A(n9378), .ZN(n9382) );
  NAND3_X1 U10398 ( .A1(n9382), .A2(n9472), .A3(n9381), .ZN(n9387) );
  INV_X1 U10399 ( .A(n9383), .ZN(n9750) );
  AOI22_X1 U10400 ( .A1(n9777), .A2(n9451), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3086), .ZN(n9384) );
  OAI21_X1 U10401 ( .B1(n9743), .B2(n9434), .A(n9384), .ZN(n9385) );
  AOI21_X1 U10402 ( .B1(n9750), .B2(n9486), .A(n9385), .ZN(n9386) );
  OAI211_X1 U10403 ( .C1(n9980), .C2(n9480), .A(n9387), .B(n9386), .ZN(
        P1_U3223) );
  OAI21_X1 U10404 ( .B1(n9390), .B2(n9389), .A(n9388), .ZN(n9391) );
  NAND2_X1 U10405 ( .A1(n9391), .A2(n9472), .ZN(n9395) );
  AOI22_X1 U10406 ( .A1(n9707), .A2(n9451), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3086), .ZN(n9392) );
  OAI21_X1 U10407 ( .B1(n9678), .B2(n9454), .A(n9392), .ZN(n9393) );
  AOI21_X1 U10408 ( .B1(n9488), .B2(n9673), .A(n9393), .ZN(n9394) );
  OAI211_X1 U10409 ( .C1(n9396), .C2(n9480), .A(n9395), .B(n9394), .ZN(
        P1_U3225) );
  XOR2_X1 U10410 ( .A(n9397), .B(n9398), .Z(n9405) );
  NAND2_X1 U10411 ( .A1(n9486), .A2(n9826), .ZN(n9401) );
  AOI21_X1 U10412 ( .B1(n9488), .B2(n9819), .A(n9399), .ZN(n9400) );
  OAI211_X1 U10413 ( .C1(n9402), .C2(n9491), .A(n9401), .B(n9400), .ZN(n9403)
         );
  AOI21_X1 U10414 ( .B1(n9830), .B2(n9494), .A(n9403), .ZN(n9404) );
  OAI21_X1 U10415 ( .B1(n9405), .B2(n9496), .A(n9404), .ZN(P1_U3226) );
  XOR2_X1 U10416 ( .A(n9408), .B(n9407), .Z(n9409) );
  XNOR2_X1 U10417 ( .A(n9406), .B(n9409), .ZN(n9417) );
  NAND2_X1 U10418 ( .A1(n9451), .A2(n9500), .ZN(n9411) );
  OAI211_X1 U10419 ( .C1(n9412), .C2(n9434), .A(n9411), .B(n9410), .ZN(n9413)
         );
  AOI21_X1 U10420 ( .B1(n9414), .B2(n9486), .A(n9413), .ZN(n9416) );
  NAND2_X1 U10421 ( .A1(n9925), .A2(n9494), .ZN(n9415) );
  OAI211_X1 U10422 ( .C1(n9417), .C2(n9496), .A(n9416), .B(n9415), .ZN(
        P1_U3228) );
  NOR3_X1 U10423 ( .A1(n9420), .A2(n5089), .A3(n9419), .ZN(n9423) );
  INV_X1 U10424 ( .A(n9421), .ZN(n9422) );
  OAI21_X1 U10425 ( .B1(n9423), .B2(n9422), .A(n9472), .ZN(n9429) );
  OAI22_X1 U10426 ( .A1(n9425), .A2(n9491), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9424), .ZN(n9427) );
  NOR2_X1 U10427 ( .A1(n9476), .A2(n9434), .ZN(n9426) );
  AOI211_X1 U10428 ( .C1(n9486), .C2(n9696), .A(n9427), .B(n9426), .ZN(n9428)
         );
  OAI211_X1 U10429 ( .C1(n9968), .C2(n9480), .A(n9429), .B(n9428), .ZN(
        P1_U3229) );
  OAI21_X1 U10430 ( .B1(n9431), .B2(n9430), .A(n9377), .ZN(n9432) );
  NAND2_X1 U10431 ( .A1(n9432), .A2(n9472), .ZN(n9438) );
  NOR2_X1 U10432 ( .A1(n9454), .A2(n9765), .ZN(n9436) );
  OAI22_X1 U10433 ( .A1(n9763), .A2(n9434), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9433), .ZN(n9435) );
  AOI211_X1 U10434 ( .C1(n9451), .C2(n9807), .A(n9436), .B(n9435), .ZN(n9437)
         );
  OAI211_X1 U10435 ( .C1(n5360), .C2(n9480), .A(n9438), .B(n9437), .ZN(
        P1_U3233) );
  XOR2_X1 U10436 ( .A(n9439), .B(n9440), .Z(n9446) );
  NAND2_X1 U10437 ( .A1(n9486), .A2(n9842), .ZN(n9442) );
  AOI22_X1 U10438 ( .A1(n9488), .A2(n9501), .B1(P1_REG3_REG_13__SCAN_IN), .B2(
        P1_U3086), .ZN(n9441) );
  OAI211_X1 U10439 ( .C1(n9443), .C2(n9491), .A(n9442), .B(n9441), .ZN(n9444)
         );
  AOI21_X1 U10440 ( .B1(n9846), .B2(n9494), .A(n9444), .ZN(n9445) );
  OAI21_X1 U10441 ( .B1(n9446), .B2(n9496), .A(n9445), .ZN(P1_U3234) );
  NAND2_X1 U10442 ( .A1(n9448), .A2(n9447), .ZN(n9449) );
  XOR2_X1 U10443 ( .A(n9450), .B(n9449), .Z(n9457) );
  NAND2_X1 U10444 ( .A1(n9726), .A2(n9488), .ZN(n9453) );
  AOI22_X1 U10445 ( .A1(n9725), .A2(n9451), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3086), .ZN(n9452) );
  OAI211_X1 U10446 ( .C1(n9454), .C2(n9732), .A(n9453), .B(n9452), .ZN(n9455)
         );
  AOI21_X1 U10447 ( .B1(n9721), .B2(n9494), .A(n9455), .ZN(n9456) );
  OAI21_X1 U10448 ( .B1(n9457), .B2(n9496), .A(n9456), .ZN(P1_U3235) );
  XOR2_X1 U10449 ( .A(n9460), .B(n9459), .Z(n9461) );
  XNOR2_X1 U10450 ( .A(n9458), .B(n9461), .ZN(n9467) );
  NAND2_X1 U10451 ( .A1(n9807), .A2(n9488), .ZN(n9462) );
  NAND2_X1 U10452 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n10364)
         );
  OAI211_X1 U10453 ( .C1(n9463), .C2(n9491), .A(n9462), .B(n10364), .ZN(n9465)
         );
  NOR2_X1 U10454 ( .A1(n9989), .A2(n9480), .ZN(n9464) );
  AOI211_X1 U10455 ( .C1(n9486), .C2(n9799), .A(n9465), .B(n9464), .ZN(n9466)
         );
  OAI21_X1 U10456 ( .B1(n9467), .B2(n9496), .A(n9466), .ZN(P1_U3238) );
  INV_X1 U10457 ( .A(n9388), .ZN(n9470) );
  OAI21_X1 U10458 ( .B1(n9470), .B2(n9469), .A(n9468), .ZN(n9473) );
  NAND3_X1 U10459 ( .A1(n9473), .A2(n9472), .A3(n9471), .ZN(n9479) );
  INV_X1 U10460 ( .A(n9474), .ZN(n9661) );
  AOI22_X1 U10461 ( .A1(n9661), .A2(n9486), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3086), .ZN(n9475) );
  OAI21_X1 U10462 ( .B1(n9476), .B2(n9491), .A(n9475), .ZN(n9477) );
  AOI21_X1 U10463 ( .B1(n9488), .B2(n9656), .A(n9477), .ZN(n9478) );
  OAI211_X1 U10464 ( .C1(n9963), .C2(n9480), .A(n9479), .B(n9478), .ZN(
        P1_U3240) );
  XNOR2_X1 U10465 ( .A(n9483), .B(n9482), .ZN(n9484) );
  XNOR2_X1 U10466 ( .A(n9481), .B(n9484), .ZN(n9497) );
  NAND2_X1 U10467 ( .A1(n9486), .A2(n9485), .ZN(n9490) );
  NAND2_X1 U10468 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n10351)
         );
  INV_X1 U10469 ( .A(n10351), .ZN(n9487) );
  AOI21_X1 U10470 ( .B1(n9488), .B2(n9500), .A(n9487), .ZN(n9489) );
  OAI211_X1 U10471 ( .C1(n9492), .C2(n9491), .A(n9490), .B(n9489), .ZN(n9493)
         );
  AOI21_X1 U10472 ( .B1(n9998), .B2(n9494), .A(n9493), .ZN(n9495) );
  OAI21_X1 U10473 ( .B1(n9497), .B2(n9496), .A(n9495), .ZN(P1_U3241) );
  MUX2_X1 U10474 ( .A(n9616), .B(P1_DATAO_REG_31__SCAN_IN), .S(n9528), .Z(
        P1_U3585) );
  MUX2_X1 U10475 ( .A(n9498), .B(P1_DATAO_REG_30__SCAN_IN), .S(n9528), .Z(
        P1_U3584) );
  MUX2_X1 U10476 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9499), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U10477 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9656), .S(P1_U3973), .Z(
        P1_U3581) );
  MUX2_X1 U10478 ( .A(n9673), .B(P1_DATAO_REG_26__SCAN_IN), .S(n9528), .Z(
        P1_U3580) );
  MUX2_X1 U10479 ( .A(n9689), .B(P1_DATAO_REG_25__SCAN_IN), .S(n9528), .Z(
        P1_U3579) );
  MUX2_X1 U10480 ( .A(n9726), .B(P1_DATAO_REG_23__SCAN_IN), .S(n9528), .Z(
        P1_U3577) );
  MUX2_X1 U10481 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9706), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U10482 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9725), .S(P1_U3973), .Z(
        P1_U3575) );
  MUX2_X1 U10483 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9777), .S(P1_U3973), .Z(
        P1_U3574) );
  MUX2_X1 U10484 ( .A(n9807), .B(P1_DATAO_REG_19__SCAN_IN), .S(n9528), .Z(
        P1_U3573) );
  MUX2_X1 U10485 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9776), .S(P1_U3973), .Z(
        P1_U3572) );
  MUX2_X1 U10486 ( .A(n9500), .B(P1_DATAO_REG_16__SCAN_IN), .S(n9528), .Z(
        P1_U3570) );
  MUX2_X1 U10487 ( .A(n9820), .B(P1_DATAO_REG_15__SCAN_IN), .S(n9528), .Z(
        P1_U3569) );
  MUX2_X1 U10488 ( .A(n9501), .B(P1_DATAO_REG_14__SCAN_IN), .S(n9528), .Z(
        P1_U3568) );
  MUX2_X1 U10489 ( .A(n9502), .B(P1_DATAO_REG_13__SCAN_IN), .S(n9528), .Z(
        P1_U3567) );
  MUX2_X1 U10490 ( .A(n9503), .B(P1_DATAO_REG_12__SCAN_IN), .S(n9528), .Z(
        P1_U3566) );
  MUX2_X1 U10491 ( .A(n9504), .B(P1_DATAO_REG_11__SCAN_IN), .S(n9528), .Z(
        P1_U3565) );
  MUX2_X1 U10492 ( .A(n9505), .B(P1_DATAO_REG_10__SCAN_IN), .S(n9528), .Z(
        P1_U3564) );
  MUX2_X1 U10493 ( .A(n9506), .B(P1_DATAO_REG_9__SCAN_IN), .S(n9528), .Z(
        P1_U3563) );
  MUX2_X1 U10494 ( .A(n9507), .B(P1_DATAO_REG_8__SCAN_IN), .S(n9528), .Z(
        P1_U3562) );
  MUX2_X1 U10495 ( .A(n9508), .B(P1_DATAO_REG_7__SCAN_IN), .S(n9528), .Z(
        P1_U3561) );
  MUX2_X1 U10496 ( .A(n9509), .B(P1_DATAO_REG_6__SCAN_IN), .S(n9528), .Z(
        P1_U3560) );
  MUX2_X1 U10497 ( .A(n9510), .B(P1_DATAO_REG_5__SCAN_IN), .S(n9528), .Z(
        P1_U3559) );
  MUX2_X1 U10498 ( .A(n9511), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9528), .Z(
        P1_U3558) );
  MUX2_X1 U10499 ( .A(n10544), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9528), .Z(
        P1_U3557) );
  MUX2_X1 U10500 ( .A(n9512), .B(P1_DATAO_REG_2__SCAN_IN), .S(n9528), .Z(
        P1_U3556) );
  MUX2_X1 U10501 ( .A(n10542), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9528), .Z(
        P1_U3555) );
  MUX2_X1 U10502 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n9513), .S(P1_U3973), .Z(
        P1_U3554) );
  OAI22_X1 U10503 ( .A1(n10394), .A2(n10224), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6364), .ZN(n9514) );
  AOI21_X1 U10504 ( .B1(n10390), .B2(n9515), .A(n9514), .ZN(n9524) );
  OAI211_X1 U10505 ( .C1(n9518), .C2(n9517), .A(n10329), .B(n9516), .ZN(n9523)
         );
  OAI211_X1 U10506 ( .C1(n9521), .C2(n9520), .A(n10334), .B(n9519), .ZN(n9522)
         );
  NAND3_X1 U10507 ( .A1(n9524), .A2(n9523), .A3(n9522), .ZN(P1_U3244) );
  NAND2_X1 U10508 ( .A1(n10013), .A2(n9525), .ZN(n9531) );
  NAND2_X1 U10509 ( .A1(n10013), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n9527) );
  XNOR2_X1 U10510 ( .A(n9527), .B(n9526), .ZN(n9529) );
  AOI21_X1 U10511 ( .B1(n9529), .B2(n9531), .A(n9528), .ZN(n9530) );
  OAI21_X1 U10512 ( .B1(n9532), .B2(n9531), .A(n9530), .ZN(n9571) );
  INV_X1 U10513 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n9533) );
  OAI22_X1 U10514 ( .A1(n10394), .A2(n9533), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6376), .ZN(n9534) );
  AOI21_X1 U10515 ( .B1(n10390), .B2(n9535), .A(n9534), .ZN(n9544) );
  OAI211_X1 U10516 ( .C1(n9538), .C2(n9537), .A(n10334), .B(n9536), .ZN(n9543)
         );
  OAI211_X1 U10517 ( .C1(n9541), .C2(n9540), .A(n10329), .B(n9539), .ZN(n9542)
         );
  NAND4_X1 U10518 ( .A1(n9571), .A2(n9544), .A3(n9543), .A4(n9542), .ZN(
        P1_U3245) );
  INV_X1 U10519 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n9546) );
  OAI21_X1 U10520 ( .B1(n10394), .B2(n9546), .A(n9545), .ZN(n9547) );
  AOI21_X1 U10521 ( .B1(n10390), .B2(n9548), .A(n9547), .ZN(n9557) );
  OAI211_X1 U10522 ( .C1(n9551), .C2(n9550), .A(n10334), .B(n9549), .ZN(n9556)
         );
  OAI211_X1 U10523 ( .C1(n9554), .C2(n9553), .A(n10329), .B(n9552), .ZN(n9555)
         );
  NAND3_X1 U10524 ( .A1(n9557), .A2(n9556), .A3(n9555), .ZN(P1_U3246) );
  INV_X1 U10525 ( .A(n9558), .ZN(n9559) );
  NOR2_X1 U10526 ( .A1(n10338), .A2(n9559), .ZN(n9560) );
  AOI211_X1 U10527 ( .C1(n9607), .C2(P1_ADDR_REG_4__SCAN_IN), .A(n9561), .B(
        n9560), .ZN(n9570) );
  OAI211_X1 U10528 ( .C1(n9564), .C2(n9563), .A(n10329), .B(n9562), .ZN(n9569)
         );
  OAI211_X1 U10529 ( .C1(n9567), .C2(n9566), .A(n10334), .B(n9565), .ZN(n9568)
         );
  NAND4_X1 U10530 ( .A1(n9571), .A2(n9570), .A3(n9569), .A4(n9568), .ZN(
        P1_U3247) );
  INV_X1 U10531 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n9573) );
  OAI21_X1 U10532 ( .B1(n10394), .B2(n9573), .A(n9572), .ZN(n9574) );
  AOI21_X1 U10533 ( .B1(n10390), .B2(n9575), .A(n9574), .ZN(n9584) );
  OAI211_X1 U10534 ( .C1(n9578), .C2(n9577), .A(n10334), .B(n9576), .ZN(n9583)
         );
  OAI211_X1 U10535 ( .C1(n9581), .C2(n9580), .A(n10329), .B(n9579), .ZN(n9582)
         );
  NAND3_X1 U10536 ( .A1(n9584), .A2(n9583), .A3(n9582), .ZN(P1_U3248) );
  INV_X1 U10537 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n9586) );
  OAI21_X1 U10538 ( .B1(n10394), .B2(n9586), .A(n9585), .ZN(n9587) );
  AOI21_X1 U10539 ( .B1(n10390), .B2(n9588), .A(n9587), .ZN(n9597) );
  OAI211_X1 U10540 ( .C1(n9591), .C2(n9590), .A(n10334), .B(n9589), .ZN(n9596)
         );
  OAI211_X1 U10541 ( .C1(n9594), .C2(n9593), .A(n10329), .B(n9592), .ZN(n9595)
         );
  NAND3_X1 U10542 ( .A1(n9597), .A2(n9596), .A3(n9595), .ZN(P1_U3249) );
  OAI21_X1 U10543 ( .B1(n9604), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9598), .ZN(
        n10360) );
  NAND2_X1 U10544 ( .A1(n10363), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9599) );
  OAI21_X1 U10545 ( .B1(n10363), .B2(P1_REG2_REG_18__SCAN_IN), .A(n9599), .ZN(
        n10359) );
  OR2_X1 U10546 ( .A1(n10360), .A2(n10359), .ZN(n10357) );
  NAND2_X1 U10547 ( .A1(n10357), .A2(n9599), .ZN(n9602) );
  INV_X1 U10548 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n9600) );
  MUX2_X1 U10549 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n9600), .S(n4926), .Z(n9601) );
  XNOR2_X1 U10550 ( .A(n9602), .B(n9601), .ZN(n9613) );
  OAI21_X1 U10551 ( .B1(P1_REG1_REG_17__SCAN_IN), .B2(n9604), .A(n9603), .ZN(
        n10355) );
  XNOR2_X1 U10552 ( .A(n10363), .B(P1_REG1_REG_18__SCAN_IN), .ZN(n10356) );
  NOR2_X1 U10553 ( .A1(n10355), .A2(n10356), .ZN(n10354) );
  AOI21_X1 U10554 ( .B1(P1_REG1_REG_18__SCAN_IN), .B2(n10363), .A(n10354), 
        .ZN(n9606) );
  XNOR2_X1 U10555 ( .A(n4926), .B(n9915), .ZN(n9605) );
  XNOR2_X1 U10556 ( .A(n9606), .B(n9605), .ZN(n9611) );
  NAND2_X1 U10557 ( .A1(n9607), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n9608) );
  OAI211_X1 U10558 ( .C1(n10338), .C2(n6738), .A(n9609), .B(n9608), .ZN(n9610)
         );
  AOI21_X1 U10559 ( .B1(n9611), .B2(n10334), .A(n9610), .ZN(n9612) );
  OAI21_X1 U10560 ( .B1(n9613), .B2(n10383), .A(n9612), .ZN(P1_U3262) );
  NOR2_X2 U10561 ( .A1(n4947), .A2(n9621), .ZN(n9620) );
  XNOR2_X1 U10562 ( .A(n9951), .B(n9620), .ZN(n9614) );
  NAND2_X1 U10563 ( .A1(n9865), .A2(n4924), .ZN(n9619) );
  AND2_X1 U10564 ( .A1(n9616), .A2(n9615), .ZN(n9868) );
  INV_X1 U10565 ( .A(n9868), .ZN(n9617) );
  NOR2_X1 U10566 ( .A1(n9617), .A2(n9800), .ZN(n9622) );
  AOI21_X1 U10567 ( .B1(n10555), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9622), .ZN(
        n9618) );
  OAI211_X1 U10568 ( .C1(n9951), .C2(n9802), .A(n9619), .B(n9618), .ZN(
        P1_U3263) );
  AOI211_X1 U10569 ( .C1(n9621), .C2(n4947), .A(n9797), .B(n9620), .ZN(n9869)
         );
  NAND2_X1 U10570 ( .A1(n9869), .A2(n4924), .ZN(n9624) );
  AOI21_X1 U10571 ( .B1(n10555), .B2(P1_REG2_REG_30__SCAN_IN), .A(n9622), .ZN(
        n9623) );
  OAI211_X1 U10572 ( .C1(n9955), .C2(n9802), .A(n9624), .B(n9623), .ZN(
        P1_U3264) );
  INV_X1 U10573 ( .A(n9625), .ZN(n9632) );
  AOI22_X1 U10574 ( .A1(n9626), .A2(n10554), .B1(P1_REG2_REG_28__SCAN_IN), 
        .B2(n9800), .ZN(n9627) );
  OAI21_X1 U10575 ( .B1(n9628), .B2(n9802), .A(n9627), .ZN(n9631) );
  NOR2_X1 U10576 ( .A1(n9629), .A2(n9836), .ZN(n9630) );
  OAI21_X1 U10577 ( .B1(n10555), .B2(n9634), .A(n9633), .ZN(P1_U3265) );
  XNOR2_X1 U10578 ( .A(n9635), .B(n9636), .ZN(n9874) );
  INV_X1 U10579 ( .A(n9874), .ZN(n9651) );
  XNOR2_X1 U10580 ( .A(n9637), .B(n9636), .ZN(n9638) );
  NAND2_X1 U10581 ( .A1(n9638), .A2(n10546), .ZN(n9643) );
  OAI22_X1 U10582 ( .A1(n9640), .A2(n9764), .B1(n9639), .B2(n9762), .ZN(n9641)
         );
  INV_X1 U10583 ( .A(n9641), .ZN(n9642) );
  NAND2_X1 U10584 ( .A1(n9643), .A2(n9642), .ZN(n9872) );
  AOI211_X1 U10585 ( .C1(n9645), .C2(n9659), .A(n9797), .B(n9644), .ZN(n9873)
         );
  NAND2_X1 U10586 ( .A1(n9873), .A2(n4924), .ZN(n9648) );
  AOI22_X1 U10587 ( .A1(n9646), .A2(n10554), .B1(P1_REG2_REG_27__SCAN_IN), 
        .B2(n10555), .ZN(n9647) );
  OAI211_X1 U10588 ( .C1(n9959), .C2(n9802), .A(n9648), .B(n9647), .ZN(n9649)
         );
  AOI21_X1 U10589 ( .B1(n10524), .B2(n9872), .A(n9649), .ZN(n9650) );
  OAI21_X1 U10590 ( .B1(n9651), .B2(n9836), .A(n9650), .ZN(P1_U3266) );
  XNOR2_X1 U10591 ( .A(n9652), .B(n5163), .ZN(n9879) );
  INV_X1 U10592 ( .A(n9879), .ZN(n9666) );
  OAI21_X1 U10593 ( .B1(n5163), .B2(n9654), .A(n9653), .ZN(n9655) );
  NAND2_X1 U10594 ( .A1(n9655), .A2(n10546), .ZN(n9658) );
  AOI22_X1 U10595 ( .A1(n9656), .A2(n10543), .B1(n9821), .B2(n9689), .ZN(n9657) );
  NAND2_X1 U10596 ( .A1(n9658), .A2(n9657), .ZN(n9877) );
  AOI211_X1 U10597 ( .C1(n9660), .C2(n9675), .A(n9797), .B(n5366), .ZN(n9878)
         );
  NAND2_X1 U10598 ( .A1(n9878), .A2(n4924), .ZN(n9663) );
  AOI22_X1 U10599 ( .A1(n9661), .A2(n10554), .B1(P1_REG2_REG_26__SCAN_IN), 
        .B2(n9800), .ZN(n9662) );
  OAI211_X1 U10600 ( .C1(n9963), .C2(n9802), .A(n9663), .B(n9662), .ZN(n9664)
         );
  AOI21_X1 U10601 ( .B1(n10524), .B2(n9877), .A(n9664), .ZN(n9665) );
  OAI21_X1 U10602 ( .B1(n9666), .B2(n9836), .A(n9665), .ZN(P1_U3267) );
  XNOR2_X1 U10603 ( .A(n9668), .B(n9667), .ZN(n9886) );
  AOI22_X1 U10604 ( .A1(n9883), .A2(n10552), .B1(P1_REG2_REG_25__SCAN_IN), 
        .B2(n10555), .ZN(n9681) );
  INV_X1 U10605 ( .A(n9669), .ZN(n9672) );
  OAI21_X1 U10606 ( .B1(n9672), .B2(n9671), .A(n9670), .ZN(n9674) );
  AOI222_X1 U10607 ( .A1(n10546), .A2(n9674), .B1(n9673), .B2(n10543), .C1(
        n9707), .C2(n10541), .ZN(n9885) );
  INV_X1 U10608 ( .A(n9675), .ZN(n9676) );
  AOI211_X1 U10609 ( .C1(n9883), .C2(n9692), .A(n9797), .B(n9676), .ZN(n9882)
         );
  NAND2_X1 U10610 ( .A1(n9882), .A2(n6738), .ZN(n9677) );
  OAI211_X1 U10611 ( .C1(n9854), .C2(n9678), .A(n9885), .B(n9677), .ZN(n9679)
         );
  NAND2_X1 U10612 ( .A1(n9679), .A2(n10524), .ZN(n9680) );
  OAI211_X1 U10613 ( .C1(n9886), .C2(n9836), .A(n9681), .B(n9680), .ZN(
        P1_U3268) );
  INV_X1 U10614 ( .A(n9682), .ZN(n9683) );
  AOI21_X1 U10615 ( .B1(n9685), .B2(n9684), .A(n9683), .ZN(n9889) );
  INV_X1 U10616 ( .A(n9889), .ZN(n9701) );
  NAND2_X1 U10617 ( .A1(n9686), .A2(n6678), .ZN(n9687) );
  NAND3_X1 U10618 ( .A1(n9688), .A2(n10546), .A3(n9687), .ZN(n9691) );
  AOI22_X1 U10619 ( .A1(n9689), .A2(n10543), .B1(n10541), .B2(n9726), .ZN(
        n9690) );
  NAND2_X1 U10620 ( .A1(n9691), .A2(n9690), .ZN(n9887) );
  INV_X1 U10621 ( .A(n9710), .ZN(n9694) );
  INV_X1 U10622 ( .A(n9692), .ZN(n9693) );
  AOI211_X1 U10623 ( .C1(n9695), .C2(n9694), .A(n9797), .B(n9693), .ZN(n9888)
         );
  NAND2_X1 U10624 ( .A1(n9888), .A2(n4924), .ZN(n9698) );
  AOI22_X1 U10625 ( .A1(n9696), .A2(n10554), .B1(P1_REG2_REG_24__SCAN_IN), 
        .B2(n9800), .ZN(n9697) );
  OAI211_X1 U10626 ( .C1(n9968), .C2(n9802), .A(n9698), .B(n9697), .ZN(n9699)
         );
  AOI21_X1 U10627 ( .B1(n10524), .B2(n9887), .A(n9699), .ZN(n9700) );
  OAI21_X1 U10628 ( .B1(n9701), .B2(n9836), .A(n9700), .ZN(P1_U3269) );
  XOR2_X1 U10629 ( .A(n9702), .B(n9703), .Z(n9894) );
  INV_X1 U10630 ( .A(n9894), .ZN(n9718) );
  XNOR2_X1 U10631 ( .A(n9704), .B(n9703), .ZN(n9705) );
  NAND2_X1 U10632 ( .A1(n9705), .A2(n10546), .ZN(n9709) );
  AOI22_X1 U10633 ( .A1(n9707), .A2(n10543), .B1(n9821), .B2(n9706), .ZN(n9708) );
  NAND2_X1 U10634 ( .A1(n9709), .A2(n9708), .ZN(n9892) );
  AOI211_X1 U10635 ( .C1(n9711), .C2(n9719), .A(n9797), .B(n9710), .ZN(n9893)
         );
  NAND2_X1 U10636 ( .A1(n9893), .A2(n4924), .ZN(n9715) );
  INV_X1 U10637 ( .A(n9712), .ZN(n9713) );
  AOI22_X1 U10638 ( .A1(n9713), .A2(n10554), .B1(P1_REG2_REG_23__SCAN_IN), 
        .B2(n10555), .ZN(n9714) );
  OAI211_X1 U10639 ( .C1(n9972), .C2(n9802), .A(n9715), .B(n9714), .ZN(n9716)
         );
  AOI21_X1 U10640 ( .B1(n10524), .B2(n9892), .A(n9716), .ZN(n9717) );
  OAI21_X1 U10641 ( .B1(n9718), .B2(n9836), .A(n9717), .ZN(P1_U3270) );
  INV_X1 U10642 ( .A(n9719), .ZN(n9720) );
  AOI211_X1 U10643 ( .C1(n9721), .C2(n9749), .A(n9797), .B(n9720), .ZN(n9898)
         );
  OAI21_X1 U10644 ( .B1(n9724), .B2(n9723), .A(n9722), .ZN(n9727) );
  AOI222_X1 U10645 ( .A1(n10546), .A2(n9727), .B1(n9726), .B2(n10543), .C1(
        n9725), .C2(n10541), .ZN(n9728) );
  INV_X1 U10646 ( .A(n9728), .ZN(n9897) );
  AOI21_X1 U10647 ( .B1(n9898), .B2(n6738), .A(n9897), .ZN(n9737) );
  OAI21_X1 U10648 ( .B1(n4957), .B2(n9731), .A(n9730), .ZN(n9899) );
  INV_X1 U10649 ( .A(n9732), .ZN(n9733) );
  AOI22_X1 U10650 ( .A1(n9733), .A2(n10554), .B1(P1_REG2_REG_22__SCAN_IN), 
        .B2(n9800), .ZN(n9734) );
  OAI21_X1 U10651 ( .B1(n9976), .B2(n9802), .A(n9734), .ZN(n9735) );
  AOI21_X1 U10652 ( .B1(n9899), .B2(n10559), .A(n9735), .ZN(n9736) );
  OAI21_X1 U10653 ( .B1(n10555), .B2(n9737), .A(n9736), .ZN(P1_U3271) );
  NAND2_X1 U10654 ( .A1(n9739), .A2(n9738), .ZN(n9740) );
  XOR2_X1 U10655 ( .A(n9747), .B(n9740), .Z(n9741) );
  OAI222_X1 U10656 ( .A1(n9764), .A2(n9743), .B1(n9762), .B2(n9742), .C1(n9741), .C2(n9759), .ZN(n9902) );
  INV_X1 U10657 ( .A(n9902), .ZN(n9755) );
  INV_X1 U10658 ( .A(n9744), .ZN(n9745) );
  AOI21_X1 U10659 ( .B1(n9747), .B2(n9746), .A(n9745), .ZN(n9904) );
  OR2_X1 U10660 ( .A1(n9980), .A2(n5002), .ZN(n9748) );
  AND3_X1 U10661 ( .A1(n9749), .A2(n9748), .A3(n10537), .ZN(n9903) );
  NAND2_X1 U10662 ( .A1(n9903), .A2(n4924), .ZN(n9752) );
  AOI22_X1 U10663 ( .A1(n9750), .A2(n10554), .B1(P1_REG2_REG_21__SCAN_IN), 
        .B2(n10555), .ZN(n9751) );
  OAI211_X1 U10664 ( .C1(n9980), .C2(n9802), .A(n9752), .B(n9751), .ZN(n9753)
         );
  AOI21_X1 U10665 ( .B1(n9904), .B2(n10559), .A(n9753), .ZN(n9754) );
  OAI21_X1 U10666 ( .B1(n10555), .B2(n9755), .A(n9754), .ZN(P1_U3272) );
  XNOR2_X1 U10667 ( .A(n9756), .B(n9757), .ZN(n9911) );
  XNOR2_X1 U10668 ( .A(n9758), .B(n9757), .ZN(n9760) );
  OAI222_X1 U10669 ( .A1(n9764), .A2(n9763), .B1(n9762), .B2(n9761), .C1(n9760), .C2(n9759), .ZN(n9907) );
  AOI211_X1 U10670 ( .C1(n9909), .C2(n9782), .A(n9797), .B(n5002), .ZN(n9908)
         );
  NAND2_X1 U10671 ( .A1(n9908), .A2(n4924), .ZN(n9768) );
  INV_X1 U10672 ( .A(n9765), .ZN(n9766) );
  AOI22_X1 U10673 ( .A1(n9800), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9766), .B2(
        n10554), .ZN(n9767) );
  OAI211_X1 U10674 ( .C1(n5360), .C2(n9802), .A(n9768), .B(n9767), .ZN(n9769)
         );
  AOI21_X1 U10675 ( .B1(n9907), .B2(n10524), .A(n9769), .ZN(n9770) );
  OAI21_X1 U10676 ( .B1(n9911), .B2(n9836), .A(n9770), .ZN(P1_U3273) );
  NAND2_X1 U10677 ( .A1(n9804), .A2(n9771), .ZN(n9772) );
  NAND2_X1 U10678 ( .A1(n9772), .A2(n9780), .ZN(n9774) );
  NAND2_X1 U10679 ( .A1(n9774), .A2(n9773), .ZN(n9775) );
  NAND2_X1 U10680 ( .A1(n9775), .A2(n10546), .ZN(n9779) );
  AOI22_X1 U10681 ( .A1(n9777), .A2(n10543), .B1(n9776), .B2(n9821), .ZN(n9778) );
  NAND2_X1 U10682 ( .A1(n9779), .A2(n9778), .ZN(n9912) );
  INV_X1 U10683 ( .A(n9912), .ZN(n9790) );
  XOR2_X1 U10684 ( .A(n9781), .B(n9780), .Z(n9914) );
  NAND2_X1 U10685 ( .A1(n9914), .A2(n10559), .ZN(n9789) );
  INV_X1 U10686 ( .A(n9782), .ZN(n9783) );
  AOI211_X1 U10687 ( .C1(n9784), .C2(n9795), .A(n9797), .B(n9783), .ZN(n9913)
         );
  INV_X1 U10688 ( .A(n9784), .ZN(n9985) );
  NOR2_X1 U10689 ( .A1(n9985), .A2(n9802), .ZN(n9787) );
  OAI22_X1 U10690 ( .A1(n10524), .A2(n9600), .B1(n9785), .B2(n9854), .ZN(n9786) );
  AOI211_X1 U10691 ( .C1(n9913), .C2(n4924), .A(n9787), .B(n9786), .ZN(n9788)
         );
  OAI211_X1 U10692 ( .C1(n10555), .C2(n9790), .A(n9789), .B(n9788), .ZN(
        P1_U3274) );
  OAI21_X1 U10693 ( .B1(n9793), .B2(n9792), .A(n9791), .ZN(n9917) );
  INV_X1 U10694 ( .A(n9794), .ZN(n9798) );
  INV_X1 U10695 ( .A(n9795), .ZN(n9796) );
  AOI211_X1 U10696 ( .C1(n5362), .C2(n9798), .A(n9797), .B(n9796), .ZN(n9919)
         );
  AOI22_X1 U10697 ( .A1(n9800), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9799), .B2(
        n10554), .ZN(n9801) );
  OAI21_X1 U10698 ( .B1(n9989), .B2(n9802), .A(n9801), .ZN(n9803) );
  AOI21_X1 U10699 ( .B1(n9919), .B2(n4924), .A(n9803), .ZN(n9811) );
  OAI211_X1 U10700 ( .C1(n9806), .C2(n9805), .A(n9804), .B(n10546), .ZN(n9809)
         );
  AOI22_X1 U10701 ( .A1(n9807), .A2(n10543), .B1(n9821), .B2(n9819), .ZN(n9808) );
  NAND2_X1 U10702 ( .A1(n9809), .A2(n9808), .ZN(n9918) );
  NAND2_X1 U10703 ( .A1(n9918), .A2(n10524), .ZN(n9810) );
  OAI211_X1 U10704 ( .C1(n9917), .C2(n9836), .A(n9811), .B(n9810), .ZN(
        P1_U3275) );
  INV_X1 U10705 ( .A(n9812), .ZN(n9815) );
  INV_X1 U10706 ( .A(n9813), .ZN(n9814) );
  OAI21_X1 U10707 ( .B1(n9815), .B2(n9814), .A(n9834), .ZN(n9816) );
  OAI211_X1 U10708 ( .C1(n9818), .C2(n9817), .A(n9816), .B(n10546), .ZN(n9823)
         );
  AOI22_X1 U10709 ( .A1(n9821), .A2(n9820), .B1(n9819), .B2(n10543), .ZN(n9822) );
  NAND2_X1 U10710 ( .A1(n9823), .A2(n9822), .ZN(n9930) );
  OAI211_X1 U10711 ( .C1(n9825), .C2(n9994), .A(n10537), .B(n9824), .ZN(n9928)
         );
  INV_X1 U10712 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n9828) );
  INV_X1 U10713 ( .A(n9826), .ZN(n9827) );
  OAI22_X1 U10714 ( .A1(n10524), .A2(n9828), .B1(n9827), .B2(n9854), .ZN(n9829) );
  AOI21_X1 U10715 ( .B1(n9830), .B2(n10552), .A(n9829), .ZN(n9831) );
  OAI21_X1 U10716 ( .B1(n9928), .B2(n9832), .A(n9831), .ZN(n9838) );
  OAI21_X1 U10717 ( .B1(n9835), .B2(n9834), .A(n9833), .ZN(n9929) );
  NOR2_X1 U10718 ( .A1(n9929), .A2(n9836), .ZN(n9837) );
  AOI211_X1 U10719 ( .C1(n10524), .C2(n9930), .A(n9838), .B(n9837), .ZN(n9839)
         );
  INV_X1 U10720 ( .A(n9839), .ZN(P1_U3277) );
  NAND2_X1 U10721 ( .A1(n9840), .A2(n10524), .ZN(n9851) );
  NAND2_X1 U10722 ( .A1(n9841), .A2(n10559), .ZN(n9850) );
  INV_X1 U10723 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n9844) );
  INV_X1 U10724 ( .A(n9842), .ZN(n9843) );
  OAI22_X1 U10725 ( .A1(n10524), .A2(n9844), .B1(n9843), .B2(n9854), .ZN(n9845) );
  AOI21_X1 U10726 ( .B1(n9846), .B2(n10552), .A(n9845), .ZN(n9849) );
  NAND2_X1 U10727 ( .A1(n9847), .A2(n4924), .ZN(n9848) );
  NAND4_X1 U10728 ( .A1(n9851), .A2(n9850), .A3(n9849), .A4(n9848), .ZN(
        P1_U3280) );
  NAND2_X1 U10729 ( .A1(n9852), .A2(n10559), .ZN(n9864) );
  INV_X1 U10730 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n9856) );
  INV_X1 U10731 ( .A(n9853), .ZN(n9855) );
  OAI22_X1 U10732 ( .A1(n10524), .A2(n9856), .B1(n9855), .B2(n9854), .ZN(n9857) );
  AOI21_X1 U10733 ( .B1(n9858), .B2(n10552), .A(n9857), .ZN(n9863) );
  NAND2_X1 U10734 ( .A1(n9859), .A2(n10524), .ZN(n9862) );
  NAND2_X1 U10735 ( .A1(n9860), .A2(n4924), .ZN(n9861) );
  NAND4_X1 U10736 ( .A1(n9864), .A2(n9863), .A3(n9862), .A4(n9861), .ZN(
        P1_U3282) );
  INV_X1 U10737 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9866) );
  NOR2_X1 U10738 ( .A1(n9865), .A2(n9868), .ZN(n9948) );
  MUX2_X1 U10739 ( .A(n9866), .B(n9948), .S(n10677), .Z(n9867) );
  OAI21_X1 U10740 ( .B1(n9951), .B2(n9934), .A(n9867), .ZN(P1_U3553) );
  INV_X1 U10741 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9870) );
  NOR2_X1 U10742 ( .A1(n9869), .A2(n9868), .ZN(n9952) );
  MUX2_X1 U10743 ( .A(n9870), .B(n9952), .S(n10677), .Z(n9871) );
  OAI21_X1 U10744 ( .B1(n9955), .B2(n9934), .A(n9871), .ZN(P1_U3552) );
  AOI211_X1 U10745 ( .C1(n9874), .C2(n10675), .A(n9873), .B(n9872), .ZN(n9956)
         );
  MUX2_X1 U10746 ( .A(n9875), .B(n9956), .S(n10677), .Z(n9876) );
  OAI21_X1 U10747 ( .B1(n9959), .B2(n9934), .A(n9876), .ZN(P1_U3549) );
  AOI211_X1 U10748 ( .C1(n9879), .C2(n10675), .A(n9878), .B(n9877), .ZN(n9960)
         );
  MUX2_X1 U10749 ( .A(n9880), .B(n9960), .S(n10677), .Z(n9881) );
  OAI21_X1 U10750 ( .B1(n9963), .B2(n9934), .A(n9881), .ZN(P1_U3548) );
  AOI21_X1 U10751 ( .B1(n10610), .B2(n9883), .A(n9882), .ZN(n9884) );
  OAI211_X1 U10752 ( .C1(n9886), .C2(n9937), .A(n9885), .B(n9884), .ZN(n9964)
         );
  MUX2_X1 U10753 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9964), .S(n10677), .Z(
        P1_U3547) );
  AOI211_X1 U10754 ( .C1(n9889), .C2(n10675), .A(n9888), .B(n9887), .ZN(n9965)
         );
  MUX2_X1 U10755 ( .A(n9890), .B(n9965), .S(n10677), .Z(n9891) );
  OAI21_X1 U10756 ( .B1(n9968), .B2(n9934), .A(n9891), .ZN(P1_U3546) );
  AOI211_X1 U10757 ( .C1(n9894), .C2(n10675), .A(n9893), .B(n9892), .ZN(n9969)
         );
  MUX2_X1 U10758 ( .A(n9895), .B(n9969), .S(n10677), .Z(n9896) );
  OAI21_X1 U10759 ( .B1(n9972), .B2(n9934), .A(n9896), .ZN(P1_U3545) );
  AOI211_X1 U10760 ( .C1(n9899), .C2(n10675), .A(n9898), .B(n9897), .ZN(n9973)
         );
  MUX2_X1 U10761 ( .A(n9900), .B(n9973), .S(n10677), .Z(n9901) );
  OAI21_X1 U10762 ( .B1(n9976), .B2(n9934), .A(n9901), .ZN(P1_U3544) );
  AOI211_X1 U10763 ( .C1(n9904), .C2(n10675), .A(n9903), .B(n9902), .ZN(n9977)
         );
  MUX2_X1 U10764 ( .A(n9905), .B(n9977), .S(n10677), .Z(n9906) );
  OAI21_X1 U10765 ( .B1(n9980), .B2(n9934), .A(n9906), .ZN(P1_U3543) );
  AOI211_X1 U10766 ( .C1(n10610), .C2(n9909), .A(n9908), .B(n9907), .ZN(n9910)
         );
  OAI21_X1 U10767 ( .B1(n9937), .B2(n9911), .A(n9910), .ZN(n9981) );
  MUX2_X1 U10768 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9981), .S(n10677), .Z(
        P1_U3542) );
  AOI211_X1 U10769 ( .C1(n9914), .C2(n10675), .A(n9913), .B(n9912), .ZN(n9982)
         );
  MUX2_X1 U10770 ( .A(n9915), .B(n9982), .S(n10677), .Z(n9916) );
  OAI21_X1 U10771 ( .B1(n9985), .B2(n9934), .A(n9916), .ZN(P1_U3541) );
  INV_X1 U10772 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9921) );
  INV_X1 U10773 ( .A(n9917), .ZN(n9920) );
  AOI211_X1 U10774 ( .C1(n9920), .C2(n10675), .A(n9919), .B(n9918), .ZN(n9986)
         );
  MUX2_X1 U10775 ( .A(n9921), .B(n9986), .S(n10677), .Z(n9922) );
  OAI21_X1 U10776 ( .B1(n9989), .B2(n9934), .A(n9922), .ZN(P1_U3540) );
  AOI211_X1 U10777 ( .C1(n10610), .C2(n9925), .A(n9924), .B(n9923), .ZN(n9926)
         );
  OAI21_X1 U10778 ( .B1(n9927), .B2(n9937), .A(n9926), .ZN(n9990) );
  MUX2_X1 U10779 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9990), .S(n10677), .Z(
        P1_U3539) );
  OAI21_X1 U10780 ( .B1(n9929), .B2(n9937), .A(n9928), .ZN(n9931) );
  NOR2_X1 U10781 ( .A1(n9931), .A2(n9930), .ZN(n9991) );
  MUX2_X1 U10782 ( .A(n9932), .B(n9991), .S(n10677), .Z(n9933) );
  OAI21_X1 U10783 ( .B1(n9994), .B2(n9934), .A(n9933), .ZN(P1_U3538) );
  OAI211_X1 U10784 ( .C1(n9938), .C2(n9937), .A(n9936), .B(n9935), .ZN(n9996)
         );
  MUX2_X1 U10785 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n9996), .S(n10677), .Z(
        n9939) );
  AOI21_X1 U10786 ( .B1(n9940), .B2(n9998), .A(n9939), .ZN(n9941) );
  INV_X1 U10787 ( .A(n9941), .ZN(P1_U3537) );
  NAND2_X1 U10788 ( .A1(n9942), .A2(n10675), .ZN(n9947) );
  NAND2_X1 U10789 ( .A1(n9943), .A2(n10610), .ZN(n9944) );
  NAND4_X1 U10790 ( .A1(n9947), .A2(n9946), .A3(n9945), .A4(n9944), .ZN(n10000) );
  MUX2_X1 U10791 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n10000), .S(n10677), .Z(
        P1_U3536) );
  INV_X1 U10792 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n9949) );
  MUX2_X1 U10793 ( .A(n9949), .B(n9948), .S(n10681), .Z(n9950) );
  OAI21_X1 U10794 ( .B1(n9951), .B2(n9995), .A(n9950), .ZN(P1_U3521) );
  INV_X1 U10795 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9953) );
  MUX2_X1 U10796 ( .A(n9953), .B(n9952), .S(n10681), .Z(n9954) );
  OAI21_X1 U10797 ( .B1(n9955), .B2(n9995), .A(n9954), .ZN(P1_U3520) );
  INV_X1 U10798 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n9957) );
  MUX2_X1 U10799 ( .A(n9957), .B(n9956), .S(n10681), .Z(n9958) );
  OAI21_X1 U10800 ( .B1(n9959), .B2(n9995), .A(n9958), .ZN(P1_U3517) );
  INV_X1 U10801 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n9961) );
  MUX2_X1 U10802 ( .A(n9961), .B(n9960), .S(n10681), .Z(n9962) );
  OAI21_X1 U10803 ( .B1(n9963), .B2(n9995), .A(n9962), .ZN(P1_U3516) );
  MUX2_X1 U10804 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9964), .S(n10681), .Z(
        P1_U3515) );
  INV_X1 U10805 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n9966) );
  MUX2_X1 U10806 ( .A(n9966), .B(n9965), .S(n10681), .Z(n9967) );
  OAI21_X1 U10807 ( .B1(n9968), .B2(n9995), .A(n9967), .ZN(P1_U3514) );
  INV_X1 U10808 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n9970) );
  MUX2_X1 U10809 ( .A(n9970), .B(n9969), .S(n10681), .Z(n9971) );
  OAI21_X1 U10810 ( .B1(n9972), .B2(n9995), .A(n9971), .ZN(P1_U3513) );
  INV_X1 U10811 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n9974) );
  MUX2_X1 U10812 ( .A(n9974), .B(n9973), .S(n10681), .Z(n9975) );
  OAI21_X1 U10813 ( .B1(n9976), .B2(n9995), .A(n9975), .ZN(P1_U3512) );
  INV_X1 U10814 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n9978) );
  MUX2_X1 U10815 ( .A(n9978), .B(n9977), .S(n10681), .Z(n9979) );
  OAI21_X1 U10816 ( .B1(n9980), .B2(n9995), .A(n9979), .ZN(P1_U3511) );
  MUX2_X1 U10817 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9981), .S(n10681), .Z(
        P1_U3510) );
  INV_X1 U10818 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n9983) );
  MUX2_X1 U10819 ( .A(n9983), .B(n9982), .S(n10681), .Z(n9984) );
  OAI21_X1 U10820 ( .B1(n9985), .B2(n9995), .A(n9984), .ZN(P1_U3509) );
  INV_X1 U10821 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n9987) );
  MUX2_X1 U10822 ( .A(n9987), .B(n9986), .S(n10681), .Z(n9988) );
  OAI21_X1 U10823 ( .B1(n9989), .B2(n9995), .A(n9988), .ZN(P1_U3507) );
  MUX2_X1 U10824 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9990), .S(n10681), .Z(
        P1_U3504) );
  INV_X1 U10825 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n9992) );
  MUX2_X1 U10826 ( .A(n9992), .B(n9991), .S(n10681), .Z(n9993) );
  OAI21_X1 U10827 ( .B1(n9994), .B2(n9995), .A(n9993), .ZN(P1_U3501) );
  MUX2_X1 U10828 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n9996), .S(n10681), .Z(
        n9997) );
  AOI21_X1 U10829 ( .B1(n6798), .B2(n9998), .A(n9997), .ZN(n9999) );
  INV_X1 U10830 ( .A(n9999), .ZN(P1_U3498) );
  MUX2_X1 U10831 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n10000), .S(n10681), .Z(
        P1_U3495) );
  NOR4_X1 U10832 ( .A1(n10001), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3086), 
        .A4(n6509), .ZN(n10002) );
  AOI21_X1 U10833 ( .B1(n10003), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n10002), 
        .ZN(n10004) );
  OAI21_X1 U10834 ( .B1(n10005), .B2(n7945), .A(n10004), .ZN(P1_U3324) );
  AOI22_X1 U10835 ( .A1(n10006), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n10012), .ZN(n10007) );
  OAI21_X1 U10836 ( .B1(n10008), .B2(n7945), .A(n10007), .ZN(P1_U3325) );
  AOI22_X1 U10837 ( .A1(n10009), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n10012), .ZN(n10010) );
  OAI21_X1 U10838 ( .B1(n10011), .B2(n7945), .A(n10010), .ZN(P1_U3326) );
  AOI22_X1 U10839 ( .A1(n10013), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n10012), .ZN(n10014) );
  OAI21_X1 U10840 ( .B1(n10015), .B2(n7945), .A(n10014), .ZN(P1_U3327) );
  INV_X1 U10841 ( .A(n10016), .ZN(n10017) );
  MUX2_X1 U10842 ( .A(n10017), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  AND2_X1 U10843 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n10018), .ZN(P1_U3323) );
  AND2_X1 U10844 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n10018), .ZN(P1_U3322) );
  AND2_X1 U10845 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n10018), .ZN(P1_U3321) );
  AND2_X1 U10846 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n10018), .ZN(P1_U3320) );
  AND2_X1 U10847 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n10018), .ZN(P1_U3319) );
  AND2_X1 U10848 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n10018), .ZN(P1_U3318) );
  AND2_X1 U10849 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n10018), .ZN(P1_U3317) );
  AND2_X1 U10850 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n10018), .ZN(P1_U3316) );
  AND2_X1 U10851 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n10018), .ZN(P1_U3315) );
  AND2_X1 U10852 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n10018), .ZN(P1_U3314) );
  AND2_X1 U10853 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n10018), .ZN(P1_U3313) );
  AND2_X1 U10854 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n10018), .ZN(P1_U3312) );
  AND2_X1 U10855 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n10018), .ZN(P1_U3311) );
  AND2_X1 U10856 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n10018), .ZN(P1_U3310) );
  AND2_X1 U10857 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n10018), .ZN(P1_U3309) );
  AND2_X1 U10858 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n10018), .ZN(P1_U3308) );
  AND2_X1 U10859 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n10018), .ZN(P1_U3307) );
  AND2_X1 U10860 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n10018), .ZN(P1_U3306) );
  AND2_X1 U10861 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n10018), .ZN(P1_U3305) );
  AND2_X1 U10862 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n10018), .ZN(P1_U3304) );
  AND2_X1 U10863 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n10018), .ZN(P1_U3303) );
  AND2_X1 U10864 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n10018), .ZN(P1_U3302) );
  AND2_X1 U10865 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n10018), .ZN(P1_U3301) );
  AND2_X1 U10866 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n10018), .ZN(P1_U3300) );
  AND2_X1 U10867 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n10018), .ZN(P1_U3299) );
  AND2_X1 U10868 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n10018), .ZN(P1_U3298) );
  AND2_X1 U10869 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n10018), .ZN(P1_U3297) );
  AND2_X1 U10870 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n10018), .ZN(P1_U3296) );
  AND2_X1 U10871 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n10018), .ZN(P1_U3295) );
  AND2_X1 U10872 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n10018), .ZN(P1_U3294) );
  INV_X1 U10873 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n10109) );
  INV_X1 U10874 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n10211) );
  OAI22_X1 U10875 ( .A1(n10211), .A2(keyinput_126), .B1(
        P2_REG3_REG_15__SCAN_IN), .B2(keyinput_127), .ZN(n10019) );
  AOI221_X1 U10876 ( .B1(n10211), .B2(keyinput_126), .C1(keyinput_127), .C2(
        P2_REG3_REG_15__SCAN_IN), .A(n10019), .ZN(n10107) );
  OAI22_X1 U10877 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(keyinput_124), .B1(
        keyinput_122), .B2(P2_REG3_REG_11__SCAN_IN), .ZN(n10020) );
  AOI221_X1 U10878 ( .B1(P2_REG3_REG_18__SCAN_IN), .B2(keyinput_124), .C1(
        P2_REG3_REG_11__SCAN_IN), .C2(keyinput_122), .A(n10020), .ZN(n10105)
         );
  OAI22_X1 U10879 ( .A1(P2_REG3_REG_20__SCAN_IN), .A2(keyinput_119), .B1(
        P2_REG3_REG_13__SCAN_IN), .B2(keyinput_120), .ZN(n10021) );
  AOI221_X1 U10880 ( .B1(P2_REG3_REG_20__SCAN_IN), .B2(keyinput_119), .C1(
        keyinput_120), .C2(P2_REG3_REG_13__SCAN_IN), .A(n10021), .ZN(n10104)
         );
  OAI22_X1 U10881 ( .A1(n10205), .A2(keyinput_121), .B1(n7300), .B2(
        keyinput_123), .ZN(n10022) );
  AOI221_X1 U10882 ( .B1(n10205), .B2(keyinput_121), .C1(keyinput_123), .C2(
        n7300), .A(n10022), .ZN(n10103) );
  INV_X1 U10883 ( .A(keyinput_118), .ZN(n10101) );
  INV_X1 U10884 ( .A(keyinput_117), .ZN(n10099) );
  INV_X1 U10885 ( .A(keyinput_116), .ZN(n10097) );
  OAI22_X1 U10886 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(keyinput_110), .B1(
        keyinput_108), .B2(P2_REG3_REG_1__SCAN_IN), .ZN(n10023) );
  AOI221_X1 U10887 ( .B1(P2_REG3_REG_12__SCAN_IN), .B2(keyinput_110), .C1(
        P2_REG3_REG_1__SCAN_IN), .C2(keyinput_108), .A(n10023), .ZN(n10087) );
  OAI22_X1 U10888 ( .A1(P2_STATE_REG_SCAN_IN), .A2(keyinput_98), .B1(
        P2_REG3_REG_7__SCAN_IN), .B2(keyinput_99), .ZN(n10024) );
  AOI221_X1 U10889 ( .B1(P2_STATE_REG_SCAN_IN), .B2(keyinput_98), .C1(
        keyinput_99), .C2(P2_REG3_REG_7__SCAN_IN), .A(n10024), .ZN(n10074) );
  OAI22_X1 U10890 ( .A1(SI_10_), .A2(keyinput_86), .B1(SI_9_), .B2(keyinput_87), .ZN(n10025) );
  AOI221_X1 U10891 ( .B1(SI_10_), .B2(keyinput_86), .C1(keyinput_87), .C2(
        SI_9_), .A(n10025), .ZN(n10055) );
  AOI22_X1 U10892 ( .A1(n10140), .A2(keyinput_80), .B1(keyinput_82), .B2(
        n10139), .ZN(n10026) );
  OAI221_X1 U10893 ( .B1(n10140), .B2(keyinput_80), .C1(n10139), .C2(
        keyinput_82), .A(n10026), .ZN(n10053) );
  AOI22_X1 U10894 ( .A1(SI_18_), .A2(keyinput_78), .B1(n10129), .B2(
        keyinput_77), .ZN(n10027) );
  OAI221_X1 U10895 ( .B1(SI_18_), .B2(keyinput_78), .C1(n10129), .C2(
        keyinput_77), .A(n10027), .ZN(n10046) );
  OAI22_X1 U10896 ( .A1(SI_21_), .A2(keyinput_75), .B1(SI_20_), .B2(
        keyinput_76), .ZN(n10028) );
  AOI221_X1 U10897 ( .B1(SI_21_), .B2(keyinput_75), .C1(keyinput_76), .C2(
        SI_20_), .A(n10028), .ZN(n10045) );
  AOI22_X1 U10898 ( .A1(SI_29_), .A2(keyinput_67), .B1(SI_27_), .B2(
        keyinput_69), .ZN(n10029) );
  OAI221_X1 U10899 ( .B1(SI_29_), .B2(keyinput_67), .C1(SI_27_), .C2(
        keyinput_69), .A(n10029), .ZN(n10040) );
  XOR2_X1 U10900 ( .A(SI_30_), .B(keyinput_66), .Z(n10034) );
  AOI22_X1 U10901 ( .A1(P2_WR_REG_SCAN_IN), .A2(keyinput_64), .B1(SI_31_), 
        .B2(keyinput_65), .ZN(n10030) );
  OAI221_X1 U10902 ( .B1(P2_WR_REG_SCAN_IN), .B2(keyinput_64), .C1(SI_31_), 
        .C2(keyinput_65), .A(n10030), .ZN(n10033) );
  OAI22_X1 U10903 ( .A1(SI_26_), .A2(keyinput_70), .B1(keyinput_68), .B2(
        SI_28_), .ZN(n10031) );
  AOI221_X1 U10904 ( .B1(SI_26_), .B2(keyinput_70), .C1(SI_28_), .C2(
        keyinput_68), .A(n10031), .ZN(n10032) );
  OAI21_X1 U10905 ( .B1(n10034), .B2(n10033), .A(n10032), .ZN(n10039) );
  OAI22_X1 U10906 ( .A1(n10121), .A2(keyinput_74), .B1(keyinput_72), .B2(
        SI_24_), .ZN(n10035) );
  AOI221_X1 U10907 ( .B1(n10121), .B2(keyinput_74), .C1(SI_24_), .C2(
        keyinput_72), .A(n10035), .ZN(n10038) );
  OAI22_X1 U10908 ( .A1(SI_25_), .A2(keyinput_71), .B1(keyinput_73), .B2(
        SI_23_), .ZN(n10036) );
  AOI221_X1 U10909 ( .B1(SI_25_), .B2(keyinput_71), .C1(SI_23_), .C2(
        keyinput_73), .A(n10036), .ZN(n10037) );
  OAI211_X1 U10910 ( .C1(n10040), .C2(n10039), .A(n10038), .B(n10037), .ZN(
        n10044) );
  OAI22_X1 U10911 ( .A1(n10133), .A2(keyinput_79), .B1(n10042), .B2(
        keyinput_81), .ZN(n10041) );
  AOI221_X1 U10912 ( .B1(n10133), .B2(keyinput_79), .C1(keyinput_81), .C2(
        n10042), .A(n10041), .ZN(n10043) );
  OAI221_X1 U10913 ( .B1(n10046), .B2(n10045), .C1(n10046), .C2(n10044), .A(
        n10043), .ZN(n10052) );
  INV_X1 U10914 ( .A(SI_13_), .ZN(n10049) );
  OAI22_X1 U10915 ( .A1(n10049), .A2(keyinput_83), .B1(n10048), .B2(
        keyinput_84), .ZN(n10047) );
  AOI221_X1 U10916 ( .B1(n10049), .B2(keyinput_83), .C1(keyinput_84), .C2(
        n10048), .A(n10047), .ZN(n10051) );
  XNOR2_X1 U10917 ( .A(SI_11_), .B(keyinput_85), .ZN(n10050) );
  OAI211_X1 U10918 ( .C1(n10053), .C2(n10052), .A(n10051), .B(n10050), .ZN(
        n10054) );
  AOI22_X1 U10919 ( .A1(SI_8_), .A2(keyinput_88), .B1(n10055), .B2(n10054), 
        .ZN(n10058) );
  AOI22_X1 U10920 ( .A1(SI_7_), .A2(keyinput_89), .B1(n5839), .B2(keyinput_91), 
        .ZN(n10056) );
  OAI221_X1 U10921 ( .B1(SI_7_), .B2(keyinput_89), .C1(n5839), .C2(keyinput_91), .A(n10056), .ZN(n10057) );
  AOI221_X1 U10922 ( .B1(SI_8_), .B2(n10058), .C1(keyinput_88), .C2(n10058), 
        .A(n10057), .ZN(n10061) );
  XNOR2_X1 U10923 ( .A(SI_4_), .B(keyinput_92), .ZN(n10060) );
  XNOR2_X1 U10924 ( .A(SI_6_), .B(keyinput_90), .ZN(n10059) );
  NAND3_X1 U10925 ( .A1(n10061), .A2(n10060), .A3(n10059), .ZN(n10064) );
  XNOR2_X1 U10926 ( .A(n10062), .B(keyinput_93), .ZN(n10063) );
  NAND2_X1 U10927 ( .A1(n10064), .A2(n10063), .ZN(n10070) );
  INV_X1 U10928 ( .A(keyinput_94), .ZN(n10065) );
  MUX2_X1 U10929 ( .A(keyinput_94), .B(n10065), .S(SI_2_), .Z(n10069) );
  XNOR2_X1 U10930 ( .A(n10066), .B(keyinput_95), .ZN(n10068) );
  XNOR2_X1 U10931 ( .A(SI_0_), .B(keyinput_96), .ZN(n10067) );
  AOI211_X1 U10932 ( .C1(n10070), .C2(n10069), .A(n10068), .B(n10067), .ZN(
        n10071) );
  AOI21_X1 U10933 ( .B1(P2_RD_REG_SCAN_IN), .B2(keyinput_97), .A(n10071), .ZN(
        n10072) );
  OAI21_X1 U10934 ( .B1(keyinput_97), .B2(P2_RD_REG_SCAN_IN), .A(n10072), .ZN(
        n10073) );
  AOI22_X1 U10935 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(keyinput_100), .B1(
        n10074), .B2(n10073), .ZN(n10077) );
  AOI22_X1 U10936 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(keyinput_101), .B1(
        P2_REG3_REG_23__SCAN_IN), .B2(keyinput_102), .ZN(n10075) );
  OAI221_X1 U10937 ( .B1(P2_REG3_REG_14__SCAN_IN), .B2(keyinput_101), .C1(
        P2_REG3_REG_23__SCAN_IN), .C2(keyinput_102), .A(n10075), .ZN(n10076)
         );
  AOI221_X1 U10938 ( .B1(P2_REG3_REG_27__SCAN_IN), .B2(n10077), .C1(
        keyinput_100), .C2(n10077), .A(n10076), .ZN(n10085) );
  INV_X1 U10939 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n10079) );
  AOI22_X1 U10940 ( .A1(n10080), .A2(keyinput_104), .B1(n10079), .B2(
        keyinput_103), .ZN(n10078) );
  OAI221_X1 U10941 ( .B1(n10080), .B2(keyinput_104), .C1(n10079), .C2(
        keyinput_103), .A(n10078), .ZN(n10084) );
  OAI22_X1 U10942 ( .A1(n5872), .A2(keyinput_107), .B1(P2_REG3_REG_19__SCAN_IN), .B2(keyinput_105), .ZN(n10081) );
  AOI221_X1 U10943 ( .B1(n5872), .B2(keyinput_107), .C1(keyinput_105), .C2(
        P2_REG3_REG_19__SCAN_IN), .A(n10081), .ZN(n10083) );
  XNOR2_X1 U10944 ( .A(P2_REG3_REG_28__SCAN_IN), .B(keyinput_106), .ZN(n10082)
         );
  OAI211_X1 U10945 ( .C1(n10085), .C2(n10084), .A(n10083), .B(n10082), .ZN(
        n10086) );
  OAI211_X1 U10946 ( .C1(P2_REG3_REG_21__SCAN_IN), .C2(keyinput_109), .A(
        n10087), .B(n10086), .ZN(n10088) );
  AOI21_X1 U10947 ( .B1(P2_REG3_REG_21__SCAN_IN), .B2(keyinput_109), .A(n10088), .ZN(n10095) );
  XOR2_X1 U10948 ( .A(n10184), .B(keyinput_111), .Z(n10094) );
  OAI22_X1 U10949 ( .A1(n10090), .A2(keyinput_112), .B1(n5816), .B2(
        keyinput_113), .ZN(n10089) );
  AOI221_X1 U10950 ( .B1(n10090), .B2(keyinput_112), .C1(keyinput_113), .C2(
        n5816), .A(n10089), .ZN(n10093) );
  OAI22_X1 U10951 ( .A1(P2_REG3_REG_24__SCAN_IN), .A2(keyinput_115), .B1(
        keyinput_114), .B2(P2_REG3_REG_17__SCAN_IN), .ZN(n10091) );
  AOI221_X1 U10952 ( .B1(P2_REG3_REG_24__SCAN_IN), .B2(keyinput_115), .C1(
        P2_REG3_REG_17__SCAN_IN), .C2(keyinput_114), .A(n10091), .ZN(n10092)
         );
  OAI211_X1 U10953 ( .C1(n10095), .C2(n10094), .A(n10093), .B(n10092), .ZN(
        n10096) );
  OAI221_X1 U10954 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(keyinput_116), .C1(
        n10193), .C2(n10097), .A(n10096), .ZN(n10098) );
  OAI221_X1 U10955 ( .B1(P2_REG3_REG_9__SCAN_IN), .B2(keyinput_117), .C1(
        n10195), .C2(n10099), .A(n10098), .ZN(n10100) );
  OAI221_X1 U10956 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(n10101), .C1(n10198), 
        .C2(keyinput_118), .A(n10100), .ZN(n10102) );
  NAND4_X1 U10957 ( .A1(n10105), .A2(n10104), .A3(n10103), .A4(n10102), .ZN(
        n10106) );
  OAI211_X1 U10958 ( .C1(n10109), .C2(keyinput_125), .A(n10107), .B(n10106), 
        .ZN(n10108) );
  AOI21_X1 U10959 ( .B1(n10109), .B2(keyinput_125), .A(n10108), .ZN(n10216) );
  XOR2_X1 U10960 ( .A(keyinput_61), .B(P2_REG3_REG_6__SCAN_IN), .Z(n10215) );
  INV_X1 U10961 ( .A(keyinput_54), .ZN(n10199) );
  INV_X1 U10962 ( .A(keyinput_53), .ZN(n10196) );
  INV_X1 U10963 ( .A(keyinput_52), .ZN(n10192) );
  INV_X1 U10964 ( .A(keyinput_47), .ZN(n10185) );
  OAI22_X1 U10965 ( .A1(n7698), .A2(keyinput_44), .B1(keyinput_46), .B2(
        P2_REG3_REG_12__SCAN_IN), .ZN(n10110) );
  AOI221_X1 U10966 ( .B1(n7698), .B2(keyinput_44), .C1(P2_REG3_REG_12__SCAN_IN), .C2(keyinput_46), .A(n10110), .ZN(n10181) );
  OAI22_X1 U10967 ( .A1(P2_STATE_REG_SCAN_IN), .A2(keyinput_34), .B1(
        keyinput_35), .B2(P2_REG3_REG_7__SCAN_IN), .ZN(n10111) );
  AOI221_X1 U10968 ( .B1(P2_STATE_REG_SCAN_IN), .B2(keyinput_34), .C1(
        P2_REG3_REG_7__SCAN_IN), .C2(keyinput_35), .A(n10111), .ZN(n10170) );
  INV_X1 U10969 ( .A(SI_29_), .ZN(n10113) );
  OAI22_X1 U10970 ( .A1(n10113), .A2(keyinput_3), .B1(keyinput_4), .B2(SI_28_), 
        .ZN(n10112) );
  AOI221_X1 U10971 ( .B1(n10113), .B2(keyinput_3), .C1(SI_28_), .C2(keyinput_4), .A(n10112), .ZN(n10127) );
  XOR2_X1 U10972 ( .A(SI_30_), .B(keyinput_2), .Z(n10118) );
  OAI22_X1 U10973 ( .A1(SI_31_), .A2(keyinput_1), .B1(P2_WR_REG_SCAN_IN), .B2(
        keyinput_0), .ZN(n10114) );
  AOI221_X1 U10974 ( .B1(SI_31_), .B2(keyinput_1), .C1(keyinput_0), .C2(
        P2_WR_REG_SCAN_IN), .A(n10114), .ZN(n10117) );
  AOI22_X1 U10975 ( .A1(SI_26_), .A2(keyinput_6), .B1(SI_27_), .B2(keyinput_5), 
        .ZN(n10115) );
  OAI221_X1 U10976 ( .B1(SI_26_), .B2(keyinput_6), .C1(SI_27_), .C2(keyinput_5), .A(n10115), .ZN(n10116) );
  AOI21_X1 U10977 ( .B1(n10118), .B2(n10117), .A(n10116), .ZN(n10126) );
  AOI22_X1 U10978 ( .A1(n10121), .A2(keyinput_10), .B1(n10120), .B2(keyinput_8), .ZN(n10119) );
  OAI221_X1 U10979 ( .B1(n10121), .B2(keyinput_10), .C1(n10120), .C2(
        keyinput_8), .A(n10119), .ZN(n10125) );
  AOI22_X1 U10980 ( .A1(SI_23_), .A2(keyinput_9), .B1(n10123), .B2(keyinput_7), 
        .ZN(n10122) );
  OAI221_X1 U10981 ( .B1(SI_23_), .B2(keyinput_9), .C1(n10123), .C2(keyinput_7), .A(n10122), .ZN(n10124) );
  AOI211_X1 U10982 ( .C1(n10127), .C2(n10126), .A(n10125), .B(n10124), .ZN(
        n10137) );
  OAI22_X1 U10983 ( .A1(n10129), .A2(keyinput_13), .B1(SI_18_), .B2(
        keyinput_14), .ZN(n10128) );
  AOI221_X1 U10984 ( .B1(n10129), .B2(keyinput_13), .C1(keyinput_14), .C2(
        SI_18_), .A(n10128), .ZN(n10136) );
  AOI22_X1 U10985 ( .A1(SI_21_), .A2(keyinput_11), .B1(n10131), .B2(
        keyinput_12), .ZN(n10130) );
  OAI221_X1 U10986 ( .B1(SI_21_), .B2(keyinput_11), .C1(n10131), .C2(
        keyinput_12), .A(n10130), .ZN(n10135) );
  AOI22_X1 U10987 ( .A1(SI_15_), .A2(keyinput_17), .B1(n10133), .B2(
        keyinput_15), .ZN(n10132) );
  OAI221_X1 U10988 ( .B1(SI_15_), .B2(keyinput_17), .C1(n10133), .C2(
        keyinput_15), .A(n10132), .ZN(n10134) );
  AOI221_X1 U10989 ( .B1(n10137), .B2(n10136), .C1(n10135), .C2(n10136), .A(
        n10134), .ZN(n10142) );
  OAI22_X1 U10990 ( .A1(n10140), .A2(keyinput_16), .B1(n10139), .B2(
        keyinput_18), .ZN(n10138) );
  AOI221_X1 U10991 ( .B1(n10140), .B2(keyinput_16), .C1(keyinput_18), .C2(
        n10139), .A(n10138), .ZN(n10141) );
  AOI22_X1 U10992 ( .A1(n10142), .A2(n10141), .B1(SI_11_), .B2(keyinput_21), 
        .ZN(n10143) );
  OAI21_X1 U10993 ( .B1(SI_11_), .B2(keyinput_21), .A(n10143), .ZN(n10149) );
  AOI22_X1 U10994 ( .A1(SI_12_), .A2(keyinput_20), .B1(SI_13_), .B2(
        keyinput_19), .ZN(n10144) );
  OAI221_X1 U10995 ( .B1(SI_12_), .B2(keyinput_20), .C1(SI_13_), .C2(
        keyinput_19), .A(n10144), .ZN(n10148) );
  OAI22_X1 U10996 ( .A1(n10146), .A2(keyinput_23), .B1(SI_10_), .B2(
        keyinput_22), .ZN(n10145) );
  AOI221_X1 U10997 ( .B1(n10146), .B2(keyinput_23), .C1(keyinput_22), .C2(
        SI_10_), .A(n10145), .ZN(n10147) );
  OAI21_X1 U10998 ( .B1(n10149), .B2(n10148), .A(n10147), .ZN(n10156) );
  XNOR2_X1 U10999 ( .A(SI_8_), .B(keyinput_24), .ZN(n10155) );
  AOI22_X1 U11000 ( .A1(SI_5_), .A2(keyinput_27), .B1(SI_7_), .B2(keyinput_25), 
        .ZN(n10150) );
  OAI221_X1 U11001 ( .B1(SI_5_), .B2(keyinput_27), .C1(SI_7_), .C2(keyinput_25), .A(n10150), .ZN(n10154) );
  XNOR2_X1 U11002 ( .A(SI_6_), .B(keyinput_26), .ZN(n10152) );
  XNOR2_X1 U11003 ( .A(SI_4_), .B(keyinput_28), .ZN(n10151) );
  NAND2_X1 U11004 ( .A1(n10152), .A2(n10151), .ZN(n10153) );
  AOI211_X1 U11005 ( .C1(n10156), .C2(n10155), .A(n10154), .B(n10153), .ZN(
        n10159) );
  INV_X1 U11006 ( .A(keyinput_29), .ZN(n10157) );
  MUX2_X1 U11007 ( .A(keyinput_29), .B(n10157), .S(SI_3_), .Z(n10158) );
  NOR2_X1 U11008 ( .A1(n10159), .A2(n10158), .ZN(n10166) );
  INV_X1 U11009 ( .A(keyinput_30), .ZN(n10160) );
  MUX2_X1 U11010 ( .A(keyinput_30), .B(n10160), .S(SI_2_), .Z(n10165) );
  AOI22_X1 U11011 ( .A1(SI_1_), .A2(keyinput_31), .B1(n10162), .B2(keyinput_32), .ZN(n10161) );
  OAI221_X1 U11012 ( .B1(SI_1_), .B2(keyinput_31), .C1(n10162), .C2(
        keyinput_32), .A(n10161), .ZN(n10163) );
  INV_X1 U11013 ( .A(n10163), .ZN(n10164) );
  OAI21_X1 U11014 ( .B1(n10166), .B2(n10165), .A(n10164), .ZN(n10168) );
  NAND2_X1 U11015 ( .A1(P2_RD_REG_SCAN_IN), .A2(keyinput_33), .ZN(n10167) );
  OAI211_X1 U11016 ( .C1(P2_RD_REG_SCAN_IN), .C2(keyinput_33), .A(n10168), .B(
        n10167), .ZN(n10169) );
  AOI22_X1 U11017 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(keyinput_36), .B1(n10170), .B2(n10169), .ZN(n10173) );
  AOI22_X1 U11018 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(keyinput_37), .B1(
        P2_REG3_REG_23__SCAN_IN), .B2(keyinput_38), .ZN(n10171) );
  OAI221_X1 U11019 ( .B1(P2_REG3_REG_14__SCAN_IN), .B2(keyinput_37), .C1(
        P2_REG3_REG_23__SCAN_IN), .C2(keyinput_38), .A(n10171), .ZN(n10172) );
  AOI221_X1 U11020 ( .B1(P2_REG3_REG_27__SCAN_IN), .B2(n10173), .C1(
        keyinput_36), .C2(n10173), .A(n10172), .ZN(n10179) );
  AOI22_X1 U11021 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(keyinput_40), .B1(
        P2_REG3_REG_10__SCAN_IN), .B2(keyinput_39), .ZN(n10174) );
  OAI221_X1 U11022 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(keyinput_40), .C1(
        P2_REG3_REG_10__SCAN_IN), .C2(keyinput_39), .A(n10174), .ZN(n10178) );
  OAI22_X1 U11023 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(keyinput_41), .B1(
        P2_REG3_REG_8__SCAN_IN), .B2(keyinput_43), .ZN(n10175) );
  AOI221_X1 U11024 ( .B1(P2_REG3_REG_19__SCAN_IN), .B2(keyinput_41), .C1(
        keyinput_43), .C2(P2_REG3_REG_8__SCAN_IN), .A(n10175), .ZN(n10177) );
  XNOR2_X1 U11025 ( .A(P2_REG3_REG_28__SCAN_IN), .B(keyinput_42), .ZN(n10176)
         );
  OAI211_X1 U11026 ( .C1(n10179), .C2(n10178), .A(n10177), .B(n10176), .ZN(
        n10180) );
  OAI211_X1 U11027 ( .C1(P2_REG3_REG_21__SCAN_IN), .C2(keyinput_45), .A(n10181), .B(n10180), .ZN(n10182) );
  AOI21_X1 U11028 ( .B1(P2_REG3_REG_21__SCAN_IN), .B2(keyinput_45), .A(n10182), 
        .ZN(n10183) );
  AOI221_X1 U11029 ( .B1(P2_REG3_REG_25__SCAN_IN), .B2(n10185), .C1(n10184), 
        .C2(keyinput_47), .A(n10183), .ZN(n10190) );
  AOI22_X1 U11030 ( .A1(P2_REG3_REG_24__SCAN_IN), .A2(keyinput_51), .B1(n8858), 
        .B2(keyinput_50), .ZN(n10186) );
  OAI221_X1 U11031 ( .B1(P2_REG3_REG_24__SCAN_IN), .B2(keyinput_51), .C1(n8858), .C2(keyinput_50), .A(n10186), .ZN(n10189) );
  AOI22_X1 U11032 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(keyinput_49), .B1(
        P2_REG3_REG_16__SCAN_IN), .B2(keyinput_48), .ZN(n10187) );
  OAI221_X1 U11033 ( .B1(P2_REG3_REG_5__SCAN_IN), .B2(keyinput_49), .C1(
        P2_REG3_REG_16__SCAN_IN), .C2(keyinput_48), .A(n10187), .ZN(n10188) );
  NOR3_X1 U11034 ( .A1(n10190), .A2(n10189), .A3(n10188), .ZN(n10191) );
  AOI221_X1 U11035 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(keyinput_52), .C1(n10193), .C2(n10192), .A(n10191), .ZN(n10194) );
  AOI221_X1 U11036 ( .B1(P2_REG3_REG_9__SCAN_IN), .B2(n10196), .C1(n10195), 
        .C2(keyinput_53), .A(n10194), .ZN(n10197) );
  AOI221_X1 U11037 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(n10199), .C1(n10198), 
        .C2(keyinput_54), .A(n10197), .ZN(n10209) );
  AOI22_X1 U11038 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(keyinput_56), .B1(
        P2_REG3_REG_18__SCAN_IN), .B2(keyinput_60), .ZN(n10200) );
  OAI221_X1 U11039 ( .B1(P2_REG3_REG_13__SCAN_IN), .B2(keyinput_56), .C1(
        P2_REG3_REG_18__SCAN_IN), .C2(keyinput_60), .A(n10200), .ZN(n10208) );
  INV_X1 U11040 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n10202) );
  AOI22_X1 U11041 ( .A1(n10203), .A2(keyinput_55), .B1(keyinput_58), .B2(
        n10202), .ZN(n10201) );
  OAI221_X1 U11042 ( .B1(n10203), .B2(keyinput_55), .C1(n10202), .C2(
        keyinput_58), .A(n10201), .ZN(n10207) );
  AOI22_X1 U11043 ( .A1(n10205), .A2(keyinput_57), .B1(keyinput_59), .B2(n7300), .ZN(n10204) );
  OAI221_X1 U11044 ( .B1(n10205), .B2(keyinput_57), .C1(n7300), .C2(
        keyinput_59), .A(n10204), .ZN(n10206) );
  NOR4_X1 U11045 ( .A1(n10209), .A2(n10208), .A3(n10207), .A4(n10206), .ZN(
        n10214) );
  AOI22_X1 U11046 ( .A1(n10212), .A2(keyinput_63), .B1(n10211), .B2(
        keyinput_62), .ZN(n10210) );
  OAI221_X1 U11047 ( .B1(n10212), .B2(keyinput_63), .C1(n10211), .C2(
        keyinput_62), .A(n10210), .ZN(n10213) );
  NOR4_X1 U11048 ( .A1(n10216), .A2(n10215), .A3(n10214), .A4(n10213), .ZN(
        n10220) );
  OAI21_X1 U11049 ( .B1(n10546), .B2(n10675), .A(n10516), .ZN(n10218) );
  AND2_X1 U11050 ( .A1(n10542), .A2(n10543), .ZN(n10523) );
  INV_X1 U11051 ( .A(n10523), .ZN(n10217) );
  OAI211_X1 U11052 ( .C1(n6883), .C2(n10518), .A(n10218), .B(n10217), .ZN(
        n10527) );
  AOI22_X1 U11053 ( .A1(n10677), .A2(n10527), .B1(P1_REG1_REG_0__SCAN_IN), 
        .B2(n10676), .ZN(n10219) );
  XNOR2_X1 U11054 ( .A(n10220), .B(n10219), .ZN(P1_U3522) );
  OAI21_X1 U11055 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(n10223), .ZN(n10221) );
  INV_X1 U11056 ( .A(n10221), .ZN(ADD_1068_U46) );
  OAI21_X1 U11057 ( .B1(n10224), .B2(n10223), .A(n10222), .ZN(n10225) );
  XNOR2_X1 U11058 ( .A(n10225), .B(P2_ADDR_REG_1__SCAN_IN), .ZN(ADD_1068_U5)
         );
  AOI21_X1 U11059 ( .B1(n10228), .B2(n10227), .A(n10226), .ZN(ADD_1068_U54) );
  AOI21_X1 U11060 ( .B1(n10231), .B2(n10230), .A(n10229), .ZN(ADD_1068_U53) );
  OAI21_X1 U11061 ( .B1(n10234), .B2(n10233), .A(n10232), .ZN(ADD_1068_U52) );
  OAI21_X1 U11062 ( .B1(n10237), .B2(n10236), .A(n10235), .ZN(ADD_1068_U51) );
  OAI21_X1 U11063 ( .B1(n10240), .B2(n10239), .A(n10238), .ZN(ADD_1068_U50) );
  OAI21_X1 U11064 ( .B1(n10243), .B2(n10242), .A(n10241), .ZN(ADD_1068_U49) );
  OAI21_X1 U11065 ( .B1(n10246), .B2(n10245), .A(n10244), .ZN(ADD_1068_U48) );
  OAI21_X1 U11066 ( .B1(n10249), .B2(n10248), .A(n10247), .ZN(ADD_1068_U47) );
  OAI21_X1 U11067 ( .B1(n10252), .B2(n10251), .A(n10250), .ZN(ADD_1068_U63) );
  OAI21_X1 U11068 ( .B1(n10255), .B2(n10254), .A(n10253), .ZN(ADD_1068_U62) );
  OAI21_X1 U11069 ( .B1(n10258), .B2(n10257), .A(n10256), .ZN(ADD_1068_U61) );
  OAI21_X1 U11070 ( .B1(n10261), .B2(n10260), .A(n10259), .ZN(ADD_1068_U60) );
  OAI21_X1 U11071 ( .B1(n10264), .B2(n10263), .A(n10262), .ZN(ADD_1068_U59) );
  OAI21_X1 U11072 ( .B1(n10267), .B2(n10266), .A(n10265), .ZN(ADD_1068_U58) );
  OAI21_X1 U11073 ( .B1(n10270), .B2(n10269), .A(n10268), .ZN(ADD_1068_U57) );
  OAI21_X1 U11074 ( .B1(n10273), .B2(n10272), .A(n10271), .ZN(ADD_1068_U56) );
  OAI21_X1 U11075 ( .B1(n10276), .B2(n10275), .A(n10274), .ZN(ADD_1068_U55) );
  AOI21_X1 U11076 ( .B1(n10279), .B2(n10278), .A(n10277), .ZN(P1_U3440) );
  INV_X1 U11077 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n10294) );
  OAI21_X1 U11078 ( .B1(n10281), .B2(n10280), .A(n10329), .ZN(n10283) );
  NOR2_X1 U11079 ( .A1(n10283), .A2(n10282), .ZN(n10290) );
  INV_X1 U11080 ( .A(n10284), .ZN(n10288) );
  INV_X1 U11081 ( .A(n10285), .ZN(n10287) );
  INV_X1 U11082 ( .A(n10334), .ZN(n10379) );
  AOI211_X1 U11083 ( .C1(n10288), .C2(n10287), .A(n10286), .B(n10379), .ZN(
        n10289) );
  AOI211_X1 U11084 ( .C1(n10390), .C2(n10291), .A(n10290), .B(n10289), .ZN(
        n10293) );
  OAI211_X1 U11085 ( .C1(n10394), .C2(n10294), .A(n10293), .B(n10292), .ZN(
        P1_U3250) );
  INV_X1 U11086 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n10311) );
  INV_X1 U11087 ( .A(n10295), .ZN(n10307) );
  AOI21_X1 U11088 ( .B1(n10298), .B2(n10297), .A(n10296), .ZN(n10299) );
  NAND2_X1 U11089 ( .A1(n10329), .A2(n10299), .ZN(n10306) );
  NAND2_X1 U11090 ( .A1(n10301), .A2(n10300), .ZN(n10304) );
  INV_X1 U11091 ( .A(n10302), .ZN(n10303) );
  NAND3_X1 U11092 ( .A1(n10334), .A2(n10304), .A3(n10303), .ZN(n10305) );
  OAI211_X1 U11093 ( .C1(n10338), .C2(n10307), .A(n10306), .B(n10305), .ZN(
        n10308) );
  INV_X1 U11094 ( .A(n10308), .ZN(n10310) );
  OAI211_X1 U11095 ( .C1(n10394), .C2(n10311), .A(n10310), .B(n10309), .ZN(
        P1_U3251) );
  INV_X1 U11096 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n10323) );
  AOI211_X1 U11097 ( .C1(n10314), .C2(n10313), .A(n10312), .B(n10383), .ZN(
        n10319) );
  AOI211_X1 U11098 ( .C1(n10317), .C2(n10316), .A(n10315), .B(n10379), .ZN(
        n10318) );
  AOI211_X1 U11099 ( .C1(n10390), .C2(n10320), .A(n10319), .B(n10318), .ZN(
        n10322) );
  OAI211_X1 U11100 ( .C1(n10394), .C2(n10323), .A(n10322), .B(n10321), .ZN(
        P1_U3254) );
  INV_X1 U11101 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n10342) );
  INV_X1 U11102 ( .A(n10324), .ZN(n10337) );
  AOI21_X1 U11103 ( .B1(n10327), .B2(n10326), .A(n10325), .ZN(n10328) );
  NAND2_X1 U11104 ( .A1(n10329), .A2(n10328), .ZN(n10336) );
  AOI21_X1 U11105 ( .B1(n10332), .B2(n10331), .A(n10330), .ZN(n10333) );
  NAND2_X1 U11106 ( .A1(n10334), .A2(n10333), .ZN(n10335) );
  OAI211_X1 U11107 ( .C1(n10338), .C2(n10337), .A(n10336), .B(n10335), .ZN(
        n10339) );
  INV_X1 U11108 ( .A(n10339), .ZN(n10341) );
  OAI211_X1 U11109 ( .C1(n10394), .C2(n10342), .A(n10341), .B(n10340), .ZN(
        P1_U3257) );
  INV_X1 U11110 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n10353) );
  AOI211_X1 U11111 ( .C1(n10345), .C2(n10344), .A(n10343), .B(n10379), .ZN(
        n10349) );
  AOI211_X1 U11112 ( .C1(n10347), .C2(n8092), .A(n10346), .B(n10383), .ZN(
        n10348) );
  AOI211_X1 U11113 ( .C1(n10390), .C2(n10350), .A(n10349), .B(n10348), .ZN(
        n10352) );
  OAI211_X1 U11114 ( .C1(n10394), .C2(n10353), .A(n10352), .B(n10351), .ZN(
        P1_U3258) );
  INV_X1 U11115 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10366) );
  AOI211_X1 U11116 ( .C1(n10356), .C2(n10355), .A(n10379), .B(n10354), .ZN(
        n10362) );
  INV_X1 U11117 ( .A(n10357), .ZN(n10358) );
  AOI211_X1 U11118 ( .C1(n10360), .C2(n10359), .A(n10383), .B(n10358), .ZN(
        n10361) );
  AOI211_X1 U11119 ( .C1(n10390), .C2(n10363), .A(n10362), .B(n10361), .ZN(
        n10365) );
  OAI211_X1 U11120 ( .C1(n10394), .C2(n10366), .A(n10365), .B(n10364), .ZN(
        P1_U3261) );
  INV_X1 U11121 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n10378) );
  AOI211_X1 U11122 ( .C1(n10369), .C2(n10368), .A(n10367), .B(n10379), .ZN(
        n10374) );
  AOI211_X1 U11123 ( .C1(n10372), .C2(n10371), .A(n10370), .B(n10383), .ZN(
        n10373) );
  AOI211_X1 U11124 ( .C1(n10390), .C2(n10375), .A(n10374), .B(n10373), .ZN(
        n10377) );
  NAND2_X1 U11125 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n10376)
         );
  OAI211_X1 U11126 ( .C1(n10394), .C2(n10378), .A(n10377), .B(n10376), .ZN(
        P1_U3256) );
  INV_X1 U11127 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n10393) );
  AOI211_X1 U11128 ( .C1(n10382), .C2(n10381), .A(n10380), .B(n10379), .ZN(
        n10388) );
  AOI211_X1 U11129 ( .C1(n10386), .C2(n10385), .A(n10384), .B(n10383), .ZN(
        n10387) );
  AOI211_X1 U11130 ( .C1(n10390), .C2(n10389), .A(n10388), .B(n10387), .ZN(
        n10392) );
  OAI211_X1 U11131 ( .C1(n10394), .C2(n10393), .A(n10392), .B(n10391), .ZN(
        P1_U3253) );
  INV_X1 U11132 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n10414) );
  AOI21_X1 U11133 ( .B1(n10397), .B2(n10396), .A(n10395), .ZN(n10405) );
  AOI21_X1 U11134 ( .B1(n10400), .B2(n10399), .A(n10398), .ZN(n10401) );
  OR2_X1 U11135 ( .A1(n10501), .A2(n10401), .ZN(n10404) );
  INV_X1 U11136 ( .A(n10402), .ZN(n10403) );
  OAI211_X1 U11137 ( .C1(n10405), .C2(n10506), .A(n10404), .B(n10403), .ZN(
        n10408) );
  NOR2_X1 U11138 ( .A1(n10507), .A2(n10406), .ZN(n10407) );
  NOR2_X1 U11139 ( .A1(n10408), .A2(n10407), .ZN(n10413) );
  OAI211_X1 U11140 ( .C1(n10411), .C2(n10410), .A(n10409), .B(n10495), .ZN(
        n10412) );
  OAI211_X1 U11141 ( .C1(n10414), .C2(n10489), .A(n10413), .B(n10412), .ZN(
        P2_U3186) );
  INV_X1 U11142 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n10432) );
  AOI21_X1 U11143 ( .B1(n10605), .B2(n10416), .A(n10415), .ZN(n10425) );
  AOI21_X1 U11144 ( .B1(n10474), .B2(n10418), .A(n10417), .ZN(n10424) );
  AOI21_X1 U11145 ( .B1(n10421), .B2(n10420), .A(n10419), .ZN(n10422) );
  OR2_X1 U11146 ( .A1(n10422), .A2(n10506), .ZN(n10423) );
  OAI211_X1 U11147 ( .C1(n10425), .C2(n10501), .A(n10424), .B(n10423), .ZN(
        n10426) );
  INV_X1 U11148 ( .A(n10426), .ZN(n10431) );
  XOR2_X1 U11149 ( .A(n10428), .B(n10427), .Z(n10429) );
  NAND2_X1 U11150 ( .A1(n10429), .A2(n10495), .ZN(n10430) );
  OAI211_X1 U11151 ( .C1(n10432), .C2(n10489), .A(n10431), .B(n10430), .ZN(
        P2_U3187) );
  AOI21_X1 U11152 ( .B1(n5026), .B2(n10434), .A(n10433), .ZN(n10436) );
  OAI22_X1 U11153 ( .A1(n10436), .A2(n10506), .B1(n10435), .B2(n10507), .ZN(
        n10437) );
  AOI21_X1 U11154 ( .B1(n10498), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n10437), .ZN(
        n10449) );
  OAI21_X1 U11155 ( .B1(n10440), .B2(n10439), .A(n10438), .ZN(n10441) );
  NAND2_X1 U11156 ( .A1(n10441), .A2(n10495), .ZN(n10447) );
  AOI21_X1 U11157 ( .B1(n10444), .B2(n10443), .A(n10442), .ZN(n10445) );
  OR2_X1 U11158 ( .A1(n10445), .A2(n10501), .ZN(n10446) );
  NAND4_X1 U11159 ( .A1(n10449), .A2(n10448), .A3(n10447), .A4(n10446), .ZN(
        P2_U3188) );
  INV_X1 U11160 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n10468) );
  AOI21_X1 U11161 ( .B1(n10626), .B2(n10451), .A(n10450), .ZN(n10460) );
  AOI21_X1 U11162 ( .B1(n10474), .B2(n10453), .A(n10452), .ZN(n10459) );
  AOI21_X1 U11163 ( .B1(n10456), .B2(n10455), .A(n10454), .ZN(n10457) );
  OR2_X1 U11164 ( .A1(n10457), .A2(n10506), .ZN(n10458) );
  OAI211_X1 U11165 ( .C1(n10460), .C2(n10501), .A(n10459), .B(n10458), .ZN(
        n10461) );
  INV_X1 U11166 ( .A(n10461), .ZN(n10467) );
  OAI21_X1 U11167 ( .B1(n10464), .B2(n10463), .A(n10462), .ZN(n10465) );
  NAND2_X1 U11168 ( .A1(n10465), .A2(n10495), .ZN(n10466) );
  OAI211_X1 U11169 ( .C1(n10468), .C2(n10489), .A(n10467), .B(n10466), .ZN(
        P2_U3189) );
  INV_X1 U11170 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n10490) );
  AOI21_X1 U11171 ( .B1(n10471), .B2(n10470), .A(n10469), .ZN(n10481) );
  AOI21_X1 U11172 ( .B1(n10474), .B2(n10473), .A(n10472), .ZN(n10480) );
  AOI21_X1 U11173 ( .B1(n10477), .B2(n10476), .A(n10475), .ZN(n10478) );
  OR2_X1 U11174 ( .A1(n10478), .A2(n10506), .ZN(n10479) );
  OAI211_X1 U11175 ( .C1(n10481), .C2(n10501), .A(n10480), .B(n10479), .ZN(
        n10482) );
  INV_X1 U11176 ( .A(n10482), .ZN(n10488) );
  NOR2_X1 U11177 ( .A1(n10484), .A2(n10483), .ZN(n10485) );
  OAI21_X1 U11178 ( .B1(n10486), .B2(n10485), .A(n10495), .ZN(n10487) );
  OAI211_X1 U11179 ( .C1(n10490), .C2(n10489), .A(n10488), .B(n10487), .ZN(
        P2_U3190) );
  INV_X1 U11180 ( .A(n10491), .ZN(n10493) );
  NAND2_X1 U11181 ( .A1(n10493), .A2(n10492), .ZN(n10509) );
  AND3_X1 U11182 ( .A1(n10509), .A2(n10495), .A3(n10494), .ZN(n10496) );
  AOI211_X1 U11183 ( .C1(n10498), .C2(P2_ADDR_REG_18__SCAN_IN), .A(n10497), 
        .B(n10496), .ZN(n10514) );
  AOI21_X1 U11184 ( .B1(n10500), .B2(n4993), .A(n10499), .ZN(n10502) );
  OAI21_X1 U11185 ( .B1(n10509), .B2(n10508), .A(n10507), .ZN(n10511) );
  NAND2_X1 U11186 ( .A1(n10511), .A2(n10510), .ZN(n10512) );
  XNOR2_X1 U11187 ( .A(P2_RD_REG_SCAN_IN), .B(P1_RD_REG_SCAN_IN), .ZN(U126) );
  INV_X1 U11188 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n10526) );
  AND2_X1 U11189 ( .A1(n10516), .A2(n10515), .ZN(n10521) );
  NOR2_X1 U11190 ( .A1(n10518), .A2(n10517), .ZN(n10520) );
  MUX2_X1 U11191 ( .A(n10521), .B(n10520), .S(n10519), .Z(n10522) );
  AOI211_X1 U11192 ( .C1(n10554), .C2(P1_REG3_REG_0__SCAN_IN), .A(n10523), .B(
        n10522), .ZN(n10525) );
  AOI22_X1 U11193 ( .A1(n10555), .A2(n10526), .B1(n10525), .B2(n10524), .ZN(
        P1_U3293) );
  MUX2_X1 U11194 ( .A(n10527), .B(P1_REG0_REG_0__SCAN_IN), .S(n10678), .Z(
        P1_U3453) );
  INV_X1 U11195 ( .A(n10613), .ZN(n10634) );
  INV_X1 U11196 ( .A(n10528), .ZN(n10529) );
  OAI21_X1 U11197 ( .B1(n6373), .B2(n10669), .A(n10529), .ZN(n10530) );
  AOI211_X1 U11198 ( .C1(n10634), .C2(n10532), .A(n10531), .B(n10530), .ZN(
        n10535) );
  AOI22_X1 U11199 ( .A1(n10677), .A2(n10535), .B1(n10533), .B2(n10676), .ZN(
        P1_U3523) );
  INV_X1 U11200 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n10534) );
  AOI22_X1 U11201 ( .A1(n10681), .A2(n10535), .B1(n10534), .B2(n10678), .ZN(
        P1_U3456) );
  OAI211_X1 U11202 ( .C1(n5025), .C2(n10538), .A(n10537), .B(n10536), .ZN(
        n10556) );
  OAI21_X1 U11203 ( .B1(n10538), .B2(n10669), .A(n10556), .ZN(n10548) );
  XOR2_X1 U11204 ( .A(n10540), .B(n10539), .Z(n10545) );
  AOI222_X1 U11205 ( .A1(n10546), .A2(n10545), .B1(n10544), .B2(n10543), .C1(
        n10542), .C2(n10541), .ZN(n10563) );
  INV_X1 U11206 ( .A(n10563), .ZN(n10547) );
  AOI211_X1 U11207 ( .C1(n10675), .C2(n10560), .A(n10548), .B(n10547), .ZN(
        n10551) );
  AOI22_X1 U11208 ( .A1(n10677), .A2(n10551), .B1(n10549), .B2(n10676), .ZN(
        P1_U3524) );
  INV_X1 U11209 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n10550) );
  AOI22_X1 U11210 ( .A1(n10681), .A2(n10551), .B1(n10550), .B2(n10678), .ZN(
        P1_U3459) );
  AOI222_X1 U11211 ( .A1(P1_REG2_REG_2__SCAN_IN), .A2(n10555), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n10554), .C1(n10553), .C2(n10552), .ZN(
        n10562) );
  INV_X1 U11212 ( .A(n10556), .ZN(n10557) );
  AOI22_X1 U11213 ( .A1(n10560), .A2(n10559), .B1(n4924), .B2(n10557), .ZN(
        n10561) );
  OAI211_X1 U11214 ( .C1(n10555), .C2(n10563), .A(n10562), .B(n10561), .ZN(
        P1_U3291) );
  AOI211_X1 U11215 ( .C1(n10749), .C2(n10566), .A(n10565), .B(n10564), .ZN(
        n10568) );
  AOI22_X1 U11216 ( .A1(n10761), .A2(n10568), .B1(n5766), .B2(n10760), .ZN(
        P2_U3461) );
  INV_X1 U11217 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10567) );
  AOI22_X1 U11218 ( .A1(n10764), .A2(n10568), .B1(n10567), .B2(n6872), .ZN(
        P2_U3396) );
  INV_X1 U11219 ( .A(n10569), .ZN(n10574) );
  OAI21_X1 U11220 ( .B1(n10571), .B2(n10669), .A(n10570), .ZN(n10573) );
  AOI211_X1 U11221 ( .C1(n10634), .C2(n10574), .A(n10573), .B(n10572), .ZN(
        n10576) );
  AOI22_X1 U11222 ( .A1(n10677), .A2(n10576), .B1(n7177), .B2(n10676), .ZN(
        P1_U3525) );
  INV_X1 U11223 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n10575) );
  AOI22_X1 U11224 ( .A1(n10681), .A2(n10576), .B1(n10575), .B2(n10678), .ZN(
        P1_U3462) );
  NOR2_X1 U11225 ( .A1(n10577), .A2(n10740), .ZN(n10579) );
  AOI211_X1 U11226 ( .C1(n10749), .C2(n10580), .A(n10579), .B(n10578), .ZN(
        n10583) );
  AOI22_X1 U11227 ( .A1(n10761), .A2(n10583), .B1(n10581), .B2(n10760), .ZN(
        P2_U3462) );
  INV_X1 U11228 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10582) );
  AOI22_X1 U11229 ( .A1(n10764), .A2(n10583), .B1(n10582), .B2(n6872), .ZN(
        P2_U3399) );
  OR2_X1 U11230 ( .A1(n10584), .A2(n10710), .ZN(n10587) );
  NAND2_X1 U11231 ( .A1(n10585), .A2(n10751), .ZN(n10586) );
  AOI22_X1 U11232 ( .A1(n10761), .A2(n10591), .B1(n10589), .B2(n10760), .ZN(
        P2_U3463) );
  INV_X1 U11233 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10590) );
  AOI22_X1 U11234 ( .A1(n10764), .A2(n10591), .B1(n10590), .B2(n6872), .ZN(
        P2_U3402) );
  OAI21_X1 U11235 ( .B1(n10593), .B2(n10669), .A(n10592), .ZN(n10595) );
  AOI211_X1 U11236 ( .C1(n10675), .C2(n10596), .A(n10595), .B(n10594), .ZN(
        n10598) );
  AOI22_X1 U11237 ( .A1(n10677), .A2(n10598), .B1(n7179), .B2(n10676), .ZN(
        P1_U3526) );
  INV_X1 U11238 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10597) );
  AOI22_X1 U11239 ( .A1(n10681), .A2(n10598), .B1(n10597), .B2(n10678), .ZN(
        P1_U3465) );
  NOR2_X1 U11240 ( .A1(n10599), .A2(n10710), .ZN(n10604) );
  OAI22_X1 U11241 ( .A1(n10601), .A2(n10754), .B1(n10600), .B2(n10740), .ZN(
        n10603) );
  AOI211_X1 U11242 ( .C1(n10604), .C2(n7662), .A(n10603), .B(n10602), .ZN(
        n10607) );
  AOI22_X1 U11243 ( .A1(n10761), .A2(n10607), .B1(n10605), .B2(n10760), .ZN(
        P2_U3464) );
  INV_X1 U11244 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10606) );
  AOI22_X1 U11245 ( .A1(n10764), .A2(n10607), .B1(n10606), .B2(n6872), .ZN(
        P2_U3405) );
  AOI21_X1 U11246 ( .B1(n10610), .B2(n10609), .A(n10608), .ZN(n10611) );
  OAI211_X1 U11247 ( .C1(n10614), .C2(n10613), .A(n10612), .B(n10611), .ZN(
        n10615) );
  INV_X1 U11248 ( .A(n10615), .ZN(n10618) );
  AOI22_X1 U11249 ( .A1(n10677), .A2(n10618), .B1(n10616), .B2(n10676), .ZN(
        P1_U3528) );
  INV_X1 U11250 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10617) );
  AOI22_X1 U11251 ( .A1(n10681), .A2(n10618), .B1(n10617), .B2(n10678), .ZN(
        P1_U3471) );
  AOI22_X1 U11252 ( .A1(n10620), .A2(n10658), .B1(n10619), .B2(n10751), .ZN(
        n10621) );
  OAI21_X1 U11253 ( .B1(n10622), .B2(n10684), .A(n10621), .ZN(n10625) );
  NOR2_X1 U11254 ( .A1(n10622), .A2(n10683), .ZN(n10624) );
  NOR3_X1 U11255 ( .A1(n10625), .A2(n10624), .A3(n10623), .ZN(n10628) );
  AOI22_X1 U11256 ( .A1(n10761), .A2(n10628), .B1(n10626), .B2(n10760), .ZN(
        P2_U3466) );
  INV_X1 U11257 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10627) );
  AOI22_X1 U11258 ( .A1(n10764), .A2(n10628), .B1(n10627), .B2(n6872), .ZN(
        P2_U3411) );
  OAI21_X1 U11259 ( .B1(n10630), .B2(n10669), .A(n10629), .ZN(n10632) );
  AOI211_X1 U11260 ( .C1(n10634), .C2(n10633), .A(n10632), .B(n10631), .ZN(
        n10636) );
  AOI22_X1 U11261 ( .A1(n10677), .A2(n10636), .B1(n7187), .B2(n10676), .ZN(
        P1_U3530) );
  INV_X1 U11262 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n10635) );
  AOI22_X1 U11263 ( .A1(n10681), .A2(n10636), .B1(n10635), .B2(n10678), .ZN(
        P1_U3477) );
  OAI21_X1 U11264 ( .B1(n5525), .B2(n10638), .A(n10637), .ZN(n10644) );
  AOI222_X1 U11265 ( .A1(n10644), .A2(n10643), .B1(n10642), .B2(n10641), .C1(
        n10640), .C2(n10639), .ZN(n10645) );
  OAI21_X1 U11266 ( .B1(n10647), .B2(n10646), .A(n10645), .ZN(P2_U3225) );
  OAI21_X1 U11267 ( .B1(n10649), .B2(n10669), .A(n10648), .ZN(n10650) );
  AOI21_X1 U11268 ( .B1(n10651), .B2(n10675), .A(n10650), .ZN(n10652) );
  AND2_X1 U11269 ( .A1(n10653), .A2(n10652), .ZN(n10656) );
  AOI22_X1 U11270 ( .A1(n10677), .A2(n10656), .B1(n10654), .B2(n10676), .ZN(
        P1_U3531) );
  INV_X1 U11271 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n10655) );
  AOI22_X1 U11272 ( .A1(n10681), .A2(n10656), .B1(n10655), .B2(n10678), .ZN(
        P1_U3480) );
  INV_X1 U11273 ( .A(n10683), .ZN(n10664) );
  AOI22_X1 U11274 ( .A1(n5895), .A2(n10751), .B1(n10658), .B2(n10657), .ZN(
        n10659) );
  OAI21_X1 U11275 ( .B1(n10660), .B2(n10684), .A(n10659), .ZN(n10662) );
  AOI211_X1 U11276 ( .C1(n10664), .C2(n10663), .A(n10662), .B(n10661), .ZN(
        n10667) );
  AOI22_X1 U11277 ( .A1(n10761), .A2(n10667), .B1(n10665), .B2(n10760), .ZN(
        P2_U3468) );
  INV_X1 U11278 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10666) );
  AOI22_X1 U11279 ( .A1(n10764), .A2(n10667), .B1(n10666), .B2(n6872), .ZN(
        P2_U3417) );
  OAI21_X1 U11280 ( .B1(n10670), .B2(n10669), .A(n10668), .ZN(n10673) );
  INV_X1 U11281 ( .A(n10671), .ZN(n10672) );
  AOI211_X1 U11282 ( .C1(n10675), .C2(n10674), .A(n10673), .B(n10672), .ZN(
        n10680) );
  AOI22_X1 U11283 ( .A1(n10677), .A2(n10680), .B1(n7352), .B2(n10676), .ZN(
        P1_U3532) );
  INV_X1 U11284 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n10679) );
  AOI22_X1 U11285 ( .A1(n10681), .A2(n10680), .B1(n10679), .B2(n10678), .ZN(
        P1_U3483) );
  AOI21_X1 U11286 ( .B1(n10684), .B2(n10683), .A(n10682), .ZN(n10689) );
  INV_X1 U11287 ( .A(n10685), .ZN(n10687) );
  OAI22_X1 U11288 ( .A1(n10687), .A2(n10740), .B1(n10686), .B2(n10754), .ZN(
        n10688) );
  NOR3_X1 U11289 ( .A1(n10690), .A2(n10689), .A3(n10688), .ZN(n10693) );
  AOI22_X1 U11290 ( .A1(n10761), .A2(n10693), .B1(n10691), .B2(n10760), .ZN(
        P2_U3469) );
  INV_X1 U11291 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10692) );
  AOI22_X1 U11292 ( .A1(n10764), .A2(n10693), .B1(n10692), .B2(n6872), .ZN(
        P2_U3420) );
  INV_X1 U11293 ( .A(n10694), .ZN(n10700) );
  INV_X1 U11294 ( .A(n10695), .ZN(n10697) );
  OAI22_X1 U11295 ( .A1(n10697), .A2(n10740), .B1(n10696), .B2(n10754), .ZN(
        n10699) );
  AOI211_X1 U11296 ( .C1(n10700), .C2(n10749), .A(n10699), .B(n10698), .ZN(
        n10703) );
  AOI22_X1 U11297 ( .A1(n10761), .A2(n10703), .B1(n10701), .B2(n10760), .ZN(
        P2_U3470) );
  INV_X1 U11298 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10702) );
  AOI22_X1 U11299 ( .A1(n10764), .A2(n10703), .B1(n10702), .B2(n6872), .ZN(
        P2_U3423) );
  NOR2_X1 U11300 ( .A1(n10704), .A2(n10710), .ZN(n10707) );
  INV_X1 U11301 ( .A(n10705), .ZN(n10706) );
  AOI211_X1 U11302 ( .C1(n10751), .C2(n10708), .A(n10707), .B(n10706), .ZN(
        n10709) );
  AOI22_X1 U11303 ( .A1(n10761), .A2(n10709), .B1(n5624), .B2(n10760), .ZN(
        P2_U3471) );
  AOI22_X1 U11304 ( .A1(n10764), .A2(n10709), .B1(n5931), .B2(n6872), .ZN(
        P2_U3426) );
  NOR2_X1 U11305 ( .A1(n10711), .A2(n10710), .ZN(n10713) );
  AOI211_X1 U11306 ( .C1(n10751), .C2(n10714), .A(n10713), .B(n10712), .ZN(
        n10717) );
  AOI22_X1 U11307 ( .A1(n10761), .A2(n10717), .B1(n10715), .B2(n10760), .ZN(
        P2_U3472) );
  INV_X1 U11308 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n10716) );
  AOI22_X1 U11309 ( .A1(n10764), .A2(n10717), .B1(n10716), .B2(n6872), .ZN(
        P2_U3429) );
  NOR2_X1 U11310 ( .A1(n10718), .A2(n10740), .ZN(n10720) );
  AOI211_X1 U11311 ( .C1(n10749), .C2(n10721), .A(n10720), .B(n10719), .ZN(
        n10723) );
  AOI22_X1 U11312 ( .A1(n10761), .A2(n10723), .B1(n5969), .B2(n10760), .ZN(
        P2_U3473) );
  INV_X1 U11313 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n10722) );
  AOI22_X1 U11314 ( .A1(n10764), .A2(n10723), .B1(n10722), .B2(n6872), .ZN(
        P2_U3432) );
  AND2_X1 U11315 ( .A1(n10724), .A2(n10749), .ZN(n10727) );
  AND2_X1 U11316 ( .A1(n10725), .A2(n10751), .ZN(n10726) );
  NOR3_X1 U11317 ( .A1(n10728), .A2(n10727), .A3(n10726), .ZN(n10731) );
  AOI22_X1 U11318 ( .A1(n10761), .A2(n10731), .B1(n10729), .B2(n10760), .ZN(
        P2_U3474) );
  INV_X1 U11319 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n10730) );
  AOI22_X1 U11320 ( .A1(n10764), .A2(n10731), .B1(n10730), .B2(n6872), .ZN(
        P2_U3435) );
  NOR2_X1 U11321 ( .A1(n10732), .A2(n10740), .ZN(n10734) );
  AOI211_X1 U11322 ( .C1(n10735), .C2(n10749), .A(n10734), .B(n10733), .ZN(
        n10738) );
  AOI22_X1 U11323 ( .A1(n10761), .A2(n10738), .B1(n10736), .B2(n10760), .ZN(
        P2_U3475) );
  INV_X1 U11324 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n10737) );
  AOI22_X1 U11325 ( .A1(n10764), .A2(n10738), .B1(n10737), .B2(n6872), .ZN(
        P2_U3438) );
  OAI22_X1 U11326 ( .A1(n10741), .A2(n10740), .B1(n10739), .B2(n10754), .ZN(
        n10744) );
  INV_X1 U11327 ( .A(n10742), .ZN(n10743) );
  AOI211_X1 U11328 ( .C1(n10745), .C2(n10749), .A(n10744), .B(n10743), .ZN(
        n10748) );
  AOI22_X1 U11329 ( .A1(n10761), .A2(n10748), .B1(n10746), .B2(n10760), .ZN(
        P2_U3476) );
  INV_X1 U11330 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n10747) );
  AOI22_X1 U11331 ( .A1(n10764), .A2(n10748), .B1(n10747), .B2(n6872), .ZN(
        P2_U3441) );
  AND2_X1 U11332 ( .A1(n10750), .A2(n10749), .ZN(n10757) );
  NAND2_X1 U11333 ( .A1(n10752), .A2(n10751), .ZN(n10753) );
  OAI21_X1 U11334 ( .B1(n10755), .B2(n10754), .A(n10753), .ZN(n10756) );
  AOI21_X1 U11335 ( .B1(n10757), .B2(n9180), .A(n10756), .ZN(n10758) );
  AND2_X1 U11336 ( .A1(n10759), .A2(n10758), .ZN(n10763) );
  AOI22_X1 U11337 ( .A1(n10761), .A2(n10763), .B1(n5643), .B2(n10760), .ZN(
        P2_U3477) );
  INV_X1 U11338 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n10762) );
  AOI22_X1 U11339 ( .A1(n10764), .A2(n10763), .B1(n10762), .B2(n6872), .ZN(
        P2_U3444) );
  XNOR2_X1 U11340 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
endmodule

