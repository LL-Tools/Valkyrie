

module b14_C_SARLock_k_64_9 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, U3352, U3351, U3350, U3349, U3348, U3347, 
        U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, U3338, U3337, 
        U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, U3328, U3327, 
        U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, U3320, U3319, 
        U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, U3310, U3309, 
        U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, U3300, U3299, 
        U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, U3467, U3469, 
        U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, U3487, U3489, 
        U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, U3506, U3507, 
        U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, U3516, U3517, 
        U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, U3526, U3527, 
        U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, U3536, U3537, 
        U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, U3546, U3547, 
        U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, U3284, U3283, 
        U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, U3274, U3273, 
        U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, U3264, U3263, 
        U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, U3255, U3254, 
        U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, U3245, U3244, 
        U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, U3554, U3555, 
        U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, U3564, U3565, 
        U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, U3574, U3575, 
        U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, U3237, U3236, 
        U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, U3227, U3226, 
        U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, U3217, U3216, 
        U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, U4043 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599;

  INV_X1 U2255 ( .A(n2798), .ZN(n2626) );
  INV_X1 U2256 ( .A(n2763), .ZN(n2800) );
  AOI21_X1 U2258 ( .B1(n3038), .B2(n3039), .A(n2618), .ZN(n3047) );
  CLKBUF_X1 U2259 ( .A(n2254), .Z(n3840) );
  NAND2_X1 U2260 ( .A1(n2508), .A2(n3808), .ZN(n2603) );
  NAND3_X2 U2261 ( .A1(n4202), .A2(n4204), .A3(n4203), .ZN(n2604) );
  CLKBUF_X1 U2262 ( .A(n2217), .Z(n2349) );
  CLKBUF_X1 U2263 ( .A(n2268), .Z(n2269) );
  OR2_X1 U2264 ( .A1(n2816), .A2(n2815), .ZN(n2838) );
  NAND2_X1 U2265 ( .A1(n2524), .A2(n3726), .ZN(n3231) );
  OR2_X1 U2266 ( .A1(n3209), .A2(n3208), .ZN(n2524) );
  AND2_X1 U2267 ( .A1(n2624), .A2(n2625), .ZN(n3046) );
  NAND2_X1 U2268 ( .A1(n3706), .A2(n3703), .ZN(n2520) );
  NOR2_X1 U2269 ( .A1(n2608), .A2(n2015), .ZN(n2613) );
  AND2_X2 U2270 ( .A1(n2594), .A2(n4590), .ZN(n3035) );
  OAI21_X1 U2271 ( .B1(n3021), .B2(n2999), .A(n3000), .ZN(n3191) );
  OR2_X1 U2272 ( .A1(n4383), .A2(n3134), .ZN(n2280) );
  OAI21_X1 U2273 ( .B1(n2799), .B2(n3060), .A(n2111), .ZN(n2110) );
  AND4_X2 U2274 ( .A1(n2266), .A2(n2265), .A3(n2264), .A4(n2263), .ZN(n3138)
         );
  NAND4_X2 U2275 ( .A1(n2277), .A2(n2276), .A3(n2275), .A4(n2274), .ZN(n4383)
         );
  INV_X1 U2276 ( .A(n2254), .ZN(n3015) );
  XNOR2_X1 U2277 ( .A(n2996), .B(n2984), .ZN(n2995) );
  INV_X1 U2278 ( .A(n2802), .ZN(n2774) );
  NAND2_X1 U2279 ( .A1(n3006), .A2(n2982), .ZN(n2996) );
  CLKBUF_X3 U2280 ( .A(n2262), .Z(n3668) );
  NOR2_X1 U2281 ( .A1(n2799), .A2(n2053), .ZN(n2131) );
  INV_X1 U2282 ( .A(n2602), .ZN(n3060) );
  AND2_X1 U2283 ( .A1(n2239), .A2(n2240), .ZN(n2262) );
  NAND2_X2 U2284 ( .A1(n2604), .A2(n2603), .ZN(n2798) );
  AND2_X1 U2285 ( .A1(n2231), .A2(n3505), .ZN(n2924) );
  XNOR2_X1 U2286 ( .A(n2233), .B(IR_REG_30__SCAN_IN), .ZN(n4200) );
  MUX2_X1 U2287 ( .A(IR_REG_31__SCAN_IN), .B(n2230), .S(IR_REG_29__SCAN_IN), 
        .Z(n2231) );
  XNOR2_X1 U2288 ( .A(n2565), .B(IR_REG_26__SCAN_IN), .ZN(n4202) );
  OAI21_X1 U2289 ( .B1(n2228), .B2(IR_REG_26__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2598) );
  OR2_X1 U2290 ( .A1(n2228), .A2(n2183), .ZN(n2517) );
  XNOR2_X1 U2291 ( .A(n2506), .B(IR_REG_21__SCAN_IN), .ZN(n3808) );
  NAND2_X1 U2292 ( .A1(n2228), .A2(IR_REG_31__SCAN_IN), .ZN(n2565) );
  AND2_X1 U2293 ( .A1(n2504), .A2(n2186), .ZN(n2560) );
  AND2_X1 U2294 ( .A1(n2013), .A2(n2034), .ZN(n2104) );
  NOR2_X1 U2295 ( .A1(IR_REG_11__SCAN_IN), .A2(IR_REG_14__SCAN_IN), .ZN(n2207)
         );
  NOR2_X1 U2296 ( .A1(IR_REG_15__SCAN_IN), .A2(IR_REG_13__SCAN_IN), .ZN(n2206)
         );
  NOR2_X1 U2297 ( .A1(IR_REG_12__SCAN_IN), .A2(IR_REG_16__SCAN_IN), .ZN(n2205)
         );
  INV_X1 U2298 ( .A(IR_REG_20__SCAN_IN), .ZN(n2502) );
  INV_X1 U2299 ( .A(IR_REG_19__SCAN_IN), .ZN(n2448) );
  INV_X1 U2300 ( .A(IR_REG_5__SCAN_IN), .ZN(n2301) );
  INV_X4 U2301 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  INV_X1 U2302 ( .A(IR_REG_4__SCAN_IN), .ZN(n2297) );
  INV_X1 U2303 ( .A(IR_REG_10__SCAN_IN), .ZN(n2362) );
  OAI211_X1 U2304 ( .C1(n2970), .C2(n4222), .A(n2089), .B(1'b1), .ZN(n2086) );
  OAI21_X1 U2306 ( .B1(n2158), .B2(n2155), .A(n2042), .ZN(n2154) );
  INV_X1 U2307 ( .A(n2458), .ZN(n2155) );
  NAND4_X1 U2308 ( .A1(n2203), .A2(n2202), .A3(n2301), .A4(n2297), .ZN(n2204)
         );
  INV_X1 U2309 ( .A(IR_REG_6__SCAN_IN), .ZN(n2202) );
  NOR2_X1 U2310 ( .A1(IR_REG_8__SCAN_IN), .A2(IR_REG_7__SCAN_IN), .ZN(n2203)
         );
  INV_X1 U2311 ( .A(n3331), .ZN(n2116) );
  AND2_X1 U2312 ( .A1(n2605), .A2(n2603), .ZN(n2763) );
  OR2_X1 U2313 ( .A1(n2802), .A2(n3015), .ZN(n2111) );
  XNOR2_X1 U2314 ( .A(n2606), .B(n2763), .ZN(n2617) );
  OAI21_X1 U2315 ( .B1(n3060), .B2(n2798), .A(n2147), .ZN(n2606) );
  NAND2_X1 U2316 ( .A1(n2254), .A2(n2134), .ZN(n2147) );
  CLKBUF_X1 U2317 ( .A(n2246), .Z(n2255) );
  CLKBUF_X1 U2318 ( .A(n2245), .Z(n2823) );
  AND4_X1 U2319 ( .A1(n2412), .A2(n2411), .A3(n2410), .A4(n2409), .ZN(n3575)
         );
  NAND2_X1 U2320 ( .A1(n2182), .A2(n2181), .ZN(n2180) );
  INV_X1 U2321 ( .A(IR_REG_29__SCAN_IN), .ZN(n2181) );
  INV_X1 U2322 ( .A(n2183), .ZN(n2182) );
  OAI21_X1 U2323 ( .B1(n2520), .B2(n2151), .A(n2281), .ZN(n2150) );
  NAND2_X1 U2324 ( .A1(n3558), .A2(n2129), .ZN(n2128) );
  INV_X1 U2325 ( .A(n3557), .ZN(n2129) );
  INV_X1 U2326 ( .A(n3558), .ZN(n2130) );
  OAI21_X1 U2327 ( .B1(n3860), .B2(n2094), .A(n2960), .ZN(n2967) );
  INV_X1 U2328 ( .A(n3859), .ZN(n2094) );
  INV_X1 U2329 ( .A(n2268), .ZN(n2201) );
  NAND2_X1 U2330 ( .A1(n2089), .A2(n4222), .ZN(n2082) );
  NAND2_X1 U2331 ( .A1(n4210), .A2(REG2_REG_5__SCAN_IN), .ZN(n2091) );
  INV_X1 U2332 ( .A(n2084), .ZN(n2081) );
  NAND2_X1 U2333 ( .A1(n2091), .A2(n2085), .ZN(n2084) );
  INV_X1 U2334 ( .A(n2992), .ZN(n2078) );
  OR2_X1 U2335 ( .A1(n3869), .A2(n2061), .ZN(n2060) );
  AND2_X1 U2336 ( .A1(n4207), .A2(REG1_REG_11__SCAN_IN), .ZN(n2061) );
  INV_X1 U2337 ( .A(n2159), .ZN(n2157) );
  NOR2_X1 U2338 ( .A1(n3579), .A2(n3648), .ZN(n2106) );
  NAND2_X1 U2339 ( .A1(n3413), .A2(n3391), .ZN(n2384) );
  NOR2_X1 U2340 ( .A1(n2376), .A2(n2043), .ZN(n2163) );
  AND2_X1 U2341 ( .A1(n3429), .A2(n2187), .ZN(n2178) );
  INV_X1 U2342 ( .A(n3180), .ZN(n3318) );
  AND2_X1 U2343 ( .A1(n2218), .A2(n2219), .ZN(n2186) );
  NOR2_X1 U2344 ( .A1(IR_REG_18__SCAN_IN), .A2(IR_REG_9__SCAN_IN), .ZN(n2146)
         );
  OR2_X1 U2345 ( .A1(n2657), .A2(n3143), .ZN(n3169) );
  NAND2_X1 U2346 ( .A1(n2696), .A2(n2695), .ZN(n2699) );
  AND2_X1 U2347 ( .A1(n3573), .A2(n2140), .ZN(n2139) );
  NAND2_X1 U2348 ( .A1(n2698), .A2(n3639), .ZN(n2140) );
  OR2_X1 U2349 ( .A1(n3159), .A2(n3160), .ZN(n2145) );
  AOI21_X1 U2350 ( .B1(n2030), .B2(n3259), .A(n2016), .ZN(n2119) );
  INV_X1 U2351 ( .A(n3619), .ZN(n2740) );
  NOR2_X1 U2352 ( .A1(n2354), .A2(n3251), .ZN(n2365) );
  AOI21_X1 U2353 ( .B1(n3832), .B2(n2774), .A(n2132), .ZN(n2675) );
  INV_X1 U2354 ( .A(n2110), .ZN(n2616) );
  NAND2_X1 U2355 ( .A1(n3559), .A2(n3557), .ZN(n2126) );
  AND4_X1 U2356 ( .A1(n2370), .A2(n2369), .A3(n2368), .A4(n2367), .ZN(n2679)
         );
  XNOR2_X1 U2357 ( .A(n4211), .B(REG2_REG_2__SCAN_IN), .ZN(n3860) );
  NAND2_X1 U2358 ( .A1(n3862), .A2(n2955), .ZN(n2974) );
  NOR2_X1 U2359 ( .A1(n2075), .A2(n3290), .ZN(n2072) );
  NAND2_X1 U2360 ( .A1(n2078), .A2(n3192), .ZN(n2076) );
  AND2_X1 U2361 ( .A1(n4208), .A2(REG2_REG_7__SCAN_IN), .ZN(n2992) );
  NOR2_X1 U2362 ( .A1(n3025), .A2(n3024), .ZN(n3023) );
  INV_X1 U2363 ( .A(n2057), .ZN(n3197) );
  OAI21_X1 U2364 ( .B1(n3195), .B2(n4231), .A(n2055), .ZN(n2057) );
  INV_X1 U2365 ( .A(n2056), .ZN(n2055) );
  OAI21_X1 U2366 ( .B1(n3194), .B2(n4231), .A(n2047), .ZN(n2056) );
  NOR2_X1 U2367 ( .A1(n3201), .A2(n3200), .ZN(n3869) );
  NAND2_X1 U2368 ( .A1(n3882), .A2(n3883), .ZN(n3884) );
  XNOR2_X1 U2369 ( .A(n2060), .B(n3885), .ZN(n4251) );
  NOR2_X1 U2370 ( .A1(n4251), .A2(n4252), .ZN(n4250) );
  XNOR2_X1 U2371 ( .A(n3890), .B(n3875), .ZN(n4298) );
  NOR2_X1 U2372 ( .A1(n4286), .A2(n2095), .ZN(n3890) );
  AND2_X1 U2373 ( .A1(n4347), .A2(REG2_REG_15__SCAN_IN), .ZN(n2095) );
  NAND2_X1 U2374 ( .A1(n4298), .A2(n4297), .ZN(n4296) );
  NAND2_X1 U2375 ( .A1(n4299), .A2(n3877), .ZN(n4311) );
  NAND2_X1 U2376 ( .A1(n4311), .A2(n4312), .ZN(n4310) );
  NAND2_X1 U2377 ( .A1(n3921), .A2(n3920), .ZN(n4110) );
  AND3_X1 U2378 ( .A1(n2786), .A2(n2785), .A3(n2784), .ZN(n3761) );
  NAND2_X1 U2379 ( .A1(n2160), .A2(n2020), .ZN(n2158) );
  NAND2_X1 U2380 ( .A1(n2162), .A2(n2020), .ZN(n2159) );
  AND4_X1 U2381 ( .A1(n2464), .A2(n2463), .A3(n2462), .A4(n2461), .ZN(n4029)
         );
  NAND2_X1 U2382 ( .A1(n4064), .A2(n4071), .ZN(n4063) );
  AOI21_X1 U2383 ( .B1(n3455), .B2(n2417), .A(n2416), .ZN(n3471) );
  INV_X1 U2384 ( .A(n3833), .ZN(n3345) );
  AND2_X1 U2385 ( .A1(n2525), .A2(n3725), .ZN(n3770) );
  OR2_X1 U2386 ( .A1(n3230), .A2(n2317), .ZN(n2185) );
  INV_X1 U2387 ( .A(n3232), .ZN(n3238) );
  INV_X1 U2388 ( .A(n4373), .ZN(n2586) );
  NOR2_X1 U2389 ( .A1(n3214), .A2(n3215), .ZN(n3239) );
  AND2_X1 U2390 ( .A1(n2555), .A2(n2554), .ZN(n3031) );
  NOR2_X1 U2391 ( .A1(n2027), .A2(n3760), .ZN(n3516) );
  NOR3_X1 U2392 ( .A1(n4034), .A2(n2108), .A3(n2109), .ZN(n3953) );
  NAND2_X1 U2393 ( .A1(n3978), .A2(n3955), .ZN(n2108) );
  AND2_X1 U2394 ( .A1(n4066), .A2(n4069), .ZN(n4067) );
  NOR2_X1 U2395 ( .A1(n3306), .A2(n3312), .ZN(n3348) );
  NAND2_X1 U2396 ( .A1(n4380), .A2(n4414), .ZN(n4400) );
  OR2_X1 U2397 ( .A1(n3014), .A2(n4206), .ZN(n4413) );
  AND2_X1 U2398 ( .A1(n2604), .A2(n4340), .ZN(n2927) );
  INV_X1 U2399 ( .A(IR_REG_25__SCAN_IN), .ZN(n2221) );
  INV_X1 U2400 ( .A(n2562), .ZN(n2222) );
  XNOR2_X1 U2401 ( .A(n2503), .B(n2502), .ZN(n2508) );
  NAND2_X1 U2402 ( .A1(n2501), .A2(IR_REG_31__SCAN_IN), .ZN(n2503) );
  NAND2_X1 U2403 ( .A1(n2559), .A2(n2102), .ZN(n2101) );
  NOR2_X1 U2404 ( .A1(IR_REG_0__SCAN_IN), .A2(IR_REG_1__SCAN_IN), .ZN(n2267)
         );
  NAND2_X1 U2405 ( .A1(n2064), .A2(n2063), .ZN(n2062) );
  NAND2_X1 U2406 ( .A1(IR_REG_0__SCAN_IN), .A2(IR_REG_31__SCAN_IN), .ZN(n2063)
         );
  NAND2_X1 U2407 ( .A1(n3843), .A2(n3844), .ZN(n3842) );
  XNOR2_X1 U2408 ( .A(n4211), .B(n2952), .ZN(n3864) );
  NAND2_X1 U2409 ( .A1(n3863), .A2(n3864), .ZN(n3862) );
  XNOR2_X1 U2410 ( .A(n3184), .B(n4249), .ZN(n4246) );
  NAND2_X1 U2411 ( .A1(n3189), .A2(n3188), .ZN(n3882) );
  AND2_X1 U2412 ( .A1(n2945), .A2(n2940), .ZN(n4320) );
  NAND2_X1 U2413 ( .A1(n4110), .A2(n3922), .ZN(n4117) );
  OR2_X1 U2414 ( .A1(n3921), .A2(n3920), .ZN(n3922) );
  XNOR2_X1 U2415 ( .A(n2175), .B(n2174), .ZN(n4116) );
  INV_X1 U2416 ( .A(n3910), .ZN(n2174) );
  AOI21_X1 U2417 ( .B1(n2170), .B2(n2173), .A(n2046), .ZN(n2168) );
  XNOR2_X1 U2418 ( .A(n3906), .B(n3905), .ZN(n3521) );
  NAND2_X1 U2419 ( .A1(n2169), .A2(n2854), .ZN(n3906) );
  AOI21_X1 U2420 ( .B1(n2842), .B2(n2872), .A(n2871), .ZN(n2874) );
  XNOR2_X1 U2421 ( .A(n2499), .B(n3785), .ZN(n3936) );
  NAND2_X1 U2422 ( .A1(n2491), .A2(n2845), .ZN(n2499) );
  INV_X1 U2423 ( .A(IR_REG_17__SCAN_IN), .ZN(n2213) );
  XNOR2_X1 U2424 ( .A(n2619), .B(n2763), .ZN(n2623) );
  OAI22_X1 U2425 ( .A1(n3138), .A2(n2799), .B1(n3052), .B2(n2798), .ZN(n2619)
         );
  INV_X1 U2426 ( .A(n4265), .ZN(n2093) );
  AOI21_X1 U2427 ( .B1(n4351), .B2(REG1_REG_13__SCAN_IN), .A(n4260), .ZN(n3873) );
  NOR2_X1 U2428 ( .A1(n4284), .A2(n3874), .ZN(n3876) );
  AND2_X1 U2429 ( .A1(n4347), .A2(REG1_REG_15__SCAN_IN), .ZN(n3874) );
  INV_X1 U2430 ( .A(n3579), .ZN(n2701) );
  NAND2_X1 U2431 ( .A1(n3840), .A2(n3060), .ZN(n3699) );
  NAND2_X1 U2432 ( .A1(n3015), .A2(n2602), .ZN(n3702) );
  OR2_X1 U2433 ( .A1(n4004), .A2(n3996), .ZN(n2109) );
  OAI21_X1 U2434 ( .B1(n3067), .B2(n2149), .A(n2148), .ZN(n4371) );
  NAND2_X1 U2435 ( .A1(n2280), .A2(n2273), .ZN(n2149) );
  NAND2_X1 U2436 ( .A1(n2150), .A2(n2280), .ZN(n2148) );
  NAND2_X1 U2437 ( .A1(n4371), .A2(n4375), .ZN(n4370) );
  NAND2_X1 U2438 ( .A1(n2184), .A2(n2229), .ZN(n2183) );
  INV_X1 U2439 ( .A(n2227), .ZN(n2184) );
  OAI22_X1 U2440 ( .A1(n3462), .A2(n2802), .B1(n2799), .B2(n2408), .ZN(n3356)
         );
  OR2_X1 U2441 ( .A1(n2893), .A2(n2128), .ZN(n2127) );
  NAND2_X1 U2442 ( .A1(n2253), .A2(n2252), .ZN(n2602) );
  NAND2_X1 U2443 ( .A1(n2939), .A2(DATAI_1_), .ZN(n2253) );
  NAND2_X1 U2444 ( .A1(n2251), .A2(n4212), .ZN(n2252) );
  INV_X1 U2445 ( .A(n2939), .ZN(n2251) );
  OAI22_X1 U2446 ( .A1(n2643), .A2(n2799), .B1(n2798), .B2(n2645), .ZN(n2644)
         );
  XNOR2_X1 U2447 ( .A(n2629), .B(n2800), .ZN(n2631) );
  NAND2_X1 U2448 ( .A1(n3159), .A2(n3160), .ZN(n2144) );
  AND2_X1 U2449 ( .A1(n2452), .A2(REG3_REG_20__SCAN_IN), .ZN(n2459) );
  NOR2_X1 U2450 ( .A1(n2441), .A2(n2440), .ZN(n2452) );
  NAND2_X1 U2451 ( .A1(n3606), .A2(n3607), .ZN(n3605) );
  NAND2_X1 U2452 ( .A1(n2459), .A2(REG3_REG_21__SCAN_IN), .ZN(n2467) );
  INV_X1 U2453 ( .A(n2698), .ZN(n2137) );
  INV_X1 U2454 ( .A(n2699), .ZN(n2138) );
  OR2_X1 U2455 ( .A1(n2598), .A2(IR_REG_27__SCAN_IN), .ZN(n2225) );
  AOI21_X1 U2456 ( .B1(n2598), .B2(IR_REG_28__SCAN_IN), .A(n2194), .ZN(n2224)
         );
  NAND4_X1 U2457 ( .A1(n2250), .A2(n2249), .A3(n2248), .A4(n2247), .ZN(n2254)
         );
  XNOR2_X1 U2458 ( .A(n2970), .B(n2977), .ZN(n4217) );
  OAI211_X1 U2459 ( .C1(n2970), .C2(n2080), .A(n2079), .B(n2031), .ZN(n2989)
         );
  AOI21_X1 U2460 ( .B1(n2082), .B2(n2091), .A(n2081), .ZN(n2080) );
  INV_X1 U2461 ( .A(n2076), .ZN(n2066) );
  AND2_X1 U2462 ( .A1(n2349), .A2(n2212), .ZN(n2436) );
  INV_X1 U2463 ( .A(REG3_REG_10__SCAN_IN), .ZN(n3251) );
  NOR2_X1 U2464 ( .A1(n3198), .A2(n4240), .ZN(n3201) );
  OR3_X1 U2465 ( .A1(n2394), .A2(IR_REG_11__SCAN_IN), .A3(IR_REG_12__SCAN_IN), 
        .ZN(n2396) );
  INV_X1 U2466 ( .A(n2060), .ZN(n3870) );
  NOR2_X1 U2467 ( .A1(n2396), .A2(IR_REG_13__SCAN_IN), .ZN(n2414) );
  OAI22_X1 U2468 ( .A1(n4274), .A2(n2058), .B1(n2024), .B2(n4285), .ZN(n4284)
         );
  OR2_X1 U2469 ( .A1(n4285), .A2(n4275), .ZN(n2058) );
  OR2_X1 U2470 ( .A1(n4274), .A2(n4275), .ZN(n2059) );
  NAND2_X1 U2471 ( .A1(n4310), .A2(n2054), .ZN(n4323) );
  NAND2_X1 U2472 ( .A1(n2447), .A2(IR_REG_31__SCAN_IN), .ZN(n2449) );
  NOR2_X1 U2473 ( .A1(n4323), .A2(n4322), .ZN(n4324) );
  NOR2_X1 U2474 ( .A1(n4110), .A2(n4113), .ZN(n4109) );
  NOR2_X1 U2475 ( .A1(n2172), .A2(n2171), .ZN(n2170) );
  INV_X1 U2476 ( .A(n3905), .ZN(n2171) );
  NOR2_X1 U2477 ( .A1(n2853), .A2(n2173), .ZN(n2172) );
  INV_X1 U2478 ( .A(n2854), .ZN(n2173) );
  AND3_X1 U2479 ( .A1(n2797), .A2(n2796), .A3(n2795), .ZN(n3916) );
  INV_X1 U2480 ( .A(n2152), .ZN(n4001) );
  NAND2_X1 U2481 ( .A1(n2157), .A2(n2458), .ZN(n2156) );
  INV_X1 U2482 ( .A(n2154), .ZN(n2153) );
  AND4_X1 U2483 ( .A1(n2473), .A2(n2472), .A3(n2471), .A4(n2470), .ZN(n4007)
         );
  NAND2_X1 U2484 ( .A1(n2429), .A2(REG3_REG_17__SCAN_IN), .ZN(n2431) );
  CLKBUF_X1 U2485 ( .A(n4020), .Z(n4085) );
  NAND2_X1 U2486 ( .A1(n2177), .A2(n2176), .ZN(n3455) );
  AOI21_X1 U2487 ( .B1(n2178), .B2(n2197), .A(n2045), .ZN(n2176) );
  OR2_X1 U2488 ( .A1(n2388), .A2(n2235), .ZN(n2400) );
  NOR2_X1 U2489 ( .A1(n2400), .A2(n4485), .ZN(n2418) );
  NAND2_X1 U2490 ( .A1(n2365), .A2(REG3_REG_11__SCAN_IN), .ZN(n2388) );
  AND2_X1 U2491 ( .A1(n2200), .A2(n2352), .ZN(n2165) );
  AND2_X1 U2492 ( .A1(n2374), .A2(n3364), .ZN(n3365) );
  AND4_X1 U2493 ( .A1(n2333), .A2(n2332), .A3(n2331), .A4(n2330), .ZN(n3319)
         );
  AND4_X1 U2494 ( .A1(n2325), .A2(n2324), .A3(n2323), .A4(n2322), .ZN(n3286)
         );
  INV_X1 U2495 ( .A(n4387), .ZN(n4049) );
  OR2_X1 U2496 ( .A1(n2320), .A2(n2319), .ZN(n2343) );
  INV_X1 U2497 ( .A(REG3_REG_5__SCAN_IN), .ZN(n2289) );
  NOR2_X1 U2498 ( .A1(n2290), .A2(n2289), .ZN(n2309) );
  AND4_X1 U2499 ( .A1(n2285), .A2(n2284), .A3(n2283), .A4(n2282), .ZN(n3211)
         );
  NAND2_X1 U2500 ( .A1(n3067), .A2(n2520), .ZN(n3068) );
  OR2_X1 U2501 ( .A1(n4413), .A2(n4592), .ZN(n2607) );
  INV_X1 U2502 ( .A(n4379), .ZN(n4089) );
  OR2_X1 U2503 ( .A1(n2956), .A2(n2811), .ZN(n4093) );
  INV_X1 U2504 ( .A(n4112), .ZN(n4377) );
  AND2_X1 U2505 ( .A1(n2807), .A2(n2199), .ZN(n2591) );
  NOR3_X1 U2506 ( .A1(n2589), .A2(n3904), .A3(n2107), .ZN(n3921) );
  OR2_X1 U2507 ( .A1(n2899), .A2(n3760), .ZN(n2107) );
  NOR3_X1 U2508 ( .A1(n4034), .A2(n2109), .A3(n3971), .ZN(n3976) );
  OR2_X1 U2509 ( .A1(n4056), .A2(n3802), .ZN(n4034) );
  NAND2_X1 U2510 ( .A1(n4067), .A2(n4057), .ZN(n4056) );
  AND2_X1 U2511 ( .A1(n2106), .A2(n4096), .ZN(n2105) );
  NAND2_X1 U2512 ( .A1(n2179), .A2(n2178), .ZN(n3428) );
  OR2_X1 U2513 ( .A1(n3405), .A2(n2197), .ZN(n2179) );
  NOR2_X1 U2514 ( .A1(n3418), .A2(n3411), .ZN(n3419) );
  NAND2_X1 U2515 ( .A1(n3375), .A2(n3374), .ZN(n3390) );
  OR2_X1 U2516 ( .A1(n3390), .A2(n3385), .ZN(n3418) );
  AND2_X1 U2517 ( .A1(n3348), .A2(n2133), .ZN(n3375) );
  NAND2_X1 U2518 ( .A1(n3239), .A2(n2044), .ZN(n3306) );
  NAND2_X1 U2519 ( .A1(n3239), .A2(n2022), .ZN(n3317) );
  INV_X1 U2520 ( .A(n4400), .ZN(n4406) );
  NOR2_X1 U2521 ( .A1(n3076), .A2(n2272), .ZN(n3096) );
  NOR2_X1 U2522 ( .A1(IR_REG_24__SCAN_IN), .A2(IR_REG_23__SCAN_IN), .ZN(n2220)
         );
  INV_X1 U2523 ( .A(IR_REG_21__SCAN_IN), .ZN(n2218) );
  AND2_X1 U2524 ( .A1(n2286), .A2(n2279), .ZN(n2973) );
  AND2_X1 U2525 ( .A1(n2658), .A2(n3169), .ZN(n2659) );
  AOI21_X1 U2526 ( .B1(n2014), .B2(n2115), .A(n2050), .ZN(n2114) );
  INV_X1 U2527 ( .A(n2025), .ZN(n2115) );
  AND2_X1 U2528 ( .A1(n3532), .A2(n3530), .ZN(n2750) );
  AND2_X1 U2529 ( .A1(n3248), .A2(n3249), .ZN(n2673) );
  NAND2_X1 U2530 ( .A1(n2143), .A2(n2141), .ZN(n3220) );
  NOR2_X1 U2531 ( .A1(n3223), .A2(n2142), .ZN(n2141) );
  INV_X1 U2532 ( .A(n2144), .ZN(n2142) );
  NAND2_X1 U2533 ( .A1(n2615), .A2(n2614), .ZN(n3039) );
  NAND2_X1 U2534 ( .A1(n3605), .A2(n3608), .ZN(n3550) );
  NAND2_X1 U2535 ( .A1(n2684), .A2(n3268), .ZN(n3261) );
  AND4_X1 U2536 ( .A1(n2490), .A2(n2489), .A3(n2488), .A4(n2487), .ZN(n3565)
         );
  INV_X1 U2537 ( .A(n2645), .ZN(n3215) );
  AND4_X1 U2538 ( .A1(n2423), .A2(n2422), .A3(n2421), .A4(n2420), .ZN(n4094)
         );
  AOI21_X1 U2539 ( .B1(n2139), .B2(n2023), .A(n2041), .ZN(n2135) );
  INV_X1 U2540 ( .A(n2139), .ZN(n2136) );
  NAND2_X1 U2541 ( .A1(n2143), .A2(n2144), .ZN(n3222) );
  OAI21_X1 U2542 ( .B1(n2939), .B2(n2112), .A(n2260), .ZN(n3085) );
  INV_X1 U2543 ( .A(n3642), .ZN(n3630) );
  INV_X1 U2544 ( .A(n4035), .ZN(n3802) );
  NAND2_X1 U2545 ( .A1(n2117), .A2(n2119), .ZN(n3333) );
  NAND2_X1 U2546 ( .A1(n2118), .A2(n2025), .ZN(n2117) );
  INV_X1 U2547 ( .A(n2684), .ZN(n2118) );
  OAI21_X1 U2548 ( .B1(n3606), .B2(n2124), .A(n2121), .ZN(n3618) );
  AOI21_X1 U2549 ( .B1(n2123), .B2(n2122), .A(n2038), .ZN(n2121) );
  INV_X1 U2550 ( .A(n3607), .ZN(n2122) );
  NOR2_X1 U2551 ( .A1(n2820), .A2(n2813), .ZN(n3609) );
  INV_X1 U2552 ( .A(n3644), .ZN(n3601) );
  NAND2_X1 U2553 ( .A1(n2126), .A2(n3558), .ZN(n2896) );
  AND3_X1 U2554 ( .A1(n2511), .A2(n2510), .A3(n2509), .ZN(n2512) );
  OAI211_X1 U2555 ( .C1(n3561), .C2(n2794), .A(n2497), .B(n2496), .ZN(n3949)
         );
  INV_X1 U2556 ( .A(n3565), .ZN(n3972) );
  INV_X1 U2557 ( .A(n4007), .ZN(n3823) );
  INV_X1 U2558 ( .A(n4075), .ZN(n3825) );
  INV_X1 U2559 ( .A(n3575), .ZN(n3827) );
  NAND4_X1 U2560 ( .A1(n2360), .A2(n2359), .A3(n2358), .A4(n2357), .ZN(n3832)
         );
  NAND4_X1 U2561 ( .A1(n2348), .A2(n2347), .A3(n2346), .A4(n2345), .ZN(n3833)
         );
  INV_X1 U2562 ( .A(n3319), .ZN(n3834) );
  INV_X1 U2563 ( .A(n3286), .ZN(n3835) );
  NAND2_X1 U2564 ( .A1(n2315), .A2(n2314), .ZN(n3836) );
  AND3_X1 U2565 ( .A1(n2313), .A2(n2312), .A3(n2311), .ZN(n2315) );
  AND2_X1 U2566 ( .A1(n2945), .A2(n2944), .ZN(n2957) );
  NAND2_X1 U2567 ( .A1(n3842), .A2(n2954), .ZN(n3863) );
  XNOR2_X1 U2568 ( .A(n2974), .B(n2965), .ZN(n2972) );
  AND2_X1 U2569 ( .A1(n2088), .A2(n2087), .ZN(n3004) );
  INV_X1 U2570 ( .A(n2090), .ZN(n2088) );
  NAND2_X1 U2571 ( .A1(n4217), .A2(REG2_REG_4__SCAN_IN), .ZN(n2087) );
  NOR2_X1 U2572 ( .A1(n2090), .A2(REG2_REG_4__SCAN_IN), .ZN(n2083) );
  NAND2_X1 U2573 ( .A1(n2998), .A2(n2997), .ZN(n3021) );
  NAND2_X1 U2574 ( .A1(n2067), .A2(n2066), .ZN(n2073) );
  OAI211_X1 U2575 ( .C1(n3023), .C2(n2070), .A(n2069), .B(n2068), .ZN(n4236)
         );
  NAND2_X1 U2576 ( .A1(n2992), .A2(n2077), .ZN(n2069) );
  NAND2_X1 U2577 ( .A1(n2072), .A2(n2076), .ZN(n2070) );
  NOR2_X1 U2578 ( .A1(n4232), .A2(n4231), .ZN(n4230) );
  AND2_X1 U2579 ( .A1(n3195), .A2(n3194), .ZN(n4232) );
  XNOR2_X1 U2580 ( .A(n3197), .B(n4249), .ZN(n4241) );
  NOR2_X1 U2581 ( .A1(n4241), .A2(n4242), .ZN(n4240) );
  NAND2_X1 U2582 ( .A1(n4245), .A2(n3185), .ZN(n3189) );
  XNOR2_X1 U2583 ( .A(n3884), .B(n4353), .ZN(n4257) );
  XNOR2_X1 U2584 ( .A(n3887), .B(n4350), .ZN(n4277) );
  NOR2_X1 U2585 ( .A1(n4277), .A2(n3440), .ZN(n4276) );
  NAND2_X1 U2586 ( .A1(n4296), .A2(n3891), .ZN(n4308) );
  AND2_X1 U2587 ( .A1(n2957), .A2(n3851), .ZN(n4314) );
  NOR2_X1 U2588 ( .A1(n4333), .A2(n2099), .ZN(n2098) );
  NAND2_X1 U2589 ( .A1(n4337), .A2(n4336), .ZN(n2099) );
  OAI21_X1 U2590 ( .B1(n2449), .B2(n2448), .A(n2501), .ZN(n3898) );
  AOI21_X1 U2591 ( .B1(n4331), .B2(REG1_REG_18__SCAN_IN), .A(n4324), .ZN(n3879) );
  INV_X1 U2592 ( .A(n4314), .ZN(n4321) );
  AND2_X1 U2593 ( .A1(n2783), .A2(n2792), .ZN(n3514) );
  OAI21_X1 U2594 ( .B1(n4064), .B2(n2159), .A(n2158), .ZN(n4019) );
  NAND2_X1 U2595 ( .A1(n4063), .A2(n2162), .ZN(n4043) );
  NAND2_X1 U2596 ( .A1(n2927), .A2(n2593), .ZN(n4590) );
  INV_X1 U2597 ( .A(n3770), .ZN(n2328) );
  NAND2_X1 U2598 ( .A1(n2185), .A2(n2318), .ZN(n3325) );
  OR2_X1 U2599 ( .A1(n3035), .A2(n2607), .ZN(n4101) );
  INV_X1 U2600 ( .A(n3085), .ZN(n2585) );
  OR2_X1 U2601 ( .A1(n4117), .A2(n4413), .ZN(n4119) );
  OR2_X1 U2602 ( .A1(n2232), .A2(n2559), .ZN(n2233) );
  AND2_X1 U2603 ( .A1(n2937), .A2(STATE_REG_SCAN_IN), .ZN(n4340) );
  INV_X1 U2604 ( .A(n3898), .ZN(n4592) );
  AND2_X1 U2605 ( .A1(n2381), .A2(n2373), .ZN(n4207) );
  INV_X1 U2606 ( .A(IR_REG_8__SCAN_IN), .ZN(n2337) );
  NOR2_X1 U2607 ( .A1(n2271), .A2(n2270), .ZN(n4211) );
  OAI21_X1 U2608 ( .B1(n2103), .B2(n2267), .A(n2101), .ZN(n2271) );
  NAND2_X1 U2609 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_2__SCAN_IN), .ZN(n2103)
         );
  NAND2_X1 U2610 ( .A1(n2100), .A2(n2096), .ZN(U3258) );
  INV_X1 U2611 ( .A(n2097), .ZN(n2096) );
  NAND2_X1 U2612 ( .A1(n4334), .A2(n4335), .ZN(n2100) );
  OAI21_X1 U2613 ( .B1(n4330), .B2(n4329), .A(n2098), .ZN(n2097) );
  MUX2_X1 U2614 ( .A(REG1_REG_28__SCAN_IN), .B(n2867), .S(n4433), .Z(n2863) );
  OR2_X1 U2615 ( .A1(n3931), .A2(n4159), .ZN(n2886) );
  MUX2_X1 U2616 ( .A(REG1_REG_26__SCAN_IN), .B(n2888), .S(n4433), .Z(n2883) );
  MUX2_X1 U2617 ( .A(n4127), .B(n4126), .S(n4433), .Z(n4128) );
  MUX2_X1 U2618 ( .A(REG0_REG_28__SCAN_IN), .B(n2867), .S(n4419), .Z(n2868) );
  OR2_X1 U2619 ( .A1(n3931), .A2(n4197), .ZN(n2890) );
  MUX2_X1 U2620 ( .A(REG0_REG_26__SCAN_IN), .B(n2888), .S(n4419), .Z(n2889) );
  OR2_X1 U2621 ( .A1(n4129), .A2(n4197), .ZN(n2587) );
  NOR2_X1 U2622 ( .A1(n2216), .A2(IR_REG_18__SCAN_IN), .ZN(n2013) );
  AND2_X1 U2623 ( .A1(n2119), .A2(n2116), .ZN(n2014) );
  INV_X1 U2624 ( .A(n2255), .ZN(n2308) );
  AND2_X1 U2625 ( .A1(n3841), .A2(n2134), .ZN(n2015) );
  AND2_X1 U2626 ( .A1(n3258), .A2(n2120), .ZN(n2016) );
  INV_X1 U2627 ( .A(IR_REG_9__SCAN_IN), .ZN(n2212) );
  AND2_X1 U2628 ( .A1(n2215), .A2(n2214), .ZN(n2017) );
  OR2_X1 U2629 ( .A1(n2072), .A2(n2077), .ZN(n2018) );
  INV_X1 U2630 ( .A(n2036), .ZN(n2089) );
  AND2_X1 U2631 ( .A1(n2328), .A2(n2318), .ZN(n2019) );
  NAND2_X1 U2632 ( .A1(n2138), .A2(n2137), .ZN(n3570) );
  OR2_X1 U2633 ( .A1(n4073), .A2(n3543), .ZN(n2020) );
  AND2_X1 U2634 ( .A1(n2164), .A2(n2166), .ZN(n2021) );
  AND2_X1 U2635 ( .A1(n3238), .A2(n3318), .ZN(n2022) );
  NOR2_X1 U2636 ( .A1(n2698), .A2(n3639), .ZN(n2023) );
  NAND2_X1 U2637 ( .A1(n3437), .A2(n3464), .ZN(n3463) );
  OR2_X1 U2638 ( .A1(n3873), .A2(n4350), .ZN(n2024) );
  AND4_X1 U2639 ( .A1(n2295), .A2(n2294), .A3(n2293), .A4(n2292), .ZN(n2643)
         );
  AOI21_X1 U2640 ( .B1(n3961), .B2(n2484), .A(n2483), .ZN(n2842) );
  OR2_X1 U2641 ( .A1(n3258), .A2(n3259), .ZN(n2025) );
  XOR2_X1 U2642 ( .A(n3191), .B(n3192), .Z(n2026) );
  XNOR2_X1 U2643 ( .A(n2287), .B(IR_REG_4__SCAN_IN), .ZN(n4222) );
  OR2_X1 U2644 ( .A1(n2589), .A2(n2899), .ZN(n2027) );
  AND4_X1 U2645 ( .A1(n2207), .A2(n2206), .A3(n2205), .A4(n2362), .ZN(n2215)
         );
  AND2_X1 U2646 ( .A1(n3840), .A2(n2602), .ZN(n2028) );
  INV_X1 U2647 ( .A(n3268), .ZN(n2120) );
  OR2_X1 U2648 ( .A1(n2897), .A2(n3650), .ZN(n2029) );
  OR2_X1 U2649 ( .A1(n2120), .A2(n3258), .ZN(n2030) );
  INV_X2 U2650 ( .A(n2799), .ZN(n2134) );
  OR2_X1 U2651 ( .A1(n2084), .A2(n4222), .ZN(n2031) );
  INV_X1 U2652 ( .A(n2273), .ZN(n2151) );
  INV_X1 U2653 ( .A(n2075), .ZN(n2074) );
  NOR2_X1 U2654 ( .A1(n2078), .A2(n3192), .ZN(n2075) );
  AND3_X1 U2655 ( .A1(n2017), .A2(n2217), .A3(n2013), .ZN(n2504) );
  NAND2_X1 U2656 ( .A1(n2504), .A2(n2218), .ZN(n2032) );
  INV_X1 U2657 ( .A(IR_REG_31__SCAN_IN), .ZN(n2559) );
  AND2_X1 U2658 ( .A1(n3886), .A2(n2093), .ZN(n2033) );
  AND2_X1 U2659 ( .A1(n2186), .A2(n2220), .ZN(n2034) );
  AND2_X1 U2660 ( .A1(n2059), .A2(n2024), .ZN(n2035) );
  INV_X1 U2661 ( .A(IR_REG_2__SCAN_IN), .ZN(n2102) );
  INV_X1 U2662 ( .A(IR_REG_1__SCAN_IN), .ZN(n2064) );
  NOR2_X1 U2663 ( .A1(n4034), .A2(n2109), .ZN(n3975) );
  NAND2_X1 U2664 ( .A1(n2353), .A2(n2352), .ZN(n3346) );
  XNOR2_X1 U2665 ( .A(n2338), .B(n2337), .ZN(n3192) );
  INV_X1 U2666 ( .A(n3192), .ZN(n2077) );
  OAI21_X1 U2667 ( .B1(n3629), .B2(n3626), .A(n3625), .ZN(n3539) );
  OAI21_X1 U2668 ( .B1(n2699), .B2(n2136), .A(n2135), .ZN(n3582) );
  INV_X1 U2669 ( .A(n3342), .ZN(n2133) );
  OR2_X1 U2670 ( .A1(n3548), .A2(n3547), .ZN(n2037) );
  AND2_X1 U2671 ( .A1(n3548), .A2(n3547), .ZN(n2038) );
  AND2_X1 U2672 ( .A1(n2179), .A2(n2187), .ZN(n2039) );
  OR2_X1 U2673 ( .A1(n4034), .A2(n4004), .ZN(n2040) );
  INV_X1 U2674 ( .A(n2663), .ZN(n3288) );
  NAND2_X1 U2675 ( .A1(n2062), .A2(n2065), .ZN(n2958) );
  INV_X1 U2676 ( .A(n3648), .ZN(n3464) );
  AND2_X1 U2677 ( .A1(n2704), .A2(n2703), .ZN(n2041) );
  OR2_X1 U2678 ( .A1(n3552), .A2(n4035), .ZN(n2042) );
  NOR2_X1 U2679 ( .A1(n3413), .A2(n3391), .ZN(n2043) );
  INV_X1 U2680 ( .A(n3462), .ZN(n3828) );
  AND4_X1 U2681 ( .A1(n2406), .A2(n2405), .A3(n2404), .A4(n2403), .ZN(n3462)
         );
  AND2_X1 U2682 ( .A1(n2022), .A2(n2663), .ZN(n2044) );
  AND2_X1 U2683 ( .A1(n3462), .A2(n2408), .ZN(n2045) );
  AND2_X1 U2684 ( .A1(n3903), .A2(n3904), .ZN(n2046) );
  NAND2_X1 U2685 ( .A1(n3196), .A2(REG1_REG_9__SCAN_IN), .ZN(n2047) );
  INV_X1 U2686 ( .A(n2124), .ZN(n2123) );
  NAND2_X1 U2687 ( .A1(n3608), .A2(n2037), .ZN(n2124) );
  NAND2_X1 U2688 ( .A1(n2699), .A2(n2698), .ZN(n3569) );
  AND2_X1 U2689 ( .A1(n3437), .A2(n2105), .ZN(n4066) );
  OAI21_X1 U2690 ( .B1(n4071), .B2(n2161), .A(n2451), .ZN(n2160) );
  INV_X1 U2691 ( .A(n2162), .ZN(n2161) );
  OR2_X1 U2692 ( .A1(n4090), .A2(n4072), .ZN(n2162) );
  NOR2_X1 U2693 ( .A1(n2893), .A2(n2130), .ZN(n2048) );
  AND2_X1 U2694 ( .A1(n2127), .A2(n2892), .ZN(n2049) );
  NAND2_X1 U2695 ( .A1(n2586), .A2(n4378), .ZN(n3214) );
  AOI21_X1 U2696 ( .B1(n3280), .B2(n2340), .A(n2339), .ZN(n3305) );
  NAND2_X1 U2697 ( .A1(n3324), .A2(n2329), .ZN(n3280) );
  AND2_X1 U2698 ( .A1(n3239), .A2(n3238), .ZN(n3240) );
  NAND2_X1 U2699 ( .A1(n3437), .A2(n2106), .ZN(n3479) );
  AND2_X1 U2700 ( .A1(n2690), .A2(n2689), .ZN(n2050) );
  AND2_X1 U2701 ( .A1(n3419), .A2(n2408), .ZN(n3437) );
  AOI21_X1 U2702 ( .B1(n2519), .B2(n3054), .A(n2028), .ZN(n3067) );
  OR2_X1 U2703 ( .A1(n4351), .A2(REG2_REG_13__SCAN_IN), .ZN(n2051) );
  AND2_X1 U2704 ( .A1(n2970), .A2(n4222), .ZN(n2090) );
  XNOR2_X1 U2705 ( .A(n2617), .B(n2110), .ZN(n3038) );
  NAND2_X1 U2706 ( .A1(n3068), .A2(n2273), .ZN(n3088) );
  NOR2_X1 U2707 ( .A1(n2228), .A2(n2227), .ZN(n2514) );
  NOR2_X1 U2708 ( .A1(n2086), .A2(n2083), .ZN(n2052) );
  NAND2_X1 U2709 ( .A1(n4340), .A2(n2821), .ZN(n2053) );
  OR2_X1 U2710 ( .A1(n3892), .A2(REG1_REG_17__SCAN_IN), .ZN(n2054) );
  INV_X1 U2711 ( .A(REG2_REG_4__SCAN_IN), .ZN(n2085) );
  INV_X1 U2712 ( .A(n2059), .ZN(n4273) );
  NAND3_X1 U2713 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .A3(
        IR_REG_1__SCAN_IN), .ZN(n2065) );
  INV_X2 U2714 ( .A(IR_REG_0__SCAN_IN), .ZN(n2112) );
  XNOR2_X1 U2715 ( .A(n3876), .B(n3875), .ZN(n4301) );
  NAND2_X1 U2716 ( .A1(n3023), .A2(n2018), .ZN(n2068) );
  NAND2_X1 U2717 ( .A1(n3023), .A2(n2077), .ZN(n2071) );
  INV_X1 U2718 ( .A(n3023), .ZN(n2067) );
  NAND3_X1 U2719 ( .A1(n2073), .A2(n2074), .A3(n2071), .ZN(n3183) );
  NAND2_X1 U2720 ( .A1(n4236), .A2(n4237), .ZN(n4235) );
  NAND3_X1 U2721 ( .A1(n2036), .A2(n2091), .A3(n2970), .ZN(n2079) );
  NAND2_X1 U2722 ( .A1(n4256), .A2(n2033), .ZN(n2092) );
  NAND2_X1 U2723 ( .A1(n2092), .A2(n2051), .ZN(n3887) );
  NAND2_X1 U2724 ( .A1(n4256), .A2(n3886), .ZN(n4268) );
  NAND3_X1 U2725 ( .A1(n2104), .A2(n2217), .A3(n2017), .ZN(n2562) );
  NOR2_X2 U2726 ( .A1(n2296), .A2(n2204), .ZN(n2217) );
  NAND3_X1 U2727 ( .A1(n2112), .A2(n2064), .A3(n2102), .ZN(n2268) );
  NAND2_X1 U2728 ( .A1(n2684), .A2(n2014), .ZN(n2113) );
  NAND2_X1 U2729 ( .A1(n2113), .A2(n2114), .ZN(n3354) );
  INV_X1 U2730 ( .A(n3618), .ZN(n2741) );
  NAND3_X1 U2731 ( .A1(n2760), .A2(n3593), .A3(n2048), .ZN(n2125) );
  NAND2_X1 U2732 ( .A1(n2760), .A2(n3593), .ZN(n3559) );
  NAND2_X1 U2733 ( .A1(n2125), .A2(n2049), .ZN(n2906) );
  NAND2_X1 U2734 ( .A1(n3760), .A2(n2134), .ZN(n2789) );
  AOI21_X1 U2735 ( .B1(n3085), .B2(n2134), .A(n2611), .ZN(n2612) );
  NAND2_X1 U2736 ( .A1(n2899), .A2(n2134), .ZN(n2775) );
  NAND2_X1 U2737 ( .A1(n3232), .A2(n2134), .ZN(n2641) );
  NAND2_X1 U2738 ( .A1(n3802), .A2(n2134), .ZN(n2731) );
  NAND2_X1 U2739 ( .A1(n3836), .A2(n2134), .ZN(n2639) );
  NAND2_X1 U2740 ( .A1(n4072), .A2(n2134), .ZN(n2713) );
  NAND2_X1 U2741 ( .A1(n4383), .A2(n2134), .ZN(n2628) );
  NAND2_X1 U2742 ( .A1(n3833), .A2(n2134), .ZN(n2666) );
  NAND2_X1 U2743 ( .A1(n4090), .A2(n2134), .ZN(n2711) );
  NAND2_X1 U2744 ( .A1(n3832), .A2(n2134), .ZN(n2669) );
  AOI22_X1 U2745 ( .A1(n2774), .A2(n4383), .B1(n2134), .B2(n3134), .ZN(n2632)
         );
  AOI22_X1 U2746 ( .A1(n2774), .A2(n3833), .B1(n2134), .B2(n3312), .ZN(n2671)
         );
  NOR2_X1 U2747 ( .A1(n2133), .A2(n2799), .ZN(n2132) );
  NAND2_X1 U2748 ( .A1(n4073), .A2(n2134), .ZN(n2720) );
  NAND2_X1 U2749 ( .A1(n4052), .A2(n2134), .ZN(n2729) );
  NAND2_X1 U2750 ( .A1(n3989), .A2(n2134), .ZN(n2743) );
  NAND2_X1 U2751 ( .A1(n3949), .A2(n2134), .ZN(n2762) );
  NAND2_X1 U2752 ( .A1(n3822), .A2(n2134), .ZN(n2772) );
  NAND2_X4 U2753 ( .A1(n2601), .A2(n2604), .ZN(n2799) );
  NAND2_X1 U2754 ( .A1(n3158), .A2(n2145), .ZN(n2143) );
  NAND3_X1 U2755 ( .A1(n2349), .A2(n2208), .A3(n2212), .ZN(n2210) );
  NAND3_X1 U2756 ( .A1(n2349), .A2(n2208), .A3(n2146), .ZN(n2447) );
  OAI21_X1 U2757 ( .B1(n4064), .B2(n2156), .A(n2153), .ZN(n2152) );
  NAND2_X1 U2758 ( .A1(n2353), .A2(n2165), .ZN(n2164) );
  NAND2_X1 U2759 ( .A1(n2164), .A2(n2163), .ZN(n2385) );
  INV_X1 U2760 ( .A(n2376), .ZN(n2166) );
  NAND2_X1 U2761 ( .A1(n3507), .A2(n2170), .ZN(n2167) );
  NAND2_X1 U2762 ( .A1(n2167), .A2(n2168), .ZN(n2175) );
  NAND2_X1 U2763 ( .A1(n3507), .A2(n2853), .ZN(n2169) );
  NAND2_X1 U2764 ( .A1(n3405), .A2(n2178), .ZN(n2177) );
  NOR2_X1 U2765 ( .A1(n2228), .A2(n2180), .ZN(n2232) );
  NAND2_X1 U2766 ( .A1(n2185), .A2(n2019), .ZN(n3324) );
  NOR2_X1 U2767 ( .A1(n2906), .A2(n2904), .ZN(n2816) );
  NAND2_X1 U2768 ( .A1(n4200), .A2(n2240), .ZN(n2246) );
  AND2_X1 U2769 ( .A1(n2957), .A2(n3855), .ZN(n4316) );
  OR2_X1 U2770 ( .A1(n3432), .A2(n3420), .ZN(n2187) );
  INV_X1 U2771 ( .A(n3420), .ZN(n3411) );
  INV_X1 U2772 ( .A(n3391), .ZN(n3385) );
  INV_X1 U2773 ( .A(n2520), .ZN(n3792) );
  NAND2_X1 U2774 ( .A1(n3647), .A2(n2899), .ZN(n2188) );
  AND2_X1 U2775 ( .A1(n4029), .A2(n4010), .ZN(n2189) );
  OR2_X1 U2776 ( .A1(n4094), .A2(n2701), .ZN(n2190) );
  OR2_X1 U2777 ( .A1(n3526), .A2(n4159), .ZN(n2191) );
  OR2_X1 U2778 ( .A1(n3526), .A2(n4197), .ZN(n2192) );
  INV_X1 U2779 ( .A(n3430), .ZN(n2408) );
  AND2_X1 U2780 ( .A1(n2817), .A2(n3609), .ZN(n2193) );
  AND2_X1 U2781 ( .A1(n2229), .A2(IR_REG_27__SCAN_IN), .ZN(n2194) );
  INV_X1 U2782 ( .A(n3413), .ZN(n3830) );
  AND4_X1 U2783 ( .A1(n2380), .A2(n2379), .A3(n2378), .A4(n2377), .ZN(n3413)
         );
  AND2_X1 U2784 ( .A1(n2836), .A2(n2835), .ZN(n2195) );
  AND2_X1 U2785 ( .A1(n3825), .A2(n4088), .ZN(n2196) );
  AND2_X1 U2786 ( .A1(n3432), .A2(n3420), .ZN(n2197) );
  INV_X1 U2787 ( .A(n3432), .ZN(n3829) );
  AND4_X1 U2788 ( .A1(n2393), .A2(n2392), .A3(n2391), .A4(n2390), .ZN(n3432)
         );
  NAND2_X2 U2789 ( .A1(n2924), .A2(n4200), .ZN(n2469) );
  OR2_X1 U2790 ( .A1(n3644), .A2(n2898), .ZN(n2198) );
  AND2_X1 U2791 ( .A1(n2927), .A2(n2831), .ZN(n2199) );
  NOR2_X1 U2792 ( .A1(n3363), .A2(n2375), .ZN(n2200) );
  NAND2_X1 U2793 ( .A1(n2530), .A2(n3733), .ZN(n3370) );
  AND2_X1 U2794 ( .A1(n2213), .A2(n2212), .ZN(n2214) );
  AND2_X1 U2795 ( .A1(n3943), .A2(n3779), .ZN(n3756) );
  NAND2_X1 U2796 ( .A1(n2529), .A2(n3720), .ZN(n3340) );
  NAND2_X1 U2797 ( .A1(n2541), .A2(n3745), .ZN(n4020) );
  INV_X1 U2798 ( .A(n2675), .ZN(n2676) );
  OR3_X1 U2799 ( .A1(n2782), .A2(n4571), .A3(n2781), .ZN(n2792) );
  INV_X1 U2800 ( .A(IR_REG_22__SCAN_IN), .ZN(n2219) );
  AND2_X1 U2801 ( .A1(n2418), .A2(n2236), .ZN(n2429) );
  OR2_X1 U2802 ( .A1(n2467), .A2(n2466), .ZN(n2476) );
  AND2_X1 U2803 ( .A1(n2485), .A2(REG3_REG_24__SCAN_IN), .ZN(n2492) );
  INV_X1 U2804 ( .A(n2924), .ZN(n2240) );
  INV_X1 U2805 ( .A(n4346), .ZN(n3875) );
  OR2_X1 U2806 ( .A1(n2431), .A2(n2237), .ZN(n2441) );
  OR2_X1 U2807 ( .A1(n2343), .A2(n2234), .ZN(n2354) );
  INV_X1 U2808 ( .A(n3271), .ZN(n3374) );
  INV_X1 U2809 ( .A(n3134), .ZN(n3095) );
  INV_X1 U2810 ( .A(REG3_REG_7__SCAN_IN), .ZN(n2319) );
  NOR2_X1 U2811 ( .A1(n2476), .A2(n2475), .ZN(n2485) );
  NAND2_X1 U2812 ( .A1(n3174), .A2(n2662), .ZN(n3158) );
  NAND2_X1 U2813 ( .A1(n2939), .A2(DATAI_0_), .ZN(n2260) );
  OR2_X1 U2814 ( .A1(n2830), .A2(n2822), .ZN(n3632) );
  OR2_X1 U2815 ( .A1(n2830), .A2(n2935), .ZN(n2820) );
  NAND2_X1 U2816 ( .A1(n2492), .A2(REG3_REG_25__SCAN_IN), .ZN(n2782) );
  INV_X2 U2817 ( .A(n2255), .ZN(n2478) );
  NOR2_X1 U2818 ( .A1(n3871), .A2(n4250), .ZN(n4262) );
  NOR2_X1 U2819 ( .A1(n3888), .A2(n4276), .ZN(n4288) );
  AND2_X1 U2820 ( .A1(n4332), .A2(n4331), .ZN(n4333) );
  INV_X1 U2821 ( .A(n2870), .ZN(n2871) );
  AOI21_X1 U2822 ( .B1(n4083), .B2(n2439), .A(n2196), .ZN(n4064) );
  AND2_X1 U2823 ( .A1(n3575), .A2(n3464), .ZN(n2416) );
  NAND2_X1 U2824 ( .A1(n3953), .A2(n2765), .ZN(n2589) );
  OR2_X1 U2825 ( .A1(n2326), .A2(IR_REG_6__SCAN_IN), .ZN(n2327) );
  INV_X1 U2826 ( .A(n4057), .ZN(n3543) );
  INV_X1 U2827 ( .A(n4069), .ZN(n4072) );
  INV_X1 U2828 ( .A(n3053), .ZN(n3647) );
  INV_X1 U2829 ( .A(n2823), .ZN(n2794) );
  AND4_X1 U2830 ( .A1(n2435), .A2(n2434), .A3(n2433), .A4(n2432), .ZN(n4075)
         );
  NAND2_X1 U2831 ( .A1(n2026), .A2(REG1_REG_8__SCAN_IN), .ZN(n3195) );
  NAND2_X1 U2832 ( .A1(n4246), .A2(REG2_REG_10__SCAN_IN), .ZN(n4245) );
  AND2_X1 U2833 ( .A1(n2957), .A2(n2956), .ZN(n4332) );
  AND2_X1 U2834 ( .A1(n3381), .A2(n3383), .ZN(n3791) );
  INV_X1 U2835 ( .A(n4101), .ZN(n4213) );
  AND2_X1 U2836 ( .A1(n4119), .A2(n4118), .ZN(n4120) );
  INV_X1 U2837 ( .A(n3948), .ZN(n3955) );
  INV_X1 U2838 ( .A(n4004), .ZN(n4010) );
  INV_X1 U2839 ( .A(n4088), .ZN(n4096) );
  INV_X1 U2840 ( .A(n3419), .ZN(n3436) );
  INV_X1 U2841 ( .A(n4413), .ZN(n4411) );
  AND2_X1 U2842 ( .A1(n2580), .A2(n2591), .ZN(n2862) );
  INV_X1 U2843 ( .A(n4249), .ZN(n4354) );
  INV_X1 U2844 ( .A(n2272), .ZN(n3052) );
  INV_X1 U2845 ( .A(n3609), .ZN(n3650) );
  NAND2_X1 U2846 ( .A1(n2513), .A2(n2512), .ZN(n3822) );
  NAND4_X1 U2847 ( .A1(n2244), .A2(n2243), .A3(n2242), .A4(n2241), .ZN(n4090)
         );
  INV_X1 U2848 ( .A(n3211), .ZN(n3838) );
  INV_X1 U2849 ( .A(n2973), .ZN(n2965) );
  OR2_X1 U2850 ( .A1(n2364), .A2(n2363), .ZN(n4249) );
  INV_X1 U2851 ( .A(n4332), .ZN(n4319) );
  INV_X1 U2852 ( .A(n3397), .ZN(n4104) );
  OR2_X1 U2853 ( .A1(n3035), .A2(n3030), .ZN(n3445) );
  INV_X1 U2854 ( .A(n4433), .ZN(n4431) );
  INV_X1 U2855 ( .A(n4419), .ZN(n4418) );
  INV_X1 U2856 ( .A(n4204), .ZN(n2930) );
  XNOR2_X1 U2857 ( .A(n2561), .B(IR_REG_24__SCAN_IN), .ZN(n4204) );
  INV_X1 U2858 ( .A(n3885), .ZN(n4353) );
  XNOR2_X1 U2859 ( .A(n2335), .B(IR_REG_7__SCAN_IN), .ZN(n4208) );
  INV_X1 U2860 ( .A(REG0_REG_25__SCAN_IN), .ZN(n2584) );
  NAND2_X1 U2861 ( .A1(n2201), .A2(n4525), .ZN(n2296) );
  AND2_X1 U2862 ( .A1(n2215), .A2(n2213), .ZN(n2208) );
  NAND2_X1 U2863 ( .A1(n2210), .A2(IR_REG_31__SCAN_IN), .ZN(n2209) );
  MUX2_X1 U2864 ( .A(IR_REG_31__SCAN_IN), .B(n2209), .S(IR_REG_18__SCAN_IN), 
        .Z(n2211) );
  AND2_X1 U2865 ( .A1(n2211), .A2(n2447), .ZN(n4331) );
  INV_X1 U2866 ( .A(n4331), .ZN(n4342) );
  INV_X1 U2867 ( .A(DATAI_18_), .ZN(n4341) );
  NAND2_X1 U2868 ( .A1(n2448), .A2(n2502), .ZN(n2216) );
  NAND2_X1 U2869 ( .A1(n2222), .A2(n2221), .ZN(n2228) );
  INV_X1 U2870 ( .A(IR_REG_26__SCAN_IN), .ZN(n2223) );
  INV_X1 U2871 ( .A(IR_REG_28__SCAN_IN), .ZN(n2229) );
  NAND2_X4 U2872 ( .A1(n2225), .A2(n2224), .ZN(n2939) );
  MUX2_X1 U2873 ( .A(n4342), .B(n4341), .S(n2939), .Z(n4069) );
  INV_X1 U2874 ( .A(IR_REG_27__SCAN_IN), .ZN(n2226) );
  NAND2_X1 U2875 ( .A1(n2223), .A2(n2226), .ZN(n2227) );
  NAND2_X1 U2876 ( .A1(n2517), .A2(IR_REG_31__SCAN_IN), .ZN(n2230) );
  INV_X1 U2877 ( .A(n2232), .ZN(n3505) );
  NAND2_X1 U2878 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .ZN(
        n2290) );
  NAND2_X1 U2879 ( .A1(n2309), .A2(REG3_REG_6__SCAN_IN), .ZN(n2320) );
  NAND2_X1 U2880 ( .A1(REG3_REG_8__SCAN_IN), .A2(REG3_REG_9__SCAN_IN), .ZN(
        n2234) );
  NAND2_X1 U2881 ( .A1(REG3_REG_12__SCAN_IN), .A2(REG3_REG_13__SCAN_IN), .ZN(
        n2235) );
  INV_X1 U2882 ( .A(REG3_REG_14__SCAN_IN), .ZN(n4485) );
  AND2_X1 U2883 ( .A1(REG3_REG_16__SCAN_IN), .A2(REG3_REG_15__SCAN_IN), .ZN(
        n2236) );
  INV_X1 U2884 ( .A(REG3_REG_18__SCAN_IN), .ZN(n2237) );
  NAND2_X1 U2885 ( .A1(n2431), .A2(n2237), .ZN(n2238) );
  NAND2_X1 U2886 ( .A1(n2441), .A2(n2238), .ZN(n4078) );
  OR2_X1 U2887 ( .A1(n2469), .A2(n4078), .ZN(n2244) );
  INV_X1 U2888 ( .A(n4200), .ZN(n2239) );
  AND2_X2 U2889 ( .A1(n2239), .A2(n2924), .ZN(n2261) );
  NAND2_X1 U2890 ( .A1(n3667), .A2(REG1_REG_18__SCAN_IN), .ZN(n2243) );
  NAND2_X1 U2891 ( .A1(n3668), .A2(REG0_REG_18__SCAN_IN), .ZN(n2242) );
  NAND2_X1 U2892 ( .A1(n2478), .A2(REG2_REG_18__SCAN_IN), .ZN(n2241) );
  INV_X1 U2893 ( .A(n2469), .ZN(n2245) );
  NAND2_X1 U2894 ( .A1(n2245), .A2(REG3_REG_1__SCAN_IN), .ZN(n2250) );
  NAND2_X1 U2895 ( .A1(n2262), .A2(REG0_REG_1__SCAN_IN), .ZN(n2249) );
  NAND2_X1 U2896 ( .A1(n2261), .A2(REG1_REG_1__SCAN_IN), .ZN(n2248) );
  INV_X1 U2897 ( .A(REG2_REG_1__SCAN_IN), .ZN(n3062) );
  OR2_X1 U2898 ( .A1(n2246), .A2(n3062), .ZN(n2247) );
  INV_X1 U2899 ( .A(n2958), .ZN(n4212) );
  NAND2_X1 U2900 ( .A1(n3699), .A2(n3702), .ZN(n2519) );
  NAND2_X1 U2901 ( .A1(n2245), .A2(REG3_REG_0__SCAN_IN), .ZN(n2259) );
  NAND2_X1 U2902 ( .A1(n2262), .A2(REG0_REG_0__SCAN_IN), .ZN(n2258) );
  NAND2_X1 U2903 ( .A1(n2308), .A2(REG2_REG_0__SCAN_IN), .ZN(n2257) );
  NAND2_X1 U2904 ( .A1(n2261), .A2(REG1_REG_0__SCAN_IN), .ZN(n2256) );
  NAND4_X2 U2905 ( .A1(n2259), .A2(n2258), .A3(n2257), .A4(n2256), .ZN(n3841)
         );
  AND2_X1 U2906 ( .A1(n3841), .A2(n3085), .ZN(n3054) );
  NAND2_X1 U2907 ( .A1(n2261), .A2(REG1_REG_2__SCAN_IN), .ZN(n2266) );
  NAND2_X1 U2908 ( .A1(n2308), .A2(REG2_REG_2__SCAN_IN), .ZN(n2265) );
  NAND2_X1 U2909 ( .A1(n2262), .A2(REG0_REG_2__SCAN_IN), .ZN(n2264) );
  NAND2_X1 U2910 ( .A1(n2245), .A2(REG3_REG_2__SCAN_IN), .ZN(n2263) );
  INV_X1 U2911 ( .A(n3138), .ZN(n3839) );
  INV_X1 U2912 ( .A(n2269), .ZN(n2270) );
  MUX2_X1 U2913 ( .A(n4211), .B(DATAI_2_), .S(n2939), .Z(n2272) );
  NAND2_X1 U2914 ( .A1(n3839), .A2(n3052), .ZN(n3706) );
  NAND2_X1 U2915 ( .A1(n3138), .A2(n2272), .ZN(n3703) );
  NAND2_X1 U2916 ( .A1(n3138), .A2(n3052), .ZN(n2273) );
  OR2_X1 U2917 ( .A1(n2469), .A2(REG3_REG_3__SCAN_IN), .ZN(n2277) );
  NAND2_X1 U2918 ( .A1(n3668), .A2(REG0_REG_3__SCAN_IN), .ZN(n2276) );
  NAND2_X1 U2919 ( .A1(n2478), .A2(REG2_REG_3__SCAN_IN), .ZN(n2275) );
  NAND2_X1 U2920 ( .A1(n2261), .A2(REG1_REG_3__SCAN_IN), .ZN(n2274) );
  NAND2_X1 U2921 ( .A1(n2269), .A2(IR_REG_31__SCAN_IN), .ZN(n2278) );
  INV_X1 U2922 ( .A(IR_REG_3__SCAN_IN), .ZN(n4525) );
  NAND2_X1 U2923 ( .A1(n2278), .A2(n4525), .ZN(n2286) );
  OR2_X1 U2924 ( .A1(n2278), .A2(n4525), .ZN(n2279) );
  MUX2_X1 U2925 ( .A(n2973), .B(DATAI_3_), .S(n2939), .Z(n3134) );
  NAND2_X1 U2926 ( .A1(n4383), .A2(n3134), .ZN(n2281) );
  NAND2_X1 U2927 ( .A1(n2261), .A2(REG1_REG_4__SCAN_IN), .ZN(n2285) );
  NAND2_X1 U2928 ( .A1(n3668), .A2(REG0_REG_4__SCAN_IN), .ZN(n2284) );
  NAND2_X1 U2929 ( .A1(n2308), .A2(REG2_REG_4__SCAN_IN), .ZN(n2283) );
  OAI21_X1 U2930 ( .B1(REG3_REG_3__SCAN_IN), .B2(REG3_REG_4__SCAN_IN), .A(
        n2290), .ZN(n4589) );
  OR2_X1 U2931 ( .A1(n2469), .A2(n4589), .ZN(n2282) );
  NAND2_X1 U2932 ( .A1(n2286), .A2(IR_REG_31__SCAN_IN), .ZN(n2287) );
  MUX2_X1 U2933 ( .A(n4222), .B(DATAI_4_), .S(n2939), .Z(n4372) );
  NAND2_X1 U2934 ( .A1(n3211), .A2(n4372), .ZN(n3709) );
  INV_X1 U2935 ( .A(n4372), .ZN(n4378) );
  NAND2_X1 U2936 ( .A1(n3838), .A2(n4378), .ZN(n3713) );
  NAND2_X1 U2937 ( .A1(n3709), .A2(n3713), .ZN(n4375) );
  NAND2_X1 U2938 ( .A1(n3838), .A2(n4372), .ZN(n2288) );
  NAND2_X1 U2939 ( .A1(n4370), .A2(n2288), .ZN(n3207) );
  NAND2_X1 U2940 ( .A1(n2478), .A2(REG2_REG_5__SCAN_IN), .ZN(n2295) );
  NAND2_X1 U2941 ( .A1(n2261), .A2(REG1_REG_5__SCAN_IN), .ZN(n2294) );
  AND2_X1 U2942 ( .A1(n2290), .A2(n2289), .ZN(n2291) );
  OR2_X1 U2943 ( .A1(n2291), .A2(n2309), .ZN(n3216) );
  OR2_X1 U2944 ( .A1(n2469), .A2(n3216), .ZN(n2293) );
  NAND2_X1 U2945 ( .A1(n3668), .A2(REG0_REG_5__SCAN_IN), .ZN(n2292) );
  INV_X1 U2946 ( .A(n2296), .ZN(n2298) );
  NAND2_X1 U2947 ( .A1(n2298), .A2(n2297), .ZN(n2300) );
  NAND2_X1 U2948 ( .A1(n2300), .A2(IR_REG_31__SCAN_IN), .ZN(n2299) );
  MUX2_X1 U2949 ( .A(n2299), .B(IR_REG_31__SCAN_IN), .S(n2301), .Z(n2303) );
  INV_X1 U2950 ( .A(n2300), .ZN(n2302) );
  NAND2_X1 U2951 ( .A1(n2302), .A2(n2301), .ZN(n2326) );
  NAND2_X1 U2952 ( .A1(n2303), .A2(n2326), .ZN(n3011) );
  INV_X1 U2953 ( .A(DATAI_5_), .ZN(n2304) );
  MUX2_X1 U2954 ( .A(n3011), .B(n2304), .S(n2939), .Z(n2645) );
  NAND2_X1 U2955 ( .A1(n2643), .A2(n2645), .ZN(n2305) );
  NAND2_X1 U2956 ( .A1(n3207), .A2(n2305), .ZN(n2307) );
  INV_X1 U2957 ( .A(n2643), .ZN(n3837) );
  NAND2_X1 U2958 ( .A1(n3837), .A2(n3215), .ZN(n2306) );
  NAND2_X1 U2959 ( .A1(n2307), .A2(n2306), .ZN(n3230) );
  NAND2_X1 U2960 ( .A1(n2261), .A2(REG1_REG_6__SCAN_IN), .ZN(n2313) );
  NAND2_X1 U2961 ( .A1(n2308), .A2(REG2_REG_6__SCAN_IN), .ZN(n2312) );
  OR2_X1 U2962 ( .A1(n2309), .A2(REG3_REG_6__SCAN_IN), .ZN(n2310) );
  NAND2_X1 U2963 ( .A1(n2320), .A2(n2310), .ZN(n3241) );
  OR2_X1 U2964 ( .A1(n2469), .A2(n3241), .ZN(n2311) );
  NAND2_X1 U2965 ( .A1(n3668), .A2(REG0_REG_6__SCAN_IN), .ZN(n2314) );
  NAND2_X1 U2966 ( .A1(n2326), .A2(IR_REG_31__SCAN_IN), .ZN(n2316) );
  XNOR2_X1 U2967 ( .A(n2316), .B(IR_REG_6__SCAN_IN), .ZN(n4209) );
  MUX2_X1 U2968 ( .A(n4209), .B(DATAI_6_), .S(n2939), .Z(n3232) );
  AND2_X1 U2969 ( .A1(n3836), .A2(n3232), .ZN(n2317) );
  INV_X1 U2970 ( .A(n3836), .ZN(n3178) );
  NAND2_X1 U2971 ( .A1(n3178), .A2(n3238), .ZN(n2318) );
  NAND2_X1 U2972 ( .A1(n3667), .A2(REG1_REG_7__SCAN_IN), .ZN(n2325) );
  NAND2_X1 U2973 ( .A1(n3668), .A2(REG0_REG_7__SCAN_IN), .ZN(n2324) );
  NAND2_X1 U2974 ( .A1(n2478), .A2(REG2_REG_7__SCAN_IN), .ZN(n2323) );
  NAND2_X1 U2975 ( .A1(n2320), .A2(n2319), .ZN(n2321) );
  NAND2_X1 U2976 ( .A1(n2343), .A2(n2321), .ZN(n3326) );
  OR2_X1 U2977 ( .A1(n2469), .A2(n3326), .ZN(n2322) );
  NAND2_X1 U2978 ( .A1(n2327), .A2(IR_REG_31__SCAN_IN), .ZN(n2335) );
  MUX2_X1 U2979 ( .A(n4208), .B(DATAI_7_), .S(n2939), .Z(n3180) );
  NAND2_X1 U2980 ( .A1(n3286), .A2(n3180), .ZN(n2525) );
  NAND2_X1 U2981 ( .A1(n3835), .A2(n3318), .ZN(n3725) );
  NAND2_X1 U2982 ( .A1(n3835), .A2(n3180), .ZN(n2329) );
  NAND2_X1 U2983 ( .A1(n3667), .A2(REG1_REG_8__SCAN_IN), .ZN(n2333) );
  NAND2_X1 U2984 ( .A1(n3668), .A2(REG0_REG_8__SCAN_IN), .ZN(n2332) );
  NAND2_X1 U2985 ( .A1(n2478), .A2(REG2_REG_8__SCAN_IN), .ZN(n2331) );
  INV_X1 U2986 ( .A(REG3_REG_8__SCAN_IN), .ZN(n2342) );
  XNOR2_X1 U2987 ( .A(n2343), .B(n2342), .ZN(n3289) );
  OR2_X1 U2988 ( .A1(n2469), .A2(n3289), .ZN(n2330) );
  INV_X1 U2989 ( .A(IR_REG_7__SCAN_IN), .ZN(n2334) );
  NAND2_X1 U2990 ( .A1(n2335), .A2(n2334), .ZN(n2336) );
  NAND2_X1 U2991 ( .A1(n2336), .A2(IR_REG_31__SCAN_IN), .ZN(n2338) );
  INV_X1 U2992 ( .A(DATAI_8_), .ZN(n2920) );
  MUX2_X1 U2993 ( .A(n3192), .B(n2920), .S(n2939), .Z(n2663) );
  NAND2_X1 U2994 ( .A1(n3319), .A2(n2663), .ZN(n2340) );
  AND2_X1 U2995 ( .A1(n3834), .A2(n3288), .ZN(n2339) );
  INV_X1 U2996 ( .A(REG3_REG_9__SCAN_IN), .ZN(n2341) );
  OAI21_X1 U2997 ( .B1(n2343), .B2(n2342), .A(n2341), .ZN(n2344) );
  NAND2_X1 U2998 ( .A1(n2344), .A2(n2354), .ZN(n3307) );
  OR2_X1 U2999 ( .A1(n2469), .A2(n3307), .ZN(n2348) );
  NAND2_X1 U3000 ( .A1(n3667), .A2(REG1_REG_9__SCAN_IN), .ZN(n2347) );
  NAND2_X1 U3001 ( .A1(n3668), .A2(REG0_REG_9__SCAN_IN), .ZN(n2346) );
  NAND2_X1 U3002 ( .A1(n2478), .A2(REG2_REG_9__SCAN_IN), .ZN(n2345) );
  OR2_X1 U3003 ( .A1(n2349), .A2(n2559), .ZN(n2350) );
  XNOR2_X1 U3004 ( .A(n2350), .B(IR_REG_9__SCAN_IN), .ZN(n3196) );
  MUX2_X1 U3005 ( .A(n3196), .B(DATAI_9_), .S(n2939), .Z(n3312) );
  NAND2_X1 U3006 ( .A1(n3833), .A2(n3312), .ZN(n2351) );
  NAND2_X1 U3007 ( .A1(n3305), .A2(n2351), .ZN(n2353) );
  INV_X1 U3008 ( .A(n3312), .ZN(n2528) );
  NAND2_X1 U3009 ( .A1(n3345), .A2(n2528), .ZN(n2352) );
  INV_X1 U3010 ( .A(n2365), .ZN(n2356) );
  NAND2_X1 U3011 ( .A1(n2354), .A2(n3251), .ZN(n2355) );
  NAND2_X1 U3012 ( .A1(n2356), .A2(n2355), .ZN(n3250) );
  OR2_X1 U3013 ( .A1(n2469), .A2(n3250), .ZN(n2360) );
  NAND2_X1 U3014 ( .A1(n3667), .A2(REG1_REG_10__SCAN_IN), .ZN(n2359) );
  NAND2_X1 U3015 ( .A1(n3668), .A2(REG0_REG_10__SCAN_IN), .ZN(n2358) );
  NAND2_X1 U3016 ( .A1(n2478), .A2(REG2_REG_10__SCAN_IN), .ZN(n2357) );
  NOR2_X1 U3017 ( .A1(n2436), .A2(n2559), .ZN(n2361) );
  MUX2_X1 U3018 ( .A(n2559), .B(n2361), .S(IR_REG_10__SCAN_IN), .Z(n2364) );
  NAND2_X1 U3019 ( .A1(n2436), .A2(n2362), .ZN(n2394) );
  INV_X1 U3020 ( .A(n2394), .ZN(n2363) );
  MUX2_X1 U3021 ( .A(n4354), .B(DATAI_10_), .S(n2939), .Z(n3342) );
  NOR2_X1 U3022 ( .A1(n3832), .A2(n3342), .ZN(n3363) );
  NAND2_X1 U3023 ( .A1(n3667), .A2(REG1_REG_11__SCAN_IN), .ZN(n2370) );
  NAND2_X1 U3024 ( .A1(n3668), .A2(REG0_REG_11__SCAN_IN), .ZN(n2369) );
  NAND2_X1 U3025 ( .A1(n2478), .A2(REG2_REG_11__SCAN_IN), .ZN(n2368) );
  OR2_X1 U3026 ( .A1(n2365), .A2(REG3_REG_11__SCAN_IN), .ZN(n2366) );
  NAND2_X1 U3027 ( .A1(n2388), .A2(n2366), .ZN(n3376) );
  OR2_X1 U3028 ( .A1(n2469), .A2(n3376), .ZN(n2367) );
  NAND2_X1 U3029 ( .A1(n2394), .A2(IR_REG_31__SCAN_IN), .ZN(n2372) );
  INV_X1 U3030 ( .A(IR_REG_11__SCAN_IN), .ZN(n2371) );
  NAND2_X1 U3031 ( .A1(n2372), .A2(n2371), .ZN(n2381) );
  OR2_X1 U3032 ( .A1(n2372), .A2(n2371), .ZN(n2373) );
  MUX2_X1 U3033 ( .A(n4207), .B(DATAI_11_), .S(n2939), .Z(n3271) );
  AND2_X1 U3034 ( .A1(n2679), .A2(n3374), .ZN(n2375) );
  NAND2_X1 U3035 ( .A1(n2679), .A2(n3271), .ZN(n3381) );
  INV_X1 U3036 ( .A(n2679), .ZN(n3831) );
  NAND2_X1 U3037 ( .A1(n3831), .A2(n3374), .ZN(n3383) );
  INV_X1 U3038 ( .A(n3791), .ZN(n2374) );
  NAND2_X1 U3039 ( .A1(n3832), .A2(n3342), .ZN(n3364) );
  NOR2_X1 U3040 ( .A1(n2375), .A2(n3365), .ZN(n2376) );
  NAND2_X1 U3041 ( .A1(n3667), .A2(REG1_REG_12__SCAN_IN), .ZN(n2380) );
  NAND2_X1 U3042 ( .A1(n3668), .A2(REG0_REG_12__SCAN_IN), .ZN(n2379) );
  NAND2_X1 U3043 ( .A1(n2478), .A2(REG2_REG_12__SCAN_IN), .ZN(n2378) );
  INV_X1 U3044 ( .A(REG3_REG_12__SCAN_IN), .ZN(n2387) );
  XNOR2_X1 U3045 ( .A(n2388), .B(n2387), .ZN(n3393) );
  OR2_X1 U3046 ( .A1(n2794), .A2(n3393), .ZN(n2377) );
  NAND2_X1 U3047 ( .A1(n2381), .A2(IR_REG_31__SCAN_IN), .ZN(n2382) );
  XNOR2_X1 U3048 ( .A(n2382), .B(IR_REG_12__SCAN_IN), .ZN(n3885) );
  INV_X1 U3049 ( .A(DATAI_12_), .ZN(n2383) );
  MUX2_X1 U3050 ( .A(n4353), .B(n2383), .S(n2939), .Z(n3391) );
  NAND2_X1 U3051 ( .A1(n2385), .A2(n2384), .ZN(n3405) );
  NAND2_X1 U3052 ( .A1(n3667), .A2(REG1_REG_13__SCAN_IN), .ZN(n2393) );
  NAND2_X1 U3053 ( .A1(n3668), .A2(REG0_REG_13__SCAN_IN), .ZN(n2392) );
  NAND2_X1 U3054 ( .A1(n2478), .A2(REG2_REG_13__SCAN_IN), .ZN(n2391) );
  INV_X1 U3055 ( .A(REG3_REG_13__SCAN_IN), .ZN(n2386) );
  OAI21_X1 U3056 ( .B1(n2388), .B2(n2387), .A(n2386), .ZN(n2389) );
  NAND2_X1 U3057 ( .A1(n2389), .A2(n2400), .ZN(n3334) );
  OR2_X1 U3058 ( .A1(n2794), .A2(n3334), .ZN(n2390) );
  NAND2_X1 U3059 ( .A1(n2396), .A2(IR_REG_31__SCAN_IN), .ZN(n2395) );
  MUX2_X1 U3060 ( .A(IR_REG_31__SCAN_IN), .B(n2395), .S(IR_REG_13__SCAN_IN), 
        .Z(n2398) );
  INV_X1 U3061 ( .A(n2414), .ZN(n2397) );
  NAND2_X1 U3062 ( .A1(n2398), .A2(n2397), .ZN(n4272) );
  INV_X1 U3063 ( .A(DATAI_13_), .ZN(n2399) );
  MUX2_X1 U3064 ( .A(n4272), .B(n2399), .S(n2939), .Z(n3420) );
  NAND2_X1 U3065 ( .A1(n3667), .A2(REG1_REG_14__SCAN_IN), .ZN(n2406) );
  NAND2_X1 U3066 ( .A1(n3668), .A2(REG0_REG_14__SCAN_IN), .ZN(n2405) );
  NAND2_X1 U3067 ( .A1(n2478), .A2(REG2_REG_14__SCAN_IN), .ZN(n2404) );
  INV_X1 U3068 ( .A(n2418), .ZN(n2402) );
  NAND2_X1 U3069 ( .A1(n2400), .A2(n4485), .ZN(n2401) );
  NAND2_X1 U3070 ( .A1(n2402), .A2(n2401), .ZN(n3439) );
  OR2_X1 U3071 ( .A1(n2794), .A2(n3439), .ZN(n2403) );
  OR2_X1 U3072 ( .A1(n2414), .A2(n2559), .ZN(n2407) );
  XNOR2_X1 U3073 ( .A(n2407), .B(IR_REG_14__SCAN_IN), .ZN(n4280) );
  MUX2_X1 U3074 ( .A(n4280), .B(DATAI_14_), .S(n2939), .Z(n3430) );
  NAND2_X1 U3075 ( .A1(n3462), .A2(n3430), .ZN(n3652) );
  NAND2_X1 U3076 ( .A1(n3828), .A2(n2408), .ZN(n3653) );
  NAND2_X1 U3077 ( .A1(n3652), .A2(n3653), .ZN(n3429) );
  NAND2_X1 U3078 ( .A1(n3667), .A2(REG1_REG_15__SCAN_IN), .ZN(n2412) );
  NAND2_X1 U3079 ( .A1(n3668), .A2(REG0_REG_15__SCAN_IN), .ZN(n2411) );
  NAND2_X1 U3080 ( .A1(n2478), .A2(REG2_REG_15__SCAN_IN), .ZN(n2410) );
  XNOR2_X1 U3081 ( .A(n2418), .B(REG3_REG_15__SCAN_IN), .ZN(n3643) );
  OR2_X1 U3082 ( .A1(n2469), .A2(n3643), .ZN(n2409) );
  INV_X1 U3083 ( .A(IR_REG_14__SCAN_IN), .ZN(n2413) );
  NAND2_X1 U3084 ( .A1(n2414), .A2(n2413), .ZN(n2415) );
  NAND2_X1 U3085 ( .A1(n2415), .A2(IR_REG_31__SCAN_IN), .ZN(n2425) );
  XNOR2_X1 U3086 ( .A(n2425), .B(IR_REG_15__SCAN_IN), .ZN(n4347) );
  MUX2_X1 U3087 ( .A(n4347), .B(DATAI_15_), .S(n2939), .Z(n3648) );
  NAND2_X1 U3088 ( .A1(n3827), .A2(n3648), .ZN(n2417) );
  NAND2_X1 U3089 ( .A1(n3667), .A2(REG1_REG_16__SCAN_IN), .ZN(n2423) );
  NAND2_X1 U3090 ( .A1(n3668), .A2(REG0_REG_16__SCAN_IN), .ZN(n2422) );
  NAND2_X1 U3091 ( .A1(n2478), .A2(REG2_REG_16__SCAN_IN), .ZN(n2421) );
  AOI21_X1 U3092 ( .B1(n2418), .B2(REG3_REG_15__SCAN_IN), .A(
        REG3_REG_16__SCAN_IN), .ZN(n2419) );
  OR2_X1 U3093 ( .A1(n2429), .A2(n2419), .ZN(n3576) );
  OR2_X1 U3094 ( .A1(n2794), .A2(n3576), .ZN(n2420) );
  INV_X1 U3095 ( .A(IR_REG_15__SCAN_IN), .ZN(n2424) );
  NAND2_X1 U3096 ( .A1(n2425), .A2(n2424), .ZN(n2426) );
  NAND2_X1 U3097 ( .A1(n2426), .A2(IR_REG_31__SCAN_IN), .ZN(n2428) );
  INV_X1 U3098 ( .A(IR_REG_16__SCAN_IN), .ZN(n2427) );
  XNOR2_X1 U3099 ( .A(n2428), .B(n2427), .ZN(n4346) );
  MUX2_X1 U3100 ( .A(n3875), .B(DATAI_16_), .S(n2939), .Z(n3579) );
  NAND2_X1 U3101 ( .A1(n4094), .A2(n3579), .ZN(n3748) );
  INV_X1 U3102 ( .A(n4094), .ZN(n3826) );
  NAND2_X1 U3103 ( .A1(n3826), .A2(n2701), .ZN(n3745) );
  NAND2_X1 U3104 ( .A1(n3748), .A2(n3745), .ZN(n3472) );
  NAND2_X1 U3105 ( .A1(n3471), .A2(n3472), .ZN(n3470) );
  NAND2_X1 U3106 ( .A1(n3470), .A2(n2190), .ZN(n4083) );
  NAND2_X1 U3107 ( .A1(n3667), .A2(REG1_REG_17__SCAN_IN), .ZN(n2435) );
  NAND2_X1 U3108 ( .A1(n3668), .A2(REG0_REG_17__SCAN_IN), .ZN(n2434) );
  NAND2_X1 U3109 ( .A1(n2478), .A2(REG2_REG_17__SCAN_IN), .ZN(n2433) );
  OR2_X1 U3110 ( .A1(n2429), .A2(REG3_REG_17__SCAN_IN), .ZN(n2430) );
  NAND2_X1 U3111 ( .A1(n2431), .A2(n2430), .ZN(n3586) );
  OR2_X1 U3112 ( .A1(n2794), .A2(n3586), .ZN(n2432) );
  NAND2_X1 U3113 ( .A1(n2436), .A2(n2215), .ZN(n2437) );
  NAND2_X1 U3114 ( .A1(n2437), .A2(IR_REG_31__SCAN_IN), .ZN(n2438) );
  XNOR2_X1 U3115 ( .A(n2438), .B(IR_REG_17__SCAN_IN), .ZN(n3892) );
  MUX2_X1 U3116 ( .A(n3892), .B(DATAI_17_), .S(n2939), .Z(n4088) );
  NAND2_X1 U3117 ( .A1(n4075), .A2(n4096), .ZN(n2439) );
  INV_X1 U3118 ( .A(n4090), .ZN(n4055) );
  NAND2_X1 U3119 ( .A1(n4055), .A2(n4072), .ZN(n4044) );
  NAND2_X1 U3120 ( .A1(n4090), .A2(n4069), .ZN(n4045) );
  NAND2_X1 U3121 ( .A1(n4044), .A2(n4045), .ZN(n4071) );
  INV_X1 U3122 ( .A(REG3_REG_19__SCAN_IN), .ZN(n2440) );
  AND2_X1 U3123 ( .A1(n2441), .A2(n2440), .ZN(n2442) );
  NOR2_X1 U3124 ( .A1(n2452), .A2(n2442), .ZN(n4058) );
  NAND2_X1 U3125 ( .A1(n2823), .A2(n4058), .ZN(n2446) );
  NAND2_X1 U3126 ( .A1(n3667), .A2(REG1_REG_19__SCAN_IN), .ZN(n2445) );
  NAND2_X1 U3127 ( .A1(n3668), .A2(REG0_REG_19__SCAN_IN), .ZN(n2444) );
  NAND2_X1 U3128 ( .A1(n2478), .A2(REG2_REG_19__SCAN_IN), .ZN(n2443) );
  NAND4_X1 U3129 ( .A1(n2446), .A2(n2445), .A3(n2444), .A4(n2443), .ZN(n4073)
         );
  NAND2_X1 U3130 ( .A1(n2449), .A2(n2448), .ZN(n2501) );
  INV_X1 U3131 ( .A(DATAI_19_), .ZN(n2450) );
  MUX2_X1 U3132 ( .A(n3898), .B(n2450), .S(n2939), .Z(n4057) );
  NAND2_X1 U3133 ( .A1(n4073), .A2(n3543), .ZN(n2451) );
  NOR2_X1 U3134 ( .A1(n2452), .A2(REG3_REG_20__SCAN_IN), .ZN(n2453) );
  OR2_X1 U3135 ( .A1(n2459), .A2(n2453), .ZN(n4037) );
  OR2_X1 U3136 ( .A1(n2794), .A2(n4037), .ZN(n2457) );
  NAND2_X1 U3137 ( .A1(n3667), .A2(REG1_REG_20__SCAN_IN), .ZN(n2456) );
  NAND2_X1 U3138 ( .A1(n3668), .A2(REG0_REG_20__SCAN_IN), .ZN(n2455) );
  NAND2_X1 U3139 ( .A1(n2478), .A2(REG2_REG_20__SCAN_IN), .ZN(n2454) );
  NAND4_X1 U3140 ( .A1(n2457), .A2(n2456), .A3(n2455), .A4(n2454), .ZN(n4052)
         );
  INV_X1 U3141 ( .A(n4052), .ZN(n3552) );
  NAND2_X1 U3142 ( .A1(n2939), .A2(DATAI_20_), .ZN(n4035) );
  NAND2_X1 U3143 ( .A1(n3552), .A2(n4035), .ZN(n2458) );
  NAND2_X1 U3144 ( .A1(n2261), .A2(REG1_REG_21__SCAN_IN), .ZN(n2464) );
  NAND2_X1 U3145 ( .A1(n3668), .A2(REG0_REG_21__SCAN_IN), .ZN(n2463) );
  NAND2_X1 U3146 ( .A1(n2478), .A2(REG2_REG_21__SCAN_IN), .ZN(n2462) );
  OR2_X1 U3147 ( .A1(n2459), .A2(REG3_REG_21__SCAN_IN), .ZN(n2460) );
  NAND2_X1 U31480 ( .A1(n2467), .A2(n2460), .ZN(n4012) );
  OR2_X1 U31490 ( .A1(n2469), .A2(n4012), .ZN(n2461) );
  INV_X1 U3150 ( .A(n4029), .ZN(n3824) );
  AND2_X1 U3151 ( .A1(n2939), .A2(DATAI_21_), .ZN(n4004) );
  NAND2_X1 U3152 ( .A1(n3824), .A2(n4004), .ZN(n2465) );
  AOI21_X1 U3153 ( .B1(n4001), .B2(n2465), .A(n2189), .ZN(n3986) );
  NAND2_X1 U3154 ( .A1(n3668), .A2(REG0_REG_22__SCAN_IN), .ZN(n2473) );
  NAND2_X1 U3155 ( .A1(n2478), .A2(REG2_REG_22__SCAN_IN), .ZN(n2472) );
  NAND2_X1 U3156 ( .A1(n3667), .A2(REG1_REG_22__SCAN_IN), .ZN(n2471) );
  INV_X1 U3157 ( .A(REG3_REG_22__SCAN_IN), .ZN(n2466) );
  NAND2_X1 U3158 ( .A1(n2467), .A2(n2466), .ZN(n2468) );
  NAND2_X1 U3159 ( .A1(n2476), .A2(n2468), .ZN(n3994) );
  OR2_X1 U3160 ( .A1(n2469), .A2(n3994), .ZN(n2470) );
  AND2_X1 U3161 ( .A1(n2939), .A2(DATAI_22_), .ZN(n3996) );
  NAND2_X1 U3162 ( .A1(n4007), .A2(n3996), .ZN(n2545) );
  INV_X1 U3163 ( .A(n3996), .ZN(n2739) );
  NAND2_X1 U3164 ( .A1(n3823), .A2(n2739), .ZN(n2547) );
  NAND2_X1 U3165 ( .A1(n2545), .A2(n2547), .ZN(n3985) );
  NAND2_X1 U3166 ( .A1(n3986), .A2(n3985), .ZN(n3984) );
  NAND2_X1 U3167 ( .A1(n3823), .A2(n3996), .ZN(n2474) );
  NAND2_X1 U3168 ( .A1(n3984), .A2(n2474), .ZN(n3961) );
  INV_X1 U3169 ( .A(REG3_REG_23__SCAN_IN), .ZN(n2475) );
  AND2_X1 U3170 ( .A1(n2476), .A2(n2475), .ZN(n2477) );
  NOR2_X1 U3171 ( .A1(n2485), .A2(n2477), .ZN(n3979) );
  NAND2_X1 U3172 ( .A1(n2823), .A2(n3979), .ZN(n2482) );
  NAND2_X1 U3173 ( .A1(n3667), .A2(REG1_REG_23__SCAN_IN), .ZN(n2481) );
  NAND2_X1 U3174 ( .A1(n3668), .A2(REG0_REG_23__SCAN_IN), .ZN(n2480) );
  NAND2_X1 U3175 ( .A1(n2478), .A2(REG2_REG_23__SCAN_IN), .ZN(n2479) );
  NAND4_X1 U3176 ( .A1(n2482), .A2(n2481), .A3(n2480), .A4(n2479), .ZN(n3989)
         );
  INV_X1 U3177 ( .A(n3989), .ZN(n3952) );
  NAND2_X1 U3178 ( .A1(n2939), .A2(DATAI_23_), .ZN(n3978) );
  NAND2_X1 U3179 ( .A1(n3952), .A2(n3978), .ZN(n2484) );
  NOR2_X1 U3180 ( .A1(n3952), .A2(n3978), .ZN(n2483) );
  NAND2_X1 U3181 ( .A1(n3667), .A2(REG1_REG_24__SCAN_IN), .ZN(n2490) );
  NOR2_X1 U3182 ( .A1(n2485), .A2(REG3_REG_24__SCAN_IN), .ZN(n2486) );
  OR2_X1 U3183 ( .A1(n2492), .A2(n2486), .ZN(n3597) );
  OR2_X1 U3184 ( .A1(n3597), .A2(n2794), .ZN(n2489) );
  NAND2_X1 U3185 ( .A1(n3668), .A2(REG0_REG_24__SCAN_IN), .ZN(n2488) );
  NAND2_X1 U3186 ( .A1(n2478), .A2(REG2_REG_24__SCAN_IN), .ZN(n2487) );
  AND2_X1 U3187 ( .A1(n2939), .A2(DATAI_24_), .ZN(n3948) );
  NAND2_X1 U3188 ( .A1(n3972), .A2(n3948), .ZN(n2839) );
  NAND2_X1 U3189 ( .A1(n2842), .A2(n2839), .ZN(n2491) );
  NAND2_X1 U3190 ( .A1(n3565), .A2(n3955), .ZN(n2845) );
  OR2_X1 U3191 ( .A1(n2492), .A2(REG3_REG_25__SCAN_IN), .ZN(n2493) );
  NAND2_X1 U3192 ( .A1(n2782), .A2(n2493), .ZN(n3561) );
  NAND2_X1 U3193 ( .A1(n3667), .A2(REG1_REG_25__SCAN_IN), .ZN(n2495) );
  NAND2_X1 U3194 ( .A1(n3668), .A2(REG0_REG_25__SCAN_IN), .ZN(n2494) );
  AND2_X1 U3195 ( .A1(n2495), .A2(n2494), .ZN(n2497) );
  NAND2_X1 U3196 ( .A1(n2478), .A2(REG2_REG_25__SCAN_IN), .ZN(n2496) );
  INV_X1 U3197 ( .A(n3949), .ZN(n2498) );
  NAND2_X1 U3198 ( .A1(n2939), .A2(DATAI_25_), .ZN(n2765) );
  INV_X1 U3199 ( .A(n2765), .ZN(n3562) );
  NAND2_X1 U3200 ( .A1(n2498), .A2(n3562), .ZN(n2875) );
  NAND2_X1 U3201 ( .A1(n3949), .A2(n2765), .ZN(n2855) );
  NAND2_X1 U3202 ( .A1(n2875), .A2(n2855), .ZN(n3785) );
  NAND2_X1 U3203 ( .A1(n2032), .A2(IR_REG_31__SCAN_IN), .ZN(n2500) );
  XNOR2_X1 U3204 ( .A(n2500), .B(IR_REG_22__SCAN_IN), .ZN(n4205) );
  INV_X1 U3205 ( .A(n2504), .ZN(n2505) );
  NAND2_X1 U3206 ( .A1(n2505), .A2(IR_REG_31__SCAN_IN), .ZN(n2506) );
  XNOR2_X1 U3207 ( .A(n4205), .B(n2603), .ZN(n2507) );
  NAND2_X1 U3208 ( .A1(n2507), .A2(n3898), .ZN(n4380) );
  INV_X1 U3209 ( .A(n4205), .ZN(n2555) );
  NAND3_X1 U32100 ( .A1(n2555), .A2(n4592), .A3(n2508), .ZN(n4414) );
  XNOR2_X1 U32110 ( .A(n2782), .B(REG3_REG_26__SCAN_IN), .ZN(n3929) );
  NAND2_X1 U32120 ( .A1(n3929), .A2(n2823), .ZN(n2513) );
  NAND2_X1 U32130 ( .A1(n2478), .A2(REG2_REG_26__SCAN_IN), .ZN(n2511) );
  NAND2_X1 U32140 ( .A1(n3667), .A2(REG1_REG_26__SCAN_IN), .ZN(n2510) );
  NAND2_X1 U32150 ( .A1(n3668), .A2(REG0_REG_26__SCAN_IN), .ZN(n2509) );
  INV_X1 U32160 ( .A(n3822), .ZN(n2849) );
  NOR2_X1 U32170 ( .A1(n2514), .A2(n2559), .ZN(n2515) );
  MUX2_X1 U32180 ( .A(n2559), .B(n2515), .S(IR_REG_28__SCAN_IN), .Z(n2516) );
  INV_X1 U32190 ( .A(n2516), .ZN(n2518) );
  NAND2_X1 U32200 ( .A1(n2518), .A2(n2517), .ZN(n2956) );
  NAND2_X1 U32210 ( .A1(n4205), .A2(n3808), .ZN(n2811) );
  INV_X1 U32220 ( .A(n2811), .ZN(n2936) );
  NAND2_X1 U32230 ( .A1(n2956), .A2(n2936), .ZN(n4379) );
  INV_X1 U32240 ( .A(n2519), .ZN(n3774) );
  NOR2_X1 U32250 ( .A1(n3841), .A2(n2585), .ZN(n3701) );
  NAND2_X1 U32260 ( .A1(n3774), .A2(n3701), .ZN(n3070) );
  NAND2_X1 U32270 ( .A1(n3070), .A2(n3702), .ZN(n2521) );
  NAND2_X1 U32280 ( .A1(n2521), .A2(n3792), .ZN(n3072) );
  NAND2_X1 U32290 ( .A1(n3072), .A2(n3703), .ZN(n3090) );
  INV_X1 U32300 ( .A(n4383), .ZN(n3126) );
  NAND2_X1 U32310 ( .A1(n3126), .A2(n3134), .ZN(n3708) );
  NAND2_X1 U32320 ( .A1(n4383), .A2(n3095), .ZN(n3705) );
  AND2_X2 U32330 ( .A1(n3708), .A2(n3705), .ZN(n3789) );
  NAND2_X1 U32340 ( .A1(n3090), .A2(n3789), .ZN(n3089) );
  NAND2_X1 U32350 ( .A1(n3089), .A2(n3708), .ZN(n4376) );
  INV_X1 U32360 ( .A(n3709), .ZN(n2522) );
  OR2_X1 U32370 ( .A1(n4376), .A2(n2522), .ZN(n2523) );
  NAND2_X1 U32380 ( .A1(n2523), .A2(n3713), .ZN(n3209) );
  AND2_X1 U32390 ( .A1(n3837), .A2(n2645), .ZN(n3208) );
  NAND2_X1 U32400 ( .A1(n2643), .A2(n3215), .ZN(n3726) );
  NAND2_X1 U32410 ( .A1(n3836), .A2(n3238), .ZN(n3712) );
  NOR2_X1 U32420 ( .A1(n3836), .A2(n3238), .ZN(n3715) );
  AOI21_X1 U32430 ( .B1(n3231), .B2(n3712), .A(n3715), .ZN(n3320) );
  NAND2_X1 U32440 ( .A1(n3320), .A2(n2525), .ZN(n2526) );
  NAND2_X1 U32450 ( .A1(n2526), .A2(n3725), .ZN(n3281) );
  NAND2_X1 U32460 ( .A1(n3319), .A2(n3288), .ZN(n3719) );
  NAND2_X1 U32470 ( .A1(n3281), .A2(n3719), .ZN(n2527) );
  NAND2_X1 U32480 ( .A1(n3834), .A2(n2663), .ZN(n3729) );
  NAND2_X1 U32490 ( .A1(n2527), .A2(n3729), .ZN(n3310) );
  AND2_X1 U32500 ( .A1(n3833), .A2(n2528), .ZN(n3723) );
  OR2_X2 U32510 ( .A1(n3310), .A2(n3723), .ZN(n2529) );
  NAND2_X1 U32520 ( .A1(n3345), .A2(n3312), .ZN(n3720) );
  NAND2_X1 U32530 ( .A1(n3832), .A2(n2133), .ZN(n3735) );
  NAND2_X1 U32540 ( .A1(n3340), .A2(n3735), .ZN(n2530) );
  INV_X1 U32550 ( .A(n3832), .ZN(n3275) );
  NAND2_X1 U32560 ( .A1(n3275), .A2(n3342), .ZN(n3733) );
  NAND2_X1 U32570 ( .A1(n3830), .A2(n3391), .ZN(n3406) );
  NAND2_X1 U32580 ( .A1(n3829), .A2(n3420), .ZN(n2531) );
  NAND2_X1 U32590 ( .A1(n3406), .A2(n2531), .ZN(n2533) );
  INV_X1 U32600 ( .A(n3383), .ZN(n2532) );
  NOR2_X1 U32610 ( .A1(n2533), .A2(n2532), .ZN(n3736) );
  NAND2_X1 U32620 ( .A1(n3370), .A2(n3736), .ZN(n2537) );
  NAND2_X1 U32630 ( .A1(n3413), .A2(n3385), .ZN(n3408) );
  NAND2_X1 U32640 ( .A1(n3381), .A2(n3408), .ZN(n2536) );
  INV_X1 U32650 ( .A(n2533), .ZN(n2535) );
  NOR2_X1 U32660 ( .A1(n3829), .A2(n3420), .ZN(n2534) );
  AOI21_X1 U32670 ( .B1(n2536), .B2(n2535), .A(n2534), .ZN(n3739) );
  NAND2_X1 U32680 ( .A1(n2537), .A2(n3739), .ZN(n3656) );
  INV_X1 U32690 ( .A(n3429), .ZN(n3772) );
  NAND2_X1 U32700 ( .A1(n3656), .A2(n3772), .ZN(n3456) );
  NAND2_X1 U32710 ( .A1(n3575), .A2(n3648), .ZN(n3655) );
  NAND2_X1 U32720 ( .A1(n3827), .A2(n3464), .ZN(n3654) );
  NAND2_X1 U32730 ( .A1(n3655), .A2(n3654), .ZN(n3457) );
  INV_X1 U32740 ( .A(n3652), .ZN(n2538) );
  NOR2_X1 U32750 ( .A1(n3457), .A2(n2538), .ZN(n2539) );
  NAND2_X1 U32760 ( .A1(n3456), .A2(n2539), .ZN(n2540) );
  NAND2_X1 U32770 ( .A1(n2540), .A2(n3654), .ZN(n3473) );
  INV_X1 U32780 ( .A(n3472), .ZN(n3771) );
  NAND2_X1 U32790 ( .A1(n3473), .A2(n3771), .ZN(n2541) );
  NAND2_X1 U32800 ( .A1(n4073), .A2(n4057), .ZN(n3781) );
  NAND2_X1 U32810 ( .A1(n3781), .A2(n4045), .ZN(n2542) );
  INV_X1 U32820 ( .A(n2542), .ZN(n4025) );
  NAND2_X1 U32830 ( .A1(n3825), .A2(n4096), .ZN(n4021) );
  NAND2_X1 U32840 ( .A1(n4025), .A2(n4021), .ZN(n3747) );
  INV_X1 U32850 ( .A(n4073), .ZN(n4033) );
  NAND2_X1 U32860 ( .A1(n4033), .A2(n3543), .ZN(n3782) );
  OAI21_X1 U32870 ( .B1(n2542), .B2(n4044), .A(n3782), .ZN(n4024) );
  NAND2_X1 U32880 ( .A1(n4075), .A2(n4088), .ZN(n4022) );
  OAI22_X1 U32890 ( .A1(n2542), .A2(n4022), .B1(n4035), .B2(n4052), .ZN(n2543)
         );
  OR2_X1 U32900 ( .A1(n4024), .A2(n2543), .ZN(n3751) );
  INV_X1 U32910 ( .A(n3751), .ZN(n3660) );
  OAI21_X1 U32920 ( .B1(n4020), .B2(n3747), .A(n3660), .ZN(n2544) );
  NAND2_X1 U32930 ( .A1(n4052), .A2(n4035), .ZN(n3750) );
  NAND2_X1 U32940 ( .A1(n2544), .A2(n3750), .ZN(n4003) );
  NAND2_X1 U32950 ( .A1(n4029), .A2(n4004), .ZN(n3965) );
  NAND2_X1 U32960 ( .A1(n2545), .A2(n3965), .ZN(n3664) );
  INV_X1 U32970 ( .A(n3664), .ZN(n3755) );
  NAND2_X1 U32980 ( .A1(n4003), .A2(n3755), .ZN(n2550) );
  NAND2_X1 U32990 ( .A1(n3824), .A2(n4010), .ZN(n3963) );
  INV_X1 U33000 ( .A(n2545), .ZN(n3967) );
  OR2_X1 U33010 ( .A1(n3963), .A2(n3967), .ZN(n2549) );
  NAND2_X1 U33020 ( .A1(n3989), .A2(n3978), .ZN(n2546) );
  NAND2_X1 U33030 ( .A1(n2547), .A2(n2546), .ZN(n3753) );
  INV_X1 U33040 ( .A(n3753), .ZN(n2548) );
  AND2_X1 U33050 ( .A1(n2549), .A2(n2548), .ZN(n3662) );
  NAND2_X1 U33060 ( .A1(n2550), .A2(n3662), .ZN(n3944) );
  OR2_X1 U33070 ( .A1(n3989), .A2(n3978), .ZN(n3943) );
  NAND2_X1 U33080 ( .A1(n3565), .A2(n3948), .ZN(n3779) );
  NAND2_X1 U33090 ( .A1(n3944), .A2(n3756), .ZN(n2856) );
  NAND2_X1 U33100 ( .A1(n3972), .A2(n3955), .ZN(n3780) );
  NAND2_X1 U33110 ( .A1(n2856), .A2(n3780), .ZN(n2551) );
  XNOR2_X1 U33120 ( .A(n2551), .B(n3785), .ZN(n2553) );
  NAND2_X1 U33130 ( .A1(n4205), .A2(n4592), .ZN(n2552) );
  INV_X1 U33140 ( .A(n2508), .ZN(n4206) );
  NAND2_X1 U33150 ( .A1(n4206), .A2(n3808), .ZN(n3691) );
  NAND2_X1 U33160 ( .A1(n2552), .A2(n3691), .ZN(n4086) );
  NAND2_X1 U33170 ( .A1(n2553), .A2(n4086), .ZN(n2558) );
  INV_X1 U33180 ( .A(n3808), .ZN(n2554) );
  AND2_X2 U33190 ( .A1(n3031), .A2(n4206), .ZN(n4112) );
  OAI22_X1 U33200 ( .A1(n3565), .A2(n4093), .B1(n2765), .B2(n4377), .ZN(n2556)
         );
  INV_X1 U33210 ( .A(n2556), .ZN(n2557) );
  OAI211_X1 U33220 ( .C1(n2849), .C2(n4379), .A(n2558), .B(n2557), .ZN(n3940)
         );
  AOI21_X1 U33230 ( .B1(n3936), .B2(n4400), .A(n3940), .ZN(n4126) );
  OR2_X1 U33240 ( .A1(n2560), .A2(n2559), .ZN(n2579) );
  INV_X1 U33250 ( .A(IR_REG_23__SCAN_IN), .ZN(n2578) );
  NAND2_X1 U33260 ( .A1(n2579), .A2(n2578), .ZN(n2577) );
  NAND2_X1 U33270 ( .A1(n2577), .A2(IR_REG_31__SCAN_IN), .ZN(n2561) );
  NAND2_X1 U33280 ( .A1(n2562), .A2(IR_REG_31__SCAN_IN), .ZN(n2563) );
  XNOR2_X1 U33290 ( .A(n2563), .B(IR_REG_25__SCAN_IN), .ZN(n4203) );
  INV_X1 U33300 ( .A(n4203), .ZN(n2932) );
  NAND2_X1 U33310 ( .A1(n2930), .A2(n2932), .ZN(n2564) );
  MUX2_X1 U33320 ( .A(n2930), .B(n2564), .S(B_REG_SCAN_IN), .Z(n2566) );
  NAND2_X1 U33330 ( .A1(n2566), .A2(n4202), .ZN(n2928) );
  OAI22_X1 U33340 ( .A1(n2928), .A2(D_REG_1__SCAN_IN), .B1(n4203), .B2(n4202), 
        .ZN(n2590) );
  OR2_X1 U33350 ( .A1(n4414), .A2(n3808), .ZN(n2829) );
  AND2_X1 U33360 ( .A1(n2590), .A2(n2829), .ZN(n2580) );
  INV_X1 U33370 ( .A(n2928), .ZN(n2583) );
  NOR4_X1 U33380 ( .A1(D_REG_16__SCAN_IN), .A2(D_REG_20__SCAN_IN), .A3(
        D_REG_30__SCAN_IN), .A4(D_REG_7__SCAN_IN), .ZN(n2575) );
  NOR4_X1 U33390 ( .A1(D_REG_11__SCAN_IN), .A2(D_REG_3__SCAN_IN), .A3(
        D_REG_4__SCAN_IN), .A4(D_REG_5__SCAN_IN), .ZN(n2574) );
  INV_X1 U33400 ( .A(D_REG_2__SCAN_IN), .ZN(n4526) );
  INV_X1 U33410 ( .A(D_REG_23__SCAN_IN), .ZN(n4532) );
  INV_X1 U33420 ( .A(D_REG_17__SCAN_IN), .ZN(n4531) );
  INV_X1 U33430 ( .A(D_REG_12__SCAN_IN), .ZN(n4535) );
  NAND4_X1 U33440 ( .A1(n4526), .A2(n4532), .A3(n4531), .A4(n4535), .ZN(n2572)
         );
  NOR4_X1 U33450 ( .A1(D_REG_13__SCAN_IN), .A2(D_REG_14__SCAN_IN), .A3(
        D_REG_15__SCAN_IN), .A4(D_REG_18__SCAN_IN), .ZN(n2570) );
  NOR4_X1 U33460 ( .A1(D_REG_9__SCAN_IN), .A2(D_REG_6__SCAN_IN), .A3(
        D_REG_8__SCAN_IN), .A4(D_REG_10__SCAN_IN), .ZN(n2569) );
  NOR4_X1 U33470 ( .A1(D_REG_25__SCAN_IN), .A2(D_REG_26__SCAN_IN), .A3(
        D_REG_27__SCAN_IN), .A4(D_REG_31__SCAN_IN), .ZN(n2568) );
  NOR4_X1 U33480 ( .A1(D_REG_19__SCAN_IN), .A2(D_REG_21__SCAN_IN), .A3(
        D_REG_22__SCAN_IN), .A4(D_REG_24__SCAN_IN), .ZN(n2567) );
  NAND4_X1 U33490 ( .A1(n2570), .A2(n2569), .A3(n2568), .A4(n2567), .ZN(n2571)
         );
  NOR4_X1 U33500 ( .A1(D_REG_28__SCAN_IN), .A2(D_REG_29__SCAN_IN), .A3(n2572), 
        .A4(n2571), .ZN(n2573) );
  NAND3_X1 U33510 ( .A1(n2575), .A2(n2574), .A3(n2573), .ZN(n2576) );
  NAND2_X1 U33520 ( .A1(n2583), .A2(n2576), .ZN(n2807) );
  OAI21_X1 U3353 ( .B1(n2579), .B2(n2578), .A(n2577), .ZN(n2937) );
  AND2_X1 U33540 ( .A1(n2508), .A2(n3898), .ZN(n2809) );
  OR2_X1 U3355 ( .A1(n2809), .A2(n2811), .ZN(n2831) );
  INV_X1 U3356 ( .A(D_REG_0__SCAN_IN), .ZN(n2931) );
  INV_X1 U3357 ( .A(n4202), .ZN(n2581) );
  AND2_X1 U3358 ( .A1(n2581), .A2(n2930), .ZN(n2582) );
  AOI21_X1 U3359 ( .B1(n2583), .B2(n2931), .A(n2582), .ZN(n2861) );
  INV_X1 U3360 ( .A(n2861), .ZN(n2592) );
  AND2_X2 U3361 ( .A1(n2862), .A2(n2592), .ZN(n4419) );
  MUX2_X1 U3362 ( .A(n2584), .B(n4126), .S(n4419), .Z(n2588) );
  NAND2_X1 U3363 ( .A1(n3060), .A2(n2585), .ZN(n3076) );
  NAND2_X1 U3364 ( .A1(n3096), .A2(n3095), .ZN(n4373) );
  OAI21_X1 U3365 ( .B1(n3953), .B2(n2765), .A(n2589), .ZN(n4129) );
  INV_X1 U3366 ( .A(n3031), .ZN(n3014) );
  NAND2_X1 U3367 ( .A1(n4419), .A2(n4411), .ZN(n4197) );
  NAND2_X1 U3368 ( .A1(n2588), .A2(n2587), .ZN(U3511) );
  NAND2_X1 U3369 ( .A1(n2939), .A2(DATAI_26_), .ZN(n2884) );
  INV_X1 U3370 ( .A(n2884), .ZN(n2899) );
  AND2_X1 U3371 ( .A1(n2939), .A2(DATAI_27_), .ZN(n3760) );
  AND2_X1 U3372 ( .A1(n2939), .A2(DATAI_28_), .ZN(n3904) );
  INV_X1 U3373 ( .A(n3904), .ZN(n2865) );
  NAND2_X1 U3374 ( .A1(n2939), .A2(DATAI_29_), .ZN(n3920) );
  AND2_X1 U3375 ( .A1(n2939), .A2(DATAI_30_), .ZN(n4113) );
  NAND2_X1 U3376 ( .A1(n2939), .A2(DATAI_31_), .ZN(n3694) );
  INV_X1 U3377 ( .A(n3694), .ZN(n3689) );
  XNOR2_X1 U3378 ( .A(n4109), .B(n3689), .ZN(n4106) );
  INV_X1 U3379 ( .A(n2590), .ZN(n2808) );
  NAND3_X1 U3380 ( .A1(n2592), .A2(n2591), .A3(n2808), .ZN(n2594) );
  INV_X1 U3381 ( .A(n2829), .ZN(n2593) );
  AOI22_X1 U3382 ( .A1(n4106), .A2(n4213), .B1(n3035), .B2(
        REG2_REG_31__SCAN_IN), .ZN(n2600) );
  NAND2_X1 U3383 ( .A1(n3667), .A2(REG1_REG_31__SCAN_IN), .ZN(n2597) );
  NAND2_X1 U3384 ( .A1(n2478), .A2(REG2_REG_31__SCAN_IN), .ZN(n2596) );
  NAND2_X1 U3385 ( .A1(n3668), .A2(REG0_REG_31__SCAN_IN), .ZN(n2595) );
  NAND3_X1 U3386 ( .A1(n2597), .A2(n2596), .A3(n2595), .ZN(n3819) );
  XNOR2_X1 U3387 ( .A(n2598), .B(IR_REG_27__SCAN_IN), .ZN(n2946) );
  AOI21_X1 U3388 ( .B1(n2946), .B2(B_REG_SCAN_IN), .A(n4379), .ZN(n3913) );
  AND2_X1 U3389 ( .A1(n3819), .A2(n3913), .ZN(n4111) );
  AOI21_X1 U3390 ( .B1(n3689), .B2(n4112), .A(n4111), .ZN(n4164) );
  OR2_X1 U3391 ( .A1(n4164), .A2(n3035), .ZN(n2599) );
  NAND2_X1 U3392 ( .A1(n2600), .A2(n2599), .ZN(U3260) );
  INV_X1 U3393 ( .A(n2603), .ZN(n2601) );
  AND2_X1 U3394 ( .A1(n4205), .A2(n3898), .ZN(n2821) );
  INV_X1 U3395 ( .A(n2821), .ZN(n2605) );
  NAND2_X4 U3396 ( .A1(n2626), .A2(n2607), .ZN(n2802) );
  AND2_X1 U3397 ( .A1(n3085), .A2(n2626), .ZN(n2608) );
  INV_X1 U3398 ( .A(n2604), .ZN(n2609) );
  NAND2_X1 U3399 ( .A1(n2609), .A2(REG1_REG_0__SCAN_IN), .ZN(n2610) );
  NAND2_X1 U3400 ( .A1(n2613), .A2(n2610), .ZN(n3083) );
  INV_X1 U3401 ( .A(n3841), .ZN(n3055) );
  NOR2_X1 U3402 ( .A1(n2604), .A2(n2112), .ZN(n2611) );
  OAI21_X1 U3403 ( .B1(n3055), .B2(n2802), .A(n2612), .ZN(n3082) );
  NAND2_X1 U3404 ( .A1(n3083), .A2(n3082), .ZN(n2615) );
  NAND2_X1 U3405 ( .A1(n2613), .A2(n2763), .ZN(n2614) );
  NOR2_X1 U3406 ( .A1(n2617), .A2(n2616), .ZN(n2618) );
  INV_X1 U3407 ( .A(n2623), .ZN(n2620) );
  OAI22_X1 U3408 ( .A1(n3138), .A2(n2802), .B1(n3052), .B2(n2799), .ZN(n2621)
         );
  NAND2_X1 U3409 ( .A1(n2620), .A2(n2621), .ZN(n2624) );
  INV_X1 U3410 ( .A(n2621), .ZN(n2622) );
  NAND2_X1 U3411 ( .A1(n2623), .A2(n2622), .ZN(n2625) );
  NAND2_X1 U3412 ( .A1(n3047), .A2(n3046), .ZN(n3045) );
  NAND2_X1 U3413 ( .A1(n3045), .A2(n2625), .ZN(n3132) );
  NAND2_X1 U3414 ( .A1(n3134), .A2(n2626), .ZN(n2627) );
  NAND2_X1 U3415 ( .A1(n2628), .A2(n2627), .ZN(n2629) );
  XNOR2_X1 U3416 ( .A(n2631), .B(n2632), .ZN(n3133) );
  NAND2_X1 U3417 ( .A1(n3132), .A2(n3133), .ZN(n3121) );
  OAI22_X1 U3418 ( .A1(n3211), .A2(n2799), .B1(n2798), .B2(n4378), .ZN(n2630)
         );
  XNOR2_X1 U3419 ( .A(n2630), .B(n2763), .ZN(n2635) );
  OAI22_X1 U3420 ( .A1(n3211), .A2(n2802), .B1(n2799), .B2(n4378), .ZN(n2636)
         );
  XNOR2_X1 U3421 ( .A(n2635), .B(n2636), .ZN(n3122) );
  INV_X1 U3422 ( .A(n2631), .ZN(n2633) );
  NAND2_X1 U3423 ( .A1(n2633), .A2(n2632), .ZN(n3123) );
  AND2_X1 U3424 ( .A1(n3122), .A2(n3123), .ZN(n2634) );
  NAND2_X1 U3425 ( .A1(n3121), .A2(n2634), .ZN(n3103) );
  INV_X1 U3426 ( .A(n2635), .ZN(n2637) );
  NAND2_X1 U3427 ( .A1(n2637), .A2(n2636), .ZN(n3104) );
  NAND2_X1 U3428 ( .A1(n3232), .A2(n2626), .ZN(n2638) );
  NAND2_X1 U3429 ( .A1(n2639), .A2(n2638), .ZN(n2640) );
  XNOR2_X1 U3430 ( .A(n2640), .B(n2800), .ZN(n2650) );
  NAND2_X1 U3431 ( .A1(n3836), .A2(n2774), .ZN(n2642) );
  NAND2_X1 U3432 ( .A1(n2642), .A2(n2641), .ZN(n2651) );
  AND2_X1 U3433 ( .A1(n2650), .A2(n2651), .ZN(n3147) );
  INV_X1 U3434 ( .A(n3147), .ZN(n2647) );
  XNOR2_X1 U3435 ( .A(n2644), .B(n2763), .ZN(n2656) );
  INV_X1 U3436 ( .A(n2656), .ZN(n2646) );
  OAI22_X1 U3437 ( .A1(n2643), .A2(n2802), .B1(n2799), .B2(n2645), .ZN(n2655)
         );
  NAND2_X1 U3438 ( .A1(n2646), .A2(n2655), .ZN(n3145) );
  NAND2_X1 U3439 ( .A1(n2647), .A2(n3145), .ZN(n2657) );
  INV_X1 U3440 ( .A(n2657), .ZN(n2648) );
  AND2_X1 U3441 ( .A1(n3104), .A2(n2648), .ZN(n2649) );
  NAND2_X1 U3442 ( .A1(n3103), .A2(n2649), .ZN(n3168) );
  INV_X1 U3443 ( .A(n2650), .ZN(n2653) );
  INV_X1 U3444 ( .A(n2651), .ZN(n2652) );
  NAND2_X1 U3445 ( .A1(n2653), .A2(n2652), .ZN(n3170) );
  INV_X1 U3446 ( .A(n3170), .ZN(n3148) );
  OAI22_X1 U3447 ( .A1(n3286), .A2(n2799), .B1(n2798), .B2(n3318), .ZN(n2654)
         );
  XNOR2_X1 U3448 ( .A(n2654), .B(n2800), .ZN(n2661) );
  OAI22_X1 U3449 ( .A1(n3286), .A2(n2802), .B1(n2799), .B2(n3318), .ZN(n2660)
         );
  XNOR2_X1 U3450 ( .A(n2661), .B(n2660), .ZN(n3172) );
  NOR2_X1 U3451 ( .A1(n3148), .A2(n3172), .ZN(n2658) );
  XNOR2_X1 U3452 ( .A(n2656), .B(n2655), .ZN(n3143) );
  NAND2_X1 U3453 ( .A1(n3168), .A2(n2659), .ZN(n3174) );
  NAND2_X1 U3454 ( .A1(n2661), .A2(n2660), .ZN(n2662) );
  OAI22_X1 U3455 ( .A1(n3319), .A2(n2802), .B1(n2799), .B2(n2663), .ZN(n3160)
         );
  OAI22_X1 U3456 ( .A1(n3319), .A2(n2799), .B1(n2798), .B2(n2663), .ZN(n2664)
         );
  XNOR2_X1 U3457 ( .A(n2664), .B(n2800), .ZN(n3159) );
  NAND2_X1 U34580 ( .A1(n3312), .A2(n2626), .ZN(n2665) );
  NAND2_X1 U34590 ( .A1(n2666), .A2(n2665), .ZN(n2667) );
  XNOR2_X1 U3460 ( .A(n2667), .B(n2763), .ZN(n2672) );
  XNOR2_X1 U3461 ( .A(n2672), .B(n2671), .ZN(n3223) );
  NAND2_X1 U3462 ( .A1(n3342), .A2(n2626), .ZN(n2668) );
  NAND2_X1 U3463 ( .A1(n2669), .A2(n2668), .ZN(n2670) );
  XNOR2_X1 U3464 ( .A(n2670), .B(n2800), .ZN(n2674) );
  XNOR2_X1 U3465 ( .A(n2674), .B(n2675), .ZN(n3248) );
  NAND2_X1 U3466 ( .A1(n2672), .A2(n2671), .ZN(n3249) );
  NAND2_X1 U34670 ( .A1(n3220), .A2(n2673), .ZN(n3247) );
  NAND2_X1 U3468 ( .A1(n2674), .A2(n2676), .ZN(n2677) );
  NAND2_X1 U34690 ( .A1(n3247), .A2(n2677), .ZN(n3269) );
  OAI22_X1 U3470 ( .A1(n2679), .A2(n2799), .B1(n2798), .B2(n3374), .ZN(n2678)
         );
  XNOR2_X1 U34710 ( .A(n2678), .B(n2763), .ZN(n2681) );
  OAI22_X1 U3472 ( .A1(n2679), .A2(n2802), .B1(n2799), .B2(n3374), .ZN(n2682)
         );
  INV_X1 U34730 ( .A(n2682), .ZN(n2680) );
  NAND2_X1 U3474 ( .A1(n2681), .A2(n2680), .ZN(n3267) );
  NAND2_X1 U34750 ( .A1(n3269), .A2(n3267), .ZN(n2684) );
  INV_X1 U3476 ( .A(n2681), .ZN(n2683) );
  NAND2_X1 U34770 ( .A1(n2683), .A2(n2682), .ZN(n3268) );
  OAI22_X1 U3478 ( .A1(n3413), .A2(n2799), .B1(n2798), .B2(n3391), .ZN(n2685)
         );
  XNOR2_X1 U34790 ( .A(n2685), .B(n2800), .ZN(n3258) );
  OAI22_X1 U3480 ( .A1(n3413), .A2(n2802), .B1(n2799), .B2(n3391), .ZN(n3259)
         );
  OAI22_X1 U34810 ( .A1(n3432), .A2(n2799), .B1(n2798), .B2(n3420), .ZN(n2686)
         );
  XNOR2_X1 U3482 ( .A(n2686), .B(n2800), .ZN(n2687) );
  OAI22_X1 U34830 ( .A1(n3432), .A2(n2802), .B1(n2799), .B2(n3420), .ZN(n2688)
         );
  AND2_X1 U3484 ( .A1(n2687), .A2(n2688), .ZN(n3331) );
  INV_X1 U34850 ( .A(n2687), .ZN(n2690) );
  INV_X1 U3486 ( .A(n2688), .ZN(n2689) );
  OAI22_X1 U34870 ( .A1(n3462), .A2(n2799), .B1(n2798), .B2(n2408), .ZN(n2691)
         );
  XNOR2_X1 U3488 ( .A(n2691), .B(n2763), .ZN(n3355) );
  NAND2_X1 U34890 ( .A1(n3354), .A2(n3355), .ZN(n2692) );
  NAND2_X1 U3490 ( .A1(n2692), .A2(n3356), .ZN(n2696) );
  INV_X1 U34910 ( .A(n3354), .ZN(n2694) );
  INV_X1 U3492 ( .A(n3355), .ZN(n2693) );
  NAND2_X1 U34930 ( .A1(n2694), .A2(n2693), .ZN(n2695) );
  OAI22_X1 U3494 ( .A1(n3575), .A2(n2799), .B1(n2798), .B2(n3464), .ZN(n2697)
         );
  XNOR2_X1 U34950 ( .A(n2697), .B(n2800), .ZN(n2698) );
  OAI22_X1 U3496 ( .A1(n3575), .A2(n2802), .B1(n2799), .B2(n3464), .ZN(n3639)
         );
  OAI22_X1 U34970 ( .A1(n4094), .A2(n2799), .B1(n2701), .B2(n2798), .ZN(n2700)
         );
  XNOR2_X1 U3498 ( .A(n2700), .B(n2763), .ZN(n2704) );
  OAI22_X1 U34990 ( .A1(n4094), .A2(n2802), .B1(n2701), .B2(n2799), .ZN(n2702)
         );
  XNOR2_X1 U3500 ( .A(n2704), .B(n2702), .ZN(n3573) );
  INV_X1 U35010 ( .A(n2702), .ZN(n2703) );
  OAI22_X1 U3502 ( .A1(n4075), .A2(n2799), .B1(n4096), .B2(n2798), .ZN(n2705)
         );
  XNOR2_X1 U35030 ( .A(n2705), .B(n2763), .ZN(n3584) );
  OAI22_X1 U3504 ( .A1(n4075), .A2(n2802), .B1(n4096), .B2(n2799), .ZN(n2706)
         );
  INV_X1 U35050 ( .A(n2706), .ZN(n3583) );
  AND2_X1 U35060 ( .A1(n3584), .A2(n3583), .ZN(n2709) );
  INV_X1 U35070 ( .A(n3584), .ZN(n2707) );
  NAND2_X1 U35080 ( .A1(n2707), .A2(n2706), .ZN(n2708) );
  OAI21_X1 U35090 ( .B1(n3582), .B2(n2709), .A(n2708), .ZN(n3629) );
  NAND2_X1 U35100 ( .A1(n4072), .A2(n2626), .ZN(n2710) );
  NAND2_X1 U35110 ( .A1(n2711), .A2(n2710), .ZN(n2712) );
  XNOR2_X1 U35120 ( .A(n2712), .B(n2800), .ZN(n2715) );
  NAND2_X1 U35130 ( .A1(n4090), .A2(n2774), .ZN(n2714) );
  NAND2_X1 U35140 ( .A1(n2714), .A2(n2713), .ZN(n2716) );
  AND2_X1 U35150 ( .A1(n2715), .A2(n2716), .ZN(n3626) );
  INV_X1 U35160 ( .A(n2715), .ZN(n2718) );
  INV_X1 U35170 ( .A(n2716), .ZN(n2717) );
  NAND2_X1 U35180 ( .A1(n2718), .A2(n2717), .ZN(n3625) );
  NAND2_X1 U35190 ( .A1(n3543), .A2(n2626), .ZN(n2719) );
  NAND2_X1 U35200 ( .A1(n2720), .A2(n2719), .ZN(n2721) );
  XNOR2_X1 U35210 ( .A(n2721), .B(n2800), .ZN(n2723) );
  NOR2_X1 U35220 ( .A1(n4057), .A2(n2799), .ZN(n2722) );
  AOI21_X1 U35230 ( .B1(n4073), .B2(n2774), .A(n2722), .ZN(n2724) );
  XNOR2_X1 U35240 ( .A(n2723), .B(n2724), .ZN(n3540) );
  NAND2_X1 U35250 ( .A1(n3539), .A2(n3540), .ZN(n2727) );
  INV_X1 U35260 ( .A(n2723), .ZN(n2725) );
  NAND2_X1 U35270 ( .A1(n2725), .A2(n2724), .ZN(n2726) );
  NAND2_X1 U35280 ( .A1(n2727), .A2(n2726), .ZN(n3606) );
  NAND2_X1 U35290 ( .A1(n3802), .A2(n2626), .ZN(n2728) );
  NAND2_X1 U35300 ( .A1(n2729), .A2(n2728), .ZN(n2730) );
  XNOR2_X1 U35310 ( .A(n2730), .B(n2800), .ZN(n2733) );
  NAND2_X1 U35320 ( .A1(n4052), .A2(n2774), .ZN(n2732) );
  NAND2_X1 U35330 ( .A1(n2732), .A2(n2731), .ZN(n2734) );
  NAND2_X1 U35340 ( .A1(n2733), .A2(n2734), .ZN(n3607) );
  INV_X1 U35350 ( .A(n2733), .ZN(n2736) );
  INV_X1 U35360 ( .A(n2734), .ZN(n2735) );
  NAND2_X1 U35370 ( .A1(n2736), .A2(n2735), .ZN(n3608) );
  OAI22_X1 U35380 ( .A1(n4029), .A2(n2799), .B1(n4010), .B2(n2798), .ZN(n2737)
         );
  XNOR2_X1 U35390 ( .A(n2737), .B(n2800), .ZN(n3548) );
  OAI22_X1 U35400 ( .A1(n4029), .A2(n2802), .B1(n4010), .B2(n2799), .ZN(n3547)
         );
  OAI22_X1 U35410 ( .A1(n4007), .A2(n2799), .B1(n2739), .B2(n2798), .ZN(n2738)
         );
  XNOR2_X1 U35420 ( .A(n2738), .B(n2800), .ZN(n2746) );
  OAI22_X1 U35430 ( .A1(n4007), .A2(n2802), .B1(n2739), .B2(n2799), .ZN(n2747)
         );
  XNOR2_X1 U35440 ( .A(n2746), .B(n2747), .ZN(n3619) );
  NAND2_X1 U35450 ( .A1(n2741), .A2(n2740), .ZN(n3616) );
  INV_X1 U35460 ( .A(n3978), .ZN(n3971) );
  NAND2_X1 U35470 ( .A1(n3971), .A2(n2626), .ZN(n2742) );
  NAND2_X1 U35480 ( .A1(n2743), .A2(n2742), .ZN(n2744) );
  XNOR2_X1 U35490 ( .A(n2744), .B(n2800), .ZN(n2753) );
  NOR2_X1 U35500 ( .A1(n3978), .A2(n2799), .ZN(n2745) );
  AOI21_X1 U35510 ( .B1(n3989), .B2(n2774), .A(n2745), .ZN(n2751) );
  XNOR2_X1 U35520 ( .A(n2753), .B(n2751), .ZN(n3532) );
  INV_X1 U35530 ( .A(n2746), .ZN(n2749) );
  INV_X1 U35540 ( .A(n2747), .ZN(n2748) );
  NAND2_X1 U35550 ( .A1(n2749), .A2(n2748), .ZN(n3530) );
  NAND2_X1 U35560 ( .A1(n3616), .A2(n2750), .ZN(n3531) );
  INV_X1 U35570 ( .A(n2751), .ZN(n2752) );
  NAND2_X1 U35580 ( .A1(n2753), .A2(n2752), .ZN(n2757) );
  OAI22_X1 U35590 ( .A1(n3565), .A2(n2802), .B1(n2799), .B2(n3955), .ZN(n2758)
         );
  INV_X1 U35600 ( .A(n2758), .ZN(n2754) );
  AND2_X1 U35610 ( .A1(n2757), .A2(n2754), .ZN(n2755) );
  NAND2_X1 U35620 ( .A1(n3531), .A2(n2755), .ZN(n3594) );
  OAI22_X1 U35630 ( .A1(n3565), .A2(n2799), .B1(n2798), .B2(n3955), .ZN(n2756)
         );
  XNOR2_X1 U35640 ( .A(n2756), .B(n2800), .ZN(n3596) );
  NAND2_X1 U35650 ( .A1(n3594), .A2(n3596), .ZN(n2760) );
  NAND2_X1 U35660 ( .A1(n3531), .A2(n2757), .ZN(n2759) );
  NAND2_X1 U35670 ( .A1(n2759), .A2(n2758), .ZN(n3593) );
  NAND2_X1 U35680 ( .A1(n3562), .A2(n2626), .ZN(n2761) );
  NAND2_X1 U35690 ( .A1(n2762), .A2(n2761), .ZN(n2764) );
  XNOR2_X1 U35700 ( .A(n2764), .B(n2763), .ZN(n2767) );
  NOR2_X1 U35710 ( .A1(n2765), .A2(n2799), .ZN(n2766) );
  AOI21_X1 U35720 ( .B1(n3949), .B2(n2774), .A(n2766), .ZN(n2768) );
  NAND2_X1 U35730 ( .A1(n2767), .A2(n2768), .ZN(n3557) );
  INV_X1 U35740 ( .A(n2767), .ZN(n2770) );
  INV_X1 U35750 ( .A(n2768), .ZN(n2769) );
  NAND2_X1 U35760 ( .A1(n2770), .A2(n2769), .ZN(n3558) );
  NAND2_X1 U35770 ( .A1(n2899), .A2(n2626), .ZN(n2771) );
  NAND2_X1 U35780 ( .A1(n2772), .A2(n2771), .ZN(n2773) );
  XNOR2_X1 U35790 ( .A(n2773), .B(n2800), .ZN(n2777) );
  NAND2_X1 U35800 ( .A1(n3822), .A2(n2774), .ZN(n2776) );
  NAND2_X1 U35810 ( .A1(n2776), .A2(n2775), .ZN(n2778) );
  AND2_X1 U3582 ( .A1(n2777), .A2(n2778), .ZN(n2893) );
  INV_X1 U3583 ( .A(n2777), .ZN(n2780) );
  INV_X1 U3584 ( .A(n2778), .ZN(n2779) );
  NAND2_X1 U3585 ( .A1(n2780), .A2(n2779), .ZN(n2892) );
  INV_X1 U3586 ( .A(REG3_REG_26__SCAN_IN), .ZN(n2781) );
  INV_X1 U3587 ( .A(REG3_REG_27__SCAN_IN), .ZN(n4571) );
  OAI21_X1 U3588 ( .B1(n2782), .B2(n2781), .A(n4571), .ZN(n2783) );
  NAND2_X1 U3589 ( .A1(n3514), .A2(n2823), .ZN(n2786) );
  AOI22_X1 U3590 ( .A1(n3667), .A2(REG1_REG_27__SCAN_IN), .B1(n3668), .B2(
        REG0_REG_27__SCAN_IN), .ZN(n2785) );
  NAND2_X1 U3591 ( .A1(n2478), .A2(REG2_REG_27__SCAN_IN), .ZN(n2784) );
  INV_X1 U3592 ( .A(n3760), .ZN(n2787) );
  OAI22_X1 U3593 ( .A1(n3761), .A2(n2799), .B1(n2798), .B2(n2787), .ZN(n2788)
         );
  XNOR2_X1 U3594 ( .A(n2788), .B(n2800), .ZN(n2806) );
  OR2_X1 U3595 ( .A1(n3761), .A2(n2802), .ZN(n2790) );
  NAND2_X1 U3596 ( .A1(n2790), .A2(n2789), .ZN(n2805) );
  XNOR2_X1 U3597 ( .A(n2806), .B(n2805), .ZN(n2904) );
  INV_X1 U3598 ( .A(n2792), .ZN(n2791) );
  NAND2_X1 U3599 ( .A1(n2791), .A2(REG3_REG_28__SCAN_IN), .ZN(n3919) );
  INV_X1 U3600 ( .A(REG3_REG_28__SCAN_IN), .ZN(n4471) );
  NAND2_X1 U3601 ( .A1(n2792), .A2(n4471), .ZN(n2793) );
  NAND2_X1 U3602 ( .A1(n3919), .A2(n2793), .ZN(n3523) );
  OR2_X1 U3603 ( .A1(n3523), .A2(n2794), .ZN(n2797) );
  AOI22_X1 U3604 ( .A1(n3667), .A2(REG1_REG_28__SCAN_IN), .B1(n3668), .B2(
        REG0_REG_28__SCAN_IN), .ZN(n2796) );
  NAND2_X1 U3605 ( .A1(n2478), .A2(REG2_REG_28__SCAN_IN), .ZN(n2795) );
  OAI22_X1 U3606 ( .A1(n3916), .A2(n2799), .B1(n2865), .B2(n2798), .ZN(n2801)
         );
  XNOR2_X1 U3607 ( .A(n2801), .B(n2800), .ZN(n2804) );
  OAI22_X1 U3608 ( .A1(n3916), .A2(n2802), .B1(n2865), .B2(n2799), .ZN(n2803)
         );
  XNOR2_X1 U3609 ( .A(n2804), .B(n2803), .ZN(n2819) );
  INV_X1 U3610 ( .A(n2819), .ZN(n2814) );
  NAND2_X1 U3611 ( .A1(n2806), .A2(n2805), .ZN(n2817) );
  NAND3_X1 U3612 ( .A1(n2808), .A2(n2861), .A3(n2807), .ZN(n2830) );
  INV_X1 U3613 ( .A(n2927), .ZN(n2935) );
  INV_X1 U3614 ( .A(n2809), .ZN(n2810) );
  NAND2_X1 U3615 ( .A1(n3031), .A2(n2810), .ZN(n2812) );
  NAND2_X1 U3616 ( .A1(n2812), .A2(n2811), .ZN(n2813) );
  NAND2_X1 U3617 ( .A1(n2814), .A2(n2193), .ZN(n2815) );
  NAND3_X1 U3618 ( .A1(n2816), .A2(n3609), .A3(n2819), .ZN(n2837) );
  INV_X1 U3619 ( .A(n2817), .ZN(n2818) );
  NAND3_X1 U3620 ( .A1(n2819), .A2(n3609), .A3(n2818), .ZN(n2836) );
  OAI21_X1 U3621 ( .B1(n2820), .B2(n4377), .A(n4590), .ZN(n3635) );
  INV_X1 U3622 ( .A(n2956), .ZN(n4201) );
  NAND2_X1 U3623 ( .A1(n2131), .A2(n4201), .ZN(n2822) );
  INV_X1 U3624 ( .A(REG2_REG_29__SCAN_IN), .ZN(n3923) );
  INV_X1 U3625 ( .A(n3919), .ZN(n2824) );
  NAND2_X1 U3626 ( .A1(n2824), .A2(n2823), .ZN(n2826) );
  AOI22_X1 U3627 ( .A1(REG1_REG_29__SCAN_IN), .A2(n3667), .B1(n3668), .B2(
        REG0_REG_29__SCAN_IN), .ZN(n2825) );
  OAI211_X1 U3628 ( .C1(n2255), .C2(n3923), .A(n2826), .B(n2825), .ZN(n3820)
         );
  NAND2_X1 U3629 ( .A1(n2131), .A2(n2956), .ZN(n2827) );
  OR2_X1 U3630 ( .A1(n2830), .A2(n2827), .ZN(n3642) );
  AOI22_X1 U3631 ( .A1(n3820), .A2(n3630), .B1(REG3_REG_28__SCAN_IN), .B2(
        U3149), .ZN(n2828) );
  OAI21_X1 U3632 ( .B1(n3761), .B2(n3632), .A(n2828), .ZN(n2834) );
  NAND2_X1 U3633 ( .A1(n2830), .A2(n2829), .ZN(n3040) );
  NAND4_X1 U3634 ( .A1(n3040), .A2(n2831), .A3(n2937), .A4(n2604), .ZN(n2832)
         );
  NAND2_X1 U3635 ( .A1(n2832), .A2(STATE_REG_SCAN_IN), .ZN(n3644) );
  NOR2_X1 U3636 ( .A1(n3644), .A2(n3523), .ZN(n2833) );
  AOI211_X1 U3637 ( .C1(n3904), .C2(n3635), .A(n2834), .B(n2833), .ZN(n2835)
         );
  NAND3_X1 U3638 ( .A1(n2838), .A2(n2837), .A3(n2195), .ZN(U3217) );
  NAND2_X1 U3639 ( .A1(n3949), .A2(n3562), .ZN(n2843) );
  AND2_X1 U3640 ( .A1(n2839), .A2(n2843), .ZN(n2872) );
  NOR2_X1 U3641 ( .A1(n2849), .A2(n2884), .ZN(n2848) );
  INV_X1 U3642 ( .A(n2848), .ZN(n2840) );
  AND2_X1 U3643 ( .A1(n2872), .A2(n2840), .ZN(n2841) );
  NAND2_X1 U3644 ( .A1(n2842), .A2(n2841), .ZN(n3507) );
  INV_X1 U3645 ( .A(n2843), .ZN(n2847) );
  OR2_X1 U3646 ( .A1(n3949), .A2(n3562), .ZN(n2844) );
  AND2_X1 U3647 ( .A1(n2845), .A2(n2844), .ZN(n2846) );
  OR2_X1 U3648 ( .A1(n2847), .A2(n2846), .ZN(n2870) );
  OR2_X1 U3649 ( .A1(n2848), .A2(n2870), .ZN(n2851) );
  NAND2_X1 U3650 ( .A1(n2849), .A2(n2884), .ZN(n2850) );
  AND2_X1 U3651 ( .A1(n2851), .A2(n2850), .ZN(n3506) );
  INV_X1 U3652 ( .A(n3761), .ZN(n3821) );
  OR2_X1 U3653 ( .A1(n3821), .A2(n3760), .ZN(n2852) );
  AND2_X1 U3654 ( .A1(n3506), .A2(n2852), .ZN(n2853) );
  NAND2_X1 U3655 ( .A1(n3821), .A2(n3760), .ZN(n2854) );
  INV_X1 U3656 ( .A(n3916), .ZN(n3903) );
  NAND2_X1 U3657 ( .A1(n3903), .A2(n2865), .ZN(n3908) );
  NAND2_X1 U3658 ( .A1(n3916), .A2(n3904), .ZN(n3677) );
  NAND2_X1 U3659 ( .A1(n3908), .A2(n3677), .ZN(n3905) );
  AND2_X1 U3660 ( .A1(n3780), .A2(n2855), .ZN(n3757) );
  NAND2_X1 U3661 ( .A1(n2856), .A2(n3757), .ZN(n2876) );
  OR2_X1 U3662 ( .A1(n3822), .A2(n2884), .ZN(n2873) );
  AND2_X1 U3663 ( .A1(n2875), .A2(n2873), .ZN(n3765) );
  NAND2_X1 U3664 ( .A1(n2876), .A2(n3765), .ZN(n2857) );
  NAND2_X1 U3665 ( .A1(n3822), .A2(n2884), .ZN(n3676) );
  NAND2_X1 U3666 ( .A1(n2857), .A2(n3676), .ZN(n3509) );
  XNOR2_X1 U3667 ( .A(n3761), .B(n3760), .ZN(n3804) );
  NAND2_X1 U3668 ( .A1(n3761), .A2(n3760), .ZN(n3678) );
  OAI21_X1 U3669 ( .B1(n3509), .B2(n3804), .A(n3678), .ZN(n3909) );
  XOR2_X1 U3670 ( .A(n3905), .B(n3909), .Z(n2860) );
  INV_X1 U3671 ( .A(n4086), .ZN(n4387) );
  AOI22_X1 U3672 ( .A1(n3820), .A2(n4089), .B1(n4112), .B2(n3904), .ZN(n2858)
         );
  OAI21_X1 U3673 ( .B1(n3761), .B2(n4093), .A(n2858), .ZN(n2859) );
  AOI21_X1 U3674 ( .B1(n2860), .B2(n4049), .A(n2859), .ZN(n3522) );
  OAI21_X1 U3675 ( .B1(n3521), .B2(n4406), .A(n3522), .ZN(n2867) );
  AND2_X2 U3676 ( .A1(n2862), .A2(n2861), .ZN(n4433) );
  INV_X1 U3677 ( .A(n2863), .ZN(n2866) );
  INV_X1 U3678 ( .A(n3921), .ZN(n2864) );
  OAI21_X1 U3679 ( .B1(n3516), .B2(n2865), .A(n2864), .ZN(n3526) );
  NAND2_X1 U3680 ( .A1(n4433), .A2(n4411), .ZN(n4159) );
  NAND2_X1 U3681 ( .A1(n2866), .A2(n2191), .ZN(U3546) );
  INV_X1 U3682 ( .A(n2868), .ZN(n2869) );
  NAND2_X1 U3683 ( .A1(n2869), .A2(n2192), .ZN(U3514) );
  NAND2_X1 U3684 ( .A1(n2873), .A2(n3676), .ZN(n3803) );
  XNOR2_X1 U3685 ( .A(n2874), .B(n3803), .ZN(n3935) );
  NAND2_X1 U3686 ( .A1(n2876), .A2(n2875), .ZN(n2878) );
  INV_X1 U3687 ( .A(n3803), .ZN(n2877) );
  XNOR2_X1 U3688 ( .A(n2878), .B(n2877), .ZN(n2882) );
  NAND2_X1 U3689 ( .A1(n2899), .A2(n4112), .ZN(n2880) );
  INV_X1 U3690 ( .A(n4093), .ZN(n4384) );
  NAND2_X1 U3691 ( .A1(n3949), .A2(n4384), .ZN(n2879) );
  OAI211_X1 U3692 ( .C1(n3761), .C2(n4379), .A(n2880), .B(n2879), .ZN(n2881)
         );
  AOI21_X1 U3693 ( .B1(n2882), .B2(n4049), .A(n2881), .ZN(n3928) );
  OAI21_X1 U3694 ( .B1(n3935), .B2(n4406), .A(n3928), .ZN(n2888) );
  INV_X1 U3695 ( .A(n2883), .ZN(n2887) );
  INV_X1 U3696 ( .A(n2589), .ZN(n2885) );
  OAI21_X1 U3697 ( .B1(n2885), .B2(n2884), .A(n2027), .ZN(n3931) );
  NAND2_X1 U3698 ( .A1(n2887), .A2(n2886), .ZN(U3544) );
  INV_X1 U3699 ( .A(n2889), .ZN(n2891) );
  NAND2_X1 U3700 ( .A1(n2891), .A2(n2890), .ZN(U3512) );
  INV_X1 U3701 ( .A(n2892), .ZN(n2894) );
  NOR2_X1 U3702 ( .A1(n2894), .A2(n2893), .ZN(n2895) );
  XNOR2_X1 U3703 ( .A(n2896), .B(n2895), .ZN(n2897) );
  INV_X1 U3704 ( .A(n3929), .ZN(n2898) );
  INV_X1 U3705 ( .A(n3635), .ZN(n3053) );
  NAND2_X1 U3706 ( .A1(U3149), .A2(REG3_REG_26__SCAN_IN), .ZN(n2901) );
  INV_X1 U3707 ( .A(n3632), .ZN(n3640) );
  NAND2_X1 U3708 ( .A1(n3640), .A2(n3949), .ZN(n2900) );
  OAI211_X1 U3709 ( .C1(n3761), .C2(n3642), .A(n2901), .B(n2900), .ZN(n2902)
         );
  INV_X1 U3710 ( .A(n2902), .ZN(n2903) );
  NAND4_X1 U3711 ( .A1(n2029), .A2(n2198), .A3(n2188), .A4(n2903), .ZN(U3237)
         );
  INV_X1 U3712 ( .A(n2904), .ZN(n2905) );
  XNOR2_X1 U3713 ( .A(n2906), .B(n2905), .ZN(n2907) );
  NAND2_X1 U3714 ( .A1(n2907), .A2(n3609), .ZN(n2916) );
  NAND2_X1 U3715 ( .A1(U3149), .A2(REG3_REG_27__SCAN_IN), .ZN(n2909) );
  NAND2_X1 U3716 ( .A1(n3640), .A2(n3822), .ZN(n2908) );
  OAI211_X1 U3717 ( .C1(n3916), .C2(n3642), .A(n2909), .B(n2908), .ZN(n2911)
         );
  AND2_X1 U3718 ( .A1(n3647), .A2(n3760), .ZN(n2910) );
  NOR2_X1 U3719 ( .A1(n2911), .A2(n2910), .ZN(n2914) );
  INV_X1 U3720 ( .A(n3514), .ZN(n2912) );
  OR2_X1 U3721 ( .A1(n2912), .A2(n3644), .ZN(n2913) );
  AND2_X1 U3722 ( .A1(n2914), .A2(n2913), .ZN(n2915) );
  NAND2_X1 U3723 ( .A1(n2916), .A2(n2915), .ZN(U3211) );
  INV_X1 U3724 ( .A(n4340), .ZN(n2929) );
  NOR2_X1 U3725 ( .A1(n2604), .A2(n2929), .ZN(U4043) );
  INV_X1 U3726 ( .A(DATAI_21_), .ZN(n4555) );
  NAND2_X1 U3727 ( .A1(n3808), .A2(STATE_REG_SCAN_IN), .ZN(n2917) );
  OAI21_X1 U3728 ( .B1(STATE_REG_SCAN_IN), .B2(n4555), .A(n2917), .ZN(U3331)
         );
  INV_X1 U3729 ( .A(DATAI_3_), .ZN(n2918) );
  MUX2_X1 U3730 ( .A(n2965), .B(n2918), .S(U3149), .Z(n2919) );
  INV_X1 U3731 ( .A(n2919), .ZN(U3349) );
  MUX2_X1 U3732 ( .A(n2920), .B(n3192), .S(STATE_REG_SCAN_IN), .Z(n2921) );
  INV_X1 U3733 ( .A(n2921), .ZN(U3344) );
  INV_X1 U3734 ( .A(DATAI_27_), .ZN(n2923) );
  NAND2_X1 U3735 ( .A1(n2946), .A2(STATE_REG_SCAN_IN), .ZN(n2922) );
  OAI21_X1 U3736 ( .B1(STATE_REG_SCAN_IN), .B2(n2923), .A(n2922), .ZN(U3325)
         );
  INV_X1 U3737 ( .A(DATAI_29_), .ZN(n2926) );
  NAND2_X1 U3738 ( .A1(n2924), .A2(STATE_REG_SCAN_IN), .ZN(n2925) );
  OAI21_X1 U3739 ( .B1(STATE_REG_SCAN_IN), .B2(n2926), .A(n2925), .ZN(U3323)
         );
  NAND2_X1 U3740 ( .A1(n2928), .A2(n2927), .ZN(n4338) );
  NOR2_X1 U3741 ( .A1(n2929), .A2(n4202), .ZN(n2933) );
  AOI22_X1 U3742 ( .A1(n4338), .A2(n2931), .B1(n2933), .B2(n2930), .ZN(U3458)
         );
  INV_X1 U3743 ( .A(D_REG_1__SCAN_IN), .ZN(n4491) );
  AOI22_X1 U3744 ( .A1(n4338), .A2(n4491), .B1(n2933), .B2(n2932), .ZN(U3459)
         );
  INV_X1 U3745 ( .A(n2937), .ZN(n2934) );
  NAND2_X1 U3746 ( .A1(n2934), .A2(STATE_REG_SCAN_IN), .ZN(n3817) );
  NAND2_X1 U3747 ( .A1(n2935), .A2(n3817), .ZN(n2945) );
  NAND2_X1 U3748 ( .A1(n2937), .A2(n2936), .ZN(n2938) );
  AND2_X1 U3749 ( .A1(n2939), .A2(n2938), .ZN(n2944) );
  INV_X1 U3750 ( .A(n2944), .ZN(n2940) );
  NOR2_X1 U3751 ( .A1(n4320), .A2(U4043), .ZN(U3148) );
  INV_X1 U3752 ( .A(REG2_REG_0__SCAN_IN), .ZN(n2941) );
  AND2_X1 U3753 ( .A1(n2946), .A2(n2941), .ZN(n2942) );
  NOR2_X1 U3754 ( .A1(n2956), .A2(n2942), .ZN(n3858) );
  OAI21_X1 U3755 ( .B1(REG1_REG_0__SCAN_IN), .B2(n2946), .A(n3858), .ZN(n2943)
         );
  MUX2_X1 U3756 ( .A(n2943), .B(n3858), .S(IR_REG_0__SCAN_IN), .Z(n2951) );
  INV_X1 U3757 ( .A(n2957), .ZN(n2950) );
  INV_X1 U3758 ( .A(n2946), .ZN(n3851) );
  INV_X1 U3759 ( .A(REG1_REG_0__SCAN_IN), .ZN(n2947) );
  NAND3_X1 U3760 ( .A1(n4314), .A2(IR_REG_0__SCAN_IN), .A3(n2947), .ZN(n2949)
         );
  AOI22_X1 U3761 ( .A1(n4320), .A2(ADDR_REG_0__SCAN_IN), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n2948) );
  OAI211_X1 U3762 ( .C1(n2951), .C2(n2950), .A(n2949), .B(n2948), .ZN(U3240)
         );
  INV_X1 U3763 ( .A(REG1_REG_2__SCAN_IN), .ZN(n2952) );
  INV_X1 U3764 ( .A(REG1_REG_1__SCAN_IN), .ZN(n2953) );
  MUX2_X1 U3765 ( .A(n2953), .B(REG1_REG_1__SCAN_IN), .S(n2958), .Z(n3843) );
  AND2_X1 U3766 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n3844)
         );
  NAND2_X1 U3767 ( .A1(n4212), .A2(REG1_REG_1__SCAN_IN), .ZN(n2954) );
  NAND2_X1 U3768 ( .A1(n4211), .A2(REG1_REG_2__SCAN_IN), .ZN(n2955) );
  XOR2_X1 U3769 ( .A(REG1_REG_3__SCAN_IN), .B(n2972), .Z(n2962) );
  NOR2_X1 U3770 ( .A1(n2956), .A2(n3851), .ZN(n3855) );
  XNOR2_X1 U3771 ( .A(n2958), .B(REG2_REG_1__SCAN_IN), .ZN(n3846) );
  AND2_X1 U3772 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n3854)
         );
  NAND2_X1 U3773 ( .A1(n3846), .A2(n3854), .ZN(n3845) );
  NAND2_X1 U3774 ( .A1(n4212), .A2(REG2_REG_1__SCAN_IN), .ZN(n2959) );
  NAND2_X1 U3775 ( .A1(n3845), .A2(n2959), .ZN(n3859) );
  NAND2_X1 U3776 ( .A1(n4211), .A2(REG2_REG_2__SCAN_IN), .ZN(n2960) );
  XNOR2_X1 U3777 ( .A(n2967), .B(n2965), .ZN(n2966) );
  XOR2_X1 U3778 ( .A(n2966), .B(REG2_REG_3__SCAN_IN), .Z(n2961) );
  AOI22_X1 U3779 ( .A1(n4314), .A2(n2962), .B1(n4316), .B2(n2961), .ZN(n2964)
         );
  INV_X1 U3780 ( .A(REG3_REG_3__SCAN_IN), .ZN(n3097) );
  NOR2_X1 U3781 ( .A1(STATE_REG_SCAN_IN), .A2(n3097), .ZN(n3135) );
  AOI21_X1 U3782 ( .B1(n4320), .B2(ADDR_REG_3__SCAN_IN), .A(n3135), .ZN(n2963)
         );
  OAI211_X1 U3783 ( .C1(n2965), .C2(n4319), .A(n2964), .B(n2963), .ZN(U3243)
         );
  INV_X1 U3784 ( .A(n3011), .ZN(n4210) );
  NAND2_X1 U3785 ( .A1(n2966), .A2(REG2_REG_3__SCAN_IN), .ZN(n2969) );
  NAND2_X1 U3786 ( .A1(n2967), .A2(n2973), .ZN(n2968) );
  NAND2_X1 U3787 ( .A1(n2969), .A2(n2968), .ZN(n2970) );
  INV_X1 U3788 ( .A(n4222), .ZN(n2977) );
  INV_X1 U3789 ( .A(REG2_REG_5__SCAN_IN), .ZN(n2971) );
  MUX2_X1 U3790 ( .A(REG2_REG_5__SCAN_IN), .B(n2971), .S(n3011), .Z(n2036) );
  XNOR2_X1 U3791 ( .A(n2989), .B(n4209), .ZN(n2991) );
  XNOR2_X1 U3792 ( .A(n2991), .B(REG2_REG_6__SCAN_IN), .ZN(n2988) );
  INV_X1 U3793 ( .A(n4316), .ZN(n4327) );
  NAND2_X1 U3794 ( .A1(n2972), .A2(REG1_REG_3__SCAN_IN), .ZN(n2976) );
  NAND2_X1 U3795 ( .A1(n2974), .A2(n2973), .ZN(n2975) );
  NAND2_X1 U3796 ( .A1(n2976), .A2(n2975), .ZN(n2978) );
  XNOR2_X1 U3797 ( .A(n2978), .B(n2977), .ZN(n4220) );
  NAND2_X1 U3798 ( .A1(n4220), .A2(REG1_REG_4__SCAN_IN), .ZN(n2980) );
  NAND2_X1 U3799 ( .A1(n2978), .A2(n4222), .ZN(n2979) );
  NAND2_X1 U3800 ( .A1(n2980), .A2(n2979), .ZN(n3007) );
  INV_X1 U3801 ( .A(REG1_REG_5__SCAN_IN), .ZN(n2981) );
  MUX2_X1 U3802 ( .A(n2981), .B(REG1_REG_5__SCAN_IN), .S(n3011), .Z(n3008) );
  NAND2_X1 U3803 ( .A1(n3007), .A2(n3008), .ZN(n3006) );
  NAND2_X1 U3804 ( .A1(n4210), .A2(REG1_REG_5__SCAN_IN), .ZN(n2982) );
  INV_X1 U3805 ( .A(n4209), .ZN(n2984) );
  XOR2_X1 U3806 ( .A(n2995), .B(REG1_REG_6__SCAN_IN), .Z(n2986) );
  AND2_X1 U3807 ( .A1(U3149), .A2(REG3_REG_6__SCAN_IN), .ZN(n3151) );
  AOI21_X1 U3808 ( .B1(n4320), .B2(ADDR_REG_6__SCAN_IN), .A(n3151), .ZN(n2983)
         );
  OAI21_X1 U3809 ( .B1(n4319), .B2(n2984), .A(n2983), .ZN(n2985) );
  AOI21_X1 U3810 ( .B1(n4314), .B2(n2986), .A(n2985), .ZN(n2987) );
  OAI21_X1 U3811 ( .B1(n2988), .B2(n4327), .A(n2987), .ZN(U3246) );
  INV_X1 U3812 ( .A(n2989), .ZN(n2990) );
  AOI22_X1 U3813 ( .A1(n2991), .A2(REG2_REG_6__SCAN_IN), .B1(n4209), .B2(n2990), .ZN(n3025) );
  INV_X1 U3814 ( .A(REG2_REG_7__SCAN_IN), .ZN(n4492) );
  MUX2_X1 U3815 ( .A(n4492), .B(REG2_REG_7__SCAN_IN), .S(n4208), .Z(n3024) );
  INV_X1 U3816 ( .A(REG2_REG_8__SCAN_IN), .ZN(n3290) );
  XNOR2_X1 U3817 ( .A(n3183), .B(n3290), .ZN(n3003) );
  NAND2_X1 U3818 ( .A1(REG3_REG_8__SCAN_IN), .A2(U3149), .ZN(n3162) );
  INV_X1 U3819 ( .A(n3162), .ZN(n2994) );
  NOR2_X1 U3820 ( .A1(n4319), .A2(n3192), .ZN(n2993) );
  AOI211_X1 U3821 ( .C1(n4320), .C2(ADDR_REG_8__SCAN_IN), .A(n2994), .B(n2993), 
        .ZN(n3002) );
  NAND2_X1 U3822 ( .A1(n2995), .A2(REG1_REG_6__SCAN_IN), .ZN(n2998) );
  NAND2_X1 U3823 ( .A1(n2996), .A2(n4209), .ZN(n2997) );
  AND2_X1 U3824 ( .A1(n4208), .A2(REG1_REG_7__SCAN_IN), .ZN(n2999) );
  OR2_X1 U3825 ( .A1(n4208), .A2(REG1_REG_7__SCAN_IN), .ZN(n3000) );
  OAI211_X1 U3826 ( .C1(n2026), .C2(REG1_REG_8__SCAN_IN), .A(n3195), .B(n4314), 
        .ZN(n3001) );
  OAI211_X1 U3827 ( .C1(n3003), .C2(n4327), .A(n3002), .B(n3001), .ZN(U3248)
         );
  AOI211_X1 U3828 ( .C1(n3004), .C2(n2036), .A(n2052), .B(n4327), .ZN(n3013)
         );
  NAND2_X1 U3829 ( .A1(U3149), .A2(REG3_REG_5__SCAN_IN), .ZN(n3105) );
  INV_X1 U3830 ( .A(n3105), .ZN(n3005) );
  AOI21_X1 U3831 ( .B1(n4320), .B2(ADDR_REG_5__SCAN_IN), .A(n3005), .ZN(n3010)
         );
  OAI211_X1 U3832 ( .C1(n3008), .C2(n3007), .A(n4314), .B(n3006), .ZN(n3009)
         );
  OAI211_X1 U3833 ( .C1(n4319), .C2(n3011), .A(n3010), .B(n3009), .ZN(n3012)
         );
  OR2_X1 U3834 ( .A1(n3013), .A2(n3012), .ZN(U3245) );
  AND2_X1 U3835 ( .A1(n3841), .A2(n2585), .ZN(n3698) );
  OR2_X1 U3836 ( .A1(n3698), .A2(n3701), .ZN(n3016) );
  INV_X1 U3837 ( .A(n3016), .ZN(n3776) );
  OAI22_X1 U3838 ( .A1(n3776), .A2(n4414), .B1(n2585), .B2(n3014), .ZN(n3018)
         );
  INV_X1 U3839 ( .A(n4380), .ZN(n3075) );
  OAI21_X1 U3840 ( .B1(n3075), .B2(n4086), .A(n3016), .ZN(n3017) );
  OAI21_X1 U3841 ( .B1(n3015), .B2(n4379), .A(n3017), .ZN(n3034) );
  NOR2_X1 U3842 ( .A1(n3018), .A2(n3034), .ZN(n4359) );
  NAND2_X1 U3843 ( .A1(n4431), .A2(REG1_REG_0__SCAN_IN), .ZN(n3019) );
  OAI21_X1 U3844 ( .B1(n4359), .B2(n4431), .A(n3019), .ZN(U3518) );
  INV_X1 U3845 ( .A(REG1_REG_7__SCAN_IN), .ZN(n4427) );
  XNOR2_X1 U3846 ( .A(n4208), .B(n4427), .ZN(n3020) );
  XNOR2_X1 U3847 ( .A(n3021), .B(n3020), .ZN(n3029) );
  NAND2_X1 U3848 ( .A1(n4320), .A2(ADDR_REG_7__SCAN_IN), .ZN(n3022) );
  NAND2_X1 U3849 ( .A1(U3149), .A2(REG3_REG_7__SCAN_IN), .ZN(n3176) );
  NAND2_X1 U3850 ( .A1(n3022), .A2(n3176), .ZN(n3027) );
  AOI211_X1 U3851 ( .C1(n3025), .C2(n3024), .A(n4327), .B(n3023), .ZN(n3026)
         );
  AOI211_X1 U3852 ( .C1(n4332), .C2(n4208), .A(n3027), .B(n3026), .ZN(n3028)
         );
  OAI21_X1 U3853 ( .B1(n4321), .B2(n3029), .A(n3028), .ZN(U3247) );
  OR2_X1 U3854 ( .A1(n2603), .A2(n3898), .ZN(n3030) );
  AOI21_X1 U3855 ( .B1(n3031), .B2(n3898), .A(n4112), .ZN(n3032) );
  NOR2_X1 U3856 ( .A1(n2585), .A2(n3032), .ZN(n3033) );
  INV_X2 U3857 ( .A(n3035), .ZN(n4595) );
  OAI21_X1 U3858 ( .B1(n3034), .B2(n3033), .A(n4595), .ZN(n3037) );
  INV_X1 U3859 ( .A(n4590), .ZN(n4098) );
  AOI22_X1 U3860 ( .A1(n3035), .A2(REG2_REG_0__SCAN_IN), .B1(
        REG3_REG_0__SCAN_IN), .B2(n4098), .ZN(n3036) );
  OAI211_X1 U3861 ( .C1(n3776), .C2(n3445), .A(n3037), .B(n3036), .ZN(U3290)
         );
  XNOR2_X1 U3862 ( .A(n3038), .B(n3039), .ZN(n3044) );
  NAND2_X1 U3863 ( .A1(n3040), .A2(n2199), .ZN(n3084) );
  OAI22_X1 U3864 ( .A1(n3055), .A2(n3632), .B1(n3642), .B2(n3138), .ZN(n3042)
         );
  NOR2_X1 U3865 ( .A1(n3053), .A2(n3060), .ZN(n3041) );
  AOI211_X1 U3866 ( .C1(REG3_REG_1__SCAN_IN), .C2(n3084), .A(n3042), .B(n3041), 
        .ZN(n3043) );
  OAI21_X1 U3867 ( .B1(n3044), .B2(n3650), .A(n3043), .ZN(U3219) );
  OAI21_X1 U3868 ( .B1(n3047), .B2(n3046), .A(n3045), .ZN(n3048) );
  NAND2_X1 U3869 ( .A1(n3048), .A2(n3609), .ZN(n3051) );
  OAI22_X1 U3870 ( .A1(n3126), .A2(n3642), .B1(n3632), .B2(n3015), .ZN(n3049)
         );
  AOI21_X1 U3871 ( .B1(REG3_REG_2__SCAN_IN), .B2(n3084), .A(n3049), .ZN(n3050)
         );
  OAI211_X1 U3872 ( .C1(n3053), .C2(n3052), .A(n3051), .B(n3050), .ZN(U3234)
         );
  XNOR2_X1 U3873 ( .A(n3054), .B(n2519), .ZN(n4361) );
  OAI21_X1 U3874 ( .B1(n3774), .B2(n3701), .A(n3070), .ZN(n3058) );
  NOR2_X1 U3875 ( .A1(n3055), .A2(n4093), .ZN(n3057) );
  OAI22_X1 U3876 ( .A1(n3138), .A2(n4379), .B1(n4377), .B2(n3060), .ZN(n3056)
         );
  AOI211_X1 U3877 ( .C1(n3058), .C2(n4086), .A(n3057), .B(n3056), .ZN(n3059)
         );
  OAI21_X1 U3878 ( .B1(n4361), .B2(n4380), .A(n3059), .ZN(n4363) );
  NAND2_X1 U3879 ( .A1(n4363), .A2(n4595), .ZN(n3066) );
  OAI21_X1 U3880 ( .B1(n2585), .B2(n3060), .A(n3076), .ZN(n4360) );
  INV_X1 U3881 ( .A(n4360), .ZN(n3064) );
  INV_X1 U3882 ( .A(REG3_REG_1__SCAN_IN), .ZN(n3061) );
  OAI22_X1 U3883 ( .A1(n4595), .A2(n3062), .B1(n3061), .B2(n4590), .ZN(n3063)
         );
  AOI21_X1 U3884 ( .B1(n4213), .B2(n3064), .A(n3063), .ZN(n3065) );
  OAI211_X1 U3885 ( .C1(n4361), .C2(n3445), .A(n3066), .B(n3065), .ZN(U3289)
         );
  OAI21_X1 U3886 ( .B1(n3067), .B2(n2520), .A(n3068), .ZN(n3111) );
  AOI22_X1 U3887 ( .A1(n4383), .A2(n4089), .B1(n2272), .B2(n4112), .ZN(n3069)
         );
  OAI21_X1 U3888 ( .B1(n3015), .B2(n4093), .A(n3069), .ZN(n3074) );
  NAND3_X1 U3889 ( .A1(n3070), .A2(n2520), .A3(n3702), .ZN(n3071) );
  AOI21_X1 U3890 ( .B1(n3072), .B2(n3071), .A(n4387), .ZN(n3073) );
  AOI211_X1 U3891 ( .C1(n3075), .C2(n3111), .A(n3074), .B(n3073), .ZN(n3112)
         );
  INV_X1 U3892 ( .A(n3445), .ZN(n3425) );
  INV_X1 U3893 ( .A(n3096), .ZN(n3078) );
  NAND2_X1 U3894 ( .A1(n3076), .A2(n2272), .ZN(n3077) );
  NAND2_X1 U3895 ( .A1(n3078), .A2(n3077), .ZN(n3117) );
  AOI22_X1 U3896 ( .A1(n3035), .A2(REG2_REG_2__SCAN_IN), .B1(
        REG3_REG_2__SCAN_IN), .B2(n4098), .ZN(n3079) );
  OAI21_X1 U3897 ( .B1(n4101), .B2(n3117), .A(n3079), .ZN(n3080) );
  AOI21_X1 U3898 ( .B1(n3111), .B2(n3425), .A(n3080), .ZN(n3081) );
  OAI21_X1 U3899 ( .B1(n3112), .B2(n3035), .A(n3081), .ZN(U3288) );
  XNOR2_X1 U3900 ( .A(n3083), .B(n3082), .ZN(n3852) );
  AOI22_X1 U3901 ( .A1(n3630), .A2(n3840), .B1(n3084), .B2(REG3_REG_0__SCAN_IN), .ZN(n3087) );
  NAND2_X1 U3902 ( .A1(n3647), .A2(n3085), .ZN(n3086) );
  OAI211_X1 U3903 ( .C1(n3852), .C2(n3650), .A(n3087), .B(n3086), .ZN(U3229)
         );
  XNOR2_X1 U3904 ( .A(n3088), .B(n3789), .ZN(n4366) );
  OAI21_X1 U3905 ( .B1(n3789), .B2(n3090), .A(n3089), .ZN(n3093) );
  AOI22_X1 U3906 ( .A1(n3838), .A2(n4089), .B1(n4112), .B2(n3134), .ZN(n3091)
         );
  OAI21_X1 U3907 ( .B1(n3138), .B2(n4093), .A(n3091), .ZN(n3092) );
  AOI21_X1 U3908 ( .B1(n3093), .B2(n4086), .A(n3092), .ZN(n3094) );
  OAI21_X1 U3909 ( .B1(n4366), .B2(n4380), .A(n3094), .ZN(n4368) );
  INV_X1 U3910 ( .A(n4368), .ZN(n3102) );
  INV_X1 U3911 ( .A(n4366), .ZN(n3100) );
  OAI21_X1 U3912 ( .B1(n3096), .B2(n3095), .A(n4373), .ZN(n4365) );
  AOI22_X1 U3913 ( .A1(n3035), .A2(REG2_REG_3__SCAN_IN), .B1(n4098), .B2(n3097), .ZN(n3098) );
  OAI21_X1 U3914 ( .B1(n4365), .B2(n4101), .A(n3098), .ZN(n3099) );
  AOI21_X1 U3915 ( .B1(n3100), .B2(n3425), .A(n3099), .ZN(n3101) );
  OAI21_X1 U3916 ( .B1(n3102), .B2(n3035), .A(n3101), .ZN(U3287) );
  NAND2_X1 U3917 ( .A1(n3103), .A2(n3104), .ZN(n3144) );
  XNOR2_X1 U3918 ( .A(n3144), .B(n3143), .ZN(n3110) );
  NAND2_X1 U3919 ( .A1(n3640), .A2(n3838), .ZN(n3106) );
  OAI211_X1 U3920 ( .C1(n3178), .C2(n3642), .A(n3106), .B(n3105), .ZN(n3108)
         );
  NOR2_X1 U3921 ( .A1(n3644), .A2(n3216), .ZN(n3107) );
  AOI211_X1 U3922 ( .C1(n3215), .C2(n3647), .A(n3108), .B(n3107), .ZN(n3109)
         );
  OAI21_X1 U3923 ( .B1(n3110), .B2(n3650), .A(n3109), .ZN(U3224) );
  INV_X1 U3924 ( .A(n3111), .ZN(n3113) );
  OAI21_X1 U3925 ( .B1(n3113), .B2(n4414), .A(n3112), .ZN(n3119) );
  OAI22_X1 U3926 ( .A1(n4159), .A2(n3117), .B1(n4433), .B2(n2952), .ZN(n3114)
         );
  AOI21_X1 U3927 ( .B1(n3119), .B2(n4433), .A(n3114), .ZN(n3115) );
  INV_X1 U3928 ( .A(n3115), .ZN(U3520) );
  INV_X1 U3929 ( .A(REG0_REG_2__SCAN_IN), .ZN(n3116) );
  OAI22_X1 U3930 ( .A1(n4197), .A2(n3117), .B1(n4419), .B2(n3116), .ZN(n3118)
         );
  AOI21_X1 U3931 ( .B1(n3119), .B2(n4419), .A(n3118), .ZN(n3120) );
  INV_X1 U3932 ( .A(n3120), .ZN(U3471) );
  NAND2_X1 U3933 ( .A1(n3103), .A2(n3609), .ZN(n3131) );
  AOI21_X1 U3934 ( .B1(n3121), .B2(n3123), .A(n3122), .ZN(n3130) );
  INV_X1 U3935 ( .A(n4589), .ZN(n3128) );
  NAND2_X1 U3936 ( .A1(n3647), .A2(n4372), .ZN(n3125) );
  AND2_X1 U3937 ( .A1(U3149), .A2(REG3_REG_4__SCAN_IN), .ZN(n4223) );
  AOI21_X1 U3938 ( .B1(n3630), .B2(n3837), .A(n4223), .ZN(n3124) );
  OAI211_X1 U3939 ( .C1(n3126), .C2(n3632), .A(n3125), .B(n3124), .ZN(n3127)
         );
  AOI21_X1 U3940 ( .B1(n3128), .B2(n3601), .A(n3127), .ZN(n3129) );
  OAI21_X1 U3941 ( .B1(n3131), .B2(n3130), .A(n3129), .ZN(U3227) );
  OAI21_X1 U3942 ( .B1(n3133), .B2(n3132), .A(n3121), .ZN(n3141) );
  NOR2_X1 U3943 ( .A1(n3644), .A2(REG3_REG_3__SCAN_IN), .ZN(n3140) );
  NAND2_X1 U3944 ( .A1(n3647), .A2(n3134), .ZN(n3137) );
  AOI21_X1 U3945 ( .B1(n3630), .B2(n3838), .A(n3135), .ZN(n3136) );
  OAI211_X1 U3946 ( .C1(n3138), .C2(n3632), .A(n3137), .B(n3136), .ZN(n3139)
         );
  AOI211_X1 U3947 ( .C1(n3141), .C2(n3609), .A(n3140), .B(n3139), .ZN(n3142)
         );
  INV_X1 U3948 ( .A(n3142), .ZN(U3215) );
  NAND2_X1 U3949 ( .A1(n3144), .A2(n3143), .ZN(n3146) );
  NAND2_X1 U3950 ( .A1(n3146), .A2(n3145), .ZN(n3150) );
  NOR2_X1 U3951 ( .A1(n3148), .A2(n3147), .ZN(n3149) );
  XNOR2_X1 U3952 ( .A(n3150), .B(n3149), .ZN(n3157) );
  INV_X1 U3953 ( .A(n3241), .ZN(n3155) );
  NAND2_X1 U3954 ( .A1(n3647), .A2(n3232), .ZN(n3153) );
  AOI21_X1 U3955 ( .B1(n3630), .B2(n3835), .A(n3151), .ZN(n3152) );
  OAI211_X1 U3956 ( .C1(n2643), .C2(n3632), .A(n3153), .B(n3152), .ZN(n3154)
         );
  AOI21_X1 U3957 ( .B1(n3155), .B2(n3601), .A(n3154), .ZN(n3156) );
  OAI21_X1 U3958 ( .B1(n3157), .B2(n3650), .A(n3156), .ZN(U3236) );
  XOR2_X1 U3959 ( .A(n3160), .B(n3159), .Z(n3161) );
  XNOR2_X1 U3960 ( .A(n3158), .B(n3161), .ZN(n3167) );
  NAND2_X1 U3961 ( .A1(n3640), .A2(n3835), .ZN(n3163) );
  OAI211_X1 U3962 ( .C1(n3345), .C2(n3642), .A(n3163), .B(n3162), .ZN(n3165)
         );
  NOR2_X1 U3963 ( .A1(n3644), .A2(n3289), .ZN(n3164) );
  AOI211_X1 U3964 ( .C1(n3288), .C2(n3635), .A(n3165), .B(n3164), .ZN(n3166)
         );
  OAI21_X1 U3965 ( .B1(n3167), .B2(n3650), .A(n3166), .ZN(U3218) );
  AND2_X1 U3966 ( .A1(n3168), .A2(n3169), .ZN(n3171) );
  NAND2_X1 U3967 ( .A1(n3171), .A2(n3170), .ZN(n3173) );
  AOI21_X1 U3968 ( .B1(n3173), .B2(n3172), .A(n3650), .ZN(n3175) );
  NAND2_X1 U3969 ( .A1(n3175), .A2(n3174), .ZN(n3182) );
  NAND2_X1 U3970 ( .A1(n3630), .A2(n3834), .ZN(n3177) );
  OAI211_X1 U3971 ( .C1(n3178), .C2(n3632), .A(n3177), .B(n3176), .ZN(n3179)
         );
  AOI21_X1 U3972 ( .B1(n3180), .B2(n3647), .A(n3179), .ZN(n3181) );
  OAI211_X1 U3973 ( .C1(n3644), .C2(n3326), .A(n3182), .B(n3181), .ZN(U3210)
         );
  INV_X1 U3974 ( .A(n4207), .ZN(n3205) );
  INV_X1 U3975 ( .A(REG2_REG_9__SCAN_IN), .ZN(n3308) );
  INV_X1 U3976 ( .A(n3196), .ZN(n4356) );
  AOI22_X1 U3977 ( .A1(n3196), .A2(REG2_REG_9__SCAN_IN), .B1(n3308), .B2(n4356), .ZN(n4237) );
  OAI21_X1 U3978 ( .B1(n3308), .B2(n4356), .A(n4235), .ZN(n3184) );
  NAND2_X1 U3979 ( .A1(n4354), .A2(n3184), .ZN(n3185) );
  INV_X1 U3980 ( .A(REG2_REG_11__SCAN_IN), .ZN(n3186) );
  MUX2_X1 U3981 ( .A(n3186), .B(REG2_REG_11__SCAN_IN), .S(n4207), .Z(n3187) );
  INV_X1 U3982 ( .A(n3187), .ZN(n3188) );
  OAI211_X1 U3983 ( .C1(n3189), .C2(n3188), .A(n4316), .B(n3882), .ZN(n3204)
         );
  INV_X1 U3984 ( .A(REG3_REG_11__SCAN_IN), .ZN(n3190) );
  NOR2_X1 U3985 ( .A1(STATE_REG_SCAN_IN), .A2(n3190), .ZN(n3272) );
  INV_X1 U3986 ( .A(n3191), .ZN(n3193) );
  NAND2_X1 U3987 ( .A1(n3193), .A2(n2077), .ZN(n3194) );
  INV_X1 U3988 ( .A(REG1_REG_9__SCAN_IN), .ZN(n4429) );
  AOI22_X1 U3989 ( .A1(n3196), .A2(n4429), .B1(REG1_REG_9__SCAN_IN), .B2(n4356), .ZN(n4231) );
  NOR2_X1 U3990 ( .A1(n3197), .A2(n4249), .ZN(n3198) );
  INV_X1 U3991 ( .A(REG1_REG_10__SCAN_IN), .ZN(n4242) );
  INV_X1 U3992 ( .A(REG1_REG_11__SCAN_IN), .ZN(n3199) );
  MUX2_X1 U3993 ( .A(n3199), .B(REG1_REG_11__SCAN_IN), .S(n4207), .Z(n3200) );
  AOI211_X1 U3994 ( .C1(n3201), .C2(n3200), .A(n3869), .B(n4321), .ZN(n3202)
         );
  AOI211_X1 U3995 ( .C1(n4320), .C2(ADDR_REG_11__SCAN_IN), .A(n3272), .B(n3202), .ZN(n3203) );
  OAI211_X1 U3996 ( .C1(n4319), .C2(n3205), .A(n3204), .B(n3203), .ZN(U3251)
         );
  OR2_X1 U3997 ( .A1(n3035), .A2(n4380), .ZN(n3206) );
  NAND2_X1 U3998 ( .A1(n3445), .A2(n3206), .ZN(n3397) );
  INV_X1 U3999 ( .A(n3208), .ZN(n3711) );
  NAND2_X1 U4000 ( .A1(n3711), .A2(n3726), .ZN(n3788) );
  XNOR2_X1 U4001 ( .A(n3207), .B(n3788), .ZN(n4390) );
  XNOR2_X1 U4002 ( .A(n3209), .B(n3788), .ZN(n3213) );
  AOI22_X1 U4003 ( .A1(n3836), .A2(n4089), .B1(n4112), .B2(n3215), .ZN(n3210)
         );
  OAI21_X1 U4004 ( .B1(n3211), .B2(n4093), .A(n3210), .ZN(n3212) );
  AOI21_X1 U4005 ( .B1(n3213), .B2(n4086), .A(n3212), .ZN(n4391) );
  MUX2_X1 U4006 ( .A(n2971), .B(n4391), .S(n4595), .Z(n3219) );
  AOI21_X1 U4007 ( .B1(n3215), .B2(n3214), .A(n3239), .ZN(n4394) );
  INV_X1 U4008 ( .A(n3216), .ZN(n3217) );
  AOI22_X1 U4009 ( .A1(n4394), .A2(n4213), .B1(n3217), .B2(n4098), .ZN(n3218)
         );
  OAI211_X1 U4010 ( .C1(n4104), .C2(n4390), .A(n3219), .B(n3218), .ZN(U3285)
         );
  INV_X1 U4011 ( .A(n3220), .ZN(n3221) );
  AOI21_X1 U4012 ( .B1(n3223), .B2(n3222), .A(n3221), .ZN(n3229) );
  INV_X1 U4013 ( .A(n3307), .ZN(n3227) );
  NAND2_X1 U4014 ( .A1(n3647), .A2(n3312), .ZN(n3225) );
  AND2_X1 U4015 ( .A1(U3149), .A2(REG3_REG_9__SCAN_IN), .ZN(n4234) );
  AOI21_X1 U4016 ( .B1(n3630), .B2(n3832), .A(n4234), .ZN(n3224) );
  OAI211_X1 U4017 ( .C1(n3319), .C2(n3632), .A(n3225), .B(n3224), .ZN(n3226)
         );
  AOI21_X1 U4018 ( .B1(n3227), .B2(n3601), .A(n3226), .ZN(n3228) );
  OAI21_X1 U4019 ( .B1(n3229), .B2(n3650), .A(n3228), .ZN(U3228) );
  INV_X1 U4020 ( .A(n3712), .ZN(n3727) );
  NOR2_X1 U4021 ( .A1(n3715), .A2(n3727), .ZN(n3794) );
  XOR2_X1 U4022 ( .A(n3230), .B(n3794), .Z(n3237) );
  XNOR2_X1 U4023 ( .A(n3231), .B(n3794), .ZN(n3235) );
  AOI22_X1 U4024 ( .A1(n3835), .A2(n4089), .B1(n4112), .B2(n3232), .ZN(n3233)
         );
  OAI21_X1 U4025 ( .B1(n2643), .B2(n4093), .A(n3233), .ZN(n3234) );
  AOI21_X1 U4026 ( .B1(n3235), .B2(n4086), .A(n3234), .ZN(n3236) );
  OAI21_X1 U4027 ( .B1(n3237), .B2(n4380), .A(n3236), .ZN(n4396) );
  INV_X1 U4028 ( .A(n4396), .ZN(n3246) );
  INV_X1 U4029 ( .A(n3237), .ZN(n4399) );
  NOR2_X1 U4030 ( .A1(n3239), .A2(n3238), .ZN(n4395) );
  NOR3_X1 U4031 ( .A1(n4395), .A2(n3240), .A3(n4101), .ZN(n3244) );
  INV_X1 U4032 ( .A(REG2_REG_6__SCAN_IN), .ZN(n3242) );
  OAI22_X1 U4033 ( .A1(n4595), .A2(n3242), .B1(n3241), .B2(n4590), .ZN(n3243)
         );
  AOI211_X1 U4034 ( .C1(n4399), .C2(n3425), .A(n3244), .B(n3243), .ZN(n3245)
         );
  OAI21_X1 U4035 ( .B1(n3246), .B2(n3035), .A(n3245), .ZN(U3284) );
  NAND2_X1 U4036 ( .A1(n3247), .A2(n3609), .ZN(n3257) );
  AOI21_X1 U4037 ( .B1(n3220), .B2(n3249), .A(n3248), .ZN(n3256) );
  INV_X1 U4038 ( .A(n3250), .ZN(n3349) );
  NAND2_X1 U4039 ( .A1(n3647), .A2(n3342), .ZN(n3253) );
  NOR2_X1 U4040 ( .A1(STATE_REG_SCAN_IN), .A2(n3251), .ZN(n4243) );
  AOI21_X1 U4041 ( .B1(n3630), .B2(n3831), .A(n4243), .ZN(n3252) );
  OAI211_X1 U4042 ( .C1(n3345), .C2(n3632), .A(n3253), .B(n3252), .ZN(n3254)
         );
  AOI21_X1 U40430 ( .B1(n3349), .B2(n3601), .A(n3254), .ZN(n3255) );
  OAI21_X1 U4044 ( .B1(n3257), .B2(n3256), .A(n3255), .ZN(U3214) );
  XOR2_X1 U4045 ( .A(n3259), .B(n3258), .Z(n3260) );
  XNOR2_X1 U4046 ( .A(n3261), .B(n3260), .ZN(n3266) );
  NAND2_X1 U4047 ( .A1(n3640), .A2(n3831), .ZN(n3262) );
  NAND2_X1 U4048 ( .A1(REG3_REG_12__SCAN_IN), .A2(U3149), .ZN(n4253) );
  OAI211_X1 U4049 ( .C1(n3432), .C2(n3642), .A(n3262), .B(n4253), .ZN(n3264)
         );
  NOR2_X1 U4050 ( .A1(n3644), .A2(n3393), .ZN(n3263) );
  AOI211_X1 U4051 ( .C1(n3385), .C2(n3647), .A(n3264), .B(n3263), .ZN(n3265)
         );
  OAI21_X1 U4052 ( .B1(n3266), .B2(n3650), .A(n3265), .ZN(U3221) );
  NAND2_X1 U4053 ( .A1(n3268), .A2(n3267), .ZN(n3270) );
  XOR2_X1 U4054 ( .A(n3270), .B(n3269), .Z(n3279) );
  INV_X1 U4055 ( .A(n3376), .ZN(n3277) );
  NAND2_X1 U4056 ( .A1(n3647), .A2(n3271), .ZN(n3274) );
  AOI21_X1 U4057 ( .B1(n3630), .B2(n3830), .A(n3272), .ZN(n3273) );
  OAI211_X1 U4058 ( .C1(n3275), .C2(n3632), .A(n3274), .B(n3273), .ZN(n3276)
         );
  AOI21_X1 U4059 ( .B1(n3277), .B2(n3601), .A(n3276), .ZN(n3278) );
  OAI21_X1 U4060 ( .B1(n3279), .B2(n3650), .A(n3278), .ZN(U3233) );
  AND2_X1 U4061 ( .A1(n3719), .A2(n3729), .ZN(n3793) );
  XNOR2_X1 U4062 ( .A(n3280), .B(n3793), .ZN(n3296) );
  INV_X1 U4063 ( .A(n3296), .ZN(n3294) );
  CLKBUF_X1 U4064 ( .A(n3281), .Z(n3282) );
  XOR2_X1 U4065 ( .A(n3793), .B(n3282), .Z(n3283) );
  NAND2_X1 U4066 ( .A1(n3283), .A2(n4049), .ZN(n3285) );
  AOI22_X1 U4067 ( .A1(n3833), .A2(n4089), .B1(n4112), .B2(n3288), .ZN(n3284)
         );
  OAI211_X1 U4068 ( .C1(n3286), .C2(n4093), .A(n3285), .B(n3284), .ZN(n3295)
         );
  NAND2_X1 U4069 ( .A1(n3295), .A2(n4595), .ZN(n3293) );
  INV_X1 U4070 ( .A(n3306), .ZN(n3287) );
  AOI21_X1 U4071 ( .B1(n3288), .B2(n3317), .A(n3287), .ZN(n3302) );
  OAI22_X1 U4072 ( .A1(n4595), .A2(n3290), .B1(n3289), .B2(n4590), .ZN(n3291)
         );
  AOI21_X1 U4073 ( .B1(n3302), .B2(n4213), .A(n3291), .ZN(n3292) );
  OAI211_X1 U4074 ( .C1(n4104), .C2(n3294), .A(n3293), .B(n3292), .ZN(U3282)
         );
  AOI21_X1 U4075 ( .B1(n3296), .B2(n4400), .A(n3295), .ZN(n3304) );
  INV_X1 U4076 ( .A(n4197), .ZN(n3299) );
  INV_X1 U4077 ( .A(REG0_REG_8__SCAN_IN), .ZN(n3297) );
  NOR2_X1 U4078 ( .A1(n4419), .A2(n3297), .ZN(n3298) );
  AOI21_X1 U4079 ( .B1(n3302), .B2(n3299), .A(n3298), .ZN(n3300) );
  OAI21_X1 U4080 ( .B1(n3304), .B2(n4418), .A(n3300), .ZN(U3483) );
  INV_X1 U4081 ( .A(n4159), .ZN(n3301) );
  AOI22_X1 U4082 ( .A1(n3302), .A2(n3301), .B1(n4431), .B2(REG1_REG_8__SCAN_IN), .ZN(n3303) );
  OAI21_X1 U4083 ( .B1(n3304), .B2(n4431), .A(n3303), .ZN(U3526) );
  INV_X1 U4084 ( .A(n3723), .ZN(n3730) );
  NAND2_X1 U4085 ( .A1(n3730), .A2(n3720), .ZN(n3795) );
  XOR2_X1 U4086 ( .A(n3795), .B(n3305), .Z(n4407) );
  AOI21_X1 U4087 ( .B1(n3312), .B2(n3306), .A(n3348), .ZN(n4410) );
  OAI22_X1 U4088 ( .A1(n4595), .A2(n3308), .B1(n3307), .B2(n4590), .ZN(n3309)
         );
  AOI21_X1 U4089 ( .B1(n4410), .B2(n4213), .A(n3309), .ZN(n3316) );
  XNOR2_X1 U4090 ( .A(n3310), .B(n3795), .ZN(n3311) );
  NAND2_X1 U4091 ( .A1(n3311), .A2(n4049), .ZN(n3314) );
  AOI22_X1 U4092 ( .A1(n3832), .A2(n4089), .B1(n4112), .B2(n3312), .ZN(n3313)
         );
  OAI211_X1 U4093 ( .C1(n3319), .C2(n4093), .A(n3314), .B(n3313), .ZN(n4409)
         );
  NAND2_X1 U4094 ( .A1(n4409), .A2(n4595), .ZN(n3315) );
  OAI211_X1 U4095 ( .C1(n4407), .C2(n4104), .A(n3316), .B(n3315), .ZN(U3281)
         );
  OAI211_X1 U4096 ( .C1(n3240), .C2(n3318), .A(n4411), .B(n3317), .ZN(n4403)
         );
  OAI22_X1 U4097 ( .A1(n3319), .A2(n4379), .B1(n3318), .B2(n4377), .ZN(n3323)
         );
  XNOR2_X1 U4098 ( .A(n3320), .B(n3770), .ZN(n3321) );
  NOR2_X1 U4099 ( .A1(n3321), .A2(n4387), .ZN(n3322) );
  AOI211_X1 U4100 ( .C1(n4384), .C2(n3836), .A(n3323), .B(n3322), .ZN(n4404)
         );
  OAI21_X1 U4101 ( .B1(n4592), .B2(n4403), .A(n4404), .ZN(n3329) );
  NAND2_X1 U4102 ( .A1(n3325), .A2(n3770), .ZN(n4401) );
  AND3_X1 U4103 ( .A1(n3324), .A2(n3397), .A3(n4401), .ZN(n3328) );
  OAI22_X1 U4104 ( .A1(n4595), .A2(n4492), .B1(n3326), .B2(n4590), .ZN(n3327)
         );
  AOI211_X1 U4105 ( .C1(n3329), .C2(n4595), .A(n3328), .B(n3327), .ZN(n3330)
         );
  INV_X1 U4106 ( .A(n3330), .ZN(U3283) );
  NOR2_X1 U4107 ( .A1(n2050), .A2(n3331), .ZN(n3332) );
  XNOR2_X1 U4108 ( .A(n3333), .B(n3332), .ZN(n3339) );
  INV_X1 U4109 ( .A(n3334), .ZN(n3422) );
  NAND2_X1 U4110 ( .A1(n3647), .A2(n3411), .ZN(n3336) );
  AND2_X1 U4111 ( .A1(U3149), .A2(REG3_REG_13__SCAN_IN), .ZN(n4264) );
  AOI21_X1 U4112 ( .B1(n3630), .B2(n3828), .A(n4264), .ZN(n3335) );
  OAI211_X1 U4113 ( .C1(n3413), .C2(n3632), .A(n3336), .B(n3335), .ZN(n3337)
         );
  AOI21_X1 U4114 ( .B1(n3422), .B2(n3601), .A(n3337), .ZN(n3338) );
  OAI21_X1 U4115 ( .B1(n3339), .B2(n3650), .A(n3338), .ZN(U3231) );
  NAND2_X1 U4116 ( .A1(n3733), .A2(n3735), .ZN(n3786) );
  XOR2_X1 U4117 ( .A(n3340), .B(n3786), .Z(n3341) );
  NAND2_X1 U4118 ( .A1(n3341), .A2(n4086), .ZN(n3344) );
  AOI22_X1 U4119 ( .A1(n3831), .A2(n4089), .B1(n4112), .B2(n3342), .ZN(n3343)
         );
  OAI211_X1 U4120 ( .C1(n3345), .C2(n4093), .A(n3344), .B(n3343), .ZN(n3399)
         );
  INV_X1 U4121 ( .A(n3399), .ZN(n3353) );
  XNOR2_X1 U4122 ( .A(n3346), .B(n3786), .ZN(n3400) );
  INV_X1 U4123 ( .A(n3375), .ZN(n3347) );
  OAI21_X1 U4124 ( .B1(n3348), .B2(n2133), .A(n3347), .ZN(n3404) );
  AOI22_X1 U4125 ( .A1(n3035), .A2(REG2_REG_10__SCAN_IN), .B1(n3349), .B2(
        n4098), .ZN(n3350) );
  OAI21_X1 U4126 ( .B1(n3404), .B2(n4101), .A(n3350), .ZN(n3351) );
  AOI21_X1 U4127 ( .B1(n3400), .B2(n3397), .A(n3351), .ZN(n3352) );
  OAI21_X1 U4128 ( .B1(n3353), .B2(n3035), .A(n3352), .ZN(U3280) );
  XOR2_X1 U4129 ( .A(n3356), .B(n3355), .Z(n3357) );
  XNOR2_X1 U4130 ( .A(n3354), .B(n3357), .ZN(n3362) );
  NAND2_X1 U4131 ( .A1(n3630), .A2(n3827), .ZN(n3358) );
  NAND2_X1 U4132 ( .A1(REG3_REG_14__SCAN_IN), .A2(U3149), .ZN(n4281) );
  OAI211_X1 U4133 ( .C1(n3432), .C2(n3632), .A(n3358), .B(n4281), .ZN(n3360)
         );
  NOR2_X1 U4134 ( .A1(n3644), .A2(n3439), .ZN(n3359) );
  AOI211_X1 U4135 ( .C1(n3430), .C2(n3635), .A(n3360), .B(n3359), .ZN(n3361)
         );
  OAI21_X1 U4136 ( .B1(n3362), .B2(n3650), .A(n3361), .ZN(U3212) );
  OR2_X1 U4137 ( .A1(n3346), .A2(n3363), .ZN(n3366) );
  NAND2_X1 U4138 ( .A1(n3366), .A2(n3364), .ZN(n3368) );
  AND2_X1 U4139 ( .A1(n3366), .A2(n3365), .ZN(n3367) );
  AOI21_X1 U4140 ( .B1(n3791), .B2(n3368), .A(n3367), .ZN(n4415) );
  OAI22_X1 U4141 ( .A1(n3413), .A2(n4379), .B1(n3374), .B2(n4377), .ZN(n3369)
         );
  AOI21_X1 U4142 ( .B1(n4384), .B2(n3832), .A(n3369), .ZN(n3373) );
  XNOR2_X1 U4143 ( .A(n3370), .B(n3791), .ZN(n3371) );
  NAND2_X1 U4144 ( .A1(n3371), .A2(n4049), .ZN(n3372) );
  OAI211_X1 U4145 ( .C1(n4415), .C2(n4380), .A(n3373), .B(n3372), .ZN(n4417)
         );
  NAND2_X1 U4146 ( .A1(n4417), .A2(n4595), .ZN(n3380) );
  OAI21_X1 U4147 ( .B1(n3375), .B2(n3374), .A(n3390), .ZN(n4412) );
  INV_X1 U4148 ( .A(n4412), .ZN(n3378) );
  OAI22_X1 U4149 ( .A1(n4595), .A2(n3186), .B1(n3376), .B2(n4590), .ZN(n3377)
         );
  AOI21_X1 U4150 ( .B1(n3378), .B2(n4213), .A(n3377), .ZN(n3379) );
  OAI211_X1 U4151 ( .C1(n4415), .C2(n3445), .A(n3380), .B(n3379), .ZN(U3279)
         );
  INV_X1 U4152 ( .A(n3381), .ZN(n3382) );
  OR2_X1 U4153 ( .A1(n3370), .A2(n3382), .ZN(n3384) );
  NAND2_X1 U4154 ( .A1(n3384), .A2(n3383), .ZN(n3409) );
  NAND2_X1 U4155 ( .A1(n3408), .A2(n3406), .ZN(n3787) );
  XNOR2_X1 U4156 ( .A(n3409), .B(n3787), .ZN(n3389) );
  NAND2_X1 U4157 ( .A1(n3831), .A2(n4384), .ZN(n3387) );
  NAND2_X1 U4158 ( .A1(n3385), .A2(n4112), .ZN(n3386) );
  OAI211_X1 U4159 ( .C1(n3432), .C2(n4379), .A(n3387), .B(n3386), .ZN(n3388)
         );
  AOI21_X1 U4160 ( .B1(n3389), .B2(n4086), .A(n3388), .ZN(n3449) );
  XNOR2_X1 U4161 ( .A(n2021), .B(n3787), .ZN(n3447) );
  INV_X1 U4162 ( .A(n3390), .ZN(n3392) );
  OAI21_X1 U4163 ( .B1(n3392), .B2(n3391), .A(n3418), .ZN(n3454) );
  NOR2_X1 U4164 ( .A1(n3454), .A2(n4101), .ZN(n3396) );
  INV_X1 U4165 ( .A(REG2_REG_12__SCAN_IN), .ZN(n3394) );
  OAI22_X1 U4166 ( .A1(n4595), .A2(n3394), .B1(n3393), .B2(n4590), .ZN(n3395)
         );
  AOI211_X1 U4167 ( .C1(n3447), .C2(n3397), .A(n3396), .B(n3395), .ZN(n3398)
         );
  OAI21_X1 U4168 ( .B1(n3035), .B2(n3449), .A(n3398), .ZN(U3278) );
  INV_X1 U4169 ( .A(REG0_REG_10__SCAN_IN), .ZN(n4510) );
  AOI21_X1 U4170 ( .B1(n4400), .B2(n3400), .A(n3399), .ZN(n3402) );
  MUX2_X1 U4171 ( .A(n4510), .B(n3402), .S(n4419), .Z(n3401) );
  OAI21_X1 U4172 ( .B1(n3404), .B2(n4197), .A(n3401), .ZN(U3487) );
  MUX2_X1 U4173 ( .A(n4242), .B(n3402), .S(n4433), .Z(n3403) );
  OAI21_X1 U4174 ( .B1(n3404), .B2(n4159), .A(n3403), .ZN(U3528) );
  XNOR2_X1 U4175 ( .A(n3432), .B(n3411), .ZN(n3806) );
  XOR2_X1 U4176 ( .A(n3806), .B(n3405), .Z(n3417) );
  INV_X1 U4177 ( .A(n3406), .ZN(n3407) );
  AOI21_X1 U4178 ( .B1(n3409), .B2(n3408), .A(n3407), .ZN(n3410) );
  XOR2_X1 U4179 ( .A(n3806), .B(n3410), .Z(n3415) );
  AOI22_X1 U4180 ( .A1(n3828), .A2(n4089), .B1(n4112), .B2(n3411), .ZN(n3412)
         );
  OAI21_X1 U4181 ( .B1(n3413), .B2(n4093), .A(n3412), .ZN(n3414) );
  AOI21_X1 U4182 ( .B1(n3415), .B2(n4049), .A(n3414), .ZN(n3416) );
  OAI21_X1 U4183 ( .B1(n3417), .B2(n4380), .A(n3416), .ZN(n3497) );
  INV_X1 U4184 ( .A(n3497), .ZN(n3427) );
  INV_X1 U4185 ( .A(n3417), .ZN(n3498) );
  INV_X1 U4186 ( .A(n3418), .ZN(n3421) );
  OAI21_X1 U4187 ( .B1(n3421), .B2(n3420), .A(n3436), .ZN(n3502) );
  AOI22_X1 U4188 ( .A1(n3035), .A2(REG2_REG_13__SCAN_IN), .B1(n3422), .B2(
        n4098), .ZN(n3423) );
  OAI21_X1 U4189 ( .B1(n3502), .B2(n4101), .A(n3423), .ZN(n3424) );
  AOI21_X1 U4190 ( .B1(n3498), .B2(n3425), .A(n3424), .ZN(n3426) );
  OAI21_X1 U4191 ( .B1(n3427), .B2(n3035), .A(n3426), .ZN(U3277) );
  OAI21_X1 U4192 ( .B1(n2039), .B2(n3429), .A(n3428), .ZN(n3491) );
  INV_X1 U4193 ( .A(n3491), .ZN(n3446) );
  OAI21_X1 U4194 ( .B1(n3772), .B2(n3656), .A(n3456), .ZN(n3434) );
  AOI22_X1 U4195 ( .A1(n3827), .A2(n4089), .B1(n3430), .B2(n4112), .ZN(n3431)
         );
  OAI21_X1 U4196 ( .B1(n3432), .B2(n4093), .A(n3431), .ZN(n3433) );
  AOI21_X1 U4197 ( .B1(n3434), .B2(n4049), .A(n3433), .ZN(n3435) );
  OAI21_X1 U4198 ( .B1(n3446), .B2(n4380), .A(n3435), .ZN(n3490) );
  NAND2_X1 U4199 ( .A1(n3490), .A2(n4595), .ZN(n3444) );
  INV_X1 U4200 ( .A(n3437), .ZN(n3438) );
  OAI21_X1 U4201 ( .B1(n3419), .B2(n2408), .A(n3438), .ZN(n3496) );
  INV_X1 U4202 ( .A(n3496), .ZN(n3442) );
  INV_X1 U4203 ( .A(REG2_REG_14__SCAN_IN), .ZN(n3440) );
  OAI22_X1 U4204 ( .A1(n4595), .A2(n3440), .B1(n3439), .B2(n4590), .ZN(n3441)
         );
  AOI21_X1 U4205 ( .B1(n3442), .B2(n4213), .A(n3441), .ZN(n3443) );
  OAI211_X1 U4206 ( .C1(n3446), .C2(n3445), .A(n3444), .B(n3443), .ZN(U3276)
         );
  NAND2_X1 U4207 ( .A1(n3447), .A2(n4400), .ZN(n3448) );
  AND2_X1 U4208 ( .A1(n3449), .A2(n3448), .ZN(n3452) );
  INV_X1 U4209 ( .A(REG0_REG_12__SCAN_IN), .ZN(n3450) );
  MUX2_X1 U4210 ( .A(n3452), .B(n3450), .S(n4418), .Z(n3451) );
  OAI21_X1 U4211 ( .B1(n3454), .B2(n4197), .A(n3451), .ZN(U3491) );
  INV_X1 U4212 ( .A(REG1_REG_12__SCAN_IN), .ZN(n4252) );
  MUX2_X1 U4213 ( .A(n4252), .B(n3452), .S(n4433), .Z(n3453) );
  OAI21_X1 U4214 ( .B1(n3454), .B2(n4159), .A(n3453), .ZN(U3530) );
  XNOR2_X1 U4215 ( .A(n3455), .B(n3457), .ZN(n3485) );
  INV_X1 U4216 ( .A(n3485), .ZN(n3469) );
  NAND2_X1 U4217 ( .A1(n3456), .A2(n3652), .ZN(n3458) );
  INV_X1 U4218 ( .A(n3457), .ZN(n3773) );
  XNOR2_X1 U4219 ( .A(n3458), .B(n3773), .ZN(n3459) );
  NAND2_X1 U4220 ( .A1(n3459), .A2(n4086), .ZN(n3461) );
  AOI22_X1 U4221 ( .A1(n3826), .A2(n4089), .B1(n4112), .B2(n3648), .ZN(n3460)
         );
  OAI211_X1 U4222 ( .C1(n3462), .C2(n4093), .A(n3461), .B(n3460), .ZN(n3484)
         );
  OAI21_X1 U4223 ( .B1(n3437), .B2(n3464), .A(n3463), .ZN(n3489) );
  NOR2_X1 U4224 ( .A1(n3489), .A2(n4101), .ZN(n3467) );
  INV_X1 U4225 ( .A(REG2_REG_15__SCAN_IN), .ZN(n3465) );
  OAI22_X1 U4226 ( .A1(n4595), .A2(n3465), .B1(n3643), .B2(n4590), .ZN(n3466)
         );
  AOI211_X1 U4227 ( .C1(n3484), .C2(n4595), .A(n3467), .B(n3466), .ZN(n3468)
         );
  OAI21_X1 U4228 ( .B1(n3469), .B2(n4104), .A(n3468), .ZN(U3275) );
  OAI21_X1 U4229 ( .B1(n3471), .B2(n3472), .A(n3470), .ZN(n4163) );
  XNOR2_X1 U4230 ( .A(n3473), .B(n3472), .ZN(n3477) );
  NAND2_X1 U4231 ( .A1(n3825), .A2(n4089), .ZN(n3475) );
  NAND2_X1 U4232 ( .A1(n3579), .A2(n4112), .ZN(n3474) );
  OAI211_X1 U4233 ( .C1(n3575), .C2(n4093), .A(n3475), .B(n3474), .ZN(n3476)
         );
  AOI21_X1 U4234 ( .B1(n3477), .B2(n4086), .A(n3476), .ZN(n4162) );
  NOR2_X1 U4235 ( .A1(n4590), .A2(n3576), .ZN(n3478) );
  AOI21_X1 U4236 ( .B1(n3035), .B2(REG2_REG_16__SCAN_IN), .A(n3478), .ZN(n3481) );
  NAND2_X1 U4237 ( .A1(n3463), .A2(n3579), .ZN(n4160) );
  NAND3_X1 U4238 ( .A1(n3479), .A2(n4213), .A3(n4160), .ZN(n3480) );
  OAI211_X1 U4239 ( .C1(n4162), .C2(n3035), .A(n3481), .B(n3480), .ZN(n3482)
         );
  INV_X1 U4240 ( .A(n3482), .ZN(n3483) );
  OAI21_X1 U4241 ( .B1(n4163), .B2(n4104), .A(n3483), .ZN(U3274) );
  INV_X1 U4242 ( .A(REG0_REG_15__SCAN_IN), .ZN(n4507) );
  AOI21_X1 U4243 ( .B1(n3485), .B2(n4400), .A(n3484), .ZN(n3487) );
  MUX2_X1 U4244 ( .A(n4507), .B(n3487), .S(n4419), .Z(n3486) );
  OAI21_X1 U4245 ( .B1(n3489), .B2(n4197), .A(n3486), .ZN(U3497) );
  INV_X1 U4246 ( .A(REG1_REG_15__SCAN_IN), .ZN(n4494) );
  MUX2_X1 U4247 ( .A(n4494), .B(n3487), .S(n4433), .Z(n3488) );
  OAI21_X1 U4248 ( .B1(n4159), .B2(n3489), .A(n3488), .ZN(U3533) );
  INV_X1 U4249 ( .A(REG0_REG_14__SCAN_IN), .ZN(n3492) );
  INV_X1 U4250 ( .A(n4414), .ZN(n4398) );
  AOI21_X1 U4251 ( .B1(n4398), .B2(n3491), .A(n3490), .ZN(n3494) );
  MUX2_X1 U4252 ( .A(n3492), .B(n3494), .S(n4419), .Z(n3493) );
  OAI21_X1 U4253 ( .B1(n3496), .B2(n4197), .A(n3493), .ZN(U3495) );
  INV_X1 U4254 ( .A(REG1_REG_14__SCAN_IN), .ZN(n4275) );
  MUX2_X1 U4255 ( .A(n4275), .B(n3494), .S(n4433), .Z(n3495) );
  OAI21_X1 U4256 ( .B1(n4159), .B2(n3496), .A(n3495), .ZN(U3532) );
  INV_X1 U4257 ( .A(REG0_REG_13__SCAN_IN), .ZN(n4504) );
  AOI21_X1 U4258 ( .B1(n4398), .B2(n3498), .A(n3497), .ZN(n3500) );
  MUX2_X1 U4259 ( .A(n4504), .B(n3500), .S(n4419), .Z(n3499) );
  OAI21_X1 U4260 ( .B1(n3502), .B2(n4197), .A(n3499), .ZN(U3493) );
  INV_X1 U4261 ( .A(REG1_REG_13__SCAN_IN), .ZN(n3872) );
  MUX2_X1 U4262 ( .A(n3872), .B(n3500), .S(n4433), .Z(n3501) );
  OAI21_X1 U4263 ( .B1(n4159), .B2(n3502), .A(n3501), .ZN(U3531) );
  INV_X1 U4264 ( .A(IR_REG_30__SCAN_IN), .ZN(n3503) );
  NAND3_X1 U4265 ( .A1(n3503), .A2(IR_REG_31__SCAN_IN), .A3(STATE_REG_SCAN_IN), 
        .ZN(n3504) );
  INV_X1 U4266 ( .A(DATAI_31_), .ZN(n4558) );
  OAI22_X1 U4267 ( .A1(n3505), .A2(n3504), .B1(STATE_REG_SCAN_IN), .B2(n4558), 
        .ZN(U3321) );
  NAND2_X1 U4268 ( .A1(n3507), .A2(n3506), .ZN(n3508) );
  XOR2_X1 U4269 ( .A(n3804), .B(n3508), .Z(n4125) );
  XNOR2_X1 U4270 ( .A(n3509), .B(n3804), .ZN(n3513) );
  NAND2_X1 U4271 ( .A1(n3760), .A2(n4112), .ZN(n3511) );
  NAND2_X1 U4272 ( .A1(n3822), .A2(n4384), .ZN(n3510) );
  OAI211_X1 U4273 ( .C1(n3916), .C2(n4379), .A(n3511), .B(n3510), .ZN(n3512)
         );
  AOI21_X1 U4274 ( .B1(n3513), .B2(n4049), .A(n3512), .ZN(n4124) );
  AOI22_X1 U4275 ( .A1(n3035), .A2(REG2_REG_27__SCAN_IN), .B1(n3514), .B2(
        n4098), .ZN(n3518) );
  AND2_X1 U4276 ( .A1(n2027), .A2(n3760), .ZN(n3515) );
  NOR2_X1 U4277 ( .A1(n3516), .A2(n3515), .ZN(n4122) );
  NAND2_X1 U4278 ( .A1(n4122), .A2(n4213), .ZN(n3517) );
  OAI211_X1 U4279 ( .C1(n4124), .C2(n3035), .A(n3518), .B(n3517), .ZN(n3519)
         );
  INV_X1 U4280 ( .A(n3519), .ZN(n3520) );
  OAI21_X1 U4281 ( .B1(n4125), .B2(n4104), .A(n3520), .ZN(U3263) );
  INV_X1 U4282 ( .A(n3522), .ZN(n3528) );
  INV_X1 U4283 ( .A(n3523), .ZN(n3524) );
  AOI22_X1 U4284 ( .A1(n3524), .A2(n4098), .B1(n3035), .B2(
        REG2_REG_28__SCAN_IN), .ZN(n3525) );
  OAI21_X1 U4285 ( .B1(n3526), .B2(n4101), .A(n3525), .ZN(n3527) );
  AOI21_X1 U4286 ( .B1(n3528), .B2(n4595), .A(n3527), .ZN(n3529) );
  OAI21_X1 U4287 ( .B1(n3521), .B2(n4104), .A(n3529), .ZN(U3262) );
  INV_X1 U4288 ( .A(n3979), .ZN(n3538) );
  AND2_X1 U4289 ( .A1(n3616), .A2(n3530), .ZN(n3533) );
  OAI211_X1 U4290 ( .C1(n3533), .C2(n3532), .A(n3609), .B(n3531), .ZN(n3537)
         );
  AOI22_X1 U4291 ( .A1(n3630), .A2(n3972), .B1(REG3_REG_23__SCAN_IN), .B2(
        U3149), .ZN(n3534) );
  OAI21_X1 U4292 ( .B1(n4007), .B2(n3632), .A(n3534), .ZN(n3535) );
  AOI21_X1 U4293 ( .B1(n3971), .B2(n3647), .A(n3535), .ZN(n3536) );
  OAI211_X1 U4294 ( .C1(n3644), .C2(n3538), .A(n3537), .B(n3536), .ZN(U3213)
         );
  XOR2_X1 U4295 ( .A(n3540), .B(n3539), .Z(n3546) );
  NAND2_X1 U4296 ( .A1(n3640), .A2(n4090), .ZN(n3541) );
  NAND2_X1 U4297 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n3897) );
  OAI211_X1 U4298 ( .C1(n3552), .C2(n3642), .A(n3541), .B(n3897), .ZN(n3542)
         );
  AOI21_X1 U4299 ( .B1(n3543), .B2(n3647), .A(n3542), .ZN(n3545) );
  NAND2_X1 U4300 ( .A1(n3601), .A2(n4058), .ZN(n3544) );
  OAI211_X1 U4301 ( .C1(n3546), .C2(n3650), .A(n3545), .B(n3544), .ZN(U3216)
         );
  XNOR2_X1 U4302 ( .A(n3548), .B(n3547), .ZN(n3549) );
  XNOR2_X1 U4303 ( .A(n3550), .B(n3549), .ZN(n3556) );
  AOI22_X1 U4304 ( .A1(n3630), .A2(n3823), .B1(REG3_REG_21__SCAN_IN), .B2(
        U3149), .ZN(n3551) );
  OAI21_X1 U4305 ( .B1(n3552), .B2(n3632), .A(n3551), .ZN(n3554) );
  NOR2_X1 U4306 ( .A1(n3644), .A2(n4012), .ZN(n3553) );
  AOI211_X1 U4307 ( .C1(n4004), .C2(n3635), .A(n3554), .B(n3553), .ZN(n3555)
         );
  OAI21_X1 U4308 ( .B1(n3556), .B2(n3650), .A(n3555), .ZN(U3220) );
  NAND2_X1 U4309 ( .A1(n3558), .A2(n3557), .ZN(n3560) );
  XOR2_X1 U4310 ( .A(n3560), .B(n3559), .Z(n3568) );
  INV_X1 U4311 ( .A(n3561), .ZN(n3937) );
  NAND2_X1 U4312 ( .A1(n3635), .A2(n3562), .ZN(n3564) );
  AOI22_X1 U4313 ( .A1(n3630), .A2(n3822), .B1(REG3_REG_25__SCAN_IN), .B2(
        U3149), .ZN(n3563) );
  OAI211_X1 U4314 ( .C1(n3565), .C2(n3632), .A(n3564), .B(n3563), .ZN(n3566)
         );
  AOI21_X1 U4315 ( .B1(n3937), .B2(n3601), .A(n3566), .ZN(n3567) );
  OAI21_X1 U4316 ( .B1(n3568), .B2(n3650), .A(n3567), .ZN(U3222) );
  INV_X1 U4317 ( .A(n3569), .ZN(n3571) );
  OAI21_X1 U4318 ( .B1(n3571), .B2(n3639), .A(n3570), .ZN(n3572) );
  XOR2_X1 U4319 ( .A(n3573), .B(n3572), .Z(n3581) );
  NAND2_X1 U4320 ( .A1(n3630), .A2(n3825), .ZN(n3574) );
  NAND2_X1 U4321 ( .A1(REG3_REG_16__SCAN_IN), .A2(U3149), .ZN(n4294) );
  OAI211_X1 U4322 ( .C1(n3575), .C2(n3632), .A(n3574), .B(n4294), .ZN(n3578)
         );
  NOR2_X1 U4323 ( .A1(n3644), .A2(n3576), .ZN(n3577) );
  AOI211_X1 U4324 ( .C1(n3579), .C2(n3647), .A(n3578), .B(n3577), .ZN(n3580)
         );
  OAI21_X1 U4325 ( .B1(n3581), .B2(n3650), .A(n3580), .ZN(U3223) );
  XNOR2_X1 U4326 ( .A(n3584), .B(n3583), .ZN(n3585) );
  XNOR2_X1 U4327 ( .A(n3582), .B(n3585), .ZN(n3592) );
  INV_X1 U4328 ( .A(n3586), .ZN(n4099) );
  NAND2_X1 U4329 ( .A1(n3635), .A2(n4088), .ZN(n3589) );
  INV_X1 U4330 ( .A(REG3_REG_17__SCAN_IN), .ZN(n3587) );
  NOR2_X1 U4331 ( .A1(STATE_REG_SCAN_IN), .A2(n3587), .ZN(n4306) );
  AOI21_X1 U4332 ( .B1(n3630), .B2(n4090), .A(n4306), .ZN(n3588) );
  OAI211_X1 U4333 ( .C1(n4094), .C2(n3632), .A(n3589), .B(n3588), .ZN(n3590)
         );
  AOI21_X1 U4334 ( .B1(n4099), .B2(n3601), .A(n3590), .ZN(n3591) );
  OAI21_X1 U4335 ( .B1(n3592), .B2(n3650), .A(n3591), .ZN(U3225) );
  NAND2_X1 U4336 ( .A1(n3593), .A2(n3594), .ZN(n3595) );
  XOR2_X1 U4337 ( .A(n3596), .B(n3595), .Z(n3603) );
  INV_X1 U4338 ( .A(n3597), .ZN(n3956) );
  NAND2_X1 U4339 ( .A1(n3635), .A2(n3948), .ZN(n3599) );
  AOI22_X1 U4340 ( .A1(n3630), .A2(n3949), .B1(REG3_REG_24__SCAN_IN), .B2(
        U3149), .ZN(n3598) );
  OAI211_X1 U4341 ( .C1(n3952), .C2(n3632), .A(n3599), .B(n3598), .ZN(n3600)
         );
  AOI21_X1 U4342 ( .B1(n3956), .B2(n3601), .A(n3600), .ZN(n3602) );
  OAI21_X1 U4343 ( .B1(n3603), .B2(n3650), .A(n3602), .ZN(U3226) );
  INV_X1 U4344 ( .A(n3608), .ZN(n3604) );
  NOR2_X1 U4345 ( .A1(n3605), .A2(n3604), .ZN(n3611) );
  AOI21_X1 U4346 ( .B1(n3608), .B2(n3607), .A(n3606), .ZN(n3610) );
  OAI21_X1 U4347 ( .B1(n3611), .B2(n3610), .A(n3609), .ZN(n3615) );
  AOI22_X1 U4348 ( .A1(n3630), .A2(n3824), .B1(REG3_REG_20__SCAN_IN), .B2(
        U3149), .ZN(n3612) );
  OAI21_X1 U4349 ( .B1(n4033), .B2(n3632), .A(n3612), .ZN(n3613) );
  AOI21_X1 U4350 ( .B1(n3802), .B2(n3635), .A(n3613), .ZN(n3614) );
  OAI211_X1 U4351 ( .C1(n3644), .C2(n4037), .A(n3615), .B(n3614), .ZN(U3230)
         );
  INV_X1 U4352 ( .A(n3616), .ZN(n3617) );
  AOI21_X1 U4353 ( .B1(n3619), .B2(n3618), .A(n3617), .ZN(n3624) );
  AOI22_X1 U4354 ( .A1(n3630), .A2(n3989), .B1(REG3_REG_22__SCAN_IN), .B2(
        U3149), .ZN(n3620) );
  OAI21_X1 U4355 ( .B1(n4029), .B2(n3632), .A(n3620), .ZN(n3622) );
  NOR2_X1 U4356 ( .A1(n3644), .A2(n3994), .ZN(n3621) );
  AOI211_X1 U4357 ( .C1(n3996), .C2(n3635), .A(n3622), .B(n3621), .ZN(n3623)
         );
  OAI21_X1 U4358 ( .B1(n3624), .B2(n3650), .A(n3623), .ZN(U3232) );
  INV_X1 U4359 ( .A(n3625), .ZN(n3627) );
  NOR2_X1 U4360 ( .A1(n3627), .A2(n3626), .ZN(n3628) );
  XNOR2_X1 U4361 ( .A(n3629), .B(n3628), .ZN(n3637) );
  NAND2_X1 U4362 ( .A1(n3630), .A2(n4073), .ZN(n3631) );
  NAND2_X1 U4363 ( .A1(REG3_REG_18__SCAN_IN), .A2(U3149), .ZN(n4336) );
  OAI211_X1 U4364 ( .C1(n4075), .C2(n3632), .A(n3631), .B(n4336), .ZN(n3634)
         );
  NOR2_X1 U4365 ( .A1(n3644), .A2(n4078), .ZN(n3633) );
  AOI211_X1 U4366 ( .C1(n4072), .C2(n3635), .A(n3634), .B(n3633), .ZN(n3636)
         );
  OAI21_X1 U4367 ( .B1(n3637), .B2(n3650), .A(n3636), .ZN(U3235) );
  NAND2_X1 U4368 ( .A1(n3570), .A2(n3569), .ZN(n3638) );
  XOR2_X1 U4369 ( .A(n3639), .B(n3638), .Z(n3651) );
  NAND2_X1 U4370 ( .A1(n3640), .A2(n3828), .ZN(n3641) );
  NAND2_X1 U4371 ( .A1(REG3_REG_15__SCAN_IN), .A2(U3149), .ZN(n4291) );
  OAI211_X1 U4372 ( .C1(n4094), .C2(n3642), .A(n3641), .B(n4291), .ZN(n3646)
         );
  NOR2_X1 U4373 ( .A1(n3644), .A2(n3643), .ZN(n3645) );
  AOI211_X1 U4374 ( .C1(n3648), .C2(n3647), .A(n3646), .B(n3645), .ZN(n3649)
         );
  OAI21_X1 U4375 ( .B1(n3651), .B2(n3650), .A(n3649), .ZN(U3238) );
  NAND2_X1 U4376 ( .A1(n3652), .A2(n3655), .ZN(n3741) );
  NAND2_X1 U4377 ( .A1(n3654), .A2(n3653), .ZN(n3722) );
  NAND2_X1 U4378 ( .A1(n3722), .A2(n3655), .ZN(n3740) );
  OAI21_X1 U4379 ( .B1(n3656), .B2(n3741), .A(n3740), .ZN(n3657) );
  NAND2_X1 U4380 ( .A1(n3657), .A2(n3748), .ZN(n3658) );
  NAND4_X1 U4381 ( .A1(n3658), .A2(n4025), .A3(n3745), .A4(n4021), .ZN(n3661)
         );
  INV_X1 U4382 ( .A(n3750), .ZN(n3659) );
  AOI21_X1 U4383 ( .B1(n3661), .B2(n3660), .A(n3659), .ZN(n3663) );
  OAI21_X1 U4384 ( .B1(n3664), .B2(n3663), .A(n3662), .ZN(n3665) );
  NAND2_X1 U4385 ( .A1(n3665), .A2(n3756), .ZN(n3675) );
  INV_X1 U4386 ( .A(n3820), .ZN(n3666) );
  INV_X1 U4387 ( .A(n3920), .ZN(n3912) );
  NAND2_X1 U4388 ( .A1(n3666), .A2(n3912), .ZN(n3681) );
  NAND4_X1 U4389 ( .A1(n3765), .A2(n3681), .A3(n3677), .A4(n3678), .ZN(n3674)
         );
  NAND2_X1 U4390 ( .A1(n3667), .A2(REG1_REG_30__SCAN_IN), .ZN(n3671) );
  NAND2_X1 U4391 ( .A1(n2478), .A2(REG2_REG_30__SCAN_IN), .ZN(n3670) );
  NAND2_X1 U4392 ( .A1(n3668), .A2(REG0_REG_30__SCAN_IN), .ZN(n3669) );
  NAND3_X1 U4393 ( .A1(n3671), .A2(n3670), .A3(n3669), .ZN(n3914) );
  INV_X1 U4394 ( .A(n3914), .ZN(n3672) );
  AND2_X1 U4395 ( .A1(n3819), .A2(n3694), .ZN(n3769) );
  AOI21_X1 U4396 ( .B1(n4113), .B2(n3672), .A(n3769), .ZN(n3775) );
  INV_X1 U4397 ( .A(n3775), .ZN(n3673) );
  AOI211_X1 U4398 ( .C1(n3675), .C2(n3757), .A(n3674), .B(n3673), .ZN(n3687)
         );
  INV_X1 U4399 ( .A(n3804), .ZN(n3685) );
  NAND2_X1 U4400 ( .A1(n3820), .A2(n3920), .ZN(n3680) );
  NAND3_X1 U4401 ( .A1(n3680), .A2(n3908), .A3(n3676), .ZN(n3762) );
  INV_X1 U4402 ( .A(n3762), .ZN(n3684) );
  INV_X1 U4403 ( .A(n3677), .ZN(n3907) );
  INV_X1 U4404 ( .A(n3678), .ZN(n3679) );
  NOR2_X1 U4405 ( .A1(n3907), .A2(n3679), .ZN(n3683) );
  NAND2_X1 U4406 ( .A1(n3680), .A2(n3908), .ZN(n3682) );
  OAI211_X1 U4407 ( .C1(n3683), .C2(n3682), .A(n3775), .B(n3681), .ZN(n3766)
         );
  AOI21_X1 U4408 ( .B1(n3685), .B2(n3684), .A(n3766), .ZN(n3686) );
  INV_X1 U4409 ( .A(n4113), .ZN(n3688) );
  OAI22_X1 U4410 ( .A1(n3687), .A2(n3686), .B1(n3819), .B2(n3688), .ZN(n3693)
         );
  AND2_X1 U4411 ( .A1(n3914), .A2(n3688), .ZN(n3695) );
  INV_X1 U4412 ( .A(n3819), .ZN(n3690) );
  OAI21_X1 U4413 ( .B1(n3695), .B2(n3690), .A(n3689), .ZN(n3692) );
  AOI21_X1 U4414 ( .B1(n3693), .B2(n3692), .A(n3691), .ZN(n3813) );
  OR2_X1 U4415 ( .A1(n3819), .A2(n3694), .ZN(n3697) );
  INV_X1 U4416 ( .A(n3695), .ZN(n3696) );
  AND2_X1 U4417 ( .A1(n3697), .A2(n3696), .ZN(n3783) );
  INV_X1 U4418 ( .A(n3698), .ZN(n3700) );
  OAI211_X1 U4419 ( .C1(n3701), .C2(n3808), .A(n3700), .B(n3699), .ZN(n3704)
         );
  NAND3_X1 U4420 ( .A1(n3704), .A2(n3703), .A3(n3702), .ZN(n3707) );
  NAND3_X1 U4421 ( .A1(n3707), .A2(n3706), .A3(n3705), .ZN(n3710) );
  NAND3_X1 U4422 ( .A1(n3710), .A2(n3709), .A3(n3708), .ZN(n3714) );
  NAND4_X1 U4423 ( .A1(n3714), .A2(n3713), .A3(n3712), .A4(n3711), .ZN(n3717)
         );
  INV_X1 U4424 ( .A(n3715), .ZN(n3716) );
  NAND3_X1 U4425 ( .A1(n3717), .A2(n3770), .A3(n3716), .ZN(n3718) );
  NAND3_X1 U4426 ( .A1(n3718), .A2(n3725), .A3(n3729), .ZN(n3721) );
  AND3_X1 U4427 ( .A1(n3721), .A2(n3720), .A3(n3719), .ZN(n3724) );
  NOR3_X1 U4428 ( .A1(n3724), .A2(n3723), .A3(n3722), .ZN(n3738) );
  INV_X1 U4429 ( .A(n3725), .ZN(n3728) );
  NOR3_X1 U4430 ( .A1(n3728), .A2(n3727), .A3(n3726), .ZN(n3731) );
  NAND3_X1 U4431 ( .A1(n3731), .A2(n3730), .A3(n3729), .ZN(n3734) );
  INV_X1 U4432 ( .A(n3740), .ZN(n3732) );
  AOI21_X1 U4433 ( .B1(n3734), .B2(n3733), .A(n3732), .ZN(n3737) );
  OAI211_X1 U4434 ( .C1(n3738), .C2(n3737), .A(n3736), .B(n3735), .ZN(n3744)
         );
  INV_X1 U4435 ( .A(n3739), .ZN(n3742) );
  OAI21_X1 U4436 ( .B1(n3742), .B2(n3741), .A(n3740), .ZN(n3743) );
  NAND2_X1 U4437 ( .A1(n3744), .A2(n3743), .ZN(n3746) );
  NAND2_X1 U4438 ( .A1(n3746), .A2(n3745), .ZN(n3749) );
  AOI21_X1 U4439 ( .B1(n3749), .B2(n3748), .A(n3747), .ZN(n3752) );
  OAI211_X1 U4440 ( .C1(n3752), .C2(n3751), .A(n3750), .B(n3963), .ZN(n3754)
         );
  AOI21_X1 U4441 ( .B1(n3755), .B2(n3754), .A(n3753), .ZN(n3759) );
  INV_X1 U4442 ( .A(n3756), .ZN(n3758) );
  OAI21_X1 U4443 ( .B1(n3759), .B2(n3758), .A(n3757), .ZN(n3764) );
  NOR2_X1 U4444 ( .A1(n3761), .A2(n3760), .ZN(n3763) );
  AOI211_X1 U4445 ( .C1(n3765), .C2(n3764), .A(n3763), .B(n3762), .ZN(n3767)
         );
  OR2_X1 U4446 ( .A1(n3767), .A2(n3766), .ZN(n3768) );
  OAI21_X1 U4447 ( .B1(n3769), .B2(n3783), .A(n3768), .ZN(n3811) );
  INV_X1 U4448 ( .A(n3985), .ZN(n3987) );
  NAND4_X1 U4449 ( .A1(n3987), .A2(n3772), .A3(n3771), .A4(n3770), .ZN(n3778)
         );
  NAND4_X1 U4450 ( .A1(n3776), .A2(n3775), .A3(n3774), .A4(n3773), .ZN(n3777)
         );
  XNOR2_X1 U4451 ( .A(n3820), .B(n3920), .ZN(n3910) );
  XNOR2_X1 U4452 ( .A(n3989), .B(n3971), .ZN(n3962) );
  INV_X1 U4453 ( .A(n3962), .ZN(n3968) );
  NOR4_X1 U4454 ( .A1(n3778), .A2(n3777), .A3(n3910), .A4(n3968), .ZN(n3801)
         );
  NAND2_X1 U4455 ( .A1(n3780), .A2(n3779), .ZN(n3946) );
  NAND2_X1 U4456 ( .A1(n3782), .A2(n3781), .ZN(n4047) );
  INV_X1 U4457 ( .A(n3783), .ZN(n3784) );
  NOR4_X1 U4458 ( .A1(n3946), .A2(n3785), .A3(n4047), .A4(n3784), .ZN(n3800)
         );
  NOR4_X1 U4459 ( .A1(n4071), .A2(n3788), .A3(n3787), .A4(n3786), .ZN(n3799)
         );
  INV_X1 U4460 ( .A(n4375), .ZN(n3790) );
  NAND4_X1 U4461 ( .A1(n3792), .A2(n3791), .A3(n3790), .A4(n3789), .ZN(n3797)
         );
  NAND2_X1 U4462 ( .A1(n3794), .A2(n3793), .ZN(n3796) );
  NAND2_X1 U4463 ( .A1(n4021), .A2(n4022), .ZN(n4084) );
  NOR4_X1 U4464 ( .A1(n3797), .A2(n3796), .A3(n4084), .A4(n3795), .ZN(n3798)
         );
  NAND4_X1 U4465 ( .A1(n3801), .A2(n3800), .A3(n3799), .A4(n3798), .ZN(n3807)
         );
  XNOR2_X1 U4466 ( .A(n4052), .B(n3802), .ZN(n4018) );
  INV_X1 U4467 ( .A(n4018), .ZN(n4026) );
  NAND2_X1 U4468 ( .A1(n3963), .A2(n3965), .ZN(n4002) );
  OR4_X1 U4469 ( .A1(n3905), .A2(n3804), .A3(n3803), .A4(n4002), .ZN(n3805) );
  NOR4_X1 U4470 ( .A1(n3807), .A2(n4026), .A3(n3806), .A4(n3805), .ZN(n3809)
         );
  NOR2_X1 U4471 ( .A1(n3809), .A2(n3808), .ZN(n3810) );
  MUX2_X1 U4472 ( .A(n3811), .B(n3810), .S(n4206), .Z(n3812) );
  NOR2_X1 U4473 ( .A1(n3813), .A2(n3812), .ZN(n3814) );
  XNOR2_X1 U4474 ( .A(n3814), .B(n4592), .ZN(n3818) );
  NAND2_X1 U4475 ( .A1(n3855), .A2(n2131), .ZN(n3815) );
  OAI211_X1 U4476 ( .C1(n4205), .C2(n3817), .A(n3815), .B(B_REG_SCAN_IN), .ZN(
        n3816) );
  OAI21_X1 U4477 ( .B1(n3818), .B2(n3817), .A(n3816), .ZN(U3239) );
  INV_X2 U4478 ( .A(U4043), .ZN(n3853) );
  MUX2_X1 U4479 ( .A(n3819), .B(DATAO_REG_31__SCAN_IN), .S(n3853), .Z(U3581)
         );
  MUX2_X1 U4480 ( .A(n3914), .B(DATAO_REG_30__SCAN_IN), .S(n3853), .Z(U3580)
         );
  MUX2_X1 U4481 ( .A(n3820), .B(DATAO_REG_29__SCAN_IN), .S(n3853), .Z(U3579)
         );
  MUX2_X1 U4482 ( .A(n3903), .B(DATAO_REG_28__SCAN_IN), .S(n3853), .Z(U3578)
         );
  MUX2_X1 U4483 ( .A(DATAO_REG_27__SCAN_IN), .B(n3821), .S(U4043), .Z(U3577)
         );
  MUX2_X1 U4484 ( .A(DATAO_REG_26__SCAN_IN), .B(n3822), .S(U4043), .Z(U3576)
         );
  MUX2_X1 U4485 ( .A(n3949), .B(DATAO_REG_25__SCAN_IN), .S(n3853), .Z(U3575)
         );
  MUX2_X1 U4486 ( .A(n3972), .B(DATAO_REG_24__SCAN_IN), .S(n3853), .Z(U3574)
         );
  MUX2_X1 U4487 ( .A(n3989), .B(DATAO_REG_23__SCAN_IN), .S(n3853), .Z(U3573)
         );
  MUX2_X1 U4488 ( .A(n3823), .B(DATAO_REG_22__SCAN_IN), .S(n3853), .Z(U3572)
         );
  MUX2_X1 U4489 ( .A(n3824), .B(DATAO_REG_21__SCAN_IN), .S(n3853), .Z(U3571)
         );
  MUX2_X1 U4490 ( .A(n4052), .B(DATAO_REG_20__SCAN_IN), .S(n3853), .Z(U3570)
         );
  MUX2_X1 U4491 ( .A(n4073), .B(DATAO_REG_19__SCAN_IN), .S(n3853), .Z(U3569)
         );
  MUX2_X1 U4492 ( .A(n4090), .B(DATAO_REG_18__SCAN_IN), .S(n3853), .Z(U3568)
         );
  MUX2_X1 U4493 ( .A(n3825), .B(DATAO_REG_17__SCAN_IN), .S(n3853), .Z(U3567)
         );
  MUX2_X1 U4494 ( .A(n3826), .B(DATAO_REG_16__SCAN_IN), .S(n3853), .Z(U3566)
         );
  MUX2_X1 U4495 ( .A(n3827), .B(DATAO_REG_15__SCAN_IN), .S(n3853), .Z(U3565)
         );
  MUX2_X1 U4496 ( .A(n3828), .B(DATAO_REG_14__SCAN_IN), .S(n3853), .Z(U3564)
         );
  MUX2_X1 U4497 ( .A(n3829), .B(DATAO_REG_13__SCAN_IN), .S(n3853), .Z(U3563)
         );
  MUX2_X1 U4498 ( .A(n3830), .B(DATAO_REG_12__SCAN_IN), .S(n3853), .Z(U3562)
         );
  MUX2_X1 U4499 ( .A(n3831), .B(DATAO_REG_11__SCAN_IN), .S(n3853), .Z(U3561)
         );
  MUX2_X1 U4500 ( .A(n3832), .B(DATAO_REG_10__SCAN_IN), .S(n3853), .Z(U3560)
         );
  MUX2_X1 U4501 ( .A(n3833), .B(DATAO_REG_9__SCAN_IN), .S(n3853), .Z(U3559) );
  MUX2_X1 U4502 ( .A(n3834), .B(DATAO_REG_8__SCAN_IN), .S(n3853), .Z(U3558) );
  MUX2_X1 U4503 ( .A(n3835), .B(DATAO_REG_7__SCAN_IN), .S(n3853), .Z(U3557) );
  MUX2_X1 U4504 ( .A(n3836), .B(DATAO_REG_6__SCAN_IN), .S(n3853), .Z(U3556) );
  MUX2_X1 U4505 ( .A(n3837), .B(DATAO_REG_5__SCAN_IN), .S(n3853), .Z(U3555) );
  MUX2_X1 U4506 ( .A(n3838), .B(DATAO_REG_4__SCAN_IN), .S(n3853), .Z(U3554) );
  MUX2_X1 U4507 ( .A(n4383), .B(DATAO_REG_3__SCAN_IN), .S(n3853), .Z(U3553) );
  MUX2_X1 U4508 ( .A(n3839), .B(DATAO_REG_2__SCAN_IN), .S(n3853), .Z(U3552) );
  MUX2_X1 U4509 ( .A(n3840), .B(DATAO_REG_1__SCAN_IN), .S(n3853), .Z(U3551) );
  MUX2_X1 U4510 ( .A(n3841), .B(DATAO_REG_0__SCAN_IN), .S(n3853), .Z(U3550) );
  OAI211_X1 U4511 ( .C1(n3844), .C2(n3843), .A(n4314), .B(n3842), .ZN(n3850)
         );
  OAI211_X1 U4512 ( .C1(n3846), .C2(n3854), .A(n4316), .B(n3845), .ZN(n3849)
         );
  AOI22_X1 U4513 ( .A1(n4320), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n3848) );
  NAND2_X1 U4514 ( .A1(n4332), .A2(n4212), .ZN(n3847) );
  NAND4_X1 U4515 ( .A1(n3850), .A2(n3849), .A3(n3848), .A4(n3847), .ZN(U3241)
         );
  NAND3_X1 U4516 ( .A1(n3852), .A2(n4201), .A3(n3851), .ZN(n3857) );
  AOI21_X1 U4517 ( .B1(n3855), .B2(n3854), .A(n3853), .ZN(n3856) );
  OAI211_X1 U4518 ( .C1(IR_REG_0__SCAN_IN), .C2(n3858), .A(n3857), .B(n3856), 
        .ZN(n4228) );
  AOI22_X1 U4519 ( .A1(ADDR_REG_2__SCAN_IN), .A2(n4320), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n3867) );
  XNOR2_X1 U4520 ( .A(n3860), .B(n3859), .ZN(n3861) );
  AOI22_X1 U4521 ( .A1(n4211), .A2(n4332), .B1(n4316), .B2(n3861), .ZN(n3866)
         );
  OAI211_X1 U4522 ( .C1(n3864), .C2(n3863), .A(n4314), .B(n3862), .ZN(n3865)
         );
  NAND4_X1 U4523 ( .A1(n4228), .A2(n3867), .A3(n3866), .A4(n3865), .ZN(U3242)
         );
  INV_X1 U4524 ( .A(REG1_REG_18__SCAN_IN), .ZN(n3868) );
  AOI22_X1 U4525 ( .A1(REG1_REG_18__SCAN_IN), .A2(n4342), .B1(n4331), .B2(
        n3868), .ZN(n4322) );
  INV_X1 U4526 ( .A(REG1_REG_17__SCAN_IN), .ZN(n4157) );
  INV_X1 U4527 ( .A(n3892), .ZN(n4344) );
  AOI22_X1 U4528 ( .A1(n3892), .A2(REG1_REG_17__SCAN_IN), .B1(n4157), .B2(
        n4344), .ZN(n4312) );
  INV_X1 U4529 ( .A(n4280), .ZN(n4350) );
  INV_X1 U4530 ( .A(n4272), .ZN(n4351) );
  NOR2_X1 U4531 ( .A1(n3870), .A2(n4353), .ZN(n3871) );
  AOI22_X1 U4532 ( .A1(REG1_REG_13__SCAN_IN), .A2(n4272), .B1(n4351), .B2(
        n3872), .ZN(n4261) );
  NOR2_X1 U4533 ( .A1(n4262), .A2(n4261), .ZN(n4260) );
  XNOR2_X1 U4534 ( .A(n4350), .B(n3873), .ZN(n4274) );
  INV_X1 U4535 ( .A(n4347), .ZN(n3889) );
  AOI22_X1 U4536 ( .A1(REG1_REG_15__SCAN_IN), .A2(n3889), .B1(n4347), .B2(
        n4494), .ZN(n4285) );
  NAND2_X1 U4537 ( .A1(n3876), .A2(n4346), .ZN(n3877) );
  INV_X1 U4538 ( .A(REG1_REG_16__SCAN_IN), .ZN(n4300) );
  NAND2_X1 U4539 ( .A1(n4301), .A2(n4300), .ZN(n4299) );
  XNOR2_X1 U4540 ( .A(n4592), .B(REG1_REG_19__SCAN_IN), .ZN(n3878) );
  XNOR2_X1 U4541 ( .A(n3879), .B(n3878), .ZN(n3902) );
  NAND2_X1 U4542 ( .A1(REG2_REG_18__SCAN_IN), .A2(n4331), .ZN(n3880) );
  OAI21_X1 U4543 ( .B1(REG2_REG_18__SCAN_IN), .B2(n4331), .A(n3880), .ZN(n4325) );
  NOR2_X1 U4544 ( .A1(n3892), .A2(REG2_REG_17__SCAN_IN), .ZN(n3881) );
  AOI21_X1 U4545 ( .B1(REG2_REG_17__SCAN_IN), .B2(n3892), .A(n3881), .ZN(n4309) );
  NAND2_X1 U4546 ( .A1(n4207), .A2(REG2_REG_11__SCAN_IN), .ZN(n3883) );
  NAND2_X1 U4547 ( .A1(REG2_REG_12__SCAN_IN), .A2(n4257), .ZN(n4256) );
  NAND2_X1 U4548 ( .A1(n3885), .A2(n3884), .ZN(n3886) );
  INV_X1 U4549 ( .A(REG2_REG_13__SCAN_IN), .ZN(n4266) );
  NOR2_X1 U4550 ( .A1(n4266), .A2(n4272), .ZN(n4265) );
  NOR2_X1 U4551 ( .A1(n4350), .A2(n3887), .ZN(n3888) );
  AOI22_X1 U4552 ( .A1(REG2_REG_15__SCAN_IN), .A2(n3889), .B1(n4347), .B2(
        n3465), .ZN(n4287) );
  NOR2_X1 U4553 ( .A1(n4288), .A2(n4287), .ZN(n4286) );
  NAND2_X1 U4554 ( .A1(n3890), .A2(n4346), .ZN(n3891) );
  INV_X1 U4555 ( .A(REG2_REG_16__SCAN_IN), .ZN(n4297) );
  NAND2_X1 U4556 ( .A1(n4309), .A2(n4308), .ZN(n4307) );
  OAI21_X1 U4557 ( .B1(n3892), .B2(REG2_REG_17__SCAN_IN), .A(n4307), .ZN(n4326) );
  NOR2_X1 U4558 ( .A1(n4325), .A2(n4326), .ZN(n4329) );
  AOI21_X1 U4559 ( .B1(n4331), .B2(REG2_REG_18__SCAN_IN), .A(n4329), .ZN(n3895) );
  INV_X1 U4560 ( .A(REG2_REG_19__SCAN_IN), .ZN(n3893) );
  MUX2_X1 U4561 ( .A(n3893), .B(REG2_REG_19__SCAN_IN), .S(n3898), .Z(n3894) );
  XNOR2_X1 U4562 ( .A(n3895), .B(n3894), .ZN(n3900) );
  NAND2_X1 U4563 ( .A1(n4320), .A2(ADDR_REG_19__SCAN_IN), .ZN(n3896) );
  OAI211_X1 U4564 ( .C1(n4319), .C2(n3898), .A(n3897), .B(n3896), .ZN(n3899)
         );
  AOI21_X1 U4565 ( .B1(n3900), .B2(n4316), .A(n3899), .ZN(n3901) );
  OAI21_X1 U4566 ( .B1(n3902), .B2(n4321), .A(n3901), .ZN(U3259) );
  INV_X1 U4567 ( .A(n4116), .ZN(n3927) );
  AOI21_X1 U4568 ( .B1(n3909), .B2(n3908), .A(n3907), .ZN(n3911) );
  XNOR2_X1 U4569 ( .A(n3911), .B(n3910), .ZN(n3918) );
  AOI22_X1 U4570 ( .A1(n3914), .A2(n3913), .B1(n3912), .B2(n4112), .ZN(n3915)
         );
  OAI21_X1 U4571 ( .B1(n3916), .B2(n4093), .A(n3915), .ZN(n3917) );
  AOI21_X2 U4572 ( .B1(n3918), .B2(n4049), .A(n3917), .ZN(n4118) );
  OAI21_X1 U4573 ( .B1(n3919), .B2(n4590), .A(n4118), .ZN(n3925) );
  OAI22_X1 U4574 ( .A1(n4117), .A2(n4101), .B1(n3923), .B2(n4595), .ZN(n3924)
         );
  AOI21_X1 U4575 ( .B1(n3925), .B2(n4595), .A(n3924), .ZN(n3926) );
  OAI21_X1 U4576 ( .B1(n3927), .B2(n4104), .A(n3926), .ZN(U3354) );
  INV_X1 U4577 ( .A(n3928), .ZN(n3933) );
  AOI22_X1 U4578 ( .A1(n3035), .A2(REG2_REG_26__SCAN_IN), .B1(n3929), .B2(
        n4098), .ZN(n3930) );
  OAI21_X1 U4579 ( .B1(n3931), .B2(n4101), .A(n3930), .ZN(n3932) );
  AOI21_X1 U4580 ( .B1(n3933), .B2(n4595), .A(n3932), .ZN(n3934) );
  OAI21_X1 U4581 ( .B1(n3935), .B2(n4104), .A(n3934), .ZN(U3264) );
  INV_X1 U4582 ( .A(n3936), .ZN(n3942) );
  AOI22_X1 U4583 ( .A1(n3035), .A2(REG2_REG_25__SCAN_IN), .B1(n3937), .B2(
        n4098), .ZN(n3938) );
  OAI21_X1 U4584 ( .B1(n4129), .B2(n4101), .A(n3938), .ZN(n3939) );
  AOI21_X1 U4585 ( .B1(n3940), .B2(n4595), .A(n3939), .ZN(n3941) );
  OAI21_X1 U4586 ( .B1(n3942), .B2(n4104), .A(n3941), .ZN(U3265) );
  XNOR2_X1 U4587 ( .A(n2842), .B(n3946), .ZN(n4131) );
  INV_X1 U4588 ( .A(n4131), .ZN(n3960) );
  NAND2_X1 U4589 ( .A1(n3944), .A2(n3943), .ZN(n3945) );
  XOR2_X1 U4590 ( .A(n3946), .B(n3945), .Z(n3947) );
  NAND2_X1 U4591 ( .A1(n3947), .A2(n4086), .ZN(n3951) );
  AOI22_X1 U4592 ( .A1(n3949), .A2(n4089), .B1(n4112), .B2(n3948), .ZN(n3950)
         );
  OAI211_X1 U4593 ( .C1(n3952), .C2(n4093), .A(n3951), .B(n3950), .ZN(n4130)
         );
  INV_X1 U4594 ( .A(n3953), .ZN(n3954) );
  OAI21_X1 U4595 ( .B1(n3976), .B2(n3955), .A(n3954), .ZN(n4175) );
  AOI22_X1 U4596 ( .A1(n3035), .A2(REG2_REG_24__SCAN_IN), .B1(n3956), .B2(
        n4098), .ZN(n3957) );
  OAI21_X1 U4597 ( .B1(n4175), .B2(n4101), .A(n3957), .ZN(n3958) );
  AOI21_X1 U4598 ( .B1(n4130), .B2(n4595), .A(n3958), .ZN(n3959) );
  OAI21_X1 U4599 ( .B1(n3960), .B2(n4104), .A(n3959), .ZN(U3266) );
  XNOR2_X1 U4600 ( .A(n3961), .B(n3962), .ZN(n4134) );
  INV_X1 U4601 ( .A(n4134), .ZN(n3983) );
  INV_X1 U4602 ( .A(n3963), .ZN(n3964) );
  OR2_X1 U4603 ( .A1(n4003), .A2(n3964), .ZN(n3966) );
  NAND2_X1 U4604 ( .A1(n3966), .A2(n3965), .ZN(n3988) );
  AOI21_X1 U4605 ( .B1(n3988), .B2(n3987), .A(n3967), .ZN(n3969) );
  XNOR2_X1 U4606 ( .A(n3969), .B(n3968), .ZN(n3970) );
  NAND2_X1 U4607 ( .A1(n3970), .A2(n4049), .ZN(n3974) );
  AOI22_X1 U4608 ( .A1(n3972), .A2(n4089), .B1(n4112), .B2(n3971), .ZN(n3973)
         );
  OAI211_X1 U4609 ( .C1(n4007), .C2(n4093), .A(n3974), .B(n3973), .ZN(n4133)
         );
  INV_X1 U4610 ( .A(n3976), .ZN(n3977) );
  OAI21_X1 U4611 ( .B1(n3975), .B2(n3978), .A(n3977), .ZN(n4179) );
  AOI22_X1 U4612 ( .A1(n3035), .A2(REG2_REG_23__SCAN_IN), .B1(n3979), .B2(
        n4098), .ZN(n3980) );
  OAI21_X1 U4613 ( .B1(n4179), .B2(n4101), .A(n3980), .ZN(n3981) );
  AOI21_X1 U4614 ( .B1(n4133), .B2(n4595), .A(n3981), .ZN(n3982) );
  OAI21_X1 U4615 ( .B1(n3983), .B2(n4104), .A(n3982), .ZN(U3267) );
  OAI21_X1 U4616 ( .B1(n3986), .B2(n3985), .A(n3984), .ZN(n4140) );
  XNOR2_X1 U4617 ( .A(n3988), .B(n3987), .ZN(n3993) );
  NAND2_X1 U4618 ( .A1(n3989), .A2(n4089), .ZN(n3991) );
  NAND2_X1 U4619 ( .A1(n3996), .A2(n4112), .ZN(n3990) );
  OAI211_X1 U4620 ( .C1(n4029), .C2(n4093), .A(n3991), .B(n3990), .ZN(n3992)
         );
  AOI21_X1 U4621 ( .B1(n3993), .B2(n4049), .A(n3992), .ZN(n4139) );
  NOR2_X1 U4622 ( .A1(n4590), .A2(n3994), .ZN(n3995) );
  AOI21_X1 U4623 ( .B1(n3035), .B2(REG2_REG_22__SCAN_IN), .A(n3995), .ZN(n3998) );
  INV_X1 U4624 ( .A(n3975), .ZN(n4137) );
  NAND2_X1 U4625 ( .A1(n2040), .A2(n3996), .ZN(n4136) );
  NAND3_X1 U4626 ( .A1(n4137), .A2(n4213), .A3(n4136), .ZN(n3997) );
  OAI211_X1 U4627 ( .C1(n4139), .C2(n3035), .A(n3998), .B(n3997), .ZN(n3999)
         );
  INV_X1 U4628 ( .A(n3999), .ZN(n4000) );
  OAI21_X1 U4629 ( .B1(n4140), .B2(n4104), .A(n4000), .ZN(U3268) );
  XOR2_X1 U4630 ( .A(n4002), .B(n4001), .Z(n4142) );
  XNOR2_X1 U4631 ( .A(n4003), .B(n4002), .ZN(n4009) );
  NAND2_X1 U4632 ( .A1(n4004), .A2(n4112), .ZN(n4006) );
  NAND2_X1 U4633 ( .A1(n4052), .A2(n4384), .ZN(n4005) );
  OAI211_X1 U4634 ( .C1(n4007), .C2(n4379), .A(n4006), .B(n4005), .ZN(n4008)
         );
  AOI21_X1 U4635 ( .B1(n4009), .B2(n4049), .A(n4008), .ZN(n4141) );
  INV_X1 U4636 ( .A(n4141), .ZN(n4016) );
  INV_X1 U4637 ( .A(n4034), .ZN(n4011) );
  OAI21_X1 U4638 ( .B1(n4011), .B2(n4010), .A(n2040), .ZN(n4184) );
  INV_X1 U4639 ( .A(n4012), .ZN(n4013) );
  AOI22_X1 U4640 ( .A1(n3035), .A2(REG2_REG_21__SCAN_IN), .B1(n4013), .B2(
        n4098), .ZN(n4014) );
  OAI21_X1 U4641 ( .B1(n4184), .B2(n4101), .A(n4014), .ZN(n4015) );
  AOI21_X1 U4642 ( .B1(n4016), .B2(n4595), .A(n4015), .ZN(n4017) );
  OAI21_X1 U4643 ( .B1(n4142), .B2(n4104), .A(n4017), .ZN(U3269) );
  XNOR2_X1 U4644 ( .A(n4019), .B(n4018), .ZN(n4146) );
  INV_X1 U4645 ( .A(n4146), .ZN(n4042) );
  INV_X1 U4646 ( .A(n4021), .ZN(n4023) );
  OAI21_X1 U4647 ( .B1(n4085), .B2(n4023), .A(n4022), .ZN(n4070) );
  AOI21_X1 U4648 ( .B1(n4070), .B2(n4025), .A(n4024), .ZN(n4027) );
  XNOR2_X1 U4649 ( .A(n4027), .B(n4026), .ZN(n4028) );
  NAND2_X1 U4650 ( .A1(n4028), .A2(n4086), .ZN(n4032) );
  OAI22_X1 U4651 ( .A1(n4029), .A2(n4379), .B1(n4377), .B2(n4035), .ZN(n4030)
         );
  INV_X1 U4652 ( .A(n4030), .ZN(n4031) );
  OAI211_X1 U4653 ( .C1(n4033), .C2(n4093), .A(n4032), .B(n4031), .ZN(n4145)
         );
  INV_X1 U4654 ( .A(n4056), .ZN(n4036) );
  OAI21_X1 U4655 ( .B1(n4036), .B2(n4035), .A(n4034), .ZN(n4188) );
  INV_X1 U4656 ( .A(n4037), .ZN(n4038) );
  AOI22_X1 U4657 ( .A1(n3035), .A2(REG2_REG_20__SCAN_IN), .B1(n4038), .B2(
        n4098), .ZN(n4039) );
  OAI21_X1 U4658 ( .B1(n4188), .B2(n4101), .A(n4039), .ZN(n4040) );
  AOI21_X1 U4659 ( .B1(n4145), .B2(n4595), .A(n4040), .ZN(n4041) );
  OAI21_X1 U4660 ( .B1(n4042), .B2(n4104), .A(n4041), .ZN(U3270) );
  XNOR2_X1 U4661 ( .A(n4043), .B(n4047), .ZN(n4150) );
  INV_X1 U4662 ( .A(n4150), .ZN(n4062) );
  INV_X1 U4663 ( .A(n4044), .ZN(n4046) );
  OAI21_X1 U4664 ( .B1(n4070), .B2(n4046), .A(n4045), .ZN(n4048) );
  XNOR2_X1 U4665 ( .A(n4048), .B(n4047), .ZN(n4050) );
  NAND2_X1 U4666 ( .A1(n4050), .A2(n4049), .ZN(n4054) );
  NOR2_X1 U4667 ( .A1(n4057), .A2(n4377), .ZN(n4051) );
  AOI21_X1 U4668 ( .B1(n4052), .B2(n4089), .A(n4051), .ZN(n4053) );
  OAI211_X1 U4669 ( .C1(n4055), .C2(n4093), .A(n4054), .B(n4053), .ZN(n4149)
         );
  OAI21_X1 U4670 ( .B1(n4067), .B2(n4057), .A(n4056), .ZN(n4192) );
  AOI22_X1 U4671 ( .A1(n3035), .A2(REG2_REG_19__SCAN_IN), .B1(n4058), .B2(
        n4098), .ZN(n4059) );
  OAI21_X1 U4672 ( .B1(n4192), .B2(n4101), .A(n4059), .ZN(n4060) );
  AOI21_X1 U4673 ( .B1(n4149), .B2(n4595), .A(n4060), .ZN(n4061) );
  OAI21_X1 U4674 ( .B1(n4062), .B2(n4104), .A(n4061), .ZN(U3271) );
  OAI21_X1 U4675 ( .B1(n4064), .B2(n4071), .A(n4063), .ZN(n4065) );
  INV_X1 U4676 ( .A(n4065), .ZN(n4154) );
  INV_X1 U4677 ( .A(n4067), .ZN(n4068) );
  OAI211_X1 U4678 ( .C1(n4066), .C2(n4069), .A(n4068), .B(n4411), .ZN(n4152)
         );
  XOR2_X1 U4679 ( .A(n4071), .B(n4070), .Z(n4077) );
  AOI22_X1 U4680 ( .A1(n4073), .A2(n4089), .B1(n4072), .B2(n4112), .ZN(n4074)
         );
  OAI21_X1 U4681 ( .B1(n4075), .B2(n4093), .A(n4074), .ZN(n4076) );
  AOI21_X1 U4682 ( .B1(n4077), .B2(n4086), .A(n4076), .ZN(n4153) );
  OAI21_X1 U4683 ( .B1(n4592), .B2(n4152), .A(n4153), .ZN(n4081) );
  INV_X1 U4684 ( .A(REG2_REG_18__SCAN_IN), .ZN(n4079) );
  OAI22_X1 U4685 ( .A1(n4595), .A2(n4079), .B1(n4078), .B2(n4590), .ZN(n4080)
         );
  AOI21_X1 U4686 ( .B1(n4081), .B2(n4595), .A(n4080), .ZN(n4082) );
  OAI21_X1 U4687 ( .B1(n4154), .B2(n4104), .A(n4082), .ZN(U3272) );
  XOR2_X1 U4688 ( .A(n4084), .B(n4083), .Z(n4156) );
  INV_X1 U4689 ( .A(n4156), .ZN(n4105) );
  XNOR2_X1 U4690 ( .A(n4085), .B(n4084), .ZN(n4087) );
  NAND2_X1 U4691 ( .A1(n4087), .A2(n4086), .ZN(n4092) );
  AOI22_X1 U4692 ( .A1(n4090), .A2(n4089), .B1(n4112), .B2(n4088), .ZN(n4091)
         );
  OAI211_X1 U4693 ( .C1(n4094), .C2(n4093), .A(n4092), .B(n4091), .ZN(n4155)
         );
  INV_X1 U4694 ( .A(n3479), .ZN(n4097) );
  INV_X1 U4695 ( .A(n4066), .ZN(n4095) );
  OAI21_X1 U4696 ( .B1(n4097), .B2(n4096), .A(n4095), .ZN(n4198) );
  AOI22_X1 U4697 ( .A1(n3035), .A2(REG2_REG_17__SCAN_IN), .B1(n4099), .B2(
        n4098), .ZN(n4100) );
  OAI21_X1 U4698 ( .B1(n4198), .B2(n4101), .A(n4100), .ZN(n4102) );
  AOI21_X1 U4699 ( .B1(n4155), .B2(n4595), .A(n4102), .ZN(n4103) );
  OAI21_X1 U4700 ( .B1(n4105), .B2(n4104), .A(n4103), .ZN(U3273) );
  INV_X1 U4701 ( .A(n4106), .ZN(n4166) );
  INV_X1 U4702 ( .A(REG1_REG_31__SCAN_IN), .ZN(n4107) );
  MUX2_X1 U4703 ( .A(n4107), .B(n4164), .S(n4433), .Z(n4108) );
  OAI21_X1 U4704 ( .B1(n4166), .B2(n4159), .A(n4108), .ZN(U3549) );
  AOI21_X1 U4705 ( .B1(n4113), .B2(n4110), .A(n4109), .ZN(n4214) );
  INV_X1 U4706 ( .A(n4214), .ZN(n4169) );
  INV_X1 U4707 ( .A(REG1_REG_30__SCAN_IN), .ZN(n4114) );
  AOI21_X1 U4708 ( .B1(n4113), .B2(n4112), .A(n4111), .ZN(n4216) );
  MUX2_X1 U4709 ( .A(n4114), .B(n4216), .S(n4433), .Z(n4115) );
  OAI21_X1 U4710 ( .B1(n4169), .B2(n4159), .A(n4115), .ZN(U3548) );
  NAND2_X1 U4711 ( .A1(n4116), .A2(n4400), .ZN(n4121) );
  NAND2_X1 U4712 ( .A1(n4121), .A2(n4120), .ZN(n4170) );
  MUX2_X1 U4713 ( .A(REG1_REG_29__SCAN_IN), .B(n4170), .S(n4433), .Z(U3547) );
  NAND2_X1 U4714 ( .A1(n4122), .A2(n4411), .ZN(n4123) );
  OAI211_X1 U4715 ( .C1(n4125), .C2(n4406), .A(n4124), .B(n4123), .ZN(n4171)
         );
  MUX2_X1 U4716 ( .A(REG1_REG_27__SCAN_IN), .B(n4171), .S(n4433), .Z(U3545) );
  INV_X1 U4717 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4127) );
  OAI21_X1 U4718 ( .B1(n4159), .B2(n4129), .A(n4128), .ZN(U3543) );
  INV_X1 U4719 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4546) );
  AOI21_X1 U4720 ( .B1(n4131), .B2(n4400), .A(n4130), .ZN(n4172) );
  MUX2_X1 U4721 ( .A(n4546), .B(n4172), .S(n4433), .Z(n4132) );
  OAI21_X1 U4722 ( .B1(n4159), .B2(n4175), .A(n4132), .ZN(U3542) );
  INV_X1 U4723 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4544) );
  AOI21_X1 U4724 ( .B1(n4134), .B2(n4400), .A(n4133), .ZN(n4176) );
  MUX2_X1 U4725 ( .A(n4544), .B(n4176), .S(n4433), .Z(n4135) );
  OAI21_X1 U4726 ( .B1(n4159), .B2(n4179), .A(n4135), .ZN(U3541) );
  NAND3_X1 U4727 ( .A1(n4137), .A2(n4411), .A3(n4136), .ZN(n4138) );
  OAI211_X1 U4728 ( .C1(n4140), .C2(n4406), .A(n4139), .B(n4138), .ZN(n4180)
         );
  MUX2_X1 U4729 ( .A(REG1_REG_22__SCAN_IN), .B(n4180), .S(n4433), .Z(U3540) );
  OAI21_X1 U4730 ( .B1(n4142), .B2(n4406), .A(n4141), .ZN(n4181) );
  MUX2_X1 U4731 ( .A(REG1_REG_21__SCAN_IN), .B(n4181), .S(n4433), .Z(n4143) );
  INV_X1 U4732 ( .A(n4143), .ZN(n4144) );
  OAI21_X1 U4733 ( .B1(n4159), .B2(n4184), .A(n4144), .ZN(U3539) );
  INV_X1 U4734 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4147) );
  AOI21_X1 U4735 ( .B1(n4146), .B2(n4400), .A(n4145), .ZN(n4185) );
  MUX2_X1 U4736 ( .A(n4147), .B(n4185), .S(n4433), .Z(n4148) );
  OAI21_X1 U4737 ( .B1(n4159), .B2(n4188), .A(n4148), .ZN(U3538) );
  INV_X1 U4738 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4466) );
  AOI21_X1 U4739 ( .B1(n4150), .B2(n4400), .A(n4149), .ZN(n4189) );
  MUX2_X1 U4740 ( .A(n4466), .B(n4189), .S(n4433), .Z(n4151) );
  OAI21_X1 U4741 ( .B1(n4159), .B2(n4192), .A(n4151), .ZN(U3537) );
  OAI211_X1 U4742 ( .C1(n4154), .C2(n4406), .A(n4153), .B(n4152), .ZN(n4193)
         );
  MUX2_X1 U4743 ( .A(REG1_REG_18__SCAN_IN), .B(n4193), .S(n4433), .Z(U3536) );
  AOI21_X1 U4744 ( .B1(n4156), .B2(n4400), .A(n4155), .ZN(n4194) );
  MUX2_X1 U4745 ( .A(n4157), .B(n4194), .S(n4433), .Z(n4158) );
  OAI21_X1 U4746 ( .B1(n4159), .B2(n4198), .A(n4158), .ZN(U3535) );
  NAND3_X1 U4747 ( .A1(n3479), .A2(n4411), .A3(n4160), .ZN(n4161) );
  OAI211_X1 U4748 ( .C1(n4163), .C2(n4406), .A(n4162), .B(n4161), .ZN(n4199)
         );
  MUX2_X1 U4749 ( .A(REG1_REG_16__SCAN_IN), .B(n4199), .S(n4433), .Z(U3534) );
  INV_X1 U4750 ( .A(REG0_REG_31__SCAN_IN), .ZN(n4524) );
  MUX2_X1 U4751 ( .A(n4524), .B(n4164), .S(n4419), .Z(n4165) );
  OAI21_X1 U4752 ( .B1(n4166), .B2(n4197), .A(n4165), .ZN(U3517) );
  INV_X1 U4753 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4167) );
  MUX2_X1 U4754 ( .A(n4167), .B(n4216), .S(n4419), .Z(n4168) );
  OAI21_X1 U4755 ( .B1(n4169), .B2(n4197), .A(n4168), .ZN(U3516) );
  MUX2_X1 U4756 ( .A(REG0_REG_29__SCAN_IN), .B(n4170), .S(n4419), .Z(U3515) );
  MUX2_X1 U4757 ( .A(REG0_REG_27__SCAN_IN), .B(n4171), .S(n4419), .Z(U3513) );
  INV_X1 U4758 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4173) );
  MUX2_X1 U4759 ( .A(n4173), .B(n4172), .S(n4419), .Z(n4174) );
  OAI21_X1 U4760 ( .B1(n4175), .B2(n4197), .A(n4174), .ZN(U3510) );
  INV_X1 U4761 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4177) );
  MUX2_X1 U4762 ( .A(n4177), .B(n4176), .S(n4419), .Z(n4178) );
  OAI21_X1 U4763 ( .B1(n4179), .B2(n4197), .A(n4178), .ZN(U3509) );
  MUX2_X1 U4764 ( .A(REG0_REG_22__SCAN_IN), .B(n4180), .S(n4419), .Z(U3508) );
  MUX2_X1 U4765 ( .A(REG0_REG_21__SCAN_IN), .B(n4181), .S(n4419), .Z(n4182) );
  INV_X1 U4766 ( .A(n4182), .ZN(n4183) );
  OAI21_X1 U4767 ( .B1(n4184), .B2(n4197), .A(n4183), .ZN(U3507) );
  INV_X1 U4768 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4186) );
  MUX2_X1 U4769 ( .A(n4186), .B(n4185), .S(n4419), .Z(n4187) );
  OAI21_X1 U4770 ( .B1(n4188), .B2(n4197), .A(n4187), .ZN(U3506) );
  INV_X1 U4771 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4190) );
  MUX2_X1 U4772 ( .A(n4190), .B(n4189), .S(n4419), .Z(n4191) );
  OAI21_X1 U4773 ( .B1(n4192), .B2(n4197), .A(n4191), .ZN(U3505) );
  MUX2_X1 U4774 ( .A(REG0_REG_18__SCAN_IN), .B(n4193), .S(n4419), .Z(U3503) );
  INV_X1 U4775 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4195) );
  MUX2_X1 U4776 ( .A(n4195), .B(n4194), .S(n4419), .Z(n4196) );
  OAI21_X1 U4777 ( .B1(n4198), .B2(n4197), .A(n4196), .ZN(U3501) );
  MUX2_X1 U4778 ( .A(REG0_REG_16__SCAN_IN), .B(n4199), .S(n4419), .Z(U3499) );
  MUX2_X1 U4779 ( .A(n4200), .B(DATAI_30_), .S(U3149), .Z(U3322) );
  MUX2_X1 U4780 ( .A(DATAI_28_), .B(n4201), .S(STATE_REG_SCAN_IN), .Z(U3324)
         );
  MUX2_X1 U4781 ( .A(n4202), .B(DATAI_26_), .S(U3149), .Z(U3326) );
  MUX2_X1 U4782 ( .A(n4203), .B(DATAI_25_), .S(U3149), .Z(U3327) );
  MUX2_X1 U4783 ( .A(n4204), .B(DATAI_24_), .S(U3149), .Z(U3328) );
  MUX2_X1 U4784 ( .A(n4205), .B(DATAI_22_), .S(U3149), .Z(U3330) );
  MUX2_X1 U4785 ( .A(DATAI_20_), .B(n4206), .S(STATE_REG_SCAN_IN), .Z(U3332)
         );
  MUX2_X1 U4786 ( .A(n4592), .B(DATAI_19_), .S(U3149), .Z(U3333) );
  MUX2_X1 U4787 ( .A(n4207), .B(DATAI_11_), .S(U3149), .Z(U3341) );
  MUX2_X1 U4788 ( .A(n4208), .B(DATAI_7_), .S(U3149), .Z(U3345) );
  MUX2_X1 U4789 ( .A(DATAI_6_), .B(n4209), .S(STATE_REG_SCAN_IN), .Z(U3346) );
  MUX2_X1 U4790 ( .A(n4210), .B(DATAI_5_), .S(U3149), .Z(U3347) );
  MUX2_X1 U4791 ( .A(DATAI_4_), .B(n4222), .S(STATE_REG_SCAN_IN), .Z(U3348) );
  MUX2_X1 U4792 ( .A(DATAI_2_), .B(n4211), .S(STATE_REG_SCAN_IN), .Z(U3350) );
  MUX2_X1 U4793 ( .A(n4212), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  AOI22_X1 U4794 ( .A1(n4214), .A2(n4213), .B1(REG2_REG_30__SCAN_IN), .B2(
        n3035), .ZN(n4215) );
  OAI21_X1 U4795 ( .B1(n3035), .B2(n4216), .A(n4215), .ZN(U3261) );
  XNOR2_X1 U4796 ( .A(n4217), .B(n2085), .ZN(n4218) );
  NAND2_X1 U4797 ( .A1(n4316), .A2(n4218), .ZN(n4227) );
  INV_X1 U4798 ( .A(REG1_REG_4__SCAN_IN), .ZN(n4219) );
  XNOR2_X1 U4799 ( .A(n4220), .B(n4219), .ZN(n4221) );
  NAND2_X1 U4800 ( .A1(n4314), .A2(n4221), .ZN(n4226) );
  NAND2_X1 U4801 ( .A1(n4332), .A2(n4222), .ZN(n4225) );
  AOI21_X1 U4802 ( .B1(n4320), .B2(ADDR_REG_4__SCAN_IN), .A(n4223), .ZN(n4224)
         );
  AND4_X1 U4803 ( .A1(n4227), .A2(n4226), .A3(n4225), .A4(n4224), .ZN(n4229)
         );
  NAND2_X1 U4804 ( .A1(n4229), .A2(n4228), .ZN(U3244) );
  AOI211_X1 U4805 ( .C1(n4232), .C2(n4231), .A(n4230), .B(n4321), .ZN(n4233)
         );
  AOI211_X1 U4806 ( .C1(n4320), .C2(ADDR_REG_9__SCAN_IN), .A(n4234), .B(n4233), 
        .ZN(n4239) );
  OAI211_X1 U4807 ( .C1(n4237), .C2(n4236), .A(n4316), .B(n4235), .ZN(n4238)
         );
  OAI211_X1 U4808 ( .C1(n4319), .C2(n4356), .A(n4239), .B(n4238), .ZN(U3249)
         );
  AOI211_X1 U4809 ( .C1(n4242), .C2(n4241), .A(n4240), .B(n4321), .ZN(n4244)
         );
  AOI211_X1 U4810 ( .C1(n4320), .C2(ADDR_REG_10__SCAN_IN), .A(n4244), .B(n4243), .ZN(n4248) );
  OAI211_X1 U4811 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4246), .A(n4316), .B(n4245), .ZN(n4247) );
  OAI211_X1 U4812 ( .C1(n4319), .C2(n4249), .A(n4248), .B(n4247), .ZN(U3250)
         );
  AOI211_X1 U4813 ( .C1(n4252), .C2(n4251), .A(n4250), .B(n4321), .ZN(n4255)
         );
  INV_X1 U4814 ( .A(n4253), .ZN(n4254) );
  AOI211_X1 U4815 ( .C1(n4320), .C2(ADDR_REG_12__SCAN_IN), .A(n4255), .B(n4254), .ZN(n4259) );
  OAI211_X1 U4816 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4257), .A(n4316), .B(n4256), .ZN(n4258) );
  OAI211_X1 U4817 ( .C1(n4319), .C2(n4353), .A(n4259), .B(n4258), .ZN(U3252)
         );
  AOI211_X1 U4818 ( .C1(n4262), .C2(n4261), .A(n4260), .B(n4321), .ZN(n4263)
         );
  AOI211_X1 U4819 ( .C1(n4320), .C2(ADDR_REG_13__SCAN_IN), .A(n4264), .B(n4263), .ZN(n4271) );
  AOI21_X1 U4820 ( .B1(n4266), .B2(n4272), .A(n4265), .ZN(n4269) );
  AOI21_X1 U4821 ( .B1(n4269), .B2(n4268), .A(n4327), .ZN(n4267) );
  OAI21_X1 U4822 ( .B1(n4269), .B2(n4268), .A(n4267), .ZN(n4270) );
  OAI211_X1 U4823 ( .C1(n4319), .C2(n4272), .A(n4271), .B(n4270), .ZN(U3253)
         );
  NAND2_X1 U4824 ( .A1(ADDR_REG_14__SCAN_IN), .A2(n4320), .ZN(n4283) );
  AOI211_X1 U4825 ( .C1(n4275), .C2(n4274), .A(n4273), .B(n4321), .ZN(n4279)
         );
  AOI211_X1 U4826 ( .C1(n3440), .C2(n4277), .A(n4276), .B(n4327), .ZN(n4278)
         );
  AOI211_X1 U4827 ( .C1(n4332), .C2(n4280), .A(n4279), .B(n4278), .ZN(n4282)
         );
  NAND3_X1 U4828 ( .A1(n4283), .A2(n4282), .A3(n4281), .ZN(U3254) );
  INV_X1 U4829 ( .A(n4320), .ZN(n4293) );
  INV_X1 U4830 ( .A(ADDR_REG_15__SCAN_IN), .ZN(n4484) );
  AOI211_X1 U4831 ( .C1(n2035), .C2(n4285), .A(n4284), .B(n4321), .ZN(n4290)
         );
  AOI211_X1 U4832 ( .C1(n4288), .C2(n4287), .A(n4286), .B(n4327), .ZN(n4289)
         );
  AOI211_X1 U4833 ( .C1(n4332), .C2(n4347), .A(n4290), .B(n4289), .ZN(n4292)
         );
  OAI211_X1 U4834 ( .C1(n4293), .C2(n4484), .A(n4292), .B(n4291), .ZN(U3255)
         );
  INV_X1 U4835 ( .A(n4294), .ZN(n4295) );
  AOI21_X1 U4836 ( .B1(n4320), .B2(ADDR_REG_16__SCAN_IN), .A(n4295), .ZN(n4305) );
  OAI21_X1 U4837 ( .B1(n4298), .B2(n4297), .A(n4296), .ZN(n4303) );
  OAI21_X1 U4838 ( .B1(n4301), .B2(n4300), .A(n4299), .ZN(n4302) );
  AOI22_X1 U4839 ( .A1(n4316), .A2(n4303), .B1(n4314), .B2(n4302), .ZN(n4304)
         );
  OAI211_X1 U4840 ( .C1(n4346), .C2(n4319), .A(n4305), .B(n4304), .ZN(U3256)
         );
  AOI21_X1 U4841 ( .B1(n4320), .B2(ADDR_REG_17__SCAN_IN), .A(n4306), .ZN(n4318) );
  OAI21_X1 U4842 ( .B1(n4309), .B2(n4308), .A(n4307), .ZN(n4315) );
  OAI21_X1 U4843 ( .B1(n4312), .B2(n4311), .A(n4310), .ZN(n4313) );
  AOI22_X1 U4844 ( .A1(n4316), .A2(n4315), .B1(n4314), .B2(n4313), .ZN(n4317)
         );
  OAI211_X1 U4845 ( .C1(n4344), .C2(n4319), .A(n4318), .B(n4317), .ZN(U3257)
         );
  NAND2_X1 U4846 ( .A1(ADDR_REG_18__SCAN_IN), .A2(n4320), .ZN(n4337) );
  AOI21_X1 U4847 ( .B1(n4323), .B2(n4322), .A(n4321), .ZN(n4335) );
  INV_X1 U4848 ( .A(n4324), .ZN(n4334) );
  NAND2_X1 U4849 ( .A1(n4326), .A2(n4325), .ZN(n4328) );
  NAND2_X1 U4850 ( .A1(n4328), .A2(n4316), .ZN(n4330) );
  AND2_X1 U4851 ( .A1(D_REG_31__SCAN_IN), .A2(n4338), .ZN(U3291) );
  INV_X1 U4852 ( .A(n4338), .ZN(n4339) );
  INV_X1 U4853 ( .A(D_REG_30__SCAN_IN), .ZN(n4568) );
  NOR2_X1 U4854 ( .A1(n4339), .A2(n4568), .ZN(U3292) );
  AND2_X1 U4855 ( .A1(D_REG_29__SCAN_IN), .A2(n4338), .ZN(U3293) );
  AND2_X1 U4856 ( .A1(D_REG_28__SCAN_IN), .A2(n4338), .ZN(U3294) );
  AND2_X1 U4857 ( .A1(D_REG_27__SCAN_IN), .A2(n4338), .ZN(U3295) );
  AND2_X1 U4858 ( .A1(D_REG_26__SCAN_IN), .A2(n4338), .ZN(U3296) );
  AND2_X1 U4859 ( .A1(D_REG_25__SCAN_IN), .A2(n4338), .ZN(U3297) );
  AND2_X1 U4860 ( .A1(D_REG_24__SCAN_IN), .A2(n4338), .ZN(U3298) );
  NOR2_X1 U4861 ( .A1(n4339), .A2(n4532), .ZN(U3299) );
  AND2_X1 U4862 ( .A1(D_REG_22__SCAN_IN), .A2(n4338), .ZN(U3300) );
  AND2_X1 U4863 ( .A1(D_REG_21__SCAN_IN), .A2(n4338), .ZN(U3301) );
  INV_X1 U4864 ( .A(D_REG_20__SCAN_IN), .ZN(n4569) );
  NOR2_X1 U4865 ( .A1(n4339), .A2(n4569), .ZN(U3302) );
  AND2_X1 U4866 ( .A1(D_REG_19__SCAN_IN), .A2(n4338), .ZN(U3303) );
  AND2_X1 U4867 ( .A1(D_REG_18__SCAN_IN), .A2(n4338), .ZN(U3304) );
  NOR2_X1 U4868 ( .A1(n4339), .A2(n4531), .ZN(U3305) );
  INV_X1 U4869 ( .A(D_REG_16__SCAN_IN), .ZN(n4534) );
  NOR2_X1 U4870 ( .A1(n4339), .A2(n4534), .ZN(U3306) );
  AND2_X1 U4871 ( .A1(D_REG_15__SCAN_IN), .A2(n4338), .ZN(U3307) );
  AND2_X1 U4872 ( .A1(D_REG_14__SCAN_IN), .A2(n4338), .ZN(U3308) );
  AND2_X1 U4873 ( .A1(D_REG_13__SCAN_IN), .A2(n4338), .ZN(U3309) );
  NOR2_X1 U4874 ( .A1(n4339), .A2(n4535), .ZN(U3310) );
  INV_X1 U4875 ( .A(D_REG_11__SCAN_IN), .ZN(n4462) );
  NOR2_X1 U4876 ( .A1(n4339), .A2(n4462), .ZN(U3311) );
  AND2_X1 U4877 ( .A1(D_REG_10__SCAN_IN), .A2(n4338), .ZN(U3312) );
  AND2_X1 U4878 ( .A1(D_REG_9__SCAN_IN), .A2(n4338), .ZN(U3313) );
  AND2_X1 U4879 ( .A1(D_REG_8__SCAN_IN), .A2(n4338), .ZN(U3314) );
  INV_X1 U4880 ( .A(D_REG_7__SCAN_IN), .ZN(n4575) );
  NOR2_X1 U4881 ( .A1(n4339), .A2(n4575), .ZN(U3315) );
  AND2_X1 U4882 ( .A1(D_REG_6__SCAN_IN), .A2(n4338), .ZN(U3316) );
  AND2_X1 U4883 ( .A1(D_REG_5__SCAN_IN), .A2(n4338), .ZN(U3317) );
  AND2_X1 U4884 ( .A1(D_REG_4__SCAN_IN), .A2(n4338), .ZN(U3318) );
  AND2_X1 U4885 ( .A1(D_REG_3__SCAN_IN), .A2(n4338), .ZN(U3319) );
  NOR2_X1 U4886 ( .A1(n4339), .A2(n4526), .ZN(U3320) );
  INV_X1 U4887 ( .A(DATAI_23_), .ZN(n4559) );
  AOI21_X1 U4888 ( .B1(U3149), .B2(n4559), .A(n4340), .ZN(U3329) );
  AOI22_X1 U4889 ( .A1(STATE_REG_SCAN_IN), .A2(n4342), .B1(n4341), .B2(U3149), 
        .ZN(U3334) );
  INV_X1 U4890 ( .A(DATAI_17_), .ZN(n4343) );
  AOI22_X1 U4891 ( .A1(STATE_REG_SCAN_IN), .A2(n4344), .B1(n4343), .B2(U3149), 
        .ZN(U3335) );
  INV_X1 U4892 ( .A(DATAI_16_), .ZN(n4345) );
  AOI22_X1 U4893 ( .A1(STATE_REG_SCAN_IN), .A2(n4346), .B1(n4345), .B2(U3149), 
        .ZN(U3336) );
  OAI22_X1 U4894 ( .A1(U3149), .A2(n4347), .B1(DATAI_15_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4348) );
  INV_X1 U4895 ( .A(n4348), .ZN(U3337) );
  INV_X1 U4896 ( .A(DATAI_14_), .ZN(n4349) );
  AOI22_X1 U4897 ( .A1(STATE_REG_SCAN_IN), .A2(n4350), .B1(n4349), .B2(U3149), 
        .ZN(U3338) );
  OAI22_X1 U4898 ( .A1(U3149), .A2(n4351), .B1(DATAI_13_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4352) );
  INV_X1 U4899 ( .A(n4352), .ZN(U3339) );
  AOI22_X1 U4900 ( .A1(STATE_REG_SCAN_IN), .A2(n4353), .B1(n2383), .B2(U3149), 
        .ZN(U3340) );
  OAI22_X1 U4901 ( .A1(U3149), .A2(n4354), .B1(DATAI_10_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4355) );
  INV_X1 U4902 ( .A(n4355), .ZN(U3342) );
  INV_X1 U4903 ( .A(DATAI_9_), .ZN(n4503) );
  AOI22_X1 U4904 ( .A1(STATE_REG_SCAN_IN), .A2(n4356), .B1(n4503), .B2(U3149), 
        .ZN(U3343) );
  OAI22_X1 U4905 ( .A1(U3149), .A2(IR_REG_0__SCAN_IN), .B1(DATAI_0_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4357) );
  INV_X1 U4906 ( .A(n4357), .ZN(U3352) );
  INV_X1 U4907 ( .A(REG0_REG_0__SCAN_IN), .ZN(n4358) );
  AOI22_X1 U4908 ( .A1(n4419), .A2(n4359), .B1(n4358), .B2(n4418), .ZN(U3467)
         );
  OAI22_X1 U4909 ( .A1(n4361), .A2(n4414), .B1(n4413), .B2(n4360), .ZN(n4362)
         );
  NOR2_X1 U4910 ( .A1(n4363), .A2(n4362), .ZN(n4420) );
  INV_X1 U4911 ( .A(REG0_REG_1__SCAN_IN), .ZN(n4364) );
  AOI22_X1 U4912 ( .A1(n4419), .A2(n4420), .B1(n4364), .B2(n4418), .ZN(U3469)
         );
  OAI22_X1 U4913 ( .A1(n4366), .A2(n4414), .B1(n4413), .B2(n4365), .ZN(n4367)
         );
  NOR2_X1 U4914 ( .A1(n4368), .A2(n4367), .ZN(n4422) );
  INV_X1 U4915 ( .A(REG0_REG_3__SCAN_IN), .ZN(n4369) );
  AOI22_X1 U4916 ( .A1(n4419), .A2(n4422), .B1(n4369), .B2(n4418), .ZN(U3473)
         );
  OAI21_X1 U4917 ( .B1(n4371), .B2(n4375), .A(n4370), .ZN(n4591) );
  INV_X1 U4918 ( .A(n4591), .ZN(n4388) );
  AOI21_X1 U4919 ( .B1(n4373), .B2(n4372), .A(n4413), .ZN(n4374) );
  AND2_X1 U4920 ( .A1(n4374), .A2(n3214), .ZN(n4594) );
  XNOR2_X1 U4921 ( .A(n4376), .B(n4375), .ZN(n4386) );
  OAI22_X1 U4922 ( .A1(n2643), .A2(n4379), .B1(n4378), .B2(n4377), .ZN(n4382)
         );
  NOR2_X1 U4923 ( .A1(n4591), .A2(n4380), .ZN(n4381) );
  AOI211_X1 U4924 ( .C1(n4384), .C2(n4383), .A(n4382), .B(n4381), .ZN(n4385)
         );
  OAI21_X1 U4925 ( .B1(n4387), .B2(n4386), .A(n4385), .ZN(n4587) );
  AOI211_X1 U4926 ( .C1(n4398), .C2(n4388), .A(n4594), .B(n4587), .ZN(n4423)
         );
  INV_X1 U4927 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4389) );
  AOI22_X1 U4928 ( .A1(n4419), .A2(n4423), .B1(n4389), .B2(n4418), .ZN(U3475)
         );
  NOR2_X1 U4929 ( .A1(n4390), .A2(n4406), .ZN(n4393) );
  INV_X1 U4930 ( .A(n4391), .ZN(n4392) );
  AOI211_X1 U4931 ( .C1(n4411), .C2(n4394), .A(n4393), .B(n4392), .ZN(n4424)
         );
  INV_X1 U4932 ( .A(REG0_REG_5__SCAN_IN), .ZN(n4523) );
  AOI22_X1 U4933 ( .A1(n4419), .A2(n4424), .B1(n4523), .B2(n4418), .ZN(U3477)
         );
  NOR3_X1 U4934 ( .A1(n4395), .A2(n3240), .A3(n4413), .ZN(n4397) );
  AOI211_X1 U4935 ( .C1(n4399), .C2(n4398), .A(n4397), .B(n4396), .ZN(n4426)
         );
  INV_X1 U4936 ( .A(REG0_REG_6__SCAN_IN), .ZN(n4506) );
  AOI22_X1 U4937 ( .A1(n4419), .A2(n4426), .B1(n4506), .B2(n4418), .ZN(U3479)
         );
  NAND3_X1 U4938 ( .A1(n3324), .A2(n4401), .A3(n4400), .ZN(n4402) );
  AND3_X1 U4939 ( .A1(n4404), .A2(n4403), .A3(n4402), .ZN(n4428) );
  INV_X1 U4940 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4405) );
  AOI22_X1 U4941 ( .A1(n4419), .A2(n4428), .B1(n4405), .B2(n4418), .ZN(U3481)
         );
  NOR2_X1 U4942 ( .A1(n4407), .A2(n4406), .ZN(n4408) );
  AOI211_X1 U4943 ( .C1(n4411), .C2(n4410), .A(n4409), .B(n4408), .ZN(n4430)
         );
  INV_X1 U4944 ( .A(REG0_REG_9__SCAN_IN), .ZN(n4511) );
  AOI22_X1 U4945 ( .A1(n4419), .A2(n4430), .B1(n4511), .B2(n4418), .ZN(U3485)
         );
  OAI22_X1 U4946 ( .A1(n4415), .A2(n4414), .B1(n4413), .B2(n4412), .ZN(n4416)
         );
  NOR2_X1 U4947 ( .A1(n4417), .A2(n4416), .ZN(n4432) );
  INV_X1 U4948 ( .A(REG0_REG_11__SCAN_IN), .ZN(n4509) );
  AOI22_X1 U4949 ( .A1(n4419), .A2(n4432), .B1(n4509), .B2(n4418), .ZN(U3489)
         );
  AOI22_X1 U4950 ( .A1(n4433), .A2(n4420), .B1(n2953), .B2(n4431), .ZN(U3519)
         );
  INV_X1 U4951 ( .A(REG1_REG_3__SCAN_IN), .ZN(n4421) );
  AOI22_X1 U4952 ( .A1(n4433), .A2(n4422), .B1(n4421), .B2(n4431), .ZN(U3521)
         );
  AOI22_X1 U4953 ( .A1(n4433), .A2(n4423), .B1(n4219), .B2(n4431), .ZN(U3522)
         );
  AOI22_X1 U4954 ( .A1(n4433), .A2(n4424), .B1(n2981), .B2(n4431), .ZN(U3523)
         );
  INV_X1 U4955 ( .A(REG1_REG_6__SCAN_IN), .ZN(n4425) );
  AOI22_X1 U4956 ( .A1(n4433), .A2(n4426), .B1(n4425), .B2(n4431), .ZN(U3524)
         );
  AOI22_X1 U4957 ( .A1(n4433), .A2(n4428), .B1(n4427), .B2(n4431), .ZN(U3525)
         );
  AOI22_X1 U4958 ( .A1(n4433), .A2(n4430), .B1(n4429), .B2(n4431), .ZN(U3527)
         );
  AOI22_X1 U4959 ( .A1(n4433), .A2(n4432), .B1(n3199), .B2(n4431), .ZN(U3529)
         );
  NOR2_X1 U4960 ( .A1(keyinput43), .A2(keyinput30), .ZN(n4434) );
  NAND3_X1 U4961 ( .A1(keyinput54), .A2(keyinput1), .A3(n4434), .ZN(n4439) );
  NAND3_X1 U4962 ( .A1(keyinput6), .A2(keyinput4), .A3(keyinput57), .ZN(n4438)
         );
  NOR3_X1 U4963 ( .A1(keyinput10), .A2(keyinput11), .A3(keyinput27), .ZN(n4436) );
  NOR3_X1 U4964 ( .A1(keyinput50), .A2(keyinput46), .A3(keyinput2), .ZN(n4435)
         );
  NAND4_X1 U4965 ( .A1(keyinput51), .A2(n4436), .A3(keyinput31), .A4(n4435), 
        .ZN(n4437) );
  NOR4_X1 U4966 ( .A1(keyinput12), .A2(n4439), .A3(n4438), .A4(n4437), .ZN(
        n4460) );
  NOR2_X1 U4967 ( .A1(keyinput29), .A2(keyinput26), .ZN(n4440) );
  NAND3_X1 U4968 ( .A1(keyinput5), .A2(keyinput15), .A3(n4440), .ZN(n4452) );
  NAND2_X1 U4969 ( .A1(keyinput17), .A2(keyinput55), .ZN(n4443) );
  NOR2_X1 U4970 ( .A1(keyinput34), .A2(keyinput56), .ZN(n4441) );
  NAND3_X1 U4971 ( .A1(keyinput52), .A2(keyinput61), .A3(n4441), .ZN(n4442) );
  NOR4_X1 U4972 ( .A1(keyinput14), .A2(keyinput53), .A3(n4443), .A4(n4442), 
        .ZN(n4444) );
  NAND4_X1 U4973 ( .A1(keyinput18), .A2(keyinput49), .A3(keyinput25), .A4(
        n4444), .ZN(n4451) );
  NOR3_X1 U4974 ( .A1(keyinput0), .A2(keyinput48), .A3(keyinput40), .ZN(n4446)
         );
  NOR3_X1 U4975 ( .A1(keyinput45), .A2(keyinput33), .A3(keyinput37), .ZN(n4445) );
  NAND4_X1 U4976 ( .A1(keyinput42), .A2(n4446), .A3(keyinput24), .A4(n4445), 
        .ZN(n4450) );
  NOR3_X1 U4977 ( .A1(keyinput63), .A2(keyinput60), .A3(keyinput9), .ZN(n4448)
         );
  NOR3_X1 U4978 ( .A1(keyinput28), .A2(keyinput22), .A3(keyinput62), .ZN(n4447) );
  NAND4_X1 U4979 ( .A1(keyinput32), .A2(n4448), .A3(keyinput3), .A4(n4447), 
        .ZN(n4449) );
  NOR4_X1 U4980 ( .A1(n4452), .A2(n4451), .A3(n4450), .A4(n4449), .ZN(n4459)
         );
  NAND3_X1 U4981 ( .A1(keyinput19), .A2(keyinput36), .A3(keyinput21), .ZN(
        n4457) );
  NAND4_X1 U4982 ( .A1(keyinput7), .A2(keyinput39), .A3(keyinput59), .A4(
        keyinput8), .ZN(n4456) );
  NOR3_X1 U4983 ( .A1(keyinput47), .A2(keyinput16), .A3(keyinput44), .ZN(n4454) );
  NOR3_X1 U4984 ( .A1(keyinput41), .A2(keyinput35), .A3(keyinput58), .ZN(n4453) );
  NAND4_X1 U4985 ( .A1(keyinput38), .A2(n4454), .A3(keyinput23), .A4(n4453), 
        .ZN(n4455) );
  NOR4_X1 U4986 ( .A1(keyinput20), .A2(n4457), .A3(n4456), .A4(n4455), .ZN(
        n4458) );
  NAND3_X1 U4987 ( .A1(n4460), .A2(n4459), .A3(n4458), .ZN(n4461) );
  NAND2_X1 U4988 ( .A1(n4461), .A2(keyinput13), .ZN(n4586) );
  INV_X1 U4989 ( .A(REG2_REG_25__SCAN_IN), .ZN(n4464) );
  AOI22_X1 U4990 ( .A1(keyinput18), .A2(n4464), .B1(keyinput13), .B2(n4462), 
        .ZN(n4463) );
  OAI21_X1 U4991 ( .B1(n4464), .B2(keyinput18), .A(n4463), .ZN(n4475) );
  INV_X1 U4992 ( .A(REG2_REG_17__SCAN_IN), .ZN(n4467) );
  AOI22_X1 U4993 ( .A1(n4467), .A2(keyinput49), .B1(n4466), .B2(keyinput29), 
        .ZN(n4465) );
  OAI221_X1 U4994 ( .B1(n4467), .B2(keyinput49), .C1(n4466), .C2(keyinput29), 
        .A(n4465), .ZN(n4474) );
  INV_X1 U4995 ( .A(keyinput5), .ZN(n4469) );
  AOI22_X1 U4996 ( .A1(U3149), .A2(keyinput26), .B1(DATAO_REG_1__SCAN_IN), 
        .B2(n4469), .ZN(n4468) );
  OAI221_X1 U4997 ( .B1(U3149), .B2(keyinput26), .C1(n4469), .C2(
        DATAO_REG_1__SCAN_IN), .A(n4468), .ZN(n4473) );
  AOI22_X1 U4998 ( .A1(n3923), .A2(keyinput15), .B1(keyinput17), .B2(n4471), 
        .ZN(n4470) );
  OAI221_X1 U4999 ( .B1(n3923), .B2(keyinput15), .C1(n4471), .C2(keyinput17), 
        .A(n4470), .ZN(n4472) );
  NOR4_X1 U5000 ( .A1(n4475), .A2(n4474), .A3(n4473), .A4(n4472), .ZN(n4521)
         );
  INV_X1 U5001 ( .A(REG2_REG_23__SCAN_IN), .ZN(n4478) );
  INV_X1 U5002 ( .A(keyinput55), .ZN(n4477) );
  AOI22_X1 U5003 ( .A1(n4478), .A2(keyinput14), .B1(ADDR_REG_1__SCAN_IN), .B2(
        n4477), .ZN(n4476) );
  OAI221_X1 U5004 ( .B1(n4478), .B2(keyinput14), .C1(n4477), .C2(
        ADDR_REG_1__SCAN_IN), .A(n4476), .ZN(n4489) );
  INV_X1 U5005 ( .A(keyinput34), .ZN(n4480) );
  AOI22_X1 U5006 ( .A1(n4219), .A2(keyinput53), .B1(ADDR_REG_4__SCAN_IN), .B2(
        n4480), .ZN(n4479) );
  OAI221_X1 U5007 ( .B1(n4219), .B2(keyinput53), .C1(n4480), .C2(
        ADDR_REG_4__SCAN_IN), .A(n4479), .ZN(n4488) );
  INV_X1 U5008 ( .A(keyinput61), .ZN(n4482) );
  AOI22_X1 U5009 ( .A1(n3242), .A2(keyinput52), .B1(ADDR_REG_9__SCAN_IN), .B2(
        n4482), .ZN(n4481) );
  OAI221_X1 U5010 ( .B1(n3242), .B2(keyinput52), .C1(n4482), .C2(
        ADDR_REG_9__SCAN_IN), .A(n4481), .ZN(n4487) );
  AOI22_X1 U5011 ( .A1(n4485), .A2(keyinput56), .B1(keyinput43), .B2(n4484), 
        .ZN(n4483) );
  OAI221_X1 U5012 ( .B1(n4485), .B2(keyinput56), .C1(n4484), .C2(keyinput43), 
        .A(n4483), .ZN(n4486) );
  NOR4_X1 U5013 ( .A1(n4489), .A2(n4488), .A3(n4487), .A4(n4486), .ZN(n4520)
         );
  AOI22_X1 U5014 ( .A1(n4492), .A2(keyinput51), .B1(n4491), .B2(keyinput6), 
        .ZN(n4490) );
  OAI221_X1 U5015 ( .B1(n4492), .B2(keyinput51), .C1(n4491), .C2(keyinput6), 
        .A(n4490), .ZN(n4501) );
  AOI22_X1 U5016 ( .A1(n4494), .A2(keyinput30), .B1(n2112), .B2(keyinput54), 
        .ZN(n4493) );
  OAI221_X1 U5017 ( .B1(n4494), .B2(keyinput30), .C1(n2112), .C2(keyinput54), 
        .A(n4493), .ZN(n4500) );
  XNOR2_X1 U5018 ( .A(REG1_REG_0__SCAN_IN), .B(keyinput1), .ZN(n4498) );
  XNOR2_X1 U5019 ( .A(REG2_REG_1__SCAN_IN), .B(keyinput11), .ZN(n4497) );
  XNOR2_X1 U5020 ( .A(REG2_REG_2__SCAN_IN), .B(keyinput27), .ZN(n4496) );
  XNOR2_X1 U5021 ( .A(keyinput10), .B(REG1_REG_5__SCAN_IN), .ZN(n4495) );
  NAND4_X1 U5022 ( .A1(n4498), .A2(n4497), .A3(n4496), .A4(n4495), .ZN(n4499)
         );
  NOR3_X1 U5023 ( .A1(n4501), .A2(n4500), .A3(n4499), .ZN(n4519) );
  AOI22_X1 U5024 ( .A1(n4504), .A2(keyinput2), .B1(keyinput20), .B2(n4503), 
        .ZN(n4502) );
  OAI221_X1 U5025 ( .B1(n4504), .B2(keyinput2), .C1(n4503), .C2(keyinput20), 
        .A(n4502), .ZN(n4517) );
  AOI22_X1 U5026 ( .A1(n4507), .A2(keyinput12), .B1(keyinput4), .B2(n4506), 
        .ZN(n4505) );
  OAI221_X1 U5027 ( .B1(n4507), .B2(keyinput12), .C1(n4506), .C2(keyinput4), 
        .A(n4505), .ZN(n4516) );
  AOI22_X1 U5028 ( .A1(n4510), .A2(keyinput46), .B1(n4509), .B2(keyinput31), 
        .ZN(n4508) );
  OAI221_X1 U5029 ( .B1(n4510), .B2(keyinput46), .C1(n4509), .C2(keyinput31), 
        .A(n4508), .ZN(n4515) );
  XOR2_X1 U5030 ( .A(n4511), .B(keyinput50), .Z(n4513) );
  XNOR2_X1 U5031 ( .A(REG3_REG_7__SCAN_IN), .B(keyinput57), .ZN(n4512) );
  NAND2_X1 U5032 ( .A1(n4513), .A2(n4512), .ZN(n4514) );
  NOR4_X1 U5033 ( .A1(n4517), .A2(n4516), .A3(n4515), .A4(n4514), .ZN(n4518)
         );
  NAND4_X1 U5034 ( .A1(n4521), .A2(n4520), .A3(n4519), .A4(n4518), .ZN(n4585)
         );
  AOI22_X1 U5035 ( .A1(n4524), .A2(keyinput39), .B1(n4523), .B2(keyinput59), 
        .ZN(n4522) );
  OAI221_X1 U5036 ( .B1(n4524), .B2(keyinput39), .C1(n4523), .C2(keyinput59), 
        .A(n4522), .ZN(n4529) );
  XNOR2_X1 U5037 ( .A(n4525), .B(keyinput8), .ZN(n4528) );
  XNOR2_X1 U5038 ( .A(n4526), .B(keyinput41), .ZN(n4527) );
  OR3_X1 U5039 ( .A1(n4529), .A2(n4528), .A3(n4527), .ZN(n4538) );
  AOI22_X1 U5040 ( .A1(n4532), .A2(keyinput23), .B1(keyinput35), .B2(n4531), 
        .ZN(n4530) );
  OAI221_X1 U5041 ( .B1(n4532), .B2(keyinput23), .C1(n4531), .C2(keyinput35), 
        .A(n4530), .ZN(n4537) );
  AOI22_X1 U5042 ( .A1(n4535), .A2(keyinput58), .B1(keyinput63), .B2(n4534), 
        .ZN(n4533) );
  OAI221_X1 U5043 ( .B1(n4535), .B2(keyinput58), .C1(n4534), .C2(keyinput63), 
        .A(n4533), .ZN(n4536) );
  NOR3_X1 U5044 ( .A1(n4538), .A2(n4537), .A3(n4536), .ZN(n4583) );
  INV_X1 U5045 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4541) );
  INV_X1 U5046 ( .A(keyinput44), .ZN(n4540) );
  AOI22_X1 U5047 ( .A1(n4541), .A2(keyinput7), .B1(DATAO_REG_25__SCAN_IN), 
        .B2(n4540), .ZN(n4539) );
  OAI221_X1 U5048 ( .B1(n4541), .B2(keyinput7), .C1(n4540), .C2(
        DATAO_REG_25__SCAN_IN), .A(n4539), .ZN(n4553) );
  INV_X1 U5049 ( .A(keyinput21), .ZN(n4543) );
  AOI22_X1 U5050 ( .A1(n4544), .A2(keyinput38), .B1(DATAO_REG_23__SCAN_IN), 
        .B2(n4543), .ZN(n4542) );
  OAI221_X1 U5051 ( .B1(n4544), .B2(keyinput38), .C1(n4543), .C2(
        DATAO_REG_23__SCAN_IN), .A(n4542), .ZN(n4552) );
  INV_X1 U5052 ( .A(REG2_REG_24__SCAN_IN), .ZN(n4547) );
  AOI22_X1 U5053 ( .A1(n4547), .A2(keyinput47), .B1(n4546), .B2(keyinput16), 
        .ZN(n4545) );
  OAI221_X1 U5054 ( .B1(n4547), .B2(keyinput47), .C1(n4546), .C2(keyinput16), 
        .A(n4545), .ZN(n4551) );
  XNOR2_X1 U5055 ( .A(REG0_REG_17__SCAN_IN), .B(keyinput36), .ZN(n4549) );
  XNOR2_X1 U5056 ( .A(IR_REG_11__SCAN_IN), .B(keyinput19), .ZN(n4548) );
  NAND2_X1 U5057 ( .A1(n4549), .A2(n4548), .ZN(n4550) );
  NOR4_X1 U5058 ( .A1(n4553), .A2(n4552), .A3(n4551), .A4(n4550), .ZN(n4582)
         );
  INV_X1 U5059 ( .A(DATAI_25_), .ZN(n4556) );
  AOI22_X1 U5060 ( .A1(n4556), .A2(keyinput40), .B1(keyinput24), .B2(n4555), 
        .ZN(n4554) );
  OAI221_X1 U5061 ( .B1(n4556), .B2(keyinput40), .C1(n4555), .C2(keyinput24), 
        .A(n4554), .ZN(n4566) );
  AOI22_X1 U5062 ( .A1(n4559), .A2(keyinput0), .B1(keyinput48), .B2(n4558), 
        .ZN(n4557) );
  OAI221_X1 U5063 ( .B1(n4559), .B2(keyinput0), .C1(n4558), .C2(keyinput48), 
        .A(n4557), .ZN(n4565) );
  XNOR2_X1 U5064 ( .A(DATAI_14_), .B(keyinput25), .ZN(n4563) );
  XNOR2_X1 U5065 ( .A(IR_REG_29__SCAN_IN), .B(keyinput37), .ZN(n4562) );
  XNOR2_X1 U5066 ( .A(IR_REG_22__SCAN_IN), .B(keyinput33), .ZN(n4561) );
  XNOR2_X1 U5067 ( .A(keyinput45), .B(DATAI_4_), .ZN(n4560) );
  NAND4_X1 U5068 ( .A1(n4563), .A2(n4562), .A3(n4561), .A4(n4560), .ZN(n4564)
         );
  NOR3_X1 U5069 ( .A1(n4566), .A2(n4565), .A3(n4564), .ZN(n4581) );
  AOI22_X1 U5070 ( .A1(n4569), .A2(keyinput32), .B1(keyinput60), .B2(n4568), 
        .ZN(n4567) );
  OAI221_X1 U5071 ( .B1(n4569), .B2(keyinput32), .C1(n4568), .C2(keyinput60), 
        .A(n4567), .ZN(n4579) );
  AOI22_X1 U5072 ( .A1(n4571), .A2(keyinput62), .B1(keyinput42), .B2(n2383), 
        .ZN(n4570) );
  OAI221_X1 U5073 ( .B1(n4571), .B2(keyinput62), .C1(n2383), .C2(keyinput42), 
        .A(n4570), .ZN(n4578) );
  XNOR2_X1 U5074 ( .A(IR_REG_19__SCAN_IN), .B(keyinput28), .ZN(n4574) );
  XNOR2_X1 U5075 ( .A(IR_REG_30__SCAN_IN), .B(keyinput22), .ZN(n4573) );
  XNOR2_X1 U5076 ( .A(keyinput3), .B(DATAI_19_), .ZN(n4572) );
  NAND3_X1 U5077 ( .A1(n4574), .A2(n4573), .A3(n4572), .ZN(n4577) );
  XNOR2_X1 U5078 ( .A(n4575), .B(keyinput9), .ZN(n4576) );
  NOR4_X1 U5079 ( .A1(n4579), .A2(n4578), .A3(n4577), .A4(n4576), .ZN(n4580)
         );
  NAND4_X1 U5080 ( .A1(n4583), .A2(n4582), .A3(n4581), .A4(n4580), .ZN(n4584)
         );
  AOI211_X1 U5081 ( .C1(D_REG_11__SCAN_IN), .C2(n4586), .A(n4585), .B(n4584), 
        .ZN(n4599) );
  INV_X1 U5082 ( .A(n4587), .ZN(n4588) );
  OAI211_X1 U5083 ( .C1(n4590), .C2(n4589), .A(n4588), .B(n4595), .ZN(n4597)
         );
  NOR2_X1 U5084 ( .A1(n4591), .A2(n2603), .ZN(n4593) );
  MUX2_X1 U5085 ( .A(n4594), .B(n4593), .S(n4592), .Z(n4596) );
  OAI22_X1 U5086 ( .A1(n4597), .A2(n4596), .B1(REG2_REG_4__SCAN_IN), .B2(n4595), .ZN(n4598) );
  XNOR2_X1 U5087 ( .A(n4599), .B(n4598), .ZN(U3286) );
  CLKBUF_X1 U2257 ( .A(n2261), .Z(n3667) );
endmodule

