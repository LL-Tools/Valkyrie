

module b17_C_2inp_gates_syn ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, 
        DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, 
        DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, 
        DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, 
        DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, 
        DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, 
        READY1, READY2, P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN, 
        P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN, 
        P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN, 
        P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN, 
        P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN, 
        P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN, 
        P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN, 
        P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN, 
        P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN, 
        P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN, 
        P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN, 
        P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN, 
        P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN, 
        P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN, 
        P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN, 
        P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN, 
        P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN, 
        P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, 
        P1_REIP_REG_6__SCAN_IN, P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, 
        P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, 
        P1_REIP_REG_0__SCAN_IN, P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, 
        P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, 
        P1_EBX_REG_26__SCAN_IN, P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, 
        P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, 
        P1_EBX_REG_20__SCAN_IN, P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, 
        P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, 
        P1_EBX_REG_14__SCAN_IN, P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, 
        P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, 
        P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, 
        P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, 
        P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, 
        P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, 
        P1_EAX_REG_28__SCAN_IN, P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, 
        P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, 
        P1_EAX_REG_22__SCAN_IN, P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, 
        P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, 
        P1_EAX_REG_16__SCAN_IN, P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, 
        P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, 
        P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, 
        P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, 
        P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, 
        P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, U355, 
        U356, U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, 
        U369, U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, 
        U352, U353, U354, U365, U376, U247, U246, U245, U244, U243, U242, U241, 
        U240, U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, 
        U228, U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, 
        U216, U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, 
        U262, U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, 
        U274, U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, 
        U214, P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, 
        P3_U3059, P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, 
        P3_U3052, P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, 
        P3_U3045, P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, 
        P3_U3038, P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, 
        P3_U3031, P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, 
        P3_U3026, P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, 
        P3_U3019, P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, 
        P3_U3012, P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, 
        P3_U3005, P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, 
        P3_U3282, P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, 
        P3_U2992, P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, 
        P3_U2985, P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, 
        P3_U2978, P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, 
        P3_U2971, P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, 
        P3_U2964, P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, 
        P3_U2957, P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, 
        P3_U2950, P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, 
        P3_U2943, P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, 
        P3_U2936, P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, 
        P3_U2929, P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, 
        P3_U2922, P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, 
        P3_U2915, P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, 
        P3_U2908, P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, 
        P3_U2901, P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, 
        P3_U2894, P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, 
        P3_U2887, P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, 
        P3_U2880, P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, 
        P3_U2873, P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, 
        P3_U3285, P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, 
        P3_U2864, P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, 
        P3_U2857, P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, 
        P3_U2850, P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, 
        P3_U2843, P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, 
        P3_U2836, P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, 
        P3_U2829, P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, 
        P3_U2822, P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, 
        P3_U2815, P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, 
        P3_U2808, P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, 
        P3_U2801, P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, 
        P3_U2794, P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, 
        P3_U2787, P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, 
        P3_U2780, P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, 
        P3_U2773, P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, 
        P3_U2766, P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, 
        P3_U2759, P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, 
        P3_U2752, P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, 
        P3_U2745, P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, 
        P3_U2738, P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, 
        P3_U2731, P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, 
        P3_U2724, P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, 
        P3_U2717, P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, 
        P3_U2710, P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, 
        P3_U2703, P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, 
        P3_U2696, P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, 
        P3_U2689, P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, 
        P3_U2682, P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, 
        P3_U2675, P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, 
        P3_U2668, P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, 
        P3_U2661, P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, 
        P3_U2654, P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, 
        P3_U2647, P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, 
        P3_U2640, P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, 
        P3_U3295, P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, 
        P3_U3298, P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, 
        P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, 
        P2_U3179, P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, 
        P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, 
        P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, 
        P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, 
        P2_U3152, P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, 
        P2_U3145, P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, 
        P2_U3138, P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, 
        P2_U3131, P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, 
        P2_U3124, P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, 
        P2_U3117, P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, 
        P2_U3110, P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, 
        P2_U3103, P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, 
        P2_U3096, P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, 
        P2_U3089, P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, 
        P2_U3082, P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, 
        P2_U3075, P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, 
        P2_U3068, P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, 
        P2_U3061, P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, 
        P2_U3054, P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, 
        P2_U3595, P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, 
        P2_U3603, P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, 
        P2_U3042, P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, 
        P2_U3035, P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, 
        P2_U3028, P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, 
        P2_U3021, P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, 
        P2_U3014, P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, 
        P2_U3007, P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, 
        P2_U3000, P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, 
        P2_U2993, P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, 
        P2_U2986, P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, 
        P2_U2979, P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, 
        P2_U2972, P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, 
        P2_U2965, P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, 
        P2_U2958, P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, 
        P2_U2951, P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, 
        P2_U2944, P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, 
        P2_U2937, P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, 
        P2_U2930, P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, 
        P2_U2923, P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, 
        P2_U2916, P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, 
        P2_U2909, P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, 
        P2_U2902, P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, 
        P2_U2895, P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, 
        P2_U2888, P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, 
        P2_U2881, P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, 
        P2_U2874, P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, 
        P2_U2867, P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, 
        P2_U2860, P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, 
        P2_U2853, P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, 
        P2_U2846, P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, 
        P2_U2839, P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, 
        P2_U2832, P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, 
        P2_U2825, P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, 
        P2_U2819, P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, 
        P2_U2815, P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, 
        P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, 
        P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, 
        P1_U3212, P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, 
        P1_U3205, P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, 
        P1_U3198, P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, 
        P1_U3193, P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, 
        P1_U3186, P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, 
        P1_U3179, P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, 
        P1_U3172, P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, 
        P1_U3165, P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, 
        P1_U3159, P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, 
        P1_U3152, P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, 
        P1_U3145, P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, 
        P1_U3138, P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, 
        P1_U3131, P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, 
        P1_U3124, P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, 
        P1_U3117, P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, 
        P1_U3110, P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, 
        P1_U3103, P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, 
        P1_U3096, P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, 
        P1_U3089, P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, 
        P1_U3082, P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, 
        P1_U3075, P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, 
        P1_U3068, P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, 
        P1_U3061, P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, 
        P1_U3054, P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, 
        P1_U3047, P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, 
        P1_U3040, P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, 
        P1_U3033, P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, 
        P1_U3475, P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, 
        P1_U3028, P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, 
        P1_U3021, P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, 
        P1_U3014, P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, 
        P1_U3007, P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, 
        P1_U3000, P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, 
        P1_U2993, P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, 
        P1_U2986, P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, 
        P1_U2979, P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, 
        P1_U2972, P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, 
        P1_U2965, P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, 
        P1_U2958, P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, 
        P1_U2951, P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, 
        P1_U2944, P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, 
        P1_U2937, P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, 
        P1_U2930, P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, 
        P1_U2923, P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, 
        P1_U2916, P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, 
        P1_U2909, P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, 
        P1_U2902, P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, 
        P1_U2895, P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, 
        P1_U2888, P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, 
        P1_U2881, P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, 
        P1_U2874, P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, 
        P1_U2867, P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, 
        P1_U2860, P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, 
        P1_U2853, P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, 
        P1_U2846, P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, 
        P1_U2839, P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, 
        P1_U2832, P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, 
        P1_U2825, P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, 
        P1_U2818, P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, 
        P1_U2811, P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, 
        P1_U3483, P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, 
        P1_U2803, P1_U2802, P1_U3487, P1_U2801, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput0, keyinput1, keyinput2,
         keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8,
         keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685,
         n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695,
         n9696, n9697, n9698, n9699, n9701, n9702, n9703, n9704, n9705, n9706,
         n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716,
         n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726,
         n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736,
         n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746,
         n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756,
         n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766,
         n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776,
         n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786,
         n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796,
         n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806,
         n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816,
         n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826,
         n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836,
         n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846,
         n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856,
         n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866,
         n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876,
         n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886,
         n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896,
         n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906,
         n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916,
         n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926,
         n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936,
         n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946,
         n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956,
         n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966,
         n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976,
         n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986,
         n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996,
         n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005,
         n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013,
         n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021,
         n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029,
         n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037,
         n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045,
         n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053,
         n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061,
         n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069,
         n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077,
         n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085,
         n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093,
         n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101,
         n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109,
         n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117,
         n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125,
         n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133,
         n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141,
         n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149,
         n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157,
         n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165,
         n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173,
         n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181,
         n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189,
         n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197,
         n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205,
         n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213,
         n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221,
         n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229,
         n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237,
         n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245,
         n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253,
         n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261,
         n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269,
         n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277,
         n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285,
         n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293,
         n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301,
         n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309,
         n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317,
         n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325,
         n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333,
         n10334, n10335, n10336, n10337, n10338, n10339, n10340, n10341,
         n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349,
         n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357,
         n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365,
         n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373,
         n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381,
         n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389,
         n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397,
         n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405,
         n10406, n10407, n10408, n10409, n10410, n10411, n10412, n10413,
         n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421,
         n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429,
         n10430, n10431, n10432, n10433, n10434, n10435, n10436, n10437,
         n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445,
         n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453,
         n10454, n10455, n10456, n10457, n10458, n10459, n10460, n10461,
         n10462, n10463, n10464, n10465, n10466, n10467, n10468, n10469,
         n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477,
         n10478, n10479, n10480, n10481, n10482, n10483, n10484, n10485,
         n10486, n10487, n10488, n10489, n10490, n10491, n10492, n10493,
         n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501,
         n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509,
         n10510, n10511, n10512, n10513, n10514, n10515, n10516, n10517,
         n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525,
         n10526, n10527, n10528, n10529, n10530, n10531, n10532, n10533,
         n10534, n10535, n10536, n10537, n10538, n10539, n10540, n10541,
         n10542, n10543, n10544, n10545, n10546, n10547, n10548, n10549,
         n10550, n10551, n10552, n10553, n10554, n10555, n10556, n10557,
         n10558, n10559, n10560, n10561, n10562, n10563, n10564, n10565,
         n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10573,
         n10574, n10575, n10576, n10577, n10578, n10579, n10580, n10581,
         n10582, n10583, n10584, n10585, n10586, n10587, n10588, n10589,
         n10590, n10591, n10592, n10593, n10594, n10595, n10596, n10597,
         n10598, n10599, n10600, n10601, n10602, n10603, n10604, n10605,
         n10606, n10607, n10608, n10609, n10610, n10611, n10612, n10613,
         n10614, n10615, n10616, n10617, n10618, n10619, n10620, n10621,
         n10622, n10623, n10624, n10625, n10626, n10627, n10628, n10629,
         n10630, n10631, n10632, n10633, n10634, n10635, n10636, n10637,
         n10638, n10639, n10640, n10641, n10642, n10644, n10645, n10646,
         n10647, n10648, n10649, n10650, n10651, n10652, n10653, n10654,
         n10655, n10656, n10657, n10658, n10659, n10660, n10661, n10662,
         n10663, n10664, n10665, n10666, n10667, n10668, n10669, n10670,
         n10671, n10672, n10673, n10674, n10675, n10676, n10677, n10678,
         n10679, n10680, n10681, n10682, n10683, n10684, n10685, n10686,
         n10687, n10688, n10689, n10690, n10691, n10692, n10693, n10694,
         n10695, n10696, n10697, n10698, n10699, n10700, n10701, n10702,
         n10703, n10704, n10705, n10706, n10707, n10708, n10709, n10710,
         n10711, n10712, n10713, n10714, n10715, n10716, n10717, n10718,
         n10719, n10720, n10721, n10722, n10723, n10724, n10725, n10726,
         n10727, n10728, n10729, n10730, n10731, n10732, n10733, n10734,
         n10735, n10736, n10737, n10738, n10739, n10740, n10741, n10742,
         n10743, n10744, n10745, n10746, n10747, n10748, n10749, n10750,
         n10751, n10752, n10753, n10754, n10755, n10756, n10757, n10758,
         n10759, n10760, n10761, n10762, n10763, n10764, n10765, n10766,
         n10767, n10768, n10769, n10770, n10771, n10772, n10773, n10774,
         n10775, n10776, n10777, n10778, n10779, n10780, n10781, n10782,
         n10783, n10784, n10785, n10786, n10787, n10788, n10789, n10790,
         n10791, n10792, n10793, n10794, n10795, n10796, n10797, n10798,
         n10799, n10800, n10801, n10802, n10803, n10804, n10805, n10806,
         n10807, n10808, n10809, n10810, n10811, n10812, n10813, n10814,
         n10815, n10816, n10817, n10818, n10819, n10820, n10821, n10822,
         n10823, n10824, n10825, n10826, n10827, n10828, n10829, n10830,
         n10831, n10832, n10833, n10834, n10835, n10836, n10837, n10838,
         n10839, n10840, n10841, n10842, n10843, n10844, n10845, n10846,
         n10847, n10848, n10849, n10850, n10851, n10852, n10853, n10854,
         n10855, n10856, n10857, n10858, n10859, n10860, n10861, n10862,
         n10863, n10864, n10865, n10866, n10867, n10868, n10869, n10870,
         n10871, n10872, n10873, n10874, n10875, n10876, n10877, n10878,
         n10879, n10880, n10881, n10882, n10883, n10884, n10885, n10886,
         n10887, n10888, n10889, n10890, n10891, n10892, n10893, n10894,
         n10895, n10896, n10897, n10898, n10899, n10900, n10901, n10902,
         n10903, n10904, n10905, n10906, n10907, n10908, n10909, n10910,
         n10911, n10912, n10913, n10914, n10915, n10916, n10917, n10918,
         n10919, n10920, n10921, n10922, n10923, n10924, n10925, n10926,
         n10927, n10928, n10929, n10930, n10931, n10932, n10933, n10934,
         n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942,
         n10943, n10944, n10945, n10946, n10947, n10948, n10949, n10950,
         n10951, n10952, n10953, n10954, n10955, n10956, n10957, n10958,
         n10959, n10960, n10961, n10962, n10963, n10964, n10965, n10966,
         n10967, n10968, n10969, n10970, n10971, n10972, n10973, n10974,
         n10975, n10976, n10977, n10978, n10979, n10980, n10981, n10982,
         n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990,
         n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998,
         n10999, n11000, n11001, n11002, n11003, n11004, n11005, n11006,
         n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014,
         n11015, n11016, n11017, n11018, n11019, n11020, n11021, n11022,
         n11023, n11024, n11025, n11026, n11027, n11028, n11029, n11030,
         n11031, n11032, n11033, n11034, n11035, n11036, n11037, n11038,
         n11039, n11040, n11041, n11042, n11043, n11044, n11045, n11046,
         n11047, n11048, n11049, n11050, n11051, n11052, n11053, n11054,
         n11055, n11056, n11057, n11058, n11059, n11060, n11061, n11062,
         n11063, n11064, n11065, n11066, n11067, n11068, n11069, n11070,
         n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078,
         n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086,
         n11087, n11088, n11089, n11090, n11091, n11092, n11093, n11094,
         n11095, n11096, n11097, n11098, n11099, n11100, n11101, n11102,
         n11103, n11104, n11105, n11106, n11107, n11108, n11109, n11110,
         n11111, n11112, n11113, n11114, n11115, n11116, n11117, n11118,
         n11119, n11120, n11121, n11122, n11123, n11124, n11125, n11126,
         n11127, n11128, n11129, n11130, n11131, n11132, n11133, n11134,
         n11135, n11136, n11137, n11138, n11139, n11140, n11141, n11142,
         n11143, n11144, n11145, n11146, n11147, n11148, n11149, n11150,
         n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11158,
         n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166,
         n11167, n11168, n11169, n11170, n11171, n11172, n11173, n11174,
         n11175, n11176, n11177, n11178, n11179, n11180, n11181, n11182,
         n11183, n11184, n11185, n11186, n11187, n11188, n11189, n11190,
         n11191, n11192, n11193, n11194, n11195, n11196, n11197, n11198,
         n11199, n11200, n11201, n11202, n11203, n11204, n11205, n11206,
         n11207, n11208, n11209, n11210, n11211, n11212, n11213, n11214,
         n11215, n11216, n11217, n11218, n11219, n11220, n11221, n11222,
         n11223, n11224, n11225, n11226, n11227, n11228, n11229, n11230,
         n11231, n11232, n11233, n11234, n11235, n11236, n11237, n11238,
         n11239, n11240, n11241, n11242, n11243, n11244, n11245, n11246,
         n11247, n11248, n11249, n11250, n11251, n11252, n11253, n11254,
         n11255, n11256, n11257, n11258, n11259, n11260, n11261, n11262,
         n11263, n11264, n11265, n11266, n11267, n11268, n11269, n11270,
         n11271, n11272, n11273, n11274, n11275, n11276, n11277, n11278,
         n11279, n11280, n11281, n11282, n11283, n11284, n11285, n11286,
         n11287, n11288, n11289, n11290, n11291, n11292, n11293, n11294,
         n11295, n11296, n11297, n11298, n11299, n11300, n11301, n11302,
         n11303, n11304, n11305, n11306, n11307, n11308, n11309, n11310,
         n11311, n11312, n11313, n11314, n11315, n11316, n11317, n11318,
         n11319, n11320, n11321, n11322, n11323, n11324, n11325, n11326,
         n11327, n11328, n11329, n11330, n11331, n11332, n11333, n11334,
         n11335, n11336, n11337, n11338, n11339, n11340, n11341, n11342,
         n11343, n11344, n11345, n11346, n11347, n11348, n11349, n11350,
         n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358,
         n11359, n11360, n11361, n11362, n11363, n11364, n11365, n11366,
         n11367, n11368, n11369, n11370, n11371, n11372, n11373, n11374,
         n11375, n11376, n11377, n11378, n11379, n11380, n11381, n11382,
         n11383, n11384, n11385, n11386, n11387, n11388, n11389, n11390,
         n11391, n11392, n11393, n11394, n11395, n11396, n11397, n11398,
         n11399, n11400, n11401, n11402, n11403, n11404, n11405, n11406,
         n11407, n11408, n11409, n11410, n11411, n11412, n11413, n11414,
         n11415, n11416, n11417, n11418, n11419, n11420, n11421, n11422,
         n11423, n11424, n11425, n11426, n11427, n11428, n11429, n11430,
         n11431, n11432, n11433, n11434, n11435, n11436, n11437, n11438,
         n11439, n11440, n11441, n11442, n11443, n11444, n11445, n11446,
         n11447, n11448, n11449, n11450, n11451, n11452, n11453, n11454,
         n11455, n11456, n11457, n11458, n11459, n11460, n11461, n11462,
         n11463, n11464, n11465, n11466, n11467, n11468, n11469, n11470,
         n11471, n11472, n11473, n11474, n11475, n11476, n11477, n11478,
         n11479, n11480, n11481, n11482, n11483, n11484, n11485, n11486,
         n11487, n11488, n11489, n11490, n11491, n11492, n11493, n11494,
         n11495, n11496, n11497, n11498, n11499, n11500, n11501, n11502,
         n11503, n11504, n11505, n11506, n11507, n11508, n11509, n11510,
         n11511, n11512, n11513, n11514, n11515, n11516, n11517, n11518,
         n11519, n11520, n11521, n11522, n11523, n11524, n11525, n11526,
         n11527, n11528, n11529, n11530, n11531, n11532, n11533, n11534,
         n11535, n11536, n11537, n11538, n11539, n11540, n11541, n11542,
         n11543, n11544, n11545, n11546, n11547, n11548, n11549, n11550,
         n11551, n11552, n11553, n11554, n11555, n11556, n11557, n11558,
         n11559, n11560, n11561, n11562, n11563, n11564, n11565, n11566,
         n11567, n11568, n11569, n11570, n11571, n11572, n11573, n11574,
         n11575, n11576, n11577, n11578, n11579, n11580, n11581, n11582,
         n11583, n11584, n11585, n11586, n11587, n11588, n11589, n11590,
         n11591, n11592, n11593, n11594, n11595, n11596, n11597, n11598,
         n11599, n11600, n11601, n11602, n11603, n11604, n11605, n11606,
         n11607, n11608, n11609, n11610, n11611, n11612, n11613, n11614,
         n11615, n11616, n11617, n11618, n11619, n11620, n11621, n11622,
         n11623, n11624, n11625, n11626, n11627, n11628, n11629, n11630,
         n11631, n11632, n11633, n11634, n11635, n11636, n11637, n11638,
         n11639, n11640, n11641, n11642, n11643, n11644, n11645, n11646,
         n11647, n11648, n11649, n11650, n11651, n11652, n11653, n11654,
         n11655, n11656, n11657, n11658, n11659, n11660, n11661, n11662,
         n11663, n11664, n11665, n11666, n11667, n11668, n11669, n11670,
         n11671, n11672, n11673, n11674, n11675, n11676, n11677, n11678,
         n11679, n11680, n11681, n11682, n11683, n11684, n11685, n11686,
         n11687, n11688, n11689, n11690, n11691, n11692, n11693, n11694,
         n11695, n11696, n11697, n11698, n11699, n11700, n11701, n11702,
         n11703, n11704, n11705, n11706, n11707, n11708, n11709, n11710,
         n11711, n11712, n11713, n11714, n11715, n11716, n11717, n11718,
         n11719, n11720, n11721, n11722, n11723, n11724, n11725, n11726,
         n11727, n11728, n11729, n11730, n11731, n11732, n11733, n11734,
         n11735, n11736, n11737, n11738, n11739, n11740, n11741, n11742,
         n11743, n11744, n11745, n11746, n11747, n11748, n11749, n11750,
         n11751, n11752, n11753, n11754, n11755, n11756, n11757, n11758,
         n11759, n11760, n11761, n11762, n11763, n11764, n11765, n11766,
         n11767, n11768, n11769, n11770, n11771, n11772, n11773, n11774,
         n11775, n11776, n11777, n11778, n11779, n11780, n11781, n11782,
         n11783, n11784, n11785, n11786, n11787, n11788, n11789, n11790,
         n11791, n11792, n11793, n11794, n11795, n11796, n11797, n11798,
         n11799, n11800, n11801, n11802, n11803, n11804, n11805, n11806,
         n11807, n11808, n11809, n11810, n11811, n11812, n11813, n11814,
         n11815, n11816, n11817, n11818, n11819, n11820, n11821, n11822,
         n11823, n11824, n11825, n11826, n11827, n11828, n11829, n11830,
         n11831, n11832, n11833, n11834, n11835, n11836, n11837, n11838,
         n11839, n11840, n11841, n11842, n11843, n11844, n11845, n11846,
         n11847, n11848, n11849, n11850, n11851, n11852, n11853, n11854,
         n11855, n11856, n11857, n11858, n11859, n11860, n11861, n11862,
         n11863, n11864, n11865, n11866, n11867, n11868, n11869, n11870,
         n11871, n11872, n11873, n11874, n11875, n11876, n11877, n11878,
         n11879, n11880, n11881, n11882, n11883, n11884, n11885, n11886,
         n11887, n11888, n11889, n11890, n11891, n11892, n11893, n11894,
         n11895, n11896, n11897, n11898, n11899, n11900, n11901, n11902,
         n11903, n11904, n11905, n11906, n11907, n11908, n11909, n11910,
         n11911, n11912, n11913, n11914, n11915, n11916, n11917, n11918,
         n11919, n11920, n11921, n11922, n11923, n11924, n11925, n11926,
         n11927, n11928, n11929, n11930, n11931, n11932, n11933, n11934,
         n11935, n11936, n11937, n11938, n11939, n11940, n11941, n11942,
         n11943, n11944, n11945, n11946, n11947, n11948, n11949, n11950,
         n11951, n11952, n11953, n11954, n11955, n11956, n11957, n11958,
         n11959, n11960, n11961, n11962, n11963, n11964, n11965, n11966,
         n11967, n11968, n11969, n11970, n11971, n11972, n11973, n11974,
         n11975, n11976, n11977, n11978, n11979, n11980, n11981, n11982,
         n11983, n11984, n11985, n11986, n11987, n11988, n11989, n11990,
         n11991, n11992, n11993, n11994, n11995, n11996, n11997, n11998,
         n11999, n12000, n12001, n12002, n12003, n12004, n12005, n12006,
         n12007, n12008, n12009, n12010, n12011, n12012, n12013, n12014,
         n12015, n12016, n12017, n12018, n12019, n12020, n12021, n12022,
         n12023, n12024, n12025, n12026, n12027, n12028, n12029, n12030,
         n12031, n12032, n12033, n12034, n12035, n12036, n12037, n12038,
         n12039, n12040, n12041, n12042, n12043, n12044, n12045, n12046,
         n12047, n12048, n12049, n12050, n12051, n12052, n12053, n12054,
         n12055, n12056, n12057, n12058, n12059, n12060, n12061, n12062,
         n12063, n12064, n12065, n12066, n12067, n12068, n12069, n12070,
         n12071, n12072, n12073, n12074, n12075, n12076, n12077, n12078,
         n12079, n12080, n12081, n12082, n12083, n12084, n12085, n12086,
         n12087, n12088, n12089, n12090, n12091, n12092, n12093, n12094,
         n12095, n12096, n12097, n12098, n12099, n12100, n12101, n12102,
         n12103, n12104, n12105, n12106, n12107, n12108, n12109, n12110,
         n12111, n12112, n12113, n12114, n12115, n12116, n12117, n12118,
         n12119, n12120, n12121, n12122, n12123, n12124, n12125, n12126,
         n12127, n12128, n12129, n12130, n12131, n12132, n12133, n12134,
         n12135, n12136, n12137, n12138, n12139, n12140, n12141, n12142,
         n12143, n12144, n12145, n12146, n12147, n12148, n12149, n12150,
         n12151, n12152, n12153, n12154, n12155, n12156, n12157, n12158,
         n12159, n12160, n12161, n12162, n12163, n12164, n12165, n12166,
         n12167, n12168, n12169, n12170, n12171, n12172, n12173, n12174,
         n12175, n12176, n12177, n12178, n12179, n12180, n12181, n12182,
         n12183, n12184, n12185, n12186, n12187, n12188, n12189, n12190,
         n12191, n12192, n12193, n12194, n12195, n12196, n12197, n12198,
         n12199, n12200, n12201, n12202, n12203, n12204, n12205, n12206,
         n12207, n12208, n12209, n12210, n12211, n12212, n12213, n12214,
         n12215, n12216, n12217, n12218, n12219, n12220, n12221, n12222,
         n12223, n12224, n12225, n12226, n12227, n12228, n12229, n12230,
         n12231, n12232, n12233, n12234, n12235, n12236, n12237, n12238,
         n12239, n12240, n12241, n12242, n12243, n12244, n12245, n12246,
         n12247, n12248, n12249, n12250, n12251, n12252, n12253, n12254,
         n12255, n12256, n12257, n12258, n12259, n12260, n12261, n12262,
         n12263, n12264, n12265, n12266, n12267, n12268, n12269, n12270,
         n12271, n12272, n12273, n12274, n12275, n12276, n12277, n12278,
         n12279, n12280, n12281, n12282, n12283, n12284, n12285, n12286,
         n12287, n12288, n12289, n12290, n12291, n12292, n12293, n12294,
         n12295, n12296, n12297, n12298, n12299, n12300, n12301, n12302,
         n12303, n12304, n12305, n12306, n12307, n12308, n12309, n12310,
         n12311, n12312, n12313, n12314, n12315, n12316, n12317, n12318,
         n12319, n12320, n12321, n12322, n12323, n12324, n12325, n12326,
         n12327, n12328, n12329, n12330, n12331, n12332, n12333, n12334,
         n12335, n12336, n12337, n12338, n12339, n12340, n12341, n12342,
         n12343, n12344, n12345, n12346, n12347, n12348, n12349, n12350,
         n12351, n12352, n12353, n12354, n12355, n12356, n12357, n12358,
         n12359, n12360, n12361, n12362, n12363, n12364, n12365, n12366,
         n12367, n12368, n12369, n12370, n12371, n12372, n12373, n12374,
         n12375, n12376, n12377, n12378, n12379, n12380, n12381, n12382,
         n12383, n12384, n12385, n12386, n12387, n12388, n12389, n12390,
         n12391, n12392, n12393, n12394, n12395, n12396, n12397, n12398,
         n12399, n12400, n12401, n12402, n12403, n12404, n12405, n12406,
         n12407, n12408, n12409, n12410, n12411, n12412, n12413, n12414,
         n12415, n12416, n12417, n12418, n12419, n12420, n12421, n12422,
         n12423, n12424, n12425, n12426, n12427, n12428, n12429, n12430,
         n12431, n12432, n12433, n12434, n12435, n12436, n12437, n12438,
         n12439, n12440, n12441, n12442, n12443, n12444, n12445, n12446,
         n12447, n12448, n12449, n12450, n12451, n12452, n12453, n12454,
         n12455, n12456, n12457, n12458, n12459, n12460, n12461, n12462,
         n12463, n12464, n12465, n12466, n12467, n12468, n12469, n12470,
         n12471, n12472, n12473, n12474, n12475, n12476, n12477, n12478,
         n12479, n12480, n12481, n12482, n12483, n12484, n12485, n12486,
         n12487, n12488, n12489, n12490, n12491, n12492, n12493, n12494,
         n12495, n12496, n12497, n12498, n12499, n12500, n12501, n12502,
         n12503, n12504, n12505, n12506, n12507, n12508, n12509, n12510,
         n12511, n12512, n12513, n12514, n12515, n12516, n12517, n12518,
         n12519, n12520, n12521, n12522, n12523, n12524, n12525, n12526,
         n12527, n12528, n12529, n12530, n12531, n12532, n12533, n12534,
         n12535, n12536, n12537, n12538, n12539, n12540, n12541, n12542,
         n12543, n12544, n12545, n12546, n12547, n12548, n12549, n12550,
         n12551, n12552, n12553, n12554, n12555, n12556, n12557, n12558,
         n12559, n12560, n12561, n12562, n12563, n12564, n12565, n12566,
         n12567, n12568, n12569, n12570, n12571, n12572, n12573, n12574,
         n12575, n12576, n12577, n12578, n12579, n12580, n12581, n12582,
         n12583, n12584, n12585, n12586, n12587, n12588, n12589, n12590,
         n12591, n12592, n12593, n12594, n12595, n12596, n12597, n12598,
         n12599, n12600, n12601, n12602, n12603, n12604, n12605, n12606,
         n12607, n12608, n12609, n12610, n12611, n12612, n12613, n12614,
         n12615, n12616, n12617, n12618, n12619, n12620, n12621, n12622,
         n12623, n12624, n12625, n12626, n12627, n12628, n12629, n12630,
         n12631, n12632, n12633, n12634, n12635, n12636, n12637, n12638,
         n12639, n12640, n12641, n12642, n12643, n12644, n12645, n12646,
         n12647, n12648, n12649, n12650, n12651, n12652, n12653, n12654,
         n12655, n12656, n12657, n12658, n12659, n12660, n12661, n12662,
         n12663, n12664, n12665, n12666, n12667, n12668, n12669, n12670,
         n12671, n12672, n12673, n12674, n12675, n12676, n12677, n12678,
         n12679, n12680, n12681, n12682, n12683, n12684, n12685, n12686,
         n12687, n12688, n12689, n12690, n12691, n12692, n12693, n12694,
         n12695, n12696, n12697, n12698, n12699, n12700, n12701, n12702,
         n12703, n12704, n12705, n12706, n12707, n12708, n12709, n12710,
         n12711, n12712, n12713, n12714, n12715, n12716, n12717, n12718,
         n12719, n12720, n12721, n12722, n12723, n12724, n12725, n12726,
         n12727, n12728, n12729, n12730, n12731, n12732, n12733, n12734,
         n12735, n12736, n12737, n12738, n12739, n12740, n12741, n12742,
         n12743, n12744, n12745, n12746, n12747, n12748, n12749, n12750,
         n12751, n12752, n12753, n12754, n12755, n12756, n12757, n12758,
         n12759, n12760, n12761, n12762, n12763, n12764, n12765, n12766,
         n12767, n12768, n12769, n12770, n12771, n12772, n12773, n12774,
         n12775, n12776, n12778, n12779, n12780, n12781, n12782, n12783,
         n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791,
         n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799,
         n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807,
         n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815,
         n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823,
         n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831,
         n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839,
         n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847,
         n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855,
         n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863,
         n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871,
         n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879,
         n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887,
         n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895,
         n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903,
         n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911,
         n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919,
         n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927,
         n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935,
         n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943,
         n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951,
         n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959,
         n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967,
         n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975,
         n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983,
         n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991,
         n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999,
         n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007,
         n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015,
         n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023,
         n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031,
         n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039,
         n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047,
         n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055,
         n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063,
         n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071,
         n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079,
         n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087,
         n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095,
         n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103,
         n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111,
         n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119,
         n13120, n13121, n13122, n13123, n13124, n13125, n13126, n13127,
         n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13135,
         n13136, n13137, n13138, n13139, n13140, n13141, n13142, n13143,
         n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151,
         n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159,
         n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167,
         n13168, n13169, n13170, n13171, n13172, n13173, n13174, n13175,
         n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183,
         n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191,
         n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199,
         n13200, n13201, n13202, n13203, n13204, n13205, n13206, n13207,
         n13208, n13209, n13210, n13211, n13212, n13213, n13214, n13215,
         n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223,
         n13224, n13225, n13226, n13227, n13228, n13229, n13230, n13231,
         n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239,
         n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247,
         n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255,
         n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263,
         n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271,
         n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279,
         n13280, n13281, n13282, n13283, n13284, n13285, n13286, n13287,
         n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295,
         n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303,
         n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311,
         n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319,
         n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327,
         n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335,
         n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343,
         n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351,
         n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359,
         n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367,
         n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375,
         n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383,
         n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391,
         n13392, n13393, n13394, n13395, n13396, n13397, n13398, n13399,
         n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13407,
         n13408, n13409, n13410, n13411, n13412, n13413, n13414, n13415,
         n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423,
         n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431,
         n13432, n13433, n13434, n13435, n13436, n13438, n13439, n13440,
         n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448,
         n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456,
         n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464,
         n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472,
         n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480,
         n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488,
         n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496,
         n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504,
         n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512,
         n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520,
         n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528,
         n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536,
         n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544,
         n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552,
         n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560,
         n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568,
         n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576,
         n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584,
         n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592,
         n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600,
         n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608,
         n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616,
         n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624,
         n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632,
         n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640,
         n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648,
         n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656,
         n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664,
         n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672,
         n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680,
         n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688,
         n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696,
         n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704,
         n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712,
         n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720,
         n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728,
         n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736,
         n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744,
         n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752,
         n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760,
         n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768,
         n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776,
         n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784,
         n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792,
         n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800,
         n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808,
         n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816,
         n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824,
         n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832,
         n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840,
         n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848,
         n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856,
         n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864,
         n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872,
         n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880,
         n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888,
         n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896,
         n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904,
         n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912,
         n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920,
         n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928,
         n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936,
         n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944,
         n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952,
         n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960,
         n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968,
         n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976,
         n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984,
         n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992,
         n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000,
         n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008,
         n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016,
         n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024,
         n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032,
         n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040,
         n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048,
         n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056,
         n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064,
         n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072,
         n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080,
         n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088,
         n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096,
         n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104,
         n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112,
         n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120,
         n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128,
         n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136,
         n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144,
         n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152,
         n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160,
         n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168,
         n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176,
         n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184,
         n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192,
         n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200,
         n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208,
         n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216,
         n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224,
         n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232,
         n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240,
         n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248,
         n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256,
         n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264,
         n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272,
         n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280,
         n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288,
         n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296,
         n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304,
         n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312,
         n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320,
         n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328,
         n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336,
         n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344,
         n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352,
         n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360,
         n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368,
         n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376,
         n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384,
         n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392,
         n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400,
         n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408,
         n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416,
         n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424,
         n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432,
         n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440,
         n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448,
         n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456,
         n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464,
         n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472,
         n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480,
         n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488,
         n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496,
         n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504,
         n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512,
         n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520,
         n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528,
         n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536,
         n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544,
         n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552,
         n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560,
         n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568,
         n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576,
         n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584,
         n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592,
         n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600,
         n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608,
         n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616,
         n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624,
         n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632,
         n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640,
         n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648,
         n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656,
         n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664,
         n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672,
         n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680,
         n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688,
         n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696,
         n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704,
         n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712,
         n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720,
         n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728,
         n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736,
         n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744,
         n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752,
         n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760,
         n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768,
         n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776,
         n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784,
         n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792,
         n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800,
         n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808,
         n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816,
         n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824,
         n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832,
         n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840,
         n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848,
         n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856,
         n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864,
         n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872,
         n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880,
         n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888,
         n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896,
         n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904,
         n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912,
         n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920,
         n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928,
         n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936,
         n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944,
         n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952,
         n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960,
         n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968,
         n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976,
         n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984,
         n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992,
         n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000,
         n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008,
         n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016,
         n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024,
         n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032,
         n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040,
         n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048,
         n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056,
         n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064,
         n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072,
         n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080,
         n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088,
         n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096,
         n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104,
         n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112,
         n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120,
         n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128,
         n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136,
         n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144,
         n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152,
         n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160,
         n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168,
         n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176,
         n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184,
         n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192,
         n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200,
         n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208,
         n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216,
         n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224,
         n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232,
         n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240,
         n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248,
         n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256,
         n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264,
         n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272,
         n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280,
         n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288,
         n15289, n15290, n15291, n15292, n15293, n15294, n15295, n15296,
         n15297, n15298, n15299, n15300, n15301, n15302, n15303, n15304,
         n15305, n15306, n15307, n15308, n15309, n15310, n15311, n15312,
         n15313, n15314, n15315, n15316, n15317, n15318, n15319, n15320,
         n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328,
         n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336,
         n15337, n15338, n15339, n15340, n15341, n15342, n15343, n15344,
         n15345, n15346, n15347, n15348, n15349, n15350, n15351, n15352,
         n15353, n15354, n15355, n15356, n15357, n15358, n15359, n15360,
         n15361, n15362, n15363, n15364, n15365, n15366, n15367, n15368,
         n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376,
         n15377, n15378, n15379, n15380, n15381, n15382, n15383, n15384,
         n15385, n15386, n15387, n15388, n15389, n15390, n15391, n15392,
         n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400,
         n15401, n15402, n15403, n15404, n15405, n15406, n15407, n15408,
         n15409, n15410, n15411, n15412, n15413, n15414, n15415, n15416,
         n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15424,
         n15425, n15426, n15427, n15428, n15429, n15430, n15431, n15432,
         n15433, n15434, n15435, n15436, n15437, n15438, n15439, n15440,
         n15441, n15442, n15443, n15444, n15445, n15446, n15447, n15448,
         n15449, n15450, n15451, n15452, n15453, n15454, n15455, n15456,
         n15457, n15458, n15459, n15460, n15461, n15462, n15463, n15464,
         n15465, n15466, n15467, n15468, n15469, n15470, n15471, n15472,
         n15473, n15474, n15475, n15476, n15477, n15478, n15479, n15480,
         n15481, n15482, n15483, n15484, n15485, n15486, n15487, n15488,
         n15489, n15490, n15491, n15492, n15493, n15494, n15495, n15496,
         n15497, n15498, n15499, n15500, n15501, n15502, n15503, n15504,
         n15505, n15506, n15507, n15508, n15509, n15510, n15511, n15512,
         n15513, n15514, n15515, n15516, n15517, n15518, n15519, n15520,
         n15521, n15522, n15523, n15524, n15525, n15526, n15527, n15528,
         n15529, n15530, n15531, n15532, n15533, n15534, n15535, n15536,
         n15537, n15538, n15539, n15540, n15541, n15542, n15543, n15544,
         n15545, n15546, n15547, n15548, n15549, n15550, n15551, n15552,
         n15553, n15554, n15555, n15556, n15557, n15558, n15559, n15560,
         n15561, n15562, n15563, n15564, n15565, n15566, n15567, n15568,
         n15569, n15570, n15571, n15572, n15573, n15574, n15575, n15576,
         n15577, n15578, n15579, n15580, n15581, n15582, n15583, n15584,
         n15585, n15586, n15587, n15588, n15589, n15590, n15591, n15592,
         n15593, n15594, n15595, n15596, n15597, n15598, n15599, n15600,
         n15601, n15602, n15603, n15604, n15605, n15606, n15607, n15608,
         n15609, n15610, n15611, n15612, n15613, n15614, n15615, n15616,
         n15617, n15618, n15619, n15620, n15621, n15622, n15623, n15624,
         n15625, n15626, n15627, n15628, n15629, n15630, n15631, n15632,
         n15633, n15634, n15635, n15636, n15637, n15638, n15639, n15640,
         n15641, n15642, n15643, n15644, n15645, n15646, n15647, n15648,
         n15649, n15650, n15651, n15652, n15653, n15654, n15655, n15656,
         n15657, n15658, n15659, n15660, n15661, n15662, n15663, n15664,
         n15665, n15666, n15667, n15668, n15669, n15670, n15671, n15672,
         n15673, n15674, n15675, n15676, n15677, n15678, n15679, n15680,
         n15681, n15682, n15683, n15684, n15685, n15686, n15687, n15688,
         n15689, n15690, n15691, n15692, n15693, n15694, n15695, n15696,
         n15697, n15698, n15699, n15700, n15701, n15702, n15703, n15704,
         n15705, n15706, n15707, n15708, n15709, n15710, n15711, n15712,
         n15713, n15714, n15715, n15716, n15717, n15718, n15719, n15720,
         n15721, n15722, n15723, n15724, n15725, n15726, n15727, n15728,
         n15729, n15730, n15731, n15732, n15733, n15734, n15735, n15736,
         n15737, n15738, n15739, n15740, n15741, n15742, n15743, n15744,
         n15745, n15746, n15747, n15748, n15749, n15750, n15751, n15752,
         n15753, n15754, n15755, n15756, n15757, n15758, n15759, n15760,
         n15761, n15762, n15763, n15764, n15765, n15766, n15767, n15768,
         n15769, n15770, n15771, n15772, n15773, n15774, n15775, n15776,
         n15777, n15778, n15779, n15780, n15781, n15782, n15783, n15784,
         n15785, n15786, n15787, n15788, n15789, n15790, n15791, n15792,
         n15793, n15794, n15795, n15796, n15797, n15798, n15799, n15800,
         n15801, n15802, n15803, n15804, n15805, n15806, n15807, n15808,
         n15809, n15810, n15811, n15812, n15813, n15814, n15815, n15816,
         n15817, n15818, n15819, n15820, n15821, n15822, n15823, n15824,
         n15825, n15826, n15827, n15828, n15829, n15830, n15831, n15832,
         n15833, n15834, n15835, n15836, n15837, n15838, n15839, n15840,
         n15841, n15842, n15843, n15844, n15845, n15846, n15847, n15848,
         n15849, n15850, n15851, n15852, n15853, n15854, n15855, n15856,
         n15857, n15858, n15859, n15860, n15861, n15862, n15863, n15864,
         n15865, n15866, n15867, n15868, n15869, n15870, n15871, n15872,
         n15873, n15874, n15875, n15876, n15877, n15878, n15879, n15880,
         n15881, n15882, n15883, n15884, n15885, n15886, n15887, n15888,
         n15889, n15890, n15891, n15892, n15893, n15894, n15895, n15896,
         n15897, n15898, n15899, n15900, n15901, n15902, n15903, n15904,
         n15905, n15906, n15907, n15908, n15909, n15910, n15911, n15912,
         n15913, n15914, n15915, n15916, n15917, n15918, n15919, n15920,
         n15921, n15922, n15923, n15924, n15925, n15926, n15927, n15928,
         n15929, n15930, n15931, n15932, n15933, n15934, n15935, n15936,
         n15937, n15938, n15939, n15940, n15941, n15942, n15943, n15944,
         n15945, n15946, n15947, n15948, n15949, n15950, n15951, n15952,
         n15953, n15954, n15955, n15956, n15957, n15958, n15959, n15960,
         n15961, n15962, n15963, n15964, n15965, n15966, n15967, n15968,
         n15969, n15970, n15971, n15972, n15973, n15974, n15975, n15976,
         n15977, n15978, n15979, n15980, n15981, n15982, n15983, n15984,
         n15985, n15986, n15987, n15988, n15989, n15990, n15991, n15992,
         n15993, n15994, n15995, n15996, n15997, n15998, n15999, n16000,
         n16001, n16002, n16003, n16004, n16005, n16006, n16007, n16008,
         n16009, n16010, n16011, n16012, n16013, n16014, n16015, n16016,
         n16017, n16018, n16019, n16020, n16021, n16022, n16023, n16024,
         n16025, n16026, n16027, n16028, n16029, n16030, n16031, n16032,
         n16033, n16034, n16035, n16036, n16037, n16038, n16039, n16040,
         n16041, n16042, n16043, n16044, n16045, n16046, n16047, n16048,
         n16049, n16050, n16051, n16052, n16053, n16054, n16055, n16056,
         n16057, n16058, n16059, n16060, n16061, n16062, n16063, n16064,
         n16065, n16066, n16067, n16068, n16069, n16070, n16071, n16072,
         n16073, n16074, n16075, n16076, n16077, n16078, n16079, n16080,
         n16081, n16082, n16083, n16084, n16085, n16086, n16087, n16088,
         n16089, n16090, n16091, n16092, n16093, n16094, n16095, n16096,
         n16097, n16098, n16099, n16100, n16101, n16102, n16103, n16104,
         n16105, n16106, n16107, n16108, n16109, n16110, n16111, n16112,
         n16113, n16114, n16115, n16116, n16117, n16118, n16119, n16120,
         n16121, n16122, n16123, n16124, n16125, n16126, n16127, n16128,
         n16129, n16130, n16131, n16132, n16133, n16134, n16135, n16136,
         n16137, n16138, n16139, n16140, n16141, n16142, n16143, n16144,
         n16145, n16146, n16147, n16148, n16149, n16150, n16151, n16152,
         n16153, n16154, n16155, n16156, n16157, n16158, n16159, n16160,
         n16161, n16162, n16163, n16164, n16165, n16166, n16167, n16168,
         n16169, n16170, n16171, n16172, n16173, n16174, n16175, n16176,
         n16177, n16178, n16179, n16180, n16181, n16182, n16183, n16184,
         n16185, n16186, n16187, n16188, n16189, n16190, n16191, n16192,
         n16193, n16194, n16195, n16196, n16197, n16198, n16199, n16200,
         n16201, n16202, n16203, n16204, n16205, n16206, n16207, n16208,
         n16209, n16210, n16211, n16212, n16213, n16214, n16215, n16216,
         n16217, n16218, n16219, n16220, n16221, n16222, n16223, n16224,
         n16225, n16226, n16227, n16228, n16229, n16230, n16231, n16232,
         n16233, n16234, n16235, n16236, n16237, n16238, n16239, n16240,
         n16241, n16242, n16243, n16244, n16245, n16246, n16247, n16248,
         n16249, n16250, n16251, n16252, n16253, n16254, n16255, n16256,
         n16257, n16258, n16259, n16260, n16261, n16262, n16263, n16264,
         n16265, n16266, n16267, n16268, n16269, n16270, n16271, n16272,
         n16273, n16274, n16275, n16276, n16277, n16278, n16279, n16280,
         n16281, n16282, n16283, n16284, n16285, n16286, n16287, n16288,
         n16289, n16290, n16291, n16292, n16293, n16294, n16295, n16296,
         n16297, n16298, n16299, n16300, n16301, n16302, n16303, n16304,
         n16305, n16306, n16307, n16308, n16309, n16310, n16311, n16312,
         n16313, n16314, n16315, n16316, n16317, n16318, n16319, n16320,
         n16321, n16322, n16323, n16324, n16325, n16326, n16327, n16328,
         n16329, n16330, n16331, n16332, n16333, n16334, n16335, n16336,
         n16337, n16338, n16339, n16340, n16341, n16342, n16343, n16344,
         n16345, n16346, n16347, n16348, n16349, n16350, n16351, n16352,
         n16353, n16354, n16355, n16356, n16357, n16358, n16359, n16360,
         n16361, n16362, n16363, n16364, n16365, n16366, n16367, n16368,
         n16369, n16370, n16371, n16372, n16373, n16374, n16375, n16376,
         n16377, n16378, n16379, n16380, n16381, n16382, n16383, n16384,
         n16385, n16386, n16387, n16388, n16389, n16390, n16391, n16392,
         n16393, n16394, n16395, n16396, n16397, n16398, n16399, n16400,
         n16401, n16402, n16403, n16404, n16405, n16406, n16407, n16408,
         n16409, n16410, n16411, n16412, n16413, n16414, n16415, n16416,
         n16417, n16418, n16419, n16420, n16421, n16422, n16423, n16424,
         n16425, n16426, n16427, n16428, n16429, n16430, n16431, n16432,
         n16433, n16434, n16435, n16436, n16437, n16438, n16439, n16440,
         n16441, n16442, n16443, n16444, n16445, n16446, n16447, n16448,
         n16449, n16450, n16451, n16452, n16453, n16454, n16455, n16456,
         n16457, n16458, n16459, n16460, n16461, n16462, n16463, n16464,
         n16465, n16466, n16467, n16468, n16469, n16470, n16471, n16472,
         n16473, n16475, n16476, n16477, n16478, n16479, n16480, n16481,
         n16482, n16483, n16484, n16485, n16486, n16487, n16488, n16489,
         n16490, n16491, n16492, n16493, n16494, n16495, n16496, n16497,
         n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505,
         n16506, n16507, n16508, n16509, n16510, n16511, n16512, n16513,
         n16514, n16515, n16516, n16517, n16518, n16519, n16520, n16521,
         n16522, n16523, n16524, n16525, n16526, n16527, n16528, n16529,
         n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537,
         n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545,
         n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553,
         n16554, n16555, n16556, n16557, n16558, n16559, n16560, n16561,
         n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569,
         n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577,
         n16578, n16579, n16580, n16581, n16582, n16583, n16584, n16585,
         n16586, n16587, n16588, n16589, n16590, n16591, n16592, n16593,
         n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601,
         n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609,
         n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617,
         n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625,
         n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633,
         n16634, n16635, n16636, n16637, n16638, n16639, n16640, n16641,
         n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649,
         n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657,
         n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665,
         n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673,
         n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681,
         n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689,
         n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697,
         n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705,
         n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713,
         n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721,
         n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729,
         n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737,
         n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745,
         n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753,
         n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761,
         n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769,
         n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777,
         n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785,
         n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793,
         n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801,
         n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809,
         n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817,
         n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825,
         n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833,
         n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841,
         n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849,
         n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857,
         n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865,
         n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873,
         n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881,
         n16882, n16883, n16884, n16885, n16886, n16887, n16888, n16889,
         n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897,
         n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905,
         n16906, n16907, n16908, n16909, n16910, n16911, n16912, n16913,
         n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921,
         n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929,
         n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937,
         n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945,
         n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953,
         n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961,
         n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969,
         n16970, n16971, n16972, n16973, n16974, n16975, n16976, n16977,
         n16978, n16979, n16980, n16981, n16982, n16983, n16984, n16985,
         n16986, n16987, n16988, n16989, n16990, n16991, n16992, n16993,
         n16994, n16995, n16996, n16997, n16998, n16999, n17000, n17001,
         n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009,
         n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017,
         n17018, n17019, n17020, n17021, n17022, n17023, n17024, n17025,
         n17026, n17027, n17028, n17029, n17030, n17031, n17032, n17033,
         n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17041,
         n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049,
         n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057,
         n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065,
         n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073,
         n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081,
         n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089,
         n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097,
         n17098, n17099, n17100, n17101, n17102, n17103, n17104, n17105,
         n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113,
         n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121,
         n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129,
         n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137,
         n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145,
         n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153,
         n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161,
         n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169,
         n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177,
         n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185,
         n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193,
         n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201,
         n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209,
         n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217,
         n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225,
         n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233,
         n17234, n17235, n17236, n17237, n17238, n17239, n17240, n17241,
         n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249,
         n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257,
         n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265,
         n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273,
         n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281,
         n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289,
         n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297,
         n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305,
         n17306, n17307, n17308, n17309, n17310, n17311, n17312, n17313,
         n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321,
         n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329,
         n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337,
         n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345,
         n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353,
         n17354, n17355, n17356, n17357, n17358, n17359, n17360, n17361,
         n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369,
         n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377,
         n17378, n17379, n17380, n17381, n17382, n17383, n17384, n17385,
         n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17393,
         n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401,
         n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409,
         n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417,
         n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17425,
         n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433,
         n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441,
         n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449,
         n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457,
         n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465,
         n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473,
         n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481,
         n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489,
         n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497,
         n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505,
         n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513,
         n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521,
         n17522, n17523, n17524, n17525, n17526, n17527, n17528, n17529,
         n17530, n17531, n17532, n17533, n17534, n17535, n17536, n17537,
         n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545,
         n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553,
         n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561,
         n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569,
         n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577,
         n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585,
         n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593,
         n17594, n17595, n17596, n17597, n17598, n17599, n17600, n17601,
         n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609,
         n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617,
         n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625,
         n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633,
         n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641,
         n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649,
         n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657,
         n17658, n17659, n17660, n17661, n17662, n17663, n17664, n17665,
         n17666, n17667, n17668, n17669, n17670, n17671, n17672, n17673,
         n17674, n17675, n17676, n17677, n17678, n17679, n17680, n17681,
         n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689,
         n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697,
         n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705,
         n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713,
         n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721,
         n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729,
         n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737,
         n17738, n17739, n17740, n17741, n17742, n17743, n17744, n17745,
         n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753,
         n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761,
         n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769,
         n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777,
         n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785,
         n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793,
         n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801,
         n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809,
         n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817,
         n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825,
         n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833,
         n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841,
         n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849,
         n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857,
         n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865,
         n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873,
         n17874, n17875, n17876, n17877, n17878, n17879, n17880, n17881,
         n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17889,
         n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897,
         n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905,
         n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913,
         n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921,
         n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929,
         n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937,
         n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945,
         n17946, n17947, n17948, n17949, n17950, n17951, n17952, n17953,
         n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961,
         n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969,
         n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977,
         n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985,
         n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993,
         n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001,
         n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009,
         n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017,
         n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025,
         n18026, n18027, n18028, n18029, n18030, n18031, n18032, n18033,
         n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041,
         n18042, n18043, n18044, n18045, n18046, n18047, n18048, n18049,
         n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057,
         n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065,
         n18066, n18067, n18068, n18069, n18070, n18071, n18072, n18073,
         n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18081,
         n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089,
         n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097,
         n18098, n18099, n18100, n18101, n18102, n18103, n18104, n18105,
         n18106, n18107, n18108, n18109, n18110, n18111, n18112, n18113,
         n18114, n18115, n18116, n18117, n18118, n18119, n18120, n18121,
         n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129,
         n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137,
         n18138, n18139, n18140, n18141, n18142, n18143, n18144, n18145,
         n18146, n18147, n18148, n18149, n18150, n18151, n18152, n18153,
         n18154, n18155, n18156, n18157, n18158, n18159, n18160, n18161,
         n18162, n18163, n18164, n18165, n18166, n18167, n18168, n18169,
         n18170, n18171, n18173, n18174, n18175, n18176, n18177, n18178,
         n18179, n18180, n18181, n18182, n18183, n18184, n18185, n18186,
         n18187, n18188, n18189, n18190, n18191, n18192, n18193, n18194,
         n18195, n18196, n18197, n18198, n18199, n18200, n18201, n18202,
         n18203, n18204, n18205, n18206, n18207, n18208, n18209, n18210,
         n18211, n18212, n18213, n18214, n18215, n18216, n18217, n18218,
         n18219, n18220, n18221, n18222, n18223, n18224, n18225, n18226,
         n18227, n18228, n18229, n18230, n18231, n18232, n18233, n18234,
         n18235, n18236, n18237, n18238, n18239, n18240, n18241, n18242,
         n18243, n18244, n18245, n18246, n18247, n18248, n18249, n18250,
         n18251, n18252, n18253, n18254, n18255, n18256, n18257, n18258,
         n18259, n18260, n18261, n18262, n18263, n18264, n18265, n18266,
         n18267, n18268, n18269, n18270, n18271, n18272, n18273, n18274,
         n18275, n18276, n18277, n18278, n18279, n18280, n18281, n18282,
         n18283, n18284, n18285, n18286, n18287, n18288, n18289, n18290,
         n18291, n18292, n18293, n18294, n18295, n18296, n18297, n18298,
         n18299, n18300, n18301, n18302, n18303, n18304, n18305, n18306,
         n18307, n18308, n18309, n18310, n18311, n18312, n18313, n18314,
         n18315, n18316, n18317, n18318, n18319, n18320, n18321, n18322,
         n18323, n18324, n18325, n18326, n18327, n18328, n18329, n18330,
         n18331, n18332, n18333, n18334, n18335, n18336, n18337, n18338,
         n18339, n18340, n18341, n18342, n18343, n18344, n18345, n18346,
         n18347, n18348, n18349, n18350, n18351, n18352, n18353, n18354,
         n18355, n18356, n18357, n18358, n18359, n18360, n18361, n18362,
         n18363, n18364, n18365, n18366, n18367, n18368, n18369, n18370,
         n18371, n18372, n18373, n18374, n18375, n18376, n18377, n18378,
         n18379, n18380, n18381, n18382, n18383, n18384, n18385, n18386,
         n18387, n18388, n18389, n18390, n18391, n18392, n18393, n18394,
         n18395, n18396, n18397, n18398, n18399, n18400, n18401, n18402,
         n18403, n18404, n18405, n18406, n18407, n18408, n18409, n18410,
         n18411, n18412, n18413, n18414, n18415, n18416, n18417, n18418,
         n18419, n18420, n18421, n18422, n18423, n18424, n18425, n18426,
         n18427, n18428, n18429, n18430, n18431, n18432, n18433, n18434,
         n18435, n18436, n18437, n18438, n18439, n18440, n18441, n18442,
         n18443, n18444, n18445, n18446, n18447, n18448, n18449, n18450,
         n18451, n18452, n18453, n18454, n18455, n18456, n18457, n18458,
         n18459, n18460, n18461, n18462, n18463, n18464, n18465, n18466,
         n18467, n18468, n18469, n18470, n18471, n18472, n18473, n18474,
         n18475, n18476, n18477, n18478, n18479, n18480, n18481, n18482,
         n18483, n18484, n18485, n18486, n18487, n18488, n18489, n18490,
         n18491, n18492, n18493, n18494, n18495, n18496, n18497, n18498,
         n18499, n18500, n18501, n18502, n18503, n18504, n18505, n18506,
         n18507, n18508, n18509, n18510, n18511, n18512, n18513, n18514,
         n18515, n18516, n18517, n18518, n18519, n18520, n18521, n18522,
         n18523, n18524, n18525, n18526, n18527, n18528, n18529, n18530,
         n18531, n18532, n18533, n18534, n18535, n18536, n18537, n18538,
         n18539, n18540, n18541, n18542, n18543, n18544, n18545, n18546,
         n18547, n18548, n18549, n18550, n18551, n18552, n18553, n18554,
         n18555, n18556, n18557, n18558, n18559, n18560, n18561, n18562,
         n18563, n18564, n18565, n18566, n18567, n18568, n18569, n18570,
         n18571, n18572, n18573, n18574, n18575, n18576, n18577, n18578,
         n18579, n18580, n18581, n18582, n18583, n18584, n18585, n18586,
         n18587, n18588, n18589, n18590, n18591, n18592, n18593, n18594,
         n18595, n18596, n18597, n18598, n18599, n18600, n18601, n18602,
         n18603, n18604, n18605, n18606, n18607, n18608, n18609, n18610,
         n18611, n18612, n18613, n18614, n18615, n18616, n18617, n18618,
         n18619, n18620, n18621, n18622, n18623, n18624, n18625, n18626,
         n18627, n18628, n18629, n18630, n18631, n18632, n18633, n18634,
         n18635, n18636, n18637, n18638, n18639, n18640, n18641, n18642,
         n18643, n18644, n18645, n18646, n18647, n18648, n18649, n18650,
         n18651, n18652, n18653, n18654, n18655, n18656, n18657, n18658,
         n18659, n18660, n18661, n18662, n18663, n18664, n18665, n18666,
         n18667, n18668, n18669, n18670, n18671, n18672, n18673, n18674,
         n18675, n18676, n18677, n18678, n18679, n18680, n18681, n18682,
         n18683, n18684, n18685, n18686, n18687, n18688, n18689, n18690,
         n18691, n18692, n18693, n18694, n18695, n18696, n18697, n18698,
         n18699, n18700, n18701, n18702, n18703, n18704, n18705, n18706,
         n18707, n18708, n18709, n18710, n18711, n18712, n18713, n18714,
         n18715, n18716, n18717, n18718, n18719, n18720, n18721, n18722,
         n18723, n18724, n18725, n18726, n18727, n18728, n18729, n18730,
         n18731, n18732, n18733, n18734, n18735, n18736, n18737, n18738,
         n18739, n18740, n18741, n18742, n18743, n18744, n18745, n18746,
         n18747, n18748, n18749, n18750, n18751, n18752, n18753, n18754,
         n18755, n18756, n18757, n18758, n18759, n18760, n18761, n18762,
         n18763, n18764, n18765, n18766, n18767, n18768, n18769, n18770,
         n18771, n18772, n18773, n18774, n18775, n18776, n18777, n18778,
         n18779, n18780, n18781, n18782, n18783, n18784, n18785, n18786,
         n18787, n18788, n18789, n18790, n18791, n18792, n18793, n18794,
         n18795, n18796, n18797, n18798, n18799, n18800, n18801, n18802,
         n18803, n18804, n18805, n18806, n18807, n18808, n18809, n18810,
         n18811, n18812, n18813, n18814, n18815, n18816, n18817, n18818,
         n18819, n18820, n18821, n18822, n18823, n18824, n18825, n18826,
         n18827, n18828, n18829, n18830, n18831, n18832, n18833, n18834,
         n18835, n18836, n18837, n18838, n18839, n18840, n18841, n18842,
         n18843, n18844, n18845, n18846, n18847, n18848, n18849, n18850,
         n18851, n18852, n18853, n18854, n18855, n18856, n18857, n18858,
         n18859, n18860, n18861, n18862, n18863, n18864, n18865, n18866,
         n18867, n18868, n18869, n18870, n18871, n18872, n18873, n18874,
         n18875, n18876, n18877, n18878, n18879, n18880, n18881, n18882,
         n18883, n18884, n18885, n18886, n18887, n18888, n18889, n18890,
         n18891, n18892, n18893, n18894, n18895, n18896, n18897, n18898,
         n18899, n18900, n18901, n18902, n18903, n18904, n18905, n18906,
         n18907, n18908, n18909, n18910, n18911, n18912, n18913, n18914,
         n18915, n18916, n18917, n18918, n18919, n18920, n18921, n18922,
         n18923, n18924, n18925, n18926, n18927, n18928, n18929, n18930,
         n18931, n18932, n18933, n18934, n18935, n18936, n18937, n18938,
         n18939, n18940, n18941, n18942, n18943, n18944, n18945, n18946,
         n18947, n18948, n18949, n18950, n18951, n18952, n18953, n18954,
         n18955, n18956, n18957, n18958, n18959, n18960, n18961, n18962,
         n18963, n18964, n18965, n18966, n18967, n18968, n18969, n18970,
         n18971, n18972, n18973, n18974, n18975, n18976, n18977, n18978,
         n18979, n18980, n18981, n18982, n18983, n18984, n18985, n18986,
         n18987, n18988, n18989, n18990, n18991, n18992, n18993, n18994,
         n18995, n18996, n18997, n18998, n18999, n19000, n19001, n19002,
         n19003, n19004, n19005, n19006, n19007, n19008, n19009, n19010,
         n19011, n19012, n19013, n19014, n19015, n19016, n19017, n19018,
         n19019, n19020, n19021, n19022, n19023, n19024, n19025, n19026,
         n19027, n19028, n19029, n19030, n19031, n19032, n19033, n19034,
         n19035, n19036, n19037, n19038, n19039, n19040, n19041, n19042,
         n19043, n19044, n19045, n19046, n19047, n19048, n19049, n19050,
         n19051, n19052, n19053, n19054, n19055, n19056, n19057, n19058,
         n19059, n19060, n19061, n19062, n19063, n19064, n19065, n19066,
         n19067, n19068, n19069, n19070, n19071, n19072, n19073, n19074,
         n19075, n19076, n19077, n19078, n19079, n19080, n19081, n19082,
         n19083, n19084, n19085, n19086, n19087, n19088, n19089, n19090,
         n19091, n19092, n19093, n19094, n19095, n19096, n19097, n19098,
         n19099, n19100, n19101, n19102, n19103, n19104, n19105, n19106,
         n19107, n19108, n19109, n19110, n19111, n19112, n19113, n19114,
         n19115, n19116, n19117, n19118, n19119, n19120, n19121, n19122,
         n19123, n19124, n19125, n19126, n19127, n19128, n19129, n19130,
         n19131, n19132, n19133, n19134, n19135, n19136, n19137, n19138,
         n19139, n19140, n19141, n19142, n19143, n19144, n19145, n19146,
         n19147, n19148, n19149, n19150, n19151, n19152, n19153, n19154,
         n19155, n19156, n19157, n19158, n19159, n19160, n19161, n19162,
         n19163, n19164, n19165, n19166, n19167, n19168, n19169, n19170,
         n19171, n19172, n19173, n19174, n19175, n19176, n19177, n19178,
         n19179, n19180, n19181, n19182, n19183, n19184, n19185, n19186,
         n19187, n19188, n19189, n19190, n19191, n19192, n19193, n19194,
         n19195, n19196, n19197, n19198, n19199, n19200, n19201, n19202,
         n19203, n19204, n19205, n19206, n19207, n19208, n19209, n19210,
         n19211, n19212, n19213, n19214, n19215, n19216, n19217, n19218,
         n19219, n19220, n19221, n19222, n19223, n19224, n19225, n19226,
         n19227, n19228, n19229, n19230, n19231, n19232, n19233, n19234,
         n19235, n19236, n19237, n19238, n19239, n19240, n19241, n19242,
         n19243, n19244, n19245, n19246, n19247, n19248, n19249, n19250,
         n19251, n19252, n19253, n19254, n19255, n19256, n19257, n19258,
         n19259, n19260, n19261, n19262, n19263, n19264, n19265, n19266,
         n19267, n19268, n19269, n19270, n19271, n19272, n19273, n19274,
         n19275, n19276, n19277, n19278, n19279, n19280, n19281, n19282,
         n19283, n19284, n19285, n19286, n19287, n19288, n19289, n19290,
         n19291, n19292, n19293, n19294, n19295, n19296, n19297, n19298,
         n19299, n19300, n19301, n19302, n19303, n19304, n19305, n19306,
         n19307, n19308, n19309, n19310, n19311, n19312, n19313, n19314,
         n19315, n19316, n19317, n19318, n19319, n19320, n19321, n19322,
         n19323, n19324, n19325, n19326, n19327, n19328, n19329, n19330,
         n19331, n19332, n19333, n19334, n19335, n19336, n19337, n19338,
         n19339, n19340, n19341, n19342, n19343, n19344, n19345, n19346,
         n19347, n19348, n19349, n19350, n19351, n19352, n19353, n19354,
         n19355, n19356, n19357, n19358, n19359, n19360, n19361, n19362,
         n19363, n19364, n19365, n19366, n19367, n19368, n19369, n19370,
         n19371, n19372, n19373, n19374, n19375, n19376, n19377, n19378,
         n19379, n19380, n19381, n19382, n19383, n19384, n19385, n19386,
         n19387, n19388, n19389, n19390, n19391, n19392, n19393, n19394,
         n19395, n19396, n19397, n19398, n19399, n19400, n19401, n19402,
         n19403, n19404, n19405, n19406, n19407, n19408, n19409, n19410,
         n19411, n19412, n19413, n19414, n19415, n19416, n19417, n19418,
         n19419, n19420, n19421, n19422, n19423, n19424, n19425, n19426,
         n19427, n19428, n19429, n19430, n19431, n19432, n19433, n19434,
         n19435, n19436, n19437, n19438, n19439, n19440, n19441, n19442,
         n19443, n19444, n19445, n19446, n19447, n19448, n19449, n19450,
         n19451, n19452, n19453, n19454, n19455, n19456, n19457, n19458,
         n19459, n19460, n19461, n19462, n19463, n19464, n19465, n19466,
         n19467, n19468, n19469, n19470, n19471, n19472, n19473, n19474,
         n19475, n19476, n19477, n19478, n19479, n19480, n19481, n19482,
         n19483, n19484, n19485, n19486, n19487, n19488, n19489, n19490,
         n19491, n19492, n19493, n19494, n19495, n19496, n19497, n19498,
         n19499, n19500, n19501, n19502, n19503, n19504, n19505, n19506,
         n19507, n19508, n19509, n19510, n19511, n19512, n19513, n19514,
         n19515, n19516, n19517, n19518, n19519, n19520, n19521, n19522,
         n19523, n19524, n19525, n19526, n19527, n19528, n19529, n19530,
         n19531, n19532, n19533, n19534, n19535, n19536, n19537, n19538,
         n19539, n19540, n19541, n19542, n19543, n19544, n19545, n19546,
         n19547, n19548, n19549, n19550, n19551, n19552, n19553, n19554,
         n19555, n19556, n19557, n19558, n19559, n19560, n19561, n19562,
         n19563, n19564, n19565, n19566, n19567, n19568, n19569, n19570,
         n19571, n19572, n19573, n19574, n19575, n19576, n19577, n19578,
         n19579, n19580, n19581, n19582, n19583, n19584, n19585, n19586,
         n19587, n19588, n19589, n19590, n19591, n19592, n19593, n19594,
         n19595, n19596, n19597, n19598, n19599, n19600, n19601, n19602,
         n19603, n19604, n19605, n19606, n19607, n19608, n19609, n19610,
         n19611, n19612, n19613, n19614, n19615, n19616, n19617, n19618,
         n19619, n19620, n19621, n19622, n19623, n19624, n19625, n19626,
         n19627, n19628, n19629, n19630, n19631, n19632, n19633, n19634,
         n19635, n19636, n19637, n19638, n19639, n19640, n19641, n19642,
         n19643, n19644, n19645, n19646, n19647, n19648, n19649, n19650,
         n19651, n19652, n19653, n19654, n19655, n19656, n19657, n19658,
         n19659, n19660, n19661, n19662, n19663, n19664, n19665, n19666,
         n19667, n19668, n19669, n19670, n19671, n19672, n19673, n19674,
         n19675, n19676, n19677, n19678, n19679, n19680, n19681, n19682,
         n19683, n19684, n19685, n19686, n19687, n19688, n19689, n19690,
         n19691, n19692, n19693, n19694, n19695, n19696, n19697, n19698,
         n19699, n19700, n19701, n19702, n19703, n19704, n19705, n19706,
         n19707, n19708, n19709, n19710, n19711, n19712, n19713, n19714,
         n19715, n19716, n19717, n19718, n19719, n19720, n19721, n19722,
         n19723, n19724, n19725, n19726, n19727, n19728, n19729, n19730,
         n19731, n19732, n19733, n19734, n19735, n19736, n19737, n19738,
         n19739, n19740, n19741, n19742, n19743, n19744, n19745, n19746,
         n19747, n19748, n19749, n19750, n19751, n19752, n19753, n19754,
         n19755, n19756, n19757, n19758, n19759, n19760, n19761, n19762,
         n19763, n19764, n19765, n19766, n19767, n19768, n19769, n19770,
         n19771, n19772, n19773, n19774, n19775, n19776, n19777, n19778,
         n19779, n19780, n19781, n19782, n19783, n19784, n19785, n19786,
         n19787, n19788, n19789, n19790, n19791, n19792, n19793, n19794,
         n19795, n19796, n19797, n19798, n19799, n19800, n19801, n19802,
         n19803, n19804, n19805, n19806, n19807, n19808, n19809, n19810,
         n19811, n19812, n19813, n19814, n19815, n19816, n19817, n19818,
         n19819, n19820, n19821, n19822, n19823, n19824, n19825, n19826,
         n19827, n19828, n19829, n19830, n19831, n19832, n19833, n19834,
         n19835, n19836, n19837, n19838, n19839, n19840, n19841, n19842,
         n19843, n19844, n19845, n19846, n19847, n19848, n19849, n19850,
         n19851, n19852, n19853, n19854, n19855, n19856, n19857, n19858,
         n19859, n19860, n19861, n19862, n19863, n19864, n19865, n19866,
         n19867, n19868, n19869, n19870, n19871, n19872, n19873, n19874,
         n19875, n19876, n19877, n19878, n19879, n19880, n19881, n19882,
         n19883, n19884, n19885, n19886, n19887, n19888, n19889, n19890,
         n19891, n19892, n19893, n19894, n19895, n19896, n19897, n19898,
         n19899, n19900, n19901, n19902, n19903, n19904, n19905, n19906,
         n19907, n19908, n19909, n19910, n19911, n19912, n19913, n19914,
         n19915, n19916, n19917, n19918, n19919, n19920, n19921, n19922,
         n19923, n19924, n19925, n19926, n19927, n19928, n19929, n19930,
         n19931, n19932, n19933, n19934, n19935, n19936, n19937, n19938,
         n19939, n19940, n19941, n19942, n19943, n19944, n19945, n19946,
         n19947, n19948, n19949, n19950, n19951, n19952, n19953, n19954,
         n19955, n19956, n19957, n19958, n19959, n19960, n19961, n19962,
         n19963, n19964, n19965, n19966, n19967, n19968, n19969, n19970,
         n19971, n19972, n19973, n19974, n19975, n19976, n19977, n19978,
         n19979, n19980, n19981, n19982, n19983, n19984, n19985, n19986,
         n19987, n19988, n19989, n19990, n19991, n19992, n19993, n19994,
         n19995, n19996, n19997, n19998, n19999, n20000, n20001, n20002,
         n20003, n20004, n20005, n20006, n20007, n20008, n20009, n20010,
         n20011, n20012, n20013, n20014, n20015, n20016, n20017, n20018,
         n20019, n20020, n20021, n20022, n20023, n20024, n20025, n20026,
         n20027, n20028, n20029, n20030, n20031, n20032, n20033, n20034,
         n20035, n20036, n20037, n20038, n20039, n20040, n20041, n20042,
         n20043, n20044, n20045, n20046, n20047, n20048, n20049, n20050,
         n20051, n20052, n20053, n20054, n20055, n20056, n20057, n20058,
         n20059, n20060, n20061, n20062, n20063, n20064, n20065, n20066,
         n20067, n20068, n20069, n20070, n20071, n20072, n20073, n20074,
         n20075, n20076, n20077, n20078, n20079, n20080, n20081, n20082,
         n20083, n20084, n20085, n20086, n20087, n20088, n20089, n20090,
         n20091, n20092, n20093, n20094, n20095, n20096, n20097, n20098,
         n20099, n20100, n20101, n20102, n20103, n20104, n20105, n20106,
         n20107, n20108, n20109, n20110, n20111, n20112, n20113, n20114,
         n20115, n20116, n20117, n20118, n20119, n20120, n20121, n20122,
         n20123, n20124, n20125, n20126, n20127, n20128, n20129, n20130,
         n20131, n20132, n20133, n20134, n20135, n20136, n20137, n20138,
         n20139, n20140, n20141, n20142, n20143, n20144, n20145, n20146,
         n20147, n20148, n20149, n20150, n20151, n20152, n20153, n20154,
         n20155, n20156, n20157, n20158, n20159, n20160, n20161, n20162,
         n20163, n20164, n20165, n20166, n20167, n20168, n20169, n20170,
         n20171, n20172, n20173, n20174, n20175, n20176, n20177, n20178,
         n20179, n20180, n20181, n20182, n20183, n20184, n20185, n20186,
         n20187, n20188, n20189, n20190, n20191, n20192, n20193, n20194,
         n20195, n20196, n20197, n20198, n20199, n20200, n20201, n20202,
         n20203, n20204, n20205, n20206, n20207, n20208, n20209, n20210,
         n20211, n20212, n20213, n20214, n20215, n20216, n20217, n20218,
         n20219, n20220, n20221, n20222, n20223, n20224, n20225, n20226,
         n20227, n20228, n20229, n20230, n20231, n20232, n20233, n20234,
         n20235, n20236, n20237, n20238, n20239, n20240, n20241, n20242,
         n20243, n20244, n20245, n20246, n20247, n20248, n20249, n20250,
         n20251, n20252, n20253, n20254, n20255, n20256, n20257, n20258,
         n20259, n20260, n20261, n20262, n20263, n20264, n20265, n20266,
         n20267, n20268, n20269, n20270, n20271, n20272, n20273, n20274,
         n20275, n20276, n20277, n20278, n20279, n20280, n20281, n20282,
         n20283, n20284, n20285, n20286, n20287, n20288, n20289, n20290,
         n20291, n20292, n20293, n20294, n20295, n20296, n20297, n20298,
         n20299, n20300, n20301, n20302, n20303, n20304, n20305, n20306,
         n20307, n20308, n20309, n20310, n20311, n20312, n20313, n20314,
         n20315, n20316, n20317, n20318, n20319, n20320, n20321, n20322,
         n20323, n20324, n20325, n20326, n20327, n20328, n20329, n20330,
         n20331, n20332, n20333, n20334, n20335, n20336, n20337, n20338,
         n20339, n20340, n20341, n20342, n20343, n20344, n20345, n20346,
         n20347, n20348, n20349, n20350, n20351, n20352, n20353, n20354,
         n20355, n20356, n20357, n20358, n20359, n20360, n20361, n20362,
         n20363, n20364, n20365, n20366, n20367, n20368, n20369, n20370,
         n20371, n20372, n20373, n20374, n20375, n20376, n20377, n20378,
         n20379, n20380, n20381, n20382, n20383, n20384, n20385, n20386,
         n20387, n20388, n20389, n20390, n20391, n20392, n20393, n20394,
         n20395, n20396, n20397, n20398, n20399, n20400, n20401, n20402,
         n20403, n20404, n20405, n20406, n20407, n20408, n20409, n20410,
         n20411, n20412, n20413, n20414, n20415, n20416, n20417, n20418,
         n20419, n20420, n20421, n20422, n20423, n20424, n20425, n20426,
         n20427, n20428, n20429, n20430, n20431, n20432, n20433, n20434,
         n20435, n20436, n20437, n20438, n20439, n20440, n20441, n20442,
         n20443, n20444, n20445, n20446, n20447, n20448, n20449, n20450,
         n20451, n20452, n20453, n20454, n20455, n20456, n20457, n20458,
         n20459, n20460, n20461, n20462, n20463, n20464, n20465, n20466,
         n20467, n20468, n20469, n20470, n20471, n20472, n20473, n20474,
         n20475, n20476, n20477, n20478, n20479, n20480, n20481, n20482,
         n20483, n20484, n20485, n20486, n20487, n20488, n20489, n20490,
         n20491, n20492, n20493, n20494, n20495, n20496, n20497, n20498,
         n20499, n20500, n20501, n20502, n20503, n20504, n20505, n20506,
         n20507, n20508, n20509, n20510, n20511, n20512, n20513, n20514,
         n20515, n20516, n20517, n20518, n20519, n20520, n20521, n20522,
         n20523, n20524, n20525, n20526, n20527, n20528, n20529, n20530,
         n20531, n20532, n20533, n20534, n20535, n20536, n20537, n20538,
         n20539, n20540, n20541, n20542, n20543, n20544, n20545, n20546,
         n20547, n20548, n20549, n20550, n20551, n20552, n20553, n20554,
         n20555, n20556, n20557, n20558, n20559, n20560, n20561, n20562,
         n20563, n20564, n20565, n20566, n20567, n20568, n20569, n20570,
         n20571, n20572, n20573, n20574, n20575, n20576, n20577, n20578,
         n20579, n20580, n20581, n20582, n20583, n20584, n20585, n20586,
         n20587, n20588, n20589, n20590, n20591, n20592, n20593, n20594,
         n20595, n20596, n20597, n20598, n20599, n20600, n20601, n20602,
         n20603, n20604, n20605, n20606, n20607, n20608, n20609, n20610,
         n20611, n20612, n20613, n20614, n20615, n20616, n20617, n20618,
         n20619, n20620, n20621, n20622, n20623, n20624, n20625, n20626,
         n20627, n20628, n20629, n20630, n20631, n20632, n20633, n20634,
         n20635, n20636, n20637, n20638, n20639, n20640, n20641, n20642,
         n20643, n20644, n20645, n20646, n20647, n20648, n20649, n20650,
         n20651, n20652, n20653, n20654, n20655, n20656, n20657, n20658,
         n20659, n20660, n20661, n20662, n20663, n20664, n20665, n20666,
         n20667, n20668, n20669, n20670, n20671, n20672, n20673, n20674,
         n20675, n20676, n20677, n20678, n20679, n20680, n20681, n20682,
         n20683, n20684, n20685, n20686, n20687, n20688, n20689, n20690,
         n20691, n20692, n20693, n20694, n20695, n20696, n20697, n20698,
         n20699, n20700, n20701, n20702, n20703, n20704, n20705, n20706,
         n20707, n20708, n20709, n20710, n20711, n20712, n20713, n20714,
         n20715, n20716, n20717, n20718, n20719, n20720, n20721, n20722,
         n20723, n20724, n20725, n20726, n20727, n20728, n20729, n20730,
         n20731, n20732, n20733, n20734, n20735, n20736, n20737, n20738,
         n20739, n20740, n20741, n20742, n20743, n20744, n20745, n20746,
         n20747, n20748, n20749, n20750, n20751, n20752, n20753, n20754,
         n20755, n20756, n20757, n20758, n20759, n20760, n20761, n20762,
         n20763, n20764, n20765, n20766, n20767, n20768, n20769, n20770,
         n20771, n20772, n20773, n20774, n20775, n20776, n20777, n20778,
         n20779, n20780, n20781, n20782, n20783, n20784, n20785, n20786,
         n20787, n20788, n20789, n20790, n20791, n20792, n20793, n20794,
         n20795, n20796, n20797, n20798, n20799, n20800, n20801, n20802,
         n20803, n20804, n20805, n20806, n20807, n20808, n20809, n20810,
         n20811, n20812, n20813, n20814, n20815, n20816, n20817, n20818,
         n20819, n20820, n20821, n20822, n20823, n20824, n20825, n20826,
         n20827, n20828, n20829, n20830, n20831, n20832, n20833, n20834,
         n20835, n20836, n20837, n20838, n20839, n20840, n20841, n20842,
         n20843, n20844, n20845, n20846, n20847, n20848, n20849, n20850,
         n20851, n20852, n20853, n20854, n20855, n20856, n20857, n20858,
         n20859, n20860, n20861, n20862, n20863, n20864, n20865, n20866,
         n20867, n20868, n20869, n20870, n20871, n20872, n20873, n20874,
         n20875, n20876, n20877, n20878, n20879, n20880, n20881, n20882,
         n20883, n20884, n20885, n20886, n20887, n20888, n20889, n20890,
         n20891, n20892, n20893, n20894, n20895, n20896, n20897, n20898,
         n20899, n20900, n20901, n20902, n20903, n20904, n20905, n20906,
         n20907, n20908, n20909, n20910, n20911, n20912, n20913, n20914,
         n20915, n20916, n20917, n20918, n20919, n20920, n20921, n20922,
         n20923, n20924, n20925, n20926, n20927, n20928, n20929, n20930,
         n20931, n20932, n20933, n20934, n20935, n20936, n20937, n20938,
         n20939, n20940, n20941, n20942, n20943, n20944, n20945, n20946,
         n20947, n20948, n20949, n20950, n20951, n20952, n20953, n20954,
         n20955, n20956, n20957, n20958, n20959, n20960, n20961, n20962,
         n20963, n20964, n20965, n20966, n20967, n20968, n20969, n20970,
         n20971, n20972, n20973, n20974, n20975, n20976, n20977, n20978,
         n20979, n20980, n20981, n20982, n20983, n20984, n20985, n20986,
         n20987, n20988, n20989, n20990, n20991, n20992, n20993, n20994,
         n20995, n20996, n20997, n20998, n20999, n21000, n21001, n21002,
         n21003, n21004, n21005, n21006, n21007, n21008, n21009, n21010,
         n21011, n21012, n21013, n21014, n21015, n21016, n21017, n21018,
         n21019, n21020, n21021, n21022, n21023, n21024, n21025, n21026,
         n21027, n21028, n21029, n21030, n21031, n21032, n21033, n21034,
         n21035, n21036, n21037, n21038, n21039, n21040, n21041, n21042,
         n21043, n21044, n21045, n21046, n21047, n21048, n21049, n21050,
         n21051, n21052, n21053, n21054, n21055, n21056, n21057, n21058,
         n21059, n21060, n21061, n21062, n21063, n21064, n21065, n21066,
         n21067, n21068, n21069, n21070, n21071, n21072, n21073, n21074,
         n21075, n21076, n21077, n21078, n21079, n21080, n21081, n21082,
         n21083, n21084, n21085, n21086, n21087, n21088, n21089, n21090,
         n21091, n21092, n21093, n21094, n21095, n21096, n21097, n21098,
         n21099, n21100, n21101, n21102, n21103, n21104, n21105, n21106,
         n21107, n21108, n21109, n21110, n21111, n21112, n21113, n21114,
         n21115, n21116, n21117, n21118, n21119, n21120, n21121, n21122,
         n21123, n21124, n21125, n21126, n21127, n21128, n21129, n21130,
         n21131, n21132, n21133, n21134, n21135, n21136, n21137, n21138,
         n21139, n21140, n21141, n21142, n21143, n21144, n21145, n21146,
         n21147, n21148, n21149, n21150, n21151, n21152, n21153, n21154,
         n21155, n21156, n21157, n21158, n21159, n21160, n21161, n21162,
         n21163, n21164, n21165, n21166, n21167, n21168, n21169, n21170,
         n21171, n21172, n21173, n21174, n21175, n21176, n21177, n21178,
         n21179, n21180, n21181, n21182, n21183, n21184, n21185, n21186,
         n21187, n21188, n21189, n21190, n21191, n21192, n21193, n21194,
         n21195, n21196, n21197, n21198, n21199, n21200, n21201, n21202,
         n21203, n21204, n21205, n21206, n21207, n21208, n21209, n21210,
         n21211, n21212, n21213, n21214, n21215, n21216, n21217, n21218,
         n21219, n21220, n21221, n21222, n21223, n21224, n21225, n21226,
         n21227, n21228, n21229, n21230, n21231, n21232, n21233, n21234,
         n21235, n21236, n21237, n21238, n21239, n21240, n21241, n21242,
         n21243, n21244, n21245, n21246, n21247, n21248, n21249, n21250,
         n21251, n21252, n21253, n21254, n21255, n21256, n21257, n21258,
         n21259, n21260, n21261, n21262, n21263, n21264, n21265, n21266,
         n21267, n21268, n21269, n21270, n21271, n21272, n21273, n21274,
         n21275, n21276, n21277, n21278, n21279, n21280, n21281, n21282,
         n21283, n21284, n21285, n21286, n21287, n21288, n21289, n21290,
         n21291, n21292, n21293, n21294, n21295, n21296, n21297, n21298,
         n21299, n21300, n21301, n21302, n21303, n21304, n21305, n21306,
         n21307, n21308, n21309, n21310, n21311, n21312, n21313, n21314,
         n21315, n21316, n21317, n21318, n21319, n21320, n21321, n21322,
         n21323, n21324, n21325, n21326, n21327, n21328, n21329, n21330,
         n21331, n21332, n21333, n21334, n21335, n21336, n21337, n21338,
         n21339, n21340, n21341, n21342, n21343, n21344, n21345, n21346,
         n21347, n21348, n21349, n21350, n21351, n21352, n21353, n21354,
         n21355, n21356, n21357, n21358, n21359, n21360, n21361, n21362,
         n21363, n21364, n21365, n21366, n21367, n21368, n21369, n21370,
         n21371, n21372, n21373, n21374, n21375, n21376, n21377, n21378,
         n21379, n21380, n21381, n21382, n21383, n21384, n21385, n21386,
         n21387, n21388, n21389, n21390, n21391, n21392, n21393, n21394,
         n21395, n21396, n21397, n21398, n21399, n21400, n21401, n21402,
         n21403, n21404, n21405, n21406, n21407, n21408, n21409, n21410,
         n21411, n21412, n21413, n21414, n21415, n21416, n21417, n21418,
         n21419, n21420, n21421, n21422, n21423, n21424, n21425, n21426,
         n21427, n21428, n21429, n21430, n21431, n21432, n21433, n21434,
         n21435, n21436, n21437, n21438, n21439, n21440, n21441, n21442,
         n21443, n21444, n21445, n21446, n21447, n21448, n21449, n21450,
         n21451, n21452, n21453, n21454, n21455, n21456, n21457, n21458,
         n21459, n21460, n21461, n21462, n21463, n21464, n21465, n21466,
         n21467, n21468, n21469, n21470, n21471, n21472, n21473, n21474,
         n21475, n21476, n21477, n21478, n21479, n21480, n21481, n21482,
         n21483, n21484, n21485, n21486, n21487, n21488, n21489, n21490,
         n21491, n21492, n21493, n21494, n21495, n21496, n21497, n21498,
         n21499, n21500, n21501, n21502, n21503, n21504, n21505, n21506,
         n21507, n21508, n21509, n21510, n21511, n21512, n21513, n21514,
         n21515, n21516, n21517, n21518, n21519, n21520, n21521, n21522,
         n21523, n21524, n21525, n21526, n21527, n21528, n21529, n21530,
         n21531, n21532, n21533, n21534, n21535, n21536, n21537, n21538,
         n21539, n21540, n21541, n21542, n21543, n21544, n21545, n21546,
         n21547, n21548, n21549, n21550, n21551, n21552, n21553, n21554,
         n21555, n21556, n21557, n21558, n21559, n21560, n21561, n21562,
         n21563, n21564, n21565, n21566, n21567, n21568, n21569, n21570,
         n21571, n21572, n21573, n21574, n21575, n21576, n21577, n21578,
         n21579, n21580, n21581, n21582, n21583, n21584, n21585, n21586,
         n21587, n21588, n21589, n21590, n21591, n21592, n21593, n21594,
         n21595, n21596, n21597, n21598, n21599, n21600, n21601, n21602,
         n21603, n21604, n21605, n21606, n21607, n21608, n21609, n21610,
         n21611, n21612, n21613, n21614, n21615, n21616, n21617, n21618,
         n21619, n21620, n21621, n21622, n21623, n21624, n21625, n21626,
         n21627, n21628, n21629, n21630, n21631, n21632, n21633, n21634,
         n21635, n21636, n21637, n21638, n21639, n21640, n21641, n21642,
         n21643, n21644, n21645, n21646, n21647, n21648, n21649, n21650,
         n21651, n21652, n21653, n21654, n21655, n21656, n21657, n21658,
         n21659, n21660, n21661, n21662, n21663, n21664, n21665, n21666,
         n21667, n21668, n21669, n21670, n21671, n21672, n21673, n21674,
         n21675, n21676, n21677, n21678, n21679, n21680, n21681, n21682,
         n21683, n21684, n21685, n21686, n21687, n21688, n21689, n21690,
         n21691, n21692, n21693, n21694, n21695, n21696, n21697, n21698,
         n21699, n21700, n21701, n21702, n21703, n21704, n21705, n21706,
         n21707, n21708, n21709, n21710, n21711, n21712, n21713, n21714,
         n21715, n21716, n21717, n21718, n21719, n21720, n21721, n21722,
         n21723, n21724, n21725, n21726, n21727, n21728, n21729, n21730,
         n21731, n21732, n21733, n21734, n21735, n21736, n21737, n21738,
         n21739, n21740, n21741, n21742, n21743, n21744, n21745, n21746,
         n21747, n21748, n21749, n21750, n21751, n21752, n21753, n21754,
         n21755, n21756, n21757, n21758, n21759, n21760, n21761, n21762,
         n21763, n21764, n21765, n21766, n21767, n21768, n21769, n21770,
         n21771, n21772, n21773, n21774, n21775, n21776, n21777, n21778,
         n21779, n21780, n21781, n21782, n21783, n21784, n21785, n21786,
         n21787, n21788, n21789, n21790, n21791, n21792, n21793, n21794,
         n21795, n21796, n21797, n21798, n21799, n21800, n21801, n21802,
         n21803, n21804, n21805, n21806, n21807, n21808, n21809, n21810,
         n21811, n21812, n21813, n21814, n21815, n21816, n21817, n21818,
         n21819, n21820, n21821, n21822, n21823, n21824, n21825, n21826,
         n21827, n21828, n21829, n21830, n21831, n21832, n21833, n21834,
         n21835, n21836, n21837, n21838, n21839, n21840, n21841, n21842,
         n21843, n21844, n21845, n21846, n21847, n21848, n21849, n21850,
         n21851, n21852, n21853, n21854, n21855, n21856, n21857, n21858,
         n21859, n21860, n21861, n21862, n21863, n21864, n21865, n21866,
         n21867, n21868, n21869, n21870, n21871, n21872, n21873, n21874,
         n21875, n21876, n21877, n21878, n21879, n21880, n21881, n21882,
         n21883, n21884, n21885, n21886, n21887, n21888, n21889, n21890,
         n21891, n21892, n21893, n21894, n21895, n21896, n21897, n21898,
         n21899, n21900, n21901, n21902, n21903, n21904, n21905, n21906,
         n21907, n21908, n21909, n21910, n21911, n21912, n21913, n21914,
         n21915, n21916, n21917, n21918, n21919, n21920, n21921, n21922,
         n21923, n21924, n21925, n21926, n21927, n21928, n21929, n21930,
         n21931, n21932, n21933, n21934, n21935, n21936, n21937, n21938,
         n21939;

  INV_X1 U11120 ( .A(n21098), .ZN(n15507) );
  AND2_X1 U11121 ( .A1(n21233), .A2(n21267), .ZN(n21226) );
  AND2_X1 U11122 ( .A1(n21233), .A2(n21202), .ZN(n21262) );
  INV_X1 U11123 ( .A(n16210), .ZN(n17999) );
  CLKBUF_X1 U11124 ( .A(n14253), .Z(n9682) );
  NAND2_X1 U11125 ( .A1(n10054), .A2(n10055), .ZN(n10112) );
  OR2_X1 U11126 ( .A1(n21016), .A2(n15153), .ZN(n20970) );
  OR2_X1 U11127 ( .A1(n13023), .A2(n13012), .ZN(n16043) );
  OR3_X1 U11128 ( .A1(n13473), .A2(n13472), .A3(n21119), .ZN(n15656) );
  AND2_X1 U11129 ( .A1(n14365), .A2(n14368), .ZN(n15792) );
  NAND2_X1 U11130 ( .A1(n10305), .A2(n10304), .ZN(n16065) );
  NAND2_X1 U11131 ( .A1(n15074), .A2(n10524), .ZN(n15011) );
  INV_X1 U11132 ( .A(n20164), .ZN(n20144) );
  AND2_X1 U11133 ( .A1(n10806), .A2(n10820), .ZN(n17616) );
  OR2_X1 U11134 ( .A1(n14362), .A2(n10537), .ZN(n10536) );
  INV_X2 U11135 ( .A(n12775), .ZN(n11243) );
  NAND2_X1 U11136 ( .A1(n10798), .A2(n10801), .ZN(n10869) );
  NAND2_X1 U11137 ( .A1(n13353), .A2(n19580), .ZN(n11691) );
  BUF_X1 U11138 ( .A(n14068), .Z(n20281) );
  OR2_X1 U11139 ( .A1(n12638), .A2(n12726), .ZN(n12725) );
  INV_X1 U11140 ( .A(n11712), .ZN(n19565) );
  INV_X1 U11141 ( .A(n11223), .ZN(n11261) );
  CLKBUF_X2 U11142 ( .A(n12650), .Z(n12714) );
  INV_X1 U11143 ( .A(n10372), .ZN(n19583) );
  CLKBUF_X2 U11144 ( .A(n12075), .Z(n12395) );
  CLKBUF_X2 U11145 ( .A(n11996), .Z(n9689) );
  CLKBUF_X2 U11146 ( .A(n11792), .Z(n9707) );
  CLKBUF_X2 U11147 ( .A(n11797), .Z(n12488) );
  CLKBUF_X2 U11148 ( .A(n11837), .Z(n12526) );
  CLKBUF_X2 U11149 ( .A(n11936), .Z(n9711) );
  CLKBUF_X2 U11150 ( .A(n11849), .Z(n12527) );
  CLKBUF_X1 U11152 ( .A(n11995), .Z(n12544) );
  CLKBUF_X2 U11153 ( .A(n11823), .Z(n9690) );
  AND2_X1 U11154 ( .A1(n10753), .A2(n17986), .ZN(n9892) );
  NOR2_X1 U11155 ( .A1(n10514), .A2(n10358), .ZN(n15147) );
  AND2_X2 U11156 ( .A1(n16448), .A2(n10265), .ZN(n16438) );
  CLKBUF_X1 U11157 ( .A(n13734), .Z(n18703) );
  NAND2_X1 U11158 ( .A1(n11472), .A2(n11009), .ZN(n11471) );
  CLKBUF_X1 U11159 ( .A(n10733), .Z(n17537) );
  CLKBUF_X3 U11160 ( .A(n10809), .Z(n9710) );
  AND2_X2 U11161 ( .A1(n10696), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11190) );
  CLKBUF_X2 U11162 ( .A(n13273), .Z(n9681) );
  AND2_X2 U11163 ( .A1(n16593), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10841) );
  AND2_X1 U11164 ( .A1(n10731), .A2(n10720), .ZN(n10345) );
  AND2_X1 U11165 ( .A1(n9959), .A2(n9958), .ZN(n10732) );
  AND2_X1 U11166 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14720) );
  NAND2_X2 U11167 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n14732) );
  AND2_X1 U11168 ( .A1(n10320), .A2(n13950), .ZN(n11824) );
  INV_X1 U11169 ( .A(n11928), .ZN(n11995) );
  AND2_X2 U11170 ( .A1(n11743), .A2(n11742), .ZN(n11996) );
  NAND2_X1 U11171 ( .A1(n13949), .A2(n14443), .ZN(n11950) );
  AND2_X2 U11172 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13950) );
  AND2_X2 U11173 ( .A1(n10265), .A2(n11000), .ZN(n9685) );
  NAND3_X1 U11174 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n17480) );
  AND2_X1 U11175 ( .A1(n13603), .A2(n9710), .ZN(n9676) );
  OAI22_X1 U11176 ( .A1(n10869), .A2(n10799), .B1(n20740), .B2(n10803), .ZN(
        n9894) );
  AND2_X1 U11177 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n14443) );
  NOR2_X1 U11178 ( .A1(n10743), .A2(n10724), .ZN(n10758) );
  INV_X1 U11179 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14023) );
  NAND2_X1 U11180 ( .A1(n11011), .A2(n10733), .ZN(n9971) );
  NAND2_X1 U11181 ( .A1(n12968), .A2(n10722), .ZN(n10740) );
  INV_X1 U11182 ( .A(n11950), .ZN(n9691) );
  CLKBUF_X2 U11183 ( .A(n11824), .Z(n9713) );
  INV_X1 U11184 ( .A(n12614), .ZN(n12594) );
  AND2_X2 U11185 ( .A1(n10265), .A2(n11000), .ZN(n16613) );
  OR2_X1 U11187 ( .A1(n10816), .A2(n14079), .ZN(n10954) );
  INV_X1 U11188 ( .A(n18704), .ZN(n18728) );
  INV_X1 U11189 ( .A(n9815), .ZN(n12456) );
  NAND2_X1 U11190 ( .A1(n15742), .A2(n21117), .ZN(n21137) );
  NAND2_X1 U11191 ( .A1(n10556), .A2(n11960), .ZN(n10323) );
  OR2_X1 U11192 ( .A1(n11064), .A2(n13022), .ZN(n13001) );
  OR2_X1 U11194 ( .A1(n10819), .A2(n10806), .ZN(n17544) );
  AND2_X1 U11195 ( .A1(n10806), .A2(n10807), .ZN(n20504) );
  NAND2_X1 U11196 ( .A1(n10173), .A2(n14079), .ZN(n20606) );
  INV_X2 U11197 ( .A(n13146), .ZN(n10358) );
  NOR2_X2 U11198 ( .A1(n15092), .A2(n15072), .ZN(n15074) );
  NAND2_X1 U11199 ( .A1(n11110), .A2(n13001), .ZN(n11113) );
  NAND2_X1 U11201 ( .A1(n11163), .A2(n11162), .ZN(n17651) );
  INV_X1 U11202 ( .A(n11543), .ZN(n14596) );
  AND4_X1 U11203 ( .A1(n13192), .A2(n13191), .A3(n13190), .A4(n13189), .ZN(
        n13197) );
  INV_X1 U11204 ( .A(n13963), .ZN(n19571) );
  INV_X1 U11205 ( .A(n21003), .ZN(n21024) );
  AND2_X1 U11206 ( .A1(n15134), .A2(n15119), .ZN(n15121) );
  AND2_X2 U11207 ( .A1(n14864), .A2(n14865), .ZN(n13150) );
  INV_X1 U11208 ( .A(n10514), .ZN(n13450) );
  NAND2_X1 U11209 ( .A1(n14261), .A2(n12102), .ZN(n14412) );
  INV_X1 U11210 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n20750) );
  INV_X1 U11211 ( .A(n12943), .ZN(n16336) );
  INV_X1 U11212 ( .A(n14068), .ZN(n14079) );
  NAND2_X1 U11213 ( .A1(n16018), .A2(n16019), .ZN(n16004) );
  INV_X1 U11214 ( .A(n14033), .ZN(n10091) );
  OR2_X1 U11215 ( .A1(n17184), .A2(n10412), .ZN(n9805) );
  NOR2_X2 U11216 ( .A1(n20439), .A2(n20666), .ZN(n20430) );
  NOR2_X1 U11217 ( .A1(n20476), .A2(n20666), .ZN(n20440) );
  OR2_X1 U11218 ( .A1(n11655), .A2(n11654), .ZN(n18787) );
  INV_X1 U11219 ( .A(n18787), .ZN(n19588) );
  OR2_X1 U11220 ( .A1(n13184), .A2(n13183), .ZN(n13368) );
  INV_X1 U11221 ( .A(n19281), .ZN(n19243) );
  AND2_X1 U11222 ( .A1(n10021), .A2(n13549), .ZN(n17742) );
  OR2_X1 U11223 ( .A1(n13150), .A2(n10279), .ZN(n15322) );
  OR2_X1 U11224 ( .A1(n14129), .A2(n15950), .ZN(n20943) );
  INV_X1 U11225 ( .A(n20316), .ZN(n20348) );
  INV_X1 U11226 ( .A(n20597), .ZN(n20633) );
  NAND2_X1 U11227 ( .A1(n18192), .A2(n20024), .ZN(n18193) );
  INV_X1 U11228 ( .A(n18551), .ZN(n18574) );
  XOR2_X1 U11229 ( .A(n10436), .B(n16985), .Z(n9677) );
  OR2_X1 U11230 ( .A1(n16065), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n9678) );
  INV_X1 U11231 ( .A(n11594), .ZN(n9704) );
  INV_X2 U11232 ( .A(n10618), .ZN(n10267) );
  NOR2_X4 U11233 ( .A1(n14992), .A2(n9745), .ZN(n14913) );
  NAND3_X1 U11234 ( .A1(n11465), .A2(n9892), .A3(n17682), .ZN(n10315) );
  AND2_X1 U11235 ( .A1(n11000), .A2(n17469), .ZN(n9679) );
  AND2_X1 U11236 ( .A1(n11000), .A2(n17469), .ZN(n9680) );
  AND2_X2 U11237 ( .A1(n11000), .A2(n17469), .ZN(n9705) );
  AND2_X2 U11238 ( .A1(n11000), .A2(n17469), .ZN(n16445) );
  NAND2_X1 U11239 ( .A1(n14764), .A2(n10252), .ZN(n13273) );
  OR2_X2 U11240 ( .A1(n15519), .A2(n21139), .ZN(n9941) );
  AOI21_X1 U11241 ( .B1(n14322), .B2(n14156), .A(n20047), .ZN(n14253) );
  NAND2_X2 U11242 ( .A1(n14333), .A2(n11560), .ZN(n14603) );
  INV_X1 U11243 ( .A(n19271), .ZN(n19237) );
  BUF_X2 U11244 ( .A(n13734), .Z(n9683) );
  AND2_X1 U11245 ( .A1(n11554), .A2(n14719), .ZN(n13734) );
  AND2_X1 U11246 ( .A1(n10265), .A2(n11000), .ZN(n9684) );
  CLKBUF_X3 U11247 ( .A(n16484), .Z(n16447) );
  CLKBUF_X3 U11248 ( .A(n16484), .Z(n16593) );
  NOR3_X2 U11249 ( .A1(n17178), .A2(n13057), .A3(n17188), .ZN(n17163) );
  AND2_X4 U11250 ( .A1(n17481), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n16446) );
  CLKBUF_X1 U11251 ( .A(n16446), .Z(n9708) );
  AND2_X4 U11253 ( .A1(n14731), .A2(n11556), .ZN(n13279) );
  NAND2_X2 U11254 ( .A1(n10070), .A2(n17667), .ZN(n17986) );
  AND2_X1 U11255 ( .A1(n16896), .A2(n10319), .ZN(n17195) );
  AOI211_X1 U11256 ( .C1(n20277), .C2(n17305), .A(n17304), .B(n17303), .ZN(
        n17308) );
  NAND2_X1 U11257 ( .A1(n17021), .A2(n10402), .ZN(n17295) );
  INV_X2 U11258 ( .A(n15317), .ZN(n10370) );
  NOR2_X1 U11259 ( .A1(n13027), .A2(n9858), .ZN(n16940) );
  NAND3_X1 U11260 ( .A1(n10329), .A2(n16913), .A3(n10330), .ZN(n16917) );
  OR2_X1 U11261 ( .A1(n16637), .A2(n16636), .ZN(n10467) );
  INV_X1 U11262 ( .A(n11511), .ZN(n9686) );
  AND2_X1 U11263 ( .A1(n17789), .A2(n19030), .ZN(n19017) );
  INV_X1 U11264 ( .A(n11516), .ZN(n9687) );
  INV_X4 U11265 ( .A(n15394), .ZN(n10056) );
  NAND2_X1 U11266 ( .A1(n14229), .A2(n14285), .ZN(n20535) );
  NOR2_X2 U11267 ( .A1(n19385), .A2(n19290), .ZN(n19032) );
  BUF_X4 U11268 ( .A(n13139), .Z(n9688) );
  AND3_X1 U11269 ( .A1(n9876), .A2(n10366), .A3(n9806), .ZN(n10365) );
  OR3_X1 U11270 ( .A1(n21611), .A2(n15496), .A3(n12633), .ZN(n15158) );
  NAND2_X1 U11271 ( .A1(n13430), .A2(n13429), .ZN(n13469) );
  INV_X1 U11272 ( .A(n20021), .ZN(n19543) );
  NAND2_X1 U11273 ( .A1(n10257), .A2(n10255), .ZN(n13314) );
  NOR2_X1 U11274 ( .A1(n11066), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n11080) );
  INV_X4 U11275 ( .A(n11385), .ZN(n12840) );
  OR2_X1 U11276 ( .A1(n11056), .A2(n10596), .ZN(n11064) );
  NAND2_X1 U11277 ( .A1(n13294), .A2(n10016), .ZN(n13295) );
  AND2_X1 U11278 ( .A1(n11686), .A2(n13356), .ZN(n13353) );
  AND2_X1 U11279 ( .A1(n11927), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12568) );
  INV_X4 U11280 ( .A(n13010), .ZN(n11012) );
  NAND3_X1 U11281 ( .A1(n10728), .A2(n9991), .A3(n10721), .ZN(n10750) );
  AND2_X1 U11282 ( .A1(n16743), .A2(n14026), .ZN(n11223) );
  OR2_X2 U11283 ( .A1(n11581), .A2(n11580), .ZN(n20150) );
  CLKBUF_X2 U11284 ( .A(n11873), .Z(n14403) );
  NOR2_X1 U11285 ( .A1(n9696), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n14026) );
  OR2_X1 U11286 ( .A1(n11759), .A2(n11758), .ZN(n14385) );
  INV_X1 U11288 ( .A(n11212), .ZN(n10809) );
  AND2_X1 U11289 ( .A1(n9773), .A2(n11782), .ZN(n11871) );
  INV_X4 U11290 ( .A(n14603), .ZN(n18739) );
  BUF_X2 U11291 ( .A(n11818), .Z(n12550) );
  BUF_X2 U11292 ( .A(n12131), .Z(n12378) );
  INV_X2 U11293 ( .A(n12502), .ZN(n12019) );
  AND2_X1 U11294 ( .A1(n11734), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11743) );
  INV_X4 U11296 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10252) );
  NOR2_X1 U11297 ( .A1(n10005), .A2(n11524), .ZN(n11525) );
  AOI21_X1 U11298 ( .B1(n20267), .B2(n17195), .A(n17194), .ZN(n17196) );
  NOR2_X1 U11299 ( .A1(n9761), .A2(n14786), .ZN(n14787) );
  AND2_X1 U11300 ( .A1(n12867), .A2(n12866), .ZN(n10515) );
  NAND2_X1 U11301 ( .A1(n9924), .A2(n13032), .ZN(n13058) );
  OAI21_X1 U11302 ( .B1(n16993), .B2(n10163), .A(n10162), .ZN(n10161) );
  AND2_X1 U11303 ( .A1(n9955), .A2(n9954), .ZN(n17324) );
  OAI211_X1 U11304 ( .C1(n17021), .C2(n17385), .A(n10239), .B(n10176), .ZN(
        n17380) );
  XNOR2_X1 U11305 ( .A(n9934), .B(n12871), .ZN(n13166) );
  XNOR2_X1 U11306 ( .A(n16886), .B(n13036), .ZN(n16881) );
  OAI21_X1 U11307 ( .B1(n15322), .B2(n15511), .A(n10278), .ZN(n10277) );
  OAI21_X1 U11308 ( .B1(n17021), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n17066), .ZN(n17404) );
  NAND2_X1 U11309 ( .A1(n16976), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n16969) );
  NAND2_X1 U11310 ( .A1(n16905), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16896) );
  NAND2_X1 U11311 ( .A1(n10235), .A2(n13414), .ZN(n13415) );
  NAND2_X1 U11312 ( .A1(n16940), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n16923) );
  NAND2_X1 U11313 ( .A1(n16944), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n16943) );
  INV_X1 U11314 ( .A(n16940), .ZN(n10072) );
  NAND2_X1 U11315 ( .A1(n10094), .A2(n10415), .ZN(n13478) );
  AND2_X1 U11316 ( .A1(n10467), .A2(n9988), .ZN(n16771) );
  AND2_X1 U11317 ( .A1(n10464), .A2(n10463), .ZN(n16623) );
  AND2_X1 U11318 ( .A1(n15054), .A2(n15033), .ZN(n15034) );
  NAND2_X1 U11319 ( .A1(n13003), .A2(n16927), .ZN(n10330) );
  AND2_X1 U11320 ( .A1(n17171), .A2(n17170), .ZN(n17174) );
  AND2_X1 U11321 ( .A1(n15326), .A2(n10105), .ZN(n15302) );
  NAND2_X1 U11322 ( .A1(n15326), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n13411) );
  INV_X1 U11323 ( .A(n16633), .ZN(n17183) );
  AOI211_X1 U11324 ( .C1(n16633), .C2(n16354), .A(n16016), .B(n16015), .ZN(
        n16017) );
  NOR2_X1 U11325 ( .A1(n15987), .A2(n12967), .ZN(n12845) );
  NAND2_X1 U11326 ( .A1(n10050), .A2(n10051), .ZN(n15326) );
  OR2_X1 U11327 ( .A1(n16038), .A2(n16037), .ZN(n17205) );
  INV_X1 U11328 ( .A(n10293), .ZN(n10619) );
  OAI21_X1 U11329 ( .B1(n9869), .B2(n9870), .A(n9866), .ZN(n16926) );
  NAND2_X1 U11330 ( .A1(n9874), .A2(n15646), .ZN(n10104) );
  AND2_X1 U11331 ( .A1(n10620), .A2(n17240), .ZN(n10410) );
  INV_X1 U11332 ( .A(n15425), .ZN(n15464) );
  CLKBUF_X1 U11333 ( .A(n13061), .Z(n16022) );
  NAND2_X1 U11334 ( .A1(n9947), .A2(n9945), .ZN(n10293) );
  NAND3_X1 U11335 ( .A1(n17082), .A2(n9950), .A3(n10607), .ZN(n9870) );
  CLKBUF_X1 U11336 ( .A(n16020), .Z(n16021) );
  AND2_X1 U11337 ( .A1(n10623), .A2(n17079), .ZN(n10620) );
  NAND2_X1 U11338 ( .A1(n17080), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n17082) );
  NAND2_X1 U11339 ( .A1(n9719), .A2(n15100), .ZN(n15021) );
  INV_X1 U11340 ( .A(n11513), .ZN(n10269) );
  OR2_X1 U11341 ( .A1(n16542), .A2(n16540), .ZN(n16641) );
  OAI211_X1 U11342 ( .C1(n11518), .C2(n9966), .A(n9964), .B(n9960), .ZN(n17079) );
  NAND2_X1 U11343 ( .A1(n10624), .A2(n18055), .ZN(n10623) );
  NAND2_X1 U11344 ( .A1(n9930), .A2(n17436), .ZN(n17107) );
  NAND2_X1 U11345 ( .A1(n16062), .A2(n12818), .ZN(n16052) );
  NAND2_X1 U11346 ( .A1(n9796), .A2(n10325), .ZN(n17109) );
  OAI21_X1 U11347 ( .B1(n11518), .B2(n9832), .A(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n9949) );
  NAND2_X1 U11348 ( .A1(n10363), .A2(n10395), .ZN(n15475) );
  AOI21_X1 U11349 ( .B1(n10227), .B2(n10383), .A(n10225), .ZN(n10224) );
  NAND2_X1 U11350 ( .A1(n9686), .A2(n10010), .ZN(n10011) );
  AOI21_X1 U11351 ( .B1(n10049), .B2(n10113), .A(n15394), .ZN(n10050) );
  INV_X1 U11352 ( .A(n11517), .ZN(n11518) );
  INV_X1 U11353 ( .A(n20556), .ZN(n20577) );
  NAND2_X1 U11354 ( .A1(n10270), .A2(n11516), .ZN(n10204) );
  AND2_X1 U11355 ( .A1(n16892), .A2(n13014), .ZN(n13015) );
  NOR2_X1 U11356 ( .A1(n16735), .A2(n16699), .ZN(n16736) );
  NAND3_X1 U11357 ( .A1(n12111), .A2(n14412), .A3(n14411), .ZN(n14410) );
  AOI21_X1 U11358 ( .B1(n10598), .B2(n9868), .A(n9867), .ZN(n9866) );
  NOR2_X1 U11359 ( .A1(n16004), .A2(n10574), .ZN(n16000) );
  AND2_X1 U11360 ( .A1(n10605), .A2(n9687), .ZN(n10010) );
  AOI21_X1 U11361 ( .B1(n10390), .B2(n10384), .A(n10382), .ZN(n10381) );
  NAND2_X1 U11362 ( .A1(n16410), .A2(n9989), .ZN(n16669) );
  NAND3_X1 U11363 ( .A1(n10053), .A2(n9882), .A3(n10052), .ZN(n18023) );
  XNOR2_X1 U11364 ( .A(n12961), .B(n12780), .ZN(n13033) );
  NAND2_X1 U11365 ( .A1(n20890), .A2(n17543), .ZN(n20667) );
  AND2_X1 U11366 ( .A1(n12994), .A2(n9751), .ZN(n10598) );
  AND2_X1 U11367 ( .A1(n16018), .A2(n10572), .ZN(n12961) );
  AND2_X1 U11368 ( .A1(n11058), .A2(n11251), .ZN(n10605) );
  NOR2_X1 U11369 ( .A1(n10385), .A2(n11102), .ZN(n10384) );
  NAND2_X1 U11370 ( .A1(n20890), .A2(n20914), .ZN(n20690) );
  AND2_X1 U11371 ( .A1(n17542), .A2(n20536), .ZN(n20316) );
  AND2_X1 U11372 ( .A1(n10635), .A2(n15658), .ZN(n10541) );
  NAND2_X1 U11373 ( .A1(n16367), .A2(n14286), .ZN(n14506) );
  INV_X1 U11374 ( .A(n10388), .ZN(n10385) );
  NOR2_X1 U11375 ( .A1(n16011), .A2(n11073), .ZN(n13054) );
  AND2_X1 U11376 ( .A1(n10950), .A2(n10949), .ZN(n11058) );
  NAND2_X1 U11377 ( .A1(n11439), .A2(n11438), .ZN(n16181) );
  NOR2_X1 U11378 ( .A1(n10423), .A2(n10422), .ZN(n10421) );
  NAND2_X1 U11379 ( .A1(n10987), .A2(n10986), .ZN(n11516) );
  OR2_X1 U11380 ( .A1(n10131), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15493) );
  AOI21_X1 U11381 ( .B1(n10430), .B2(n10432), .A(n10389), .ZN(n10388) );
  OAI21_X1 U11382 ( .B1(n16936), .B2(n16946), .A(n9751), .ZN(n10597) );
  OR4_X1 U11383 ( .A1(n15957), .A2(n15956), .A3(n15955), .A4(n15954), .ZN(
        n15967) );
  AND2_X1 U11384 ( .A1(n13077), .A2(n13076), .ZN(n13141) );
  NOR2_X2 U11385 ( .A1(n21355), .A2(n21354), .ZN(n21930) );
  OR2_X1 U11386 ( .A1(n13009), .A2(n13004), .ZN(n13018) );
  AOI21_X1 U11387 ( .B1(n10431), .B2(n10433), .A(n9795), .ZN(n10430) );
  OR2_X1 U11388 ( .A1(n14227), .A2(n14228), .ZN(n14229) );
  NAND2_X1 U11389 ( .A1(n10591), .A2(n13001), .ZN(n13023) );
  NOR2_X2 U11390 ( .A1(n11383), .A2(n11384), .ZN(n12763) );
  AND3_X1 U11391 ( .A1(n10802), .A2(n9908), .A3(n9907), .ZN(n10828) );
  INV_X1 U11392 ( .A(n20970), .ZN(n20968) );
  AND2_X1 U11393 ( .A1(n9897), .A2(n9895), .ZN(n9908) );
  CLKBUF_X1 U11394 ( .A(n10915), .Z(n20541) );
  AND2_X1 U11395 ( .A1(n9909), .A2(n9896), .ZN(n9895) );
  CLKBUF_X2 U11396 ( .A(n13097), .Z(n9709) );
  NAND2_X1 U11397 ( .A1(n14095), .A2(n14094), .ZN(n14262) );
  NOR2_X1 U11398 ( .A1(n18567), .A2(n18209), .ZN(n18214) );
  NAND2_X1 U11399 ( .A1(n12074), .A2(n12073), .ZN(n14095) );
  NAND2_X1 U11400 ( .A1(n14230), .A2(n10810), .ZN(n10929) );
  INV_X1 U11401 ( .A(n12980), .ZN(n10433) );
  AND2_X1 U11402 ( .A1(n11116), .A2(n11118), .ZN(n16138) );
  AND2_X1 U11403 ( .A1(n11121), .A2(n9767), .ZN(n16122) );
  NAND2_X1 U11404 ( .A1(n9910), .A2(n9901), .ZN(n20467) );
  OR2_X2 U11405 ( .A1(n10808), .A2(n16313), .ZN(n20385) );
  NOR2_X1 U11406 ( .A1(n10365), .A2(n12061), .ZN(n10537) );
  INV_X1 U11407 ( .A(n12996), .ZN(n10305) );
  NAND2_X1 U11408 ( .A1(n9910), .A2(n9906), .ZN(n20352) );
  XNOR2_X1 U11409 ( .A(n14215), .B(n14216), .ZN(n20896) );
  NAND2_X1 U11410 ( .A1(n10264), .A2(n19030), .ZN(n17815) );
  NOR2_X2 U11411 ( .A1(n18193), .A2(n20150), .ZN(n19275) );
  NAND2_X1 U11412 ( .A1(n13471), .A2(n13470), .ZN(n21119) );
  INV_X1 U11413 ( .A(n21019), .ZN(n21001) );
  NOR2_X2 U11414 ( .A1(n18193), .A2(n19568), .ZN(n19277) );
  NAND2_X1 U11415 ( .A1(n12945), .A2(n12985), .ZN(n12996) );
  OR2_X1 U11416 ( .A1(n9752), .A2(n10260), .ZN(n10264) );
  NOR2_X1 U11417 ( .A1(n18865), .A2(n18997), .ZN(n18860) );
  NAND2_X1 U11418 ( .A1(n12987), .A2(n13001), .ZN(n12945) );
  NAND2_X1 U11419 ( .A1(n15158), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15149) );
  AND2_X1 U11420 ( .A1(n15611), .A2(n15589), .ZN(n15742) );
  NAND2_X1 U11421 ( .A1(n10246), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n13387) );
  NAND2_X1 U11422 ( .A1(n12069), .A2(n10323), .ZN(n12061) );
  OR2_X1 U11423 ( .A1(n11115), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n11118) );
  NOR2_X1 U11424 ( .A1(n14040), .A2(n10804), .ZN(n10801) );
  NOR2_X1 U11425 ( .A1(n20281), .A2(n10790), .ZN(n9906) );
  NAND2_X1 U11426 ( .A1(n19204), .A2(n13315), .ZN(n13318) );
  NAND2_X1 U11427 ( .A1(n13469), .A2(n15937), .ZN(n15611) );
  OR2_X1 U11428 ( .A1(n10804), .A2(n17467), .ZN(n10808) );
  NAND2_X1 U11429 ( .A1(n13469), .A2(n13444), .ZN(n21117) );
  OR2_X1 U11430 ( .A1(n13469), .A2(n15496), .ZN(n13470) );
  NAND2_X1 U11431 ( .A1(n11113), .A2(n11112), .ZN(n11115) );
  NAND2_X1 U11432 ( .A1(n13469), .A2(n13460), .ZN(n15589) );
  AOI21_X1 U11433 ( .B1(n17467), .B2(n14217), .A(n14039), .ZN(n14074) );
  NAND2_X1 U11434 ( .A1(n14070), .A2(n14069), .ZN(n14072) );
  NAND2_X1 U11435 ( .A1(n20943), .A2(n13154), .ZN(n15504) );
  NAND2_X1 U11436 ( .A1(n14089), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13093) );
  OR2_X2 U11437 ( .A1(n15195), .A2(n14815), .ZN(n15206) );
  AND2_X1 U11438 ( .A1(n17054), .A2(n17071), .ZN(n11079) );
  NAND2_X1 U11439 ( .A1(n14044), .A2(n13732), .ZN(n21611) );
  NAND2_X1 U11440 ( .A1(n10401), .A2(n10610), .ZN(n10380) );
  OAI21_X1 U11441 ( .B1(n14364), .B2(n13092), .A(n13091), .ZN(n14089) );
  OR2_X1 U11442 ( .A1(n14129), .A2(n13428), .ZN(n13429) );
  AOI21_X1 U11443 ( .B1(n15936), .B2(n12254), .A(n12097), .ZN(n12098) );
  OAI21_X1 U11444 ( .B1(n14033), .B2(n14037), .A(n14024), .ZN(n14036) );
  OR2_X1 U11445 ( .A1(n14129), .A2(n12622), .ZN(n14044) );
  NAND2_X1 U11446 ( .A1(n10797), .A2(n10796), .ZN(n14033) );
  INV_X1 U11447 ( .A(n11990), .ZN(n9878) );
  NAND2_X1 U11448 ( .A1(n10088), .A2(n10797), .ZN(n10160) );
  NAND2_X1 U11449 ( .A1(n15971), .A2(n20935), .ZN(n14129) );
  NAND2_X1 U11450 ( .A1(n14316), .A2(n13976), .ZN(n19532) );
  NAND2_X1 U11451 ( .A1(n11082), .A2(n11081), .ZN(n16224) );
  AOI21_X2 U11452 ( .B1(n11208), .B2(n11207), .A(n17696), .ZN(n11523) );
  NAND2_X2 U11453 ( .A1(n12621), .A2(n12620), .ZN(n15971) );
  INV_X2 U11454 ( .A(n18916), .ZN(n18923) );
  NAND2_X1 U11455 ( .A1(n19223), .A2(n13381), .ZN(n13383) );
  NAND2_X2 U11456 ( .A1(n17517), .A2(n17516), .ZN(n20748) );
  OR2_X1 U11457 ( .A1(n10477), .A2(n10475), .ZN(n10474) );
  AND2_X1 U11458 ( .A1(n10611), .A2(n10610), .ZN(n10779) );
  AND2_X1 U11459 ( .A1(n11966), .A2(n11967), .ZN(n11988) );
  OAI21_X1 U11460 ( .B1(n10013), .B2(n10489), .A(n13309), .ZN(n10256) );
  XNOR2_X1 U11461 ( .A(n10782), .B(n10090), .ZN(n10794) );
  OR3_X2 U11462 ( .A1(n14576), .A2(n14575), .A3(n14574), .ZN(n15132) );
  XNOR2_X1 U11463 ( .A(n10777), .B(n11392), .ZN(n10778) );
  NAND2_X1 U11464 ( .A1(n11904), .A2(n11903), .ZN(n11961) );
  AND2_X1 U11465 ( .A1(n9980), .A2(n12617), .ZN(n9979) );
  NAND2_X1 U11466 ( .A1(n10521), .A2(n10520), .ZN(n14576) );
  AND3_X1 U11467 ( .A1(n10523), .A2(n14416), .A3(n12648), .ZN(n10520) );
  NAND2_X1 U11468 ( .A1(n17498), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10064) );
  CLKBUF_X1 U11469 ( .A(n11888), .Z(n12623) );
  AOI21_X1 U11470 ( .B1(n10315), .B2(n10314), .A(n9891), .ZN(n10313) );
  INV_X2 U11471 ( .A(n12843), .ZN(n12833) );
  AND3_X1 U11472 ( .A1(n10581), .A2(n11032), .A3(n11037), .ZN(n11028) );
  AND3_X1 U11473 ( .A1(n11902), .A2(n11907), .A3(n13441), .ZN(n11882) );
  OAI21_X1 U11474 ( .B1(n12725), .B2(P1_EBX_REG_1__SCAN_IN), .A(n12642), .ZN(
        n12643) );
  NAND2_X1 U11475 ( .A1(n11015), .A2(n11014), .ZN(n11032) );
  AND3_X1 U11476 ( .A1(n13147), .A2(n11877), .A3(n10358), .ZN(n11906) );
  INV_X1 U11477 ( .A(n10773), .ZN(n12843) );
  NAND2_X1 U11478 ( .A1(n10752), .A2(n10751), .ZN(n9942) );
  NAND2_X1 U11479 ( .A1(n9990), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12614) );
  NAND2_X1 U11480 ( .A1(n10583), .A2(n10582), .ZN(n11037) );
  INV_X2 U11481 ( .A(n11536), .ZN(n18518) );
  AND2_X2 U11482 ( .A1(n10758), .A2(n12848), .ZN(n10773) );
  AND2_X1 U11483 ( .A1(n11868), .A2(n13448), .ZN(n11902) );
  OAI21_X1 U11484 ( .B1(n11261), .B2(n20829), .A(n11226), .ZN(n11233) );
  OAI21_X1 U11485 ( .B1(n10726), .B2(n20183), .A(n10764), .ZN(n9891) );
  NAND4_X1 U11486 ( .A1(n9814), .A2(n9953), .A3(n10345), .A4(n9861), .ZN(
        n10726) );
  INV_X1 U11487 ( .A(n12649), .ZN(n14100) );
  NAND2_X1 U11488 ( .A1(n13290), .A2(n13366), .ZN(n13300) );
  AND2_X1 U11489 ( .A1(n10718), .A2(n10723), .ZN(n12783) );
  CLKBUF_X1 U11490 ( .A(n11187), .Z(n17668) );
  AND2_X1 U11491 ( .A1(n19571), .A2(n17706), .ZN(n13966) );
  AND2_X1 U11492 ( .A1(n19583), .A2(n11677), .ZN(n14310) );
  AND2_X1 U11493 ( .A1(n13439), .A2(n11866), .ZN(n11868) );
  INV_X1 U11494 ( .A(n13296), .ZN(n14235) );
  INV_X1 U11495 ( .A(n20150), .ZN(n19568) );
  CLKBUF_X1 U11496 ( .A(n12086), .Z(n13435) );
  INV_X1 U11497 ( .A(n12638), .ZN(n12649) );
  OAI22_X1 U11498 ( .A1(n10428), .A2(n10740), .B1(n11227), .B2(n10741), .ZN(
        n10069) );
  INV_X1 U11499 ( .A(n10740), .ZN(n9861) );
  INV_X1 U11500 ( .A(n17706), .ZN(n19580) );
  AND2_X1 U11501 ( .A1(n10345), .A2(n10721), .ZN(n10727) );
  INV_X1 U11502 ( .A(n11861), .ZN(n10321) );
  CLKBUF_X3 U11503 ( .A(n12968), .Z(n13010) );
  NAND2_X1 U11504 ( .A1(n10717), .A2(n10809), .ZN(n11472) );
  OR2_X1 U11505 ( .A1(n11614), .A2(n11613), .ZN(n17706) );
  AND2_X1 U11506 ( .A1(n10734), .A2(n17575), .ZN(n10429) );
  OR2_X1 U11507 ( .A1(n13211), .A2(n13210), .ZN(n13366) );
  NAND2_X1 U11508 ( .A1(n14045), .A2(n11872), .ZN(n11890) );
  OR2_X1 U11509 ( .A1(n11670), .A2(n11669), .ZN(n13963) );
  NAND2_X1 U11510 ( .A1(n11170), .A2(n20750), .ZN(n12775) );
  NAND2_X2 U11511 ( .A1(n11769), .A2(n11768), .ZN(n11874) );
  NAND2_X2 U11512 ( .A1(n11844), .A2(n11843), .ZN(n11873) );
  OR2_X1 U11513 ( .A1(n10854), .A2(n10853), .ZN(n11500) );
  OR2_X1 U11514 ( .A1(n10840), .A2(n10839), .ZN(n11499) );
  NAND2_X1 U11515 ( .A1(n10243), .A2(n10242), .ZN(n14161) );
  NAND2_X2 U11516 ( .A1(n9772), .A2(n9722), .ZN(n11872) );
  INV_X1 U11517 ( .A(n11011), .ZN(n12968) );
  INV_X1 U11518 ( .A(n10731), .ZN(n10741) );
  OR2_X1 U11520 ( .A1(n11566), .A2(n11565), .ZN(n11712) );
  AND4_X1 U11521 ( .A1(n11836), .A2(n11835), .A3(n11834), .A4(n11833), .ZN(
        n11844) );
  INV_X1 U11522 ( .A(n14390), .ZN(n14045) );
  NAND4_X2 U11523 ( .A1(n11806), .A2(n11805), .A3(n11804), .A4(n11803), .ZN(
        n11869) );
  AND4_X1 U11524 ( .A1(n11848), .A2(n11847), .A3(n11846), .A4(n11845), .ZN(
        n9772) );
  NOR2_X1 U11525 ( .A1(n13284), .A2(n10244), .ZN(n10243) );
  AND4_X1 U11526 ( .A1(n11763), .A2(n11762), .A3(n11761), .A4(n11760), .ZN(
        n11769) );
  AND4_X2 U11527 ( .A1(n11832), .A2(n11831), .A3(n11830), .A4(n11829), .ZN(
        n14390) );
  AND4_X1 U11528 ( .A1(n11787), .A2(n11786), .A3(n11785), .A4(n11784), .ZN(
        n11806) );
  NAND2_X1 U11529 ( .A1(n10351), .A2(n10350), .ZN(n10074) );
  NAND2_X1 U11530 ( .A1(n10353), .A2(n10352), .ZN(n10075) );
  AND3_X1 U11531 ( .A1(n10650), .A2(n17650), .A3(n10652), .ZN(n10352) );
  AND3_X1 U11532 ( .A1(n10648), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n10649), .ZN(n10350) );
  AND4_X1 U11533 ( .A1(n11767), .A2(n11766), .A3(n11765), .A4(n11764), .ZN(
        n11768) );
  NAND2_X2 U11534 ( .A1(n20144), .A2(n20072), .ZN(n20117) );
  AND4_X1 U11535 ( .A1(n11747), .A2(n11746), .A3(n11745), .A4(n11744), .ZN(
        n11748) );
  AND4_X1 U11536 ( .A1(n11828), .A2(n11827), .A3(n11826), .A4(n11825), .ZN(
        n11829) );
  AND4_X1 U11537 ( .A1(n11822), .A2(n11821), .A3(n11820), .A4(n11819), .ZN(
        n11830) );
  AND4_X1 U11538 ( .A1(n11816), .A2(n11815), .A3(n11814), .A4(n11813), .ZN(
        n11831) );
  AND4_X1 U11539 ( .A1(n11810), .A2(n11809), .A3(n11808), .A4(n11807), .ZN(
        n11832) );
  AND4_X1 U11540 ( .A1(n11802), .A2(n11801), .A3(n11800), .A4(n11799), .ZN(
        n11803) );
  AND4_X1 U11541 ( .A1(n11796), .A2(n11795), .A3(n11794), .A4(n11793), .ZN(
        n11804) );
  AND4_X1 U11542 ( .A1(n11791), .A2(n11790), .A3(n11789), .A4(n11788), .ZN(
        n11805) );
  AND4_X1 U11543 ( .A1(n11842), .A2(n11841), .A3(n11840), .A4(n11839), .ZN(
        n11843) );
  INV_X2 U11544 ( .A(n19442), .ZN(n19494) );
  BUF_X2 U11545 ( .A(n11838), .Z(n12373) );
  INV_X2 U11546 ( .A(n13229), .ZN(n13795) );
  OR2_X1 U11547 ( .A1(n11928), .A2(n11817), .ZN(n11822) );
  BUF_X2 U11548 ( .A(n11928), .Z(n9701) );
  AND2_X1 U11549 ( .A1(n10646), .A2(n10647), .ZN(n10351) );
  AND2_X2 U11550 ( .A1(n16445), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10842) );
  NAND2_X2 U11551 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n20930), .ZN(n20873) );
  NAND2_X2 U11552 ( .A1(n20930), .A2(n20827), .ZN(n20876) );
  AND2_X1 U11553 ( .A1(n10651), .A2(n10653), .ZN(n10353) );
  INV_X2 U11554 ( .A(n11594), .ZN(n9703) );
  NOR2_X1 U11555 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n18541), .ZN(n18513) );
  INV_X2 U11556 ( .A(n18181), .ZN(n18183) );
  CLKBUF_X1 U11557 ( .A(n11798), .Z(n12545) );
  AND2_X2 U11558 ( .A1(n10320), .A2(n13949), .ZN(n11837) );
  OR2_X1 U11559 ( .A1(n12502), .A2(n11812), .ZN(n11813) );
  AND2_X2 U11560 ( .A1(n11743), .A2(n14443), .ZN(n12131) );
  INV_X2 U11561 ( .A(n12631), .ZN(n12058) );
  NOR2_X1 U11562 ( .A1(n17497), .A2(n17650), .ZN(n11191) );
  AND2_X2 U11563 ( .A1(n17468), .A2(n16448), .ZN(n10847) );
  AND2_X2 U11564 ( .A1(n17500), .A2(n17650), .ZN(n17505) );
  AND2_X2 U11565 ( .A1(n9698), .A2(n17650), .ZN(n16473) );
  NAND2_X1 U11566 ( .A1(n11554), .A2(n14720), .ZN(n14594) );
  AND2_X2 U11567 ( .A1(n10833), .A2(n17650), .ZN(n16472) );
  AND2_X2 U11568 ( .A1(n10833), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n16471) );
  AND2_X2 U11569 ( .A1(n17469), .A2(n16448), .ZN(n10848) );
  AND2_X2 U11570 ( .A1(n17482), .A2(n14023), .ZN(n16614) );
  NOR2_X2 U11571 ( .A1(n20062), .A2(P3_STATE_REG_0__SCAN_IN), .ZN(n20121) );
  AND2_X2 U11572 ( .A1(n17482), .A2(n14023), .ZN(n9699) );
  NAND2_X1 U11573 ( .A1(n11559), .A2(n14720), .ZN(n14591) );
  AND2_X1 U11574 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10473) );
  NOR3_X2 U11575 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n16484) );
  NOR2_X2 U11576 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n17481) );
  AND2_X1 U11577 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11555) );
  NOR2_X1 U11578 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n16448) );
  NOR3_X2 U11579 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n18545) );
  CLKBUF_X1 U11580 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n15783) );
  NOR2_X1 U11581 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20888) );
  NAND2_X1 U11582 ( .A1(n9994), .A2(n17140), .ZN(n18085) );
  CLKBUF_X1 U11583 ( .A(n9884), .Z(n9692) );
  NAND2_X1 U11584 ( .A1(n10112), .A2(n10111), .ZN(n9693) );
  INV_X1 U11585 ( .A(n9884), .ZN(n9694) );
  NAND2_X1 U11586 ( .A1(n10112), .A2(n10111), .ZN(n15346) );
  OAI21_X1 U11587 ( .B1(n14524), .B2(n13092), .A(n10044), .ZN(n15501) );
  INV_X2 U11588 ( .A(n14570), .ZN(n12125) );
  NAND2_X1 U11589 ( .A1(n10183), .A2(n10182), .ZN(n11517) );
  XNOR2_X1 U11590 ( .A(n11911), .B(n11914), .ZN(n11944) );
  NOR2_X2 U11591 ( .A1(n14435), .A2(n14403), .ZN(n13945) );
  INV_X4 U11592 ( .A(n11869), .ZN(n13146) );
  NOR2_X2 U11593 ( .A1(n14290), .A2(n14289), .ZN(n14288) );
  AND3_X1 U11594 ( .A1(n11058), .A2(n11251), .A3(n10236), .ZN(n10182) );
  NOR2_X2 U11595 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n18409), .ZN(n18389) );
  AOI21_X1 U11596 ( .B1(n10771), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n10776), .ZN(n11392) );
  NAND2_X1 U11598 ( .A1(n11209), .A2(n10723), .ZN(n11465) );
  NAND2_X4 U11599 ( .A1(n11749), .A2(n11748), .ZN(n11861) );
  AND2_X1 U11600 ( .A1(n13031), .A2(n10174), .ZN(n16886) );
  AND2_X1 U11601 ( .A1(n10765), .A2(n10767), .ZN(n10312) );
  INV_X1 U11602 ( .A(n9971), .ZN(n10728) );
  NAND2_X1 U11603 ( .A1(n10064), .A2(n9826), .ZN(n10754) );
  NAND2_X1 U11604 ( .A1(n15385), .A2(n15384), .ZN(n15360) );
  NOR2_X2 U11605 ( .A1(n14749), .A2(n14760), .ZN(n14759) );
  AND2_X2 U11606 ( .A1(n10720), .A2(n10741), .ZN(n10723) );
  AND2_X1 U11607 ( .A1(n14442), .A2(n13950), .ZN(n9695) );
  AND2_X1 U11608 ( .A1(n14442), .A2(n13950), .ZN(n11798) );
  NOR3_X4 U11609 ( .A1(n16102), .A2(n10484), .A3(n10485), .ZN(n16062) );
  OAI21_X2 U11610 ( .B1(n11919), .B2(n13958), .A(n11905), .ZN(n11911) );
  NAND2_X1 U11611 ( .A1(n10086), .A2(n10084), .ZN(n9696) );
  INV_X2 U11612 ( .A(n11009), .ZN(n9953) );
  NOR2_X2 U11613 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n18293), .ZN(n18275) );
  NOR2_X2 U11614 ( .A1(n10805), .A2(n10808), .ZN(n9911) );
  NAND2_X2 U11615 ( .A1(n10805), .A2(n9903), .ZN(n10926) );
  AND2_X1 U11616 ( .A1(n11741), .A2(n14442), .ZN(n9697) );
  NAND2_X1 U11617 ( .A1(n9926), .A2(n10410), .ZN(n10409) );
  OAI22_X2 U11618 ( .A1(n16860), .A2(n16298), .B1(n11260), .B2(n9702), .ZN(
        n14048) );
  NAND3_X2 U11619 ( .A1(n9731), .A2(n14352), .A3(n11255), .ZN(n16860) );
  AND2_X1 U11620 ( .A1(n17482), .A2(n14023), .ZN(n9698) );
  NAND2_X1 U11622 ( .A1(n14719), .A2(n11555), .ZN(n11594) );
  NAND2_X2 U11623 ( .A1(n11913), .A2(n11912), .ZN(n11945) );
  NOR2_X2 U11624 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n18270), .ZN(n18253) );
  AOI211_X2 U11625 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n18260), .A(n18235), 
        .B(n18234), .ZN(n18238) );
  INV_X2 U11626 ( .A(n19067), .ZN(n19159) );
  NOR2_X2 U11627 ( .A1(n19067), .A2(n19082), .ZN(n19281) );
  NOR2_X2 U11628 ( .A1(n19278), .A2(n20049), .ZN(n19067) );
  AOI21_X1 U11629 ( .B1(n11921), .B2(n15783), .A(n11920), .ZN(n11966) );
  XNOR2_X1 U11630 ( .A(n12565), .B(n12564), .ZN(n14818) );
  OR2_X1 U11631 ( .A1(n10370), .A2(n9738), .ZN(n10119) );
  OAI21_X1 U11632 ( .B1(n13415), .B2(n14808), .A(n13416), .ZN(n14793) );
  NOR2_X2 U11633 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n18247), .ZN(n18230) );
  NAND2_X2 U11634 ( .A1(n13062), .A2(n15988), .ZN(n15987) );
  NOR2_X4 U11635 ( .A1(n13061), .A2(n13063), .ZN(n13062) );
  NAND2_X2 U11636 ( .A1(n12281), .A2(n12280), .ZN(n14992) );
  AOI21_X2 U11637 ( .B1(n10771), .B2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n10756), .ZN(n10783) );
  XNOR2_X1 U11638 ( .A(n9877), .B(n10365), .ZN(n13097) );
  AND2_X2 U11639 ( .A1(n12763), .A2(n9834), .ZN(n16048) );
  NOR2_X2 U11640 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n18485), .ZN(n18464) );
  NAND2_X2 U11641 ( .A1(n14367), .A2(n14366), .ZN(n14365) );
  NOR2_X2 U11642 ( .A1(n16181), .A2(n10479), .ZN(n16134) );
  AND2_X1 U11643 ( .A1(n11741), .A2(n14442), .ZN(n11936) );
  AND2_X1 U11644 ( .A1(n11741), .A2(n10320), .ZN(n9712) );
  INV_X1 U11645 ( .A(n9713), .ZN(n9714) );
  AND2_X2 U11646 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n17482) );
  AND2_X1 U11647 ( .A1(n10320), .A2(n11743), .ZN(n9715) );
  AND2_X1 U11648 ( .A1(n10320), .A2(n11743), .ZN(n11849) );
  OR2_X1 U11649 ( .A1(n13160), .A2(n20196), .ZN(n10487) );
  NAND2_X1 U11650 ( .A1(n13069), .A2(n13071), .ZN(n13139) );
  XNOR2_X2 U11651 ( .A(n14826), .B(n12852), .ZN(n14806) );
  NAND2_X2 U11652 ( .A1(n13150), .A2(n10558), .ZN(n14826) );
  AND2_X1 U11653 ( .A1(n11742), .A2(n13950), .ZN(n9716) );
  AND2_X1 U11654 ( .A1(n11742), .A2(n13950), .ZN(n9717) );
  AND2_X1 U11655 ( .A1(n11742), .A2(n13950), .ZN(n11818) );
  NOR2_X1 U11656 ( .A1(n14524), .A2(n9709), .ZN(n15848) );
  AND3_X1 U11657 ( .A1(n21181), .A2(n9709), .A3(n14362), .ZN(n21419) );
  XNOR2_X2 U11658 ( .A(n14365), .B(n14457), .ZN(n14439) );
  NAND2_X1 U11659 ( .A1(n10029), .A2(n10326), .ZN(n9950) );
  NAND2_X1 U11660 ( .A1(n10328), .A2(n9827), .ZN(n10326) );
  AND2_X1 U11661 ( .A1(n10381), .A2(n10228), .ZN(n10227) );
  INV_X1 U11662 ( .A(n16990), .ZN(n10228) );
  NAND2_X1 U11663 ( .A1(n9931), .A2(n10742), .ZN(n10763) );
  NAND2_X1 U11664 ( .A1(n9875), .A2(n9784), .ZN(n9874) );
  NAND2_X1 U11665 ( .A1(n15475), .A2(n10541), .ZN(n9875) );
  NAND2_X1 U11666 ( .A1(n9873), .A2(n9781), .ZN(n9872) );
  NAND2_X1 U11667 ( .A1(n10361), .A2(n10635), .ZN(n9873) );
  AND2_X1 U11668 ( .A1(n10358), .A2(n11874), .ZN(n11927) );
  NAND2_X1 U11669 ( .A1(n13411), .A2(n10152), .ZN(n10535) );
  AND2_X1 U11670 ( .A1(n15394), .A2(n15531), .ZN(n10152) );
  NAND2_X1 U11671 ( .A1(n9879), .A2(n9878), .ZN(n9876) );
  NAND2_X1 U11672 ( .A1(n10202), .A2(n17650), .ZN(n10082) );
  NAND2_X1 U11673 ( .A1(n10201), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10083) );
  OR2_X1 U11674 ( .A1(n16171), .A2(n11108), .ZN(n12989) );
  NAND2_X1 U11675 ( .A1(n11518), .A2(n9946), .ZN(n9945) );
  NOR2_X1 U11676 ( .A1(n11073), .A2(n9966), .ZN(n9946) );
  NOR2_X1 U11677 ( .A1(n10606), .A2(n10914), .ZN(n10604) );
  AND2_X1 U11678 ( .A1(n11709), .A2(n11711), .ZN(n13350) );
  OR2_X1 U11679 ( .A1(n13348), .A2(n11705), .ZN(n11709) );
  INV_X1 U11680 ( .A(n10219), .ZN(n10218) );
  NAND2_X1 U11681 ( .A1(n10609), .A2(n9777), .ZN(n10222) );
  OAI21_X1 U11682 ( .B1(n10221), .B2(n10220), .A(n12982), .ZN(n10219) );
  NAND2_X2 U11683 ( .A1(n9997), .A2(n9995), .ZN(n9926) );
  NAND2_X1 U11684 ( .A1(n9996), .A2(n10269), .ZN(n9995) );
  NAND2_X1 U11685 ( .A1(n17096), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n9997) );
  NAND2_X1 U11686 ( .A1(n10617), .A2(n17109), .ZN(n9996) );
  NAND2_X1 U11687 ( .A1(n9953), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10743) );
  NOR2_X1 U11688 ( .A1(n10793), .A2(n10789), .ZN(n10159) );
  NAND2_X1 U11689 ( .A1(n9825), .A2(n15959), .ZN(n10044) );
  INV_X1 U11690 ( .A(n9983), .ZN(n9982) );
  OAI21_X1 U11691 ( .B1(n12591), .B2(n9758), .A(n12607), .ZN(n9983) );
  NAND2_X1 U11692 ( .A1(n12568), .A2(n13127), .ZN(n12608) );
  NAND2_X1 U11693 ( .A1(n9999), .A2(n9998), .ZN(n10749) );
  NAND2_X1 U11694 ( .A1(n10002), .A2(n11000), .ZN(n9998) );
  NOR2_X1 U11695 ( .A1(n10640), .A2(n10608), .ZN(n10422) );
  NAND2_X1 U11696 ( .A1(n9792), .A2(n10645), .ZN(n10423) );
  AND2_X1 U11697 ( .A1(n10550), .A2(n10549), .ZN(n10548) );
  INV_X1 U11698 ( .A(n14876), .ZN(n10549) );
  AND2_X1 U11699 ( .A1(n10555), .A2(n9824), .ZN(n10280) );
  AND2_X1 U11700 ( .A1(n9831), .A2(n15100), .ZN(n10555) );
  INV_X1 U11701 ( .A(n12048), .ZN(n10140) );
  NAND2_X1 U11702 ( .A1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n12048) );
  NOR2_X1 U11703 ( .A1(n10368), .A2(n10114), .ZN(n10543) );
  NOR2_X1 U11704 ( .A1(n10533), .A2(n14932), .ZN(n10532) );
  INV_X1 U11705 ( .A(n14923), .ZN(n10533) );
  INV_X1 U11706 ( .A(n14271), .ZN(n10523) );
  NAND2_X1 U11707 ( .A1(n10322), .A2(n10514), .ZN(n13088) );
  NAND2_X1 U11708 ( .A1(n15165), .A2(n9937), .ZN(n9936) );
  NAND2_X1 U11709 ( .A1(n11874), .A2(n14385), .ZN(n11855) );
  AND2_X2 U11710 ( .A1(n12086), .A2(n11873), .ZN(n13440) );
  NAND2_X1 U11711 ( .A1(n11962), .A2(n11961), .ZN(n10539) );
  OR2_X1 U11712 ( .A1(n12610), .A2(n12609), .ZN(n12612) );
  MUX2_X1 U11713 ( .A(n11246), .B(n11197), .S(n12958), .Z(n11148) );
  AOI21_X1 U11714 ( .B1(n16065), .B2(n13001), .A(n10589), .ZN(n10588) );
  OAI21_X1 U11715 ( .B1(n10592), .B2(n10590), .A(n13006), .ZN(n10589) );
  INV_X1 U11716 ( .A(n10593), .ZN(n10590) );
  OAI21_X1 U11717 ( .B1(n11148), .B2(n13010), .A(n11005), .ZN(n11030) );
  OR2_X1 U11718 ( .A1(n11012), .A2(n11004), .ZN(n11005) );
  INV_X1 U11719 ( .A(n9978), .ZN(n9973) );
  NAND2_X1 U11720 ( .A1(n12916), .A2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12920) );
  NAND2_X1 U11721 ( .A1(n10780), .A2(n10779), .ZN(n10401) );
  NAND2_X1 U11722 ( .A1(n9929), .A2(n10606), .ZN(n10603) );
  NAND2_X2 U11723 ( .A1(n10086), .A2(n10084), .ZN(n11212) );
  NAND2_X1 U11724 ( .A1(n10087), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10086) );
  INV_X1 U11725 ( .A(n10262), .ZN(n10261) );
  NAND2_X1 U11726 ( .A1(n21349), .A2(n21468), .ZN(n12631) );
  INV_X1 U11727 ( .A(n12739), .ZN(n10519) );
  INV_X1 U11728 ( .A(n12157), .ZN(n12158) );
  NAND2_X1 U11729 ( .A1(n10123), .A2(n15394), .ZN(n10122) );
  INV_X1 U11730 ( .A(n13411), .ZN(n10123) );
  NAND2_X1 U11731 ( .A1(n14439), .A2(n20939), .ZN(n10538) );
  INV_X1 U11732 ( .A(n12061), .ZN(n9877) );
  XNOR2_X1 U11733 ( .A(n12970), .B(n12969), .ZN(n13020) );
  NAND2_X1 U11734 ( .A1(n11089), .A2(n9787), .ZN(n11110) );
  NAND2_X1 U11735 ( .A1(n13031), .A2(n10271), .ZN(n9934) );
  NOR2_X1 U11736 ( .A1(n9852), .A2(n10272), .ZN(n10271) );
  INV_X1 U11737 ( .A(n13030), .ZN(n10272) );
  NAND2_X1 U11738 ( .A1(n11072), .A2(n11012), .ZN(n13022) );
  AND2_X1 U11739 ( .A1(n13479), .A2(n16884), .ZN(n10644) );
  AND2_X1 U11740 ( .A1(n13013), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n16916) );
  INV_X1 U11741 ( .A(n10329), .ZN(n13002) );
  AND2_X1 U11742 ( .A1(n16974), .A2(n13497), .ZN(n16960) );
  NOR2_X1 U11743 ( .A1(n11123), .A2(n10393), .ZN(n10392) );
  INV_X1 U11744 ( .A(n16973), .ZN(n10393) );
  INV_X1 U11745 ( .A(n12989), .ZN(n10225) );
  INV_X1 U11746 ( .A(n10227), .ZN(n10226) );
  NAND2_X1 U11747 ( .A1(n10293), .A2(n10403), .ZN(n10292) );
  NOR2_X1 U11748 ( .A1(n10411), .A2(n10296), .ZN(n10295) );
  NAND2_X1 U11749 ( .A1(n17021), .A2(n11521), .ZN(n17022) );
  OAI211_X1 U11750 ( .C1(n10237), .C2(n10618), .A(n10269), .B(n17109), .ZN(
        n10268) );
  AND4_X1 U11751 ( .A1(n17458), .A2(n13059), .A3(n11206), .A4(n11205), .ZN(
        n11207) );
  NAND2_X1 U11752 ( .A1(n12871), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12872) );
  OR3_X1 U11753 ( .A1(n13348), .A2(n13347), .A3(n13346), .ZN(n13349) );
  AND2_X1 U11754 ( .A1(n9736), .A2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n10495) );
  INV_X1 U11755 ( .A(n18887), .ZN(n17908) );
  INV_X1 U11756 ( .A(n13295), .ZN(n10015) );
  NAND2_X1 U11757 ( .A1(n13295), .A2(n21791), .ZN(n10014) );
  AND2_X1 U11758 ( .A1(n12750), .A2(n12740), .ZN(n20992) );
  AOI21_X1 U11759 ( .B1(n13063), .B2(n16022), .A(n13062), .ZN(n16633) );
  NAND2_X1 U11760 ( .A1(n18060), .A2(n20246), .ZN(n17146) );
  NAND2_X1 U11761 ( .A1(n10288), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n10285) );
  INV_X1 U11762 ( .A(n20436), .ZN(n10288) );
  NOR2_X1 U11763 ( .A1(n14079), .A2(n10791), .ZN(n9902) );
  AND2_X1 U11764 ( .A1(n10820), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n10283) );
  NAND2_X1 U11765 ( .A1(n9911), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n9914) );
  NAND2_X1 U11766 ( .A1(n20900), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11002) );
  INV_X1 U11767 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n10545) );
  AND2_X1 U11768 ( .A1(n12054), .A2(n12112), .ZN(n10547) );
  INV_X1 U11769 ( .A(n11872), .ZN(n11870) );
  AND2_X1 U11770 ( .A1(n13147), .A2(n13149), .ZN(n13454) );
  INV_X1 U11771 ( .A(n11927), .ZN(n9990) );
  NAND2_X1 U11772 ( .A1(n10763), .A2(n10744), .ZN(n10745) );
  NOR2_X1 U11773 ( .A1(n14053), .A2(n17703), .ZN(n10314) );
  NAND2_X1 U11774 ( .A1(n10739), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10767) );
  NAND2_X1 U11775 ( .A1(n10762), .A2(n17667), .ZN(n10180) );
  OAI22_X1 U11776 ( .A1(n10881), .A2(n20606), .B1(n20740), .B2(n10880), .ZN(
        n10885) );
  NAND2_X1 U11777 ( .A1(n16097), .A2(n13049), .ZN(n11134) );
  AND2_X1 U11778 ( .A1(n10414), .A2(n11073), .ZN(n10203) );
  AND3_X1 U11779 ( .A1(n9733), .A2(n10948), .A3(n9799), .ZN(n11022) );
  INV_X1 U11780 ( .A(n19210), .ZN(n10489) );
  NOR2_X1 U11781 ( .A1(n10489), .A2(n10259), .ZN(n10258) );
  NAND2_X1 U11782 ( .A1(n13241), .A2(n13240), .ZN(n13306) );
  NAND2_X1 U11783 ( .A1(n14161), .A2(n14167), .ZN(n13369) );
  NOR2_X1 U11784 ( .A1(n11874), .A2(n11873), .ZN(n14097) );
  NAND2_X1 U11785 ( .A1(n15934), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12537) );
  INV_X1 U11786 ( .A(n15130), .ZN(n10281) );
  NOR2_X2 U11787 ( .A1(n11861), .A2(n21349), .ZN(n12254) );
  AND2_X1 U11788 ( .A1(n15404), .A2(n9854), .ZN(n10057) );
  OR2_X1 U11789 ( .A1(n9688), .A2(n13140), .ZN(n15436) );
  NOR2_X1 U11790 ( .A1(n18018), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10047) );
  INV_X1 U11791 ( .A(n12725), .ZN(n12727) );
  NAND2_X1 U11792 ( .A1(n10041), .A2(n10040), .ZN(n10043) );
  AOI21_X1 U11793 ( .B1(n10044), .B2(n13092), .A(n21114), .ZN(n10040) );
  NAND2_X1 U11794 ( .A1(n14524), .A2(n10044), .ZN(n10041) );
  NAND2_X1 U11795 ( .A1(n13080), .A2(n13127), .ZN(n10110) );
  NOR2_X1 U11796 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n21144), .ZN(
        n10100) );
  INV_X1 U11797 ( .A(n14304), .ZN(n10098) );
  AND2_X1 U11798 ( .A1(n13096), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10097) );
  OR2_X1 U11799 ( .A1(n11959), .A2(n11958), .ZN(n13084) );
  AND2_X1 U11800 ( .A1(n11924), .A2(n14404), .ZN(n15852) );
  AOI21_X1 U11801 ( .B1(n16336), .B2(n10190), .A(n10189), .ZN(n10188) );
  INV_X1 U11802 ( .A(n16925), .ZN(n10189) );
  NOR2_X1 U11803 ( .A1(n12915), .A2(n12919), .ZN(n10200) );
  NOR2_X1 U11804 ( .A1(n9735), .A2(n10309), .ZN(n10308) );
  INV_X1 U11805 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n10584) );
  INV_X1 U11806 ( .A(n11120), .ZN(n10585) );
  NAND2_X1 U11807 ( .A1(n11023), .A2(n11061), .ZN(n10596) );
  CLKBUF_X1 U11808 ( .A(n10696), .Z(n16612) );
  NAND2_X1 U11809 ( .A1(n16422), .A2(n10452), .ZN(n10451) );
  INV_X1 U11810 ( .A(n16673), .ZN(n10452) );
  INV_X1 U11811 ( .A(n16691), .ZN(n10449) );
  AND2_X1 U11812 ( .A1(n14284), .A2(n14283), .ZN(n9978) );
  NAND2_X1 U11813 ( .A1(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n10439) );
  NOR2_X1 U11814 ( .A1(n21656), .A2(n10448), .ZN(n10447) );
  NOR2_X1 U11815 ( .A1(n12899), .A2(n12903), .ZN(n12902) );
  NAND2_X1 U11816 ( .A1(n11411), .A2(n10478), .ZN(n10477) );
  INV_X1 U11817 ( .A(n16267), .ZN(n10478) );
  NAND2_X1 U11818 ( .A1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10444) );
  NAND2_X1 U11819 ( .A1(n10748), .A2(n10749), .ZN(n10610) );
  NAND2_X1 U11820 ( .A1(n10613), .A2(n10612), .ZN(n10780) );
  NAND2_X1 U11821 ( .A1(n10026), .A2(n10599), .ZN(n13003) );
  AOI21_X1 U11822 ( .B1(n16936), .B2(n9751), .A(n10600), .ZN(n10599) );
  NAND2_X1 U11823 ( .A1(n16931), .A2(n10598), .ZN(n10026) );
  NAND2_X1 U11824 ( .A1(n10601), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n10600) );
  NAND2_X1 U11825 ( .A1(n10576), .A2(n10575), .ZN(n10574) );
  INV_X1 U11826 ( .A(n16001), .ZN(n10576) );
  INV_X1 U11827 ( .A(n16005), .ZN(n10575) );
  NAND2_X1 U11828 ( .A1(n13049), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10303) );
  INV_X1 U11829 ( .A(n16075), .ZN(n10561) );
  AND2_X1 U11830 ( .A1(n10571), .A2(n10570), .ZN(n10569) );
  INV_X1 U11831 ( .A(n14782), .ZN(n10570) );
  NOR2_X1 U11832 ( .A1(n10471), .A2(n10470), .ZN(n10469) );
  INV_X1 U11833 ( .A(n16203), .ZN(n10470) );
  NAND2_X1 U11834 ( .A1(n11333), .A2(n10567), .ZN(n10566) );
  INV_X1 U11835 ( .A(n14755), .ZN(n10567) );
  INV_X1 U11836 ( .A(n14515), .ZN(n11333) );
  NAND2_X1 U11837 ( .A1(n10639), .A2(n10578), .ZN(n10577) );
  INV_X1 U11838 ( .A(n14244), .ZN(n10578) );
  NOR2_X1 U11839 ( .A1(n11073), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n9963) );
  NAND3_X1 U11840 ( .A1(n10325), .A2(n10093), .A3(n10603), .ZN(n10092) );
  AND2_X1 U11841 ( .A1(n11073), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10093) );
  NAND2_X1 U11842 ( .A1(n10027), .A2(n10028), .ZN(n10618) );
  NAND2_X1 U11843 ( .A1(n18085), .A2(n9730), .ZN(n10027) );
  INV_X1 U11844 ( .A(n11022), .ZN(n11256) );
  OR2_X1 U11845 ( .A1(n10913), .A2(n10912), .ZN(n11251) );
  AND2_X1 U11846 ( .A1(n11169), .A2(n11476), .ZN(n11470) );
  OAI21_X1 U11847 ( .B1(n10734), .B2(n11215), .A(n20750), .ZN(n11216) );
  INV_X1 U11848 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10404) );
  NAND2_X1 U11849 ( .A1(n14022), .A2(n20750), .ZN(n14221) );
  NAND2_X1 U11850 ( .A1(n14072), .A2(n14071), .ZN(n14214) );
  NOR2_X1 U11851 ( .A1(n14079), .A2(n10089), .ZN(n10810) );
  NOR2_X1 U11852 ( .A1(n10790), .A2(n14079), .ZN(n9901) );
  INV_X1 U11853 ( .A(n10819), .ZN(n10820) );
  AND2_X1 U11854 ( .A1(n9739), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n10505) );
  AND2_X1 U11855 ( .A1(n14728), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11548) );
  AND2_X1 U11856 ( .A1(n14747), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11558) );
  OAI21_X1 U11857 ( .B1(n11691), .B2(n13691), .A(n17978), .ZN(n14153) );
  INV_X1 U11858 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n17834) );
  NOR2_X1 U11859 ( .A1(n19218), .A2(n10512), .ZN(n10511) );
  INV_X1 U11860 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n10512) );
  NOR2_X1 U11861 ( .A1(n13352), .A2(n18185), .ZN(n14321) );
  OAI21_X1 U11862 ( .B1(n11672), .B2(n14310), .A(n11671), .ZN(n11686) );
  INV_X1 U11863 ( .A(n13966), .ZN(n11671) );
  XNOR2_X1 U11864 ( .A(n13300), .B(n14235), .ZN(n13297) );
  NAND2_X1 U11865 ( .A1(n13981), .A2(n14312), .ZN(n14313) );
  OR2_X1 U11866 ( .A1(n11641), .A2(n11640), .ZN(n11687) );
  NOR2_X1 U11867 ( .A1(n12623), .A2(n12624), .ZN(n13866) );
  INV_X1 U11868 ( .A(n14262), .ZN(n12100) );
  NAND2_X1 U11869 ( .A1(n11921), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n9938) );
  NAND2_X1 U11870 ( .A1(n11894), .A2(n11893), .ZN(n11904) );
  NOR2_X1 U11871 ( .A1(n14877), .A2(n14861), .ZN(n10529) );
  INV_X1 U11872 ( .A(n10531), .ZN(n10526) );
  INV_X2 U11873 ( .A(n12649), .ZN(n14098) );
  INV_X1 U11874 ( .A(n15223), .ZN(n14801) );
  INV_X1 U11875 ( .A(n12062), .ZN(n12563) );
  NAND2_X1 U11876 ( .A1(n12540), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12566) );
  AND2_X1 U11877 ( .A1(n10559), .A2(n13152), .ZN(n10558) );
  AND2_X1 U11878 ( .A1(n10560), .A2(n14827), .ZN(n10559) );
  INV_X1 U11879 ( .A(n14838), .ZN(n10560) );
  NAND2_X1 U11880 ( .A1(n12441), .A2(n9749), .ZN(n12481) );
  OR2_X1 U11881 ( .A1(n12300), .A2(n12299), .ZN(n12332) );
  INV_X1 U11882 ( .A(n15009), .ZN(n12280) );
  NOR2_X1 U11883 ( .A1(n15025), .A2(n10150), .ZN(n10149) );
  NOR2_X1 U11884 ( .A1(n12208), .A2(n12207), .ZN(n12244) );
  OR2_X1 U11885 ( .A1(n12225), .A2(n15451), .ZN(n12208) );
  NOR2_X1 U11886 ( .A1(n10156), .A2(n10155), .ZN(n10154) );
  NAND2_X1 U11887 ( .A1(n12158), .A2(n10153), .ZN(n12225) );
  AND2_X1 U11888 ( .A1(n10154), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n10153) );
  NOR2_X1 U11889 ( .A1(n15138), .A2(n10138), .ZN(n10137) );
  INV_X1 U11890 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n15138) );
  NAND2_X1 U11891 ( .A1(n10057), .A2(n10130), .ZN(n15359) );
  NAND2_X1 U11892 ( .A1(n10045), .A2(n18018), .ZN(n13125) );
  NAND2_X1 U11893 ( .A1(n18017), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13124) );
  NAND2_X1 U11894 ( .A1(n10107), .A2(n10310), .ZN(n10045) );
  INV_X1 U11895 ( .A(n14266), .ZN(n10521) );
  NOR2_X1 U11896 ( .A1(n11874), .A2(n20939), .ZN(n12089) );
  AND3_X1 U11897 ( .A1(n14381), .A2(n13146), .A3(n14390), .ZN(n11854) );
  NOR2_X1 U11898 ( .A1(n15796), .A2(n21460), .ZN(n21386) );
  OAI22_X1 U11899 ( .A1(n15763), .A2(n21619), .B1(P1_STATE2_REG_0__SCAN_IN), 
        .B2(n21594), .ZN(n15818) );
  INV_X1 U11900 ( .A(n15818), .ZN(n15796) );
  NAND2_X1 U11901 ( .A1(n12619), .A2(n12618), .ZN(n12620) );
  NAND2_X1 U11902 ( .A1(n9981), .A2(n9979), .ZN(n12621) );
  INV_X1 U11903 ( .A(n15961), .ZN(n15966) );
  OR2_X1 U11904 ( .A1(n13018), .A2(n13017), .ZN(n12970) );
  AND2_X1 U11905 ( .A1(n13009), .A2(n13008), .ZN(n16026) );
  NAND2_X1 U11906 ( .A1(n16039), .A2(n16336), .ZN(n10193) );
  INV_X1 U11907 ( .A(n11083), .ZN(n11082) );
  NAND2_X1 U11908 ( .A1(n11032), .A2(n11037), .ZN(n11029) );
  OR2_X1 U11909 ( .A1(n16637), .A2(n10461), .ZN(n10464) );
  NAND2_X1 U11910 ( .A1(n9820), .A2(n10462), .ZN(n10461) );
  INV_X1 U11911 ( .A(n16636), .ZN(n10462) );
  INV_X1 U11912 ( .A(n16604), .ZN(n10460) );
  NAND2_X1 U11913 ( .A1(n10457), .A2(n10456), .ZN(n10455) );
  NAND2_X1 U11914 ( .A1(n10457), .A2(n10454), .ZN(n10453) );
  INV_X1 U11915 ( .A(n16660), .ZN(n10456) );
  NOR2_X1 U11916 ( .A1(n16669), .A2(n16503), .ZN(n10458) );
  OR2_X1 U11917 ( .A1(n16444), .A2(n16443), .ZN(n16668) );
  AND2_X1 U11918 ( .A1(n12968), .A2(n10734), .ZN(n16743) );
  AND2_X1 U11919 ( .A1(n12917), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12916) );
  INV_X1 U11920 ( .A(n16904), .ZN(n10037) );
  NAND2_X1 U11921 ( .A1(n16892), .A2(n16895), .ZN(n10036) );
  NAND2_X1 U11922 ( .A1(n13031), .A2(n13030), .ZN(n10175) );
  INV_X1 U11923 ( .A(n10598), .ZN(n9869) );
  INV_X1 U11924 ( .A(n10597), .ZN(n9867) );
  OR2_X1 U11925 ( .A1(n10482), .A2(n10480), .ZN(n10479) );
  INV_X1 U11926 ( .A(n16153), .ZN(n10480) );
  AND2_X1 U11927 ( .A1(n10403), .A2(n13507), .ZN(n10402) );
  INV_X1 U11928 ( .A(n16181), .ZN(n10481) );
  INV_X1 U11929 ( .A(n10609), .ZN(n10387) );
  INV_X1 U11930 ( .A(n17011), .ZN(n10389) );
  AOI21_X1 U11931 ( .B1(n10411), .B2(n10619), .A(n10296), .ZN(n10291) );
  NOR2_X1 U11932 ( .A1(n10300), .A2(n10240), .ZN(n10012) );
  AND3_X1 U11933 ( .A1(n11306), .A2(n11305), .A3(n11304), .ZN(n14358) );
  NAND2_X1 U11934 ( .A1(n17021), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n17066) );
  NAND2_X1 U11935 ( .A1(n10325), .A2(n10603), .ZN(n9930) );
  INV_X1 U11936 ( .A(n9942), .ZN(n9944) );
  NAND2_X1 U11937 ( .A1(n10181), .A2(n11202), .ZN(n11210) );
  INV_X1 U11938 ( .A(n14774), .ZN(n17419) );
  OR2_X1 U11939 ( .A1(n20896), .A2(n20903), .ZN(n20666) );
  OR2_X1 U11940 ( .A1(n20896), .A2(n17513), .ZN(n20747) );
  NAND2_X1 U11941 ( .A1(n17685), .A2(n17703), .ZN(n17517) );
  INV_X1 U11942 ( .A(n13965), .ZN(n20018) );
  OAI22_X2 U11943 ( .A1(n13357), .A2(n20016), .B1(n20022), .B2(n19543), .ZN(
        n20024) );
  NAND2_X1 U11944 ( .A1(n10499), .A2(n10498), .ZN(n18286) );
  AND2_X1 U11945 ( .A1(n10501), .A2(n10503), .ZN(n10498) );
  INV_X1 U11946 ( .A(n13279), .ZN(n13761) );
  AND2_X1 U11947 ( .A1(n19002), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17778) );
  INV_X1 U11948 ( .A(n19055), .ZN(n10496) );
  NAND2_X1 U11949 ( .A1(n17819), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n17810) );
  NAND2_X1 U11950 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n19238) );
  NAND2_X1 U11951 ( .A1(n10023), .A2(n9732), .ZN(n10021) );
  NAND2_X1 U11952 ( .A1(n17815), .A2(n10017), .ZN(n17800) );
  INV_X1 U11953 ( .A(n10018), .ZN(n10017) );
  OAI21_X1 U11954 ( .B1(n19325), .B2(n10019), .A(n9785), .ZN(n10018) );
  OR2_X1 U11955 ( .A1(n13310), .A2(n17908), .ZN(n19030) );
  NAND2_X1 U11956 ( .A1(n9846), .A2(n10263), .ZN(n10262) );
  INV_X1 U11957 ( .A(n10493), .ZN(n10492) );
  NAND2_X1 U11958 ( .A1(n19204), .A2(n9780), .ZN(n10253) );
  NAND2_X1 U11959 ( .A1(n13384), .A2(n19215), .ZN(n19201) );
  NAND2_X1 U11960 ( .A1(n19226), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13305) );
  XNOR2_X1 U11961 ( .A(n13297), .B(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n19234) );
  INV_X1 U11962 ( .A(n13293), .ZN(n10016) );
  NOR2_X1 U11963 ( .A1(n13350), .A2(n13335), .ZN(n13965) );
  NOR2_X2 U11964 ( .A1(n20168), .A2(n14320), .ZN(n20023) );
  INV_X1 U11965 ( .A(n20047), .ZN(n18192) );
  INV_X1 U11966 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n20049) );
  NOR2_X1 U11967 ( .A1(n20156), .A2(n20151), .ZN(n20159) );
  INV_X1 U11968 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n21468) );
  NOR2_X1 U11969 ( .A1(n10147), .A2(n10146), .ZN(n10145) );
  AOI21_X1 U11970 ( .B1(n21029), .B2(n14277), .A(n21030), .ZN(n10146) );
  NOR2_X1 U11971 ( .A1(n21026), .A2(n21124), .ZN(n10147) );
  AND2_X1 U11972 ( .A1(n14812), .A2(n12860), .ZN(n21027) );
  NAND2_X1 U11973 ( .A1(n10517), .A2(n12737), .ZN(n15512) );
  NAND2_X1 U11974 ( .A1(n10519), .A2(n10518), .ZN(n10517) );
  INV_X1 U11975 ( .A(n12738), .ZN(n10518) );
  XNOR2_X1 U11976 ( .A(n10157), .B(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14812) );
  NOR2_X1 U11977 ( .A1(n14790), .A2(n12566), .ZN(n10157) );
  NOR2_X1 U11978 ( .A1(n14875), .A2(n14865), .ZN(n10279) );
  INV_X1 U11979 ( .A(n15512), .ZN(n10133) );
  XNOR2_X1 U11980 ( .A(n10134), .B(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n15519) );
  NAND2_X1 U11981 ( .A1(n10369), .A2(n14809), .ZN(n10134) );
  NAND2_X1 U11982 ( .A1(n9986), .A2(n14789), .ZN(n9985) );
  OR2_X1 U11983 ( .A1(n14807), .A2(n21125), .ZN(n9986) );
  OR2_X1 U11984 ( .A1(n10370), .A2(n10056), .ZN(n10115) );
  NAND2_X1 U11985 ( .A1(n10122), .A2(n10124), .ZN(n10121) );
  INV_X1 U11986 ( .A(n15346), .ZN(n15335) );
  NOR2_X2 U11987 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n21376) );
  AND2_X1 U11988 ( .A1(n14471), .A2(n9709), .ZN(n21268) );
  NAND2_X1 U11989 ( .A1(n15990), .A2(n16210), .ZN(n15999) );
  NAND2_X1 U11990 ( .A1(n12943), .A2(n20204), .ZN(n16210) );
  INV_X1 U11991 ( .A(n20192), .ZN(n16348) );
  AND2_X1 U11992 ( .A1(n13686), .A2(n17640), .ZN(n20195) );
  NAND2_X1 U11993 ( .A1(n13623), .A2(n12953), .ZN(n16351) );
  XNOR2_X1 U11994 ( .A(n12845), .B(n12844), .ZN(n13160) );
  NAND2_X1 U11995 ( .A1(n12963), .A2(n10641), .ZN(n16752) );
  NAND2_X1 U11996 ( .A1(n12799), .A2(n12798), .ZN(n16850) );
  NAND2_X2 U11997 ( .A1(n12785), .A2(n20180), .ZN(n16867) );
  INV_X1 U11998 ( .A(n20914), .ZN(n17543) );
  INV_X1 U11999 ( .A(n16872), .ZN(n16852) );
  AND2_X1 U12000 ( .A1(n13603), .A2(n9710), .ZN(n13686) );
  NAND2_X1 U12001 ( .A1(n10338), .A2(n10336), .ZN(n10335) );
  NAND2_X1 U12002 ( .A1(n10337), .A2(n10340), .ZN(n10336) );
  NAND2_X1 U12003 ( .A1(n10339), .A2(n10344), .ZN(n10338) );
  INV_X1 U12004 ( .A(n10344), .ZN(n10337) );
  NAND2_X1 U12005 ( .A1(n9871), .A2(n9789), .ZN(n10333) );
  INV_X1 U12006 ( .A(n10342), .ZN(n10341) );
  NAND2_X1 U12007 ( .A1(n16958), .A2(n20252), .ZN(n9970) );
  INV_X1 U12008 ( .A(n16957), .ZN(n9969) );
  AND2_X1 U12009 ( .A1(n13027), .A2(n10356), .ZN(n10355) );
  NAND2_X1 U12010 ( .A1(n11522), .A2(n10357), .ZN(n10356) );
  AOI21_X1 U12011 ( .B1(n16997), .B2(n10357), .A(n20256), .ZN(n9919) );
  NAND2_X1 U12012 ( .A1(n17295), .A2(n17155), .ZN(n10163) );
  NAND2_X1 U12013 ( .A1(n20182), .A2(n13064), .ZN(n18060) );
  INV_X1 U12014 ( .A(n17146), .ZN(n18063) );
  INV_X1 U12015 ( .A(n18060), .ZN(n20247) );
  NAND2_X1 U12016 ( .A1(n13033), .A2(n20277), .ZN(n9933) );
  OAI21_X1 U12017 ( .B1(n13478), .B2(n13481), .A(n10644), .ZN(n13026) );
  NAND2_X1 U12018 ( .A1(n16896), .A2(n13057), .ZN(n9923) );
  NOR2_X1 U12019 ( .A1(n9925), .A2(n18091), .ZN(n10412) );
  NAND2_X1 U12020 ( .A1(n16917), .A2(n9778), .ZN(n10334) );
  INV_X1 U12021 ( .A(n10213), .ZN(n10212) );
  OAI21_X1 U12022 ( .B1(n9792), .B2(n10216), .A(n10214), .ZN(n10213) );
  NAND2_X1 U12023 ( .A1(n10638), .A2(n10215), .ZN(n10214) );
  INV_X1 U12024 ( .A(n16961), .ZN(n10215) );
  NAND2_X1 U12025 ( .A1(n10007), .A2(n10006), .ZN(n10005) );
  NAND2_X1 U12026 ( .A1(n16813), .A2(n20277), .ZN(n10006) );
  NAND2_X1 U12027 ( .A1(n10355), .A2(n10008), .ZN(n10007) );
  AOI21_X1 U12028 ( .B1(n10009), .B2(n10357), .A(n9737), .ZN(n10008) );
  NAND2_X1 U12029 ( .A1(n10207), .A2(n10206), .ZN(n10209) );
  INV_X1 U12030 ( .A(n10216), .ZN(n10206) );
  NOR2_X1 U12031 ( .A1(n10211), .A2(n10217), .ZN(n10210) );
  INV_X1 U12032 ( .A(n9792), .ZN(n10211) );
  NAND2_X1 U12033 ( .A1(n10009), .A2(n11495), .ZN(n10169) );
  NAND2_X1 U12034 ( .A1(n17021), .A2(n9856), .ZN(n10166) );
  XNOR2_X1 U12035 ( .A(n13500), .B(n13499), .ZN(n14788) );
  INV_X1 U12036 ( .A(n16984), .ZN(n10436) );
  OAI21_X1 U12037 ( .B1(n10609), .B2(n10226), .A(n10224), .ZN(n16984) );
  NAND2_X1 U12038 ( .A1(n10068), .A2(n10067), .ZN(n17306) );
  AND2_X1 U12039 ( .A1(n17316), .A2(n9838), .ZN(n10067) );
  NAND2_X1 U12040 ( .A1(n17295), .A2(n9765), .ZN(n10068) );
  NAND2_X1 U12041 ( .A1(n10609), .A2(n10384), .ZN(n10229) );
  NAND2_X1 U12042 ( .A1(n11523), .A2(n11467), .ZN(n20259) );
  INV_X1 U12043 ( .A(n17301), .ZN(n9954) );
  NAND2_X1 U12044 ( .A1(n17022), .A2(n17015), .ZN(n9955) );
  INV_X1 U12045 ( .A(n20259), .ZN(n20280) );
  INV_X1 U12046 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20919) );
  INV_X1 U12047 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20909) );
  INV_X1 U12048 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20900) );
  INV_X1 U12049 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n21853) );
  INV_X1 U12050 ( .A(n17696), .ZN(n20180) );
  INV_X1 U12051 ( .A(n10377), .ZN(n18937) );
  INV_X1 U12052 ( .A(n18211), .ZN(n10509) );
  OR2_X1 U12053 ( .A1(n11718), .A2(n11717), .ZN(n18568) );
  INV_X1 U12054 ( .A(n18540), .ZN(n18558) );
  INV_X1 U12055 ( .A(n18568), .ZN(n18581) );
  NAND2_X1 U12056 ( .A1(n14253), .A2(n18892), .ZN(n18879) );
  NOR2_X1 U12057 ( .A1(n9783), .A2(n10249), .ZN(n10248) );
  OAI21_X1 U12058 ( .B1(n17770), .B2(n17759), .A(n10250), .ZN(n10249) );
  INV_X1 U12059 ( .A(n10540), .ZN(n10324) );
  INV_X1 U12060 ( .A(n15393), .ZN(n10364) );
  AOI21_X1 U12061 ( .B1(n10396), .B2(n10635), .A(n10360), .ZN(n10362) );
  INV_X1 U12062 ( .A(n10637), .ZN(n10360) );
  INV_X1 U12063 ( .A(n11875), .ZN(n13145) );
  AOI22_X1 U12064 ( .A1(n10696), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n16445), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10689) );
  NAND2_X1 U12065 ( .A1(n10302), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n16451) );
  NAND2_X1 U12066 ( .A1(n10302), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n16457) );
  NAND2_X1 U12067 ( .A1(n9911), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n9886) );
  NAND2_X1 U12068 ( .A1(n17520), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n9863) );
  NAND2_X1 U12069 ( .A1(n9912), .A2(n9865), .ZN(n10925) );
  OAI21_X1 U12070 ( .B1(n20385), .B2(n10923), .A(n9885), .ZN(n10924) );
  NAND2_X1 U12071 ( .A1(n10286), .A2(n10285), .ZN(n10935) );
  NAND3_X1 U12072 ( .A1(n9910), .A2(n9905), .A3(n9904), .ZN(n9909) );
  NAND2_X1 U12073 ( .A1(n9898), .A2(n9910), .ZN(n9897) );
  NAND2_X1 U12074 ( .A1(n9902), .A2(n9775), .ZN(n9900) );
  AND2_X1 U12075 ( .A1(n11002), .A2(n11001), .ZN(n11007) );
  AND2_X1 U12076 ( .A1(n20919), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11033) );
  OAI21_X1 U12077 ( .B1(n12638), .B2(P1_EBX_REG_1__SCAN_IN), .A(n12650), .ZN(
        n12639) );
  CLKBUF_X1 U12078 ( .A(n11950), .Z(n12500) );
  INV_X1 U12079 ( .A(n13116), .ZN(n10046) );
  NAND2_X1 U12080 ( .A1(n13116), .A2(n18034), .ZN(n10311) );
  OR2_X1 U12081 ( .A1(n12016), .A2(n12015), .ZN(n13118) );
  OR2_X1 U12082 ( .A1(n12002), .A2(n12001), .ZN(n13108) );
  INV_X1 U12083 ( .A(n11984), .ZN(n13098) );
  INV_X1 U12084 ( .A(n10323), .ZN(n10322) );
  AOI21_X1 U12085 ( .B1(n11969), .B2(n20939), .A(n11968), .ZN(n11990) );
  AOI22_X1 U12086 ( .A1(n11995), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9691), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11835) );
  INV_X1 U12087 ( .A(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11817) );
  NAND2_X1 U12088 ( .A1(n10302), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n16587) );
  NAND2_X1 U12089 ( .A1(n10302), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n16595) );
  NAND2_X1 U12090 ( .A1(n10302), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n16550) );
  NAND2_X1 U12091 ( .A1(n10302), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n16556) );
  NAND2_X1 U12092 ( .A1(n10302), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n16522) );
  NAND2_X1 U12093 ( .A1(n10302), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n16528) );
  NAND2_X1 U12094 ( .A1(n10302), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n16507) );
  NAND2_X1 U12095 ( .A1(n10302), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n16513) );
  NAND2_X1 U12096 ( .A1(n10302), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n16483) );
  NAND2_X1 U12097 ( .A1(n10302), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n16491) );
  NAND3_X1 U12098 ( .A1(n9728), .A2(n10125), .A3(n10629), .ZN(n11006) );
  INV_X1 U12099 ( .A(n13001), .ZN(n10592) );
  NAND2_X1 U12100 ( .A1(n12946), .A2(n10594), .ZN(n10593) );
  INV_X1 U12101 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n10594) );
  NAND2_X1 U12102 ( .A1(n9751), .A2(n16946), .ZN(n10601) );
  INV_X1 U12103 ( .A(n16985), .ZN(n10223) );
  INV_X1 U12104 ( .A(n9949), .ZN(n9948) );
  NAND2_X1 U12105 ( .A1(n11518), .A2(n9962), .ZN(n9961) );
  NOR2_X1 U12106 ( .A1(n9963), .A2(n9965), .ZN(n9962) );
  INV_X1 U12107 ( .A(n17045), .ZN(n11086) );
  INV_X1 U12108 ( .A(n10605), .ZN(n10270) );
  OAI21_X1 U12109 ( .B1(n20385), .B2(n10959), .A(n9916), .ZN(n10960) );
  NAND2_X1 U12110 ( .A1(n9887), .A2(n9864), .ZN(n10961) );
  NAND2_X1 U12111 ( .A1(n10289), .A2(n10287), .ZN(n10970) );
  INV_X1 U12112 ( .A(n10347), .ZN(n10346) );
  OAI21_X1 U12113 ( .B1(n17140), .B2(n10348), .A(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n10347) );
  NAND2_X1 U12114 ( .A1(n9914), .A2(n9913), .ZN(n10814) );
  NAND2_X1 U12115 ( .A1(n9794), .A2(n14230), .ZN(n10811) );
  NAND2_X1 U12116 ( .A1(n9764), .A2(n9889), .ZN(n9918) );
  AOI22_X1 U12117 ( .A1(n17500), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n16614), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10670) );
  XNOR2_X1 U12118 ( .A(n17650), .B(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11017) );
  AND3_X1 U12119 ( .A1(n14747), .A2(n10252), .A3(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11549) );
  NAND2_X1 U12120 ( .A1(n11549), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13229) );
  AND2_X1 U12121 ( .A1(n11692), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13332) );
  AOI21_X1 U12122 ( .B1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n19560), .A(
        n11708), .ZN(n11711) );
  INV_X1 U12123 ( .A(n14714), .ZN(n13340) );
  OR2_X1 U12124 ( .A1(n9701), .A2(n11783), .ZN(n11787) );
  INV_X1 U12125 ( .A(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11783) );
  NAND2_X1 U12126 ( .A1(n11892), .A2(n14822), .ZN(n11893) );
  AND3_X1 U12127 ( .A1(n13459), .A2(n13953), .A3(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n11900) );
  NOR2_X1 U12128 ( .A1(n14889), .A2(n10551), .ZN(n10550) );
  INV_X1 U12129 ( .A(n14903), .ZN(n10551) );
  NAND2_X1 U12130 ( .A1(n10552), .A2(n10276), .ZN(n10275) );
  INV_X1 U12131 ( .A(n14944), .ZN(n10276) );
  NOR2_X1 U12132 ( .A1(n14958), .A2(n10553), .ZN(n10552) );
  NAND2_X1 U12133 ( .A1(n12112), .A2(n10234), .ZN(n10231) );
  NAND2_X1 U12134 ( .A1(n12054), .A2(n10233), .ZN(n10232) );
  NAND2_X1 U12135 ( .A1(n12103), .A2(n12112), .ZN(n10230) );
  AND2_X1 U12136 ( .A1(n13432), .A2(n13454), .ZN(n13418) );
  NOR2_X1 U12137 ( .A1(n15548), .A2(n15547), .ZN(n10106) );
  NAND2_X1 U12138 ( .A1(n10532), .A2(n12719), .ZN(n10531) );
  NAND2_X1 U12139 ( .A1(n10367), .A2(n10056), .ZN(n10055) );
  INV_X1 U12140 ( .A(n10311), .ZN(n10310) );
  OR2_X1 U12141 ( .A1(n12029), .A2(n12028), .ZN(n13129) );
  INV_X1 U12142 ( .A(n12118), .ZN(n12032) );
  NAND2_X1 U12143 ( .A1(n10135), .A2(n10547), .ZN(n12119) );
  INV_X1 U12144 ( .A(n12103), .ZN(n10135) );
  AND2_X1 U12145 ( .A1(n12657), .A2(n12656), .ZN(n14416) );
  INV_X1 U12146 ( .A(n11874), .ZN(n12086) );
  AND2_X1 U12147 ( .A1(n10514), .A2(n14403), .ZN(n13127) );
  OR2_X1 U12148 ( .A1(n12085), .A2(n12084), .ZN(n13089) );
  OR2_X1 U12149 ( .A1(n12045), .A2(n12044), .ZN(n13131) );
  OR2_X1 U12150 ( .A1(n11942), .A2(n11941), .ZN(n13109) );
  INV_X1 U12151 ( .A(n11907), .ZN(n11908) );
  AND3_X1 U12152 ( .A1(n13458), .A2(n13457), .A3(n13456), .ZN(n13948) );
  INV_X1 U12153 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n15945) );
  AOI22_X1 U12154 ( .A1(n11818), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11792), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11755) );
  AOI21_X1 U12155 ( .B1(n12619), .B2(n12616), .A(n12615), .ZN(n12617) );
  NAND2_X1 U12156 ( .A1(n9982), .A2(n9758), .ZN(n9980) );
  OAI22_X1 U12157 ( .A1(n12614), .A2(n12629), .B1(P1_STATE2_REG_0__SCAN_IN), 
        .B2(n12613), .ZN(n12615) );
  NAND2_X1 U12158 ( .A1(n12592), .A2(n9982), .ZN(n9981) );
  INV_X1 U12159 ( .A(n12608), .ZN(n12619) );
  XNOR2_X1 U12160 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11139) );
  INV_X1 U12161 ( .A(n11094), .ZN(n11093) );
  NAND2_X1 U12162 ( .A1(n11089), .A2(n9725), .ZN(n11100) );
  OR2_X1 U12163 ( .A1(n10985), .A2(n10984), .ZN(n11025) );
  NAND2_X1 U12164 ( .A1(n10307), .A2(n10306), .ZN(n11055) );
  NAND2_X1 U12165 ( .A1(n13010), .A2(P2_EBX_REG_5__SCAN_IN), .ZN(n10306) );
  NAND2_X1 U12166 ( .A1(n11022), .A2(n11012), .ZN(n10307) );
  OAI211_X1 U12167 ( .C1(n10726), .C2(n20829), .A(n10755), .B(n9927), .ZN(
        n10756) );
  NAND2_X1 U12168 ( .A1(n10773), .A2(P2_EBX_REG_1__SCAN_IN), .ZN(n9927) );
  INV_X1 U12169 ( .A(n16536), .ZN(n16563) );
  INV_X1 U12170 ( .A(n10758), .ZN(n10316) );
  NAND3_X1 U12171 ( .A1(n10312), .A2(n10313), .A3(n10317), .ZN(n10785) );
  NAND2_X1 U12172 ( .A1(n10766), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10317) );
  CLKBUF_X1 U12173 ( .A(n16447), .Z(n16489) );
  NAND2_X1 U12174 ( .A1(n10302), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n16571) );
  NAND2_X1 U12175 ( .A1(n10302), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n16577) );
  INV_X1 U12176 ( .A(n16503), .ZN(n10454) );
  INV_X1 U12177 ( .A(n16654), .ZN(n10457) );
  INV_X1 U12178 ( .A(n10733), .ZN(n12786) );
  AND2_X1 U12179 ( .A1(n14035), .A2(n17984), .ZN(n16536) );
  NAND2_X1 U12180 ( .A1(n10632), .A2(n9742), .ZN(n12913) );
  NAND2_X1 U12181 ( .A1(n11426), .A2(n10472), .ZN(n10471) );
  INV_X1 U12182 ( .A(n16222), .ZN(n10472) );
  INV_X1 U12183 ( .A(n11006), .ZN(n11504) );
  INV_X1 U12184 ( .A(n9857), .ZN(n10625) );
  OR2_X1 U12185 ( .A1(n10997), .A2(n10996), .ZN(n11072) );
  NOR2_X1 U12186 ( .A1(n13029), .A2(n13028), .ZN(n13030) );
  NAND2_X1 U12187 ( .A1(n16926), .A2(n10602), .ZN(n10329) );
  INV_X1 U12188 ( .A(n10421), .ZN(n9868) );
  INV_X1 U12189 ( .A(n16080), .ZN(n10562) );
  OR2_X1 U12190 ( .A1(n16103), .A2(n16082), .ZN(n10484) );
  NAND2_X1 U12191 ( .A1(n10486), .A2(n16665), .ZN(n10485) );
  INV_X1 U12192 ( .A(n9845), .ZN(n10486) );
  NAND2_X1 U12193 ( .A1(n9870), .A2(n10421), .ZN(n16931) );
  NAND2_X1 U12194 ( .A1(n16140), .A2(n10568), .ZN(n11383) );
  AND2_X1 U12195 ( .A1(n10569), .A2(n10634), .ZN(n10568) );
  AND2_X1 U12196 ( .A1(n16142), .A2(n16126), .ZN(n10571) );
  INV_X1 U12197 ( .A(n10224), .ZN(n10221) );
  NAND2_X1 U12198 ( .A1(n11443), .A2(n10483), .ZN(n10482) );
  INV_X1 U12199 ( .A(n16161), .ZN(n10483) );
  INV_X1 U12200 ( .A(n16182), .ZN(n11443) );
  NOR2_X1 U12201 ( .A1(n10566), .A2(n10565), .ZN(n10564) );
  INV_X1 U12202 ( .A(n14752), .ZN(n10565) );
  NAND2_X1 U12203 ( .A1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n10300) );
  NAND2_X1 U12204 ( .A1(n9950), .A2(n17082), .ZN(n17057) );
  AND2_X1 U12205 ( .A1(n11047), .A2(n10426), .ZN(n10425) );
  NAND2_X1 U12206 ( .A1(n16314), .A2(n13049), .ZN(n10426) );
  INV_X1 U12207 ( .A(n16314), .ZN(n10427) );
  OR2_X1 U12208 ( .A1(n10901), .A2(n10900), .ZN(n11246) );
  OAI21_X1 U12209 ( .B1(n10770), .B2(n21853), .A(n10769), .ZN(n10777) );
  AND2_X1 U12210 ( .A1(n10720), .A2(n11212), .ZN(n10729) );
  OAI22_X1 U12211 ( .A1(n12775), .A2(n11224), .B1(n12774), .B2(n14054), .ZN(
        n11225) );
  AND2_X1 U12212 ( .A1(n10580), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n17468) );
  NOR2_X1 U12213 ( .A1(n10719), .A2(n11011), .ZN(n10071) );
  OR2_X1 U12214 ( .A1(n16563), .A2(n20299), .ZN(n14076) );
  NAND2_X1 U12215 ( .A1(n14068), .A2(n14217), .ZN(n14070) );
  AND2_X1 U12216 ( .A1(n16536), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n14071) );
  AND2_X1 U12217 ( .A1(n16536), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n14224) );
  AND2_X1 U12218 ( .A1(n11155), .A2(n11154), .ZN(n11175) );
  OR2_X1 U12219 ( .A1(n11153), .A2(n11152), .ZN(n11155) );
  AND3_X1 U12220 ( .A1(n11470), .A2(n9790), .A3(n11177), .ZN(n17458) );
  OR2_X1 U12221 ( .A1(n11172), .A2(n17564), .ZN(n9890) );
  NAND2_X1 U12222 ( .A1(n10801), .A2(n10805), .ZN(n20436) );
  NAND2_X1 U12223 ( .A1(n10817), .A2(n14079), .ZN(n10915) );
  INV_X1 U12224 ( .A(n10954), .ZN(n20657) );
  OR2_X1 U12225 ( .A1(n11153), .A2(n11154), .ZN(n11198) );
  XNOR2_X1 U12226 ( .A(n11535), .B(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n11536) );
  AND2_X1 U12227 ( .A1(n10505), .A2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10504) );
  NOR2_X1 U12228 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11559) );
  INV_X1 U12229 ( .A(n19192), .ZN(n17849) );
  NAND2_X1 U12230 ( .A1(n17832), .A2(n19445), .ZN(n10493) );
  NAND2_X1 U12231 ( .A1(n13386), .A2(n10247), .ZN(n19188) );
  NOR2_X1 U12232 ( .A1(n13388), .A2(n19485), .ZN(n10245) );
  INV_X1 U12233 ( .A(n10256), .ZN(n10255) );
  INV_X1 U12234 ( .A(n14313), .ZN(n13354) );
  OR2_X1 U12235 ( .A1(n11627), .A2(n11626), .ZN(n11677) );
  INV_X1 U12236 ( .A(n14802), .ZN(n14796) );
  NAND2_X1 U12237 ( .A1(n11861), .A2(n14385), .ZN(n14136) );
  INV_X1 U12238 ( .A(n14102), .ZN(n21071) );
  INV_X1 U12239 ( .A(n12539), .ZN(n12540) );
  NAND2_X1 U12240 ( .A1(n12441), .A2(n9718), .ZN(n12519) );
  NAND2_X1 U12241 ( .A1(n12518), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12539) );
  INV_X1 U12242 ( .A(n12519), .ZN(n12518) );
  NAND2_X1 U12243 ( .A1(n12460), .A2(n12459), .ZN(n14876) );
  OR2_X1 U12244 ( .A1(n15331), .A2(n12631), .ZN(n12460) );
  AND2_X1 U12245 ( .A1(n12415), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12416) );
  AND2_X1 U12246 ( .A1(n12367), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12368) );
  INV_X1 U12247 ( .A(n12366), .ZN(n12367) );
  NOR2_X1 U12248 ( .A1(n12332), .A2(n15388), .ZN(n12333) );
  NAND2_X1 U12249 ( .A1(n12333), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12366) );
  NAND2_X1 U12250 ( .A1(n14981), .A2(n10554), .ZN(n10553) );
  INV_X1 U12251 ( .A(n14994), .ZN(n10554) );
  NAND2_X1 U12252 ( .A1(n12244), .A2(n9744), .ZN(n12300) );
  INV_X1 U12253 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n12299) );
  CLKBUF_X1 U12254 ( .A(n15007), .Z(n15008) );
  AND4_X1 U12255 ( .A1(n12141), .A2(n12140), .A3(n12139), .A4(n12138), .ZN(
        n15130) );
  NOR2_X1 U12256 ( .A1(n12113), .A2(n10138), .ZN(n10136) );
  AND2_X1 U12257 ( .A1(n10139), .A2(n10141), .ZN(n12122) );
  NOR2_X1 U12258 ( .A1(n12048), .A2(n10142), .ZN(n10139) );
  CLKBUF_X1 U12259 ( .A(n14570), .Z(n14571) );
  NOR2_X1 U12260 ( .A1(n12113), .A2(n12048), .ZN(n12120) );
  NOR2_X1 U12261 ( .A1(n10535), .A2(n14810), .ZN(n10371) );
  AND2_X1 U12262 ( .A1(n10106), .A2(n13412), .ZN(n10105) );
  NOR2_X2 U12263 ( .A1(n14862), .A2(n12733), .ZN(n14844) );
  AND2_X1 U12264 ( .A1(n12722), .A2(n12721), .ZN(n14877) );
  INV_X1 U12265 ( .A(n15336), .ZN(n10061) );
  NOR2_X1 U12266 ( .A1(n14954), .A2(n10530), .ZN(n14925) );
  INV_X1 U12267 ( .A(n10532), .ZN(n10530) );
  AND2_X1 U12268 ( .A1(n12709), .A2(n12708), .ZN(n14932) );
  NOR2_X1 U12269 ( .A1(n14954), .A2(n14932), .ZN(n14934) );
  NAND2_X1 U12270 ( .A1(n21137), .A2(n15594), .ZN(n15614) );
  AND2_X1 U12271 ( .A1(n12697), .A2(n12696), .ZN(n14982) );
  AND2_X1 U12272 ( .A1(n9819), .A2(n10525), .ZN(n10524) );
  NOR2_X1 U12273 ( .A1(n15024), .A2(n15010), .ZN(n10525) );
  NAND2_X1 U12274 ( .A1(n9939), .A2(n13141), .ZN(n15415) );
  INV_X1 U12275 ( .A(n15427), .ZN(n9939) );
  NAND2_X1 U12276 ( .A1(n15074), .A2(n9819), .ZN(n15039) );
  NOR2_X1 U12277 ( .A1(n15442), .A2(n13074), .ZN(n15426) );
  AND2_X1 U12278 ( .A1(n15074), .A2(n15056), .ZN(n15057) );
  NAND2_X1 U12279 ( .A1(n13076), .A2(n13072), .ZN(n15442) );
  AND2_X1 U12280 ( .A1(n12679), .A2(n12678), .ZN(n15090) );
  OR2_X1 U12281 ( .A1(n15103), .A2(n15090), .ZN(n15092) );
  NAND2_X1 U12282 ( .A1(n15121), .A2(n15101), .ZN(n15103) );
  AND2_X1 U12283 ( .A1(n12668), .A2(n12667), .ZN(n15133) );
  NAND2_X1 U12284 ( .A1(n9694), .A2(n21104), .ZN(n10052) );
  NAND2_X1 U12285 ( .A1(n21090), .A2(n10042), .ZN(n10053) );
  AND2_X1 U12286 ( .A1(n12660), .A2(n12659), .ZN(n14575) );
  AND2_X1 U12287 ( .A1(n13953), .A2(n20939), .ZN(n13153) );
  NAND2_X1 U12288 ( .A1(n11906), .A2(n10514), .ZN(n10359) );
  AND2_X1 U12290 ( .A1(n12654), .A2(n12653), .ZN(n14271) );
  OR2_X1 U12291 ( .A1(n14266), .A2(n14265), .ZN(n14270) );
  NOR2_X1 U12292 ( .A1(n14266), .A2(n10522), .ZN(n14417) );
  NAND2_X1 U12293 ( .A1(n10523), .A2(n12648), .ZN(n10522) );
  NAND3_X1 U12294 ( .A1(n10096), .A2(n10099), .A3(n10101), .ZN(n14274) );
  INV_X1 U12295 ( .A(n12568), .ZN(n12606) );
  INV_X1 U12296 ( .A(n14363), .ZN(n21181) );
  NAND2_X1 U12297 ( .A1(n11965), .A2(n11964), .ZN(n12069) );
  NAND2_X1 U12298 ( .A1(n9936), .A2(n9935), .ZN(n11965) );
  NAND2_X1 U12299 ( .A1(n11963), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n9935) );
  INV_X1 U12300 ( .A(n13148), .ZN(n11856) );
  NOR2_X1 U12301 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n13953) );
  INV_X1 U12302 ( .A(n21354), .ZN(n21267) );
  NOR2_X1 U12303 ( .A1(n14363), .A2(n21413), .ZN(n15847) );
  AND2_X1 U12304 ( .A1(n14363), .A2(n14364), .ZN(n21202) );
  INV_X1 U12305 ( .A(n15848), .ZN(n21355) );
  INV_X1 U12306 ( .A(n14389), .ZN(n14402) );
  NOR2_X2 U12307 ( .A1(n15511), .A2(n14801), .ZN(n14401) );
  INV_X1 U12308 ( .A(n14364), .ZN(n21413) );
  NAND2_X1 U12309 ( .A1(n18052), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15961) );
  INV_X1 U12310 ( .A(n18047), .ZN(n15763) );
  INV_X1 U12311 ( .A(n12846), .ZN(n17652) );
  INV_X1 U12312 ( .A(n10192), .ZN(n10191) );
  OAI21_X1 U12313 ( .B1(n12943), .B2(n16907), .A(n16898), .ZN(n10192) );
  AOI21_X1 U12314 ( .B1(n10188), .B2(n12943), .A(n12943), .ZN(n10187) );
  OR2_X1 U12315 ( .A1(n12927), .A2(n12943), .ZN(n10186) );
  NAND2_X1 U12316 ( .A1(n10200), .A2(n16956), .ZN(n10445) );
  NAND2_X1 U12317 ( .A1(n16336), .A2(n10446), .ZN(n16093) );
  INV_X1 U12318 ( .A(n10200), .ZN(n10446) );
  NAND2_X1 U12319 ( .A1(n16093), .A2(n16956), .ZN(n17998) );
  AND2_X1 U12320 ( .A1(n11380), .A2(n11379), .ZN(n14782) );
  NOR2_X1 U12321 ( .A1(n16218), .A2(n17039), .ZN(n16212) );
  OR2_X1 U12322 ( .A1(n13523), .A2(n17050), .ZN(n16218) );
  AND2_X1 U12323 ( .A1(n16249), .A2(n17074), .ZN(n16234) );
  NOR2_X1 U12324 ( .A1(n10595), .A2(n9743), .ZN(n10301) );
  NAND2_X1 U12325 ( .A1(n10195), .A2(n10194), .ZN(n16264) );
  INV_X1 U12326 ( .A(n18062), .ZN(n10194) );
  INV_X1 U12327 ( .A(n17113), .ZN(n10197) );
  NOR2_X1 U12328 ( .A1(n20200), .A2(n20201), .ZN(n10198) );
  INV_X1 U12329 ( .A(n16351), .ZN(n20190) );
  AND2_X1 U12330 ( .A1(n17145), .A2(n16334), .ZN(n16309) );
  NAND2_X1 U12331 ( .A1(n11500), .A2(n11012), .ZN(n10583) );
  NAND2_X1 U12332 ( .A1(n13010), .A2(n11013), .ZN(n11014) );
  AND2_X1 U12333 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12878) );
  OAI21_X1 U12334 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P2_STATE2_REG_0__SCAN_IN), .A(n10199), .ZN(n16332) );
  NAND2_X1 U12335 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n10199) );
  NOR2_X1 U12336 ( .A1(n17445), .A2(n16332), .ZN(n16334) );
  OR2_X1 U12337 ( .A1(n11303), .A2(n11302), .ZN(n16362) );
  NOR2_X1 U12338 ( .A1(n10574), .A2(n10573), .ZN(n10572) );
  NAND2_X1 U12339 ( .A1(n12962), .A2(n16019), .ZN(n10573) );
  NAND2_X1 U12340 ( .A1(n10302), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n16606) );
  INV_X1 U12341 ( .A(n16631), .ZN(n10465) );
  NOR2_X1 U12342 ( .A1(n16661), .A2(n16660), .ZN(n16659) );
  AND2_X1 U12343 ( .A1(n9837), .A2(n16409), .ZN(n9989) );
  INV_X1 U12344 ( .A(n10451), .ZN(n10450) );
  AND2_X1 U12345 ( .A1(n11214), .A2(n11213), .ZN(n11384) );
  OR2_X1 U12346 ( .A1(n16398), .A2(n16397), .ZN(n16687) );
  NAND2_X1 U12347 ( .A1(n9973), .A2(n9720), .ZN(n9972) );
  INV_X1 U12348 ( .A(n10730), .ZN(n12848) );
  INV_X1 U12349 ( .A(n11161), .ZN(n13855) );
  NOR3_X1 U12350 ( .A1(n9750), .A2(n10438), .A3(n10439), .ZN(n12870) );
  NAND2_X1 U12351 ( .A1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n10438) );
  NAND2_X1 U12352 ( .A1(n10342), .A2(n10340), .ZN(n10339) );
  OR2_X1 U12353 ( .A1(n16904), .A2(n10343), .ZN(n10342) );
  INV_X1 U12354 ( .A(n13053), .ZN(n10343) );
  AND2_X1 U12355 ( .A1(n12916), .A2(n9848), .ZN(n12931) );
  NAND2_X1 U12356 ( .A1(n12916), .A2(n9741), .ZN(n12928) );
  NAND2_X1 U12357 ( .A1(n12916), .A2(n10447), .ZN(n12925) );
  AND2_X1 U12358 ( .A1(n10632), .A2(n9835), .ZN(n12917) );
  AND2_X1 U12359 ( .A1(n12902), .A2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n10632) );
  INV_X1 U12360 ( .A(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n12903) );
  NAND2_X1 U12361 ( .A1(n12900), .A2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n12899) );
  INV_X1 U12362 ( .A(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n17037) );
  NOR2_X1 U12363 ( .A1(n12897), .A2(n17037), .ZN(n12900) );
  NAND2_X1 U12364 ( .A1(n10437), .A2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n12897) );
  INV_X1 U12365 ( .A(n12893), .ZN(n10437) );
  INV_X1 U12366 ( .A(n16252), .ZN(n10475) );
  NAND2_X1 U12367 ( .A1(n10442), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10441) );
  INV_X1 U12368 ( .A(n10444), .ZN(n10442) );
  NAND2_X1 U12369 ( .A1(n10443), .A2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12886) );
  INV_X1 U12370 ( .A(n12881), .ZN(n10443) );
  INV_X1 U12371 ( .A(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n17123) );
  NAND2_X1 U12372 ( .A1(n13020), .A2(n13019), .ZN(n13479) );
  NAND2_X1 U12373 ( .A1(n13003), .A2(n9727), .ZN(n10415) );
  NOR2_X1 U12374 ( .A1(n10417), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n10095) );
  NOR2_X1 U12375 ( .A1(n13052), .A2(n16916), .ZN(n10344) );
  INV_X1 U12376 ( .A(n9760), .ZN(n10340) );
  CLKBUF_X1 U12377 ( .A(n16048), .Z(n16049) );
  NOR3_X1 U12378 ( .A1(n16102), .A2(n16103), .A3(n9845), .ZN(n12811) );
  INV_X1 U12379 ( .A(n13027), .ZN(n16944) );
  OR2_X1 U12380 ( .A1(n10403), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10354) );
  NAND2_X1 U12381 ( .A1(n10217), .A2(n16961), .ZN(n10216) );
  INV_X1 U12382 ( .A(n10638), .ZN(n10217) );
  NOR2_X1 U12383 ( .A1(n16102), .A2(n16103), .ZN(n16101) );
  CLKBUF_X1 U12384 ( .A(n11383), .Z(n16100) );
  OR2_X1 U12385 ( .A1(n9748), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n10170) );
  AND2_X1 U12386 ( .A1(n11375), .A2(n11374), .ZN(n16159) );
  INV_X1 U12387 ( .A(n16998), .ZN(n10382) );
  INV_X1 U12388 ( .A(n16192), .ZN(n11438) );
  AND2_X1 U12389 ( .A1(n17341), .A2(n14771), .ZN(n17313) );
  AND3_X1 U12390 ( .A1(n11373), .A2(n11372), .A3(n11371), .ZN(n14760) );
  CLKBUF_X1 U12391 ( .A(n14749), .Z(n14750) );
  AND2_X1 U12392 ( .A1(n17325), .A2(n17394), .ZN(n17341) );
  AND3_X1 U12393 ( .A1(n11347), .A2(n11346), .A3(n11345), .ZN(n14755) );
  NOR2_X1 U12394 ( .A1(n13526), .A2(n10566), .ZN(n14751) );
  OR2_X1 U12395 ( .A1(n10300), .A2(n17327), .ZN(n10299) );
  NAND2_X1 U12396 ( .A1(n10609), .A2(n10607), .ZN(n17033) );
  AND3_X1 U12397 ( .A1(n11332), .A2(n11331), .A3(n11330), .ZN(n14515) );
  NOR2_X1 U12398 ( .A1(n9791), .A2(n9921), .ZN(n9920) );
  INV_X1 U12399 ( .A(n14083), .ZN(n9921) );
  AND3_X1 U12400 ( .A1(n11293), .A2(n11292), .A3(n11291), .ZN(n14244) );
  OR2_X1 U12401 ( .A1(n14082), .A2(n10577), .ZN(n14359) );
  NAND2_X1 U12402 ( .A1(n11518), .A2(n9963), .ZN(n9960) );
  INV_X1 U12403 ( .A(n18056), .ZN(n10624) );
  AND2_X1 U12404 ( .A1(n11075), .A2(n18055), .ZN(n18068) );
  INV_X1 U12405 ( .A(n14509), .ZN(n10476) );
  AND2_X1 U12406 ( .A1(n10092), .A2(n9818), .ZN(n11059) );
  AND3_X1 U12407 ( .A1(n11259), .A2(n11258), .A3(n11257), .ZN(n16298) );
  NAND2_X1 U12408 ( .A1(n10063), .A2(n11512), .ZN(n17121) );
  AND3_X1 U12409 ( .A1(n11254), .A2(n11253), .A3(n11252), .ZN(n16858) );
  INV_X1 U12410 ( .A(n11216), .ZN(n11217) );
  NAND2_X1 U12411 ( .A1(n14059), .A2(n14058), .ZN(n14061) );
  XNOR2_X1 U12412 ( .A(n14036), .B(n14076), .ZN(n14075) );
  NAND2_X1 U12413 ( .A1(n14073), .A2(n14214), .ZN(n14215) );
  OR2_X1 U12414 ( .A1(n14072), .A2(n14071), .ZN(n14073) );
  NAND2_X1 U12415 ( .A1(n9975), .A2(n14214), .ZN(n14227) );
  NAND2_X1 U12416 ( .A1(n9977), .A2(n9976), .ZN(n9975) );
  INV_X1 U12417 ( .A(n14215), .ZN(n9976) );
  INV_X1 U12418 ( .A(n14216), .ZN(n9977) );
  NOR2_X1 U12419 ( .A1(n10731), .A2(n10720), .ZN(n9991) );
  NAND2_X1 U12420 ( .A1(n20896), .A2(n17513), .ZN(n20497) );
  AND2_X1 U12421 ( .A1(n20896), .A2(n20903), .ZN(n20885) );
  INV_X1 U12422 ( .A(n10720), .ZN(n17564) );
  INV_X1 U12423 ( .A(n17590), .ZN(n17591) );
  INV_X1 U12424 ( .A(n17589), .ZN(n17592) );
  NOR2_X2 U12425 ( .A1(n17525), .A2(n17547), .ZN(n17590) );
  NOR2_X2 U12426 ( .A1(n12798), .A2(n17547), .ZN(n17589) );
  AND2_X1 U12427 ( .A1(n20748), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n17588) );
  NOR2_X1 U12428 ( .A1(n20535), .A2(n20691), .ZN(n20753) );
  AND2_X1 U12429 ( .A1(n11386), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12951) );
  NAND2_X1 U12430 ( .A1(n11173), .A2(n11188), .ZN(n17682) );
  NAND2_X1 U12431 ( .A1(n19568), .A2(n11712), .ZN(n13351) );
  NOR3_X1 U12432 ( .A1(n14321), .A2(n20041), .A3(n14153), .ZN(n20019) );
  NOR2_X1 U12433 ( .A1(n18218), .A2(n18219), .ZN(n18217) );
  AND2_X1 U12434 ( .A1(n18264), .A2(n10503), .ZN(n18255) );
  AND2_X1 U12435 ( .A1(n18287), .A2(n10503), .ZN(n18277) );
  NAND2_X1 U12436 ( .A1(n18518), .A2(n19058), .ZN(n10501) );
  NAND2_X1 U12437 ( .A1(n10500), .A2(n9788), .ZN(n10499) );
  INV_X1 U12438 ( .A(n19066), .ZN(n10502) );
  OR2_X1 U12439 ( .A1(n18312), .A2(n19066), .ZN(n18310) );
  INV_X1 U12440 ( .A(n20169), .ZN(n20166) );
  NOR2_X1 U12441 ( .A1(n18957), .A2(n21680), .ZN(n10374) );
  NOR2_X1 U12442 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11560) );
  NAND2_X1 U12443 ( .A1(n14731), .A2(n11557), .ZN(n13819) );
  AND2_X1 U12444 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11557) );
  OR2_X1 U12445 ( .A1(n13254), .A2(n13253), .ZN(n13362) );
  OR2_X1 U12446 ( .A1(n13239), .A2(n13238), .ZN(n13360) );
  OR2_X1 U12447 ( .A1(n13225), .A2(n13224), .ZN(n13296) );
  INV_X2 U12448 ( .A(n13819), .ZN(n13278) );
  AND2_X1 U12449 ( .A1(n14338), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11556) );
  AND2_X1 U12450 ( .A1(n19583), .A2(n17706), .ZN(n14714) );
  AOI21_X1 U12451 ( .B1(n19067), .B2(n10503), .A(n9843), .ZN(n10250) );
  NAND2_X1 U12452 ( .A1(n17778), .A2(n9739), .ZN(n17753) );
  AND2_X1 U12453 ( .A1(n17778), .A2(n11526), .ZN(n13400) );
  NAND2_X1 U12454 ( .A1(n11533), .A2(n9762), .ZN(n19054) );
  AND2_X1 U12455 ( .A1(n19387), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n19336) );
  INV_X1 U12456 ( .A(n19149), .ZN(n10510) );
  NOR2_X1 U12457 ( .A1(n18426), .A2(n17834), .ZN(n19146) );
  NAND2_X1 U12458 ( .A1(n17848), .A2(n19146), .ZN(n19147) );
  INV_X1 U12459 ( .A(n19238), .ZN(n18516) );
  NAND2_X1 U12460 ( .A1(n10021), .A2(n10020), .ZN(n17763) );
  AND2_X1 U12461 ( .A1(n10022), .A2(n13549), .ZN(n10020) );
  AND2_X1 U12462 ( .A1(n17741), .A2(n17899), .ZN(n10022) );
  NOR2_X1 U12463 ( .A1(n17929), .A2(n17765), .ZN(n17914) );
  INV_X1 U12464 ( .A(n13331), .ZN(n10024) );
  NAND2_X1 U12465 ( .A1(n18998), .A2(n13331), .ZN(n10491) );
  NAND2_X1 U12466 ( .A1(n19032), .A2(n17856), .ZN(n17929) );
  OR2_X1 U12467 ( .A1(n19042), .A2(n13359), .ZN(n17925) );
  OR2_X1 U12468 ( .A1(n19063), .A2(n19117), .ZN(n19090) );
  NAND2_X1 U12469 ( .A1(n10261), .A2(n9844), .ZN(n10260) );
  NOR2_X1 U12470 ( .A1(n14708), .A2(n14707), .ZN(n19387) );
  INV_X1 U12471 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n14707) );
  OR2_X1 U12472 ( .A1(n19172), .A2(n10493), .ZN(n19164) );
  INV_X1 U12473 ( .A(n13355), .ZN(n13979) );
  NAND2_X1 U12474 ( .A1(n11674), .A2(n14155), .ZN(n10375) );
  INV_X1 U12475 ( .A(n14321), .ZN(n10376) );
  AND2_X1 U12476 ( .A1(n11690), .A2(n11689), .ZN(n14312) );
  OR2_X1 U12477 ( .A1(n9752), .A2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n19172) );
  XNOR2_X1 U12478 ( .A(n13383), .B(n10241), .ZN(n19216) );
  INV_X1 U12479 ( .A(n13382), .ZN(n10241) );
  NAND2_X1 U12480 ( .A1(n19240), .A2(n13380), .ZN(n19224) );
  NAND2_X1 U12481 ( .A1(n19224), .A2(n19225), .ZN(n19223) );
  INV_X1 U12482 ( .A(n19546), .ZN(n19522) );
  OR2_X1 U12483 ( .A1(n13967), .A2(n13344), .ZN(n20016) );
  NOR2_X1 U12484 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n14731) );
  INV_X1 U12485 ( .A(n11687), .ZN(n19574) );
  INV_X1 U12486 ( .A(n11677), .ZN(n19577) );
  NOR2_X1 U12487 ( .A1(n13351), .A2(n11691), .ZN(n20041) );
  INV_X1 U12488 ( .A(n20982), .ZN(n15112) );
  NAND2_X1 U12489 ( .A1(n14099), .A2(n20935), .ZN(n15195) );
  OAI22_X1 U12490 ( .A1(n15971), .A2(n14434), .B1(n14098), .B2(n14131), .ZN(
        n14099) );
  OR2_X1 U12491 ( .A1(n15195), .A2(n14385), .ZN(n15203) );
  INV_X1 U12492 ( .A(n15195), .ZN(n15204) );
  OR2_X1 U12493 ( .A1(n14796), .A2(n14801), .ZN(n15258) );
  AND2_X1 U12494 ( .A1(n14802), .A2(n14801), .ZN(n15275) );
  OR2_X1 U12495 ( .A1(n14129), .A2(n14128), .ZN(n14134) );
  AND2_X1 U12496 ( .A1(n14796), .A2(n15272), .ZN(n15296) );
  OR3_X1 U12497 ( .A1(n14129), .A2(n13991), .A3(n13990), .ZN(n21060) );
  NOR2_X1 U12498 ( .A1(n15937), .A2(n13989), .ZN(n13991) );
  OAI21_X1 U12499 ( .B1(n14825), .B2(n14827), .A(n14826), .ZN(n15306) );
  INV_X1 U12500 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n15388) );
  CLKBUF_X1 U12501 ( .A(n14992), .Z(n14993) );
  NAND2_X1 U12502 ( .A1(n12244), .A2(n10149), .ZN(n12282) );
  NAND2_X1 U12503 ( .A1(n12244), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12262) );
  INV_X1 U12504 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n15451) );
  NAND2_X1 U12505 ( .A1(n12158), .A2(n10154), .ZN(n12203) );
  NAND2_X1 U12506 ( .A1(n12158), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12184) );
  INV_X1 U12507 ( .A(n15511), .ZN(n21094) );
  XNOR2_X1 U12508 ( .A(n10398), .B(n15303), .ZN(n15520) );
  OAI21_X1 U12509 ( .B1(n15317), .B2(n10400), .A(n10399), .ZN(n10398) );
  NAND2_X1 U12510 ( .A1(n15302), .A2(n10056), .ZN(n10399) );
  NAND2_X1 U12511 ( .A1(n9734), .A2(n15394), .ZN(n10400) );
  XNOR2_X1 U12512 ( .A(n10058), .B(n15572), .ZN(n15577) );
  NAND2_X1 U12513 ( .A1(n10060), .A2(n10059), .ZN(n10058) );
  NAND2_X1 U12514 ( .A1(n15336), .A2(n10056), .ZN(n10059) );
  OAI21_X1 U12515 ( .B1(n10061), .B2(n9693), .A(n15394), .ZN(n10060) );
  AOI21_X2 U12516 ( .B1(n21137), .B2(n13475), .A(n15603), .ZN(n15579) );
  OAI21_X1 U12517 ( .B1(n15359), .B2(n13143), .A(n15394), .ZN(n15350) );
  OAI21_X1 U12518 ( .B1(n15360), .B2(n13464), .A(n10056), .ZN(n15351) );
  NAND2_X1 U12519 ( .A1(n15494), .A2(n15493), .ZN(n10394) );
  INV_X1 U12520 ( .A(n15742), .ZN(n21121) );
  INV_X1 U12521 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n21147) );
  OAI21_X1 U12522 ( .B1(n14466), .B2(n18053), .A(n15796), .ZN(n21146) );
  CLKBUF_X1 U12523 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n15788) );
  NAND2_X1 U12524 ( .A1(n15971), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n21594) );
  INV_X1 U12525 ( .A(n21599), .ZN(n21597) );
  INV_X1 U12526 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n15807) );
  INV_X1 U12527 ( .A(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11812) );
  OR2_X1 U12528 ( .A1(n14373), .A2(n14364), .ZN(n21167) );
  OAI22_X1 U12529 ( .A1(n15804), .A2(n15803), .B1(n15813), .B2(n15853), .ZN(
        n21170) );
  OAI211_X1 U12530 ( .C1(n21376), .C2(n21301), .A(n14474), .B(n21422), .ZN(
        n14499) );
  AND2_X1 U12531 ( .A1(n15855), .A2(n15854), .ZN(n15892) );
  AND2_X1 U12532 ( .A1(n21268), .A2(n15812), .ZN(n15889) );
  INV_X1 U12533 ( .A(n21390), .ZN(n21933) );
  AOI22_X1 U12534 ( .A1(n15902), .A2(n15900), .B1(n15899), .B2(n21460), .ZN(
        n15932) );
  INV_X1 U12535 ( .A(n21303), .ZN(n21465) );
  INV_X1 U12536 ( .A(n21313), .ZN(n21481) );
  INV_X1 U12537 ( .A(n21397), .ZN(n21482) );
  AND2_X1 U12538 ( .A1(n14381), .A2(n14402), .ZN(n21928) );
  AND2_X1 U12539 ( .A1(n11874), .A2(n14402), .ZN(n21497) );
  INV_X1 U12540 ( .A(n21333), .ZN(n21509) );
  OAI211_X1 U12541 ( .C1(n21475), .C2(n21515), .A(n21474), .B(n21473), .ZN(
        n21521) );
  INV_X1 U12542 ( .A(n21476), .ZN(n21520) );
  OR2_X1 U12543 ( .A1(n15271), .A2(n15796), .ZN(n21394) );
  OR2_X1 U12544 ( .A1(n15261), .A2(n15796), .ZN(n21936) );
  INV_X1 U12545 ( .A(n21491), .ZN(n21321) );
  INV_X1 U12546 ( .A(n21492), .ZN(n21400) );
  OR2_X1 U12547 ( .A1(n15251), .A2(n15796), .ZN(n21403) );
  INV_X1 U12548 ( .A(n21503), .ZN(n21329) );
  OR2_X1 U12549 ( .A1(n15246), .A2(n15796), .ZN(n21406) );
  OR2_X1 U12550 ( .A1(n15242), .A2(n15796), .ZN(n21409) );
  INV_X1 U12551 ( .A(n21516), .ZN(n21337) );
  OR2_X1 U12552 ( .A1(n15297), .A2(n15796), .ZN(n21412) );
  OAI21_X1 U12553 ( .B1(n14375), .B2(n14374), .A(n21422), .ZN(n14407) );
  INV_X1 U12554 ( .A(n21167), .ZN(n15790) );
  AND2_X1 U12555 ( .A1(n15965), .A2(n18046), .ZN(n15973) );
  INV_X1 U12556 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n18052) );
  INV_X1 U12557 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n20939) );
  INV_X1 U12558 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n20691) );
  NOR2_X1 U12559 ( .A1(n17668), .A2(n11189), .ZN(n20921) );
  INV_X1 U12560 ( .A(n15989), .ZN(n16009) );
  AND2_X1 U12561 ( .A1(n11132), .A2(n11131), .ZN(n16097) );
  NAND2_X1 U12562 ( .A1(n16336), .A2(n12915), .ZN(n16105) );
  NAND2_X1 U12563 ( .A1(n11089), .A2(n9763), .ZN(n11105) );
  NAND2_X1 U12564 ( .A1(n16234), .A2(n17062), .ZN(n13523) );
  INV_X1 U12565 ( .A(n20189), .ZN(n16178) );
  INV_X1 U12566 ( .A(n10198), .ZN(n20203) );
  NAND2_X1 U12567 ( .A1(n15982), .A2(n12950), .ZN(n20192) );
  AND2_X1 U12568 ( .A1(n16351), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20189) );
  INV_X1 U12569 ( .A(n20196), .ZN(n16354) );
  OR2_X1 U12570 ( .A1(n11343), .A2(n11342), .ZN(n16711) );
  INV_X1 U12571 ( .A(n16359), .ZN(n16715) );
  OR2_X1 U12572 ( .A1(n11316), .A2(n11315), .ZN(n16719) );
  INV_X1 U12573 ( .A(n16362), .ZN(n16724) );
  OR2_X1 U12574 ( .A1(n11276), .A2(n11275), .ZN(n16739) );
  INV_X1 U12575 ( .A(n16733), .ZN(n16737) );
  INV_X1 U12576 ( .A(n20903), .ZN(n17513) );
  INV_X2 U12577 ( .A(n16728), .ZN(n16723) );
  OR2_X1 U12578 ( .A1(n16723), .A2(n11170), .ZN(n16733) );
  NAND2_X1 U12579 ( .A1(n10466), .A2(n16631), .ZN(n16627) );
  AND2_X1 U12580 ( .A1(n16872), .A2(n16855), .ZN(n16864) );
  INV_X1 U12581 ( .A(n16855), .ZN(n16868) );
  AND2_X1 U12582 ( .A1(n13854), .A2(n20812), .ZN(n20238) );
  INV_X1 U12583 ( .A(n20241), .ZN(n20242) );
  INV_X1 U12584 ( .A(n20238), .ZN(n20245) );
  AND2_X1 U12585 ( .A1(n13603), .A2(n13600), .ZN(n13677) );
  NAND2_X1 U12586 ( .A1(n9993), .A2(n9992), .ZN(n18086) );
  INV_X1 U12587 ( .A(n17467), .ZN(n14040) );
  OR2_X1 U12588 ( .A1(n17160), .A2(n20259), .ZN(n17171) );
  XNOR2_X1 U12589 ( .A(n10128), .B(n9768), .ZN(n17175) );
  NAND2_X1 U12590 ( .A1(n10129), .A2(n13015), .ZN(n10128) );
  NAND2_X1 U12591 ( .A1(n16912), .A2(n10418), .ZN(n10129) );
  NAND2_X1 U12592 ( .A1(n10184), .A2(n17188), .ZN(n10319) );
  INV_X1 U12593 ( .A(n16905), .ZN(n10184) );
  NAND2_X1 U12594 ( .A1(n9871), .A2(n9786), .ZN(n10031) );
  NAND2_X1 U12595 ( .A1(n16917), .A2(n10032), .ZN(n10030) );
  INV_X1 U12596 ( .A(n10036), .ZN(n10032) );
  INV_X1 U12597 ( .A(n10034), .ZN(n10033) );
  OAI21_X1 U12598 ( .B1(n10036), .B2(n10037), .A(n10035), .ZN(n10034) );
  NAND2_X1 U12599 ( .A1(n16893), .A2(n10039), .ZN(n10035) );
  AND2_X1 U12600 ( .A1(n10175), .A2(n17202), .ZN(n10406) );
  NAND2_X1 U12601 ( .A1(n16943), .A2(n17239), .ZN(n10073) );
  NOR2_X1 U12602 ( .A1(n16997), .A2(n11522), .ZN(n16968) );
  NAND2_X1 U12603 ( .A1(n10391), .A2(n16960), .ZN(n16964) );
  NOR2_X1 U12604 ( .A1(n20290), .A2(n10168), .ZN(n10167) );
  INV_X1 U12605 ( .A(n10170), .ZN(n10168) );
  AND2_X1 U12606 ( .A1(n10402), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n10079) );
  NAND2_X1 U12607 ( .A1(n10386), .A2(n10388), .ZN(n17001) );
  NAND2_X1 U12608 ( .A1(n10387), .A2(n10430), .ZN(n10386) );
  NAND2_X1 U12609 ( .A1(n17021), .A2(n10298), .ZN(n10297) );
  NOR2_X1 U12610 ( .A1(n10299), .A2(n10240), .ZN(n10298) );
  NOR2_X1 U12611 ( .A1(n17066), .A2(n17385), .ZN(n17060) );
  NAND2_X1 U12612 ( .A1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n10240), .ZN(
        n10239) );
  NAND2_X1 U12613 ( .A1(n17021), .A2(n10238), .ZN(n10176) );
  NOR2_X1 U12614 ( .A1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n10240), .ZN(
        n10238) );
  CLKBUF_X1 U12615 ( .A(n17096), .Z(n17097) );
  INV_X1 U12616 ( .A(n10617), .ZN(n17106) );
  NAND2_X1 U12617 ( .A1(n14352), .A2(n11242), .ZN(n14563) );
  NAND2_X1 U12618 ( .A1(n12846), .A2(n9943), .ZN(n11211) );
  AND2_X1 U12619 ( .A1(n11523), .A2(n17653), .ZN(n20275) );
  OR2_X1 U12620 ( .A1(n20275), .A2(n17294), .ZN(n14774) );
  NAND2_X1 U12621 ( .A1(n17451), .A2(n14027), .ZN(n20914) );
  INV_X1 U12622 ( .A(n20535), .ZN(n20890) );
  INV_X1 U12623 ( .A(n14036), .ZN(n17451) );
  AND2_X1 U12624 ( .A1(n17651), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n17685) );
  INV_X1 U12625 ( .A(n17990), .ZN(n17511) );
  OR2_X1 U12626 ( .A1(n20667), .A2(n20747), .ZN(n20310) );
  OAI21_X1 U12627 ( .B1(n20324), .B2(n20692), .A(n20323), .ZN(n20343) );
  NOR2_X1 U12628 ( .A1(n20476), .A2(n20350), .ZN(n20387) );
  NOR2_X2 U12629 ( .A1(n20439), .A2(n20350), .ZN(n20377) );
  OAI21_X1 U12630 ( .B1(n20360), .B2(n20356), .A(n20355), .ZN(n20379) );
  OAI21_X1 U12631 ( .B1(n17607), .B2(n17606), .A(n17605), .ZN(n20431) );
  NAND2_X1 U12632 ( .A1(n10615), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n17605) );
  NOR2_X1 U12633 ( .A1(n20476), .A2(n20747), .ZN(n20499) );
  OAI21_X1 U12634 ( .B1(n20887), .B2(n20475), .A(n20474), .ZN(n20494) );
  NOR2_X1 U12635 ( .A1(n20501), .A2(n9917), .ZN(n20502) );
  NOR2_X2 U12636 ( .A1(n20690), .A2(n20350), .ZN(n20597) );
  NOR2_X1 U12637 ( .A1(n17614), .A2(n10290), .ZN(n17615) );
  AOI21_X1 U12638 ( .B1(n20742), .B2(n17633), .A(n17632), .ZN(n20651) );
  OAI22_X1 U12639 ( .A1(n18110), .A2(n17592), .B1(n16787), .B2(n17591), .ZN(
        n20705) );
  OAI22_X1 U12640 ( .A1(n18100), .A2(n17592), .B1(n18178), .B2(n17591), .ZN(
        n20733) );
  AND2_X1 U12641 ( .A1(n20748), .A2(n17524), .ZN(n20746) );
  INV_X1 U12642 ( .A(n20708), .ZN(n20762) );
  AND2_X1 U12643 ( .A1(n17588), .A2(n17984), .ZN(n20760) );
  AND2_X1 U12644 ( .A1(n20748), .A2(n17558), .ZN(n20761) );
  INV_X1 U12645 ( .A(n20705), .ZN(n20765) );
  INV_X1 U12646 ( .A(n20713), .ZN(n20768) );
  AND2_X1 U12647 ( .A1(n20748), .A2(n17563), .ZN(n20767) );
  AND2_X1 U12648 ( .A1(n17588), .A2(n10731), .ZN(n20772) );
  AND2_X1 U12649 ( .A1(n20748), .A2(n17569), .ZN(n20773) );
  AND2_X1 U12650 ( .A1(n20748), .A2(n17574), .ZN(n20779) );
  INV_X1 U12651 ( .A(n20720), .ZN(n20786) );
  AND2_X1 U12652 ( .A1(n17588), .A2(n11012), .ZN(n20784) );
  AND2_X1 U12653 ( .A1(n20748), .A2(n17531), .ZN(n20785) );
  INV_X1 U12654 ( .A(n20726), .ZN(n20792) );
  AND2_X1 U12655 ( .A1(n20748), .A2(n17536), .ZN(n20791) );
  INV_X1 U12656 ( .A(n20738), .ZN(n20800) );
  INV_X1 U12657 ( .A(n20310), .ZN(n20801) );
  AND2_X1 U12658 ( .A1(n20748), .A2(n17587), .ZN(n20798) );
  INV_X1 U12659 ( .A(n20733), .ZN(n20806) );
  OR2_X1 U12660 ( .A1(n13065), .A2(n12944), .ZN(n17996) );
  NAND2_X1 U12661 ( .A1(n12951), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n17696) );
  INV_X1 U12662 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n20829) );
  NOR2_X1 U12663 ( .A1(n20019), .A2(n18935), .ZN(n20169) );
  NAND2_X1 U12664 ( .A1(n18192), .A2(n20018), .ZN(n18935) );
  NOR2_X1 U12665 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n18316), .ZN(n18302) );
  NAND2_X1 U12666 ( .A1(n10499), .A2(n10501), .ZN(n18300) );
  NOR2_X1 U12667 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n18337), .ZN(n18323) );
  NOR3_X1 U12668 ( .A1(n20093), .A2(n20091), .A3(n18406), .ZN(n18377) );
  NOR2_X1 U12669 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n18434), .ZN(n18415) );
  NOR2_X2 U12670 ( .A1(n20038), .A2(n11718), .ZN(n18551) );
  NOR2_X2 U12671 ( .A1(n20134), .A2(n18576), .ZN(n18540) );
  OAI211_X1 U12672 ( .C1(n20156), .C2(n20043), .A(n18481), .B(n20166), .ZN(
        n18564) );
  INV_X1 U12673 ( .A(n18564), .ZN(n18576) );
  INV_X1 U12674 ( .A(n18633), .ZN(n18643) );
  AND2_X1 U12675 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n18655), .ZN(n18649) );
  NOR2_X1 U12676 ( .A1(n18294), .A2(n18650), .ZN(n18655) );
  INV_X1 U12677 ( .A(n18782), .ZN(n18780) );
  INV_X1 U12678 ( .A(n18749), .ZN(n18777) );
  AND2_X1 U12679 ( .A1(n18818), .A2(n10373), .ZN(n18803) );
  AND2_X1 U12680 ( .A1(n9747), .A2(P3_EAX_REG_28__SCAN_IN), .ZN(n10373) );
  NAND2_X1 U12681 ( .A1(n18818), .A2(n9747), .ZN(n18808) );
  INV_X1 U12682 ( .A(n18823), .ZN(n18818) );
  NAND2_X1 U12683 ( .A1(n18818), .A2(P3_EAX_REG_25__SCAN_IN), .ZN(n18817) );
  NOR2_X1 U12684 ( .A1(n18828), .A2(n18787), .ZN(n18824) );
  NOR2_X1 U12685 ( .A1(n18859), .A2(n10378), .ZN(n18829) );
  INV_X1 U12686 ( .A(n18786), .ZN(n10379) );
  NAND2_X1 U12687 ( .A1(n18829), .A2(P3_EAX_REG_23__SCAN_IN), .ZN(n18828) );
  NOR2_X1 U12688 ( .A1(n18859), .A2(n18787), .ZN(n18854) );
  NAND2_X1 U12689 ( .A1(n18860), .A2(P3_EAX_REG_16__SCAN_IN), .ZN(n18859) );
  INV_X1 U12690 ( .A(n18788), .ZN(n18858) );
  NAND4_X1 U12691 ( .A1(n18878), .A2(P3_EAX_REG_14__SCAN_IN), .A3(
        P3_EAX_REG_13__SCAN_IN), .A4(n14299), .ZN(n18865) );
  AND2_X1 U12692 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n17737), .ZN(n17740) );
  NOR2_X1 U12693 ( .A1(n18980), .A2(n18879), .ZN(n18878) );
  INV_X1 U12694 ( .A(n18886), .ZN(n18877) );
  INV_X1 U12695 ( .A(n13274), .ZN(n10242) );
  OR2_X1 U12696 ( .A1(n18886), .A2(n14714), .ZN(n18883) );
  AND2_X1 U12697 ( .A1(n9682), .A2(n14714), .ZN(n18888) );
  NAND2_X1 U12698 ( .A1(n18930), .A2(n18934), .ZN(n18916) );
  NOR2_X1 U12699 ( .A1(n18935), .A2(n18894), .ZN(n18928) );
  AND2_X1 U12700 ( .A1(n11533), .A2(n9810), .ZN(n19002) );
  INV_X1 U12701 ( .A(n19021), .ZN(n10494) );
  INV_X1 U12702 ( .A(n19594), .ZN(n19945) );
  NAND2_X1 U12703 ( .A1(n19227), .A2(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n19217) );
  INV_X1 U12704 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n19218) );
  NOR2_X1 U12705 ( .A1(n21869), .A2(n19238), .ZN(n19227) );
  INV_X1 U12706 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n21869) );
  INV_X1 U12707 ( .A(n19877), .ZN(n19594) );
  INV_X1 U12708 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n19272) );
  INV_X1 U12709 ( .A(n19454), .ZN(n19314) );
  INV_X1 U12710 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n20151) );
  OR2_X1 U12711 ( .A1(n9752), .A2(n10262), .ZN(n19132) );
  INV_X1 U12712 ( .A(n10246), .ZN(n19200) );
  NAND2_X1 U12713 ( .A1(n19211), .A2(n19210), .ZN(n19213) );
  NAND2_X1 U12714 ( .A1(n10254), .A2(n13295), .ZN(n19235) );
  NAND2_X1 U12715 ( .A1(n19248), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10254) );
  AND2_X1 U12716 ( .A1(n13975), .A2(n18192), .ZN(n19546) );
  INV_X1 U12717 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n14747) );
  AOI211_X1 U12718 ( .C1(n18192), .C2(n19999), .A(n14327), .B(n19564), .ZN(
        n14748) );
  AND2_X1 U12719 ( .A1(n20036), .A2(n20035), .ZN(n20048) );
  INV_X1 U12720 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n20134) );
  AND2_X1 U12721 ( .A1(n13517), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n15223)
         );
  CLKBUF_X1 U12722 ( .A(n18174), .Z(n18179) );
  NOR2_X1 U12723 ( .A1(n18144), .A2(n18099), .ZN(n18145) );
  OAI21_X1 U12724 ( .B1(n15512), .B2(n21026), .A(n12758), .ZN(n12759) );
  INV_X1 U12725 ( .A(n10143), .ZN(P1_U2838) );
  AOI21_X1 U12726 ( .B1(n21018), .B2(n21017), .A(n10144), .ZN(n10143) );
  NAND2_X1 U12727 ( .A1(n21027), .A2(n21028), .ZN(n10148) );
  NAND2_X1 U12728 ( .A1(n14793), .A2(n21095), .ZN(n14794) );
  NAND2_X1 U12729 ( .A1(n10116), .A2(n10118), .ZN(n15546) );
  INV_X1 U12730 ( .A(n10277), .ZN(n15325) );
  AOI21_X1 U12731 ( .B1(n15507), .B2(n15324), .A(n15323), .ZN(n10278) );
  NAND2_X1 U12732 ( .A1(n9941), .A2(n9940), .ZN(P1_U3000) );
  AND2_X1 U12733 ( .A1(n9800), .A2(n10132), .ZN(n9940) );
  NAND2_X1 U12734 ( .A1(n10133), .A2(n21135), .ZN(n10132) );
  OR2_X1 U12735 ( .A1(n15515), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9987) );
  NAND2_X1 U12736 ( .A1(n10117), .A2(n15545), .ZN(P1_U3004) );
  OR2_X1 U12737 ( .A1(n12966), .A2(n12965), .ZN(n12979) );
  AOI21_X1 U12738 ( .B1(n15999), .B2(n15991), .A(n15998), .ZN(n16003) );
  NAND2_X1 U12739 ( .A1(n15997), .A2(n15996), .ZN(n15998) );
  NOR2_X1 U12740 ( .A1(n16748), .A2(n16750), .ZN(n16751) );
  NAND2_X1 U12741 ( .A1(n16771), .A2(n16852), .ZN(n16777) );
  AOI21_X1 U12742 ( .B1(n17155), .B2(n16881), .A(n16880), .ZN(n16882) );
  NAND2_X1 U12743 ( .A1(n9798), .A2(n10334), .ZN(n17185) );
  NAND2_X1 U12744 ( .A1(n17219), .A2(n9770), .ZN(n16921) );
  AOI21_X1 U12745 ( .B1(n16930), .B2(n20252), .A(n16929), .ZN(n9951) );
  AOI21_X1 U12746 ( .B1(n10355), .B2(n9919), .A(n9968), .ZN(n9967) );
  NAND2_X1 U12747 ( .A1(n9970), .A2(n9969), .ZN(n9968) );
  AOI21_X1 U12748 ( .B1(n14770), .B2(n20252), .A(n13505), .ZN(n13506) );
  OAI211_X1 U12749 ( .C1(n16988), .C2(n20256), .A(n10435), .B(n10434), .ZN(
        P2_U2997) );
  AOI21_X1 U12750 ( .B1(n16987), .B2(n20252), .A(n16986), .ZN(n10434) );
  NAND2_X1 U12751 ( .A1(n9677), .A2(n18070), .ZN(n10435) );
  INV_X1 U12752 ( .A(n10161), .ZN(n16996) );
  AOI21_X1 U12753 ( .B1(n16995), .B2(n20252), .A(n16994), .ZN(n10162) );
  INV_X1 U12754 ( .A(n9932), .ZN(n13044) );
  NAND2_X1 U12755 ( .A1(n9797), .A2(n20267), .ZN(n10413) );
  NAND2_X1 U12756 ( .A1(n17219), .A2(n9769), .ZN(n17220) );
  NAND2_X1 U12757 ( .A1(n9677), .A2(n20279), .ZN(n10065) );
  OAI21_X1 U12758 ( .B1(n17306), .B2(n17297), .A(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n10066) );
  NAND2_X1 U12759 ( .A1(n17324), .A2(n20267), .ZN(n17339) );
  OR2_X1 U12760 ( .A1(n18213), .A2(n18212), .ZN(n10507) );
  NAND2_X1 U12761 ( .A1(n10251), .A2(n10248), .ZN(n17760) );
  NAND2_X1 U12762 ( .A1(n17865), .A2(n19275), .ZN(n10251) );
  AOI21_X1 U12763 ( .B1(n17773), .B2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n13409), .ZN(n13410) );
  INV_X1 U12764 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n19257) );
  INV_X2 U12765 ( .A(n9688), .ZN(n15394) );
  AND3_X1 U12766 ( .A1(n9749), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A3(
        P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n9718) );
  AND3_X1 U12767 ( .A1(n12125), .A2(n12126), .A3(n9824), .ZN(n9719) );
  NOR2_X1 U12768 ( .A1(n13151), .A2(n14838), .ZN(n14825) );
  INV_X1 U12769 ( .A(n15384), .ZN(n10114) );
  AND2_X1 U12770 ( .A1(n9726), .A2(n10449), .ZN(n9720) );
  OR2_X1 U12771 ( .A1(n11085), .A2(n10587), .ZN(n9721) );
  AND4_X1 U12772 ( .A1(n11853), .A2(n11852), .A3(n11851), .A4(n11850), .ZN(
        n9722) );
  INV_X1 U12773 ( .A(n17021), .ZN(n10009) );
  NAND2_X1 U12774 ( .A1(n12873), .A2(n12872), .ZN(n12943) );
  INV_X1 U12775 ( .A(n10771), .ZN(n11385) );
  NAND2_X1 U12776 ( .A1(n14228), .A2(n14227), .ZN(n14285) );
  BUF_X2 U12777 ( .A(n10792), .Z(n14218) );
  INV_X1 U12778 ( .A(n10806), .ZN(n9910) );
  NAND2_X1 U12780 ( .A1(n13146), .A2(n10514), .ZN(n13439) );
  NAND2_X1 U12781 ( .A1(n12125), .A2(n12126), .ZN(n15129) );
  NAND2_X1 U12782 ( .A1(n16140), .A2(n10571), .ZN(n14781) );
  OR2_X1 U12783 ( .A1(n16676), .A2(n16677), .ZN(n16672) );
  NAND2_X1 U12784 ( .A1(n11113), .A2(n10308), .ZN(n9723) );
  NAND2_X1 U12785 ( .A1(n10466), .A2(n9820), .ZN(n9724) );
  NAND2_X2 U12786 ( .A1(n10083), .A2(n10082), .ZN(n11011) );
  NOR2_X1 U12787 ( .A1(n13048), .A2(n16916), .ZN(n16892) );
  INV_X1 U12788 ( .A(n10806), .ZN(n14230) );
  AND2_X1 U12789 ( .A1(n11093), .A2(n11088), .ZN(n9725) );
  INV_X1 U12790 ( .A(n16917), .ZN(n9871) );
  AND2_X1 U12791 ( .A1(n16366), .A2(n16378), .ZN(n9726) );
  NAND2_X1 U12792 ( .A1(n17526), .A2(n11212), .ZN(n11009) );
  INV_X1 U12793 ( .A(n10089), .ZN(n9904) );
  AOI21_X1 U12794 ( .B1(n9688), .B2(n13464), .A(n10545), .ZN(n10544) );
  INV_X1 U12795 ( .A(n10544), .ZN(n10368) );
  AND2_X1 U12796 ( .A1(n13015), .A2(n16927), .ZN(n9727) );
  AND3_X1 U12797 ( .A1(n10855), .A2(n10858), .A3(n10862), .ZN(n9728) );
  AND2_X1 U12798 ( .A1(n9922), .A2(n13068), .ZN(n9729) );
  AND2_X1 U12799 ( .A1(n11510), .A2(n20264), .ZN(n9730) );
  AND2_X1 U12800 ( .A1(n11242), .A2(n11250), .ZN(n9731) );
  OR2_X1 U12801 ( .A1(n10490), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n9732) );
  AND4_X1 U12802 ( .A1(n10944), .A2(n10943), .A3(n10942), .A4(n10941), .ZN(
        n9733) );
  AND2_X1 U12803 ( .A1(n13411), .A2(n15531), .ZN(n9734) );
  NAND2_X1 U12804 ( .A1(n10585), .A2(n10584), .ZN(n9735) );
  NAND2_X1 U12805 ( .A1(n10481), .A2(n11443), .ZN(n16160) );
  NAND2_X1 U12806 ( .A1(n12763), .A2(n9817), .ZN(n16074) );
  AND2_X1 U12807 ( .A1(n9762), .A2(n10496), .ZN(n9736) );
  NAND2_X1 U12808 ( .A1(n20267), .A2(n10354), .ZN(n9737) );
  INV_X1 U12809 ( .A(n18518), .ZN(n10503) );
  INV_X1 U12810 ( .A(n10620), .ZN(n10411) );
  OR2_X1 U12811 ( .A1(n10056), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9738) );
  INV_X2 U12812 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n21349) );
  NAND2_X1 U12813 ( .A1(n14081), .A2(n14083), .ZN(n14082) );
  AND2_X1 U12814 ( .A1(n11526), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9739) );
  NAND2_X1 U12815 ( .A1(n10476), .A2(n11411), .ZN(n14518) );
  AND2_X1 U12816 ( .A1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n9740) );
  AND2_X1 U12817 ( .A1(n10447), .A2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n9741) );
  AND2_X1 U12818 ( .A1(n9740), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n9742) );
  NAND2_X1 U12819 ( .A1(n11869), .A2(n14390), .ZN(n21617) );
  INV_X1 U12820 ( .A(n21617), .ZN(n15959) );
  AND2_X1 U12821 ( .A1(n13010), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n9743) );
  AND2_X1 U12822 ( .A1(n10149), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n9744) );
  OR2_X1 U12823 ( .A1(n10275), .A2(n10273), .ZN(n9745) );
  AND2_X1 U12824 ( .A1(n17086), .A2(n17084), .ZN(n9746) );
  AND2_X1 U12825 ( .A1(n10374), .A2(P3_EAX_REG_27__SCAN_IN), .ZN(n9747) );
  AND2_X1 U12826 ( .A1(n10402), .A2(n9859), .ZN(n9748) );
  AND2_X1 U12827 ( .A1(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n9749) );
  INV_X1 U12828 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n10602) );
  OR2_X1 U12829 ( .A1(n12930), .A2(n12934), .ZN(n9750) );
  CLKBUF_X3 U12830 ( .A(n13273), .Z(n18735) );
  OR3_X1 U12831 ( .A1(n13000), .A2(n11073), .A3(n17239), .ZN(n9751) );
  AND2_X2 U12832 ( .A1(n11741), .A2(n10320), .ZN(n12075) );
  OR2_X1 U12833 ( .A1(n10253), .A2(n19184), .ZN(n9752) );
  AND2_X2 U12834 ( .A1(n9685), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10891) );
  AND4_X1 U12835 ( .A1(n13196), .A2(n13195), .A3(n13194), .A4(n13193), .ZN(
        n9753) );
  OR2_X1 U12836 ( .A1(n16004), .A2(n16005), .ZN(n9754) );
  INV_X1 U12837 ( .A(n10490), .ZN(n17920) );
  NAND2_X1 U12838 ( .A1(n10491), .A2(n17937), .ZN(n10490) );
  AOI22_X1 U12839 ( .A1(n10544), .A2(n15394), .B1(n15394), .B2(n13143), .ZN(
        n10367) );
  NOR2_X1 U12840 ( .A1(n14992), .A2(n14994), .ZN(n14980) );
  NAND2_X1 U12841 ( .A1(n14285), .A2(n9978), .ZN(n16367) );
  NOR2_X1 U12842 ( .A1(n12881), .A2(n10444), .ZN(n12885) );
  OAI21_X2 U12843 ( .B1(n15165), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n12093), 
        .ZN(n14364) );
  NAND2_X1 U12844 ( .A1(n14901), .A2(n14903), .ZN(n14887) );
  AND2_X1 U12845 ( .A1(n16140), .A2(n16142), .ZN(n16125) );
  AND3_X1 U12846 ( .A1(n12125), .A2(n12126), .A3(n10281), .ZN(n15113) );
  NAND2_X1 U12847 ( .A1(n10424), .A2(n16314), .ZN(n17116) );
  INV_X2 U12848 ( .A(n11593), .ZN(n18740) );
  NAND2_X1 U12849 ( .A1(n12763), .A2(n16805), .ZN(n16079) );
  AND2_X1 U12850 ( .A1(n16140), .A2(n10569), .ZN(n9755) );
  AND2_X1 U12851 ( .A1(n10193), .A2(n16907), .ZN(n9756) );
  AND2_X1 U12852 ( .A1(n10186), .A2(n10188), .ZN(n9757) );
  AND3_X1 U12853 ( .A1(n12595), .A2(n12594), .A3(n12627), .ZN(n9758) );
  AND2_X1 U12854 ( .A1(n18818), .A2(n10374), .ZN(n9759) );
  XOR2_X1 U12855 ( .A(n13054), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .Z(
        n9760) );
  AND3_X1 U12856 ( .A1(n10169), .A2(n10167), .A3(n10166), .ZN(n9761) );
  NAND2_X1 U12857 ( .A1(n11086), .A2(n11079), .ZN(n10608) );
  NOR2_X1 U12858 ( .A1(n12877), .A2(n17123), .ZN(n12879) );
  AND2_X1 U12859 ( .A1(n11532), .A2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n9762) );
  AND2_X1 U12860 ( .A1(n10586), .A2(n11103), .ZN(n9763) );
  NOR2_X1 U12861 ( .A1(n14992), .A2(n10275), .ZN(n14930) );
  NOR2_X1 U12862 ( .A1(n16181), .A2(n10482), .ZN(n16151) );
  INV_X1 U12863 ( .A(n10396), .ZN(n10395) );
  NAND2_X1 U12864 ( .A1(n10274), .A2(n10552), .ZN(n14943) );
  AND2_X1 U12865 ( .A1(n11171), .A2(n10734), .ZN(n9764) );
  INV_X1 U12866 ( .A(n11202), .ZN(n11173) );
  BUF_X1 U12867 ( .A(n14218), .Z(n16313) );
  NAND2_X1 U12868 ( .A1(n10609), .A2(n11079), .ZN(n17046) );
  OR2_X1 U12869 ( .A1(n20267), .A2(n20275), .ZN(n9765) );
  INV_X1 U12870 ( .A(n14226), .ZN(n14228) );
  OR3_X1 U12871 ( .A1(n16102), .A2(n10485), .A3(n16103), .ZN(n9766) );
  OR2_X1 U12872 ( .A1(n11115), .A2(n11120), .ZN(n9767) );
  INV_X1 U12873 ( .A(n10723), .ZN(n10724) );
  NAND2_X1 U12874 ( .A1(n10222), .A2(n10218), .ZN(n16972) );
  NAND2_X1 U12875 ( .A1(n10621), .A2(n10622), .ZN(n17078) );
  NAND2_X1 U12876 ( .A1(n10229), .A2(n10381), .ZN(n16989) );
  NAND2_X1 U12877 ( .A1(n10394), .A2(n15492), .ZN(n15484) );
  NOR2_X1 U12878 ( .A1(n12881), .A2(n10441), .ZN(n12888) );
  NOR2_X1 U12879 ( .A1(n17810), .A2(n17811), .ZN(n11533) );
  AND2_X1 U12880 ( .A1(n16885), .A2(n16884), .ZN(n9768) );
  AND2_X1 U12881 ( .A1(n10175), .A2(n20267), .ZN(n9769) );
  AND2_X1 U12882 ( .A1(n10175), .A2(n17155), .ZN(n9770) );
  NAND2_X1 U12883 ( .A1(n17021), .A2(n10012), .ZN(n9771) );
  AND4_X1 U12884 ( .A1(n11773), .A2(n11772), .A3(n11771), .A4(n11770), .ZN(
        n9773) );
  NAND2_X1 U12885 ( .A1(n11089), .A2(n11088), .ZN(n11091) );
  NAND2_X1 U12886 ( .A1(n12927), .A2(n16938), .ZN(n16068) );
  AND2_X1 U12887 ( .A1(n11872), .A2(n11871), .ZN(n11875) );
  OR2_X1 U12888 ( .A1(n16879), .A2(n20196), .ZN(n9774) );
  AND2_X1 U12889 ( .A1(n10159), .A2(n10088), .ZN(n9775) );
  AND2_X1 U12890 ( .A1(n19202), .A2(n19201), .ZN(n9776) );
  AND2_X1 U12891 ( .A1(n10224), .A2(n10223), .ZN(n9777) );
  AND2_X1 U12892 ( .A1(n10344), .A2(n10340), .ZN(n9778) );
  NAND2_X1 U12893 ( .A1(n10745), .A2(n10767), .ZN(n10768) );
  INV_X1 U12894 ( .A(n16895), .ZN(n10039) );
  OR2_X1 U12895 ( .A1(n14992), .A2(n10553), .ZN(n14957) );
  NOR2_X1 U12896 ( .A1(n10458), .A2(n16659), .ZN(n9779) );
  AND2_X1 U12897 ( .A1(n13315), .A2(n13316), .ZN(n9780) );
  INV_X1 U12898 ( .A(n10432), .ZN(n10431) );
  OAI21_X1 U12899 ( .B1(n10607), .B2(n10433), .A(n10636), .ZN(n10432) );
  AND2_X1 U12900 ( .A1(n10362), .A2(n10364), .ZN(n9781) );
  AND2_X1 U12901 ( .A1(n13548), .A2(n19184), .ZN(n17907) );
  NOR2_X1 U12902 ( .A1(n10368), .A2(n10114), .ZN(n10113) );
  AND2_X1 U12903 ( .A1(n14081), .A2(n9920), .ZN(n9782) );
  INV_X1 U12904 ( .A(n10608), .ZN(n10607) );
  AND2_X1 U12905 ( .A1(n17767), .A2(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n9783) );
  NAND2_X1 U12906 ( .A1(n11010), .A2(n11144), .ZN(n11178) );
  AOI21_X1 U12907 ( .B1(n16633), .B2(n20252), .A(n13067), .ZN(n13068) );
  INV_X1 U12908 ( .A(n9925), .ZN(n17176) );
  NAND2_X1 U12909 ( .A1(n9754), .A2(n16006), .ZN(n9925) );
  AND2_X1 U12910 ( .A1(n10542), .A2(n10324), .ZN(n9784) );
  INV_X1 U12911 ( .A(n10384), .ZN(n10383) );
  OR2_X1 U12912 ( .A1(n19030), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n9785) );
  AND2_X1 U12913 ( .A1(n10037), .A2(n10039), .ZN(n9786) );
  AND2_X1 U12914 ( .A1(n9763), .A2(n11104), .ZN(n9787) );
  INV_X1 U12915 ( .A(n14992), .ZN(n10274) );
  INV_X1 U12916 ( .A(n10528), .ZN(n14896) );
  NOR2_X1 U12917 ( .A1(n14954), .A2(n10531), .ZN(n10528) );
  AND2_X1 U12918 ( .A1(n10502), .A2(n19058), .ZN(n9788) );
  NOR2_X1 U12919 ( .A1(n16676), .A2(n10451), .ZN(n16667) );
  AND2_X1 U12920 ( .A1(n10341), .A2(n9760), .ZN(n9789) );
  AND2_X1 U12921 ( .A1(n9890), .A2(n9888), .ZN(n9790) );
  OR2_X1 U12922 ( .A1(n10577), .A2(n14358), .ZN(n9791) );
  INV_X1 U12923 ( .A(n12054), .ZN(n10234) );
  OAI21_X1 U12924 ( .B1(n12606), .B2(n21162), .A(n12003), .ZN(n12054) );
  AND2_X1 U12925 ( .A1(n16960), .A2(n16962), .ZN(n9792) );
  NAND2_X1 U12926 ( .A1(n15326), .A2(n10106), .ZN(n9793) );
  AND2_X1 U12927 ( .A1(n10810), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n9794) );
  INV_X1 U12928 ( .A(n10000), .ZN(n10748) );
  NAND2_X1 U12929 ( .A1(n10003), .A2(n10001), .ZN(n10000) );
  NAND2_X1 U12930 ( .A1(n17012), .A2(n17024), .ZN(n9795) );
  NAND2_X1 U12931 ( .A1(n14901), .A2(n10550), .ZN(n14874) );
  AND2_X1 U12932 ( .A1(n10603), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n9796) );
  AND2_X1 U12933 ( .A1(n13058), .A2(n9923), .ZN(n9797) );
  INV_X1 U12934 ( .A(n10430), .ZN(n10390) );
  INV_X1 U12935 ( .A(n10639), .ZN(n10579) );
  AND2_X1 U12936 ( .A1(n10333), .A2(n10335), .ZN(n9798) );
  INV_X1 U12937 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n18059) );
  AND3_X1 U12938 ( .A1(n10946), .A2(n10945), .A3(n10947), .ZN(n9799) );
  AND3_X1 U12939 ( .A1(n15518), .A2(n15517), .A3(n15516), .ZN(n9800) );
  NAND2_X1 U12940 ( .A1(n10131), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15492) );
  INV_X1 U12941 ( .A(n15492), .ZN(n10397) );
  NAND3_X1 U12942 ( .A1(n11871), .A2(n11870), .A3(n13146), .ZN(n11907) );
  AND2_X1 U12943 ( .A1(n11061), .A2(n11063), .ZN(n9801) );
  AND2_X1 U12944 ( .A1(n10511), .A2(n10510), .ZN(n9802) );
  AND2_X1 U12945 ( .A1(n10308), .A2(n11130), .ZN(n9803) );
  AND2_X1 U12946 ( .A1(n10236), .A2(n11251), .ZN(n9804) );
  NAND2_X1 U12947 ( .A1(n9872), .A2(n10056), .ZN(n10103) );
  XNOR2_X1 U12948 ( .A(n11987), .B(n11986), .ZN(n9806) );
  AND2_X1 U12949 ( .A1(n11393), .A2(n10610), .ZN(n9807) );
  AND2_X1 U12950 ( .A1(n10335), .A2(n20279), .ZN(n9808) );
  AND2_X1 U12951 ( .A1(n9952), .A2(n9951), .ZN(n9809) );
  AND2_X1 U12952 ( .A1(n10495), .A2(n10494), .ZN(n9810) );
  AND2_X1 U12953 ( .A1(n12960), .A2(n10626), .ZN(n9811) );
  INV_X1 U12954 ( .A(n10732), .ZN(n17575) );
  AND2_X1 U12955 ( .A1(n10547), .A2(n12032), .ZN(n9812) );
  OAI21_X1 U12956 ( .B1(n10417), .B2(n10418), .A(n16885), .ZN(n10416) );
  INV_X1 U12957 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14728) );
  AND2_X1 U12958 ( .A1(n10212), .A2(n20279), .ZN(n9813) );
  INV_X2 U12959 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n17650) );
  AND2_X1 U12960 ( .A1(n10721), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9814) );
  INV_X1 U12961 ( .A(n16858), .ZN(n11255) );
  OR2_X1 U12962 ( .A1(n16065), .A2(n10593), .ZN(n10591) );
  BUF_X1 U12963 ( .A(n12019), .Z(n12483) );
  INV_X1 U12964 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n10263) );
  INV_X1 U12965 ( .A(n20277), .ZN(n18091) );
  OR2_X1 U12966 ( .A1(n14385), .A2(n21349), .ZN(n9815) );
  INV_X1 U12967 ( .A(n11906), .ZN(n12622) );
  NAND2_X1 U12968 ( .A1(n9682), .A2(n18787), .ZN(n18886) );
  INV_X1 U12969 ( .A(n14170), .ZN(n14112) );
  NAND2_X1 U12970 ( .A1(n11533), .A2(n10495), .ZN(n11529) );
  AND2_X1 U12971 ( .A1(n14134), .A2(n14133), .ZN(n15286) );
  INV_X2 U12972 ( .A(n15286), .ZN(n14816) );
  NAND2_X1 U12973 ( .A1(n11523), .A2(n20923), .ZN(n17443) );
  INV_X1 U12974 ( .A(n17443), .ZN(n20279) );
  AND2_X1 U12975 ( .A1(n18060), .A2(n20902), .ZN(n20252) );
  INV_X1 U12976 ( .A(n20252), .ZN(n17126) );
  NAND2_X1 U12977 ( .A1(n14274), .A2(n14273), .ZN(n14275) );
  AND2_X1 U12978 ( .A1(n14759), .A2(n11376), .ZN(n16140) );
  OR2_X1 U12979 ( .A1(n14082), .A2(n10579), .ZN(n14116) );
  NAND2_X1 U12980 ( .A1(n16367), .A2(n16366), .ZN(n16694) );
  AND2_X2 U12981 ( .A1(n10077), .A2(n10076), .ZN(n10720) );
  AND2_X1 U12982 ( .A1(n11533), .A2(n9736), .ZN(n9816) );
  NAND2_X1 U12983 ( .A1(n12931), .A2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12930) );
  NAND2_X1 U12984 ( .A1(n9731), .A2(n14352), .ZN(n14561) );
  NAND2_X1 U12985 ( .A1(n10632), .A2(n9740), .ZN(n12910) );
  OR2_X1 U12986 ( .A1(n19201), .A2(n19202), .ZN(n10246) );
  INV_X1 U12987 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n17703) );
  NAND2_X1 U12988 ( .A1(n9974), .A2(n9972), .ZN(n16686) );
  AND2_X1 U12989 ( .A1(n10562), .A2(n16805), .ZN(n9817) );
  NOR2_X1 U12990 ( .A1(n14509), .A2(n10477), .ZN(n16251) );
  NOR2_X1 U12991 ( .A1(n9750), .A2(n16029), .ZN(n12936) );
  NAND2_X1 U12992 ( .A1(n10468), .A2(n11426), .ZN(n13530) );
  NAND2_X1 U12993 ( .A1(n10563), .A2(n11333), .ZN(n14514) );
  NAND2_X1 U12994 ( .A1(n11867), .A2(n13440), .ZN(n13448) );
  NAND2_X1 U12995 ( .A1(n16410), .A2(n16409), .ZN(n16676) );
  OR2_X1 U12996 ( .A1(n16302), .A2(n17436), .ZN(n9818) );
  AND2_X1 U12997 ( .A1(n15037), .A2(n15056), .ZN(n9819) );
  NOR2_X1 U12998 ( .A1(n16626), .A2(n10465), .ZN(n9820) );
  OR2_X1 U12999 ( .A1(n11012), .A2(n11096), .ZN(n9821) );
  NOR3_X1 U13000 ( .A1(n9750), .A2(n10440), .A3(n16029), .ZN(n12938) );
  NAND2_X1 U13001 ( .A1(n10107), .A2(n13116), .ZN(n18017) );
  NOR2_X1 U13002 ( .A1(n14509), .A2(n10474), .ZN(n16238) );
  NOR2_X1 U13003 ( .A1(n13531), .A2(n10471), .ZN(n16202) );
  AND2_X1 U13004 ( .A1(n10632), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12907) );
  INV_X1 U13005 ( .A(n16913), .ZN(n10419) );
  OR3_X1 U13006 ( .A1(n9750), .A2(n10439), .A3(n10440), .ZN(n9822) );
  INV_X1 U13007 ( .A(n11112), .ZN(n10309) );
  AND2_X1 U13008 ( .A1(n16293), .A2(n10327), .ZN(n9823) );
  NAND2_X1 U13009 ( .A1(n11265), .A2(n11264), .ZN(n14081) );
  INV_X1 U13010 ( .A(n21125), .ZN(n21135) );
  AND2_X1 U13011 ( .A1(n10281), .A2(n15114), .ZN(n9824) );
  XOR2_X1 U13012 ( .A(n13111), .B(n13109), .Z(n9825) );
  NAND2_X1 U13013 ( .A1(n9782), .A2(n13527), .ZN(n13526) );
  INV_X1 U13014 ( .A(n9965), .ZN(n9964) );
  OR2_X1 U13015 ( .A1(n10770), .A2(n20909), .ZN(n9826) );
  AND2_X1 U13016 ( .A1(n9746), .A2(n9823), .ZN(n9827) );
  INV_X1 U13017 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n17048) );
  OR2_X1 U13018 ( .A1(n10595), .A2(n11056), .ZN(n9828) );
  NAND2_X1 U13019 ( .A1(n12441), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n9829) );
  INV_X1 U13020 ( .A(n10587), .ZN(n10586) );
  NAND2_X1 U13021 ( .A1(n9725), .A2(n9821), .ZN(n10587) );
  OR2_X1 U13022 ( .A1(n19172), .A2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n9830) );
  AND3_X1 U13023 ( .A1(n15023), .A2(n12261), .A3(n15033), .ZN(n9831) );
  NAND2_X1 U13024 ( .A1(n9964), .A2(n9966), .ZN(n9832) );
  AND2_X1 U13025 ( .A1(n13083), .A2(n10109), .ZN(n9833) );
  AND2_X1 U13026 ( .A1(n9817), .A2(n10561), .ZN(n9834) );
  AND2_X1 U13027 ( .A1(n9742), .A2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n9835) );
  INV_X1 U13028 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n18562) );
  AND2_X1 U13029 ( .A1(n9862), .A2(n20750), .ZN(n9836) );
  AND2_X1 U13030 ( .A1(n10450), .A2(n16668), .ZN(n9837) );
  OR2_X1 U13031 ( .A1(n17296), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n9838) );
  AND2_X1 U13032 ( .A1(n9746), .A2(n9818), .ZN(n9839) );
  INV_X1 U13033 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n12202) );
  AND2_X1 U13034 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n9840) );
  NOR2_X4 U13035 ( .A1(n18994), .A2(n19568), .ZN(n9841) );
  INV_X1 U13036 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n10497) );
  AND2_X1 U13037 ( .A1(n17778), .A2(n10505), .ZN(n9842) );
  INV_X1 U13038 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n10155) );
  NAND2_X1 U13039 ( .A1(n13060), .A2(n20180), .ZN(n20256) );
  NAND3_X1 U13040 ( .A1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A3(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12113) );
  INV_X1 U13041 ( .A(n12113), .ZN(n10141) );
  INV_X1 U13042 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n10150) );
  AND2_X1 U13043 ( .A1(n19494), .A2(P3_REIP_REG_31__SCAN_IN), .ZN(n9843) );
  INV_X1 U13044 ( .A(n16938), .ZN(n10190) );
  AND2_X1 U13045 ( .A1(n19165), .A2(n19400), .ZN(n9844) );
  INV_X1 U13046 ( .A(n14929), .ZN(n10273) );
  INV_X1 U13047 ( .A(n17654), .ZN(n12781) );
  AND2_X1 U13048 ( .A1(n11391), .A2(n11390), .ZN(n9845) );
  INV_X1 U13049 ( .A(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n10138) );
  NAND2_X1 U13050 ( .A1(n10359), .A2(n14459), .ZN(n13433) );
  AND2_X1 U13051 ( .A1(n10492), .A2(n13317), .ZN(n9846) );
  INV_X1 U13052 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11735) );
  INV_X1 U13053 ( .A(n14265), .ZN(n12648) );
  AND2_X1 U13054 ( .A1(n18310), .A2(n10503), .ZN(n9847) );
  AND2_X1 U13055 ( .A1(n9741), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n9848) );
  AND2_X1 U13056 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n21144), .ZN(
        n9849) );
  INV_X1 U13057 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n9937) );
  INV_X1 U13058 ( .A(n11487), .ZN(n17136) );
  NOR2_X1 U13059 ( .A1(n15898), .A2(n21269), .ZN(n9850) );
  NOR2_X1 U13060 ( .A1(n15898), .A2(n21464), .ZN(n9851) );
  INV_X1 U13061 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n10019) );
  INV_X1 U13062 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n10109) );
  AND2_X1 U13063 ( .A1(n19227), .A2(n10511), .ZN(n17848) );
  INV_X1 U13064 ( .A(n20429), .ZN(n10616) );
  AND3_X1 U13065 ( .A1(n19227), .A2(n19146), .A3(n9802), .ZN(n17819) );
  INV_X1 U13066 ( .A(n10403), .ZN(n10296) );
  AND2_X1 U13067 ( .A1(n11521), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10403) );
  OR2_X1 U13068 ( .A1(n10625), .A2(n13036), .ZN(n9852) );
  OR2_X1 U13069 ( .A1(n20650), .A2(n20742), .ZN(n9853) );
  AND2_X1 U13070 ( .A1(n15637), .A2(n21743), .ZN(n9854) );
  NAND2_X1 U13071 ( .A1(n16287), .A2(n17101), .ZN(n16276) );
  INV_X1 U13072 ( .A(n16276), .ZN(n10195) );
  NOR2_X1 U13073 ( .A1(n13144), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n9855) );
  AND2_X1 U13074 ( .A1(n9748), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n9856) );
  INV_X1 U13075 ( .A(n10196), .ZN(n16287) );
  NAND2_X1 U13076 ( .A1(n10198), .A2(n10197), .ZN(n10196) );
  INV_X1 U13077 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n9966) );
  NOR2_X1 U13078 ( .A1(n11486), .A2(n11519), .ZN(n17240) );
  AND2_X1 U13079 ( .A1(n13032), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9857) );
  INV_X1 U13080 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10580) );
  INV_X1 U13081 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n10259) );
  INV_X1 U13082 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n10151) );
  INV_X1 U13083 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n21776) );
  OR2_X1 U13084 ( .A1(n17239), .A2(n13034), .ZN(n9858) );
  INV_X1 U13085 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n10357) );
  AND2_X1 U13086 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n9859) );
  INV_X1 U13087 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n10240) );
  INV_X1 U13088 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n10440) );
  INV_X1 U13089 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n10448) );
  INV_X1 U13090 ( .A(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10142) );
  AND2_X1 U13091 ( .A1(n13030), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n9860) );
  OAI21_X1 U13092 ( .B1(n16959), .B2(n20249), .A(n9967), .ZN(P2_U2993) );
  OAI211_X1 U13093 ( .C1(n14788), .C2(n20249), .A(n10349), .B(n13506), .ZN(
        P2_U2995) );
  OR2_X1 U13094 ( .A1(n13170), .A2(n20249), .ZN(n13171) );
  OR2_X1 U13095 ( .A1(n17230), .A2(n20249), .ZN(n9952) );
  OAI21_X1 U13096 ( .B1(n13477), .B2(n21139), .A(n9984), .ZN(P1_U3001) );
  NOR3_X2 U13097 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20909), .A3(
        n20741), .ZN(n20731) );
  NOR2_X4 U13098 ( .A1(n21623), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n21581) );
  INV_X1 U13099 ( .A(n21625), .ZN(n21623) );
  NOR2_X2 U13101 ( .A1(n16313), .A2(n10821), .ZN(n17520) );
  OR2_X1 U13102 ( .A1(n17520), .A2(n20742), .ZN(n9862) );
  NAND2_X1 U13103 ( .A1(n9886), .A2(n9863), .ZN(n10868) );
  NAND2_X1 U13104 ( .A1(n17520), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n9864) );
  NAND2_X1 U13105 ( .A1(n17520), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n9865) );
  AND2_X1 U13106 ( .A1(n10333), .A2(n9808), .ZN(n10332) );
  NAND2_X2 U13107 ( .A1(n10104), .A2(n10103), .ZN(n10130) );
  INV_X1 U13108 ( .A(n14367), .ZN(n9879) );
  NAND2_X2 U13109 ( .A1(n15385), .A2(n10113), .ZN(n10111) );
  OAI211_X2 U13110 ( .C1(n10107), .C2(n10047), .A(n9881), .B(n9880), .ZN(
        n10363) );
  NAND2_X1 U13111 ( .A1(n10311), .A2(n18018), .ZN(n9880) );
  AOI21_X2 U13112 ( .B1(n10046), .B2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n10397), .ZN(n9881) );
  NAND2_X2 U13113 ( .A1(n18023), .A2(n18024), .ZN(n10107) );
  XNOR2_X2 U13114 ( .A(n13115), .B(n15737), .ZN(n18024) );
  NAND2_X2 U13115 ( .A1(n13114), .A2(n13113), .ZN(n13115) );
  NAND3_X1 U13116 ( .A1(n15500), .A2(n10108), .A3(n9883), .ZN(n9882) );
  NAND2_X1 U13117 ( .A1(n9884), .A2(n21114), .ZN(n9883) );
  INV_X1 U13118 ( .A(n15501), .ZN(n9884) );
  OR2_X1 U13119 ( .A1(n9911), .A2(n9853), .ZN(n17631) );
  NAND2_X1 U13120 ( .A1(n9911), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n9885) );
  NAND2_X1 U13121 ( .A1(n9911), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n9887) );
  AND2_X1 U13122 ( .A1(n9889), .A2(n11171), .ZN(n9888) );
  NAND2_X1 U13123 ( .A1(n10405), .A2(n10732), .ZN(n9889) );
  NAND2_X2 U13124 ( .A1(n10409), .A2(n10408), .ZN(n13031) );
  NAND2_X2 U13125 ( .A1(n9893), .A2(n10236), .ZN(n11511) );
  NAND3_X1 U13126 ( .A1(n10236), .A2(n9893), .A3(n11251), .ZN(n9929) );
  AND2_X1 U13127 ( .A1(n9687), .A2(n9893), .ZN(n10183) );
  NAND2_X1 U13128 ( .A1(n9804), .A2(n9893), .ZN(n10063) );
  INV_X2 U13129 ( .A(n10614), .ZN(n9893) );
  INV_X1 U13130 ( .A(n9894), .ZN(n9907) );
  NAND3_X1 U13131 ( .A1(n10805), .A2(n10801), .A3(
        P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n9896) );
  NAND2_X1 U13132 ( .A1(n9899), .A2(n9900), .ZN(n9898) );
  NAND3_X1 U13133 ( .A1(n14079), .A2(n9775), .A3(
        P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n9899) );
  NOR2_X1 U13134 ( .A1(n20281), .A2(n10089), .ZN(n9903) );
  NOR2_X1 U13135 ( .A1(n20281), .A2(n21655), .ZN(n9905) );
  NAND3_X1 U13136 ( .A1(n10806), .A2(n10807), .A3(
        P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n9913) );
  NAND3_X1 U13137 ( .A1(n10806), .A2(n10807), .A3(
        P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n9915) );
  NAND2_X1 U13138 ( .A1(n20504), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n9912) );
  OAI21_X1 U13139 ( .B1(n20385), .B2(n10866), .A(n9915), .ZN(n10867) );
  NAND2_X1 U13140 ( .A1(n20504), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n9916) );
  OAI21_X1 U13141 ( .B1(n20504), .B2(n20742), .A(n20750), .ZN(n9917) );
  NAND2_X1 U13142 ( .A1(n9918), .A2(n10731), .ZN(n9931) );
  NAND2_X1 U13143 ( .A1(n17984), .A2(n9918), .ZN(n17449) );
  NAND2_X2 U13144 ( .A1(n9686), .A2(n10604), .ZN(n10325) );
  AND2_X2 U13145 ( .A1(n16033), .A2(n16035), .ZN(n16018) );
  AND2_X2 U13146 ( .A1(n16048), .A2(n16051), .ZN(n16033) );
  NAND2_X2 U13147 ( .A1(n14350), .A2(n14349), .ZN(n14352) );
  NAND3_X1 U13148 ( .A1(n9923), .A2(n13058), .A3(n17155), .ZN(n9922) );
  INV_X1 U13149 ( .A(n10175), .ZN(n9924) );
  NAND2_X1 U13150 ( .A1(n9926), .A2(n10620), .ZN(n9928) );
  NAND2_X1 U13151 ( .A1(n9926), .A2(n10623), .ZN(n10621) );
  NAND2_X1 U13152 ( .A1(n10295), .A2(n9926), .ZN(n10294) );
  OAI21_X1 U13153 ( .B1(n9926), .B2(n10293), .A(n10291), .ZN(n16997) );
  OAI21_X1 U13154 ( .B1(n10293), .B2(n9926), .A(n10407), .ZN(n13027) );
  XNOR2_X1 U13155 ( .A(n9926), .B(n18057), .ZN(n18084) );
  AOI21_X1 U13156 ( .B1(n16881), .B2(n20267), .A(n13492), .ZN(n13493) );
  AND2_X2 U13157 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10265) );
  AND2_X2 U13158 ( .A1(n17021), .A2(n9748), .ZN(n16976) );
  NAND2_X4 U13159 ( .A1(n9928), .A2(n10619), .ZN(n17021) );
  NAND3_X1 U13160 ( .A1(n10072), .A2(n17155), .A3(n10073), .ZN(n16941) );
  OAI21_X1 U13161 ( .B1(n13166), .B2(n20290), .A(n9933), .ZN(n9932) );
  XNOR2_X2 U13162 ( .A(n11962), .B(n11961), .ZN(n15165) );
  NAND2_X2 U13163 ( .A1(n9938), .A2(n11887), .ZN(n11962) );
  NOR2_X2 U13164 ( .A1(n15415), .A2(n15414), .ZN(n15404) );
  NAND2_X2 U13165 ( .A1(n14362), .A2(n10537), .ZN(n12103) );
  NAND3_X1 U13166 ( .A1(n14362), .A2(n10537), .A3(n9812), .ZN(n13069) );
  NAND2_X2 U13167 ( .A1(n10538), .A2(n11943), .ZN(n14362) );
  NAND2_X2 U13168 ( .A1(n9942), .A2(n10753), .ZN(n17498) );
  AND2_X1 U13169 ( .A1(n9944), .A2(n17654), .ZN(n17661) );
  AND2_X1 U13170 ( .A1(n9944), .A2(n12781), .ZN(n17655) );
  NAND2_X1 U13171 ( .A1(n9944), .A2(n17984), .ZN(n9943) );
  NAND3_X1 U13172 ( .A1(n9948), .A2(n18056), .A3(n9961), .ZN(n9947) );
  XNOR2_X2 U13173 ( .A(n11517), .B(n13049), .ZN(n18056) );
  XNOR2_X1 U13174 ( .A(n16926), .B(n16928), .ZN(n17230) );
  NAND2_X2 U13175 ( .A1(n9957), .A2(n9956), .ZN(n10734) );
  NAND2_X1 U13176 ( .A1(n10178), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9956) );
  NAND2_X1 U13177 ( .A1(n10177), .A2(n17650), .ZN(n9957) );
  NAND2_X1 U13178 ( .A1(n10165), .A2(n17650), .ZN(n9958) );
  NAND2_X1 U13179 ( .A1(n10164), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9959) );
  NAND2_X1 U13180 ( .A1(n18056), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10622) );
  NOR2_X1 U13181 ( .A1(n13049), .A2(n9966), .ZN(n9965) );
  NAND2_X1 U13182 ( .A1(n10740), .A2(n9971), .ZN(n11167) );
  NAND4_X1 U13183 ( .A1(n9971), .A2(n10733), .A3(n11170), .A4(n10732), .ZN(
        n10730) );
  AND2_X1 U13184 ( .A1(n9971), .A2(n10720), .ZN(n10735) );
  NAND3_X1 U13185 ( .A1(n14228), .A2(n9720), .A3(n14227), .ZN(n9974) );
  NAND2_X1 U13186 ( .A1(n14225), .A2(n14224), .ZN(n14284) );
  AOI21_X1 U13187 ( .B1(n15513), .B2(n9987), .A(n9985), .ZN(n9984) );
  NAND2_X1 U13188 ( .A1(n16637), .A2(n16636), .ZN(n9988) );
  OAI22_X2 U13189 ( .A1(n16661), .A2(n10455), .B1(n10453), .B2(n16669), .ZN(
        n16653) );
  XNOR2_X2 U13190 ( .A(n16669), .B(n16503), .ZN(n16661) );
  INV_X1 U13191 ( .A(n10750), .ZN(n10070) );
  NAND2_X1 U13192 ( .A1(n9994), .A2(n11073), .ZN(n10424) );
  INV_X1 U13193 ( .A(n17140), .ZN(n9992) );
  INV_X1 U13194 ( .A(n9994), .ZN(n9993) );
  OAI21_X1 U13195 ( .B1(n9994), .B2(n10427), .A(n10425), .ZN(n11054) );
  OAI21_X1 U13196 ( .B1(n9994), .B2(n10348), .A(n10346), .ZN(n10062) );
  XNOR2_X2 U13197 ( .A(n10236), .B(n10614), .ZN(n9994) );
  NAND3_X1 U13198 ( .A1(n10268), .A2(n11515), .A3(n10266), .ZN(n17096) );
  NAND3_X1 U13199 ( .A1(n10745), .A2(n10767), .A3(n10002), .ZN(n9999) );
  AND2_X2 U13200 ( .A1(n10315), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10771) );
  NAND2_X1 U13201 ( .A1(n10315), .A2(n9840), .ZN(n10001) );
  INV_X1 U13202 ( .A(n10746), .ZN(n10002) );
  AOI21_X1 U13203 ( .B1(n10773), .B2(P2_EBX_REG_2__SCAN_IN), .A(n10004), .ZN(
        n10003) );
  OAI21_X1 U13204 ( .B1(n10726), .B2(n20830), .A(n10725), .ZN(n10004) );
  NAND3_X1 U13205 ( .A1(n10203), .A2(n10204), .A3(n10011), .ZN(n10328) );
  NAND3_X1 U13206 ( .A1(n10011), .A2(n10204), .A3(n10414), .ZN(n11513) );
  NAND2_X1 U13207 ( .A1(n13305), .A2(n10013), .ZN(n19211) );
  NAND2_X1 U13208 ( .A1(n13304), .A2(n13303), .ZN(n10013) );
  OAI211_X2 U13209 ( .C1(n19248), .C2(n10015), .A(n19234), .B(n10014), .ZN(
        n19233) );
  NAND2_X2 U13210 ( .A1(n19259), .A2(n13289), .ZN(n13294) );
  AND2_X4 U13211 ( .A1(n19423), .A2(n19336), .ZN(n19325) );
  AND2_X4 U13212 ( .A1(n13318), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n19423) );
  INV_X1 U13213 ( .A(n17763), .ZN(n17743) );
  INV_X1 U13214 ( .A(n17907), .ZN(n10023) );
  NOR2_X1 U13215 ( .A1(n17937), .A2(n10024), .ZN(n10025) );
  AND2_X2 U13216 ( .A1(n18998), .A2(n10025), .ZN(n13548) );
  NAND2_X2 U13217 ( .A1(n18999), .A2(n19289), .ZN(n18998) );
  NOR2_X2 U13218 ( .A1(n13327), .A2(n19017), .ZN(n18999) );
  NAND2_X1 U13219 ( .A1(n17121), .A2(n10062), .ZN(n10028) );
  NAND2_X1 U13220 ( .A1(n10267), .A2(n17107), .ZN(n10617) );
  OAI21_X1 U13221 ( .B1(n17185), .B2(n20249), .A(n9729), .ZN(P2_U2986) );
  NAND3_X1 U13222 ( .A1(n11060), .A2(n9839), .A3(n10092), .ZN(n10029) );
  AND2_X4 U13223 ( .A1(n10864), .A2(n10863), .ZN(n10236) );
  NAND3_X1 U13224 ( .A1(n10031), .A2(n10033), .A3(n10030), .ZN(n17197) );
  NAND4_X1 U13225 ( .A1(n10031), .A2(n10033), .A3(n10030), .A4(n18070), .ZN(
        n10038) );
  NAND2_X1 U13226 ( .A1(n16902), .A2(n10038), .ZN(P2_U2987) );
  AND2_X2 U13227 ( .A1(n13031), .A2(n9860), .ZN(n16905) );
  NAND2_X1 U13228 ( .A1(n10043), .A2(n10109), .ZN(n10042) );
  NAND3_X1 U13229 ( .A1(n10122), .A2(n10115), .A3(n10048), .ZN(n10118) );
  AND2_X1 U13230 ( .A1(n10124), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n10048) );
  INV_X1 U13231 ( .A(n15404), .ZN(n10049) );
  NAND3_X1 U13232 ( .A1(n10103), .A2(n10543), .A3(n10104), .ZN(n10051) );
  NAND2_X2 U13233 ( .A1(n10130), .A2(n15404), .ZN(n15385) );
  NAND2_X1 U13234 ( .A1(n10110), .A2(n13083), .ZN(n21090) );
  NAND3_X1 U13235 ( .A1(n10130), .A2(n10057), .A3(n10367), .ZN(n10054) );
  NAND3_X1 U13236 ( .A1(n17298), .A2(n10066), .A3(n10065), .ZN(P2_U3029) );
  AND3_X2 U13237 ( .A1(n10069), .A2(n10429), .A3(n11471), .ZN(n11209) );
  NAND2_X1 U13238 ( .A1(n12783), .A2(n10071), .ZN(n10753) );
  NAND3_X1 U13239 ( .A1(n10072), .A2(n20267), .A3(n10073), .ZN(n17247) );
  AND2_X4 U13240 ( .A1(n10075), .A2(n10074), .ZN(n10731) );
  NAND2_X1 U13241 ( .A1(n10663), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10076) );
  NAND2_X1 U13242 ( .A1(n10658), .A2(n17650), .ZN(n10077) );
  NOR2_X1 U13243 ( .A1(n16976), .A2(n10078), .ZN(n17282) );
  AOI21_X1 U13244 ( .B1(n17021), .B2(n10079), .A(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n10078) );
  NAND2_X1 U13245 ( .A1(n10171), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10081) );
  NAND2_X1 U13246 ( .A1(n10172), .A2(n17650), .ZN(n10080) );
  NAND2_X2 U13247 ( .A1(n10081), .A2(n10080), .ZN(n10733) );
  NAND2_X1 U13248 ( .A1(n10085), .A2(n17650), .ZN(n10084) );
  NAND4_X1 U13249 ( .A1(n10697), .A2(n10698), .A3(n10699), .A4(n10700), .ZN(
        n10085) );
  NAND4_X1 U13250 ( .A1(n10703), .A2(n10704), .A3(n10701), .A4(n10702), .ZN(
        n10087) );
  INV_X1 U13251 ( .A(n10794), .ZN(n10088) );
  NAND2_X1 U13252 ( .A1(n10091), .A2(n10794), .ZN(n10089) );
  INV_X1 U13253 ( .A(n10783), .ZN(n10090) );
  AOI21_X1 U13254 ( .B1(n16926), .B2(n10095), .A(n10416), .ZN(n10094) );
  NAND2_X1 U13255 ( .A1(n10097), .A2(n10098), .ZN(n10096) );
  NAND2_X1 U13256 ( .A1(n14304), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n14303) );
  AOI22_X1 U13257 ( .A1(n14304), .A2(n10100), .B1(n13096), .B2(n9849), .ZN(
        n10099) );
  NAND2_X1 U13258 ( .A1(n14303), .A2(n13096), .ZN(n13105) );
  NAND2_X1 U13259 ( .A1(n10102), .A2(n21131), .ZN(n10101) );
  INV_X1 U13260 ( .A(n13096), .ZN(n10102) );
  OAI21_X1 U13261 ( .B1(n18023), .B2(n18024), .A(n10107), .ZN(n18025) );
  NAND2_X1 U13262 ( .A1(n10110), .A2(n9833), .ZN(n10108) );
  XNOR2_X2 U13263 ( .A(n12103), .B(n12054), .ZN(n13080) );
  NAND3_X2 U13264 ( .A1(n10112), .A2(n10111), .A3(n9855), .ZN(n15317) );
  NAND4_X1 U13265 ( .A1(n10118), .A2(n21110), .A3(n10120), .A4(n10119), .ZN(
        n10117) );
  AND2_X1 U13266 ( .A1(n10120), .A2(n10119), .ZN(n10116) );
  NAND2_X1 U13267 ( .A1(n9793), .A2(n9688), .ZN(n10124) );
  NAND2_X1 U13268 ( .A1(n10121), .A2(n15308), .ZN(n10120) );
  INV_X1 U13269 ( .A(n10330), .ZN(n10420) );
  NAND2_X1 U13270 ( .A1(n9953), .A2(n11006), .ZN(n11010) );
  NOR2_X1 U13271 ( .A1(n10127), .A2(n10126), .ZN(n10125) );
  INV_X1 U13272 ( .A(n10856), .ZN(n10126) );
  INV_X1 U13273 ( .A(n10857), .ZN(n10127) );
  NAND2_X1 U13274 ( .A1(n13134), .A2(n13133), .ZN(n10131) );
  NAND3_X1 U13275 ( .A1(n10136), .A2(n10140), .A3(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n12152) );
  NAND4_X1 U13276 ( .A1(n10140), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A3(
        n10137), .A4(n10141), .ZN(n12157) );
  NAND3_X1 U13277 ( .A1(n21025), .A2(n10148), .A3(n10145), .ZN(n10144) );
  INV_X1 U13278 ( .A(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n10156) );
  NOR2_X2 U13279 ( .A1(n14812), .A2(n12859), .ZN(n20982) );
  CLKBUF_X1 U13280 ( .A(n18085), .Z(n10158) );
  NAND2_X1 U13281 ( .A1(n10158), .A2(n11510), .ZN(n17120) );
  NAND2_X2 U13282 ( .A1(n10795), .A2(n10160), .ZN(n17467) );
  NAND4_X1 U13283 ( .A1(n10670), .A2(n10671), .A3(n10669), .A4(n10668), .ZN(
        n10164) );
  NAND4_X1 U13284 ( .A1(n10666), .A2(n10667), .A3(n10665), .A4(n10664), .ZN(
        n10165) );
  NAND3_X1 U13285 ( .A1(n10169), .A2(n10170), .A3(n10166), .ZN(n14769) );
  NAND4_X1 U13286 ( .A1(n10687), .A2(n10686), .A3(n10685), .A4(n10684), .ZN(
        n10171) );
  NAND4_X1 U13287 ( .A1(n10680), .A2(n10683), .A3(n10682), .A4(n10681), .ZN(
        n10172) );
  NAND2_X2 U13288 ( .A1(n10173), .A2(n20281), .ZN(n20740) );
  AND2_X2 U13289 ( .A1(n10806), .A2(n9775), .ZN(n10173) );
  AND2_X1 U13290 ( .A1(n9857), .A2(n13030), .ZN(n10174) );
  NAND4_X1 U13291 ( .A1(n10672), .A2(n10675), .A3(n10673), .A4(n10674), .ZN(
        n10177) );
  NAND4_X1 U13292 ( .A1(n10678), .A2(n10679), .A3(n10676), .A4(n10677), .ZN(
        n10178) );
  NAND3_X1 U13293 ( .A1(n10179), .A2(n11479), .A3(n10180), .ZN(n10739) );
  NAND3_X1 U13294 ( .A1(n10181), .A2(n17526), .A3(n11202), .ZN(n10179) );
  NAND2_X1 U13295 ( .A1(n11187), .A2(n10729), .ZN(n10181) );
  NAND3_X1 U13296 ( .A1(n10738), .A2(n17667), .A3(n10750), .ZN(n11479) );
  NAND2_X1 U13297 ( .A1(n10727), .A2(n10728), .ZN(n11187) );
  XNOR2_X1 U13298 ( .A(n13069), .B(n12047), .ZN(n13126) );
  NAND2_X1 U13299 ( .A1(n11859), .A2(n14385), .ZN(n11876) );
  OAI21_X1 U13300 ( .B1(n15493), .B2(n10397), .A(n13138), .ZN(n10396) );
  NOR2_X1 U13301 ( .A1(n10535), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n10534) );
  NAND2_X1 U13302 ( .A1(n10786), .A2(n10761), .ZN(n10318) );
  NOR2_X2 U13303 ( .A1(n13474), .A2(n15656), .ZN(n15627) );
  OAI21_X2 U13304 ( .B1(n15554), .B2(n15530), .A(n15528), .ZN(n15521) );
  NAND2_X1 U13305 ( .A1(n10371), .A2(n10370), .ZN(n10369) );
  NAND2_X1 U13306 ( .A1(n10185), .A2(n10187), .ZN(n12933) );
  NAND2_X1 U13307 ( .A1(n12927), .A2(n10188), .ZN(n10185) );
  NAND2_X1 U13308 ( .A1(n10193), .A2(n10191), .ZN(n16007) );
  NAND4_X1 U13309 ( .A1(n10690), .A2(n10688), .A3(n10689), .A4(n10691), .ZN(
        n10201) );
  NAND4_X1 U13310 ( .A1(n10694), .A2(n10695), .A3(n10692), .A4(n10693), .ZN(
        n10202) );
  NAND2_X1 U13311 ( .A1(n10328), .A2(n16293), .ZN(n17080) );
  NAND2_X1 U13312 ( .A1(n11525), .A2(n10205), .ZN(P2_U3025) );
  NAND3_X1 U13313 ( .A1(n10209), .A2(n9813), .A3(n10208), .ZN(n10205) );
  NAND2_X1 U13314 ( .A1(n10391), .A2(n10210), .ZN(n10208) );
  INV_X1 U13315 ( .A(n10391), .ZN(n10207) );
  NAND3_X1 U13316 ( .A1(n10209), .A2(n10212), .A3(n10208), .ZN(n16959) );
  NAND2_X1 U13317 ( .A1(n10226), .A2(n10223), .ZN(n10220) );
  OAI211_X1 U13318 ( .C1(n12103), .C2(n10232), .A(n10230), .B(n10231), .ZN(
        n13107) );
  NAND2_X1 U13319 ( .A1(n13107), .A2(n13127), .ZN(n13114) );
  INV_X1 U13320 ( .A(n12112), .ZN(n10233) );
  NAND2_X1 U13321 ( .A1(n10534), .A2(n10370), .ZN(n10235) );
  NAND2_X1 U13322 ( .A1(n10318), .A2(n10785), .ZN(n10784) );
  INV_X1 U13323 ( .A(n17107), .ZN(n10237) );
  NAND2_X1 U13324 ( .A1(n17380), .A2(n20267), .ZN(n17391) );
  NAND3_X1 U13325 ( .A1(n13277), .A2(n13275), .A3(n13276), .ZN(n10244) );
  INV_X2 U13326 ( .A(n11594), .ZN(n13185) );
  AND2_X2 U13327 ( .A1(n10252), .A2(n14728), .ZN(n14719) );
  AOI21_X1 U13328 ( .B1(n10246), .B2(n10245), .A(n9776), .ZN(n10247) );
  INV_X1 U13329 ( .A(n13387), .ZN(n13385) );
  NAND2_X2 U13330 ( .A1(n19426), .A2(n19336), .ZN(n19385) );
  NAND2_X1 U13331 ( .A1(n10252), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n13333) );
  NAND4_X1 U13332 ( .A1(n21766), .A2(n21883), .A3(n10252), .A4(
        P2_EAX_REG_5__SCAN_IN), .ZN(n21658) );
  NAND2_X1 U13333 ( .A1(n20037), .A2(n10252), .ZN(n14718) );
  NAND2_X1 U13334 ( .A1(n14736), .A2(n10252), .ZN(n14319) );
  MUX2_X1 U13335 ( .A(n19314), .B(n14722), .S(n10252), .Z(n20001) );
  NAND2_X1 U13336 ( .A1(n19185), .A2(n10253), .ZN(n19475) );
  XNOR2_X2 U13337 ( .A(n13294), .B(n13293), .ZN(n19248) );
  NAND2_X1 U13338 ( .A1(n19226), .A2(n10258), .ZN(n10257) );
  XNOR2_X2 U13339 ( .A(n13304), .B(n13302), .ZN(n19226) );
  XNOR2_X2 U13340 ( .A(n13314), .B(n13312), .ZN(n19205) );
  INV_X1 U13341 ( .A(n10265), .ZN(n17479) );
  NAND3_X1 U13342 ( .A1(n10267), .A2(n11513), .A3(n17107), .ZN(n10266) );
  INV_X1 U13343 ( .A(n10345), .ZN(n11166) );
  NAND3_X1 U13344 ( .A1(n12125), .A2(n12126), .A3(n10280), .ZN(n15007) );
  NAND2_X1 U13345 ( .A1(n10282), .A2(n10757), .ZN(n10786) );
  NAND3_X1 U13346 ( .A1(n10767), .A2(n10316), .A3(n10745), .ZN(n10282) );
  NAND2_X1 U13347 ( .A1(n10806), .A2(n10283), .ZN(n10284) );
  OAI21_X1 U13348 ( .B1(n20436), .B2(n10872), .A(n10284), .ZN(n10873) );
  NAND2_X1 U13349 ( .A1(n17616), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n10286) );
  NAND2_X1 U13350 ( .A1(n10288), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n10287) );
  NAND2_X1 U13351 ( .A1(n17616), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n10289) );
  NOR2_X1 U13352 ( .A1(n17616), .A2(n20742), .ZN(n10290) );
  NAND2_X1 U13353 ( .A1(n10294), .A2(n10292), .ZN(n17301) );
  AND2_X4 U13354 ( .A1(n10834), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10833) );
  AND2_X1 U13355 ( .A1(n10833), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n16610) );
  AND2_X2 U13356 ( .A1(n10903), .A2(n10902), .ZN(n10614) );
  NAND2_X1 U13357 ( .A1(n10297), .A2(n17348), .ZN(n17023) );
  NAND2_X1 U13358 ( .A1(n11024), .A2(n10301), .ZN(n11066) );
  NAND2_X1 U13359 ( .A1(n9801), .A2(n11023), .ZN(n10595) );
  CLKBUF_X1 U13360 ( .A(n10833), .Z(n10302) );
  NOR2_X2 U13361 ( .A1(n16043), .A2(n10303), .ZN(n13048) );
  INV_X1 U13362 ( .A(n12995), .ZN(n10304) );
  NAND2_X1 U13363 ( .A1(n11113), .A2(n9803), .ZN(n12987) );
  AND2_X2 U13364 ( .A1(n11735), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10320) );
  NAND2_X2 U13365 ( .A1(n10321), .A2(n11873), .ZN(n13148) );
  NAND2_X1 U13366 ( .A1(n14364), .A2(n10321), .ZN(n12094) );
  XNOR2_X2 U13367 ( .A(n10557), .B(n10323), .ZN(n14363) );
  NOR2_X2 U13368 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10834) );
  NAND2_X1 U13369 ( .A1(n11059), .A2(n11060), .ZN(n17081) );
  INV_X1 U13370 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n10327) );
  NAND2_X1 U13371 ( .A1(n10413), .A2(n10331), .ZN(P2_U3018) );
  AOI21_X1 U13372 ( .B1(n10332), .B2(n10334), .A(n9805), .ZN(n10331) );
  INV_X1 U13373 ( .A(n11510), .ZN(n10348) );
  OR2_X1 U13374 ( .A1(n14769), .A2(n20256), .ZN(n10349) );
  INV_X1 U13375 ( .A(n10726), .ZN(n10772) );
  AOI21_X2 U13376 ( .B1(n13058), .B2(n17162), .A(n16886), .ZN(n17172) );
  NAND2_X1 U13377 ( .A1(n13147), .A2(n11877), .ZN(n13424) );
  NAND2_X1 U13378 ( .A1(n15475), .A2(n10635), .ZN(n15392) );
  INV_X1 U13379 ( .A(n10363), .ZN(n10361) );
  NAND2_X1 U13380 ( .A1(n13079), .A2(n13078), .ZN(n15393) );
  NAND2_X1 U13381 ( .A1(n11989), .A2(n14367), .ZN(n10366) );
  NAND2_X2 U13382 ( .A1(n11945), .A2(n11918), .ZN(n14367) );
  AND2_X1 U13383 ( .A1(n10372), .A2(n17706), .ZN(n11678) );
  NAND2_X1 U13384 ( .A1(n10372), .A2(n20150), .ZN(n13344) );
  NAND2_X1 U13385 ( .A1(n19580), .A2(n10372), .ZN(n13339) );
  INV_X2 U13387 ( .A(n14594), .ZN(n14679) );
  AND2_X2 U13388 ( .A1(n14338), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11554) );
  AND3_X2 U13389 ( .A1(n10377), .A2(n10376), .A3(n10375), .ZN(n13981) );
  OR2_X2 U13390 ( .A1(n11691), .A2(n19565), .ZN(n10377) );
  NAND3_X1 U13391 ( .A1(n10379), .A2(P3_EAX_REG_22__SCAN_IN), .A3(
        P3_EAX_REG_21__SCAN_IN), .ZN(n10378) );
  XNOR2_X2 U13392 ( .A(n10380), .B(n10778), .ZN(n10792) );
  NAND2_X1 U13393 ( .A1(n16972), .A2(n16973), .ZN(n13496) );
  NAND2_X1 U13394 ( .A1(n16972), .A2(n10392), .ZN(n10391) );
  NAND2_X1 U13395 ( .A1(n13125), .A2(n13124), .ZN(n15494) );
  NAND2_X1 U13396 ( .A1(n10401), .A2(n9807), .ZN(n14290) );
  AND2_X2 U13397 ( .A1(n10404), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n17469) );
  NAND2_X1 U13398 ( .A1(n11227), .A2(n17575), .ZN(n11171) );
  NAND2_X2 U13399 ( .A1(n12786), .A2(n11011), .ZN(n11227) );
  INV_X1 U13400 ( .A(n11167), .ZN(n10405) );
  AOI21_X1 U13401 ( .B1(n10411), .B2(n10619), .A(n17238), .ZN(n10407) );
  NAND2_X1 U13402 ( .A1(n10293), .A2(n17240), .ZN(n10408) );
  NAND2_X1 U13403 ( .A1(n11511), .A2(n11516), .ZN(n10414) );
  INV_X1 U13404 ( .A(n13015), .ZN(n10417) );
  NOR2_X1 U13405 ( .A1(n13002), .A2(n10420), .ZN(n16912) );
  NOR2_X2 U13406 ( .A1(n13016), .A2(n10419), .ZN(n10418) );
  NAND2_X1 U13407 ( .A1(n17057), .A2(n10640), .ZN(n10609) );
  NAND2_X1 U13408 ( .A1(n10741), .A2(n10717), .ZN(n10428) );
  NAND2_X1 U13409 ( .A1(n17033), .A2(n12980), .ZN(n17009) );
  NAND3_X1 U13410 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A3(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12877) );
  NAND2_X1 U13411 ( .A1(n16336), .A2(n10445), .ZN(n12923) );
  NAND2_X1 U13412 ( .A1(n16367), .A2(n9726), .ZN(n16690) );
  NOR2_X2 U13413 ( .A1(n16653), .A2(n16504), .ZN(n16542) );
  INV_X1 U13414 ( .A(n16569), .ZN(n10459) );
  AOI21_X1 U13415 ( .B1(n10459), .B2(n9820), .A(n10460), .ZN(n10463) );
  NAND2_X1 U13416 ( .A1(n10467), .A2(n16569), .ZN(n10466) );
  INV_X1 U13417 ( .A(n13531), .ZN(n10468) );
  NAND2_X1 U13418 ( .A1(n10468), .A2(n10469), .ZN(n16191) );
  AND2_X2 U13419 ( .A1(n10473), .A2(n10580), .ZN(n10696) );
  NAND3_X1 U13420 ( .A1(n10488), .A2(n9811), .A3(n10487), .ZN(P2_U2824) );
  NAND2_X1 U13421 ( .A1(n12966), .A2(n16322), .ZN(n10488) );
  NAND2_X1 U13422 ( .A1(n14719), .A2(n11559), .ZN(n11593) );
  INV_X1 U13423 ( .A(n18312), .ZN(n10500) );
  NAND2_X1 U13424 ( .A1(n17778), .A2(n10504), .ZN(n11535) );
  INV_X1 U13425 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n10506) );
  AOI21_X1 U13426 ( .B1(n10508), .B2(n20050), .A(n10507), .ZN(n18216) );
  XNOR2_X1 U13427 ( .A(n18210), .B(n10509), .ZN(n10508) );
  NOR2_X1 U13428 ( .A1(n18217), .A2(n18518), .ZN(n18210) );
  NAND2_X1 U13429 ( .A1(n10513), .A2(n12649), .ZN(n12645) );
  XNOR2_X1 U13430 ( .A(n10513), .B(n14100), .ZN(n15159) );
  XNOR2_X1 U13431 ( .A(n12643), .B(n14144), .ZN(n10513) );
  INV_X2 U13432 ( .A(n11890), .ZN(n12726) );
  INV_X2 U13433 ( .A(n14390), .ZN(n10514) );
  NAND2_X1 U13434 ( .A1(n10516), .A2(n10515), .ZN(P1_U2810) );
  OR2_X1 U13435 ( .A1(n14807), .A2(n21026), .ZN(n10516) );
  XNOR2_X1 U13436 ( .A(n12857), .B(n12856), .ZN(n14807) );
  INV_X1 U13437 ( .A(n14954), .ZN(n10527) );
  NAND3_X1 U13438 ( .A1(n10527), .A2(n10526), .A3(n10529), .ZN(n14862) );
  NAND2_X2 U13439 ( .A1(n12103), .A2(n10536), .ZN(n14524) );
  INV_X1 U13440 ( .A(n10539), .ZN(n11913) );
  NAND2_X1 U13441 ( .A1(n11944), .A2(n10539), .ZN(n21174) );
  OAI21_X1 U13442 ( .B1(n10637), .B2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n15394), .ZN(n10540) );
  NAND2_X1 U13443 ( .A1(n15393), .A2(n15658), .ZN(n10542) );
  INV_X1 U13444 ( .A(n13074), .ZN(n10546) );
  NAND4_X1 U13445 ( .A1(n10546), .A2(n13076), .A3(n13072), .A4(n13075), .ZN(
        n15403) );
  OR2_X2 U13446 ( .A1(n9688), .A2(n15683), .ZN(n13076) );
  NAND3_X1 U13447 ( .A1(n13069), .A2(n13127), .A3(n13117), .ZN(n13123) );
  AND2_X2 U13448 ( .A1(n14901), .A2(n10548), .ZN(n14864) );
  INV_X1 U13449 ( .A(n15007), .ZN(n12281) );
  NAND2_X1 U13450 ( .A1(n21174), .A2(n11945), .ZN(n13944) );
  NAND3_X1 U13451 ( .A1(n21174), .A2(n11945), .A3(n9937), .ZN(n10556) );
  INV_X1 U13452 ( .A(n12069), .ZN(n10557) );
  NAND2_X1 U13453 ( .A1(n13150), .A2(n13152), .ZN(n13151) );
  INV_X1 U13454 ( .A(n13526), .ZN(n10563) );
  NAND2_X1 U13455 ( .A1(n10563), .A2(n10564), .ZN(n14749) );
  INV_X1 U13456 ( .A(n11030), .ZN(n10581) );
  NAND2_X1 U13457 ( .A1(n11028), .A2(n11044), .ZN(n11056) );
  NAND2_X1 U13458 ( .A1(n13010), .A2(n11016), .ZN(n10582) );
  INV_X1 U13459 ( .A(n10588), .ZN(n13009) );
  NAND2_X1 U13460 ( .A1(n11024), .A2(n11023), .ZN(n11062) );
  INV_X1 U13461 ( .A(n11058), .ZN(n10606) );
  NAND2_X1 U13462 ( .A1(n10000), .A2(n10747), .ZN(n10611) );
  NAND2_X1 U13463 ( .A1(n10783), .A2(n10781), .ZN(n10612) );
  OAI21_X1 U13464 ( .B1(n10783), .B2(n10781), .A(n10784), .ZN(n10613) );
  NAND2_X1 U13465 ( .A1(n10929), .A2(n10616), .ZN(n10615) );
  AND2_X1 U13466 ( .A1(n19118), .A2(n13322), .ZN(n13326) );
  INV_X4 U13467 ( .A(n14596), .ZN(n18736) );
  INV_X1 U13468 ( .A(n14732), .ZN(n14333) );
  NOR2_X1 U13469 ( .A1(n14732), .A2(n14338), .ZN(n14764) );
  AOI21_X2 U13470 ( .B1(n16969), .B2(n17259), .A(n16968), .ZN(n17270) );
  NAND2_X1 U13471 ( .A1(n16640), .A2(n16546), .ZN(n16547) );
  NAND2_X1 U13472 ( .A1(n16566), .A2(n16565), .ZN(n16569) );
  NAND2_X1 U13473 ( .A1(n16548), .A2(n16547), .ZN(n16566) );
  NAND2_X1 U13474 ( .A1(n12853), .A2(n20982), .ZN(n12867) );
  NAND2_X1 U13475 ( .A1(n12641), .A2(n12640), .ZN(n12642) );
  AND2_X1 U13476 ( .A1(n14403), .A2(n14402), .ZN(n21503) );
  NAND2_X1 U13477 ( .A1(n11896), .A2(n11872), .ZN(n11864) );
  INV_X1 U13478 ( .A(n11988), .ZN(n14366) );
  AND2_X1 U13479 ( .A1(n11988), .A2(n20939), .ZN(n11989) );
  OR2_X1 U13480 ( .A1(n9688), .A2(n21728), .ZN(n15476) );
  INV_X1 U13481 ( .A(n16681), .ZN(n16410) );
  NOR2_X1 U13482 ( .A1(n10056), .A2(n15668), .ZN(n15414) );
  OR2_X1 U13483 ( .A1(n9688), .A2(n21804), .ZN(n15439) );
  OR2_X1 U13484 ( .A1(n9688), .A2(n15677), .ZN(n13077) );
  INV_X1 U13485 ( .A(n11056), .ZN(n11024) );
  INV_X1 U13486 ( .A(n14218), .ZN(n10805) );
  AOI211_X2 U13487 ( .C1(n17195), .C2(n17155), .A(n16901), .B(n16900), .ZN(
        n16902) );
  NAND2_X1 U13488 ( .A1(n10750), .A2(n17667), .ZN(n10751) );
  INV_X1 U13489 ( .A(n16062), .ZN(n16084) );
  INV_X1 U13490 ( .A(n11465), .ZN(n10759) );
  INV_X1 U13491 ( .A(n14263), .ZN(n12101) );
  INV_X1 U13492 ( .A(n15165), .ZN(n15936) );
  NAND2_X1 U13493 ( .A1(n11202), .A2(n17526), .ZN(n10752) );
  OR2_X1 U13494 ( .A1(n13160), .A2(n17126), .ZN(n13169) );
  OR2_X1 U13495 ( .A1(n13160), .A2(n16723), .ZN(n12851) );
  AOI22_X1 U13496 ( .A1(n10696), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n9684), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10647) );
  NAND2_X1 U13497 ( .A1(n11906), .A2(n11880), .ZN(n11881) );
  AOI22_X1 U13498 ( .A1(n9715), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12019), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11840) );
  NAND2_X1 U13499 ( .A1(n14818), .A2(n14817), .ZN(n14820) );
  AOI22_X1 U13500 ( .A1(n17500), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n9699), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10678) );
  INV_X2 U13501 ( .A(n21058), .ZN(n21053) );
  AND2_X1 U13502 ( .A1(n13469), .A2(n13436), .ZN(n21110) );
  NOR2_X1 U13503 ( .A1(n12957), .A2(n12956), .ZN(n10626) );
  AND2_X1 U13504 ( .A1(n12799), .A2(n17525), .ZN(n16845) );
  OR2_X1 U13505 ( .A1(n17901), .A2(n19109), .ZN(n10627) );
  AND2_X1 U13506 ( .A1(n13169), .A2(n13168), .ZN(n10628) );
  NAND2_X2 U13507 ( .A1(n14816), .A2(n14137), .ZN(n15298) );
  AND3_X1 U13508 ( .A1(n10861), .A2(n10860), .A3(n10859), .ZN(n10629) );
  AND3_X1 U13509 ( .A1(n12241), .A2(n12240), .A3(n12239), .ZN(n10630) );
  AND3_X1 U13510 ( .A1(n12259), .A2(n12258), .A3(n12257), .ZN(n10631) );
  AND2_X1 U13511 ( .A1(n9774), .A2(n12978), .ZN(n10633) );
  NAND2_X1 U13512 ( .A1(n11382), .A2(n11381), .ZN(n10634) );
  AND2_X1 U13513 ( .A1(n15476), .A2(n15474), .ZN(n10635) );
  AND2_X1 U13514 ( .A1(n17025), .A2(n17008), .ZN(n10636) );
  NAND2_X1 U13515 ( .A1(n9688), .A2(n21728), .ZN(n10637) );
  AND2_X1 U13516 ( .A1(n12993), .A2(n12984), .ZN(n10638) );
  NAND3_X1 U13517 ( .A1(n11279), .A2(n11278), .A3(n11277), .ZN(n10639) );
  AND3_X1 U13518 ( .A1(n17055), .A2(n17069), .A3(n17056), .ZN(n10640) );
  INV_X1 U13519 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n12894) );
  INV_X1 U13520 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n12883) );
  INV_X1 U13521 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n13142) );
  OR2_X1 U13522 ( .A1(n16000), .A2(n12962), .ZN(n10641) );
  INV_X1 U13523 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n11696) );
  INV_X1 U13524 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11693) );
  INV_X1 U13525 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n19560) );
  INV_X1 U13526 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n13316) );
  AND3_X1 U13527 ( .A1(n12223), .A2(n12222), .A3(n12221), .ZN(n10642) );
  INV_X1 U13528 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n11692) );
  NOR2_X1 U13529 ( .A1(n19098), .A2(n19237), .ZN(n19082) );
  OR2_X1 U13530 ( .A1(n11732), .A2(n11731), .ZN(P3_U2640) );
  INV_X1 U13531 ( .A(n15783), .ZN(n12589) );
  NAND2_X1 U13532 ( .A1(n11890), .A2(n12650), .ZN(n12674) );
  NAND2_X1 U13533 ( .A1(n18785), .A2(n18787), .ZN(n18770) );
  AND3_X1 U13534 ( .A1(n12984), .A2(n12983), .A3(n12982), .ZN(n10645) );
  NAND2_X1 U13535 ( .A1(n14136), .A2(n11855), .ZN(n11863) );
  INV_X1 U13536 ( .A(n13440), .ZN(n12573) );
  INV_X1 U13537 ( .A(n12741), .ZN(n11879) );
  NAND2_X1 U13538 ( .A1(n13450), .A2(n11879), .ZN(n11880) );
  INV_X1 U13539 ( .A(n10743), .ZN(n10744) );
  INV_X1 U13540 ( .A(n12570), .ZN(n12586) );
  OR2_X1 U13541 ( .A1(n11982), .A2(n11981), .ZN(n11984) );
  NAND2_X1 U13542 ( .A1(n10818), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n10824) );
  NOR2_X1 U13543 ( .A1(n16945), .A2(n16933), .ZN(n12994) );
  AND2_X1 U13544 ( .A1(n21147), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n12609) );
  NAND2_X1 U13545 ( .A1(n11889), .A2(n15147), .ZN(n11894) );
  AND2_X1 U13546 ( .A1(n12031), .A2(n12030), .ZN(n12118) );
  INV_X1 U13547 ( .A(n12639), .ZN(n12640) );
  OR2_X1 U13548 ( .A1(n10773), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10757) );
  INV_X1 U13549 ( .A(n11198), .ZN(n11156) );
  INV_X1 U13550 ( .A(n10796), .ZN(n10789) );
  AND2_X1 U13551 ( .A1(n11875), .A2(n14097), .ZN(n11877) );
  AND4_X1 U13552 ( .A1(n11902), .A2(n11901), .A3(n11900), .A4(n11899), .ZN(
        n11903) );
  OR2_X1 U13553 ( .A1(n12502), .A2(n15807), .ZN(n11786) );
  AND2_X1 U13554 ( .A1(n15849), .A2(n15863), .ZN(n15857) );
  AOI22_X1 U13555 ( .A1(n11995), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12019), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11761) );
  AOI22_X1 U13556 ( .A1(n11824), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11797), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11834) );
  NAND2_X1 U13557 ( .A1(n14218), .A2(n14217), .ZN(n14223) );
  INV_X1 U13558 ( .A(n16644), .ZN(n16538) );
  INV_X1 U13559 ( .A(n16931), .ZN(n16932) );
  INV_X1 U13560 ( .A(n14562), .ZN(n11250) );
  INV_X1 U13561 ( .A(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n13701) );
  INV_X1 U13562 ( .A(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n21699) );
  AND2_X1 U13563 ( .A1(n13296), .A2(n13360), .ZN(n13240) );
  AND2_X1 U13564 ( .A1(n13368), .A2(n14167), .ZN(n13290) );
  NAND2_X1 U13565 ( .A1(n12612), .A2(n12611), .ZN(n12629) );
  INV_X1 U13566 ( .A(n12414), .ZN(n12415) );
  OAI21_X1 U13567 ( .B1(n12606), .B2(n12018), .A(n12017), .ZN(n12112) );
  INV_X1 U13568 ( .A(n11896), .ZN(n15934) );
  OR2_X1 U13569 ( .A1(n12674), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12681) );
  NAND2_X1 U13570 ( .A1(n14275), .A2(n13106), .ZN(n15500) );
  NAND2_X1 U13571 ( .A1(n11914), .A2(n11917), .ZN(n11918) );
  INV_X1 U13572 ( .A(n12629), .ZN(n12618) );
  NAND2_X1 U13573 ( .A1(n12940), .A2(n16008), .ZN(n15989) );
  INV_X1 U13574 ( .A(n11080), .ZN(n11070) );
  OR2_X1 U13575 ( .A1(n16480), .A2(n16479), .ZN(n16499) );
  INV_X1 U13576 ( .A(n16682), .ZN(n16409) );
  INV_X1 U13577 ( .A(n16159), .ZN(n11376) );
  INV_X1 U13578 ( .A(n14519), .ZN(n11411) );
  AND2_X1 U13579 ( .A1(n11711), .A2(n11710), .ZN(n13335) );
  AND2_X1 U13580 ( .A1(n18787), .A2(n11687), .ZN(n13356) );
  NOR2_X1 U13581 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n13317) );
  INV_X1 U13582 ( .A(n12537), .ZN(n12560) );
  INV_X1 U13583 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n15025) );
  AND2_X1 U13584 ( .A1(n12688), .A2(n12687), .ZN(n15037) );
  OAI21_X1 U13585 ( .B1(n9850), .B2(n15819), .A(n21473), .ZN(n15841) );
  NAND2_X1 U13586 ( .A1(n11926), .A2(n11925), .ZN(n14457) );
  INV_X1 U13587 ( .A(n11089), .ZN(n11085) );
  INV_X1 U13588 ( .A(n11062), .ZN(n11027) );
  INV_X1 U13589 ( .A(n13532), .ZN(n11426) );
  INV_X1 U13590 ( .A(n14037), .ZN(n14217) );
  OR2_X1 U13591 ( .A1(n16535), .A2(n16642), .ZN(n16564) );
  AND2_X1 U13592 ( .A1(n12767), .A2(n12766), .ZN(n16075) );
  OR2_X1 U13593 ( .A1(n11101), .A2(n17315), .ZN(n16999) );
  INV_X1 U13594 ( .A(n17237), .ZN(n17394) );
  NAND2_X1 U13595 ( .A1(n13855), .A2(n11175), .ZN(n11162) );
  INV_X1 U13596 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n11386) );
  INV_X2 U13597 ( .A(n14593), .ZN(n13718) );
  INV_X1 U13598 ( .A(n20065), .ZN(n20149) );
  INV_X1 U13599 ( .A(n19325), .ZN(n17904) );
  AND2_X1 U13600 ( .A1(n19016), .A2(n13330), .ZN(n13331) );
  AND2_X1 U13601 ( .A1(n13355), .A2(n13354), .ZN(n14316) );
  NAND2_X1 U13602 ( .A1(n12416), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12440) );
  OR2_X1 U13603 ( .A1(n20968), .A2(n20967), .ZN(n21011) );
  NOR2_X1 U13604 ( .A1(n15149), .A2(n13146), .ZN(n12750) );
  AND2_X1 U13605 ( .A1(n14816), .A2(n14138), .ZN(n14802) );
  NAND2_X1 U13606 ( .A1(n12368), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12414) );
  AND3_X1 U13607 ( .A1(n15022), .A2(n15053), .A3(n15069), .ZN(n15054) );
  OR3_X1 U13608 ( .A1(n15569), .A2(n15547), .A3(n15548), .ZN(n15540) );
  AND2_X1 U13609 ( .A1(n12712), .A2(n12711), .ZN(n14923) );
  AND2_X1 U13610 ( .A1(n12692), .A2(n12691), .ZN(n15024) );
  NAND2_X1 U13611 ( .A1(n13941), .A2(n13940), .ZN(n15939) );
  INV_X1 U13612 ( .A(n21202), .ZN(n14475) );
  AND2_X1 U13613 ( .A1(n14363), .A2(n21413), .ZN(n15812) );
  NAND2_X1 U13614 ( .A1(n21181), .A2(n21413), .ZN(n21354) );
  INV_X1 U13615 ( .A(n21455), .ZN(n15928) );
  INV_X1 U13616 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n21414) );
  INV_X1 U13617 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21681) );
  AOI21_X1 U13618 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n21414), .A(n15796), 
        .ZN(n21422) );
  INV_X1 U13619 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n16114) );
  INV_X1 U13620 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17002) );
  INV_X1 U13621 ( .A(n16739), .ZN(n16699) );
  XNOR2_X1 U13622 ( .A(n16542), .B(n16541), .ZN(n16640) );
  AND2_X1 U13623 ( .A1(n12765), .A2(n12764), .ZN(n16080) );
  INV_X1 U13624 ( .A(n13676), .ZN(n12798) );
  NOR2_X1 U13625 ( .A1(n13489), .A2(n13488), .ZN(n13490) );
  INV_X1 U13626 ( .A(n14759), .ZN(n16158) );
  AND2_X1 U13627 ( .A1(n11470), .A2(n11469), .ZN(n17653) );
  OR2_X1 U13628 ( .A1(n17684), .A2(n17515), .ZN(n17516) );
  AND2_X1 U13629 ( .A1(n20535), .A2(n20914), .ZN(n17542) );
  AND2_X1 U13630 ( .A1(n20888), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20905) );
  INV_X1 U13631 ( .A(n17542), .ZN(n20439) );
  NAND2_X1 U13632 ( .A1(n20535), .A2(n17543), .ZN(n20476) );
  INV_X1 U13633 ( .A(n20885), .ZN(n20350) );
  NOR3_X1 U13634 ( .A1(n20657), .A2(n20684), .A3(n20742), .ZN(n20660) );
  NOR2_X1 U13635 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n15981) );
  INV_X1 U13636 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n20742) );
  INV_X1 U13637 ( .A(n11727), .ZN(n11728) );
  OAI21_X1 U13638 ( .B1(n19051), .B2(n18518), .A(n18370), .ZN(n18330) );
  INV_X1 U13639 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n18353) );
  INV_X1 U13640 ( .A(n18523), .ZN(n18481) );
  INV_X1 U13641 ( .A(n18580), .ZN(n18567) );
  NAND2_X1 U13642 ( .A1(n14310), .A2(n13353), .ZN(n14320) );
  OR2_X1 U13643 ( .A1(n18886), .A2(n19583), .ZN(n18788) );
  INV_X1 U13644 ( .A(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13823) );
  OR2_X1 U13645 ( .A1(n17904), .A2(n19290), .ZN(n19042) );
  OR2_X1 U13646 ( .A1(n17925), .A2(n17765), .ZN(n17910) );
  INV_X1 U13647 ( .A(n19030), .ZN(n19184) );
  OR2_X1 U13648 ( .A1(n17936), .A2(n19522), .ZN(n19335) );
  NOR2_X1 U13649 ( .A1(n19408), .A2(n19165), .ZN(n19139) );
  INV_X1 U13650 ( .A(n17955), .ZN(n19386) );
  NOR2_X1 U13651 ( .A1(n14326), .A2(n14325), .ZN(n20026) );
  NAND2_X1 U13652 ( .A1(n13979), .A2(n13354), .ZN(n17978) );
  NAND3_X1 U13653 ( .A1(n20151), .A2(n20134), .A3(P3_STATEBS16_REG_SCAN_IN), 
        .ZN(n19905) );
  AND2_X1 U13654 ( .A1(n12796), .A2(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n13676)
         );
  AND2_X1 U13655 ( .A1(n15966), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n20935) );
  AND2_X1 U13656 ( .A1(n12539), .A2(n12520), .ZN(n15312) );
  INV_X1 U13657 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n12207) );
  AND2_X1 U13658 ( .A1(n12750), .A2(n12748), .ZN(n21016) );
  AND2_X1 U13659 ( .A1(n15158), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n21019) );
  INV_X1 U13660 ( .A(n15203), .ZN(n15196) );
  AND2_X1 U13661 ( .A1(n14816), .A2(n14815), .ZN(n14817) );
  INV_X1 U13662 ( .A(n15258), .ZN(n15274) );
  NAND2_X1 U13663 ( .A1(n14816), .A2(n14139), .ZN(n15272) );
  INV_X1 U13664 ( .A(n14170), .ZN(n21077) );
  INV_X2 U13665 ( .A(n14169), .ZN(n21084) );
  INV_X1 U13666 ( .A(n15504), .ZN(n21088) );
  INV_X1 U13667 ( .A(n20943), .ZN(n21095) );
  INV_X1 U13668 ( .A(n21376), .ZN(n21417) );
  AND2_X1 U13669 ( .A1(n18043), .A2(n13943), .ZN(n21599) );
  INV_X1 U13670 ( .A(n21201), .ZN(n21169) );
  AND2_X1 U13671 ( .A1(n14524), .A2(n15789), .ZN(n21233) );
  OAI211_X1 U13672 ( .C1(n21210), .C2(n21209), .A(n21208), .B(n21305), .ZN(
        n21227) );
  AND2_X1 U13673 ( .A1(n21233), .A2(n15812), .ZN(n21261) );
  AND2_X1 U13674 ( .A1(n21268), .A2(n15847), .ZN(n21292) );
  OAI21_X1 U13675 ( .B1(n21310), .B2(n21309), .A(n21308), .ZN(n21342) );
  NOR2_X2 U13676 ( .A1(n21273), .A2(n14475), .ZN(n21341) );
  INV_X1 U13677 ( .A(n21375), .ZN(n15894) );
  INV_X1 U13678 ( .A(n21391), .ZN(n21932) );
  OAI211_X1 U13679 ( .C1(n21376), .C2(n21384), .A(n14527), .B(n21422), .ZN(
        n14552) );
  INV_X1 U13680 ( .A(n15896), .ZN(n15930) );
  AND2_X1 U13681 ( .A1(n21419), .A2(n14364), .ZN(n21455) );
  OAI21_X1 U13682 ( .B1(n21424), .B2(n21423), .A(n21422), .ZN(n21456) );
  AND2_X1 U13683 ( .A1(n11872), .A2(n14402), .ZN(n21491) );
  AND2_X1 U13684 ( .A1(n14385), .A2(n14402), .ZN(n21516) );
  INV_X1 U13685 ( .A(n21439), .ZN(n21493) );
  INV_X1 U13686 ( .A(n21451), .ZN(n21511) );
  AND2_X1 U13687 ( .A1(n20939), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13578) );
  INV_X1 U13688 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n21527) );
  NAND2_X1 U13689 ( .A1(n21527), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n21576) );
  AND3_X1 U13690 ( .A1(n11173), .A2(n17654), .A3(n12868), .ZN(n13603) );
  AND2_X1 U13691 ( .A1(n11186), .A2(n11185), .ZN(n20927) );
  INV_X1 U13692 ( .A(n17996), .ZN(n20204) );
  AND2_X1 U13693 ( .A1(n11176), .A2(n11185), .ZN(n17654) );
  OR2_X1 U13694 ( .A1(n11289), .A2(n11288), .ZN(n16731) );
  NOR3_X1 U13695 ( .A1(n14506), .A2(n17541), .A3(n17535), .ZN(n16698) );
  XNOR2_X1 U13696 ( .A(n14075), .B(n14074), .ZN(n20903) );
  INV_X1 U13697 ( .A(n14763), .ZN(n16869) );
  INV_X1 U13698 ( .A(n12798), .ZN(n17525) );
  INV_X1 U13699 ( .A(n20256), .ZN(n17155) );
  INV_X1 U13700 ( .A(n13059), .ZN(n13060) );
  NAND2_X1 U13701 ( .A1(n14785), .A2(n14784), .ZN(n14786) );
  AND2_X1 U13702 ( .A1(n11523), .A2(n11211), .ZN(n20277) );
  INV_X1 U13703 ( .A(n20290), .ZN(n20267) );
  OAI21_X1 U13704 ( .B1(n17523), .B2(n17522), .A(n17521), .ZN(n20317) );
  NOR2_X1 U13705 ( .A1(n17514), .A2(n20692), .ZN(n17519) );
  NAND2_X1 U13706 ( .A1(n20748), .A2(n20905), .ZN(n17547) );
  OAI21_X1 U13707 ( .B1(n20360), .B2(n20359), .A(n20358), .ZN(n20378) );
  AND2_X1 U13708 ( .A1(n20445), .A2(n20438), .ZN(n20461) );
  NOR2_X2 U13709 ( .A1(n20439), .A2(n20747), .ZN(n20493) );
  OAI21_X1 U13710 ( .B1(n20507), .B2(n20506), .A(n20505), .ZN(n20530) );
  INV_X1 U13711 ( .A(n20601), .ZN(n20562) );
  OAI21_X1 U13712 ( .B1(n17615), .B2(n20595), .A(n20748), .ZN(n20598) );
  OAI21_X1 U13713 ( .B1(n20602), .B2(n17618), .A(n17617), .ZN(n20596) );
  NOR2_X2 U13714 ( .A1(n20667), .A2(n20350), .ZN(n20652) );
  NOR2_X2 U13715 ( .A1(n20690), .A2(n20666), .ZN(n20686) );
  INV_X1 U13716 ( .A(n20730), .ZN(n20732) );
  INV_X1 U13717 ( .A(n20709), .ZN(n20766) );
  INV_X1 U13718 ( .A(n20724), .ZN(n20790) );
  INV_X1 U13719 ( .A(n17687), .ZN(n20819) );
  INV_X1 U13720 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n20827) );
  NAND2_X1 U13721 ( .A1(n13350), .A2(n13349), .ZN(n20022) );
  NOR2_X1 U13722 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n18363), .ZN(n18347) );
  NOR2_X1 U13723 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n18383), .ZN(n18367) );
  INV_X1 U13724 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n18410) );
  NOR2_X1 U13725 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n18458), .ZN(n18440) );
  NOR2_X1 U13726 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n18507), .ZN(n18490) );
  NAND2_X1 U13727 ( .A1(n20169), .A2(n11712), .ZN(n11718) );
  NOR2_X1 U13728 ( .A1(n18676), .A2(n18677), .ZN(n18656) );
  NOR4_X1 U13729 ( .A1(n13833), .A2(n18364), .A3(n13832), .A4(n13831), .ZN(
        n13885) );
  INV_X1 U13730 ( .A(n18785), .ZN(n13832) );
  OAI22_X1 U13731 ( .A1(n20022), .A2(n14320), .B1(n13690), .B2(n13689), .ZN(
        n14154) );
  INV_X1 U13732 ( .A(n18863), .ZN(n18827) );
  OR2_X1 U13733 ( .A1(n13269), .A2(n13268), .ZN(n18887) );
  INV_X1 U13734 ( .A(n18883), .ZN(n18889) );
  INV_X1 U13735 ( .A(n18996), .ZN(n18987) );
  AND2_X1 U13736 ( .A1(n13559), .A2(n19594), .ZN(n19148) );
  OR2_X1 U13737 ( .A1(n19042), .A2(n19035), .ZN(n19043) );
  AND2_X1 U13738 ( .A1(n17845), .A2(n19336), .ZN(n19050) );
  AND2_X1 U13739 ( .A1(n19277), .A2(n17908), .ZN(n19141) );
  AND2_X1 U13740 ( .A1(n19277), .A2(n18887), .ZN(n19191) );
  NAND2_X1 U13741 ( .A1(n19145), .A2(n19271), .ZN(n19278) );
  OR2_X2 U13742 ( .A1(n20023), .A2(n19532), .ZN(n19467) );
  AND2_X1 U13743 ( .A1(n19545), .A2(n18887), .ZN(n19478) );
  INV_X1 U13744 ( .A(n19551), .ZN(n19527) );
  AND2_X1 U13745 ( .A1(n19546), .A2(n13983), .ZN(n19545) );
  NAND2_X1 U13746 ( .A1(n20156), .A2(n19563), .ZN(n19592) );
  CLKBUF_X1 U13747 ( .A(n19654), .Z(n19688) );
  INV_X1 U13748 ( .A(n19732), .ZN(n19734) );
  INV_X1 U13749 ( .A(n19826), .ZN(n19819) );
  NOR2_X1 U13750 ( .A1(n19592), .A2(n19905), .ZN(n19877) );
  INV_X1 U13751 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n20062) );
  INV_X1 U13752 ( .A(U212), .ZN(n18142) );
  INV_X1 U13753 ( .A(n12759), .ZN(n12760) );
  INV_X1 U13754 ( .A(n20992), .ZN(n21026) );
  INV_X1 U13755 ( .A(n21027), .ZN(n21015) );
  NAND2_X1 U13756 ( .A1(n21060), .A2(n21615), .ZN(n21058) );
  NOR2_X1 U13757 ( .A1(n14044), .A2(n14043), .ZN(n14170) );
  NAND2_X1 U13758 ( .A1(n15504), .A2(n14090), .ZN(n21098) );
  NAND2_X1 U13759 ( .A1(n13578), .A2(n14372), .ZN(n15511) );
  NAND2_X1 U13760 ( .A1(n13469), .A2(n13438), .ZN(n21125) );
  INV_X1 U13761 ( .A(n21110), .ZN(n21139) );
  INV_X1 U13762 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13958) );
  AOI21_X1 U13763 ( .B1(n15799), .B2(n15803), .A(n15798), .ZN(n21173) );
  NAND2_X1 U13764 ( .A1(n21233), .A2(n15847), .ZN(n21201) );
  AOI22_X1 U13765 ( .A1(n21204), .A2(n21209), .B1(n21382), .B2(n21299), .ZN(
        n21230) );
  AOI22_X1 U13766 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n21238), .B1(n21239), 
        .B2(n21242), .ZN(n21266) );
  INV_X1 U13767 ( .A(n21261), .ZN(n15846) );
  NAND2_X1 U13768 ( .A1(n21268), .A2(n21267), .ZN(n21339) );
  AOI22_X1 U13769 ( .A1(n21300), .A2(n21309), .B1(n21299), .B2(n21460), .ZN(
        n21345) );
  INV_X1 U13770 ( .A(n15889), .ZN(n14505) );
  NAND2_X1 U13771 ( .A1(n15848), .A2(n15847), .ZN(n21375) );
  AOI22_X1 U13772 ( .A1(n21389), .A2(n21383), .B1(n21382), .B2(n21381), .ZN(
        n21937) );
  NAND2_X1 U13773 ( .A1(n15848), .A2(n21202), .ZN(n21391) );
  OR2_X1 U13774 ( .A1(n15266), .A2(n15796), .ZN(n21397) );
  NAND2_X1 U13775 ( .A1(n21419), .A2(n21413), .ZN(n21524) );
  OR2_X1 U13776 ( .A1(n14373), .A2(n21413), .ZN(n21476) );
  INV_X1 U13777 ( .A(n21591), .ZN(n21526) );
  INV_X1 U13778 ( .A(n21576), .ZN(n21625) );
  INV_X1 U13779 ( .A(n21577), .ZN(n21583) );
  INV_X1 U13780 ( .A(n13623), .ZN(n15982) );
  AND2_X1 U13781 ( .A1(n20256), .A2(n20249), .ZN(n20182) );
  NAND2_X1 U13782 ( .A1(n15982), .A2(n12959), .ZN(n20196) );
  INV_X1 U13783 ( .A(n20195), .ZN(n17991) );
  NAND2_X1 U13784 ( .A1(n16723), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n12850) );
  AND2_X1 U13785 ( .A1(n12849), .A2(n20180), .ZN(n16728) );
  OR2_X1 U13786 ( .A1(n16867), .A2(n10734), .ZN(n16855) );
  INV_X1 U13787 ( .A(n16867), .ZN(n16744) );
  OR2_X1 U13788 ( .A1(n16867), .A2(n11227), .ZN(n16872) );
  NAND2_X1 U13789 ( .A1(n20238), .A2(n13855), .ZN(n20211) );
  OR2_X1 U13790 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n20911), .ZN(n20240) );
  OR2_X1 U13791 ( .A1(n20238), .A2(n20243), .ZN(n20241) );
  INV_X1 U13792 ( .A(n13686), .ZN(n13852) );
  NAND2_X1 U13793 ( .A1(n13056), .A2(n18013), .ZN(n20249) );
  NAND2_X1 U13794 ( .A1(n11523), .A2(n20921), .ZN(n20290) );
  INV_X1 U13795 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n17989) );
  AOI21_X1 U13796 ( .B1(n17519), .B2(n17522), .A(n17518), .ZN(n20321) );
  OAI22_X1 U13797 ( .A1(n17548), .A2(n17547), .B1(n20661), .B2(n17546), .ZN(
        n17599) );
  INV_X1 U13798 ( .A(n20387), .ZN(n20412) );
  AND2_X1 U13799 ( .A1(n17604), .A2(n17603), .ZN(n20435) );
  INV_X1 U13800 ( .A(n20440), .ZN(n20465) );
  INV_X1 U13801 ( .A(n20499), .ZN(n20534) );
  AOI21_X1 U13802 ( .B1(n20540), .B2(n20543), .A(n20537), .ZN(n20582) );
  OR2_X1 U13803 ( .A1(n20667), .A2(n20497), .ZN(n20601) );
  AOI21_X1 U13804 ( .B1(n17628), .B2(n17627), .A(n17626), .ZN(n20656) );
  INV_X1 U13805 ( .A(n20686), .ZN(n20683) );
  OR2_X1 U13806 ( .A1(n20667), .A2(n20666), .ZN(n20730) );
  OR2_X1 U13807 ( .A1(n20690), .A2(n20747), .ZN(n20805) );
  INV_X1 U13808 ( .A(n20884), .ZN(n20881) );
  INV_X1 U13809 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n20830) );
  INV_X1 U13810 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n20156) );
  INV_X1 U13811 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n18510) );
  INV_X1 U13812 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n18544) );
  NAND2_X1 U13813 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n18643), .ZN(n18638) );
  INV_X1 U13814 ( .A(n18770), .ZN(n18749) );
  AND2_X1 U13815 ( .A1(n14154), .A2(n13692), .ZN(n18785) );
  OR2_X1 U13816 ( .A1(n18886), .A2(n17706), .ZN(n18863) );
  INV_X1 U13817 ( .A(n13362), .ZN(n14243) );
  INV_X1 U13818 ( .A(n18888), .ZN(n18832) );
  INV_X1 U13819 ( .A(n18908), .ZN(n18912) );
  INV_X1 U13820 ( .A(n18928), .ZN(n18934) );
  INV_X1 U13821 ( .A(n19050), .ZN(n19123) );
  INV_X1 U13822 ( .A(n19191), .ZN(n19109) );
  INV_X1 U13823 ( .A(n19275), .ZN(n19267) );
  OAI21_X2 U13824 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n20158), .A(n18193), 
        .ZN(n19271) );
  INV_X1 U13825 ( .A(n19478), .ZN(n19364) );
  AND3_X1 U13826 ( .A1(n17958), .A2(n17957), .A3(n17956), .ZN(n19461) );
  OR2_X1 U13827 ( .A1(n19546), .A2(n19494), .ZN(n19551) );
  INV_X2 U13828 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14338) );
  INV_X1 U13829 ( .A(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n21742) );
  INV_X1 U13830 ( .A(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n19624) );
  INV_X1 U13831 ( .A(n19711), .ZN(n19709) );
  INV_X1 U13832 ( .A(n19873), .ZN(n19949) );
  INV_X1 U13833 ( .A(n19911), .ZN(n19955) );
  NAND2_X1 U13834 ( .A1(n20049), .A2(n20159), .ZN(n20047) );
  NOR2_X1 U13835 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n20154) );
  INV_X1 U13836 ( .A(n20132), .ZN(n20057) );
  INV_X1 U13837 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n20067) );
  INV_X1 U13838 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n20084) );
  INV_X1 U13839 ( .A(n20121), .ZN(n20164) );
  NOR2_X1 U13840 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n13522), .ZN(n18174)
         );
  INV_X1 U13841 ( .A(n18145), .ZN(n18148) );
  OR4_X1 U13842 ( .A1(n13538), .A2(n13537), .A3(n13536), .A4(n13535), .ZN(
        P2_U2844) );
  NAND2_X1 U13843 ( .A1(n12851), .A2(n12850), .ZN(P2_U2856) );
  NAND2_X1 U13844 ( .A1(n10627), .A2(n13410), .ZN(P3_U2801) );
  AOI22_X1 U13845 ( .A1(n9679), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10833), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10649) );
  AOI22_X1 U13846 ( .A1(n16446), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n16447), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10648) );
  INV_X4 U13847 ( .A(n17480), .ZN(n17500) );
  AOI22_X1 U13848 ( .A1(n17500), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n16614), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10646) );
  AOI22_X1 U13849 ( .A1(n17500), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n16614), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10651) );
  AOI22_X1 U13850 ( .A1(n16446), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n16447), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10650) );
  AOI22_X1 U13851 ( .A1(n10696), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n16613), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10653) );
  AOI22_X1 U13852 ( .A1(n9680), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n10833), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10652) );
  AOI22_X1 U13853 ( .A1(n9705), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n10833), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10657) );
  AOI22_X1 U13854 ( .A1(n10696), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n16447), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10656) );
  AOI22_X1 U13855 ( .A1(n16446), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n16613), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10655) );
  AOI22_X1 U13856 ( .A1(n17500), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n9699), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10654) );
  NAND4_X1 U13857 ( .A1(n10657), .A2(n10656), .A3(n10655), .A4(n10654), .ZN(
        n10658) );
  AOI22_X1 U13858 ( .A1(n10696), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n16613), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10662) );
  AOI22_X1 U13859 ( .A1(n17500), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n16614), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10661) );
  AOI22_X1 U13860 ( .A1(n9680), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10833), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10660) );
  AOI22_X1 U13861 ( .A1(n16446), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n16447), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10659) );
  NAND4_X1 U13862 ( .A1(n10662), .A2(n10661), .A3(n10660), .A4(n10659), .ZN(
        n10663) );
  AOI22_X1 U13863 ( .A1(n10833), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n9684), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10667) );
  AOI22_X1 U13864 ( .A1(n17500), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n9699), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10666) );
  AOI22_X1 U13865 ( .A1(n16445), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n16593), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10665) );
  AOI22_X1 U13866 ( .A1(n10696), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n16446), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10664) );
  AOI22_X1 U13867 ( .A1(n16447), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n9685), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10671) );
  AOI22_X1 U13868 ( .A1(n16445), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10833), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10669) );
  AOI22_X1 U13869 ( .A1(n10696), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n16446), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10668) );
  AOI22_X1 U13870 ( .A1(n10696), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n9685), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10675) );
  AOI22_X1 U13871 ( .A1(n16446), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n16593), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10674) );
  AOI22_X1 U13872 ( .A1(n9679), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n10833), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10673) );
  AOI22_X1 U13873 ( .A1(n17500), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n16614), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10672) );
  AOI22_X1 U13874 ( .A1(n10696), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n16613), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10679) );
  AOI22_X1 U13875 ( .A1(n9705), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10833), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10677) );
  AOI22_X1 U13876 ( .A1(n16446), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n16593), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10676) );
  AOI22_X1 U13877 ( .A1(n10833), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n16613), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10683) );
  AOI22_X1 U13878 ( .A1(n10696), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n16447), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10682) );
  AOI22_X1 U13879 ( .A1(n9705), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n16446), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10681) );
  AOI22_X1 U13880 ( .A1(n17500), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n9699), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10680) );
  AOI22_X1 U13881 ( .A1(n17500), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n9698), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10687) );
  AOI22_X1 U13882 ( .A1(n16446), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n9685), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10686) );
  AOI22_X1 U13883 ( .A1(n10696), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n9705), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10685) );
  AOI22_X1 U13884 ( .A1(n16447), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10833), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10684) );
  AOI22_X1 U13885 ( .A1(n16446), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10833), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10691) );
  AOI22_X1 U13886 ( .A1(n17500), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n16614), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10690) );
  AOI22_X1 U13887 ( .A1(n16447), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n9685), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10688) );
  AOI22_X1 U13888 ( .A1(n10833), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n9685), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10695) );
  AOI22_X1 U13889 ( .A1(n17500), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n16614), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10694) );
  AOI22_X1 U13890 ( .A1(n16445), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n16447), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10693) );
  AOI22_X1 U13891 ( .A1(n10696), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n16446), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10692) );
  AOI22_X1 U13892 ( .A1(n10696), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n16593), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10700) );
  AOI22_X1 U13893 ( .A1(n9680), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n16446), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10699) );
  AOI22_X1 U13894 ( .A1(n10833), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n9684), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10698) );
  AOI22_X1 U13895 ( .A1(n17500), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n9698), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10697) );
  AOI22_X1 U13896 ( .A1(n10833), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n9685), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10704) );
  AOI22_X1 U13897 ( .A1(n17500), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n9699), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10703) );
  AOI22_X1 U13898 ( .A1(n16445), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n16446), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10702) );
  AOI22_X1 U13899 ( .A1(n10696), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n16593), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10701) );
  AOI22_X1 U13900 ( .A1(n16446), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n16613), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10708) );
  AOI22_X1 U13901 ( .A1(n10696), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10833), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10707) );
  AOI22_X1 U13902 ( .A1(n9705), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n16593), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10706) );
  AOI22_X1 U13903 ( .A1(n17500), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n16614), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10705) );
  NAND4_X1 U13904 ( .A1(n10708), .A2(n10707), .A3(n10706), .A4(n10705), .ZN(
        n10709) );
  NAND2_X1 U13905 ( .A1(n10709), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10716) );
  AOI22_X1 U13906 ( .A1(n16446), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n16613), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10713) );
  AOI22_X1 U13907 ( .A1(n17500), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n16614), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10712) );
  AOI22_X1 U13908 ( .A1(n10696), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n16593), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10711) );
  AOI22_X1 U13909 ( .A1(n9679), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10833), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10710) );
  NAND4_X1 U13910 ( .A1(n10713), .A2(n10712), .A3(n10711), .A4(n10710), .ZN(
        n10714) );
  NAND2_X1 U13911 ( .A1(n10714), .A2(n17650), .ZN(n10715) );
  NAND2_X4 U13912 ( .A1(n10716), .A2(n10715), .ZN(n17526) );
  AND2_X1 U13913 ( .A1(n9710), .A2(n17526), .ZN(n11188) );
  INV_X1 U13914 ( .A(n17526), .ZN(n10717) );
  INV_X1 U13915 ( .A(n11472), .ZN(n10718) );
  NAND2_X1 U13916 ( .A1(n17537), .A2(n10734), .ZN(n10719) );
  INV_X1 U13917 ( .A(n17526), .ZN(n17667) );
  INV_X1 U13918 ( .A(n10733), .ZN(n10722) );
  NAND2_X1 U13919 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n10725) );
  NAND3_X1 U13920 ( .A1(n10730), .A2(n9710), .A3(n11227), .ZN(n10762) );
  NAND2_X1 U13921 ( .A1(n11227), .A2(n10731), .ZN(n10737) );
  MUX2_X1 U13922 ( .A(n10734), .B(n10733), .S(n10732), .Z(n10736) );
  NAND3_X1 U13923 ( .A1(n10737), .A2(n10736), .A3(n10735), .ZN(n10738) );
  NAND2_X1 U13924 ( .A1(n10730), .A2(n10741), .ZN(n10742) );
  OAI21_X1 U13925 ( .B1(n20900), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n11386), 
        .ZN(n10746) );
  INV_X1 U13926 ( .A(n10749), .ZN(n10747) );
  INV_X1 U13927 ( .A(n15981), .ZN(n10770) );
  AOI21_X2 U13928 ( .B1(n10768), .B2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n10754), .ZN(n10781) );
  NAND2_X1 U13929 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n10755) );
  NAND2_X1 U13930 ( .A1(n10759), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10787) );
  NAND2_X1 U13931 ( .A1(n15981), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n10760) );
  AND2_X1 U13932 ( .A1(n10787), .A2(n10760), .ZN(n10761) );
  INV_X1 U13933 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n14053) );
  NAND2_X1 U13934 ( .A1(n10763), .A2(n10762), .ZN(n11475) );
  INV_X1 U13935 ( .A(n11475), .ZN(n10766) );
  INV_X1 U13936 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n20183) );
  INV_X1 U13937 ( .A(n12951), .ZN(n17697) );
  OAI21_X1 U13938 ( .B1(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n11386), .A(
        n17697), .ZN(n10764) );
  NAND2_X1 U13939 ( .A1(n10773), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n10765) );
  NAND2_X1 U13940 ( .A1(n10768), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10769) );
  INV_X1 U13941 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n17135) );
  NAND2_X1 U13942 ( .A1(n10773), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n10775) );
  NAND2_X1 U13943 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n10774) );
  OAI211_X1 U13944 ( .C1(n10726), .C2(n17135), .A(n10775), .B(n10774), .ZN(
        n10776) );
  BUF_X4 U13945 ( .A(n10792), .Z(n10806) );
  XNOR2_X2 U13946 ( .A(n10780), .B(n10779), .ZN(n14068) );
  INV_X1 U13947 ( .A(n10781), .ZN(n10782) );
  INV_X1 U13949 ( .A(n10785), .ZN(n10788) );
  NAND3_X1 U13950 ( .A1(n10788), .A2(n10786), .A3(n10787), .ZN(n10796) );
  INV_X1 U13951 ( .A(n9775), .ZN(n10790) );
  INV_X1 U13952 ( .A(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10791) );
  BUF_X2 U13953 ( .A(n14218), .Z(n10798) );
  INV_X1 U13954 ( .A(n10797), .ZN(n10793) );
  NAND2_X1 U13955 ( .A1(n10794), .A2(n10793), .ZN(n10795) );
  NAND2_X1 U13956 ( .A1(n14068), .A2(n14033), .ZN(n10804) );
  INV_X1 U13957 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10799) );
  INV_X1 U13958 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n21655) );
  INV_X1 U13959 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10803) );
  NOR2_X1 U13960 ( .A1(n14068), .A2(n10091), .ZN(n10800) );
  NAND2_X1 U13961 ( .A1(n10800), .A2(n17467), .ZN(n10819) );
  INV_X1 U13962 ( .A(n17544), .ZN(n17550) );
  NAND2_X1 U13963 ( .A1(n17550), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n10802) );
  INV_X1 U13964 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n17639) );
  INV_X1 U13965 ( .A(n17467), .ZN(n14062) );
  NAND3_X1 U13966 ( .A1(n14079), .A2(n14062), .A3(n14033), .ZN(n10821) );
  INV_X1 U13967 ( .A(n10821), .ZN(n10807) );
  INV_X1 U13968 ( .A(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10812) );
  OAI211_X1 U13969 ( .C1(n20385), .C2(n10812), .A(n17984), .B(n10811), .ZN(
        n10813) );
  NOR2_X1 U13970 ( .A1(n10814), .A2(n10813), .ZN(n10827) );
  INV_X1 U13971 ( .A(n20606), .ZN(n10815) );
  NAND2_X1 U13972 ( .A1(n14218), .A2(n9904), .ZN(n10816) );
  AOI22_X1 U13973 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n10815), .B1(
        n20657), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10826) );
  INV_X1 U13974 ( .A(n10816), .ZN(n10817) );
  INV_X1 U13975 ( .A(n10915), .ZN(n10818) );
  NAND2_X1 U13976 ( .A1(n17616), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n10823) );
  NAND2_X1 U13977 ( .A1(n17520), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n10822) );
  AND3_X1 U13978 ( .A1(n10824), .A2(n10823), .A3(n10822), .ZN(n10825) );
  NAND4_X1 U13979 ( .A1(n10828), .A2(n10827), .A3(n10826), .A4(n10825), .ZN(
        n10864) );
  AND2_X2 U13980 ( .A1(n16446), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n16411) );
  AOI22_X1 U13981 ( .A1(n11190), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n16411), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10832) );
  INV_X1 U13982 ( .A(n17482), .ZN(n17497) );
  AND2_X2 U13983 ( .A1(n11191), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n16464) );
  AOI22_X1 U13984 ( .A1(n10841), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n16464), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10831) );
  AND2_X2 U13985 ( .A1(n10696), .A2(n17650), .ZN(n16466) );
  AND2_X2 U13986 ( .A1(n11191), .A2(n14023), .ZN(n16465) );
  AOI22_X1 U13987 ( .A1(n16466), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n16465), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10830) );
  AOI22_X1 U13988 ( .A1(n10842), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10891), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10829) );
  NAND4_X1 U13989 ( .A1(n10832), .A2(n10831), .A3(n10830), .A4(n10829), .ZN(
        n10840) );
  AOI22_X1 U13990 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n16472), .B1(
        n16471), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10838) );
  AOI22_X1 U13991 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n16473), .B1(
        n17505), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10837) );
  AND2_X2 U13992 ( .A1(n16448), .A2(n10834), .ZN(n16437) );
  AOI22_X1 U13993 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n10848), .B1(
        n16437), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10836) );
  AOI22_X1 U13994 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n10847), .B1(
        n16438), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10835) );
  NAND4_X1 U13995 ( .A1(n10838), .A2(n10837), .A3(n10836), .A4(n10835), .ZN(
        n10839) );
  AND2_X1 U13996 ( .A1(n9710), .A2(n11499), .ZN(n11498) );
  AOI22_X1 U13997 ( .A1(n11190), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n16466), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10846) );
  AOI22_X1 U13998 ( .A1(n10841), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n16465), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10845) );
  AOI22_X1 U13999 ( .A1(n10842), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10891), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10844) );
  AOI22_X1 U14000 ( .A1(n16411), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n16464), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10843) );
  NAND4_X1 U14001 ( .A1(n10846), .A2(n10845), .A3(n10844), .A4(n10843), .ZN(
        n10854) );
  AOI22_X1 U14002 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n16472), .B1(
        n16471), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10852) );
  AOI22_X1 U14003 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n16473), .B1(
        n17505), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10851) );
  AOI22_X1 U14004 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n10847), .B1(
        n16437), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10850) );
  AOI22_X1 U14005 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n10848), .B1(
        n16438), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10849) );
  NAND4_X1 U14006 ( .A1(n10852), .A2(n10851), .A3(n10850), .A4(n10849), .ZN(
        n10853) );
  NAND2_X1 U14007 ( .A1(n11498), .A2(n11500), .ZN(n11505) );
  AOI22_X1 U14008 ( .A1(n11190), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n16411), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10855) );
  AOI22_X1 U14009 ( .A1(n10841), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n16464), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10856) );
  AOI22_X1 U14010 ( .A1(n16466), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n16465), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10857) );
  AOI22_X1 U14011 ( .A1(n10842), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10891), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10858) );
  AOI22_X1 U14012 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n16472), .B1(
        n16471), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10862) );
  AOI22_X1 U14013 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n16473), .B1(
        n17505), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10861) );
  AOI22_X1 U14014 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n10847), .B1(
        n16438), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10860) );
  AOI22_X1 U14015 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n10848), .B1(
        n16437), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10859) );
  NAND2_X1 U14016 ( .A1(n11505), .A2(n11504), .ZN(n10863) );
  INV_X1 U14017 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n20307) );
  INV_X1 U14018 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10865) );
  INV_X1 U14019 ( .A(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10866) );
  NOR2_X1 U14020 ( .A1(n10868), .A2(n10867), .ZN(n10889) );
  INV_X1 U14021 ( .A(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10871) );
  INV_X1 U14022 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10870) );
  OAI22_X1 U14023 ( .A1(n10871), .A2(n17544), .B1(n10869), .B2(n10870), .ZN(
        n10874) );
  INV_X1 U14024 ( .A(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10872) );
  NOR2_X1 U14025 ( .A1(n10874), .A2(n10873), .ZN(n10888) );
  INV_X1 U14026 ( .A(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n20421) );
  INV_X1 U14027 ( .A(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10875) );
  OAI22_X1 U14028 ( .A1(n20421), .A2(n10929), .B1(n20352), .B2(n10875), .ZN(
        n10879) );
  INV_X1 U14029 ( .A(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10877) );
  INV_X1 U14030 ( .A(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10876) );
  OAI22_X1 U14031 ( .A1(n10877), .A2(n10926), .B1(n20467), .B2(n10876), .ZN(
        n10878) );
  NOR2_X1 U14032 ( .A1(n10879), .A2(n10878), .ZN(n10887) );
  INV_X1 U14033 ( .A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10881) );
  INV_X1 U14034 ( .A(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10880) );
  INV_X1 U14035 ( .A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10883) );
  INV_X1 U14036 ( .A(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10882) );
  OAI22_X1 U14037 ( .A1(n10954), .A2(n10883), .B1(n10882), .B2(n10915), .ZN(
        n10884) );
  NOR2_X1 U14038 ( .A1(n10885), .A2(n10884), .ZN(n10886) );
  NAND4_X1 U14039 ( .A1(n10889), .A2(n10888), .A3(n10887), .A4(n10886), .ZN(
        n10890) );
  INV_X4 U14040 ( .A(n9710), .ZN(n17984) );
  NAND2_X1 U14041 ( .A1(n10890), .A2(n17984), .ZN(n10903) );
  AOI22_X1 U14042 ( .A1(n11190), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n16411), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10895) );
  AOI22_X1 U14043 ( .A1(n10841), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n16464), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10894) );
  AOI22_X1 U14044 ( .A1(n16466), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n16465), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10893) );
  AOI22_X1 U14045 ( .A1(n10842), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10891), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10892) );
  NAND4_X1 U14046 ( .A1(n10895), .A2(n10894), .A3(n10893), .A4(n10892), .ZN(
        n10901) );
  AOI22_X1 U14047 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n16472), .B1(
        n16471), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10899) );
  AOI22_X1 U14048 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n16473), .B1(
        n17505), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10898) );
  AOI22_X1 U14049 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n10848), .B1(
        n16437), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10897) );
  AOI22_X1 U14050 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n10847), .B1(
        n16438), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10896) );
  NAND4_X1 U14051 ( .A1(n10899), .A2(n10898), .A3(n10897), .A4(n10896), .ZN(
        n10900) );
  NAND2_X1 U14052 ( .A1(n11246), .A2(n9710), .ZN(n10902) );
  AOI22_X1 U14053 ( .A1(n11190), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n16411), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10907) );
  AOI22_X1 U14054 ( .A1(n10841), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n16464), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10906) );
  AOI22_X1 U14055 ( .A1(n16466), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n16465), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10905) );
  AOI22_X1 U14056 ( .A1(n10842), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10891), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10904) );
  NAND4_X1 U14057 ( .A1(n10907), .A2(n10906), .A3(n10905), .A4(n10904), .ZN(
        n10913) );
  AOI22_X1 U14058 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n16472), .B1(
        n16471), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10911) );
  AOI22_X1 U14059 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n16473), .B1(
        n17505), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10910) );
  AOI22_X1 U14060 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n10848), .B1(
        n16437), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10909) );
  AOI22_X1 U14061 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n10847), .B1(
        n16438), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10908) );
  NAND4_X1 U14062 ( .A1(n10911), .A2(n10910), .A3(n10909), .A4(n10908), .ZN(
        n10912) );
  INV_X1 U14063 ( .A(n11251), .ZN(n10914) );
  INV_X1 U14064 ( .A(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10917) );
  INV_X1 U14065 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10916) );
  OAI22_X1 U14066 ( .A1(n10917), .A2(n20541), .B1(n20740), .B2(n10916), .ZN(
        n10921) );
  INV_X1 U14067 ( .A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10919) );
  INV_X1 U14068 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10918) );
  OAI22_X1 U14069 ( .A1(n10919), .A2(n10954), .B1(n20606), .B2(n10918), .ZN(
        n10920) );
  NOR2_X1 U14070 ( .A1(n10921), .A2(n10920), .ZN(n10940) );
  INV_X1 U14071 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17535) );
  INV_X1 U14072 ( .A(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10923) );
  INV_X1 U14073 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10922) );
  NOR2_X1 U14074 ( .A1(n10925), .A2(n10924), .ZN(n10939) );
  INV_X1 U14075 ( .A(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10928) );
  INV_X1 U14076 ( .A(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10927) );
  OAI22_X1 U14077 ( .A1(n10928), .A2(n10926), .B1(n20467), .B2(n10927), .ZN(
        n10933) );
  INV_X1 U14078 ( .A(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10931) );
  INV_X1 U14079 ( .A(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10930) );
  OAI22_X1 U14080 ( .A1(n10931), .A2(n20352), .B1(n10929), .B2(n10930), .ZN(
        n10932) );
  NOR2_X1 U14081 ( .A1(n10933), .A2(n10932), .ZN(n10938) );
  INV_X1 U14082 ( .A(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n17583) );
  INV_X1 U14083 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10934) );
  OAI22_X1 U14084 ( .A1(n17583), .A2(n17544), .B1(n10869), .B2(n10934), .ZN(
        n10936) );
  NOR2_X1 U14085 ( .A1(n10936), .A2(n10935), .ZN(n10937) );
  NAND4_X1 U14086 ( .A1(n10940), .A2(n10939), .A3(n10938), .A4(n10937), .ZN(
        n10950) );
  AOI22_X1 U14087 ( .A1(n11190), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n16411), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10944) );
  AOI22_X1 U14088 ( .A1(n10841), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n16464), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10943) );
  AOI22_X1 U14089 ( .A1(n16466), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n16465), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10942) );
  AOI22_X1 U14090 ( .A1(n10842), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10891), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10941) );
  AOI22_X1 U14091 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n16472), .B1(
        n16471), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10948) );
  AOI22_X1 U14092 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n16473), .B1(
        n17505), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10947) );
  AOI22_X1 U14093 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n10848), .B1(
        n16437), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10946) );
  AOI22_X1 U14094 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n10847), .B1(
        n16438), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10945) );
  NAND2_X1 U14095 ( .A1(n11022), .A2(n9710), .ZN(n10949) );
  INV_X1 U14096 ( .A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10952) );
  INV_X1 U14097 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10951) );
  OAI22_X1 U14098 ( .A1(n10952), .A2(n20606), .B1(n20740), .B2(n10951), .ZN(
        n10957) );
  INV_X1 U14099 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10955) );
  INV_X1 U14100 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10953) );
  OAI22_X1 U14101 ( .A1(n10955), .A2(n10954), .B1(n20541), .B2(n10953), .ZN(
        n10956) );
  NOR2_X1 U14102 ( .A1(n10957), .A2(n10956), .ZN(n10975) );
  INV_X1 U14103 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17541) );
  INV_X1 U14104 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10958) );
  INV_X1 U14105 ( .A(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10959) );
  NOR2_X1 U14106 ( .A1(n10961), .A2(n10960), .ZN(n10974) );
  INV_X1 U14107 ( .A(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10963) );
  INV_X1 U14108 ( .A(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10962) );
  OAI22_X1 U14109 ( .A1(n10963), .A2(n20352), .B1(n10929), .B2(n10962), .ZN(
        n10967) );
  INV_X1 U14110 ( .A(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10965) );
  INV_X1 U14111 ( .A(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10964) );
  OAI22_X1 U14112 ( .A1(n10965), .A2(n10926), .B1(n20467), .B2(n10964), .ZN(
        n10966) );
  NOR2_X1 U14113 ( .A1(n10967), .A2(n10966), .ZN(n10973) );
  INV_X1 U14114 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10969) );
  INV_X1 U14115 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10968) );
  OAI22_X1 U14116 ( .A1(n10969), .A2(n17544), .B1(n10869), .B2(n10968), .ZN(
        n10971) );
  NOR2_X1 U14117 ( .A1(n10971), .A2(n10970), .ZN(n10972) );
  NAND4_X1 U14118 ( .A1(n10975), .A2(n10974), .A3(n10973), .A4(n10972), .ZN(
        n10987) );
  AOI22_X1 U14119 ( .A1(n11190), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n16411), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10979) );
  AOI22_X1 U14120 ( .A1(n10841), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n16464), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10978) );
  AOI22_X1 U14121 ( .A1(n16466), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n16465), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10977) );
  AOI22_X1 U14122 ( .A1(n10842), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10891), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10976) );
  NAND4_X1 U14123 ( .A1(n10979), .A2(n10978), .A3(n10977), .A4(n10976), .ZN(
        n10985) );
  AOI22_X1 U14124 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n16472), .B1(
        n16471), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10983) );
  AOI22_X1 U14125 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n16473), .B1(
        n17505), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10982) );
  AOI22_X1 U14126 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n10848), .B1(
        n16437), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10981) );
  AOI22_X1 U14127 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n10847), .B1(
        n16438), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10980) );
  NAND4_X1 U14128 ( .A1(n10983), .A2(n10982), .A3(n10981), .A4(n10980), .ZN(
        n10984) );
  INV_X1 U14129 ( .A(n11025), .ZN(n11260) );
  NAND2_X1 U14130 ( .A1(n11260), .A2(n9710), .ZN(n10986) );
  AOI22_X1 U14131 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n16466), .B1(
        n10841), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10991) );
  AOI22_X1 U14132 ( .A1(n11190), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n16411), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10990) );
  AOI22_X1 U14133 ( .A1(n10842), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n16465), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10989) );
  AOI22_X1 U14134 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n10891), .B1(
        n16464), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10988) );
  NAND4_X1 U14135 ( .A1(n10991), .A2(n10990), .A3(n10989), .A4(n10988), .ZN(
        n10997) );
  AOI22_X1 U14136 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n16472), .B1(
        n16471), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10995) );
  AOI22_X1 U14137 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n16473), .B1(
        n17505), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10994) );
  AOI22_X1 U14138 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n10848), .B1(
        n16437), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10993) );
  AOI22_X1 U14139 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n10847), .B1(
        n16438), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10992) );
  NAND4_X1 U14140 ( .A1(n10995), .A2(n10994), .A3(n10993), .A4(n10992), .ZN(
        n10996) );
  NAND2_X1 U14141 ( .A1(n11139), .A2(n11033), .ZN(n10999) );
  NAND2_X1 U14142 ( .A1(n20909), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10998) );
  NAND2_X1 U14143 ( .A1(n10999), .A2(n10998), .ZN(n11008) );
  NAND2_X1 U14144 ( .A1(n11000), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11001) );
  NAND2_X1 U14145 ( .A1(n11008), .A2(n11007), .ZN(n11003) );
  NAND2_X1 U14146 ( .A1(n11003), .A2(n11002), .ZN(n11019) );
  XNOR2_X1 U14147 ( .A(n11019), .B(n11017), .ZN(n11197) );
  INV_X1 U14148 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n11004) );
  XNOR2_X1 U14149 ( .A(n11008), .B(n11007), .ZN(n11141) );
  INV_X1 U14150 ( .A(n11141), .ZN(n11195) );
  NAND2_X1 U14151 ( .A1(n11009), .A2(n11195), .ZN(n11144) );
  NAND2_X1 U14152 ( .A1(n11178), .A2(n11012), .ZN(n11015) );
  INV_X1 U14153 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n11013) );
  NOR2_X1 U14154 ( .A1(P2_EBX_REG_1__SCAN_IN), .A2(P2_EBX_REG_0__SCAN_IN), 
        .ZN(n11016) );
  INV_X1 U14155 ( .A(n11017), .ZN(n11018) );
  NAND2_X1 U14156 ( .A1(n11019), .A2(n11018), .ZN(n11021) );
  NAND2_X1 U14157 ( .A1(n21853), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11020) );
  NAND2_X1 U14158 ( .A1(n11021), .A2(n11020), .ZN(n11153) );
  NAND2_X1 U14159 ( .A1(n17989), .A2(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(
        n11154) );
  MUX2_X1 U14160 ( .A(n11251), .B(n11198), .S(n12958), .Z(n11147) );
  INV_X1 U14161 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n14292) );
  MUX2_X1 U14162 ( .A(n11147), .B(n14292), .S(n13010), .Z(n11044) );
  INV_X1 U14163 ( .A(n11055), .ZN(n11023) );
  INV_X1 U14164 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n11026) );
  MUX2_X1 U14165 ( .A(n11026), .B(n11025), .S(n11012), .Z(n11061) );
  XNOR2_X1 U14166 ( .A(n11027), .B(n11061), .ZN(n16293) );
  INV_X1 U14167 ( .A(n11028), .ZN(n11046) );
  NAND2_X1 U14168 ( .A1(n11030), .A2(n11029), .ZN(n11031) );
  NAND2_X1 U14169 ( .A1(n11046), .A2(n11031), .ZN(n16314) );
  XNOR2_X1 U14170 ( .A(n11032), .B(n11037), .ZN(n16328) );
  XNOR2_X1 U14171 ( .A(n16328), .B(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n17150) );
  INV_X1 U14172 ( .A(n11499), .ZN(n11035) );
  INV_X1 U14173 ( .A(n11033), .ZN(n11136) );
  NAND2_X1 U14174 ( .A1(n14023), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n11034) );
  AND2_X1 U14175 ( .A1(n11136), .A2(n11034), .ZN(n11196) );
  INV_X1 U14176 ( .A(n11196), .ZN(n11140) );
  MUX2_X1 U14177 ( .A(n11035), .B(n11140), .S(n12958), .Z(n11181) );
  INV_X1 U14178 ( .A(n11181), .ZN(n11036) );
  MUX2_X1 U14179 ( .A(n11036), .B(P2_EBX_REG_0__SCAN_IN), .S(n13010), .Z(
        n16349) );
  NAND2_X1 U14180 ( .A1(n16349), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13924) );
  INV_X1 U14181 ( .A(n11037), .ZN(n11039) );
  INV_X1 U14182 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n14041) );
  NAND3_X1 U14183 ( .A1(n13010), .A2(P2_EBX_REG_0__SCAN_IN), .A3(
        P2_EBX_REG_1__SCAN_IN), .ZN(n11038) );
  NAND2_X1 U14184 ( .A1(n11039), .A2(n11038), .ZN(n13923) );
  INV_X1 U14185 ( .A(n13923), .ZN(n16337) );
  NAND2_X1 U14186 ( .A1(n16337), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n11041) );
  INV_X1 U14187 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n14054) );
  AND2_X1 U14188 ( .A1(n13923), .A2(n14054), .ZN(n11040) );
  AOI21_X1 U14189 ( .B1(n13924), .B2(n11041), .A(n11040), .ZN(n17149) );
  NAND2_X1 U14190 ( .A1(n17150), .A2(n17149), .ZN(n17148) );
  INV_X1 U14191 ( .A(n16328), .ZN(n11042) );
  NAND2_X1 U14192 ( .A1(n11042), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11043) );
  AND2_X1 U14193 ( .A1(n17148), .A2(n11043), .ZN(n17117) );
  INV_X1 U14194 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n18096) );
  INV_X1 U14195 ( .A(n11044), .ZN(n11045) );
  XNOR2_X1 U14196 ( .A(n11046), .B(n11045), .ZN(n20193) );
  INV_X1 U14197 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n20264) );
  AND2_X1 U14198 ( .A1(n20193), .A2(n20264), .ZN(n11048) );
  AOI21_X1 U14199 ( .B1(n17117), .B2(n18096), .A(n11048), .ZN(n11047) );
  INV_X1 U14200 ( .A(n17117), .ZN(n17133) );
  INV_X1 U14201 ( .A(n11048), .ZN(n11049) );
  NAND3_X1 U14202 ( .A1(n17133), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        n11049), .ZN(n11052) );
  INV_X1 U14203 ( .A(n20193), .ZN(n11050) );
  NAND2_X1 U14204 ( .A1(n11050), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11051) );
  AND2_X1 U14205 ( .A1(n11052), .A2(n11051), .ZN(n11053) );
  NAND2_X1 U14206 ( .A1(n11054), .A2(n11053), .ZN(n17104) );
  INV_X1 U14207 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n17436) );
  NAND2_X1 U14208 ( .A1(n11056), .A2(n11055), .ZN(n11057) );
  NAND2_X1 U14209 ( .A1(n11062), .A2(n11057), .ZN(n16302) );
  MUX2_X1 U14210 ( .A(n17436), .B(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .S(
        n16302), .Z(n17105) );
  NAND2_X1 U14211 ( .A1(n17104), .A2(n17105), .ZN(n11060) );
  OAI21_X1 U14212 ( .B1(P2_EBX_REG_7__SCAN_IN), .B2(n11012), .A(n13022), .ZN(
        n11063) );
  XNOR2_X1 U14213 ( .A(n11064), .B(n11063), .ZN(n16279) );
  NAND2_X1 U14214 ( .A1(n16279), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17084) );
  NAND2_X1 U14215 ( .A1(n9828), .A2(n9743), .ZN(n11065) );
  NAND2_X1 U14216 ( .A1(n11066), .A2(n11065), .ZN(n16272) );
  NOR2_X1 U14217 ( .A1(n16272), .A2(n11073), .ZN(n11074) );
  NAND2_X1 U14218 ( .A1(n11074), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n17086) );
  NAND2_X1 U14219 ( .A1(n13010), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n11067) );
  MUX2_X1 U14220 ( .A(P2_EBX_REG_10__SCAN_IN), .B(n11067), .S(n11070), .Z(
        n11068) );
  NAND2_X1 U14221 ( .A1(n11068), .A2(n13001), .ZN(n16244) );
  INV_X1 U14222 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17385) );
  OAI21_X1 U14223 ( .B1(n16244), .B2(n11073), .A(n17385), .ZN(n17055) );
  NAND2_X1 U14224 ( .A1(n11066), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n11069) );
  MUX2_X1 U14225 ( .A(n11066), .B(n11069), .S(n13010), .Z(n11071) );
  AND2_X1 U14226 ( .A1(n11071), .A2(n11070), .ZN(n16257) );
  INV_X1 U14227 ( .A(n11072), .ZN(n11073) );
  INV_X2 U14228 ( .A(n11073), .ZN(n13049) );
  NAND2_X1 U14229 ( .A1(n16257), .A2(n13049), .ZN(n11077) );
  NAND2_X1 U14230 ( .A1(n11077), .A2(n10240), .ZN(n17069) );
  NOR2_X1 U14231 ( .A1(n11074), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n17085) );
  INV_X1 U14232 ( .A(n16279), .ZN(n11075) );
  INV_X1 U14233 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18055) );
  NOR2_X1 U14234 ( .A1(n17085), .A2(n18068), .ZN(n17056) );
  INV_X1 U14235 ( .A(n16244), .ZN(n11076) );
  NAND3_X1 U14236 ( .A1(n11076), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        n13049), .ZN(n17054) );
  INV_X1 U14237 ( .A(n11077), .ZN(n11078) );
  NAND2_X1 U14238 ( .A1(n11078), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n17071) );
  INV_X1 U14239 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n16726) );
  NAND2_X1 U14240 ( .A1(n11080), .A2(n16726), .ZN(n11083) );
  INV_X1 U14241 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n11081) );
  NAND2_X2 U14242 ( .A1(n16224), .A2(n13001), .ZN(n11089) );
  NAND3_X1 U14243 ( .A1(n11083), .A2(n13010), .A3(P2_EBX_REG_11__SCAN_IN), 
        .ZN(n11084) );
  AND2_X1 U14244 ( .A1(n11085), .A2(n11084), .ZN(n13528) );
  NAND2_X1 U14245 ( .A1(n13528), .A2(n13049), .ZN(n11087) );
  INV_X1 U14246 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17372) );
  NOR2_X1 U14247 ( .A1(n11087), .A2(n17372), .ZN(n17045) );
  NAND2_X1 U14248 ( .A1(n11087), .A2(n17372), .ZN(n17043) );
  NAND2_X1 U14249 ( .A1(n13010), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n11088) );
  NAND2_X1 U14250 ( .A1(n11091), .A2(n13049), .ZN(n17034) );
  INV_X1 U14251 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n17327) );
  NAND2_X1 U14252 ( .A1(n17034), .A2(n17327), .ZN(n11090) );
  AND2_X1 U14253 ( .A1(n17043), .A2(n11090), .ZN(n12980) );
  INV_X1 U14254 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n11092) );
  NOR2_X1 U14255 ( .A1(n11012), .A2(n11092), .ZN(n11094) );
  NAND2_X1 U14256 ( .A1(n11091), .A2(n11094), .ZN(n11095) );
  AND2_X1 U14257 ( .A1(n11100), .A2(n11095), .ZN(n16208) );
  NAND3_X1 U14258 ( .A1(n16208), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(
        n13049), .ZN(n17025) );
  OR2_X1 U14259 ( .A1(n17034), .A2(n17327), .ZN(n17008) );
  INV_X1 U14260 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n11096) );
  XNOR2_X1 U14261 ( .A(n11100), .B(n9821), .ZN(n16194) );
  NAND2_X1 U14262 ( .A1(n16194), .A2(n13049), .ZN(n11097) );
  INV_X1 U14263 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n17015) );
  NAND2_X1 U14264 ( .A1(n11097), .A2(n17015), .ZN(n17012) );
  NAND2_X1 U14265 ( .A1(n16208), .A2(n13049), .ZN(n11098) );
  INV_X1 U14266 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17348) );
  NAND2_X1 U14267 ( .A1(n11098), .A2(n17348), .ZN(n17024) );
  AND2_X1 U14268 ( .A1(n13049), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11099) );
  NAND2_X1 U14269 ( .A1(n16194), .A2(n11099), .ZN(n17011) );
  NAND2_X1 U14270 ( .A1(n13010), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n11103) );
  XNOR2_X1 U14271 ( .A(n9721), .B(n11103), .ZN(n16180) );
  NAND2_X1 U14272 ( .A1(n16180), .A2(n13049), .ZN(n11101) );
  INV_X1 U14273 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n17315) );
  INV_X1 U14274 ( .A(n16999), .ZN(n11102) );
  NAND2_X1 U14275 ( .A1(n11101), .A2(n17315), .ZN(n16998) );
  INV_X1 U14276 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n11104) );
  NAND3_X1 U14277 ( .A1(n11105), .A2(n13010), .A3(P2_EBX_REG_16__SCAN_IN), 
        .ZN(n11106) );
  NAND3_X1 U14278 ( .A1(n11110), .A2(n13001), .A3(n11106), .ZN(n16171) );
  INV_X1 U14279 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n11107) );
  OAI21_X1 U14280 ( .B1(n16171), .B2(n11073), .A(n11107), .ZN(n11109) );
  NAND2_X1 U14281 ( .A1(n13049), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11108) );
  NAND2_X1 U14282 ( .A1(n11109), .A2(n12989), .ZN(n16990) );
  NAND2_X1 U14283 ( .A1(n13010), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n11112) );
  XNOR2_X1 U14284 ( .A(n11113), .B(n10309), .ZN(n16156) );
  NAND2_X1 U14285 ( .A1(n16156), .A2(n13049), .ZN(n11111) );
  INV_X1 U14286 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17292) );
  OR2_X1 U14287 ( .A1(n11111), .A2(n17292), .ZN(n12990) );
  NAND2_X1 U14288 ( .A1(n11111), .A2(n17292), .ZN(n12982) );
  NAND2_X1 U14289 ( .A1(n12990), .A2(n12982), .ZN(n16985) );
  NAND2_X1 U14290 ( .A1(n11115), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n11114) );
  MUX2_X1 U14291 ( .A(n11115), .B(n11114), .S(n13010), .Z(n11116) );
  AND2_X1 U14292 ( .A1(n13049), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11117) );
  NAND2_X1 U14293 ( .A1(n16138), .A2(n11117), .ZN(n16973) );
  NAND3_X1 U14294 ( .A1(n11118), .A2(n13010), .A3(P2_EBX_REG_19__SCAN_IN), 
        .ZN(n11121) );
  NOR2_X1 U14295 ( .A1(P2_EBX_REG_19__SCAN_IN), .A2(P2_EBX_REG_18__SCAN_IN), 
        .ZN(n11119) );
  NOR2_X1 U14296 ( .A1(n11012), .A2(n11119), .ZN(n11120) );
  NAND2_X1 U14297 ( .A1(n16122), .A2(n13049), .ZN(n11125) );
  INV_X1 U14298 ( .A(n11125), .ZN(n11122) );
  NAND2_X1 U14299 ( .A1(n11122), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n13498) );
  INV_X1 U14300 ( .A(n13498), .ZN(n11123) );
  NAND2_X1 U14301 ( .A1(n16138), .A2(n13049), .ZN(n11124) );
  INV_X1 U14302 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n14775) );
  NAND2_X1 U14303 ( .A1(n11124), .A2(n14775), .ZN(n16974) );
  INV_X1 U14304 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n11495) );
  NAND2_X1 U14305 ( .A1(n11125), .A2(n11495), .ZN(n13497) );
  NAND2_X1 U14306 ( .A1(n9767), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n11126) );
  MUX2_X1 U14307 ( .A(n11126), .B(n9767), .S(n11012), .Z(n11127) );
  NAND2_X1 U14308 ( .A1(n11127), .A2(n9723), .ZN(n16104) );
  INV_X1 U14309 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17259) );
  OAI21_X1 U14310 ( .B1(n16104), .B2(n11073), .A(n17259), .ZN(n16962) );
  INV_X1 U14311 ( .A(n16104), .ZN(n11129) );
  AND2_X1 U14312 ( .A1(n13049), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11128) );
  NAND2_X1 U14313 ( .A1(n11129), .A2(n11128), .ZN(n16961) );
  INV_X1 U14314 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n11130) );
  INV_X1 U14315 ( .A(n12945), .ZN(n11132) );
  NAND3_X1 U14316 ( .A1(n9723), .A2(n13010), .A3(P2_EBX_REG_21__SCAN_IN), .ZN(
        n11131) );
  INV_X1 U14317 ( .A(n11134), .ZN(n11133) );
  NAND2_X1 U14318 ( .A1(n11133), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12993) );
  NAND2_X1 U14319 ( .A1(n11134), .A2(n10357), .ZN(n12984) );
  NAND2_X1 U14320 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n17687) );
  INV_X1 U14321 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n20175) );
  NOR2_X1 U14322 ( .A1(n20175), .A2(n20827), .ZN(n20820) );
  NOR2_X1 U14323 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n20807) );
  NOR3_X1 U14324 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n20820), .A3(n20807), 
        .ZN(n20812) );
  INV_X1 U14325 ( .A(n20812), .ZN(n11135) );
  NOR2_X1 U14326 ( .A1(n20819), .A2(n11135), .ZN(n17658) );
  NAND2_X1 U14327 ( .A1(n17564), .A2(n17658), .ZN(n11165) );
  XNOR2_X1 U14328 ( .A(n11139), .B(n11136), .ZN(n11174) );
  OAI21_X1 U14329 ( .B1(n17984), .B2(n11196), .A(n11174), .ZN(n11137) );
  OAI21_X1 U14330 ( .B1(n11141), .B2(n17984), .A(n11137), .ZN(n11138) );
  NAND2_X1 U14331 ( .A1(n11138), .A2(n17667), .ZN(n11146) );
  INV_X1 U14332 ( .A(n11139), .ZN(n11180) );
  OAI21_X1 U14333 ( .B1(n11180), .B2(n11140), .A(n9953), .ZN(n11145) );
  NAND2_X1 U14334 ( .A1(n17526), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11161) );
  NAND2_X1 U14335 ( .A1(n11161), .A2(n17984), .ZN(n11142) );
  NAND2_X1 U14336 ( .A1(n11142), .A2(n11141), .ZN(n11143) );
  AOI22_X1 U14337 ( .A1(n11146), .A2(n11145), .B1(n11144), .B2(n11143), .ZN(
        n11151) );
  INV_X1 U14338 ( .A(n11197), .ZN(n11150) );
  NAND2_X1 U14339 ( .A1(n11148), .A2(n11147), .ZN(n11182) );
  NAND2_X1 U14340 ( .A1(n11182), .A2(n12958), .ZN(n11149) );
  OAI21_X1 U14341 ( .B1(n11151), .B2(n11150), .A(n11149), .ZN(n11158) );
  NOR2_X1 U14342 ( .A1(n17989), .A2(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(
        n11152) );
  AOI21_X1 U14343 ( .B1(n9953), .B2(n11156), .A(n11175), .ZN(n11157) );
  NAND2_X1 U14344 ( .A1(n11158), .A2(n11157), .ZN(n11159) );
  MUX2_X1 U14345 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B(n11159), .S(
        P2_STATE2_REG_0__SCAN_IN), .Z(n11163) );
  INV_X1 U14346 ( .A(n11163), .ZN(n11160) );
  OAI21_X1 U14347 ( .B1(n11160), .B2(n17526), .A(n17575), .ZN(n11164) );
  NAND2_X1 U14348 ( .A1(n17651), .A2(n17984), .ZN(n17453) );
  MUX2_X1 U14349 ( .A(n11165), .B(n11164), .S(n17453), .Z(n11208) );
  NAND2_X1 U14350 ( .A1(n17986), .A2(n11166), .ZN(n11169) );
  NAND2_X1 U14351 ( .A1(n11167), .A2(n10734), .ZN(n11168) );
  NAND2_X1 U14352 ( .A1(n11168), .A2(n11188), .ZN(n11476) );
  NAND2_X1 U14353 ( .A1(n9710), .A2(n17575), .ZN(n11468) );
  AOI21_X1 U14354 ( .B1(n11468), .B2(n17667), .A(n11170), .ZN(n11172) );
  NAND4_X1 U14355 ( .A1(n11198), .A2(n11197), .A3(n11174), .A4(n11195), .ZN(
        n11176) );
  INV_X1 U14356 ( .A(n11175), .ZN(n11185) );
  NAND3_X1 U14357 ( .A1(n11173), .A2(n17654), .A3(n17658), .ZN(n11177) );
  INV_X1 U14358 ( .A(n11178), .ZN(n11179) );
  OAI21_X1 U14359 ( .B1(n11181), .B2(n11180), .A(n11179), .ZN(n11184) );
  INV_X1 U14360 ( .A(n11182), .ZN(n11183) );
  NAND2_X1 U14361 ( .A1(n11184), .A2(n11183), .ZN(n11186) );
  INV_X1 U14362 ( .A(n11188), .ZN(n11189) );
  NAND2_X1 U14363 ( .A1(n20927), .A2(n20921), .ZN(n13059) );
  INV_X1 U14364 ( .A(n17668), .ZN(n11201) );
  INV_X1 U14365 ( .A(n11190), .ZN(n11193) );
  INV_X1 U14366 ( .A(n11191), .ZN(n11192) );
  AND2_X1 U14367 ( .A1(n11192), .A2(n17989), .ZN(n17985) );
  NAND2_X1 U14368 ( .A1(n11193), .A2(n17985), .ZN(n11194) );
  INV_X1 U14369 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n18012) );
  NAND2_X1 U14370 ( .A1(n11194), .A2(n18012), .ZN(n20910) );
  AND4_X1 U14371 ( .A1(n11198), .A2(n11197), .A3(n11196), .A4(n11195), .ZN(
        n11199) );
  NOR2_X1 U14372 ( .A1(n12781), .A2(n11199), .ZN(n11200) );
  MUX2_X1 U14373 ( .A(n20910), .B(n11200), .S(n11386), .Z(n18013) );
  NAND3_X1 U14374 ( .A1(n11201), .A2(n18013), .A3(n17984), .ZN(n11206) );
  MUX2_X1 U14375 ( .A(n10720), .B(n11202), .S(n17984), .Z(n11204) );
  NAND2_X1 U14376 ( .A1(n17654), .A2(n17687), .ZN(n11203) );
  OR2_X1 U14377 ( .A1(n11204), .A2(n11203), .ZN(n11205) );
  NOR2_X1 U14378 ( .A1(n17668), .A2(n12958), .ZN(n20923) );
  NAND2_X1 U14379 ( .A1(n11209), .A2(n11210), .ZN(n12846) );
  NAND2_X1 U14380 ( .A1(n12779), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n11214) );
  NAND2_X1 U14381 ( .A1(n11212), .A2(n20750), .ZN(n12774) );
  INV_X2 U14382 ( .A(n12774), .ZN(n12768) );
  AOI22_X1 U14383 ( .A1(n11243), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n12768), 
        .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n11213) );
  NAND2_X1 U14384 ( .A1(n11223), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n11219) );
  NAND2_X1 U14385 ( .A1(n17984), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n11218) );
  INV_X1 U14386 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n11215) );
  NAND3_X1 U14387 ( .A1(n11219), .A2(n11218), .A3(n11217), .ZN(n13541) );
  NAND2_X1 U14388 ( .A1(n14026), .A2(n11011), .ZN(n11229) );
  NAND2_X1 U14389 ( .A1(n11370), .A2(n11499), .ZN(n11222) );
  NAND2_X1 U14390 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n11220) );
  AND2_X1 U14391 ( .A1(n12775), .A2(n11220), .ZN(n11221) );
  OR2_X1 U14392 ( .A1(n11227), .A2(n12774), .ZN(n11236) );
  NAND3_X1 U14393 ( .A1(n11222), .A2(n11221), .A3(n11236), .ZN(n13540) );
  NAND2_X1 U14394 ( .A1(n13541), .A2(n13540), .ZN(n13539) );
  INV_X1 U14395 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n11224) );
  INV_X1 U14396 ( .A(n11225), .ZN(n11226) );
  XNOR2_X1 U14397 ( .A(n13539), .B(n11233), .ZN(n14059) );
  NAND2_X1 U14398 ( .A1(n11227), .A2(n10734), .ZN(n11228) );
  MUX2_X1 U14399 ( .A(n11228), .B(n20909), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n11232) );
  INV_X1 U14400 ( .A(n11500), .ZN(n11230) );
  OR2_X1 U14401 ( .A1(n9702), .A2(n11230), .ZN(n11231) );
  AND2_X1 U14402 ( .A1(n11232), .A2(n11231), .ZN(n14058) );
  INV_X1 U14403 ( .A(n11233), .ZN(n11234) );
  NAND2_X1 U14404 ( .A1(n13539), .A2(n11234), .ZN(n11235) );
  NAND2_X1 U14405 ( .A1(n14061), .A2(n11235), .ZN(n11241) );
  OR2_X1 U14406 ( .A1(n9702), .A2(n11504), .ZN(n11237) );
  OAI211_X1 U14407 ( .C1(n20750), .C2(n20900), .A(n11237), .B(n11236), .ZN(
        n11239) );
  XNOR2_X1 U14408 ( .A(n11241), .B(n11239), .ZN(n14350) );
  INV_X1 U14409 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n21726) );
  INV_X1 U14410 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n20295) );
  OAI22_X1 U14411 ( .A1(n12775), .A2(n21726), .B1(n12774), .B2(n20295), .ZN(
        n11238) );
  AOI21_X1 U14412 ( .B1(n12779), .B2(P2_REIP_REG_2__SCAN_IN), .A(n11238), .ZN(
        n14349) );
  INV_X1 U14413 ( .A(n11239), .ZN(n11240) );
  NAND2_X1 U14414 ( .A1(n11241), .A2(n11240), .ZN(n11242) );
  NAND2_X1 U14415 ( .A1(n12779), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n11249) );
  AOI22_X1 U14416 ( .A1(n12768), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n11245) );
  NAND2_X1 U14417 ( .A1(n11243), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n11244) );
  AND2_X1 U14418 ( .A1(n11245), .A2(n11244), .ZN(n11248) );
  INV_X1 U14419 ( .A(n11229), .ZN(n11370) );
  NAND2_X1 U14420 ( .A1(n11370), .A2(n11246), .ZN(n11247) );
  AND3_X1 U14421 ( .A1(n11249), .A2(n11248), .A3(n11247), .ZN(n14562) );
  NAND2_X1 U14422 ( .A1(n12779), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n11254) );
  AOI22_X1 U14423 ( .A1(n11243), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n12768), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n11253) );
  OR2_X1 U14424 ( .A1(n9702), .A2(n10914), .ZN(n11252) );
  NAND2_X1 U14425 ( .A1(n12779), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n11259) );
  AOI22_X1 U14426 ( .A1(n11243), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n12768), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n11258) );
  NAND2_X1 U14427 ( .A1(n11370), .A2(n11256), .ZN(n11257) );
  INV_X1 U14428 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n20835) );
  AOI22_X1 U14429 ( .A1(n11243), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n12768), .B2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n11262) );
  OAI21_X1 U14430 ( .B1(n11261), .B2(n20835), .A(n11262), .ZN(n14049) );
  NAND2_X1 U14431 ( .A1(n14048), .A2(n14049), .ZN(n11265) );
  INV_X1 U14432 ( .A(n13022), .ZN(n11263) );
  NAND2_X1 U14433 ( .A1(n14026), .A2(n11263), .ZN(n11264) );
  INV_X1 U14434 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n20837) );
  AOI22_X1 U14435 ( .A1(n11243), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n12768), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n11266) );
  OAI21_X1 U14436 ( .B1(n11261), .B2(n20837), .A(n11266), .ZN(n14083) );
  NAND2_X1 U14437 ( .A1(n12779), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n11279) );
  AOI22_X1 U14438 ( .A1(n11243), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n12768), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n11278) );
  AOI22_X1 U14439 ( .A1(n11190), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n16411), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11270) );
  AOI22_X1 U14440 ( .A1(n10841), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10891), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11269) );
  AOI22_X1 U14441 ( .A1(n16466), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n16464), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11268) );
  AOI22_X1 U14442 ( .A1(n10842), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n16465), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11267) );
  NAND4_X1 U14443 ( .A1(n11270), .A2(n11269), .A3(n11268), .A4(n11267), .ZN(
        n11276) );
  AOI22_X1 U14444 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n16472), .B1(
        n16471), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11274) );
  AOI22_X1 U14445 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n17505), .B1(
        n16473), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11273) );
  AOI22_X1 U14446 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n10848), .B1(
        n16437), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11272) );
  AOI22_X1 U14447 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n10847), .B1(
        n16438), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11271) );
  NAND4_X1 U14448 ( .A1(n11274), .A2(n11273), .A3(n11272), .A4(n11271), .ZN(
        n11275) );
  OR2_X1 U14449 ( .A1(n9702), .A2(n16699), .ZN(n11277) );
  NAND2_X1 U14450 ( .A1(n12779), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n11293) );
  AOI22_X1 U14451 ( .A1(n11243), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n12768), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n11292) );
  AOI22_X1 U14452 ( .A1(n11190), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n16411), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11283) );
  AOI22_X1 U14453 ( .A1(n10841), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n16464), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11282) );
  AOI22_X1 U14454 ( .A1(n16466), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n16465), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11281) );
  AOI22_X1 U14455 ( .A1(n10842), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10891), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11280) );
  NAND4_X1 U14456 ( .A1(n11283), .A2(n11282), .A3(n11281), .A4(n11280), .ZN(
        n11289) );
  AOI22_X1 U14457 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n16472), .B1(
        n16471), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11287) );
  AOI22_X1 U14458 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n17505), .B1(
        n16473), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11286) );
  AOI22_X1 U14459 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n10848), .B1(
        n16437), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11285) );
  AOI22_X1 U14460 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n10847), .B1(
        n16438), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11284) );
  NAND4_X1 U14461 ( .A1(n11287), .A2(n11286), .A3(n11285), .A4(n11284), .ZN(
        n11288) );
  INV_X1 U14462 ( .A(n16731), .ZN(n11290) );
  OR2_X1 U14463 ( .A1(n9702), .A2(n11290), .ZN(n11291) );
  NAND2_X1 U14464 ( .A1(n12779), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n11306) );
  AOI22_X1 U14465 ( .A1(n11243), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n12768), 
        .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n11305) );
  AOI22_X1 U14466 ( .A1(n11190), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n16411), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11297) );
  AOI22_X1 U14467 ( .A1(n10841), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n16464), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11296) );
  AOI22_X1 U14468 ( .A1(n16466), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n16465), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11295) );
  AOI22_X1 U14469 ( .A1(n10842), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10891), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11294) );
  NAND4_X1 U14470 ( .A1(n11297), .A2(n11296), .A3(n11295), .A4(n11294), .ZN(
        n11303) );
  AOI22_X1 U14471 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n16472), .B1(
        n16471), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11301) );
  AOI22_X1 U14472 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n17505), .B1(
        n16473), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11300) );
  AOI22_X1 U14473 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n10848), .B1(
        n16437), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11299) );
  AOI22_X1 U14474 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n10847), .B1(
        n16438), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11298) );
  NAND4_X1 U14475 ( .A1(n11301), .A2(n11300), .A3(n11299), .A4(n11298), .ZN(
        n11302) );
  OR2_X1 U14476 ( .A1(n9702), .A2(n16724), .ZN(n11304) );
  INV_X1 U14477 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n11424) );
  AOI22_X1 U14478 ( .A1(n11243), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n12768), 
        .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n11319) );
  AOI22_X1 U14479 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n16466), .B1(
        n10841), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11310) );
  AOI22_X1 U14480 ( .A1(n11190), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n16464), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11309) );
  AOI22_X1 U14481 ( .A1(n10842), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n16465), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11308) );
  AOI22_X1 U14482 ( .A1(n16411), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10891), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11307) );
  NAND4_X1 U14483 ( .A1(n11310), .A2(n11309), .A3(n11308), .A4(n11307), .ZN(
        n11316) );
  AOI22_X1 U14484 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n16472), .B1(
        n16471), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11314) );
  AOI22_X1 U14485 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n17505), .B1(
        n16473), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11313) );
  AOI22_X1 U14486 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n10848), .B1(
        n16437), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11312) );
  AOI22_X1 U14487 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n10847), .B1(
        n16438), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11311) );
  NAND4_X1 U14488 ( .A1(n11314), .A2(n11313), .A3(n11312), .A4(n11311), .ZN(
        n11315) );
  INV_X1 U14489 ( .A(n16719), .ZN(n11317) );
  OR2_X1 U14490 ( .A1(n9702), .A2(n11317), .ZN(n11318) );
  OAI211_X1 U14491 ( .C1(n11261), .C2(n11424), .A(n11319), .B(n11318), .ZN(
        n13527) );
  NAND2_X1 U14492 ( .A1(n12779), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n11332) );
  AOI22_X1 U14493 ( .A1(n11243), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n12768), 
        .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n11331) );
  AOI22_X1 U14494 ( .A1(n11190), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n16411), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11323) );
  AOI22_X1 U14495 ( .A1(n10841), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n16464), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11322) );
  AOI22_X1 U14496 ( .A1(n16466), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n16465), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11321) );
  AOI22_X1 U14497 ( .A1(n10842), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10891), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11320) );
  NAND4_X1 U14498 ( .A1(n11323), .A2(n11322), .A3(n11321), .A4(n11320), .ZN(
        n11329) );
  AOI22_X1 U14499 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n16472), .B1(
        n16471), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11327) );
  AOI22_X1 U14500 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n17505), .B1(
        n16473), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11326) );
  AOI22_X1 U14501 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n10848), .B1(
        n16437), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11325) );
  AOI22_X1 U14502 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n10847), .B1(
        n16438), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11324) );
  NAND4_X1 U14503 ( .A1(n11327), .A2(n11326), .A3(n11325), .A4(n11324), .ZN(
        n11328) );
  OR2_X1 U14504 ( .A1(n11329), .A2(n11328), .ZN(n16359) );
  OR2_X1 U14505 ( .A1(n9702), .A2(n16715), .ZN(n11330) );
  NAND2_X1 U14506 ( .A1(n12779), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n11347) );
  AOI22_X1 U14507 ( .A1(n11243), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n12768), 
        .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n11346) );
  AOI22_X1 U14508 ( .A1(n11190), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n16411), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11337) );
  AOI22_X1 U14509 ( .A1(n10841), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n16464), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11336) );
  AOI22_X1 U14510 ( .A1(n16466), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n16465), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11335) );
  AOI22_X1 U14511 ( .A1(n10842), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10891), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11334) );
  NAND4_X1 U14512 ( .A1(n11337), .A2(n11336), .A3(n11335), .A4(n11334), .ZN(
        n11343) );
  AOI22_X1 U14513 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n16472), .B1(
        n16471), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11341) );
  AOI22_X1 U14514 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n17505), .B1(
        n16473), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11340) );
  AOI22_X1 U14515 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n10848), .B1(
        n16437), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11339) );
  AOI22_X1 U14516 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n10847), .B1(
        n16438), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11338) );
  NAND4_X1 U14517 ( .A1(n11341), .A2(n11340), .A3(n11339), .A4(n11338), .ZN(
        n11342) );
  INV_X1 U14518 ( .A(n16711), .ZN(n11344) );
  OR2_X1 U14519 ( .A1(n9702), .A2(n11344), .ZN(n11345) );
  INV_X1 U14520 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n20848) );
  AOI22_X1 U14521 ( .A1(n11243), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n12768), 
        .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n11359) );
  AOI22_X1 U14522 ( .A1(n11190), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n16411), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11351) );
  AOI22_X1 U14523 ( .A1(n10841), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n16464), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11350) );
  AOI22_X1 U14524 ( .A1(n16466), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n16465), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11349) );
  AOI22_X1 U14525 ( .A1(n10842), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10891), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11348) );
  NAND4_X1 U14526 ( .A1(n11351), .A2(n11350), .A3(n11349), .A4(n11348), .ZN(
        n11357) );
  AOI22_X1 U14527 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n16472), .B1(
        n16471), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11355) );
  AOI22_X1 U14528 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n16473), .B1(
        n17505), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11354) );
  AOI22_X1 U14529 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n10848), .B1(
        n16437), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11353) );
  AOI22_X1 U14530 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n10847), .B1(
        n16438), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11352) );
  NAND4_X1 U14531 ( .A1(n11355), .A2(n11354), .A3(n11353), .A4(n11352), .ZN(
        n11356) );
  OR2_X1 U14532 ( .A1(n11357), .A2(n11356), .ZN(n16360) );
  INV_X1 U14533 ( .A(n16360), .ZN(n16706) );
  OR2_X1 U14534 ( .A1(n9702), .A2(n16706), .ZN(n11358) );
  OAI211_X1 U14535 ( .C1(n11261), .C2(n20848), .A(n11359), .B(n11358), .ZN(
        n14752) );
  NAND2_X1 U14536 ( .A1(n12779), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n11373) );
  AOI22_X1 U14537 ( .A1(n11243), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n12768), 
        .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n11372) );
  AOI22_X1 U14538 ( .A1(n11190), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n16411), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11363) );
  AOI22_X1 U14539 ( .A1(n10841), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n16464), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11362) );
  AOI22_X1 U14540 ( .A1(n16466), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n16465), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11361) );
  AOI22_X1 U14541 ( .A1(n10842), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10891), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11360) );
  NAND4_X1 U14542 ( .A1(n11363), .A2(n11362), .A3(n11361), .A4(n11360), .ZN(
        n11369) );
  AOI22_X1 U14543 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n16472), .B1(
        n16471), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11367) );
  AOI22_X1 U14544 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n17505), .B1(
        n16473), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11366) );
  AOI22_X1 U14545 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n10848), .B1(
        n16437), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11365) );
  AOI22_X1 U14546 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n10847), .B1(
        n16438), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11364) );
  NAND4_X1 U14547 ( .A1(n11367), .A2(n11366), .A3(n11365), .A4(n11364), .ZN(
        n11368) );
  OR2_X1 U14548 ( .A1(n11369), .A2(n11368), .ZN(n16700) );
  NAND2_X1 U14549 ( .A1(n11370), .A2(n16700), .ZN(n11371) );
  NAND2_X1 U14550 ( .A1(n12779), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n11375) );
  AOI22_X1 U14551 ( .A1(n11243), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n12768), 
        .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n11374) );
  INV_X1 U14552 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n20853) );
  AOI22_X1 U14553 ( .A1(n11243), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n12768), 
        .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n11377) );
  OAI21_X1 U14554 ( .B1(n11261), .B2(n20853), .A(n11377), .ZN(n16142) );
  INV_X1 U14555 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n20855) );
  AOI22_X1 U14556 ( .A1(n11243), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n12768), 
        .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n11378) );
  OAI21_X1 U14557 ( .B1(n11261), .B2(n20855), .A(n11378), .ZN(n16126) );
  NAND2_X1 U14558 ( .A1(n12779), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n11380) );
  AOI22_X1 U14559 ( .A1(n11243), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n12768), 
        .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n11379) );
  NAND2_X1 U14560 ( .A1(n12779), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n11382) );
  AOI22_X1 U14561 ( .A1(n11243), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n12768), 
        .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n11381) );
  AOI21_X1 U14562 ( .B1(n11384), .B2(n16100), .A(n12763), .ZN(n16813) );
  OR2_X1 U14563 ( .A1(n11385), .A2(n10357), .ZN(n11391) );
  INV_X1 U14564 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n20859) );
  NAND2_X1 U14565 ( .A1(n12833), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n11388) );
  NAND2_X1 U14566 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n11387) );
  OAI211_X1 U14567 ( .C1(n12821), .C2(n20859), .A(n11388), .B(n11387), .ZN(
        n11389) );
  INV_X1 U14568 ( .A(n11389), .ZN(n11390) );
  INV_X1 U14569 ( .A(n11392), .ZN(n11393) );
  INV_X1 U14570 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n11396) );
  OR2_X1 U14571 ( .A1(n12843), .A2(n14292), .ZN(n11395) );
  NAND2_X1 U14572 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n11394) );
  OAI211_X1 U14573 ( .C1(n12821), .C2(n11396), .A(n11395), .B(n11394), .ZN(
        n11397) );
  AOI21_X1 U14574 ( .B1(n12840), .B2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A(
        n11397), .ZN(n14289) );
  OR2_X1 U14575 ( .A1(n11385), .A2(n17436), .ZN(n11402) );
  INV_X1 U14576 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n16300) );
  NAND2_X1 U14577 ( .A1(n12833), .A2(P2_EBX_REG_5__SCAN_IN), .ZN(n11399) );
  NAND2_X1 U14578 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11398) );
  OAI211_X1 U14579 ( .C1(n12821), .C2(n16300), .A(n11399), .B(n11398), .ZN(
        n11400) );
  INV_X1 U14580 ( .A(n11400), .ZN(n11401) );
  NAND2_X1 U14581 ( .A1(n11402), .A2(n11401), .ZN(n14341) );
  NAND2_X1 U14582 ( .A1(n14288), .A2(n14341), .ZN(n14340) );
  INV_X1 U14583 ( .A(n14340), .ZN(n11407) );
  NAND2_X1 U14584 ( .A1(n12833), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n11404) );
  NAND2_X1 U14585 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11403) );
  OAI211_X1 U14586 ( .C1(n12821), .C2(n20835), .A(n11404), .B(n11403), .ZN(
        n11405) );
  AOI21_X1 U14587 ( .B1(n12840), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n11405), .ZN(n14510) );
  INV_X1 U14588 ( .A(n14510), .ZN(n11406) );
  NAND2_X1 U14589 ( .A1(n11407), .A2(n11406), .ZN(n14509) );
  NAND2_X1 U14590 ( .A1(n12833), .A2(P2_EBX_REG_7__SCAN_IN), .ZN(n11409) );
  NAND2_X1 U14591 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n11408) );
  OAI211_X1 U14592 ( .C1(n12821), .C2(n20837), .A(n11409), .B(n11408), .ZN(
        n11410) );
  AOI21_X1 U14593 ( .B1(n12840), .B2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n11410), .ZN(n14519) );
  INV_X1 U14594 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n20839) );
  NAND2_X1 U14595 ( .A1(n12833), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n11413) );
  NAND2_X1 U14596 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n11412) );
  OAI211_X1 U14597 ( .C1(n12821), .C2(n20839), .A(n11413), .B(n11412), .ZN(
        n11414) );
  AOI21_X1 U14598 ( .B1(n12840), .B2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A(
        n11414), .ZN(n16267) );
  OR2_X1 U14599 ( .A1(n11385), .A2(n10240), .ZN(n11419) );
  INV_X1 U14600 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n20841) );
  NAND2_X1 U14601 ( .A1(n12833), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n11416) );
  NAND2_X1 U14602 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n11415) );
  OAI211_X1 U14603 ( .C1(n12821), .C2(n20841), .A(n11416), .B(n11415), .ZN(
        n11417) );
  INV_X1 U14604 ( .A(n11417), .ZN(n11418) );
  NAND2_X1 U14605 ( .A1(n11419), .A2(n11418), .ZN(n16252) );
  OR2_X1 U14606 ( .A1(n11385), .A2(n17385), .ZN(n11421) );
  AOI22_X1 U14607 ( .A1(n10772), .A2(P2_REIP_REG_10__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), 
        .ZN(n11420) );
  OAI211_X1 U14608 ( .C1(n16726), .C2(n12843), .A(n11421), .B(n11420), .ZN(
        n16239) );
  NAND2_X1 U14609 ( .A1(n16238), .A2(n16239), .ZN(n13531) );
  NAND2_X1 U14610 ( .A1(n12833), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n11423) );
  NAND2_X1 U14611 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n11422) );
  OAI211_X1 U14612 ( .C1(n12821), .C2(n11424), .A(n11423), .B(n11422), .ZN(
        n11425) );
  AOI21_X1 U14613 ( .B1(n12840), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n11425), .ZN(n13532) );
  INV_X1 U14614 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n16227) );
  NAND2_X1 U14615 ( .A1(n12833), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n11428) );
  NAND2_X1 U14616 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n11427) );
  OAI211_X1 U14617 ( .C1(n12821), .C2(n16227), .A(n11428), .B(n11427), .ZN(
        n11429) );
  AOI21_X1 U14618 ( .B1(n12840), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n11429), .ZN(n16222) );
  OR2_X1 U14619 ( .A1(n11385), .A2(n17348), .ZN(n11434) );
  INV_X1 U14620 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n20846) );
  NAND2_X1 U14621 ( .A1(n12833), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n11431) );
  NAND2_X1 U14622 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n11430) );
  OAI211_X1 U14623 ( .C1(n12821), .C2(n20846), .A(n11431), .B(n11430), .ZN(
        n11432) );
  INV_X1 U14624 ( .A(n11432), .ZN(n11433) );
  NAND2_X1 U14625 ( .A1(n11434), .A2(n11433), .ZN(n16203) );
  INV_X1 U14626 ( .A(n16191), .ZN(n11439) );
  NAND2_X1 U14627 ( .A1(n12833), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n11436) );
  NAND2_X1 U14628 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n11435) );
  OAI211_X1 U14629 ( .C1(n12821), .C2(n20848), .A(n11436), .B(n11435), .ZN(
        n11437) );
  AOI21_X1 U14630 ( .B1(n12840), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n11437), .ZN(n16192) );
  INV_X1 U14631 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n20849) );
  NAND2_X1 U14632 ( .A1(n12833), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n11441) );
  NAND2_X1 U14633 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n11440) );
  OAI211_X1 U14634 ( .C1(n12821), .C2(n20849), .A(n11441), .B(n11440), .ZN(
        n11442) );
  AOI21_X1 U14635 ( .B1(n12840), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n11442), .ZN(n16182) );
  INV_X1 U14636 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n20851) );
  NAND2_X1 U14637 ( .A1(n12833), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n11445) );
  NAND2_X1 U14638 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n11444) );
  OAI211_X1 U14639 ( .C1(n12821), .C2(n20851), .A(n11445), .B(n11444), .ZN(
        n11446) );
  AOI21_X1 U14640 ( .B1(n12840), .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n11446), .ZN(n16161) );
  OR2_X1 U14641 ( .A1(n11385), .A2(n17292), .ZN(n11451) );
  NAND2_X1 U14642 ( .A1(n12833), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n11448) );
  NAND2_X1 U14643 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n11447) );
  OAI211_X1 U14644 ( .C1(n12821), .C2(n20853), .A(n11448), .B(n11447), .ZN(
        n11449) );
  INV_X1 U14645 ( .A(n11449), .ZN(n11450) );
  NAND2_X1 U14646 ( .A1(n11451), .A2(n11450), .ZN(n16153) );
  OR2_X1 U14647 ( .A1(n11385), .A2(n14775), .ZN(n11456) );
  NAND2_X1 U14648 ( .A1(n12833), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n11453) );
  NAND2_X1 U14649 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n11452) );
  OAI211_X1 U14650 ( .C1(n12821), .C2(n20855), .A(n11453), .B(n11452), .ZN(
        n11454) );
  INV_X1 U14651 ( .A(n11454), .ZN(n11455) );
  NAND2_X1 U14652 ( .A1(n11456), .A2(n11455), .ZN(n16135) );
  NAND2_X1 U14653 ( .A1(n16134), .A2(n16135), .ZN(n13501) );
  INV_X1 U14654 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n21778) );
  NAND2_X1 U14655 ( .A1(n12833), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n11458) );
  NAND2_X1 U14656 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n11457) );
  OAI211_X1 U14657 ( .C1(n12821), .C2(n21778), .A(n11458), .B(n11457), .ZN(
        n11459) );
  AOI21_X1 U14658 ( .B1(n12840), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n11459), .ZN(n13503) );
  OR2_X2 U14659 ( .A1(n13501), .A2(n13503), .ZN(n16102) );
  INV_X1 U14660 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n11462) );
  NAND2_X1 U14661 ( .A1(n12833), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n11461) );
  NAND2_X1 U14662 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n11460) );
  OAI211_X1 U14663 ( .C1(n12821), .C2(n11462), .A(n11461), .B(n11460), .ZN(
        n11463) );
  AOI21_X1 U14664 ( .B1(n12840), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n11463), .ZN(n16103) );
  INV_X1 U14665 ( .A(n16101), .ZN(n11464) );
  AOI21_X1 U14666 ( .B1(n9845), .B2(n11464), .A(n12811), .ZN(n16958) );
  INV_X1 U14667 ( .A(n16958), .ZN(n16675) );
  NAND2_X1 U14668 ( .A1(n17498), .A2(n9710), .ZN(n11466) );
  NAND2_X1 U14669 ( .A1(n11466), .A2(n11465), .ZN(n11467) );
  NOR3_X1 U14670 ( .A1(n11227), .A2(n11468), .A3(n11170), .ZN(n11469) );
  OAI21_X1 U14671 ( .B1(n10730), .B2(n11472), .A(n11471), .ZN(n11473) );
  INV_X1 U14672 ( .A(n11473), .ZN(n11474) );
  NAND2_X1 U14673 ( .A1(n11475), .A2(n11474), .ZN(n11483) );
  NAND2_X1 U14674 ( .A1(n17449), .A2(n11476), .ZN(n11477) );
  NAND2_X1 U14675 ( .A1(n11477), .A2(n10731), .ZN(n11481) );
  INV_X1 U14676 ( .A(n11471), .ZN(n15978) );
  AOI22_X1 U14677 ( .A1(n15978), .A2(n17575), .B1(n17564), .B2(n17526), .ZN(
        n11478) );
  AND2_X1 U14678 ( .A1(n11479), .A2(n11478), .ZN(n11480) );
  NAND2_X1 U14679 ( .A1(n11481), .A2(n11480), .ZN(n11482) );
  AOI21_X1 U14680 ( .B1(n11483), .B2(n10723), .A(n11482), .ZN(n17447) );
  NAND2_X1 U14681 ( .A1(n17447), .A2(n10730), .ZN(n11484) );
  AND2_X1 U14682 ( .A1(n11523), .A2(n11484), .ZN(n17294) );
  NAND3_X1 U14683 ( .A1(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n17274) );
  INV_X1 U14684 ( .A(n17274), .ZN(n14773) );
  NAND4_X1 U14685 ( .A1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A4(n14773), .ZN(n11522) );
  NOR2_X1 U14686 ( .A1(n11522), .A2(n10357), .ZN(n11485) );
  AND2_X1 U14687 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17328) );
  AND2_X1 U14688 ( .A1(n17328), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n14771) );
  NAND2_X1 U14689 ( .A1(n11485), .A2(n14771), .ZN(n11486) );
  NAND3_X1 U14690 ( .A1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n11519) );
  NAND3_X1 U14691 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n11492) );
  INV_X1 U14692 ( .A(n11492), .ZN(n17418) );
  AND2_X1 U14693 ( .A1(n15981), .A2(n20888), .ZN(n11487) );
  INV_X1 U14694 ( .A(n17136), .ZN(n18058) );
  OR2_X1 U14695 ( .A1(n11523), .A2(n18058), .ZN(n14051) );
  NAND2_X1 U14696 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n14052) );
  NAND2_X1 U14697 ( .A1(n20295), .A2(n14052), .ZN(n11490) );
  INV_X1 U14698 ( .A(n11490), .ZN(n20284) );
  NAND2_X1 U14699 ( .A1(n20275), .A2(n20284), .ZN(n20288) );
  NOR2_X1 U14700 ( .A1(n20295), .A2(n14052), .ZN(n11491) );
  INV_X1 U14701 ( .A(n11491), .ZN(n11488) );
  NAND2_X1 U14702 ( .A1(n17294), .A2(n11488), .ZN(n20285) );
  NAND3_X1 U14703 ( .A1(n14051), .A2(n20288), .A3(n20285), .ZN(n17435) );
  NOR2_X1 U14704 ( .A1(n10327), .A2(n17435), .ZN(n17417) );
  NAND2_X1 U14705 ( .A1(n17418), .A2(n17417), .ZN(n18076) );
  NAND2_X1 U14706 ( .A1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n17405) );
  NOR2_X1 U14707 ( .A1(n18076), .A2(n17405), .ZN(n17326) );
  INV_X1 U14708 ( .A(n17326), .ZN(n11489) );
  NAND2_X1 U14709 ( .A1(n17419), .A2(n14051), .ZN(n20257) );
  NAND2_X1 U14710 ( .A1(n11489), .A2(n20257), .ZN(n17371) );
  OAI21_X1 U14711 ( .B1(n17419), .B2(n17240), .A(n17371), .ZN(n17252) );
  NOR2_X1 U14712 ( .A1(n17136), .A2(n20859), .ZN(n16954) );
  INV_X1 U14713 ( .A(n11519), .ZN(n17325) );
  INV_X1 U14714 ( .A(n17405), .ZN(n11494) );
  OAI211_X1 U14715 ( .C1(n20275), .C2(n11491), .A(n11490), .B(n14774), .ZN(
        n18095) );
  NOR2_X1 U14716 ( .A1(n11492), .A2(n18095), .ZN(n17421) );
  NAND2_X1 U14717 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n17421), .ZN(
        n18075) );
  INV_X1 U14718 ( .A(n18075), .ZN(n11493) );
  NAND2_X1 U14719 ( .A1(n11494), .A2(n11493), .ZN(n17237) );
  NAND3_X1 U14720 ( .A1(n17313), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n14773), .ZN(n17263) );
  NOR4_X1 U14721 ( .A1(n17263), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        n17259), .A4(n11495), .ZN(n11496) );
  AOI211_X1 U14722 ( .C1(n17252), .C2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n16954), .B(n11496), .ZN(n11497) );
  OAI21_X1 U14723 ( .B1(n16675), .B2(n20259), .A(n11497), .ZN(n11524) );
  INV_X1 U14724 ( .A(n11498), .ZN(n13543) );
  NAND2_X1 U14725 ( .A1(n13543), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13542) );
  XNOR2_X1 U14726 ( .A(n11500), .B(n11499), .ZN(n11501) );
  NOR2_X1 U14727 ( .A1(n13542), .A2(n11501), .ZN(n11503) );
  AOI21_X1 U14728 ( .B1(n13542), .B2(n11501), .A(n11503), .ZN(n11502) );
  INV_X1 U14729 ( .A(n11502), .ZN(n13927) );
  NOR2_X1 U14730 ( .A1(n14054), .A2(n13927), .ZN(n13926) );
  NOR2_X1 U14731 ( .A1(n11503), .A2(n13926), .ZN(n11507) );
  XOR2_X1 U14732 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n11507), .Z(
        n17154) );
  INV_X1 U14733 ( .A(n17154), .ZN(n11506) );
  XNOR2_X1 U14734 ( .A(n11505), .B(n11504), .ZN(n17152) );
  NAND2_X1 U14735 ( .A1(n11506), .A2(n17152), .ZN(n20287) );
  OR2_X1 U14736 ( .A1(n11507), .A2(n20295), .ZN(n11508) );
  NAND2_X1 U14737 ( .A1(n20287), .A2(n11508), .ZN(n11509) );
  XNOR2_X1 U14738 ( .A(n11509), .B(n18096), .ZN(n17140) );
  NAND2_X1 U14739 ( .A1(n11509), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11510) );
  NAND2_X1 U14740 ( .A1(n11511), .A2(n10914), .ZN(n11512) );
  INV_X1 U14741 ( .A(n17109), .ZN(n11514) );
  NAND2_X1 U14742 ( .A1(n11514), .A2(n11516), .ZN(n11515) );
  INV_X1 U14743 ( .A(n17328), .ZN(n11520) );
  NOR2_X1 U14744 ( .A1(n11520), .A2(n11519), .ZN(n11521) );
  NAND2_X1 U14745 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n19192) );
  NAND3_X1 U14746 ( .A1(n17849), .A2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n18426) );
  NAND2_X1 U14747 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n19149) );
  NAND2_X1 U14748 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17811) );
  NAND2_X1 U14749 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n19101) );
  NOR2_X1 U14750 ( .A1(n18353), .A2(n19101), .ZN(n11532) );
  NAND2_X1 U14751 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n19055) );
  NAND2_X1 U14752 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n19021) );
  NAND2_X1 U14753 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n13560) );
  INV_X1 U14754 ( .A(n13560), .ZN(n11526) );
  XNOR2_X1 U14755 ( .A(n9842), .B(n10506), .ZN(n18211) );
  INV_X1 U14756 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n18220) );
  NAND2_X1 U14757 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n13400), .ZN(
        n13394) );
  AOI21_X1 U14758 ( .B1(n18220), .B2(n13394), .A(n9842), .ZN(n18219) );
  NAND2_X1 U14759 ( .A1(n17778), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n11531) );
  INV_X1 U14760 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n18243) );
  NOR2_X1 U14761 ( .A1(n11531), .A2(n18243), .ZN(n11528) );
  OAI21_X1 U14762 ( .B1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n11528), .A(
        n13394), .ZN(n13566) );
  INV_X1 U14763 ( .A(n13566), .ZN(n18233) );
  AND2_X1 U14764 ( .A1(n11531), .A2(n18243), .ZN(n11527) );
  NOR2_X1 U14765 ( .A1(n11528), .A2(n11527), .ZN(n18242) );
  NOR2_X1 U14766 ( .A1(n18562), .A2(n11529), .ZN(n11538) );
  INV_X1 U14767 ( .A(n11538), .ZN(n11530) );
  NOR2_X1 U14768 ( .A1(n19021), .A2(n11530), .ZN(n13562) );
  OAI21_X1 U14769 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n13562), .A(
        n11531), .ZN(n19005) );
  INV_X1 U14770 ( .A(n19005), .ZN(n18256) );
  NAND2_X1 U14771 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n11538), .ZN(
        n11540) );
  OAI21_X1 U14772 ( .B1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n11538), .A(
        n11540), .ZN(n17796) );
  INV_X1 U14773 ( .A(n17796), .ZN(n18278) );
  INV_X1 U14774 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n19071) );
  INV_X1 U14775 ( .A(n11532), .ZN(n19081) );
  NAND2_X1 U14776 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n11533), .ZN(
        n17808) );
  NOR2_X1 U14777 ( .A1(n19081), .A2(n17808), .ZN(n19051) );
  NAND2_X1 U14778 ( .A1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n19051), .ZN(
        n11537) );
  NOR2_X1 U14779 ( .A1(n19071), .A2(n11537), .ZN(n11534) );
  NAND2_X1 U14780 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n9816), .ZN(
        n17795) );
  OAI21_X1 U14781 ( .B1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n11534), .A(
        n17795), .ZN(n19058) );
  INV_X1 U14782 ( .A(n19058), .ZN(n18301) );
  OAI21_X1 U14783 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n19051), .A(
        n11537), .ZN(n19083) );
  INV_X1 U14784 ( .A(n19083), .ZN(n18321) );
  NOR2_X1 U14785 ( .A1(n18562), .A2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n18547) );
  INV_X1 U14786 ( .A(n18547), .ZN(n18522) );
  NOR2_X1 U14787 ( .A1(n17810), .A2(n18522), .ZN(n18378) );
  NAND2_X1 U14788 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n18378), .ZN(
        n18342) );
  NAND2_X1 U14789 ( .A1(n11536), .A2(n18342), .ZN(n18370) );
  NOR2_X1 U14790 ( .A1(n18321), .A2(n18330), .ZN(n18320) );
  NOR2_X1 U14791 ( .A1(n18320), .A2(n18518), .ZN(n18312) );
  XOR2_X1 U14792 ( .A(n19071), .B(n11537), .Z(n19066) );
  AOI21_X1 U14793 ( .B1(n10497), .B2(n17795), .A(n11538), .ZN(n19036) );
  INV_X1 U14794 ( .A(n19036), .ZN(n11539) );
  NAND2_X1 U14795 ( .A1(n18286), .A2(n11539), .ZN(n18287) );
  NOR2_X1 U14796 ( .A1(n18278), .A2(n18277), .ZN(n18276) );
  OR2_X1 U14797 ( .A1(n18276), .A2(n18518), .ZN(n18263) );
  INV_X1 U14798 ( .A(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n11541) );
  AOI21_X1 U14799 ( .B1(n11541), .B2(n11540), .A(n13562), .ZN(n19012) );
  INV_X1 U14800 ( .A(n19012), .ZN(n11542) );
  NAND2_X1 U14801 ( .A1(n18263), .A2(n11542), .ZN(n18264) );
  NOR2_X1 U14802 ( .A1(n18256), .A2(n18255), .ZN(n18254) );
  NOR2_X1 U14803 ( .A1(n18254), .A2(n18518), .ZN(n18241) );
  NOR2_X1 U14804 ( .A1(n18242), .A2(n18241), .ZN(n18240) );
  NOR2_X1 U14805 ( .A1(n18240), .A2(n18518), .ZN(n18232) );
  NOR2_X1 U14806 ( .A1(n18233), .A2(n18232), .ZN(n18231) );
  NOR2_X1 U14807 ( .A1(n18231), .A2(n18518), .ZN(n18218) );
  NOR3_X1 U14808 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .A3(P3_STATEBS16_REG_SCAN_IN), .ZN(n20055) );
  NAND2_X1 U14809 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n20055), .ZN(n18536) );
  INV_X1 U14810 ( .A(n18536), .ZN(n20050) );
  NAND2_X1 U14811 ( .A1(n10503), .A2(n20050), .ZN(n18559) );
  NOR3_X1 U14812 ( .A1(n18211), .A2(n18210), .A3(n18559), .ZN(n11732) );
  INV_X1 U14813 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n18189) );
  NAND2_X1 U14814 ( .A1(READY22_REG_SCAN_IN), .A2(READY2), .ZN(n20161) );
  INV_X1 U14815 ( .A(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11546) );
  AND2_X2 U14816 ( .A1(n14720), .A2(n11555), .ZN(n13270) );
  NAND2_X1 U14817 ( .A1(n13270), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n11545) );
  AND2_X2 U14818 ( .A1(n11558), .A2(n14720), .ZN(n11543) );
  NAND2_X1 U14819 ( .A1(n11543), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n11544) );
  OAI211_X1 U14820 ( .C1(n18735), .C2(n11546), .A(n11545), .B(n11544), .ZN(
        n11547) );
  INV_X1 U14821 ( .A(n11547), .ZN(n11553) );
  AND2_X4 U14822 ( .A1(n11549), .A2(n14338), .ZN(n18704) );
  AOI22_X1 U14823 ( .A1(n18704), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n18703), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11552) );
  AND2_X4 U14824 ( .A1(n11554), .A2(n11548), .ZN(n18706) );
  AND2_X4 U14825 ( .A1(n11548), .A2(n11555), .ZN(n18705) );
  AOI22_X1 U14826 ( .A1(n18706), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n18705), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11551) );
  NAND2_X1 U14827 ( .A1(n13795), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n11550) );
  NAND4_X1 U14828 ( .A1(n11553), .A2(n11552), .A3(n11551), .A4(n11550), .ZN(
        n11566) );
  INV_X2 U14829 ( .A(n14594), .ZN(n13878) );
  AOI22_X1 U14830 ( .A1(n13878), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n9703), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11564) );
  AOI22_X1 U14831 ( .A1(n13279), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n13278), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11563) );
  NAND2_X2 U14832 ( .A1(n11558), .A2(n14719), .ZN(n14593) );
  INV_X2 U14833 ( .A(n14591), .ZN(n14680) );
  AOI22_X1 U14834 ( .A1(n13718), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n14680), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11562) );
  INV_X2 U14835 ( .A(n11593), .ZN(n14649) );
  AOI22_X1 U14836 ( .A1(n14649), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n18739), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11561) );
  NAND4_X1 U14837 ( .A1(n11564), .A2(n11563), .A3(n11562), .A4(n11561), .ZN(
        n11565) );
  INV_X1 U14838 ( .A(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11569) );
  NAND2_X1 U14839 ( .A1(n11543), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11568) );
  NAND2_X1 U14840 ( .A1(n13270), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11567) );
  OAI211_X1 U14841 ( .C1(n18735), .C2(n11569), .A(n11568), .B(n11567), .ZN(
        n11570) );
  INV_X1 U14842 ( .A(n11570), .ZN(n11575) );
  OAI22_X1 U14843 ( .A1(n18728), .A2(n19624), .B1(n11594), .B2(n13701), .ZN(
        n11571) );
  INV_X1 U14844 ( .A(n11571), .ZN(n11574) );
  AOI22_X1 U14845 ( .A1(n18706), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n18705), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11573) );
  NAND2_X1 U14846 ( .A1(n13795), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11572) );
  NAND4_X1 U14847 ( .A1(n11575), .A2(n11574), .A3(n11573), .A4(n11572), .ZN(
        n11581) );
  AOI22_X1 U14848 ( .A1(n18703), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n14649), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11579) );
  AOI22_X1 U14849 ( .A1(n13279), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n13278), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11578) );
  AOI22_X1 U14850 ( .A1(n13718), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n14680), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11577) );
  AOI22_X1 U14851 ( .A1(n13878), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n18739), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11576) );
  NAND4_X1 U14852 ( .A1(n11579), .A2(n11578), .A3(n11577), .A4(n11576), .ZN(
        n11580) );
  NAND2_X1 U14853 ( .A1(n19565), .A2(n20150), .ZN(n13352) );
  INV_X1 U14854 ( .A(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11584) );
  NAND2_X1 U14855 ( .A1(n13270), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n11583) );
  NAND2_X1 U14856 ( .A1(n13878), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n11582) );
  OAI211_X1 U14857 ( .C1(n18735), .C2(n11584), .A(n11583), .B(n11582), .ZN(
        n11585) );
  INV_X1 U14858 ( .A(n11585), .ZN(n11592) );
  INV_X1 U14859 ( .A(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11587) );
  INV_X1 U14860 ( .A(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11586) );
  OAI22_X1 U14861 ( .A1(n13229), .A2(n11587), .B1(n14593), .B2(n11586), .ZN(
        n11588) );
  INV_X1 U14862 ( .A(n11588), .ZN(n11591) );
  AOI22_X1 U14863 ( .A1(n18706), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n18705), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11590) );
  NAND2_X1 U14864 ( .A1(n18704), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n11589) );
  NAND4_X1 U14865 ( .A1(n11592), .A2(n11591), .A3(n11590), .A4(n11589), .ZN(
        n11600) );
  AOI22_X1 U14866 ( .A1(n18736), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n18740), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11598) );
  AOI22_X1 U14867 ( .A1(n9683), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(n9703), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11597) );
  AOI22_X1 U14868 ( .A1(n13279), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n13278), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11596) );
  INV_X2 U14869 ( .A(n14591), .ZN(n18737) );
  AOI22_X1 U14870 ( .A1(n18737), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n18739), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11595) );
  NAND4_X1 U14871 ( .A1(n11598), .A2(n11597), .A3(n11596), .A4(n11595), .ZN(
        n11599) );
  INV_X1 U14872 ( .A(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11603) );
  NAND2_X1 U14873 ( .A1(n13270), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n11602) );
  NAND2_X1 U14874 ( .A1(n18739), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n11601) );
  OAI211_X1 U14875 ( .C1(n18735), .C2(n11603), .A(n11602), .B(n11601), .ZN(
        n11604) );
  INV_X1 U14876 ( .A(n11604), .ZN(n11608) );
  AOI22_X1 U14877 ( .A1(n13795), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n14649), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11607) );
  INV_X1 U14878 ( .A(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n17710) );
  AOI22_X1 U14879 ( .A1(n18706), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n18705), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11606) );
  NAND2_X1 U14880 ( .A1(n18704), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n11605) );
  NAND4_X1 U14881 ( .A1(n11608), .A2(n11607), .A3(n11606), .A4(n11605), .ZN(
        n11614) );
  INV_X1 U14882 ( .A(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n17708) );
  AOI22_X1 U14883 ( .A1(n13718), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n9683), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11612) );
  AOI22_X1 U14884 ( .A1(n11543), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9703), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11611) );
  AOI22_X1 U14885 ( .A1(n13279), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n13278), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11610) );
  AOI22_X1 U14886 ( .A1(n13878), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n18737), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11609) );
  NAND4_X1 U14887 ( .A1(n11612), .A2(n11611), .A3(n11610), .A4(n11609), .ZN(
        n11613) );
  INV_X1 U14888 ( .A(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n21760) );
  INV_X2 U14889 ( .A(n14335), .ZN(n18732) );
  NAND2_X1 U14890 ( .A1(n18732), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n11616) );
  NAND2_X1 U14891 ( .A1(n9683), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n11615) );
  OAI211_X1 U14892 ( .C1(n18735), .C2(n21760), .A(n11616), .B(n11615), .ZN(
        n11617) );
  INV_X1 U14893 ( .A(n11617), .ZN(n11621) );
  AOI22_X1 U14894 ( .A1(n18704), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n14649), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11620) );
  AOI22_X1 U14895 ( .A1(n18706), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n13279), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11619) );
  NAND2_X1 U14896 ( .A1(n13795), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n11618) );
  NAND4_X1 U14897 ( .A1(n11621), .A2(n11620), .A3(n11619), .A4(n11618), .ZN(
        n11627) );
  AOI22_X1 U14898 ( .A1(n11543), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9703), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11625) );
  INV_X1 U14899 ( .A(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n21852) );
  INV_X1 U14900 ( .A(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n14671) );
  AOI22_X1 U14901 ( .A1(n18705), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n13278), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11624) );
  AOI22_X1 U14902 ( .A1(n13878), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n18737), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11623) );
  INV_X2 U14903 ( .A(n14593), .ZN(n18738) );
  AOI22_X1 U14904 ( .A1(n18738), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n18739), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11622) );
  NAND4_X1 U14905 ( .A1(n11625), .A2(n11624), .A3(n11623), .A4(n11622), .ZN(
        n11626) );
  NOR2_X1 U14906 ( .A1(n11677), .A2(n11712), .ZN(n11656) );
  INV_X1 U14907 ( .A(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11630) );
  NAND2_X1 U14908 ( .A1(n9703), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n11629) );
  NAND2_X1 U14909 ( .A1(n13270), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n11628) );
  OAI211_X1 U14910 ( .C1(n18735), .C2(n11630), .A(n11629), .B(n11628), .ZN(
        n11631) );
  INV_X1 U14911 ( .A(n11631), .ZN(n11635) );
  AOI22_X1 U14912 ( .A1(n18704), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n18703), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11634) );
  AOI22_X1 U14913 ( .A1(n18706), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n18705), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11633) );
  NAND2_X1 U14914 ( .A1(n13795), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n11632) );
  NAND4_X1 U14915 ( .A1(n11635), .A2(n11634), .A3(n11633), .A4(n11632), .ZN(
        n11641) );
  AOI22_X1 U14916 ( .A1(n11543), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13878), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11639) );
  INV_X1 U14917 ( .A(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n14601) );
  AOI22_X1 U14918 ( .A1(n13279), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n13278), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11638) );
  AOI22_X1 U14919 ( .A1(n13718), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n14680), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11637) );
  AOI22_X1 U14920 ( .A1(n14649), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n18739), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11636) );
  NAND4_X1 U14921 ( .A1(n11639), .A2(n11638), .A3(n11637), .A4(n11636), .ZN(
        n11640) );
  INV_X1 U14922 ( .A(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11644) );
  NAND2_X1 U14923 ( .A1(n9704), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n11643) );
  NAND2_X1 U14924 ( .A1(n13270), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n11642) );
  OAI211_X1 U14925 ( .C1(n18735), .C2(n11644), .A(n11643), .B(n11642), .ZN(
        n11645) );
  INV_X1 U14926 ( .A(n11645), .ZN(n11649) );
  AOI22_X1 U14927 ( .A1(n18704), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n9683), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11648) );
  INV_X1 U14928 ( .A(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n21670) );
  AOI22_X1 U14929 ( .A1(n18706), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n18705), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11647) );
  NAND2_X1 U14930 ( .A1(n13795), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n11646) );
  NAND4_X1 U14931 ( .A1(n11649), .A2(n11648), .A3(n11647), .A4(n11646), .ZN(
        n11655) );
  AOI22_X1 U14932 ( .A1(n11543), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n13878), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11653) );
  AOI22_X1 U14933 ( .A1(n13279), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n13278), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11652) );
  AOI22_X1 U14934 ( .A1(n14649), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n18739), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11651) );
  AOI22_X1 U14935 ( .A1(n13718), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n18737), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11650) );
  NAND4_X1 U14936 ( .A1(n11653), .A2(n11652), .A3(n11651), .A4(n11650), .ZN(
        n11654) );
  NAND4_X1 U14937 ( .A1(n11678), .A2(n11656), .A3(n19574), .A4(n18787), .ZN(
        n13355) );
  INV_X1 U14938 ( .A(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11659) );
  NAND2_X1 U14939 ( .A1(n11543), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n11658) );
  INV_X1 U14940 ( .A(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n18721) );
  NAND2_X1 U14941 ( .A1(n18732), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n11657) );
  OAI211_X1 U14942 ( .C1(n18735), .C2(n11659), .A(n11658), .B(n11657), .ZN(
        n11660) );
  INV_X1 U14943 ( .A(n11660), .ZN(n11664) );
  AOI22_X1 U14944 ( .A1(n18704), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n13878), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11663) );
  AOI22_X1 U14945 ( .A1(n18706), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n18705), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11662) );
  NAND2_X1 U14946 ( .A1(n13795), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n11661) );
  NAND4_X1 U14947 ( .A1(n11664), .A2(n11663), .A3(n11662), .A4(n11661), .ZN(
        n11670) );
  AOI22_X1 U14948 ( .A1(n18703), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n14649), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11668) );
  AOI22_X1 U14949 ( .A1(n13718), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n9703), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11667) );
  AOI22_X1 U14950 ( .A1(n13279), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n13278), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11666) );
  INV_X1 U14951 ( .A(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n18725) );
  AOI22_X1 U14952 ( .A1(n18737), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n18739), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11665) );
  NAND4_X1 U14953 ( .A1(n11668), .A2(n11667), .A3(n11666), .A4(n11665), .ZN(
        n11669) );
  NAND2_X1 U14954 ( .A1(n13979), .A2(n13963), .ZN(n18185) );
  NAND2_X1 U14955 ( .A1(n13339), .A2(n19571), .ZN(n11672) );
  NAND2_X1 U14956 ( .A1(n20150), .A2(n11712), .ZN(n13691) );
  NOR2_X1 U14957 ( .A1(n20150), .A2(n11712), .ZN(n14155) );
  INV_X1 U14958 ( .A(n13339), .ZN(n11673) );
  NOR2_X1 U14959 ( .A1(n13963), .A2(n11687), .ZN(n14311) );
  NAND2_X1 U14960 ( .A1(n11673), .A2(n14311), .ZN(n13690) );
  NOR2_X1 U14961 ( .A1(n13690), .A2(n19588), .ZN(n11674) );
  INV_X1 U14962 ( .A(n14310), .ZN(n11675) );
  OAI211_X1 U14963 ( .C1(n19583), .C2(n13966), .A(n11675), .B(n19565), .ZN(
        n11683) );
  NAND2_X1 U14964 ( .A1(n19565), .A2(n18787), .ZN(n11676) );
  AOI22_X1 U14965 ( .A1(n14714), .A2(n19577), .B1(n11676), .B2(n19574), .ZN(
        n11682) );
  OAI21_X1 U14966 ( .B1(n11678), .B2(n19588), .A(n11677), .ZN(n11681) );
  NAND2_X1 U14967 ( .A1(n13352), .A2(n19571), .ZN(n13338) );
  INV_X1 U14968 ( .A(n11678), .ZN(n11679) );
  NAND2_X1 U14969 ( .A1(n13338), .A2(n11679), .ZN(n11680) );
  NAND4_X1 U14970 ( .A1(n11683), .A2(n11682), .A3(n11681), .A4(n11680), .ZN(
        n13968) );
  INV_X1 U14971 ( .A(n13968), .ZN(n11690) );
  INV_X1 U14972 ( .A(n13351), .ZN(n11685) );
  NAND2_X1 U14973 ( .A1(n13340), .A2(n18787), .ZN(n11684) );
  NAND2_X1 U14974 ( .A1(n11685), .A2(n11684), .ZN(n13969) );
  NAND2_X1 U14975 ( .A1(n11686), .A2(n13969), .ZN(n11688) );
  NAND2_X1 U14976 ( .A1(n11688), .A2(n11687), .ZN(n11689) );
  MUX2_X1 U14977 ( .A(n11693), .B(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n13345) );
  NAND2_X1 U14978 ( .A1(n13345), .A2(n13332), .ZN(n11695) );
  NAND2_X1 U14979 ( .A1(n11693), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11694) );
  NAND2_X1 U14980 ( .A1(n11695), .A2(n11694), .ZN(n11704) );
  MUX2_X1 U14981 ( .A(n11696), .B(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .S(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n11703) );
  NAND2_X1 U14982 ( .A1(n11704), .A2(n11703), .ZN(n11698) );
  NAND2_X1 U14983 ( .A1(n11696), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11697) );
  NAND2_X1 U14984 ( .A1(n11698), .A2(n11697), .ZN(n11699) );
  OAI22_X1 U14985 ( .A1(n11699), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n19560), .ZN(n11706) );
  NAND2_X1 U14986 ( .A1(n11706), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11702) );
  NAND2_X1 U14987 ( .A1(n11699), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11707) );
  NOR2_X1 U14988 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n19560), .ZN(
        n11700) );
  NAND2_X1 U14989 ( .A1(n11707), .A2(n11700), .ZN(n11701) );
  NAND2_X1 U14990 ( .A1(n11702), .A2(n11701), .ZN(n13348) );
  XNOR2_X1 U14991 ( .A(n11704), .B(n11703), .ZN(n11705) );
  AOI21_X1 U14992 ( .B1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n11707), .A(
        n11706), .ZN(n11708) );
  XNOR2_X1 U14993 ( .A(n13345), .B(n13332), .ZN(n11710) );
  NAND2_X1 U14994 ( .A1(n20150), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n11716) );
  AOI211_X4 U14995 ( .C1(n18189), .C2(n20161), .A(n11718), .B(n11716), .ZN(
        n18580) );
  NAND2_X1 U14996 ( .A1(n18545), .A2(n18544), .ZN(n18541) );
  NAND2_X1 U14997 ( .A1(n18513), .A2(n18510), .ZN(n18507) );
  INV_X1 U14998 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n18488) );
  NAND2_X1 U14999 ( .A1(n18490), .A2(n18488), .ZN(n18485) );
  INV_X1 U15000 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n18459) );
  NAND2_X1 U15001 ( .A1(n18464), .A2(n18459), .ZN(n18458) );
  INV_X1 U15002 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n18717) );
  NAND2_X1 U15003 ( .A1(n18440), .A2(n18717), .ZN(n18434) );
  NAND2_X1 U15004 ( .A1(n18415), .A2(n18410), .ZN(n18409) );
  INV_X1 U15005 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n18384) );
  NAND2_X1 U15006 ( .A1(n18389), .A2(n18384), .ZN(n18383) );
  INV_X1 U15007 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n18364) );
  NAND2_X1 U15008 ( .A1(n18367), .A2(n18364), .ZN(n18363) );
  INV_X1 U15009 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n18340) );
  NAND2_X1 U15010 ( .A1(n18347), .A2(n18340), .ZN(n18337) );
  INV_X1 U15011 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n18676) );
  NAND2_X1 U15012 ( .A1(n18323), .A2(n18676), .ZN(n18316) );
  INV_X1 U15013 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n18294) );
  NAND2_X1 U15014 ( .A1(n18302), .A2(n18294), .ZN(n18293) );
  INV_X1 U15015 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n18271) );
  NAND2_X1 U15016 ( .A1(n18275), .A2(n18271), .ZN(n18270) );
  INV_X1 U15017 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n18248) );
  NAND2_X1 U15018 ( .A1(n18253), .A2(n18248), .ZN(n18247) );
  INV_X1 U15019 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n21826) );
  NAND2_X1 U15020 ( .A1(n18230), .A2(n21826), .ZN(n18209) );
  INV_X1 U15021 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n18621) );
  NAND2_X1 U15022 ( .A1(n18214), .A2(n18621), .ZN(n11730) );
  NAND2_X1 U15023 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n20154), .ZN(n20043) );
  NOR2_X1 U15024 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n17979) );
  NAND2_X1 U15025 ( .A1(n17979), .A2(n20151), .ZN(n20167) );
  OR2_X2 U15026 ( .A1(n20167), .A2(P3_STATE2_REG_0__SCAN_IN), .ZN(n19442) );
  NAND2_X1 U15027 ( .A1(n19442), .A2(n18536), .ZN(n18523) );
  INV_X1 U15028 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n11713) );
  NOR2_X1 U15029 ( .A1(n18558), .A2(n11713), .ZN(n11722) );
  NAND2_X2 U15030 ( .A1(n20144), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n20124) );
  NOR2_X1 U15031 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n20058) );
  INV_X1 U15032 ( .A(n20058), .ZN(n11714) );
  NAND3_X1 U15033 ( .A1(n20067), .A2(n20124), .A3(n11714), .ZN(n20065) );
  AND2_X1 U15034 ( .A1(n20161), .A2(n18189), .ZN(n11715) );
  OAI21_X1 U15035 ( .B1(n20149), .B2(n20150), .A(n11715), .ZN(n20038) );
  NAND2_X1 U15036 ( .A1(n20038), .A2(n11716), .ZN(n11717) );
  INV_X1 U15037 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n20123) );
  INV_X1 U15038 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n21849) );
  INV_X1 U15039 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n21832) );
  INV_X1 U15040 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n20108) );
  INV_X1 U15041 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n20099) );
  INV_X1 U15042 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n20093) );
  INV_X1 U15043 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n20091) );
  INV_X1 U15044 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n20087) );
  INV_X1 U15045 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n20082) );
  INV_X1 U15046 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n20077) );
  NAND2_X1 U15047 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_2__SCAN_IN), 
        .ZN(n18550) );
  NOR2_X1 U15048 ( .A1(n20077), .A2(n18550), .ZN(n18511) );
  NAND3_X1 U15049 ( .A1(n18511), .A2(P3_REIP_REG_5__SCAN_IN), .A3(
        P3_REIP_REG_4__SCAN_IN), .ZN(n18489) );
  NAND2_X1 U15050 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(P3_REIP_REG_7__SCAN_IN), 
        .ZN(n18463) );
  NOR4_X1 U15051 ( .A1(n20084), .A2(n20082), .A3(n18489), .A4(n18463), .ZN(
        n18438) );
  NAND2_X1 U15052 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(n18438), .ZN(n18431) );
  NOR2_X1 U15053 ( .A1(n20087), .A2(n18431), .ZN(n18422) );
  NAND2_X1 U15054 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n18422), .ZN(n18406) );
  NAND3_X1 U15055 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(P3_REIP_REG_15__SCAN_IN), 
        .A3(n18377), .ZN(n18358) );
  NOR2_X1 U15056 ( .A1(n20099), .A2(n18358), .ZN(n18329) );
  NAND4_X1 U15057 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(P3_REIP_REG_20__SCAN_IN), 
        .A3(P3_REIP_REG_18__SCAN_IN), .A4(n18329), .ZN(n18299) );
  NOR3_X1 U15058 ( .A1(n21832), .A2(n20108), .A3(n18299), .ZN(n18285) );
  NAND2_X1 U15059 ( .A1(P3_REIP_REG_23__SCAN_IN), .A2(n18285), .ZN(n18284) );
  NOR2_X1 U15060 ( .A1(n21849), .A2(n18284), .ZN(n18252) );
  NAND3_X1 U15061 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(P3_REIP_REG_25__SCAN_IN), 
        .A3(n18252), .ZN(n11724) );
  NOR2_X1 U15062 ( .A1(n18574), .A2(n11724), .ZN(n18246) );
  NAND4_X1 U15063 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .A4(n18246), .ZN(n11723) );
  NOR3_X1 U15064 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n20123), .A3(n11723), 
        .ZN(n11719) );
  AOI21_X1 U15065 ( .B1(n18581), .B2(P3_EBX_REG_31__SCAN_IN), .A(n11719), .ZN(
        n11720) );
  INV_X1 U15066 ( .A(n11720), .ZN(n11721) );
  NOR2_X1 U15067 ( .A1(n11722), .A2(n11721), .ZN(n11729) );
  NOR2_X1 U15068 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n11723), .ZN(n18213) );
  INV_X1 U15069 ( .A(n18213), .ZN(n11726) );
  NAND3_X1 U15070 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .ZN(n11725) );
  OR2_X1 U15071 ( .A1(n11724), .A2(n18576), .ZN(n18229) );
  NAND2_X1 U15072 ( .A1(n18574), .A2(n18564), .ZN(n18579) );
  OAI21_X1 U15073 ( .B1(n11725), .B2(n18229), .A(n18579), .ZN(n18228) );
  INV_X1 U15074 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n20120) );
  AOI21_X1 U15075 ( .B1(n11726), .B2(n18228), .A(n20120), .ZN(n11727) );
  NAND3_X1 U15076 ( .A1(n11730), .A2(n11729), .A3(n11728), .ZN(n11731) );
  INV_X1 U15077 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11733) );
  AND2_X2 U15078 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n11733), .ZN(
        n11742) );
  INV_X1 U15079 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11734) );
  NOR2_X4 U15080 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n14442) );
  AND2_X2 U15081 ( .A1(n11743), .A2(n14442), .ZN(n11792) );
  AOI22_X1 U15082 ( .A1(n11818), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11792), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11740) );
  INV_X2 U15083 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11736) );
  AND2_X4 U15084 ( .A1(n11736), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11741) );
  NOR2_X4 U15085 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13949) );
  AND2_X2 U15086 ( .A1(n11742), .A2(n13949), .ZN(n11838) );
  AOI22_X1 U15087 ( .A1(n12075), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11838), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11739) );
  NAND2_X2 U15088 ( .A1(n11741), .A2(n11742), .ZN(n11928) );
  NAND2_X4 U15089 ( .A1(n13949), .A2(n14442), .ZN(n12502) );
  AOI22_X1 U15090 ( .A1(n11995), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12019), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11738) );
  AOI22_X1 U15091 ( .A1(n11849), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n9691), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11737) );
  AND4_X2 U15092 ( .A1(n11740), .A2(n11739), .A3(n11738), .A4(n11737), .ZN(
        n11749) );
  AOI22_X1 U15093 ( .A1(n11824), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12131), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11747) );
  AOI22_X1 U15095 ( .A1(n11823), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11837), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11746) );
  AOI22_X1 U15096 ( .A1(n11936), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11797), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11745) );
  AOI22_X1 U15097 ( .A1(n11996), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11798), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11744) );
  AOI22_X1 U15098 ( .A1(n11823), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11837), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11753) );
  AOI22_X1 U15099 ( .A1(n11936), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11797), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11752) );
  AOI22_X1 U15100 ( .A1(n11824), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12131), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11751) );
  AOI22_X1 U15101 ( .A1(n11996), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11798), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11750) );
  NAND4_X1 U15102 ( .A1(n11753), .A2(n11752), .A3(n11751), .A4(n11750), .ZN(
        n11759) );
  AOI22_X1 U15103 ( .A1(n11995), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12019), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11757) );
  AOI22_X1 U15104 ( .A1(n9712), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11838), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11756) );
  AOI22_X1 U15105 ( .A1(n9715), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(n9691), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11754) );
  NAND4_X1 U15106 ( .A1(n11757), .A2(n11756), .A3(n11755), .A4(n11754), .ZN(
        n11758) );
  AOI22_X1 U15107 ( .A1(n11996), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n9697), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11763) );
  AOI22_X1 U15108 ( .A1(n12075), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11838), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11762) );
  AOI22_X1 U15109 ( .A1(n11818), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11792), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11760) );
  AOI22_X1 U15110 ( .A1(n9715), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(n9691), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11767) );
  AOI22_X1 U15111 ( .A1(n11823), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11837), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11766) );
  AOI22_X1 U15112 ( .A1(n9695), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n11797), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11765) );
  AOI22_X1 U15113 ( .A1(n11824), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12131), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11764) );
  AOI22_X1 U15114 ( .A1(n11995), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9715), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11773) );
  AOI22_X1 U15115 ( .A1(n11818), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11792), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11772) );
  AOI22_X1 U15116 ( .A1(n12131), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11797), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11771) );
  AOI22_X1 U15117 ( .A1(n11936), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n9695), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11770) );
  INV_X1 U15118 ( .A(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n21154) );
  INV_X1 U15119 ( .A(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11774) );
  OAI22_X1 U15120 ( .A1(n12502), .A2(n21154), .B1(n11950), .B2(n11774), .ZN(
        n11775) );
  INV_X1 U15121 ( .A(n11775), .ZN(n11777) );
  AOI22_X1 U15122 ( .A1(n11824), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11837), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11776) );
  NAND2_X1 U15123 ( .A1(n11777), .A2(n11776), .ZN(n11781) );
  AOI22_X1 U15124 ( .A1(n12075), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11838), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11779) );
  AOI22_X1 U15125 ( .A1(n11996), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11823), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11778) );
  NAND2_X1 U15126 ( .A1(n11779), .A2(n11778), .ZN(n11780) );
  NOR2_X1 U15127 ( .A1(n11781), .A2(n11780), .ZN(n11782) );
  INV_X2 U15128 ( .A(n11871), .ZN(n14381) );
  NAND2_X1 U15129 ( .A1(n9691), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n11785) );
  NAND2_X1 U15130 ( .A1(n11849), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n11784) );
  NAND2_X1 U15131 ( .A1(n11824), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n11791) );
  NAND2_X1 U15132 ( .A1(n12131), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n11790) );
  NAND2_X1 U15133 ( .A1(n11823), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n11789) );
  NAND2_X1 U15134 ( .A1(n11837), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n11788) );
  NAND2_X1 U15135 ( .A1(n11818), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n11796) );
  NAND2_X1 U15136 ( .A1(n11792), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n11795) );
  NAND2_X1 U15137 ( .A1(n12075), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n11794) );
  NAND2_X1 U15138 ( .A1(n11838), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n11793) );
  NAND2_X1 U15139 ( .A1(n11996), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11802) );
  NAND2_X1 U15140 ( .A1(n11936), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11801) );
  NAND2_X1 U15141 ( .A1(n11797), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n11800) );
  NAND2_X1 U15142 ( .A1(n11798), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n11799) );
  NAND2_X1 U15143 ( .A1(n11837), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n11810) );
  NAND2_X1 U15144 ( .A1(n9712), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n11809) );
  NAND2_X1 U15145 ( .A1(n12131), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11808) );
  NAND2_X1 U15146 ( .A1(n11797), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11807) );
  INV_X1 U15147 ( .A(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11811) );
  OR2_X1 U15148 ( .A1(n11950), .A2(n11811), .ZN(n11816) );
  NAND2_X1 U15149 ( .A1(n11849), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n11815) );
  NAND2_X1 U15150 ( .A1(n11838), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11814) );
  NAND2_X1 U15151 ( .A1(n11792), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11821) );
  NAND2_X1 U15152 ( .A1(n11996), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11820) );
  NAND2_X1 U15153 ( .A1(n9716), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11819) );
  NAND2_X1 U15154 ( .A1(n11823), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n11828) );
  NAND2_X1 U15155 ( .A1(n11824), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n11827) );
  NAND2_X1 U15156 ( .A1(n9697), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11826) );
  NAND2_X1 U15157 ( .A1(n9695), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n11825) );
  AOI22_X1 U15158 ( .A1(n11996), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12075), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11836) );
  AOI22_X1 U15159 ( .A1(n9697), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11798), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11833) );
  AOI22_X1 U15160 ( .A1(n11823), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11792), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11842) );
  AOI22_X1 U15161 ( .A1(n12131), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11837), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11841) );
  AOI22_X1 U15162 ( .A1(n11818), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11838), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11839) );
  AOI22_X1 U15163 ( .A1(n11995), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11838), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11848) );
  AOI22_X1 U15164 ( .A1(n11823), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9697), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11847) );
  AOI22_X1 U15165 ( .A1(n11996), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n9695), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11846) );
  AOI22_X1 U15166 ( .A1(n11824), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11837), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11845) );
  AOI22_X1 U15167 ( .A1(n12019), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12075), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11853) );
  AOI22_X1 U15168 ( .A1(n9691), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11849), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11852) );
  AOI22_X1 U15169 ( .A1(n9717), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11792), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11851) );
  AOI22_X1 U15170 ( .A1(n12131), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11797), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11850) );
  NAND2_X1 U15171 ( .A1(n13148), .A2(n11872), .ZN(n11891) );
  INV_X1 U15173 ( .A(n11855), .ZN(n11857) );
  NAND2_X2 U15174 ( .A1(n11857), .A2(n11856), .ZN(n11896) );
  NAND2_X1 U15175 ( .A1(n13148), .A2(n12634), .ZN(n11858) );
  NAND2_X1 U15176 ( .A1(n11858), .A2(n21617), .ZN(n13417) );
  INV_X1 U15177 ( .A(n11873), .ZN(n12571) );
  NAND2_X1 U15178 ( .A1(n12571), .A2(n11861), .ZN(n11859) );
  NOR2_X2 U15179 ( .A1(n11876), .A2(n11874), .ZN(n11897) );
  NAND2_X1 U15180 ( .A1(n11897), .A2(n13148), .ZN(n11895) );
  OAI21_X1 U15181 ( .B1(n11896), .B2(n13417), .A(n11895), .ZN(n11860) );
  AND2_X1 U15182 ( .A1(n14459), .A2(n11860), .ZN(n11884) );
  NAND2_X1 U15183 ( .A1(n14403), .A2(n11861), .ZN(n11862) );
  MUX2_X1 U15184 ( .A(n11862), .B(n13440), .S(n14381), .Z(n11865) );
  NAND3_X1 U15185 ( .A1(n11865), .A2(n11863), .A3(n11864), .ZN(n11888) );
  NAND2_X1 U15186 ( .A1(n11888), .A2(n13146), .ZN(n11883) );
  NAND2_X1 U15187 ( .A1(n14381), .A2(n12634), .ZN(n11866) );
  INV_X1 U15188 ( .A(n11890), .ZN(n11867) );
  NAND2_X1 U15189 ( .A1(n11870), .A2(n11869), .ZN(n12650) );
  NAND2_X1 U15190 ( .A1(n12674), .A2(n13145), .ZN(n13441) );
  INV_X1 U15191 ( .A(n11876), .ZN(n13147) );
  INV_X1 U15192 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n11878) );
  XNOR2_X1 U15193 ( .A(n11878), .B(P1_STATE_REG_2__SCAN_IN), .ZN(n12741) );
  NAND4_X1 U15194 ( .A1(n11884), .A2(n11883), .A3(n11882), .A4(n11881), .ZN(
        n11885) );
  NAND2_X1 U15195 ( .A1(n11885), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11919) );
  INV_X1 U15196 ( .A(n13153), .ZN(n11886) );
  MUX2_X1 U15197 ( .A(n11886), .B(n15966), .S(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Z(n11887) );
  INV_X1 U15198 ( .A(n12623), .ZN(n11889) );
  INV_X4 U15199 ( .A(n12726), .ZN(n14821) );
  NAND2_X1 U15200 ( .A1(n11891), .A2(n14821), .ZN(n11892) );
  NAND3_X1 U15201 ( .A1(n11895), .A2(n11896), .A3(n10514), .ZN(n11901) );
  OR2_X1 U15202 ( .A1(n11907), .A2(n11861), .ZN(n13459) );
  INV_X1 U15203 ( .A(n11897), .ZN(n11898) );
  NAND2_X1 U15204 ( .A1(n11898), .A2(n15959), .ZN(n11899) );
  NAND2_X1 U15205 ( .A1(n21414), .A2(n21681), .ZN(n15898) );
  NAND2_X1 U15206 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n14525) );
  AND2_X1 U15207 ( .A1(n15898), .A2(n14525), .ZN(n21380) );
  AND2_X1 U15208 ( .A1(n15961), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n11915) );
  AOI21_X1 U15209 ( .B1(n13153), .B2(n21380), .A(n11915), .ZN(n11905) );
  NAND2_X1 U15210 ( .A1(n11908), .A2(n13450), .ZN(n14435) );
  INV_X1 U15211 ( .A(n14136), .ZN(n14138) );
  NAND2_X1 U15212 ( .A1(n13945), .A2(n14138), .ZN(n13431) );
  OAI21_X1 U15213 ( .B1(n12622), .B2(n11879), .A(n13431), .ZN(n11909) );
  OAI21_X1 U15214 ( .B1(n11909), .B2(n13433), .A(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n11910) );
  INV_X1 U15215 ( .A(n11910), .ZN(n11914) );
  INV_X1 U15216 ( .A(n11944), .ZN(n11912) );
  INV_X1 U15217 ( .A(n11915), .ZN(n11916) );
  NAND2_X1 U15218 ( .A1(n11916), .A2(n13958), .ZN(n11917) );
  INV_X1 U15219 ( .A(n11919), .ZN(n11921) );
  AND2_X1 U15220 ( .A1(n15961), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11920) );
  XNOR2_X1 U15221 ( .A(n14525), .B(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n15802) );
  NAND2_X1 U15222 ( .A1(n13153), .A2(n15802), .ZN(n11967) );
  NAND2_X1 U15223 ( .A1(n11921), .A2(n15788), .ZN(n11926) );
  INV_X1 U15224 ( .A(n14525), .ZN(n21235) );
  INV_X1 U15225 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n15793) );
  NAND2_X1 U15226 ( .A1(n15793), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n21269) );
  INV_X1 U15227 ( .A(n21269), .ZN(n11922) );
  NAND2_X1 U15228 ( .A1(n21235), .A2(n11922), .ZN(n14500) );
  NAND2_X1 U15229 ( .A1(n14500), .A2(n15793), .ZN(n11924) );
  NAND2_X1 U15230 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n21464) );
  INV_X1 U15231 ( .A(n21464), .ZN(n11923) );
  NAND2_X1 U15232 ( .A1(n21235), .A2(n11923), .ZN(n14404) );
  AOI22_X1 U15233 ( .A1(n15852), .A2(n13153), .B1(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n15961), .ZN(n11925) );
  AOI22_X1 U15234 ( .A1(n12550), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9707), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11935) );
  AOI22_X1 U15235 ( .A1(n12395), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12373), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11934) );
  AOI22_X1 U15236 ( .A1(n9706), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12527), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11933) );
  INV_X1 U15237 ( .A(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11930) );
  INV_X1 U15238 ( .A(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11929) );
  OAI22_X1 U15239 ( .A1(n9701), .A2(n11930), .B1(n12502), .B2(n11929), .ZN(
        n11931) );
  INV_X1 U15240 ( .A(n11931), .ZN(n11932) );
  NAND4_X1 U15241 ( .A1(n11935), .A2(n11934), .A3(n11933), .A4(n11932), .ZN(
        n11942) );
  INV_X1 U15242 ( .A(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n21653) );
  AOI22_X1 U15243 ( .A1(n9713), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12378), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11940) );
  AOI22_X1 U15244 ( .A1(n9690), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11837), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11939) );
  AOI22_X1 U15245 ( .A1(n9711), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12488), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11938) );
  AOI22_X1 U15246 ( .A1(n9689), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12545), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11937) );
  NAND4_X1 U15247 ( .A1(n11940), .A2(n11939), .A3(n11938), .A4(n11937), .ZN(
        n11941) );
  AOI22_X1 U15248 ( .A1(n12568), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12594), .B2(n13109), .ZN(n11943) );
  AOI22_X1 U15249 ( .A1(n9713), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(n9690), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11949) );
  AOI22_X1 U15250 ( .A1(n12544), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12527), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11948) );
  AOI22_X1 U15251 ( .A1(n9689), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12373), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11947) );
  AOI22_X1 U15252 ( .A1(n9711), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n12488), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11946) );
  NAND4_X1 U15253 ( .A1(n11949), .A2(n11948), .A3(n11947), .A4(n11946), .ZN(
        n11959) );
  AOI22_X1 U15254 ( .A1(n12378), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12526), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11957) );
  AOI22_X1 U15255 ( .A1(n9712), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12550), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11956) );
  INV_X1 U15256 ( .A(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11952) );
  INV_X1 U15257 ( .A(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11951) );
  OAI22_X1 U15258 ( .A1(n12502), .A2(n11952), .B1(n12500), .B2(n11951), .ZN(
        n11953) );
  INV_X1 U15259 ( .A(n11953), .ZN(n11955) );
  AOI22_X1 U15260 ( .A1(n9707), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12545), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11954) );
  NAND4_X1 U15261 ( .A1(n11957), .A2(n11956), .A3(n11955), .A4(n11954), .ZN(
        n11958) );
  NAND2_X1 U15262 ( .A1(n12089), .A2(n13084), .ZN(n11960) );
  NAND2_X1 U15263 ( .A1(n13146), .A2(n13084), .ZN(n11963) );
  AOI21_X1 U15264 ( .B1(n12568), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A(
        n12089), .ZN(n11964) );
  INV_X1 U15265 ( .A(n11966), .ZN(n11969) );
  INV_X1 U15266 ( .A(n11967), .ZN(n11968) );
  AOI22_X1 U15267 ( .A1(n12550), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9707), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11976) );
  AOI22_X1 U15268 ( .A1(n12075), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12373), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11975) );
  AOI22_X1 U15269 ( .A1(n9706), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12527), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11974) );
  INV_X1 U15270 ( .A(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11971) );
  INV_X1 U15271 ( .A(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11970) );
  OAI22_X1 U15272 ( .A1(n9701), .A2(n11971), .B1(n12502), .B2(n11970), .ZN(
        n11972) );
  INV_X1 U15273 ( .A(n11972), .ZN(n11973) );
  NAND4_X1 U15274 ( .A1(n11976), .A2(n11975), .A3(n11974), .A4(n11973), .ZN(
        n11982) );
  AOI22_X1 U15275 ( .A1(n9713), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12378), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11980) );
  AOI22_X1 U15276 ( .A1(n9690), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11837), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11979) );
  AOI22_X1 U15277 ( .A1(n9711), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n12488), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11978) );
  AOI22_X1 U15278 ( .A1(n9689), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12545), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11977) );
  NAND4_X1 U15279 ( .A1(n11980), .A2(n11979), .A3(n11978), .A4(n11977), .ZN(
        n11981) );
  NAND3_X1 U15280 ( .A1(n13146), .A2(P1_STATE2_REG_0__SCAN_IN), .A3(n11984), 
        .ZN(n11983) );
  OAI21_X1 U15281 ( .B1(n12606), .B2(n21154), .A(n11983), .ZN(n11987) );
  INV_X1 U15282 ( .A(n12089), .ZN(n11985) );
  NOR2_X1 U15283 ( .A1(n13098), .A2(n11985), .ZN(n11986) );
  INV_X1 U15284 ( .A(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n21162) );
  AOI22_X1 U15285 ( .A1(n9713), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11837), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11994) );
  AOI22_X1 U15286 ( .A1(n9690), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n9711), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11993) );
  AOI22_X1 U15287 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n9706), .B1(
        n12395), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11992) );
  AOI22_X1 U15288 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n12550), .B1(
        n9707), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11991) );
  NAND4_X1 U15289 ( .A1(n11994), .A2(n11993), .A3(n11992), .A4(n11991), .ZN(
        n12002) );
  AOI22_X1 U15290 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n12483), .B1(
        n12527), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12000) );
  AOI22_X1 U15291 ( .A1(n12544), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12373), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11999) );
  AOI22_X1 U15292 ( .A1(n12378), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12488), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11998) );
  AOI22_X1 U15293 ( .A1(n9689), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12545), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11997) );
  NAND4_X1 U15294 ( .A1(n12000), .A2(n11999), .A3(n11998), .A4(n11997), .ZN(
        n12001) );
  NAND2_X1 U15295 ( .A1(n12594), .A2(n13108), .ZN(n12003) );
  INV_X1 U15296 ( .A(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12018) );
  AOI22_X1 U15297 ( .A1(n12550), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9707), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12010) );
  AOI22_X1 U15298 ( .A1(n12395), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12373), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12009) );
  AOI22_X1 U15299 ( .A1(n9706), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12527), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12008) );
  INV_X1 U15300 ( .A(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12005) );
  INV_X1 U15301 ( .A(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12004) );
  OAI22_X1 U15302 ( .A1(n9701), .A2(n12005), .B1(n12502), .B2(n12004), .ZN(
        n12006) );
  INV_X1 U15303 ( .A(n12006), .ZN(n12007) );
  NAND4_X1 U15304 ( .A1(n12010), .A2(n12009), .A3(n12008), .A4(n12007), .ZN(
        n12016) );
  AOI22_X1 U15305 ( .A1(n9713), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12378), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12014) );
  AOI22_X1 U15306 ( .A1(n9690), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12526), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12013) );
  AOI22_X1 U15307 ( .A1(n9711), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12488), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12012) );
  AOI22_X1 U15308 ( .A1(n9689), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12545), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12011) );
  NAND4_X1 U15309 ( .A1(n12014), .A2(n12013), .A3(n12012), .A4(n12011), .ZN(
        n12015) );
  NAND2_X1 U15310 ( .A1(n12594), .A2(n13118), .ZN(n12017) );
  NAND2_X1 U15311 ( .A1(n12568), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n12031) );
  AOI22_X1 U15312 ( .A1(n12378), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12526), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12023) );
  AOI22_X1 U15313 ( .A1(n9689), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9690), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12022) );
  AOI22_X1 U15314 ( .A1(n9706), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12527), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12021) );
  AOI22_X1 U15315 ( .A1(n12483), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n9707), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12020) );
  NAND4_X1 U15316 ( .A1(n12023), .A2(n12022), .A3(n12021), .A4(n12020), .ZN(
        n12029) );
  AOI22_X1 U15317 ( .A1(n12395), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12550), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12027) );
  AOI22_X1 U15318 ( .A1(n12544), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12373), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12026) );
  AOI22_X1 U15319 ( .A1(n9713), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12488), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12025) );
  AOI22_X1 U15320 ( .A1(n9711), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n12545), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12024) );
  NAND4_X1 U15321 ( .A1(n12027), .A2(n12026), .A3(n12025), .A4(n12024), .ZN(
        n12028) );
  NAND2_X1 U15322 ( .A1(n12594), .A2(n13129), .ZN(n12030) );
  INV_X1 U15323 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12046) );
  AOI22_X1 U15324 ( .A1(n12550), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9707), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12039) );
  AOI22_X1 U15325 ( .A1(n12075), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12373), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12038) );
  AOI22_X1 U15326 ( .A1(n9706), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12527), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12037) );
  INV_X1 U15327 ( .A(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12034) );
  INV_X1 U15328 ( .A(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12033) );
  OAI22_X1 U15329 ( .A1(n9701), .A2(n12034), .B1(n12502), .B2(n12033), .ZN(
        n12035) );
  INV_X1 U15330 ( .A(n12035), .ZN(n12036) );
  NAND4_X1 U15331 ( .A1(n12039), .A2(n12038), .A3(n12037), .A4(n12036), .ZN(
        n12045) );
  AOI22_X1 U15332 ( .A1(n9713), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12378), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12043) );
  AOI22_X1 U15333 ( .A1(n9690), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12526), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12042) );
  AOI22_X1 U15334 ( .A1(n9711), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n12488), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12041) );
  AOI22_X1 U15335 ( .A1(n11996), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12545), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12040) );
  NAND4_X1 U15336 ( .A1(n12043), .A2(n12042), .A3(n12041), .A4(n12040), .ZN(
        n12044) );
  INV_X1 U15337 ( .A(n13131), .ZN(n13135) );
  OAI22_X1 U15338 ( .A1(n12606), .A2(n12046), .B1(n12614), .B2(n13135), .ZN(
        n12047) );
  INV_X1 U15339 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n12052) );
  INV_X1 U15340 ( .A(n12122), .ZN(n12049) );
  NAND2_X1 U15341 ( .A1(n12049), .A2(n10138), .ZN(n12050) );
  NAND2_X1 U15342 ( .A1(n12152), .A2(n12050), .ZN(n20974) );
  NAND2_X1 U15343 ( .A1(n21349), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12062) );
  AOI22_X1 U15344 ( .A1(n20974), .A2(n12058), .B1(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n12563), .ZN(n12051) );
  OAI21_X1 U15345 ( .B1(n9815), .B2(n12052), .A(n12051), .ZN(n12053) );
  AOI21_X1 U15346 ( .B1(n13126), .B2(n12254), .A(n12053), .ZN(n15200) );
  INV_X1 U15347 ( .A(n15200), .ZN(n12126) );
  AND2_X1 U15348 ( .A1(n14138), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12070) );
  INV_X1 U15349 ( .A(n12070), .ZN(n12108) );
  INV_X1 U15350 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n12613) );
  NAND2_X1 U15351 ( .A1(n21349), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12056) );
  NAND2_X1 U15352 ( .A1(n12456), .A2(P1_EAX_REG_4__SCAN_IN), .ZN(n12055) );
  OAI211_X1 U15353 ( .C1(n12108), .C2(n12613), .A(n12056), .B(n12055), .ZN(
        n12059) );
  INV_X1 U15354 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n12057) );
  XNOR2_X1 U15355 ( .A(n12113), .B(n12057), .ZN(n21099) );
  MUX2_X1 U15356 ( .A(n12059), .B(n21099), .S(n12058), .Z(n12060) );
  AOI21_X1 U15357 ( .B1(n13080), .B2(n12254), .A(n12060), .ZN(n14413) );
  INV_X1 U15358 ( .A(n14413), .ZN(n12111) );
  NAND2_X1 U15359 ( .A1(n13097), .A2(n12254), .ZN(n12067) );
  NAND2_X1 U15360 ( .A1(n12070), .A2(n15783), .ZN(n12065) );
  INV_X1 U15361 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n14278) );
  XNOR2_X1 U15362 ( .A(n14278), .B(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n21028) );
  OAI21_X1 U15363 ( .B1(n21028), .B2(n12631), .A(n12062), .ZN(n12063) );
  AOI21_X1 U15364 ( .B1(n12456), .B2(P1_EAX_REG_2__SCAN_IN), .A(n12063), .ZN(
        n12064) );
  AND2_X1 U15365 ( .A1(n12065), .A2(n12064), .ZN(n12066) );
  NAND2_X1 U15366 ( .A1(n12067), .A2(n12066), .ZN(n12068) );
  NAND2_X1 U15367 ( .A1(n12563), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12102) );
  NAND2_X1 U15368 ( .A1(n12068), .A2(n12102), .ZN(n14263) );
  NAND2_X1 U15369 ( .A1(n14363), .A2(n12254), .ZN(n12074) );
  AOI22_X1 U15370 ( .A1(n12456), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n21349), .ZN(n12072) );
  NAND2_X1 U15371 ( .A1(n12070), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12071) );
  AND2_X1 U15372 ( .A1(n12072), .A2(n12071), .ZN(n12073) );
  AOI22_X1 U15373 ( .A1(n12544), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9712), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12079) );
  AOI22_X1 U15374 ( .A1(n9706), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12527), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12078) );
  AOI22_X1 U15375 ( .A1(n11996), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9711), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12077) );
  AOI22_X1 U15376 ( .A1(n12526), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12488), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12076) );
  NAND4_X1 U15377 ( .A1(n12079), .A2(n12078), .A3(n12077), .A4(n12076), .ZN(
        n12085) );
  AOI22_X1 U15378 ( .A1(n9713), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12378), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12083) );
  AOI22_X1 U15379 ( .A1(n12550), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n9707), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12082) );
  AOI22_X1 U15380 ( .A1(n12483), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12373), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12081) );
  AOI22_X1 U15381 ( .A1(n9690), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12545), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12080) );
  NAND4_X1 U15382 ( .A1(n12083), .A2(n12082), .A3(n12081), .A4(n12080), .ZN(
        n12084) );
  AOI21_X1 U15383 ( .B1(n13146), .B2(n13089), .A(n20939), .ZN(n12087) );
  NAND2_X1 U15384 ( .A1(n13435), .A2(n13131), .ZN(n13070) );
  OAI211_X1 U15385 ( .C1(n12606), .C2(n15807), .A(n12087), .B(n13070), .ZN(
        n12092) );
  INV_X1 U15386 ( .A(n13089), .ZN(n12088) );
  XNOR2_X1 U15387 ( .A(n12088), .B(n13131), .ZN(n12090) );
  NAND2_X1 U15388 ( .A1(n12090), .A2(n12089), .ZN(n12091) );
  XNOR2_X1 U15389 ( .A(n12092), .B(n12091), .ZN(n12093) );
  NAND2_X1 U15390 ( .A1(n12094), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n14085) );
  NAND2_X1 U15391 ( .A1(n21349), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12096) );
  NAND2_X1 U15392 ( .A1(n12456), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n12095) );
  OAI211_X1 U15393 ( .C1(n12108), .C2(n11736), .A(n12096), .B(n12095), .ZN(
        n12097) );
  OR2_X1 U15394 ( .A1(n14085), .A2(n12098), .ZN(n14086) );
  INV_X1 U15395 ( .A(n12098), .ZN(n14087) );
  OR2_X1 U15396 ( .A1(n14087), .A2(n12631), .ZN(n12099) );
  NAND2_X1 U15397 ( .A1(n14086), .A2(n12099), .ZN(n14094) );
  NAND2_X1 U15398 ( .A1(n12101), .A2(n12100), .ZN(n14261) );
  INV_X1 U15399 ( .A(n12254), .ZN(n12187) );
  INV_X1 U15400 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n15503) );
  NAND2_X1 U15401 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12104) );
  NAND2_X1 U15402 ( .A1(n15503), .A2(n12104), .ZN(n12105) );
  NAND2_X1 U15403 ( .A1(n12113), .A2(n12105), .ZN(n15148) );
  AOI22_X1 U15404 ( .A1(n12058), .A2(n15148), .B1(n12563), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n12107) );
  NAND2_X1 U15405 ( .A1(n12456), .A2(P1_EAX_REG_3__SCAN_IN), .ZN(n12106) );
  OAI211_X1 U15406 ( .C1(n12108), .C2(n11735), .A(n12107), .B(n12106), .ZN(
        n12109) );
  INV_X1 U15407 ( .A(n12109), .ZN(n12110) );
  OAI21_X2 U15408 ( .B1(n14524), .B2(n12187), .A(n12110), .ZN(n14411) );
  INV_X1 U15409 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n12116) );
  AOI21_X1 U15410 ( .B1(n10141), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n12114) );
  OR2_X1 U15411 ( .A1(n12114), .A2(n12120), .ZN(n20997) );
  AOI22_X1 U15412 ( .A1(n20997), .A2(n12058), .B1(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n12563), .ZN(n12115) );
  OAI21_X1 U15413 ( .B1(n9815), .B2(n12116), .A(n12115), .ZN(n12117) );
  AOI21_X1 U15414 ( .B1(n13107), .B2(n12254), .A(n12117), .ZN(n14427) );
  NOR2_X2 U15415 ( .A1(n14410), .A2(n14427), .ZN(n14428) );
  INV_X1 U15416 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n21045) );
  NAND2_X1 U15417 ( .A1(n12119), .A2(n12118), .ZN(n13117) );
  NAND2_X1 U15418 ( .A1(n13117), .A2(n12254), .ZN(n12124) );
  NOR2_X1 U15419 ( .A1(n12120), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12121) );
  OR2_X1 U15420 ( .A1(n12122), .A2(n12121), .ZN(n20985) );
  AOI22_X1 U15421 ( .A1(n20985), .A2(n12058), .B1(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n12563), .ZN(n12123) );
  OAI211_X1 U15422 ( .C1(n9815), .C2(n21045), .A(n12124), .B(n12123), .ZN(
        n14572) );
  NAND2_X1 U15423 ( .A1(n14428), .A2(n14572), .ZN(n14570) );
  AOI22_X1 U15424 ( .A1(n9690), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n12526), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12130) );
  AOI22_X1 U15425 ( .A1(n9706), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12527), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12129) );
  AOI22_X1 U15426 ( .A1(n12544), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12550), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12128) );
  AOI22_X1 U15427 ( .A1(n9711), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12488), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12127) );
  NAND4_X1 U15428 ( .A1(n12130), .A2(n12129), .A3(n12128), .A4(n12127), .ZN(
        n12137) );
  AOI22_X1 U15429 ( .A1(n9713), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12378), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12135) );
  AOI22_X1 U15430 ( .A1(n12395), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n9707), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12134) );
  AOI22_X1 U15431 ( .A1(n12483), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12373), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12133) );
  AOI22_X1 U15432 ( .A1(n9689), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12545), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12132) );
  NAND4_X1 U15433 ( .A1(n12135), .A2(n12134), .A3(n12133), .A4(n12132), .ZN(
        n12136) );
  OAI21_X1 U15434 ( .B1(n12137), .B2(n12136), .A(n12254), .ZN(n12141) );
  NAND2_X1 U15435 ( .A1(n12456), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n12140) );
  XNOR2_X1 U15436 ( .A(n12152), .B(n15138), .ZN(n15488) );
  NAND2_X1 U15437 ( .A1(n15488), .A2(n12058), .ZN(n12139) );
  NAND2_X1 U15438 ( .A1(n12563), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12138) );
  AOI22_X1 U15439 ( .A1(n9690), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n12526), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12145) );
  AOI22_X1 U15440 ( .A1(n12483), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12527), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12144) );
  AOI22_X1 U15441 ( .A1(n12544), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12373), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12143) );
  AOI22_X1 U15442 ( .A1(n12550), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12488), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12142) );
  NAND4_X1 U15443 ( .A1(n12145), .A2(n12144), .A3(n12143), .A4(n12142), .ZN(
        n12151) );
  AOI22_X1 U15444 ( .A1(n9713), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12378), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12149) );
  AOI22_X1 U15445 ( .A1(n9706), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12395), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12148) );
  AOI22_X1 U15446 ( .A1(n9689), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9707), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12147) );
  AOI22_X1 U15447 ( .A1(n9711), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12545), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12146) );
  NAND4_X1 U15448 ( .A1(n12149), .A2(n12148), .A3(n12147), .A4(n12146), .ZN(
        n12150) );
  OAI21_X1 U15449 ( .B1(n12151), .B2(n12150), .A(n12254), .ZN(n12156) );
  NAND2_X1 U15450 ( .A1(n12456), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n12155) );
  XNOR2_X1 U15451 ( .A(n12157), .B(n10155), .ZN(n15480) );
  NAND2_X1 U15452 ( .A1(n15480), .A2(n12058), .ZN(n12154) );
  NAND2_X1 U15453 ( .A1(n12563), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12153) );
  NAND4_X1 U15454 ( .A1(n12156), .A2(n12155), .A3(n12154), .A4(n12153), .ZN(
        n15114) );
  XNOR2_X1 U15455 ( .A(n12184), .B(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15470) );
  AOI22_X1 U15456 ( .A1(n12456), .A2(P1_EAX_REG_10__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n12563), .ZN(n12170) );
  AOI22_X1 U15457 ( .A1(n9690), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12526), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12162) );
  AOI22_X1 U15458 ( .A1(n9706), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12527), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12161) );
  AOI22_X1 U15459 ( .A1(n12544), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12550), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12160) );
  AOI22_X1 U15460 ( .A1(n9711), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12488), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12159) );
  NAND4_X1 U15461 ( .A1(n12162), .A2(n12161), .A3(n12160), .A4(n12159), .ZN(
        n12168) );
  AOI22_X1 U15462 ( .A1(n9713), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12378), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12166) );
  AOI22_X1 U15463 ( .A1(n12395), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n9707), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12165) );
  AOI22_X1 U15464 ( .A1(n12483), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12373), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12164) );
  AOI22_X1 U15465 ( .A1(n9689), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12545), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12163) );
  NAND4_X1 U15466 ( .A1(n12166), .A2(n12165), .A3(n12164), .A4(n12163), .ZN(
        n12167) );
  OAI21_X1 U15467 ( .B1(n12168), .B2(n12167), .A(n12254), .ZN(n12169) );
  OAI211_X1 U15468 ( .C1(n15470), .C2(n12631), .A(n12170), .B(n12169), .ZN(
        n15100) );
  AOI22_X1 U15469 ( .A1(n9689), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9707), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12174) );
  AOI22_X1 U15470 ( .A1(n12544), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12527), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12173) );
  AOI22_X1 U15471 ( .A1(n12395), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12373), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12172) );
  AOI22_X1 U15472 ( .A1(n12526), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12545), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12171) );
  NAND4_X1 U15473 ( .A1(n12174), .A2(n12173), .A3(n12172), .A4(n12171), .ZN(
        n12183) );
  AOI22_X1 U15474 ( .A1(n9713), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12378), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12181) );
  AOI22_X1 U15475 ( .A1(n9711), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12550), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12180) );
  INV_X1 U15476 ( .A(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12176) );
  INV_X1 U15477 ( .A(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12175) );
  OAI22_X1 U15478 ( .A1(n12502), .A2(n12176), .B1(n12500), .B2(n12175), .ZN(
        n12177) );
  INV_X1 U15479 ( .A(n12177), .ZN(n12179) );
  AOI22_X1 U15480 ( .A1(n9690), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12488), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12178) );
  NAND4_X1 U15481 ( .A1(n12181), .A2(n12180), .A3(n12179), .A4(n12178), .ZN(
        n12182) );
  NOR2_X1 U15482 ( .A1(n12183), .A2(n12182), .ZN(n12188) );
  XNOR2_X1 U15483 ( .A(n12262), .B(n15025), .ZN(n15421) );
  NAND2_X1 U15484 ( .A1(n15421), .A2(n12058), .ZN(n12186) );
  AOI22_X1 U15485 ( .A1(n12456), .A2(P1_EAX_REG_15__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n12563), .ZN(n12185) );
  OAI211_X1 U15486 ( .C1(n12188), .C2(n12187), .A(n12186), .B(n12185), .ZN(
        n15023) );
  AOI22_X1 U15487 ( .A1(n9689), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12378), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12194) );
  AOI22_X1 U15488 ( .A1(n12550), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n9707), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12193) );
  AOI22_X1 U15489 ( .A1(n12395), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12373), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12192) );
  INV_X1 U15490 ( .A(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12189) );
  INV_X1 U15491 ( .A(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12464) );
  OAI22_X1 U15492 ( .A1(n12502), .A2(n12189), .B1(n12500), .B2(n12464), .ZN(
        n12190) );
  INV_X1 U15493 ( .A(n12190), .ZN(n12191) );
  NAND4_X1 U15494 ( .A1(n12194), .A2(n12193), .A3(n12192), .A4(n12191), .ZN(
        n12200) );
  AOI22_X1 U15495 ( .A1(n12544), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12527), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12198) );
  AOI22_X1 U15496 ( .A1(n9713), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12526), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12197) );
  AOI22_X1 U15497 ( .A1(n9690), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12488), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12196) );
  AOI22_X1 U15498 ( .A1(n9711), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12545), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12195) );
  NAND4_X1 U15499 ( .A1(n12198), .A2(n12197), .A3(n12196), .A4(n12195), .ZN(
        n12199) );
  OR2_X1 U15500 ( .A1(n12200), .A2(n12199), .ZN(n12201) );
  AND2_X1 U15501 ( .A1(n12254), .A2(n12201), .ZN(n15087) );
  NAND2_X1 U15502 ( .A1(n12203), .A2(n12202), .ZN(n12204) );
  NAND2_X1 U15503 ( .A1(n12225), .A2(n12204), .ZN(n15460) );
  NAND2_X1 U15504 ( .A1(n15460), .A2(n12058), .ZN(n12206) );
  AOI22_X1 U15505 ( .A1(n12456), .A2(P1_EAX_REG_11__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n12563), .ZN(n12205) );
  NAND2_X1 U15506 ( .A1(n12206), .A2(n12205), .ZN(n15049) );
  XNOR2_X1 U15507 ( .A(n12208), .B(n12207), .ZN(n15444) );
  NAND2_X1 U15508 ( .A1(n15444), .A2(n12058), .ZN(n12224) );
  AOI22_X1 U15509 ( .A1(n12378), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12526), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12214) );
  AOI22_X1 U15510 ( .A1(n12395), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n9707), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12213) );
  INV_X1 U15511 ( .A(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12209) );
  INV_X1 U15512 ( .A(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12503) );
  OAI22_X1 U15513 ( .A1(n12502), .A2(n12209), .B1(n12500), .B2(n12503), .ZN(
        n12210) );
  INV_X1 U15514 ( .A(n12210), .ZN(n12212) );
  AOI22_X1 U15515 ( .A1(n9689), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12545), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12211) );
  NAND4_X1 U15516 ( .A1(n12214), .A2(n12213), .A3(n12212), .A4(n12211), .ZN(
        n12220) );
  AOI22_X1 U15517 ( .A1(n9713), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(n9690), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12218) );
  AOI22_X1 U15518 ( .A1(n12544), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12527), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12217) );
  AOI22_X1 U15519 ( .A1(n12550), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12373), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12216) );
  AOI22_X1 U15520 ( .A1(n9711), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12488), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12215) );
  NAND4_X1 U15521 ( .A1(n12218), .A2(n12217), .A3(n12216), .A4(n12215), .ZN(
        n12219) );
  OAI21_X1 U15522 ( .B1(n12220), .B2(n12219), .A(n12254), .ZN(n12223) );
  NAND2_X1 U15523 ( .A1(n12456), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n12222) );
  NAND2_X1 U15524 ( .A1(n12563), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n12221) );
  NAND2_X1 U15525 ( .A1(n12224), .A2(n10642), .ZN(n15053) );
  XNOR2_X1 U15526 ( .A(n12225), .B(n15451), .ZN(n15078) );
  NAND2_X1 U15527 ( .A1(n15078), .A2(n12058), .ZN(n12242) );
  AOI22_X1 U15528 ( .A1(n9690), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n12526), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12232) );
  AOI22_X1 U15529 ( .A1(n9689), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12373), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12231) );
  INV_X1 U15530 ( .A(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12227) );
  INV_X1 U15531 ( .A(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12226) );
  OAI22_X1 U15532 ( .A1(n12227), .A2(n9701), .B1(n12502), .B2(n12226), .ZN(
        n12228) );
  INV_X1 U15533 ( .A(n12228), .ZN(n12230) );
  AOI22_X1 U15534 ( .A1(n12545), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12488), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12229) );
  NAND4_X1 U15535 ( .A1(n12232), .A2(n12231), .A3(n12230), .A4(n12229), .ZN(
        n12238) );
  AOI22_X1 U15536 ( .A1(n9713), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12378), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12236) );
  AOI22_X1 U15537 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n9711), .B1(n9707), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12235) );
  AOI22_X1 U15538 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n9706), .B1(
        n12527), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12234) );
  AOI22_X1 U15539 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n12395), .B1(
        n12550), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12233) );
  NAND4_X1 U15540 ( .A1(n12236), .A2(n12235), .A3(n12234), .A4(n12233), .ZN(
        n12237) );
  OAI21_X1 U15541 ( .B1(n12238), .B2(n12237), .A(n12254), .ZN(n12241) );
  NAND2_X1 U15542 ( .A1(n12456), .A2(P1_EAX_REG_12__SCAN_IN), .ZN(n12240) );
  NAND2_X1 U15543 ( .A1(n12563), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12239) );
  NAND2_X1 U15544 ( .A1(n12242), .A2(n10630), .ZN(n15069) );
  OAI211_X1 U15545 ( .C1(n15087), .C2(n15049), .A(n15053), .B(n15069), .ZN(
        n12243) );
  INV_X1 U15546 ( .A(n12243), .ZN(n12261) );
  INV_X1 U15547 ( .A(n12244), .ZN(n12245) );
  XNOR2_X1 U15548 ( .A(n12245), .B(n10150), .ZN(n15432) );
  NAND2_X1 U15549 ( .A1(n15432), .A2(n12058), .ZN(n12260) );
  AOI22_X1 U15550 ( .A1(n9713), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(n9690), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12249) );
  AOI22_X1 U15551 ( .A1(n9689), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9711), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12248) );
  AOI22_X1 U15552 ( .A1(n12395), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n9707), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12247) );
  AOI22_X1 U15553 ( .A1(n12483), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12373), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12246) );
  NAND4_X1 U15554 ( .A1(n12249), .A2(n12248), .A3(n12247), .A4(n12246), .ZN(
        n12256) );
  AOI22_X1 U15555 ( .A1(n12378), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12526), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12253) );
  AOI22_X1 U15556 ( .A1(n9706), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12527), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12252) );
  AOI22_X1 U15557 ( .A1(n12544), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12550), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12251) );
  AOI22_X1 U15558 ( .A1(n12545), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12488), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12250) );
  NAND4_X1 U15559 ( .A1(n12253), .A2(n12252), .A3(n12251), .A4(n12250), .ZN(
        n12255) );
  OAI21_X1 U15560 ( .B1(n12256), .B2(n12255), .A(n12254), .ZN(n12259) );
  NAND2_X1 U15561 ( .A1(n12456), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n12258) );
  NAND2_X1 U15562 ( .A1(n12563), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12257) );
  NAND2_X1 U15563 ( .A1(n12260), .A2(n10631), .ZN(n15033) );
  XNOR2_X1 U15564 ( .A(n12282), .B(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15407) );
  NAND2_X1 U15565 ( .A1(n15407), .A2(n12058), .ZN(n12279) );
  AOI22_X1 U15566 ( .A1(n12483), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n9689), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12266) );
  AOI22_X1 U15567 ( .A1(n12395), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n9690), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12265) );
  AOI22_X1 U15568 ( .A1(n12378), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n9695), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12264) );
  AOI22_X1 U15569 ( .A1(n12550), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12488), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12263) );
  NAND4_X1 U15570 ( .A1(n12266), .A2(n12265), .A3(n12264), .A4(n12263), .ZN(
        n12275) );
  AOI22_X1 U15571 ( .A1(n12526), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n9707), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12273) );
  AOI22_X1 U15572 ( .A1(n12544), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9711), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12272) );
  INV_X1 U15573 ( .A(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12268) );
  NAND2_X1 U15574 ( .A1(n9713), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n12267) );
  OAI211_X1 U15575 ( .C1(n12268), .C2(n12500), .A(n12267), .B(n12631), .ZN(
        n12269) );
  INV_X1 U15576 ( .A(n12269), .ZN(n12271) );
  AOI22_X1 U15577 ( .A1(n12527), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12373), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12270) );
  NAND4_X1 U15578 ( .A1(n12273), .A2(n12272), .A3(n12271), .A4(n12270), .ZN(
        n12274) );
  NAND2_X1 U15579 ( .A1(n12537), .A2(n12631), .ZN(n12386) );
  OAI21_X1 U15580 ( .B1(n12275), .B2(n12274), .A(n12386), .ZN(n12277) );
  AOI22_X1 U15581 ( .A1(n12456), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n21349), .ZN(n12276) );
  NAND2_X1 U15582 ( .A1(n12277), .A2(n12276), .ZN(n12278) );
  NAND2_X1 U15583 ( .A1(n12279), .A2(n12278), .ZN(n15009) );
  XNOR2_X1 U15584 ( .A(n12300), .B(n12299), .ZN(n15399) );
  AOI22_X1 U15585 ( .A1(n12378), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n9690), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12286) );
  AOI22_X1 U15586 ( .A1(n12527), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12395), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12285) );
  AOI22_X1 U15587 ( .A1(n12550), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n9707), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12284) );
  AOI22_X1 U15588 ( .A1(n9689), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12488), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12283) );
  NAND4_X1 U15589 ( .A1(n12286), .A2(n12285), .A3(n12284), .A4(n12283), .ZN(
        n12295) );
  AOI22_X1 U15590 ( .A1(n9713), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12526), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12293) );
  AOI22_X1 U15591 ( .A1(n12544), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12373), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12292) );
  INV_X1 U15592 ( .A(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12288) );
  INV_X1 U15593 ( .A(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12287) );
  OAI22_X1 U15594 ( .A1(n12502), .A2(n12288), .B1(n12500), .B2(n12287), .ZN(
        n12289) );
  INV_X1 U15595 ( .A(n12289), .ZN(n12291) );
  AOI22_X1 U15596 ( .A1(n9711), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12545), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12290) );
  NAND4_X1 U15597 ( .A1(n12293), .A2(n12292), .A3(n12291), .A4(n12290), .ZN(
        n12294) );
  NOR2_X1 U15598 ( .A1(n12295), .A2(n12294), .ZN(n12297) );
  AOI22_X1 U15599 ( .A1(n12456), .A2(P1_EAX_REG_17__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n12563), .ZN(n12296) );
  OAI21_X1 U15600 ( .B1(n12537), .B2(n12297), .A(n12296), .ZN(n12298) );
  AOI21_X1 U15601 ( .B1(n15399), .B2(n12058), .A(n12298), .ZN(n14994) );
  XNOR2_X1 U15602 ( .A(n12332), .B(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15386) );
  AOI22_X1 U15603 ( .A1(n12456), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n21349), .ZN(n12315) );
  AOI22_X1 U15604 ( .A1(n9713), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12550), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12304) );
  AOI22_X1 U15605 ( .A1(n12527), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12373), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12303) );
  AOI22_X1 U15606 ( .A1(n12483), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n12526), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12302) );
  AOI22_X1 U15607 ( .A1(n12544), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12488), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12301) );
  NAND4_X1 U15608 ( .A1(n12304), .A2(n12303), .A3(n12302), .A4(n12301), .ZN(
        n12313) );
  AOI22_X1 U15609 ( .A1(n9689), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12395), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12311) );
  INV_X1 U15610 ( .A(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12306) );
  NAND2_X1 U15611 ( .A1(n9690), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n12305) );
  OAI211_X1 U15612 ( .C1(n12306), .C2(n12500), .A(n12305), .B(n12631), .ZN(
        n12307) );
  INV_X1 U15613 ( .A(n12307), .ZN(n12310) );
  AOI22_X1 U15614 ( .A1(n9711), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(n9707), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12309) );
  AOI22_X1 U15615 ( .A1(n12378), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12545), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12308) );
  NAND4_X1 U15616 ( .A1(n12311), .A2(n12310), .A3(n12309), .A4(n12308), .ZN(
        n12312) );
  OAI21_X1 U15617 ( .B1(n12313), .B2(n12312), .A(n12386), .ZN(n12314) );
  AOI22_X1 U15618 ( .A1(n15386), .A2(n12058), .B1(n12315), .B2(n12314), .ZN(
        n14981) );
  AOI22_X1 U15619 ( .A1(n12378), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n9690), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12319) );
  AOI22_X1 U15620 ( .A1(n12483), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12527), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12318) );
  AOI22_X1 U15621 ( .A1(n12395), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12373), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12317) );
  AOI22_X1 U15622 ( .A1(n9711), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12488), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12316) );
  NAND4_X1 U15623 ( .A1(n12319), .A2(n12318), .A3(n12317), .A4(n12316), .ZN(
        n12328) );
  AOI22_X1 U15624 ( .A1(n9713), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12526), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12326) );
  AOI22_X1 U15625 ( .A1(n12550), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9707), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12325) );
  INV_X1 U15626 ( .A(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12321) );
  INV_X1 U15627 ( .A(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12320) );
  OAI22_X1 U15628 ( .A1(n9701), .A2(n12321), .B1(n12500), .B2(n12320), .ZN(
        n12322) );
  INV_X1 U15629 ( .A(n12322), .ZN(n12324) );
  AOI22_X1 U15630 ( .A1(n9689), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12545), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12323) );
  NAND4_X1 U15631 ( .A1(n12326), .A2(n12325), .A3(n12324), .A4(n12323), .ZN(
        n12327) );
  OR2_X1 U15632 ( .A1(n12328), .A2(n12327), .ZN(n12331) );
  INV_X1 U15633 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n12329) );
  INV_X1 U15634 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n15378) );
  OAI22_X1 U15635 ( .A1(n9815), .A2(n12329), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n15378), .ZN(n12330) );
  AOI21_X1 U15636 ( .B1(n12560), .B2(n12331), .A(n12330), .ZN(n12336) );
  INV_X1 U15637 ( .A(n12333), .ZN(n12334) );
  NAND2_X1 U15638 ( .A1(n12334), .A2(n15378), .ZN(n12335) );
  AND2_X1 U15639 ( .A1(n12366), .A2(n12335), .ZN(n15382) );
  MUX2_X1 U15640 ( .A(n12336), .B(n15382), .S(n12058), .Z(n14958) );
  XNOR2_X1 U15641 ( .A(n12366), .B(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15374) );
  NAND2_X1 U15642 ( .A1(n15374), .A2(n12058), .ZN(n12353) );
  AOI22_X1 U15643 ( .A1(n9690), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n12373), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12340) );
  AOI22_X1 U15644 ( .A1(n12527), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n9711), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12339) );
  AOI22_X1 U15645 ( .A1(n12544), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n9695), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12338) );
  AOI22_X1 U15646 ( .A1(n9713), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12488), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12337) );
  NAND4_X1 U15647 ( .A1(n12340), .A2(n12339), .A3(n12338), .A4(n12337), .ZN(
        n12349) );
  AOI22_X1 U15648 ( .A1(n12378), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n9707), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12347) );
  AOI22_X1 U15649 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n9689), .B1(
        n12395), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12346) );
  INV_X1 U15650 ( .A(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12342) );
  NAND2_X1 U15651 ( .A1(n12526), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n12341) );
  OAI211_X1 U15652 ( .C1(n12500), .C2(n12342), .A(n12341), .B(n12631), .ZN(
        n12343) );
  INV_X1 U15653 ( .A(n12343), .ZN(n12345) );
  AOI22_X1 U15654 ( .A1(n12483), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n12550), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12344) );
  NAND4_X1 U15655 ( .A1(n12347), .A2(n12346), .A3(n12345), .A4(n12344), .ZN(
        n12348) );
  OAI21_X1 U15656 ( .B1(n12349), .B2(n12348), .A(n12386), .ZN(n12351) );
  AOI22_X1 U15657 ( .A1(n12456), .A2(P1_EAX_REG_20__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n21349), .ZN(n12350) );
  NAND2_X1 U15658 ( .A1(n12351), .A2(n12350), .ZN(n12352) );
  NAND2_X1 U15659 ( .A1(n12353), .A2(n12352), .ZN(n14944) );
  AOI22_X1 U15660 ( .A1(n9690), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12526), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12357) );
  AOI22_X1 U15661 ( .A1(n9689), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9707), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12356) );
  AOI22_X1 U15662 ( .A1(n12483), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12550), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12355) );
  AOI22_X1 U15663 ( .A1(n9711), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12488), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12354) );
  NAND4_X1 U15664 ( .A1(n12357), .A2(n12356), .A3(n12355), .A4(n12354), .ZN(
        n12363) );
  AOI22_X1 U15665 ( .A1(n9713), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12378), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12361) );
  AOI22_X1 U15666 ( .A1(n9706), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12527), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12360) );
  AOI22_X1 U15667 ( .A1(n12544), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12373), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12359) );
  AOI22_X1 U15668 ( .A1(n12395), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12545), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12358) );
  NAND4_X1 U15669 ( .A1(n12361), .A2(n12360), .A3(n12359), .A4(n12358), .ZN(
        n12362) );
  NOR2_X1 U15670 ( .A1(n12363), .A2(n12362), .ZN(n12365) );
  AOI22_X1 U15671 ( .A1(n12456), .A2(P1_EAX_REG_21__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n21349), .ZN(n12364) );
  OAI21_X1 U15672 ( .B1(n12537), .B2(n12365), .A(n12364), .ZN(n12372) );
  INV_X1 U15673 ( .A(n12368), .ZN(n12370) );
  INV_X1 U15674 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n12369) );
  NAND2_X1 U15675 ( .A1(n12370), .A2(n12369), .ZN(n12371) );
  NAND2_X1 U15676 ( .A1(n12414), .A2(n12371), .ZN(n15363) );
  MUX2_X1 U15677 ( .A(n12372), .B(n15363), .S(n12058), .Z(n14929) );
  XNOR2_X1 U15678 ( .A(n12414), .B(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15357) );
  AOI22_X1 U15679 ( .A1(n12456), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n21349), .ZN(n12390) );
  AOI22_X1 U15680 ( .A1(n12395), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n9713), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12377) );
  AOI22_X1 U15681 ( .A1(n12483), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n9707), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12376) );
  AOI22_X1 U15682 ( .A1(n9706), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12373), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12375) );
  AOI22_X1 U15683 ( .A1(n12527), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12526), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12374) );
  NAND4_X1 U15684 ( .A1(n12377), .A2(n12376), .A3(n12375), .A4(n12374), .ZN(
        n12388) );
  AOI22_X1 U15685 ( .A1(n9689), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9690), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12385) );
  AOI22_X1 U15686 ( .A1(n9711), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12550), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12384) );
  AOI22_X1 U15687 ( .A1(n12378), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12488), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12383) );
  INV_X1 U15688 ( .A(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12380) );
  NAND2_X1 U15689 ( .A1(n11798), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n12379) );
  OAI211_X1 U15690 ( .C1(n9701), .C2(n12380), .A(n12379), .B(n12631), .ZN(
        n12381) );
  INV_X1 U15691 ( .A(n12381), .ZN(n12382) );
  NAND4_X1 U15692 ( .A1(n12385), .A2(n12384), .A3(n12383), .A4(n12382), .ZN(
        n12387) );
  OAI21_X1 U15693 ( .B1(n12388), .B2(n12387), .A(n12386), .ZN(n12389) );
  AOI22_X1 U15694 ( .A1(n15357), .A2(n12058), .B1(n12390), .B2(n12389), .ZN(
        n14915) );
  AND2_X2 U15695 ( .A1(n14913), .A2(n14915), .ZN(n14901) );
  AOI22_X1 U15696 ( .A1(n9713), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12378), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12394) );
  AOI22_X1 U15697 ( .A1(n9690), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12526), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12393) );
  AOI22_X1 U15698 ( .A1(n9711), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12488), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12392) );
  AOI22_X1 U15699 ( .A1(n9689), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12545), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12391) );
  NAND4_X1 U15700 ( .A1(n12394), .A2(n12393), .A3(n12392), .A4(n12391), .ZN(
        n12401) );
  AOI22_X1 U15701 ( .A1(n12544), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12483), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12399) );
  AOI22_X1 U15702 ( .A1(n12550), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n9707), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12398) );
  AOI22_X1 U15703 ( .A1(n9706), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n12527), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12397) );
  AOI22_X1 U15704 ( .A1(n12395), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12373), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12396) );
  NAND4_X1 U15705 ( .A1(n12399), .A2(n12398), .A3(n12397), .A4(n12396), .ZN(
        n12400) );
  NOR2_X1 U15706 ( .A1(n12401), .A2(n12400), .ZN(n12421) );
  AOI22_X1 U15707 ( .A1(n9690), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12526), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12405) );
  AOI22_X1 U15708 ( .A1(n9689), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9711), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12404) );
  AOI22_X1 U15709 ( .A1(n9706), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12527), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12403) );
  AOI22_X1 U15710 ( .A1(n12395), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12550), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12402) );
  NAND4_X1 U15711 ( .A1(n12405), .A2(n12404), .A3(n12403), .A4(n12402), .ZN(
        n12411) );
  AOI22_X1 U15712 ( .A1(n12544), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12483), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12409) );
  AOI22_X1 U15713 ( .A1(n9713), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12378), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12408) );
  AOI22_X1 U15714 ( .A1(n12545), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12488), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12407) );
  AOI22_X1 U15715 ( .A1(n9707), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12373), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12406) );
  NAND4_X1 U15716 ( .A1(n12409), .A2(n12408), .A3(n12407), .A4(n12406), .ZN(
        n12410) );
  NOR2_X1 U15717 ( .A1(n12411), .A2(n12410), .ZN(n12422) );
  XNOR2_X1 U15718 ( .A(n12421), .B(n12422), .ZN(n12413) );
  AOI22_X1 U15719 ( .A1(n12456), .A2(P1_EAX_REG_23__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n21349), .ZN(n12412) );
  OAI21_X1 U15720 ( .B1(n12537), .B2(n12413), .A(n12412), .ZN(n12420) );
  INV_X1 U15721 ( .A(n12416), .ZN(n12418) );
  INV_X1 U15722 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n12417) );
  NAND2_X1 U15723 ( .A1(n12418), .A2(n12417), .ZN(n12419) );
  NAND2_X1 U15724 ( .A1(n12440), .A2(n12419), .ZN(n15343) );
  MUX2_X1 U15725 ( .A(n12420), .B(n15343), .S(n12058), .Z(n14903) );
  NOR2_X1 U15726 ( .A1(n12422), .A2(n12421), .ZN(n12444) );
  AOI22_X1 U15727 ( .A1(n12550), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n9707), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12429) );
  AOI22_X1 U15728 ( .A1(n12395), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12373), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12428) );
  AOI22_X1 U15729 ( .A1(n9706), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n12527), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12427) );
  INV_X1 U15730 ( .A(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12424) );
  INV_X1 U15731 ( .A(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12423) );
  OAI22_X1 U15732 ( .A1(n9701), .A2(n12424), .B1(n12502), .B2(n12423), .ZN(
        n12425) );
  INV_X1 U15733 ( .A(n12425), .ZN(n12426) );
  NAND4_X1 U15734 ( .A1(n12429), .A2(n12428), .A3(n12427), .A4(n12426), .ZN(
        n12435) );
  AOI22_X1 U15735 ( .A1(n9713), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12378), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12433) );
  INV_X1 U15736 ( .A(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n21759) );
  AOI22_X1 U15737 ( .A1(n9690), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12526), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12432) );
  AOI22_X1 U15738 ( .A1(n9711), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12488), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12431) );
  AOI22_X1 U15739 ( .A1(n9689), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12545), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12430) );
  NAND4_X1 U15740 ( .A1(n12433), .A2(n12432), .A3(n12431), .A4(n12430), .ZN(
        n12434) );
  OR2_X1 U15741 ( .A1(n12435), .A2(n12434), .ZN(n12443) );
  INV_X1 U15742 ( .A(n12443), .ZN(n12436) );
  XNOR2_X1 U15743 ( .A(n12444), .B(n12436), .ZN(n12438) );
  INV_X1 U15744 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n15234) );
  INV_X1 U15745 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n15339) );
  OAI22_X1 U15746 ( .A1(n9815), .A2(n15234), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n15339), .ZN(n12437) );
  AOI21_X1 U15747 ( .B1(n12438), .B2(n12560), .A(n12437), .ZN(n12439) );
  XNOR2_X1 U15748 ( .A(n12440), .B(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15337) );
  MUX2_X1 U15749 ( .A(n12439), .B(n15337), .S(n12058), .Z(n14889) );
  INV_X1 U15750 ( .A(n12440), .ZN(n12441) );
  INV_X1 U15751 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n14879) );
  NAND2_X1 U15752 ( .A1(n9829), .A2(n14879), .ZN(n12442) );
  NAND2_X1 U15753 ( .A1(n12481), .A2(n12442), .ZN(n15331) );
  NAND2_X1 U15754 ( .A1(n12444), .A2(n12443), .ZN(n12461) );
  AOI22_X1 U15755 ( .A1(n9713), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12378), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12448) );
  AOI22_X1 U15756 ( .A1(n12527), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12395), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12447) );
  AOI22_X1 U15757 ( .A1(n12550), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n9707), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12446) );
  AOI22_X1 U15758 ( .A1(n9690), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12545), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12445) );
  NAND4_X1 U15759 ( .A1(n12448), .A2(n12447), .A3(n12446), .A4(n12445), .ZN(
        n12454) );
  AOI22_X1 U15760 ( .A1(n12483), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n9706), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12452) );
  AOI22_X1 U15761 ( .A1(n9689), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9711), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12451) );
  AOI22_X1 U15762 ( .A1(n12544), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12373), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12450) );
  AOI22_X1 U15763 ( .A1(n12526), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12488), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12449) );
  NAND4_X1 U15764 ( .A1(n12452), .A2(n12451), .A3(n12450), .A4(n12449), .ZN(
        n12453) );
  NOR2_X1 U15765 ( .A1(n12454), .A2(n12453), .ZN(n12462) );
  XNOR2_X1 U15766 ( .A(n12461), .B(n12462), .ZN(n12458) );
  AOI21_X1 U15767 ( .B1(n14879), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12455) );
  AOI21_X1 U15768 ( .B1(n12456), .B2(P1_EAX_REG_25__SCAN_IN), .A(n12455), .ZN(
        n12457) );
  OAI21_X1 U15769 ( .B1(n12458), .B2(n12537), .A(n12457), .ZN(n12459) );
  XNOR2_X1 U15770 ( .A(n12481), .B(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15324) );
  NOR2_X1 U15771 ( .A1(n12462), .A2(n12461), .ZN(n12496) );
  AOI22_X1 U15772 ( .A1(n12550), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n9707), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12469) );
  AOI22_X1 U15773 ( .A1(n12395), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12373), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12468) );
  AOI22_X1 U15774 ( .A1(n9706), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12527), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12467) );
  INV_X1 U15775 ( .A(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12463) );
  OAI22_X1 U15776 ( .A1(n9701), .A2(n12464), .B1(n12502), .B2(n12463), .ZN(
        n12465) );
  INV_X1 U15777 ( .A(n12465), .ZN(n12466) );
  NAND4_X1 U15778 ( .A1(n12469), .A2(n12468), .A3(n12467), .A4(n12466), .ZN(
        n12475) );
  AOI22_X1 U15779 ( .A1(n9713), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12378), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12473) );
  AOI22_X1 U15780 ( .A1(n9690), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12526), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12472) );
  AOI22_X1 U15781 ( .A1(n9711), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12488), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12471) );
  AOI22_X1 U15782 ( .A1(n9689), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12545), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12470) );
  NAND4_X1 U15783 ( .A1(n12473), .A2(n12472), .A3(n12471), .A4(n12470), .ZN(
        n12474) );
  OR2_X1 U15784 ( .A1(n12475), .A2(n12474), .ZN(n12495) );
  INV_X1 U15785 ( .A(n12495), .ZN(n12476) );
  XNOR2_X1 U15786 ( .A(n12496), .B(n12476), .ZN(n12479) );
  INV_X1 U15787 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n15225) );
  OAI21_X1 U15788 ( .B1(n21468), .B2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n21349), .ZN(n12477) );
  OAI21_X1 U15789 ( .B1(n9815), .B2(n15225), .A(n12477), .ZN(n12478) );
  AOI21_X1 U15790 ( .B1(n12479), .B2(n12560), .A(n12478), .ZN(n12480) );
  AOI21_X1 U15791 ( .B1(n15324), .B2(n12058), .A(n12480), .ZN(n14865) );
  INV_X1 U15792 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n15321) );
  INV_X1 U15793 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n13156) );
  OAI21_X1 U15794 ( .B1(n12481), .B2(n15321), .A(n13156), .ZN(n12482) );
  NAND2_X1 U15795 ( .A1(n12482), .A2(n12519), .ZN(n14854) );
  AOI22_X1 U15796 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n12544), .B1(
        n12483), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12487) );
  AOI22_X1 U15797 ( .A1(n9713), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12378), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12486) );
  AOI22_X1 U15798 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n9689), .B1(
        n12526), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12485) );
  AOI22_X1 U15799 ( .A1(n12395), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12550), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12484) );
  NAND4_X1 U15800 ( .A1(n12487), .A2(n12486), .A3(n12485), .A4(n12484), .ZN(
        n12494) );
  AOI22_X1 U15801 ( .A1(n9706), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n12527), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12492) );
  AOI22_X1 U15802 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n12373), .B1(
        n9707), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12491) );
  AOI22_X1 U15803 ( .A1(n9690), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n12488), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12490) );
  AOI22_X1 U15804 ( .A1(n9711), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(n9695), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12489) );
  NAND4_X1 U15805 ( .A1(n12492), .A2(n12491), .A3(n12490), .A4(n12489), .ZN(
        n12493) );
  NOR2_X1 U15806 ( .A1(n12494), .A2(n12493), .ZN(n12515) );
  NAND2_X1 U15807 ( .A1(n12496), .A2(n12495), .ZN(n12514) );
  XNOR2_X1 U15808 ( .A(n12515), .B(n12514), .ZN(n12498) );
  AOI22_X1 U15809 ( .A1(n12456), .A2(P1_EAX_REG_27__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n21349), .ZN(n12497) );
  OAI21_X1 U15810 ( .B1(n12498), .B2(n12537), .A(n12497), .ZN(n12499) );
  MUX2_X1 U15811 ( .A(n14854), .B(n12499), .S(n12631), .Z(n13152) );
  NOR2_X1 U15812 ( .A1(n12500), .A2(n12018), .ZN(n12505) );
  INV_X1 U15813 ( .A(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12501) );
  OAI22_X1 U15814 ( .A1(n9701), .A2(n12503), .B1(n12502), .B2(n12501), .ZN(
        n12504) );
  AOI211_X1 U15815 ( .C1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .C2(n12527), .A(
        n12505), .B(n12504), .ZN(n12513) );
  AOI22_X1 U15816 ( .A1(n9713), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12378), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12509) );
  AOI22_X1 U15817 ( .A1(n9690), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11837), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12508) );
  AOI22_X1 U15818 ( .A1(n9711), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12488), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12507) );
  AOI22_X1 U15819 ( .A1(n9689), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9695), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12506) );
  AND4_X1 U15820 ( .A1(n12509), .A2(n12508), .A3(n12507), .A4(n12506), .ZN(
        n12512) );
  AOI22_X1 U15821 ( .A1(n12550), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n9707), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12511) );
  AOI22_X1 U15822 ( .A1(n12395), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12373), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12510) );
  NAND4_X1 U15823 ( .A1(n12513), .A2(n12512), .A3(n12511), .A4(n12510), .ZN(
        n12534) );
  NOR2_X1 U15824 ( .A1(n12515), .A2(n12514), .ZN(n12535) );
  XOR2_X1 U15825 ( .A(n12534), .B(n12535), .Z(n12517) );
  INV_X1 U15826 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n15212) );
  INV_X1 U15827 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n21683) );
  OAI22_X1 U15828 ( .A1(n9815), .A2(n15212), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n21683), .ZN(n12516) );
  AOI21_X1 U15829 ( .B1(n12517), .B2(n12560), .A(n12516), .ZN(n12521) );
  NAND2_X1 U15830 ( .A1(n12519), .A2(n21683), .ZN(n12520) );
  MUX2_X1 U15831 ( .A(n12521), .B(n15312), .S(n12058), .Z(n14838) );
  AOI22_X1 U15832 ( .A1(n12544), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12395), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12525) );
  AOI22_X1 U15833 ( .A1(n9713), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12378), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12524) );
  AOI22_X1 U15834 ( .A1(n9690), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12488), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12523) );
  AOI22_X1 U15835 ( .A1(n9707), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11798), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12522) );
  NAND4_X1 U15836 ( .A1(n12525), .A2(n12524), .A3(n12523), .A4(n12522), .ZN(
        n12533) );
  AOI22_X1 U15837 ( .A1(n12526), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n9711), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12531) );
  AOI22_X1 U15838 ( .A1(n9689), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12550), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12530) );
  AOI22_X1 U15839 ( .A1(n9706), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12527), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12529) );
  AOI22_X1 U15840 ( .A1(n12483), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12373), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12528) );
  NAND4_X1 U15841 ( .A1(n12531), .A2(n12530), .A3(n12529), .A4(n12528), .ZN(
        n12532) );
  NOR2_X1 U15842 ( .A1(n12533), .A2(n12532), .ZN(n12543) );
  NAND2_X1 U15843 ( .A1(n12535), .A2(n12534), .ZN(n12542) );
  XNOR2_X1 U15844 ( .A(n12543), .B(n12542), .ZN(n12538) );
  AOI22_X1 U15845 ( .A1(n12456), .A2(P1_EAX_REG_29__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n21349), .ZN(n12536) );
  OAI21_X1 U15846 ( .B1(n12538), .B2(n12537), .A(n12536), .ZN(n12541) );
  OAI21_X1 U15847 ( .B1(n12540), .B2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n12566), .ZN(n15300) );
  MUX2_X1 U15848 ( .A(n12541), .B(n15300), .S(n12058), .Z(n14827) );
  NOR2_X1 U15849 ( .A1(n12543), .A2(n12542), .ZN(n12558) );
  AOI22_X1 U15850 ( .A1(n12483), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n9706), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12549) );
  AOI22_X1 U15851 ( .A1(n9713), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12378), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12548) );
  AOI22_X1 U15852 ( .A1(n12544), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12373), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12547) );
  AOI22_X1 U15853 ( .A1(n9707), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11798), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12546) );
  NAND4_X1 U15854 ( .A1(n12549), .A2(n12548), .A3(n12547), .A4(n12546), .ZN(
        n12556) );
  AOI22_X1 U15855 ( .A1(n9690), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11837), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12554) );
  AOI22_X1 U15856 ( .A1(n12527), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12395), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12553) );
  AOI22_X1 U15857 ( .A1(n9689), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12550), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12552) );
  AOI22_X1 U15858 ( .A1(n9711), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12488), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12551) );
  NAND4_X1 U15859 ( .A1(n12554), .A2(n12553), .A3(n12552), .A4(n12551), .ZN(
        n12555) );
  NOR2_X1 U15860 ( .A1(n12556), .A2(n12555), .ZN(n12557) );
  XNOR2_X1 U15861 ( .A(n12558), .B(n12557), .ZN(n12561) );
  INV_X1 U15862 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n14799) );
  INV_X1 U15863 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n14790) );
  OAI22_X1 U15864 ( .A1(n9815), .A2(n14799), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n14790), .ZN(n12559) );
  AOI21_X1 U15865 ( .B1(n12561), .B2(n12560), .A(n12559), .ZN(n12562) );
  XNOR2_X1 U15866 ( .A(n12566), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14792) );
  MUX2_X1 U15867 ( .A(n12562), .B(n14792), .S(n12058), .Z(n12852) );
  NOR2_X2 U15868 ( .A1(n14826), .A2(n12852), .ZN(n12565) );
  AOI22_X1 U15869 ( .A1(n12456), .A2(P1_EAX_REG_31__SCAN_IN), .B1(n12563), 
        .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n12564) );
  INV_X1 U15870 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n12751) );
  OAI22_X1 U15871 ( .A1(n12614), .A2(n13450), .B1(n20939), .B2(n14403), .ZN(
        n12578) );
  OR2_X1 U15872 ( .A1(n12578), .A2(n13450), .ZN(n12567) );
  XNOR2_X1 U15873 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n12585) );
  NAND2_X1 U15874 ( .A1(n21414), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12570) );
  XNOR2_X1 U15875 ( .A(n12585), .B(n12586), .ZN(n12577) );
  NAND2_X1 U15876 ( .A1(n12567), .A2(n12577), .ZN(n12580) );
  INV_X1 U15877 ( .A(n12580), .ZN(n12584) );
  NAND2_X1 U15878 ( .A1(n11736), .A2(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n12569) );
  AND2_X1 U15879 ( .A1(n12570), .A2(n12569), .ZN(n12576) );
  NAND2_X1 U15880 ( .A1(n12571), .A2(n10358), .ZN(n12572) );
  NAND2_X1 U15881 ( .A1(n12572), .A2(n13450), .ZN(n12593) );
  OAI21_X1 U15882 ( .B1(n12573), .B2(n13146), .A(n12593), .ZN(n12574) );
  NAND3_X1 U15883 ( .A1(n12574), .A2(n12594), .A3(n12576), .ZN(n12575) );
  OAI21_X1 U15884 ( .B1(n12608), .B2(n12576), .A(n12575), .ZN(n12581) );
  INV_X1 U15885 ( .A(n12581), .ZN(n12583) );
  INV_X1 U15886 ( .A(n12577), .ZN(n12625) );
  NOR2_X1 U15887 ( .A1(n12606), .A2(n12625), .ZN(n12579) );
  OAI22_X1 U15888 ( .A1(n12581), .A2(n12580), .B1(n12579), .B2(n12578), .ZN(
        n12582) );
  OAI21_X1 U15889 ( .B1(n12584), .B2(n12583), .A(n12582), .ZN(n12592) );
  NAND2_X1 U15890 ( .A1(n12586), .A2(n12585), .ZN(n12588) );
  NAND2_X1 U15891 ( .A1(n21681), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12587) );
  NAND2_X1 U15892 ( .A1(n12588), .A2(n12587), .ZN(n12598) );
  XNOR2_X1 U15893 ( .A(n12589), .B(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n12596) );
  XNOR2_X1 U15894 ( .A(n12598), .B(n12596), .ZN(n12627) );
  NAND2_X1 U15895 ( .A1(n12594), .A2(n12627), .ZN(n12590) );
  OAI211_X1 U15896 ( .C1(n12606), .C2(n12627), .A(n12590), .B(n12593), .ZN(
        n12591) );
  INV_X1 U15897 ( .A(n12593), .ZN(n12595) );
  INV_X1 U15898 ( .A(n12596), .ZN(n12597) );
  NAND2_X1 U15899 ( .A1(n12598), .A2(n12597), .ZN(n12600) );
  NAND2_X1 U15900 ( .A1(n15945), .A2(n15783), .ZN(n12599) );
  NAND2_X1 U15901 ( .A1(n12600), .A2(n12599), .ZN(n12605) );
  MUX2_X1 U15902 ( .A(n15793), .B(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .S(
        n15788), .Z(n12603) );
  NAND2_X1 U15903 ( .A1(n12605), .A2(n12603), .ZN(n12602) );
  NAND2_X1 U15904 ( .A1(n15793), .A2(n15788), .ZN(n12601) );
  NAND2_X1 U15905 ( .A1(n12602), .A2(n12601), .ZN(n12610) );
  NAND2_X1 U15906 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n12613), .ZN(
        n12611) );
  OR2_X1 U15907 ( .A1(n12610), .A2(n12611), .ZN(n12628) );
  INV_X1 U15908 ( .A(n12603), .ZN(n12604) );
  XNOR2_X1 U15909 ( .A(n12605), .B(n12604), .ZN(n12626) );
  NAND2_X1 U15910 ( .A1(n12628), .A2(n12626), .ZN(n12616) );
  NAND2_X1 U15911 ( .A1(n12606), .A2(n12616), .ZN(n12607) );
  NAND2_X1 U15912 ( .A1(n13440), .A2(n13146), .ZN(n12624) );
  NAND4_X1 U15913 ( .A1(n12628), .A2(n12627), .A3(n12626), .A4(n12625), .ZN(
        n12630) );
  NAND2_X1 U15914 ( .A1(n12630), .A2(n12629), .ZN(n13865) );
  INV_X1 U15915 ( .A(n13865), .ZN(n13858) );
  NAND3_X1 U15916 ( .A1(n13866), .A2(n20935), .A3(n13858), .ZN(n13732) );
  AND2_X2 U15917 ( .A1(n13153), .A2(n21349), .ZN(n15496) );
  INV_X1 U15918 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n21719) );
  NOR3_X1 U15919 ( .A1(n21719), .A2(P1_STATE2_REG_2__SCAN_IN), .A3(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n18049) );
  NOR2_X1 U15920 ( .A1(n12631), .A2(n18052), .ZN(n12632) );
  MUX2_X1 U15921 ( .A(n18049), .B(n12632), .S(n20939), .Z(n12633) );
  NAND2_X1 U15922 ( .A1(n15158), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n12859) );
  NAND2_X1 U15923 ( .A1(n14818), .A2(n20982), .ZN(n12761) );
  NAND2_X1 U15924 ( .A1(n10514), .A2(n12634), .ZN(n12638) );
  AOI22_X1 U15925 ( .A1(P1_EBX_REG_30__SCAN_IN), .A2(n12674), .B1(n14100), 
        .B2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12856) );
  INV_X1 U15926 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n12635) );
  OR2_X1 U15927 ( .A1(n12714), .A2(n12635), .ZN(n12637) );
  NAND2_X1 U15928 ( .A1(n12726), .A2(n12635), .ZN(n12636) );
  NAND2_X1 U15929 ( .A1(n12637), .A2(n12636), .ZN(n14144) );
  NAND2_X1 U15930 ( .A1(n14821), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12641) );
  INV_X1 U15931 ( .A(n12643), .ZN(n12644) );
  NAND2_X1 U15932 ( .A1(n12645), .A2(n12644), .ZN(n14266) );
  NAND2_X1 U15933 ( .A1(n14821), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12646) );
  OAI211_X1 U15934 ( .C1(n14100), .C2(P1_EBX_REG_2__SCAN_IN), .A(n12714), .B(
        n12646), .ZN(n12647) );
  OAI21_X1 U15935 ( .B1(n12725), .B2(P1_EBX_REG_2__SCAN_IN), .A(n12647), .ZN(
        n14265) );
  INV_X1 U15936 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n21114) );
  NAND2_X1 U15937 ( .A1(n12714), .A2(n21114), .ZN(n12651) );
  OAI211_X1 U15938 ( .C1(n14098), .C2(P1_EBX_REG_3__SCAN_IN), .A(n14821), .B(
        n12651), .ZN(n12654) );
  INV_X1 U15939 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n12652) );
  NAND2_X1 U15940 ( .A1(n12726), .A2(n12652), .ZN(n12653) );
  INV_X1 U15941 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n21004) );
  NAND2_X1 U15942 ( .A1(n12727), .A2(n21004), .ZN(n12657) );
  NAND2_X1 U15943 ( .A1(n14821), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12655) );
  OAI211_X1 U15944 ( .C1(n14098), .C2(P1_EBX_REG_4__SCAN_IN), .A(n12714), .B(
        n12655), .ZN(n12656) );
  INV_X1 U15945 ( .A(n12714), .ZN(n12658) );
  OAI21_X1 U15946 ( .B1(n12658), .B2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A(
        n14100), .ZN(n12660) );
  MUX2_X1 U15947 ( .A(n14821), .B(n12714), .S(P1_EBX_REG_5__SCAN_IN), .Z(
        n12659) );
  MUX2_X1 U15948 ( .A(n12727), .B(n12726), .S(P1_EBX_REG_6__SCAN_IN), .Z(
        n12661) );
  INV_X1 U15949 ( .A(n12661), .ZN(n12664) );
  INV_X1 U15950 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n18034) );
  INV_X1 U15951 ( .A(n12674), .ZN(n12662) );
  NAND2_X1 U15952 ( .A1(n18034), .A2(n12662), .ZN(n12663) );
  NAND2_X1 U15953 ( .A1(n12664), .A2(n12663), .ZN(n14574) );
  INV_X1 U15954 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n12665) );
  NAND2_X1 U15955 ( .A1(n12727), .A2(n12665), .ZN(n12668) );
  NAND2_X1 U15956 ( .A1(n14821), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12666) );
  OAI211_X1 U15957 ( .C1(n14098), .C2(P1_EBX_REG_8__SCAN_IN), .A(n12714), .B(
        n12666), .ZN(n12667) );
  MUX2_X1 U15958 ( .A(n14821), .B(n12714), .S(P1_EBX_REG_7__SCAN_IN), .Z(
        n12670) );
  NAND2_X1 U15959 ( .A1(n14100), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12669) );
  NAND2_X1 U15960 ( .A1(n12670), .A2(n12669), .ZN(n15201) );
  NAND2_X1 U15961 ( .A1(n15133), .A2(n15201), .ZN(n12671) );
  NOR2_X2 U15962 ( .A1(n15132), .A2(n12671), .ZN(n15134) );
  MUX2_X1 U15963 ( .A(n14821), .B(n12714), .S(P1_EBX_REG_9__SCAN_IN), .Z(
        n12673) );
  NAND2_X1 U15964 ( .A1(n14100), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12672) );
  NAND2_X1 U15965 ( .A1(n12673), .A2(n12672), .ZN(n15119) );
  MUX2_X1 U15966 ( .A(n12727), .B(n12726), .S(P1_EBX_REG_10__SCAN_IN), .Z(
        n12676) );
  NOR2_X1 U15967 ( .A1(n12674), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12675) );
  NOR2_X1 U15968 ( .A1(n12676), .A2(n12675), .ZN(n15101) );
  INV_X1 U15969 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15694) );
  NAND2_X1 U15970 ( .A1(n12714), .A2(n15694), .ZN(n12677) );
  OAI211_X1 U15971 ( .C1(n14098), .C2(P1_EBX_REG_11__SCAN_IN), .A(n14821), .B(
        n12677), .ZN(n12679) );
  INV_X1 U15972 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n15192) );
  NAND2_X1 U15973 ( .A1(n12726), .A2(n15192), .ZN(n12678) );
  MUX2_X1 U15974 ( .A(n12727), .B(n12726), .S(P1_EBX_REG_12__SCAN_IN), .Z(
        n12680) );
  INV_X1 U15975 ( .A(n12680), .ZN(n12682) );
  NAND2_X1 U15976 ( .A1(n12682), .A2(n12681), .ZN(n15072) );
  INV_X1 U15977 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15683) );
  NAND2_X1 U15978 ( .A1(n12714), .A2(n15683), .ZN(n12683) );
  OAI211_X1 U15979 ( .C1(n14098), .C2(P1_EBX_REG_13__SCAN_IN), .A(n14821), .B(
        n12683), .ZN(n12685) );
  INV_X1 U15980 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n15190) );
  NAND2_X1 U15981 ( .A1(n12726), .A2(n15190), .ZN(n12684) );
  NAND2_X1 U15982 ( .A1(n12685), .A2(n12684), .ZN(n15056) );
  INV_X1 U15983 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n15041) );
  NAND2_X1 U15984 ( .A1(n12727), .A2(n15041), .ZN(n12688) );
  NAND2_X1 U15985 ( .A1(n14821), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12686) );
  OAI211_X1 U15986 ( .C1(n14098), .C2(P1_EBX_REG_14__SCAN_IN), .A(n12714), .B(
        n12686), .ZN(n12687) );
  INV_X1 U15987 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15668) );
  NAND2_X1 U15988 ( .A1(n12714), .A2(n15668), .ZN(n12689) );
  OAI211_X1 U15989 ( .C1(n14098), .C2(P1_EBX_REG_15__SCAN_IN), .A(n14821), .B(
        n12689), .ZN(n12692) );
  INV_X1 U15990 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n12690) );
  NAND2_X1 U15991 ( .A1(n12726), .A2(n12690), .ZN(n12691) );
  NAND2_X1 U15992 ( .A1(n14821), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12693) );
  OAI211_X1 U15993 ( .C1(n14098), .C2(P1_EBX_REG_16__SCAN_IN), .A(n12714), .B(
        n12693), .ZN(n12694) );
  OAI21_X1 U15994 ( .B1(n12725), .B2(P1_EBX_REG_16__SCAN_IN), .A(n12694), .ZN(
        n15010) );
  INV_X1 U15995 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n15184) );
  NAND2_X1 U15996 ( .A1(n12727), .A2(n15184), .ZN(n12697) );
  NAND2_X1 U15997 ( .A1(n14821), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12695) );
  OAI211_X1 U15998 ( .C1(n14098), .C2(P1_EBX_REG_18__SCAN_IN), .A(n12714), .B(
        n12695), .ZN(n12696) );
  MUX2_X1 U15999 ( .A(n14821), .B(n12714), .S(P1_EBX_REG_17__SCAN_IN), .Z(
        n12699) );
  NAND2_X1 U16000 ( .A1(n14100), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n12698) );
  NAND2_X1 U16001 ( .A1(n12699), .A2(n12698), .ZN(n15001) );
  NAND2_X1 U16002 ( .A1(n14982), .A2(n15001), .ZN(n12700) );
  NOR2_X2 U16003 ( .A1(n15011), .A2(n12700), .ZN(n14984) );
  MUX2_X1 U16004 ( .A(n14821), .B(n12714), .S(P1_EBX_REG_19__SCAN_IN), .Z(
        n12702) );
  NAND2_X1 U16005 ( .A1(n14100), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12701) );
  NAND2_X1 U16006 ( .A1(n12702), .A2(n12701), .ZN(n14961) );
  NAND2_X1 U16007 ( .A1(n14984), .A2(n14961), .ZN(n14960) );
  NAND2_X1 U16008 ( .A1(n14821), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12703) );
  OAI211_X1 U16009 ( .C1(n14098), .C2(P1_EBX_REG_20__SCAN_IN), .A(n12714), .B(
        n12703), .ZN(n12704) );
  OAI21_X1 U16010 ( .B1(n12725), .B2(P1_EBX_REG_20__SCAN_IN), .A(n12704), .ZN(
        n14952) );
  OR2_X2 U16011 ( .A1(n14960), .A2(n14952), .ZN(n14954) );
  INV_X1 U16012 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n12705) );
  NAND2_X1 U16013 ( .A1(n12714), .A2(n12705), .ZN(n12706) );
  OAI211_X1 U16014 ( .C1(n14098), .C2(P1_EBX_REG_21__SCAN_IN), .A(n14821), .B(
        n12706), .ZN(n12709) );
  INV_X1 U16015 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n12707) );
  NAND2_X1 U16016 ( .A1(n12726), .A2(n12707), .ZN(n12708) );
  INV_X1 U16017 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n15180) );
  NAND2_X1 U16018 ( .A1(n12727), .A2(n15180), .ZN(n12712) );
  NAND2_X1 U16019 ( .A1(n14821), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12710) );
  OAI211_X1 U16020 ( .C1(n14098), .C2(P1_EBX_REG_22__SCAN_IN), .A(n12714), .B(
        n12710), .ZN(n12711) );
  NAND2_X1 U16021 ( .A1(n14821), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12713) );
  OAI211_X1 U16022 ( .C1(n14098), .C2(P1_EBX_REG_24__SCAN_IN), .A(n12714), .B(
        n12713), .ZN(n12715) );
  OAI21_X1 U16023 ( .B1(n12725), .B2(P1_EBX_REG_24__SCAN_IN), .A(n12715), .ZN(
        n14898) );
  MUX2_X1 U16024 ( .A(n14821), .B(n12714), .S(P1_EBX_REG_23__SCAN_IN), .Z(
        n12717) );
  NAND2_X1 U16025 ( .A1(n14100), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12716) );
  NAND2_X1 U16026 ( .A1(n12717), .A2(n12716), .ZN(n14904) );
  INV_X1 U16027 ( .A(n14904), .ZN(n12718) );
  NOR2_X1 U16028 ( .A1(n14898), .A2(n12718), .ZN(n12719) );
  INV_X1 U16029 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15558) );
  NAND2_X1 U16030 ( .A1(n12714), .A2(n15558), .ZN(n12720) );
  OAI211_X1 U16031 ( .C1(n14098), .C2(P1_EBX_REG_25__SCAN_IN), .A(n14821), .B(
        n12720), .ZN(n12722) );
  INV_X1 U16032 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n21702) );
  NAND2_X1 U16033 ( .A1(n12726), .A2(n21702), .ZN(n12721) );
  NAND2_X1 U16034 ( .A1(n14821), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12723) );
  OAI211_X1 U16035 ( .C1(n14098), .C2(P1_EBX_REG_26__SCAN_IN), .A(n12714), .B(
        n12723), .ZN(n12724) );
  OAI21_X1 U16036 ( .B1(n12725), .B2(P1_EBX_REG_26__SCAN_IN), .A(n12724), .ZN(
        n14861) );
  MUX2_X1 U16037 ( .A(n12727), .B(n12726), .S(P1_EBX_REG_28__SCAN_IN), .Z(
        n12729) );
  NOR2_X1 U16038 ( .A1(n12674), .A2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12728) );
  NOR2_X1 U16039 ( .A1(n12729), .A2(n12728), .ZN(n14843) );
  INV_X1 U16040 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15308) );
  NAND2_X1 U16041 ( .A1(n12714), .A2(n15308), .ZN(n12730) );
  OAI211_X1 U16042 ( .C1(n14098), .C2(P1_EBX_REG_27__SCAN_IN), .A(n14821), .B(
        n12730), .ZN(n12732) );
  INV_X1 U16043 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n15175) );
  NAND2_X1 U16044 ( .A1(n12726), .A2(n15175), .ZN(n12731) );
  NAND2_X1 U16045 ( .A1(n12732), .A2(n12731), .ZN(n14849) );
  NAND2_X1 U16046 ( .A1(n14843), .A2(n14849), .ZN(n12733) );
  OR2_X1 U16047 ( .A1(n12674), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12735) );
  OR2_X1 U16048 ( .A1(n14100), .A2(P1_EBX_REG_29__SCAN_IN), .ZN(n12734) );
  NAND2_X1 U16049 ( .A1(n12735), .A2(n12734), .ZN(n12854) );
  INV_X1 U16050 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n15173) );
  NAND2_X1 U16051 ( .A1(n12726), .A2(n15173), .ZN(n12736) );
  OAI21_X1 U16052 ( .B1(n12854), .B2(n11867), .A(n12736), .ZN(n14829) );
  NAND2_X1 U16053 ( .A1(n14844), .A2(n14829), .ZN(n14828) );
  MUX2_X1 U16054 ( .A(n12856), .B(n14821), .S(n14828), .Z(n12739) );
  AOI22_X1 U16055 ( .A1(P1_EBX_REG_31__SCAN_IN), .A2(n12674), .B1(n14100), 
        .B2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12738) );
  OAI21_X1 U16056 ( .B1(n14828), .B2(n12856), .A(n12738), .ZN(n12737) );
  INV_X1 U16057 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n15172) );
  OR2_X1 U16058 ( .A1(n13450), .A2(n15172), .ZN(n12746) );
  NAND2_X1 U16059 ( .A1(READY11_REG_SCAN_IN), .A2(READY1), .ZN(n21532) );
  AND2_X1 U16060 ( .A1(n21532), .A2(n21468), .ZN(n15958) );
  NOR2_X1 U16061 ( .A1(n12746), .A2(n15958), .ZN(n12740) );
  NAND2_X1 U16062 ( .A1(n12741), .A2(n21527), .ZN(n13990) );
  NAND2_X1 U16063 ( .A1(n13450), .A2(n13990), .ZN(n13425) );
  AND2_X1 U16064 ( .A1(n13425), .A2(n15958), .ZN(n12748) );
  INV_X1 U16065 ( .A(n15158), .ZN(n15153) );
  NAND2_X1 U16066 ( .A1(P1_REIP_REG_29__SCAN_IN), .A2(P1_REIP_REG_30__SCAN_IN), 
        .ZN(n12755) );
  INV_X1 U16067 ( .A(n12755), .ZN(n12745) );
  INV_X1 U16068 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n14894) );
  INV_X1 U16069 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n14939) );
  INV_X1 U16070 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n21567) );
  INV_X1 U16071 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n21557) );
  INV_X1 U16072 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n21558) );
  NAND4_X1 U16073 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(P1_REIP_REG_11__SCAN_IN), 
        .A3(P1_REIP_REG_9__SCAN_IN), .A4(P1_REIP_REG_10__SCAN_IN), .ZN(n15060)
         );
  NOR3_X1 U16074 ( .A1(n21557), .A2(n21558), .A3(n15060), .ZN(n14967) );
  AND3_X1 U16075 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(P1_REIP_REG_16__SCAN_IN), 
        .A3(P1_REIP_REG_15__SCAN_IN), .ZN(n14968) );
  NAND4_X1 U16076 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(P1_REIP_REG_3__SCAN_IN), 
        .A3(P1_REIP_REG_1__SCAN_IN), .A4(P1_REIP_REG_2__SCAN_IN), .ZN(n20961)
         );
  NAND4_X1 U16077 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(P1_REIP_REG_7__SCAN_IN), 
        .A3(P1_REIP_REG_6__SCAN_IN), .A4(P1_REIP_REG_5__SCAN_IN), .ZN(n14970)
         );
  NOR2_X1 U16078 ( .A1(n20961), .A2(n14970), .ZN(n14966) );
  NAND4_X1 U16079 ( .A1(n14967), .A2(P1_REIP_REG_18__SCAN_IN), .A3(n14968), 
        .A4(n14966), .ZN(n14963) );
  NOR2_X1 U16080 ( .A1(n21567), .A2(n14963), .ZN(n14946) );
  NAND2_X1 U16081 ( .A1(P1_REIP_REG_20__SCAN_IN), .A2(n14946), .ZN(n14916) );
  NOR2_X1 U16082 ( .A1(n14939), .A2(n14916), .ZN(n12752) );
  NAND4_X1 U16083 ( .A1(n15158), .A2(n12752), .A3(P1_REIP_REG_23__SCAN_IN), 
        .A4(P1_REIP_REG_22__SCAN_IN), .ZN(n14890) );
  NOR2_X1 U16084 ( .A1(n14894), .A2(n14890), .ZN(n14880) );
  NAND3_X1 U16085 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(P1_REIP_REG_25__SCAN_IN), 
        .A3(n14880), .ZN(n14852) );
  INV_X1 U16086 ( .A(n14852), .ZN(n12743) );
  AND2_X1 U16087 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(P1_REIP_REG_27__SCAN_IN), 
        .ZN(n12742) );
  NAND2_X1 U16088 ( .A1(n12743), .A2(n12742), .ZN(n12744) );
  NAND2_X1 U16089 ( .A1(n20970), .A2(n12744), .ZN(n14842) );
  OAI21_X1 U16090 ( .B1(n20968), .B2(n12745), .A(n14842), .ZN(n12865) );
  INV_X1 U16091 ( .A(n12746), .ZN(n12747) );
  NOR2_X1 U16092 ( .A1(n12748), .A2(n12747), .ZN(n12749) );
  NAND2_X1 U16093 ( .A1(n12750), .A2(n12749), .ZN(n21003) );
  OAI22_X1 U16094 ( .A1(n21003), .A2(n15172), .B1(n12751), .B2(n21001), .ZN(
        n12757) );
  NAND2_X1 U16095 ( .A1(n21016), .A2(n12752), .ZN(n14905) );
  NAND2_X1 U16096 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(P1_REIP_REG_22__SCAN_IN), 
        .ZN(n12753) );
  NOR2_X1 U16097 ( .A1(n14905), .A2(n12753), .ZN(n14891) );
  NAND2_X1 U16098 ( .A1(n14891), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n14878) );
  NAND2_X1 U16099 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(P1_REIP_REG_25__SCAN_IN), 
        .ZN(n12754) );
  NOR2_X1 U16100 ( .A1(n14878), .A2(n12754), .ZN(n14858) );
  NAND3_X1 U16101 ( .A1(n14858), .A2(P1_REIP_REG_27__SCAN_IN), .A3(
        P1_REIP_REG_28__SCAN_IN), .ZN(n14833) );
  NOR3_X1 U16102 ( .A1(n14833), .A2(P1_REIP_REG_31__SCAN_IN), .A3(n12755), 
        .ZN(n12756) );
  AOI211_X1 U16103 ( .C1(P1_REIP_REG_31__SCAN_IN), .C2(n12865), .A(n12757), 
        .B(n12756), .ZN(n12758) );
  NAND2_X1 U16104 ( .A1(n12761), .A2(n12760), .ZN(P1_U2809) );
  INV_X1 U16105 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n16949) );
  AOI22_X1 U16106 ( .A1(n11243), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n12768), 
        .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n12762) );
  OAI21_X1 U16107 ( .B1(n11261), .B2(n16949), .A(n12762), .ZN(n16805) );
  NAND2_X1 U16108 ( .A1(n12779), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n12765) );
  AOI22_X1 U16109 ( .A1(n11243), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n12768), 
        .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n12764) );
  NAND2_X1 U16110 ( .A1(n12779), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n12767) );
  AOI22_X1 U16111 ( .A1(n11243), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n12768), 
        .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n12766) );
  INV_X1 U16112 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n20866) );
  AOI22_X1 U16113 ( .A1(n11243), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n12768), 
        .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n12769) );
  OAI21_X1 U16114 ( .B1(n11261), .B2(n20866), .A(n12769), .ZN(n16051) );
  INV_X1 U16115 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n16906) );
  AOI22_X1 U16116 ( .A1(n11243), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n12768), 
        .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n12770) );
  OAI21_X1 U16117 ( .B1(n11261), .B2(n16906), .A(n12770), .ZN(n16035) );
  INV_X1 U16118 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n20869) );
  AOI22_X1 U16119 ( .A1(n11243), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n12768), 
        .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n12771) );
  OAI21_X1 U16120 ( .B1(n11261), .B2(n20869), .A(n12771), .ZN(n16019) );
  NAND2_X1 U16121 ( .A1(n12779), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n12773) );
  AOI22_X1 U16122 ( .A1(n11243), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n12768), 
        .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n12772) );
  AND2_X1 U16123 ( .A1(n12773), .A2(n12772), .ZN(n16005) );
  INV_X1 U16124 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n21700) );
  INV_X1 U16125 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n17162) );
  OAI22_X1 U16126 ( .A1(n12775), .A2(n21700), .B1(n12774), .B2(n17162), .ZN(
        n12776) );
  AOI21_X1 U16127 ( .B1(n12779), .B2(P2_REIP_REG_29__SCAN_IN), .A(n12776), 
        .ZN(n16001) );
  INV_X1 U16128 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n12838) );
  AOI22_X1 U16129 ( .A1(n11243), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n12768), 
        .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12778) );
  OAI21_X1 U16130 ( .B1(n11261), .B2(n12838), .A(n12778), .ZN(n12962) );
  AOI222_X1 U16131 ( .A1(n12779), .A2(P2_REIP_REG_31__SCAN_IN), .B1(n11243), 
        .B2(P2_EAX_REG_31__SCAN_IN), .C1(n12768), .C2(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12780) );
  AND2_X1 U16132 ( .A1(n11471), .A2(n17687), .ZN(n17659) );
  AND2_X1 U16133 ( .A1(n17661), .A2(n17659), .ZN(n12782) );
  AOI21_X1 U16134 ( .B1(n17651), .B2(n17653), .A(n12782), .ZN(n17459) );
  NAND2_X1 U16135 ( .A1(n12848), .A2(n12783), .ZN(n12784) );
  NAND2_X1 U16136 ( .A1(n17459), .A2(n12784), .ZN(n12785) );
  NAND2_X1 U16137 ( .A1(n13033), .A2(n16868), .ZN(n12805) );
  OR2_X1 U16138 ( .A1(n16867), .A2(n11170), .ZN(n14020) );
  NOR2_X1 U16139 ( .A1(n14020), .A2(n12786), .ZN(n12799) );
  NOR2_X1 U16140 ( .A1(P2_ADDRESS_REG_11__SCAN_IN), .A2(
        P2_ADDRESS_REG_25__SCAN_IN), .ZN(n21654) );
  NOR3_X1 U16141 ( .A1(P2_ADDRESS_REG_2__SCAN_IN), .A2(
        P2_ADDRESS_REG_1__SCAN_IN), .A3(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n12789) );
  NOR4_X1 U16142 ( .A1(P2_ADDRESS_REG_24__SCAN_IN), .A2(
        P2_ADDRESS_REG_23__SCAN_IN), .A3(P2_ADDRESS_REG_22__SCAN_IN), .A4(
        P2_ADDRESS_REG_21__SCAN_IN), .ZN(n12788) );
  NOR4_X1 U16143 ( .A1(P2_ADDRESS_REG_13__SCAN_IN), .A2(
        P2_ADDRESS_REG_27__SCAN_IN), .A3(P2_ADDRESS_REG_28__SCAN_IN), .A4(
        P2_ADDRESS_REG_26__SCAN_IN), .ZN(n12787) );
  AND4_X1 U16144 ( .A1(n21654), .A2(n12789), .A3(n12788), .A4(n12787), .ZN(
        n12795) );
  NOR4_X1 U16145 ( .A1(P2_ADDRESS_REG_16__SCAN_IN), .A2(
        P2_ADDRESS_REG_15__SCAN_IN), .A3(P2_ADDRESS_REG_14__SCAN_IN), .A4(
        P2_ADDRESS_REG_12__SCAN_IN), .ZN(n12793) );
  NOR4_X1 U16146 ( .A1(P2_ADDRESS_REG_20__SCAN_IN), .A2(
        P2_ADDRESS_REG_19__SCAN_IN), .A3(P2_ADDRESS_REG_18__SCAN_IN), .A4(
        P2_ADDRESS_REG_17__SCAN_IN), .ZN(n12792) );
  NOR4_X1 U16147 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n12791) );
  NOR4_X1 U16148 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(
        P2_ADDRESS_REG_9__SCAN_IN), .A3(P2_ADDRESS_REG_8__SCAN_IN), .A4(
        P2_ADDRESS_REG_7__SCAN_IN), .ZN(n12790) );
  AND4_X1 U16149 ( .A1(n12793), .A2(n12792), .A3(n12791), .A4(n12790), .ZN(
        n12794) );
  NAND2_X1 U16150 ( .A1(n12795), .A2(n12794), .ZN(n12796) );
  INV_X1 U16151 ( .A(n16845), .ZN(n12797) );
  INV_X1 U16152 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n18100) );
  NOR2_X1 U16153 ( .A1(n12797), .A2(n18100), .ZN(n12803) );
  INV_X1 U16154 ( .A(n16850), .ZN(n12800) );
  AOI22_X1 U16155 ( .A1(n12800), .A2(BUF2_REG_31__SCAN_IN), .B1(
        P2_EAX_REG_31__SCAN_IN), .B2(n16867), .ZN(n12801) );
  INV_X1 U16156 ( .A(n12801), .ZN(n12802) );
  NOR2_X1 U16157 ( .A1(n12803), .A2(n12802), .ZN(n12804) );
  NAND2_X1 U16158 ( .A1(n12805), .A2(n12804), .ZN(P2_U2888) );
  INV_X1 U16159 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n13034) );
  OR2_X1 U16160 ( .A1(n11385), .A2(n13034), .ZN(n12810) );
  NAND2_X1 U16161 ( .A1(n12833), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n12807) );
  NAND2_X1 U16162 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n12806) );
  OAI211_X1 U16163 ( .C1(n12821), .C2(n16949), .A(n12807), .B(n12806), .ZN(
        n12808) );
  INV_X1 U16164 ( .A(n12808), .ZN(n12809) );
  NAND2_X1 U16165 ( .A1(n12810), .A2(n12809), .ZN(n16665) );
  INV_X1 U16166 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n20862) );
  NAND2_X1 U16167 ( .A1(n12833), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n12813) );
  NAND2_X1 U16168 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n12812) );
  OAI211_X1 U16169 ( .C1(n12821), .C2(n20862), .A(n12813), .B(n12812), .ZN(
        n12814) );
  AOI21_X1 U16170 ( .B1(n12840), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n12814), .ZN(n16082) );
  INV_X1 U16171 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n20864) );
  NAND2_X1 U16172 ( .A1(n12833), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n12816) );
  NAND2_X1 U16173 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n12815) );
  OAI211_X1 U16174 ( .C1(n12821), .C2(n20864), .A(n12816), .B(n12815), .ZN(
        n12817) );
  AOI21_X1 U16175 ( .B1(n12840), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n12817), .ZN(n16063) );
  INV_X1 U16176 ( .A(n16063), .ZN(n12818) );
  NAND2_X1 U16177 ( .A1(n12833), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n12820) );
  NAND2_X1 U16178 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n12819) );
  OAI211_X1 U16179 ( .C1(n12821), .C2(n20866), .A(n12820), .B(n12819), .ZN(
        n12822) );
  AOI21_X1 U16180 ( .B1(n12840), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n12822), .ZN(n16053) );
  NOR2_X2 U16181 ( .A1(n16052), .A2(n16053), .ZN(n16020) );
  INV_X1 U16182 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n17188) );
  AOI22_X1 U16183 ( .A1(n10772), .A2(P2_REIP_REG_27__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), 
        .ZN(n12824) );
  NAND2_X1 U16184 ( .A1(n12833), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n12823) );
  OAI211_X1 U16185 ( .C1(n11385), .C2(n17188), .A(n12824), .B(n12823), .ZN(
        n16023) );
  INV_X1 U16186 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17202) );
  OR2_X1 U16187 ( .A1(n11385), .A2(n17202), .ZN(n12829) );
  NAND2_X1 U16188 ( .A1(n12833), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n12826) );
  NAND2_X1 U16189 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n12825) );
  OAI211_X1 U16190 ( .C1(n12821), .C2(n16906), .A(n12826), .B(n12825), .ZN(
        n12827) );
  INV_X1 U16191 ( .A(n12827), .ZN(n12828) );
  NAND2_X1 U16192 ( .A1(n12829), .A2(n12828), .ZN(n16036) );
  AND2_X1 U16193 ( .A1(n16023), .A2(n16036), .ZN(n12830) );
  NAND2_X1 U16194 ( .A1(n16020), .A2(n12830), .ZN(n13061) );
  INV_X1 U16195 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n12947) );
  AOI22_X1 U16196 ( .A1(n10772), .A2(P2_REIP_REG_28__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), 
        .ZN(n12831) );
  OAI21_X1 U16197 ( .B1(n12843), .B2(n12947), .A(n12831), .ZN(n12832) );
  AOI21_X1 U16198 ( .B1(n12840), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n12832), .ZN(n13063) );
  AOI22_X1 U16199 ( .A1(n10772), .A2(P2_REIP_REG_29__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n12835) );
  NAND2_X1 U16200 ( .A1(n12833), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n12834) );
  OAI211_X1 U16201 ( .C1(n11385), .C2(n17162), .A(n12835), .B(n12834), .ZN(
        n15988) );
  NAND2_X1 U16202 ( .A1(n12833), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n12837) );
  NAND2_X1 U16203 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n12836) );
  OAI211_X1 U16204 ( .C1(n12821), .C2(n12838), .A(n12837), .B(n12836), .ZN(
        n12839) );
  AOI21_X1 U16205 ( .B1(n12840), .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n12839), .ZN(n12967) );
  INV_X1 U16206 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n12972) );
  NAND2_X1 U16207 ( .A1(n12840), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n12842) );
  AOI22_X1 U16208 ( .A1(n10772), .A2(P2_REIP_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n12841) );
  OAI211_X1 U16209 ( .C1(n12843), .C2(n12972), .A(n12842), .B(n12841), .ZN(
        n12844) );
  INV_X1 U16210 ( .A(n17651), .ZN(n12847) );
  NAND2_X1 U16211 ( .A1(n12847), .A2(n17652), .ZN(n17457) );
  NAND2_X1 U16212 ( .A1(n17447), .A2(n12848), .ZN(n17478) );
  NAND2_X1 U16213 ( .A1(n17457), .A2(n17478), .ZN(n12849) );
  INV_X1 U16214 ( .A(n14806), .ZN(n12853) );
  INV_X1 U16215 ( .A(n12854), .ZN(n12855) );
  AOI22_X1 U16216 ( .A1(n14828), .A2(n11867), .B1(n12855), .B2(n14844), .ZN(
        n12857) );
  INV_X1 U16217 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n21580) );
  INV_X1 U16218 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n12858) );
  OAI21_X1 U16219 ( .B1(n14833), .B2(n21580), .A(n12858), .ZN(n12864) );
  INV_X1 U16220 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n14805) );
  OAI22_X1 U16221 ( .A1(n21003), .A2(n14805), .B1(n14790), .B2(n21001), .ZN(
        n12863) );
  INV_X1 U16222 ( .A(n12859), .ZN(n12860) );
  INV_X1 U16223 ( .A(n14792), .ZN(n12861) );
  NOR2_X1 U16224 ( .A1(n21015), .A2(n12861), .ZN(n12862) );
  AOI211_X1 U16225 ( .C1(n12865), .C2(n12864), .A(n12863), .B(n12862), .ZN(
        n12866) );
  AND2_X1 U16226 ( .A1(n17526), .A2(n20180), .ZN(n12868) );
  INV_X1 U16227 ( .A(n17658), .ZN(n17454) );
  NOR2_X1 U16228 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n17454), .ZN(n17640) );
  NAND2_X1 U16229 ( .A1(n13033), .A2(n20195), .ZN(n12960) );
  NAND2_X1 U16230 ( .A1(n12879), .A2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12881) );
  NAND2_X1 U16231 ( .A1(n12888), .A2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12891) );
  INV_X1 U16232 ( .A(n12891), .ZN(n12869) );
  NAND2_X1 U16233 ( .A1(n12869), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12893) );
  INV_X1 U16234 ( .A(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n16133) );
  INV_X1 U16235 ( .A(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n21656) );
  INV_X1 U16236 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n12924) );
  INV_X1 U16237 ( .A(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n16067) );
  INV_X1 U16238 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n12934) );
  INV_X1 U16239 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n16029) );
  INV_X1 U16240 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16875) );
  INV_X1 U16241 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n12955) );
  XNOR2_X1 U16242 ( .A(n12870), .B(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n13163) );
  NAND2_X1 U16243 ( .A1(n13163), .A2(n17703), .ZN(n12873) );
  INV_X1 U16244 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12871) );
  MUX2_X1 U16245 ( .A(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .S(P2_STATE2_REG_0__SCAN_IN), .Z(
        n17445) );
  INV_X1 U16246 ( .A(n12878), .ZN(n12876) );
  INV_X1 U16247 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12874) );
  NAND2_X1 U16248 ( .A1(n21776), .A2(n12874), .ZN(n12875) );
  NAND2_X1 U16249 ( .A1(n12876), .A2(n12875), .ZN(n17145) );
  OAI21_X1 U16250 ( .B1(n12878), .B2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n12877), .ZN(n17138) );
  NAND2_X1 U16251 ( .A1(n16309), .A2(n17138), .ZN(n20200) );
  AND2_X1 U16252 ( .A1(n12877), .A2(n17123), .ZN(n12880) );
  NOR2_X1 U16253 ( .A1(n12879), .A2(n12880), .ZN(n20201) );
  OR2_X1 U16254 ( .A1(n12879), .A2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12882) );
  AND2_X1 U16255 ( .A1(n12881), .A2(n12882), .ZN(n17113) );
  NAND2_X1 U16256 ( .A1(n12881), .A2(n12883), .ZN(n12884) );
  NAND2_X1 U16257 ( .A1(n12886), .A2(n12884), .ZN(n17101) );
  AND2_X1 U16258 ( .A1(n12886), .A2(n18059), .ZN(n12887) );
  NOR2_X1 U16259 ( .A1(n12885), .A2(n12887), .ZN(n18062) );
  NOR2_X1 U16260 ( .A1(n12885), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12889) );
  OR2_X1 U16261 ( .A1(n12888), .A2(n12889), .ZN(n17092) );
  INV_X1 U16262 ( .A(n17092), .ZN(n12890) );
  NOR2_X1 U16263 ( .A1(n16264), .A2(n12890), .ZN(n16249) );
  OR2_X1 U16264 ( .A1(n12888), .A2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12892) );
  NAND2_X1 U16265 ( .A1(n12891), .A2(n12892), .ZN(n17074) );
  NAND2_X1 U16266 ( .A1(n12891), .A2(n12894), .ZN(n12895) );
  NAND2_X1 U16267 ( .A1(n12893), .A2(n12895), .ZN(n17062) );
  NAND2_X1 U16268 ( .A1(n12893), .A2(n17048), .ZN(n12896) );
  AND2_X1 U16269 ( .A1(n12897), .A2(n12896), .ZN(n17050) );
  AND2_X1 U16270 ( .A1(n12897), .A2(n17037), .ZN(n12898) );
  NOR2_X1 U16271 ( .A1(n12900), .A2(n12898), .ZN(n17039) );
  OR2_X1 U16272 ( .A1(n12900), .A2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n12901) );
  NAND2_X1 U16273 ( .A1(n12899), .A2(n12901), .ZN(n17029) );
  AND2_X1 U16274 ( .A1(n16212), .A2(n17029), .ZN(n16187) );
  INV_X1 U16275 ( .A(n12902), .ZN(n12905) );
  NAND2_X1 U16276 ( .A1(n12899), .A2(n12903), .ZN(n12904) );
  NAND2_X1 U16277 ( .A1(n12905), .A2(n12904), .ZN(n17017) );
  NAND2_X1 U16278 ( .A1(n16187), .A2(n17017), .ZN(n16174) );
  AND2_X1 U16279 ( .A1(n12905), .A2(n17002), .ZN(n12906) );
  NOR2_X1 U16280 ( .A1(n10632), .A2(n12906), .ZN(n17004) );
  OR2_X1 U16281 ( .A1(n16174), .A2(n17004), .ZN(n16164) );
  NOR2_X1 U16282 ( .A1(n10632), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12908) );
  OR2_X1 U16283 ( .A1(n12907), .A2(n12908), .ZN(n16992) );
  INV_X1 U16284 ( .A(n16992), .ZN(n12909) );
  NOR2_X1 U16285 ( .A1(n16164), .A2(n12909), .ZN(n16143) );
  OR2_X1 U16286 ( .A1(n12907), .A2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n12911) );
  NAND2_X1 U16287 ( .A1(n12910), .A2(n12911), .ZN(n16983) );
  AND2_X1 U16288 ( .A1(n16143), .A2(n16983), .ZN(n16127) );
  NAND2_X1 U16289 ( .A1(n12910), .A2(n16133), .ZN(n12912) );
  NAND2_X1 U16290 ( .A1(n12913), .A2(n12912), .ZN(n16977) );
  NAND2_X1 U16291 ( .A1(n16127), .A2(n16977), .ZN(n16116) );
  AND2_X1 U16292 ( .A1(n12913), .A2(n16114), .ZN(n12914) );
  NOR2_X1 U16293 ( .A1(n12917), .A2(n12914), .ZN(n16117) );
  OR2_X1 U16294 ( .A1(n16116), .A2(n16117), .ZN(n12915) );
  NOR2_X1 U16295 ( .A1(n12917), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12918) );
  OR2_X1 U16296 ( .A1(n12916), .A2(n12918), .ZN(n16966) );
  INV_X1 U16297 ( .A(n16966), .ZN(n12919) );
  OR2_X1 U16298 ( .A1(n12916), .A2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12921) );
  NAND2_X1 U16299 ( .A1(n12920), .A2(n12921), .ZN(n16956) );
  NAND2_X1 U16300 ( .A1(n12920), .A2(n21656), .ZN(n12922) );
  NAND2_X1 U16301 ( .A1(n12925), .A2(n12922), .ZN(n17995) );
  NAND2_X1 U16302 ( .A1(n12923), .A2(n17995), .ZN(n16085) );
  NAND2_X1 U16303 ( .A1(n16085), .A2(n16336), .ZN(n12927) );
  NAND2_X1 U16304 ( .A1(n12925), .A2(n12924), .ZN(n12926) );
  NAND2_X1 U16305 ( .A1(n12928), .A2(n12926), .ZN(n16938) );
  AND2_X1 U16306 ( .A1(n12928), .A2(n16067), .ZN(n12929) );
  OR2_X1 U16307 ( .A1(n12929), .A2(n12931), .ZN(n16925) );
  OR2_X1 U16308 ( .A1(n12931), .A2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12932) );
  NAND2_X1 U16309 ( .A1(n12930), .A2(n12932), .ZN(n16919) );
  NAND2_X1 U16310 ( .A1(n12933), .A2(n16919), .ZN(n16039) );
  NAND2_X1 U16311 ( .A1(n12930), .A2(n12934), .ZN(n12935) );
  NAND2_X1 U16312 ( .A1(n9750), .A2(n12935), .ZN(n16907) );
  AND2_X1 U16313 ( .A1(n9750), .A2(n16029), .ZN(n12937) );
  OR2_X1 U16314 ( .A1(n12937), .A2(n12936), .ZN(n16898) );
  NAND2_X1 U16315 ( .A1(n16007), .A2(n16336), .ZN(n12940) );
  NOR2_X1 U16316 ( .A1(n12936), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12939) );
  OR2_X1 U16317 ( .A1(n12938), .A2(n12939), .ZN(n16008) );
  NAND2_X1 U16318 ( .A1(n15989), .A2(n16336), .ZN(n12942) );
  OR2_X1 U16319 ( .A1(n12938), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12941) );
  NAND2_X1 U16320 ( .A1(n9822), .A2(n12941), .ZN(n16887) );
  NAND2_X1 U16321 ( .A1(n12942), .A2(n16887), .ZN(n15991) );
  XNOR2_X1 U16322 ( .A(n9822), .B(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16877) );
  AOI21_X1 U16323 ( .B1(n15991), .B2(n16336), .A(n16877), .ZN(n12966) );
  NAND2_X1 U16324 ( .A1(n20691), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n13065) );
  NAND2_X1 U16325 ( .A1(n20742), .A2(n17703), .ZN(n12944) );
  NOR2_X2 U16326 ( .A1(n12943), .A2(n17996), .ZN(n16322) );
  NAND2_X1 U16327 ( .A1(n13010), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n12985) );
  INV_X1 U16328 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n16087) );
  NOR2_X1 U16329 ( .A1(n11012), .A2(n16087), .ZN(n12995) );
  NOR2_X1 U16330 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(P2_EBX_REG_25__SCAN_IN), 
        .ZN(n12946) );
  NAND2_X1 U16331 ( .A1(n13010), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n13006) );
  NOR2_X1 U16332 ( .A1(n11012), .A2(n12947), .ZN(n13004) );
  INV_X1 U16333 ( .A(P2_EBX_REG_29__SCAN_IN), .ZN(n12948) );
  NOR2_X1 U16334 ( .A1(n11012), .A2(n12948), .ZN(n13017) );
  NAND2_X1 U16335 ( .A1(n17661), .A2(n20180), .ZN(n13623) );
  NAND2_X1 U16336 ( .A1(n17687), .A2(n20691), .ZN(n12971) );
  NAND2_X1 U16337 ( .A1(n12971), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n12949) );
  NOR2_X1 U16338 ( .A1(n12958), .A2(n12949), .ZN(n12950) );
  NOR3_X1 U16339 ( .A1(n12970), .A2(P2_EBX_REG_30__SCAN_IN), .A3(n20192), .ZN(
        n12957) );
  AND2_X1 U16340 ( .A1(n20742), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20658) );
  NAND2_X1 U16341 ( .A1(n12951), .A2(n20658), .ZN(n17689) );
  NAND2_X1 U16342 ( .A1(n17689), .A2(n17996), .ZN(n12952) );
  NOR2_X1 U16343 ( .A1(n12952), .A2(n18058), .ZN(n12953) );
  NOR2_X1 U16344 ( .A1(n13852), .A2(n17640), .ZN(n12974) );
  AOI22_X1 U16345 ( .A1(n20190), .A2(P2_REIP_REG_31__SCAN_IN), .B1(
        P2_EBX_REG_31__SCAN_IN), .B2(n12974), .ZN(n12954) );
  OAI21_X1 U16346 ( .B1(n16178), .B2(n12955), .A(n12954), .ZN(n12956) );
  NOR2_X1 U16347 ( .A1(n12958), .A2(n12971), .ZN(n12959) );
  INV_X1 U16348 ( .A(n12961), .ZN(n12963) );
  NAND2_X1 U16349 ( .A1(n15991), .A2(n16877), .ZN(n12964) );
  AOI21_X1 U16350 ( .B1(n12964), .B2(n20204), .A(n17999), .ZN(n12965) );
  XNOR2_X2 U16351 ( .A(n15987), .B(n12967), .ZN(n16879) );
  NAND2_X1 U16352 ( .A1(n13010), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n12969) );
  NAND2_X1 U16353 ( .A1(n13020), .A2(n16348), .ZN(n12976) );
  AND3_X1 U16354 ( .A1(n13603), .A2(n12972), .A3(n12971), .ZN(n12973) );
  OR2_X2 U16355 ( .A1(n12974), .A2(n12973), .ZN(n20188) );
  AOI22_X1 U16356 ( .A1(n20190), .A2(P2_REIP_REG_30__SCAN_IN), .B1(n20188), 
        .B2(P2_EBX_REG_30__SCAN_IN), .ZN(n12975) );
  OAI211_X1 U16357 ( .C1(n16178), .C2(n16875), .A(n12976), .B(n12975), .ZN(
        n12977) );
  INV_X1 U16358 ( .A(n12977), .ZN(n12978) );
  OAI211_X1 U16359 ( .C1(n16752), .C2(n17991), .A(n12979), .B(n10633), .ZN(
        P2_U2825) );
  NAND4_X1 U16360 ( .A1(n16998), .A2(n12980), .A3(n17012), .A4(n17024), .ZN(
        n12981) );
  NOR2_X1 U16361 ( .A1(n16990), .A2(n12981), .ZN(n12983) );
  INV_X1 U16362 ( .A(n12985), .ZN(n12986) );
  NAND2_X1 U16363 ( .A1(n12987), .A2(n12986), .ZN(n12988) );
  NAND2_X1 U16364 ( .A1(n12996), .A2(n12988), .ZN(n18001) );
  OR3_X1 U16365 ( .A1(n18001), .A2(n11073), .A3(n13034), .ZN(n16934) );
  INV_X1 U16366 ( .A(n16934), .ZN(n16945) );
  AND4_X1 U16367 ( .A1(n12989), .A2(n17011), .A3(n17008), .A4(n17025), .ZN(
        n12991) );
  AND4_X1 U16368 ( .A1(n13498), .A2(n12991), .A3(n16999), .A4(n12990), .ZN(
        n12992) );
  NAND4_X1 U16369 ( .A1(n12993), .A2(n12992), .A3(n16961), .A4(n16973), .ZN(
        n16933) );
  NAND2_X1 U16370 ( .A1(n12996), .A2(n12995), .ZN(n12997) );
  NAND2_X1 U16371 ( .A1(n16065), .A2(n12997), .ZN(n13000) );
  OR2_X1 U16372 ( .A1(n13000), .A2(n11073), .ZN(n12998) );
  INV_X1 U16373 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17239) );
  XNOR2_X1 U16374 ( .A(n12998), .B(n17239), .ZN(n16936) );
  INV_X1 U16375 ( .A(n18001), .ZN(n12999) );
  AOI21_X1 U16376 ( .B1(n12999), .B2(n13049), .A(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n16946) );
  NAND2_X1 U16377 ( .A1(n13001), .A2(n13049), .ZN(n16927) );
  INV_X1 U16378 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17214) );
  NAND2_X1 U16379 ( .A1(n16927), .A2(n17214), .ZN(n16913) );
  NAND2_X1 U16380 ( .A1(n13009), .A2(n13004), .ZN(n13005) );
  NAND2_X1 U16381 ( .A1(n13018), .A2(n13005), .ZN(n16011) );
  INV_X1 U16382 ( .A(n13006), .ZN(n13007) );
  NAND2_X1 U16383 ( .A1(n10591), .A2(n13007), .ZN(n13008) );
  NAND2_X1 U16384 ( .A1(n16026), .A2(n13049), .ZN(n16894) );
  NAND2_X1 U16385 ( .A1(n16894), .A2(n17188), .ZN(n13053) );
  OAI211_X1 U16386 ( .C1(n9678), .C2(P2_EBX_REG_25__SCAN_IN), .A(n13010), .B(
        P2_EBX_REG_26__SCAN_IN), .ZN(n13011) );
  INV_X1 U16387 ( .A(n13011), .ZN(n13012) );
  OAI21_X1 U16388 ( .B1(n16043), .B2(n11073), .A(n17202), .ZN(n13046) );
  OAI211_X1 U16389 ( .C1(n13054), .C2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n13053), .B(n13046), .ZN(n13016) );
  INV_X1 U16390 ( .A(n16927), .ZN(n13013) );
  OAI21_X1 U16391 ( .B1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(n13054), .ZN(n13014) );
  XNOR2_X1 U16392 ( .A(n13018), .B(n13017), .ZN(n13021) );
  OAI21_X1 U16393 ( .B1(n13021), .B2(n11073), .A(n17162), .ZN(n16885) );
  AOI21_X1 U16394 ( .B1(n13020), .B2(n13049), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n13481) );
  AND2_X1 U16395 ( .A1(n13049), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13019) );
  INV_X1 U16396 ( .A(n13021), .ZN(n15992) );
  NAND3_X1 U16397 ( .A1(n15992), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n13049), .ZN(n16884) );
  NOR2_X1 U16398 ( .A1(n13023), .A2(n13022), .ZN(n13024) );
  XOR2_X1 U16399 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n13024), .Z(
        n13025) );
  XNOR2_X1 U16400 ( .A(n13026), .B(n13025), .ZN(n13170) );
  OR2_X1 U16401 ( .A1(n13170), .A2(n17443), .ZN(n13045) );
  NAND2_X1 U16402 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n13029) );
  NAND2_X1 U16403 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n13028) );
  AND3_X1 U16404 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n13032) );
  INV_X1 U16405 ( .A(n17240), .ZN(n17238) );
  NOR3_X1 U16406 ( .A1(n17239), .A2(n13034), .A3(n17238), .ZN(n17223) );
  AND2_X1 U16407 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17223), .ZN(
        n17199) );
  INV_X1 U16408 ( .A(n17199), .ZN(n13035) );
  NOR3_X1 U16409 ( .A1(n13035), .A2(n17214), .A3(n17237), .ZN(n17203) );
  NAND2_X1 U16410 ( .A1(n17203), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17178) );
  INV_X1 U16411 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n13057) );
  INV_X1 U16412 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n13036) );
  NOR3_X1 U16413 ( .A1(n17162), .A2(n13036), .A3(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n13037) );
  INV_X1 U16414 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n20875) );
  NOR2_X1 U16415 ( .A1(n17136), .A2(n20875), .ZN(n13161) );
  AOI21_X1 U16416 ( .B1(n17163), .B2(n13037), .A(n13161), .ZN(n13041) );
  NOR3_X1 U16417 ( .A1(n17162), .A2(n13057), .A3(n17188), .ZN(n13039) );
  NAND2_X1 U16418 ( .A1(n17326), .A2(n17199), .ZN(n17225) );
  NAND2_X1 U16419 ( .A1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n13038) );
  OAI21_X1 U16420 ( .B1(n17225), .B2(n13038), .A(n20257), .ZN(n17189) );
  OAI211_X1 U16421 ( .C1(n17419), .C2(n13039), .A(n17189), .B(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n13485) );
  NAND3_X1 U16422 ( .A1(n13485), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n20257), .ZN(n13040) );
  OAI211_X1 U16423 ( .C1(n13160), .C2(n20259), .A(n13041), .B(n13040), .ZN(
        n13042) );
  INV_X1 U16424 ( .A(n13042), .ZN(n13043) );
  NAND3_X1 U16425 ( .A1(n13045), .A2(n13044), .A3(n13043), .ZN(P2_U3015) );
  INV_X1 U16426 ( .A(n13048), .ZN(n13047) );
  NAND2_X1 U16427 ( .A1(n13047), .A2(n13046), .ZN(n16904) );
  AOI21_X1 U16428 ( .B1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n13049), .A(
        n13048), .ZN(n13051) );
  INV_X1 U16429 ( .A(n16026), .ZN(n13050) );
  NOR2_X1 U16430 ( .A1(n13051), .A2(n13050), .ZN(n13052) );
  NAND2_X1 U16431 ( .A1(n9953), .A2(n20180), .ZN(n13055) );
  NOR2_X1 U16432 ( .A1(n17668), .A2(n13055), .ZN(n13056) );
  NOR2_X1 U16433 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n17491) );
  OR2_X1 U16434 ( .A1(n20888), .A2(n17491), .ZN(n20901) );
  NAND2_X1 U16435 ( .A1(n20901), .A2(n17703), .ZN(n13064) );
  AND2_X1 U16436 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20902) );
  NAND2_X1 U16437 ( .A1(n17703), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n14037) );
  NAND2_X1 U16438 ( .A1(n14037), .A2(n13065), .ZN(n20246) );
  NAND2_X1 U16439 ( .A1(n11487), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n17177) );
  NAND2_X1 U16440 ( .A1(n20247), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n13066) );
  OAI211_X1 U16441 ( .C1(n16008), .C2(n17146), .A(n17177), .B(n13066), .ZN(
        n13067) );
  INV_X1 U16442 ( .A(n13127), .ZN(n13092) );
  NOR2_X1 U16443 ( .A1(n13092), .A2(n13070), .ZN(n13071) );
  NAND2_X1 U16444 ( .A1(n9688), .A2(n15683), .ZN(n13072) );
  INV_X1 U16445 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n21804) );
  NAND2_X1 U16446 ( .A1(n13139), .A2(n21804), .ZN(n15440) );
  NAND2_X1 U16447 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n13073) );
  NAND2_X1 U16448 ( .A1(n13139), .A2(n13073), .ZN(n15438) );
  NAND2_X1 U16449 ( .A1(n15440), .A2(n15438), .ZN(n13074) );
  INV_X1 U16450 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15677) );
  NAND2_X1 U16451 ( .A1(n9688), .A2(n15677), .ZN(n13075) );
  NAND2_X1 U16452 ( .A1(n15403), .A2(n13141), .ZN(n13079) );
  XNOR2_X1 U16453 ( .A(n9688), .B(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15406) );
  NAND2_X1 U16454 ( .A1(n9688), .A2(n15668), .ZN(n15412) );
  AND2_X1 U16455 ( .A1(n15406), .A2(n15412), .ZN(n13078) );
  NAND2_X1 U16456 ( .A1(n13089), .A2(n13084), .ZN(n13099) );
  NAND2_X1 U16457 ( .A1(n13099), .A2(n13098), .ZN(n13111) );
  NAND2_X1 U16458 ( .A1(n13111), .A2(n13109), .ZN(n13081) );
  XNOR2_X1 U16459 ( .A(n13081), .B(n13108), .ZN(n13082) );
  NAND2_X1 U16460 ( .A1(n13082), .A2(n15959), .ZN(n13083) );
  XNOR2_X1 U16461 ( .A(n13089), .B(n13084), .ZN(n13085) );
  OAI211_X1 U16462 ( .C1(n13085), .C2(n21617), .A(n11875), .B(n14403), .ZN(
        n13086) );
  INV_X1 U16463 ( .A(n13086), .ZN(n13087) );
  NAND2_X1 U16464 ( .A1(n13088), .A2(n13087), .ZN(n13095) );
  NAND2_X1 U16465 ( .A1(n13146), .A2(n11872), .ZN(n13100) );
  OAI21_X1 U16466 ( .B1(n21617), .B2(n13089), .A(n13100), .ZN(n13090) );
  INV_X1 U16467 ( .A(n13090), .ZN(n13091) );
  XNOR2_X2 U16468 ( .A(n13095), .B(n13093), .ZN(n14304) );
  INV_X1 U16469 ( .A(n13093), .ZN(n13094) );
  NAND2_X1 U16470 ( .A1(n13095), .A2(n13094), .ZN(n13096) );
  INV_X1 U16471 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n21131) );
  NAND2_X1 U16472 ( .A1(n9709), .A2(n13127), .ZN(n13104) );
  XNOR2_X1 U16473 ( .A(n13099), .B(n13098), .ZN(n13102) );
  INV_X1 U16474 ( .A(n13100), .ZN(n13101) );
  AOI21_X1 U16475 ( .B1(n13102), .B2(n15959), .A(n13101), .ZN(n13103) );
  NAND2_X1 U16476 ( .A1(n13104), .A2(n13103), .ZN(n14273) );
  NAND2_X1 U16477 ( .A1(n13105), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13106) );
  AND2_X1 U16478 ( .A1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n21104) );
  AND2_X1 U16479 ( .A1(n13109), .A2(n13108), .ZN(n13110) );
  NAND2_X1 U16480 ( .A1(n13111), .A2(n13110), .ZN(n13120) );
  XNOR2_X1 U16481 ( .A(n13120), .B(n13118), .ZN(n13112) );
  NAND2_X1 U16482 ( .A1(n13112), .A2(n15959), .ZN(n13113) );
  INV_X1 U16483 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n15737) );
  NAND2_X1 U16484 ( .A1(n13115), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13116) );
  INV_X1 U16485 ( .A(n13118), .ZN(n13119) );
  OR2_X1 U16486 ( .A1(n13120), .A2(n13119), .ZN(n13128) );
  XNOR2_X1 U16487 ( .A(n13128), .B(n13129), .ZN(n13121) );
  NAND2_X1 U16488 ( .A1(n13121), .A2(n15959), .ZN(n13122) );
  NAND2_X1 U16489 ( .A1(n13123), .A2(n13122), .ZN(n18018) );
  NAND2_X1 U16490 ( .A1(n13126), .A2(n13127), .ZN(n13134) );
  INV_X1 U16491 ( .A(n13128), .ZN(n13130) );
  NAND2_X1 U16492 ( .A1(n13130), .A2(n13129), .ZN(n13136) );
  XNOR2_X1 U16493 ( .A(n13136), .B(n13131), .ZN(n13132) );
  NAND2_X1 U16494 ( .A1(n13132), .A2(n15959), .ZN(n13133) );
  OR3_X1 U16495 ( .A1(n13136), .A2(n13135), .A3(n21617), .ZN(n13137) );
  NAND2_X1 U16496 ( .A1(n9688), .A2(n13137), .ZN(n15485) );
  OR2_X1 U16497 ( .A1(n15485), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13138) );
  INV_X1 U16498 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n21728) );
  NAND2_X1 U16499 ( .A1(n15485), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n15474) );
  INV_X1 U16500 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15658) );
  INV_X1 U16501 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15646) );
  NOR2_X1 U16502 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n13140) );
  NAND2_X1 U16503 ( .A1(n15439), .A2(n15436), .ZN(n15427) );
  XNOR2_X1 U16504 ( .A(n9688), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15384) );
  AND2_X1 U16505 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15595) );
  NAND2_X1 U16506 ( .A1(n15595), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n13464) );
  NAND3_X1 U16507 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15548) );
  NAND2_X1 U16508 ( .A1(n12705), .A2(n13142), .ZN(n13143) );
  INV_X1 U16509 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15572) );
  NAND2_X1 U16510 ( .A1(n15572), .A2(n15558), .ZN(n13144) );
  AOI21_X1 U16511 ( .B1(n11896), .B2(n13146), .A(n13145), .ZN(n13432) );
  OR2_X1 U16512 ( .A1(n13148), .A2(n11874), .ZN(n13149) );
  NAND2_X1 U16513 ( .A1(n13418), .A2(n13440), .ZN(n15950) );
  OAI21_X1 U16514 ( .B1(n13150), .B2(n13152), .A(n13151), .ZN(n15222) );
  INV_X1 U16515 ( .A(n15222), .ZN(n14851) );
  AND2_X1 U16516 ( .A1(P1_STATEBS16_REG_SCAN_IN), .A2(n21376), .ZN(n14372) );
  OR2_X1 U16517 ( .A1(n13153), .A2(n21376), .ZN(n21612) );
  NAND2_X1 U16518 ( .A1(n21612), .A2(n20939), .ZN(n13154) );
  NAND2_X1 U16519 ( .A1(n20939), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15962) );
  NAND2_X1 U16520 ( .A1(n21468), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13155) );
  NAND2_X1 U16521 ( .A1(n15962), .A2(n13155), .ZN(n14090) );
  NOR2_X1 U16522 ( .A1(n14854), .A2(n21098), .ZN(n13158) );
  NAND2_X1 U16523 ( .A1(n15496), .A2(P1_REIP_REG_27__SCAN_IN), .ZN(n15539) );
  OAI21_X1 U16524 ( .B1(n15504), .B2(n13156), .A(n15539), .ZN(n13157) );
  AOI211_X1 U16525 ( .C1(n14851), .C2(n21094), .A(n13158), .B(n13157), .ZN(
        n13159) );
  OAI21_X1 U16526 ( .B1(n15546), .B2(n20943), .A(n13159), .ZN(P1_U2972) );
  AOI21_X1 U16527 ( .B1(n20247), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n13161), .ZN(n13162) );
  OAI21_X1 U16528 ( .B1(n13163), .B2(n17146), .A(n13162), .ZN(n13164) );
  INV_X1 U16529 ( .A(n13164), .ZN(n13165) );
  OAI21_X1 U16530 ( .B1(n13166), .B2(n20256), .A(n13165), .ZN(n13167) );
  INV_X1 U16531 ( .A(n13167), .ZN(n13168) );
  NAND2_X1 U16532 ( .A1(n10628), .A2(n13171), .ZN(P2_U2983) );
  NAND2_X1 U16533 ( .A1(n13185), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n13173) );
  NAND2_X1 U16534 ( .A1(n13270), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n13172) );
  OAI211_X1 U16535 ( .C1(n9681), .C2(n18721), .A(n13173), .B(n13172), .ZN(
        n13174) );
  INV_X1 U16536 ( .A(n13174), .ZN(n13178) );
  AOI22_X1 U16537 ( .A1(n18704), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n13734), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13177) );
  AOI22_X1 U16538 ( .A1(n18706), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n18705), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13176) );
  NAND2_X1 U16539 ( .A1(n13795), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n13175) );
  NAND4_X1 U16540 ( .A1(n13178), .A2(n13177), .A3(n13176), .A4(n13175), .ZN(
        n13184) );
  AOI22_X1 U16541 ( .A1(n11543), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n14679), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n13182) );
  AOI22_X1 U16542 ( .A1(n13279), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n13278), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13181) );
  AOI22_X1 U16543 ( .A1(n14649), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n18739), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13180) );
  AOI22_X1 U16544 ( .A1(n13718), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n14680), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13179) );
  NAND4_X1 U16545 ( .A1(n13182), .A2(n13181), .A3(n13180), .A4(n13179), .ZN(
        n13183) );
  INV_X1 U16546 ( .A(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13809) );
  NAND2_X1 U16547 ( .A1(n13185), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n13187) );
  NAND2_X1 U16548 ( .A1(n13270), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n13186) );
  OAI211_X1 U16549 ( .C1(n9681), .C2(n13809), .A(n13187), .B(n13186), .ZN(
        n13188) );
  INV_X1 U16550 ( .A(n13188), .ZN(n13192) );
  AOI22_X1 U16551 ( .A1(n18704), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n13734), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13191) );
  AOI22_X1 U16552 ( .A1(n18706), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n18705), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13190) );
  NAND2_X1 U16553 ( .A1(n13795), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n13189) );
  AOI22_X1 U16554 ( .A1(n14649), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n18739), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13196) );
  AOI22_X1 U16555 ( .A1(n13279), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n13278), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13195) );
  AOI22_X1 U16556 ( .A1(n11543), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n14679), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13194) );
  AOI22_X1 U16557 ( .A1(n13718), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n14680), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13193) );
  NAND2_X4 U16558 ( .A1(n13197), .A2(n9753), .ZN(n14167) );
  INV_X1 U16559 ( .A(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13200) );
  INV_X1 U16560 ( .A(n13270), .ZN(n14335) );
  INV_X2 U16561 ( .A(n14335), .ZN(n18699) );
  NAND2_X1 U16562 ( .A1(n18699), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n13199) );
  NAND2_X1 U16563 ( .A1(n13878), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n13198) );
  OAI211_X1 U16564 ( .C1(n9681), .C2(n13200), .A(n13199), .B(n13198), .ZN(
        n13201) );
  INV_X1 U16565 ( .A(n13201), .ZN(n13205) );
  AOI22_X1 U16566 ( .A1(n18704), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n14680), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13204) );
  AOI22_X1 U16567 ( .A1(n18706), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n18705), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13203) );
  NAND2_X1 U16568 ( .A1(n13795), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n13202) );
  NAND4_X1 U16569 ( .A1(n13205), .A2(n13204), .A3(n13203), .A4(n13202), .ZN(
        n13211) );
  AOI22_X1 U16570 ( .A1(n13718), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n18736), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n13209) );
  AOI22_X1 U16571 ( .A1(n13279), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n13278), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13208) );
  AOI22_X1 U16572 ( .A1(n14649), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n9703), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13207) );
  AOI22_X1 U16573 ( .A1(n18703), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n18739), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13206) );
  NAND4_X1 U16574 ( .A1(n13209), .A2(n13208), .A3(n13207), .A4(n13206), .ZN(
        n13210) );
  INV_X1 U16575 ( .A(n13300), .ZN(n13241) );
  INV_X1 U16576 ( .A(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13214) );
  NAND2_X1 U16577 ( .A1(n9703), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n13213) );
  NAND2_X1 U16578 ( .A1(n18699), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n13212) );
  OAI211_X1 U16579 ( .C1(n18735), .C2(n13214), .A(n13213), .B(n13212), .ZN(
        n13215) );
  INV_X1 U16580 ( .A(n13215), .ZN(n13219) );
  AOI22_X1 U16581 ( .A1(n18704), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n9683), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13218) );
  AOI22_X1 U16582 ( .A1(n18706), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n18705), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13217) );
  NAND2_X1 U16583 ( .A1(n13795), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n13216) );
  NAND4_X1 U16584 ( .A1(n13219), .A2(n13218), .A3(n13217), .A4(n13216), .ZN(
        n13225) );
  AOI22_X1 U16585 ( .A1(n11543), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n14679), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n13223) );
  INV_X2 U16586 ( .A(n13819), .ZN(n18596) );
  AOI22_X1 U16587 ( .A1(n13279), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n18596), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n13222) );
  AOI22_X1 U16588 ( .A1(n14649), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n18739), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13221) );
  AOI22_X1 U16589 ( .A1(n13718), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n14680), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13220) );
  NAND4_X1 U16590 ( .A1(n13223), .A2(n13222), .A3(n13221), .A4(n13220), .ZN(
        n13224) );
  INV_X1 U16591 ( .A(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n14595) );
  NAND2_X1 U16592 ( .A1(n9683), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n13227) );
  NAND2_X1 U16593 ( .A1(n18738), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n13226) );
  OAI211_X1 U16594 ( .C1(n18735), .C2(n14595), .A(n13227), .B(n13226), .ZN(
        n13228) );
  INV_X1 U16595 ( .A(n13228), .ZN(n13233) );
  AOI22_X1 U16596 ( .A1(n18704), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n14649), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13232) );
  AOI22_X1 U16597 ( .A1(n18706), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n18705), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13231) );
  INV_X2 U16598 ( .A(n13229), .ZN(n18731) );
  NAND2_X1 U16599 ( .A1(n18731), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n13230) );
  NAND4_X1 U16600 ( .A1(n13233), .A2(n13232), .A3(n13231), .A4(n13230), .ZN(
        n13239) );
  AOI22_X1 U16601 ( .A1(n11543), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n14679), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13237) );
  AOI22_X1 U16602 ( .A1(n13279), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n18596), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n13236) );
  AOI22_X1 U16603 ( .A1(n18737), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n18739), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13235) );
  AOI22_X1 U16604 ( .A1(n9704), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n18732), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13234) );
  NAND4_X1 U16605 ( .A1(n13237), .A2(n13236), .A3(n13235), .A4(n13234), .ZN(
        n13238) );
  INV_X1 U16606 ( .A(n13306), .ZN(n13255) );
  INV_X1 U16607 ( .A(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n18678) );
  NAND2_X1 U16608 ( .A1(n9703), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n13243) );
  NAND2_X1 U16609 ( .A1(n13270), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n13242) );
  OAI211_X1 U16610 ( .C1(n18735), .C2(n18678), .A(n13243), .B(n13242), .ZN(
        n13244) );
  INV_X1 U16611 ( .A(n13244), .ZN(n13248) );
  AOI22_X1 U16612 ( .A1(n18704), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n18703), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13247) );
  AOI22_X1 U16613 ( .A1(n18706), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n18705), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13246) );
  NAND2_X1 U16614 ( .A1(n18731), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n13245) );
  NAND4_X1 U16615 ( .A1(n13248), .A2(n13247), .A3(n13246), .A4(n13245), .ZN(
        n13254) );
  AOI22_X1 U16616 ( .A1(n18736), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n14679), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n13252) );
  AOI22_X1 U16617 ( .A1(n13279), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n18596), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13251) );
  AOI22_X1 U16618 ( .A1(n14649), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n18739), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13250) );
  AOI22_X1 U16619 ( .A1(n13718), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n14680), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13249) );
  NAND4_X1 U16620 ( .A1(n13252), .A2(n13251), .A3(n13250), .A4(n13249), .ZN(
        n13253) );
  NAND2_X1 U16621 ( .A1(n13255), .A2(n13362), .ZN(n13310) );
  INV_X1 U16622 ( .A(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13258) );
  NAND2_X1 U16623 ( .A1(n9703), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n13257) );
  NAND2_X1 U16624 ( .A1(n18699), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n13256) );
  OAI211_X1 U16625 ( .C1(n18735), .C2(n13258), .A(n13257), .B(n13256), .ZN(
        n13259) );
  INV_X1 U16626 ( .A(n13259), .ZN(n13263) );
  AOI22_X1 U16627 ( .A1(n18704), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n9683), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13262) );
  AOI22_X1 U16628 ( .A1(n18706), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n18705), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n13261) );
  NAND2_X1 U16629 ( .A1(n18731), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n13260) );
  NAND4_X1 U16630 ( .A1(n13263), .A2(n13262), .A3(n13261), .A4(n13260), .ZN(
        n13269) );
  AOI22_X1 U16631 ( .A1(n18736), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n14679), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n13267) );
  INV_X1 U16632 ( .A(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n19640) );
  AOI22_X1 U16633 ( .A1(n13279), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n18596), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n13266) );
  AOI22_X1 U16634 ( .A1(n18738), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n14680), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13265) );
  AOI22_X1 U16635 ( .A1(n18740), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n18739), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13264) );
  NAND4_X1 U16636 ( .A1(n13267), .A2(n13266), .A3(n13265), .A4(n13264), .ZN(
        n13268) );
  XNOR2_X2 U16637 ( .A(n14167), .B(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n14015) );
  INV_X1 U16638 ( .A(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13752) );
  NAND2_X1 U16639 ( .A1(n9703), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n13272) );
  NAND2_X1 U16640 ( .A1(n13270), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n13271) );
  OAI211_X1 U16641 ( .C1(n9681), .C2(n13752), .A(n13272), .B(n13271), .ZN(
        n13274) );
  AOI22_X1 U16642 ( .A1(n18704), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n13734), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13277) );
  AOI22_X1 U16643 ( .A1(n18706), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n18705), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13276) );
  NAND2_X1 U16644 ( .A1(n13795), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n13275) );
  AOI22_X1 U16645 ( .A1(n11543), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n14679), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n13283) );
  AOI22_X1 U16646 ( .A1(n13279), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n13278), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n13282) );
  AOI22_X1 U16647 ( .A1(n14649), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n18739), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13281) );
  AOI22_X1 U16648 ( .A1(n13718), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n14680), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13280) );
  NAND4_X1 U16649 ( .A1(n13283), .A2(n13282), .A3(n13281), .A4(n13280), .ZN(
        n13284) );
  AND2_X1 U16650 ( .A1(n14161), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n14014) );
  NAND2_X1 U16651 ( .A1(n14015), .A2(n14014), .ZN(n14013) );
  INV_X1 U16652 ( .A(n14167), .ZN(n13285) );
  NAND2_X1 U16653 ( .A1(n13285), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13286) );
  NAND2_X1 U16654 ( .A1(n14013), .A2(n13286), .ZN(n19260) );
  XNOR2_X2 U16655 ( .A(n13368), .B(n14167), .ZN(n13287) );
  XNOR2_X1 U16656 ( .A(n13287), .B(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n19261) );
  NAND2_X1 U16657 ( .A1(n19260), .A2(n19261), .ZN(n19259) );
  INV_X1 U16658 ( .A(n13287), .ZN(n13288) );
  NAND2_X1 U16659 ( .A1(n13288), .A2(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13289) );
  INV_X1 U16660 ( .A(n13290), .ZN(n13291) );
  INV_X1 U16661 ( .A(n13366), .ZN(n14295) );
  NAND2_X1 U16662 ( .A1(n13291), .A2(n14295), .ZN(n13292) );
  NAND2_X1 U16663 ( .A1(n13300), .A2(n13292), .ZN(n13293) );
  INV_X1 U16664 ( .A(n13297), .ZN(n13298) );
  NAND2_X1 U16665 ( .A1(n13298), .A2(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13299) );
  NAND2_X2 U16666 ( .A1(n19233), .A2(n13299), .ZN(n13304) );
  INV_X1 U16667 ( .A(n13360), .ZN(n14239) );
  OAI21_X1 U16668 ( .B1(n13300), .B2(n14235), .A(n14239), .ZN(n13301) );
  NAND2_X1 U16669 ( .A1(n13306), .A2(n13301), .ZN(n13302) );
  INV_X1 U16670 ( .A(n13302), .ZN(n13303) );
  XNOR2_X1 U16671 ( .A(n13306), .B(n14243), .ZN(n13307) );
  XNOR2_X1 U16672 ( .A(n13307), .B(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n19210) );
  INV_X1 U16673 ( .A(n13307), .ZN(n13308) );
  NAND2_X1 U16674 ( .A1(n13308), .A2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13309) );
  NAND2_X1 U16675 ( .A1(n13310), .A2(n17908), .ZN(n13311) );
  NAND2_X1 U16676 ( .A1(n19030), .A2(n13311), .ZN(n13312) );
  NAND2_X2 U16677 ( .A1(n19205), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n19204) );
  INV_X1 U16678 ( .A(n13312), .ZN(n13313) );
  NAND2_X1 U16679 ( .A1(n13314), .A2(n13313), .ZN(n13315) );
  INV_X1 U16680 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17832) );
  INV_X1 U16681 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n19165) );
  INV_X1 U16682 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n19400) );
  INV_X1 U16683 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n19445) );
  NOR2_X1 U16684 ( .A1(n10263), .A2(n19445), .ZN(n19432) );
  NAND2_X1 U16685 ( .A1(n19432), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n19408) );
  NAND2_X1 U16686 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n19139), .ZN(
        n14708) );
  OAI21_X2 U16687 ( .B1(n17800), .B2(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n19030), .ZN(n19026) );
  AND2_X1 U16688 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n19110) );
  INV_X1 U16689 ( .A(n19110), .ZN(n13319) );
  OR2_X2 U16690 ( .A1(n17904), .A2(n13319), .ZN(n19063) );
  NAND2_X2 U16691 ( .A1(n19026), .A2(n19063), .ZN(n19118) );
  NAND2_X1 U16692 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n19340) );
  INV_X1 U16693 ( .A(n19340), .ZN(n13321) );
  AND3_X1 U16694 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n13320) );
  NAND2_X1 U16695 ( .A1(n13321), .A2(n13320), .ZN(n19027) );
  INV_X1 U16696 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n19035) );
  OR2_X1 U16697 ( .A1(n19027), .A2(n19035), .ZN(n17949) );
  INV_X1 U16698 ( .A(n17949), .ZN(n13322) );
  INV_X1 U16699 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n19368) );
  NAND2_X1 U16700 ( .A1(n19030), .A2(n19368), .ZN(n19116) );
  NOR2_X1 U16701 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n19116), .ZN(
        n13323) );
  INV_X1 U16702 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n19315) );
  NAND2_X1 U16703 ( .A1(n13323), .A2(n19315), .ZN(n19064) );
  NOR2_X1 U16704 ( .A1(n19064), .A2(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n19047) );
  INV_X1 U16705 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n19060) );
  NAND3_X1 U16706 ( .A1(n19047), .A2(n19035), .A3(n19060), .ZN(n13324) );
  OAI21_X1 U16707 ( .B1(n19063), .B2(n17949), .A(n13324), .ZN(n13325) );
  NAND2_X1 U16708 ( .A1(n19026), .A2(n13325), .ZN(n17791) );
  OR2_X2 U16709 ( .A1(n17791), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n17789) );
  NAND2_X1 U16710 ( .A1(n13326), .A2(n17789), .ZN(n13328) );
  MUX2_X1 U16711 ( .A(n19184), .B(n13328), .S(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(n13327) );
  INV_X1 U16712 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n19289) );
  NAND2_X1 U16713 ( .A1(n13328), .A2(n19184), .ZN(n19016) );
  AND2_X1 U16714 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17926) );
  INV_X1 U16715 ( .A(n17926), .ZN(n13329) );
  NAND2_X1 U16716 ( .A1(n19184), .A2(n13329), .ZN(n13330) );
  INV_X1 U16717 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n17937) );
  INV_X1 U16718 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17893) );
  XNOR2_X1 U16719 ( .A(n19030), .B(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n17917) );
  XNOR2_X1 U16720 ( .A(n17742), .B(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n17901) );
  INV_X1 U16721 ( .A(n13332), .ZN(n13334) );
  NAND2_X1 U16722 ( .A1(n13334), .A2(n13333), .ZN(n13346) );
  NAND2_X1 U16723 ( .A1(n13335), .A2(n13346), .ZN(n13337) );
  INV_X1 U16724 ( .A(n13350), .ZN(n13336) );
  NAND2_X1 U16725 ( .A1(n13337), .A2(n13336), .ZN(n20017) );
  INV_X1 U16726 ( .A(n20017), .ZN(n13357) );
  INV_X1 U16727 ( .A(n13338), .ZN(n13343) );
  NAND2_X1 U16728 ( .A1(n13339), .A2(n19577), .ZN(n13341) );
  NAND2_X1 U16729 ( .A1(n13341), .A2(n13340), .ZN(n13342) );
  NAND3_X1 U16730 ( .A1(n13343), .A2(n13356), .A3(n13342), .ZN(n13967) );
  INV_X1 U16731 ( .A(n13345), .ZN(n13347) );
  NAND2_X1 U16732 ( .A1(n13352), .A2(n13351), .ZN(n20168) );
  NOR2_X1 U16733 ( .A1(n13356), .A2(n19568), .ZN(n14309) );
  NOR2_X1 U16734 ( .A1(n14311), .A2(n14309), .ZN(n13976) );
  NOR2_X4 U16735 ( .A1(n19467), .A2(n20150), .ZN(n20021) );
  INV_X1 U16736 ( .A(n19141), .ZN(n19189) );
  INV_X1 U16737 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n19341) );
  NOR2_X1 U16738 ( .A1(n19340), .A2(n19341), .ZN(n19317) );
  NAND2_X1 U16739 ( .A1(n19110), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n19337) );
  INV_X1 U16740 ( .A(n19337), .ZN(n13358) );
  AND2_X1 U16741 ( .A1(n19317), .A2(n13358), .ZN(n19326) );
  NAND2_X1 U16742 ( .A1(n19326), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n19290) );
  NAND2_X1 U16743 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n19291) );
  INV_X1 U16744 ( .A(n19291), .ZN(n19296) );
  AND2_X1 U16745 ( .A1(n17926), .A2(n19296), .ZN(n17856) );
  INV_X1 U16746 ( .A(n17856), .ZN(n13359) );
  NAND2_X1 U16747 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17765) );
  INV_X1 U16748 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n17899) );
  NOR2_X1 U16749 ( .A1(n17910), .A2(n17899), .ZN(n17884) );
  OR2_X1 U16750 ( .A1(n19189), .A2(n17884), .ZN(n13391) );
  INV_X1 U16751 ( .A(n13368), .ZN(n14260) );
  NAND2_X1 U16752 ( .A1(n13369), .A2(n14260), .ZN(n13367) );
  NAND2_X1 U16753 ( .A1(n13367), .A2(n13366), .ZN(n13376) );
  NOR2_X1 U16754 ( .A1(n13376), .A2(n14235), .ZN(n13364) );
  NAND2_X1 U16755 ( .A1(n13364), .A2(n13360), .ZN(n13363) );
  NOR2_X1 U16756 ( .A1(n13363), .A2(n14243), .ZN(n13361) );
  AND2_X1 U16757 ( .A1(n13361), .A2(n18887), .ZN(n13388) );
  XNOR2_X1 U16758 ( .A(n13361), .B(n17908), .ZN(n19202) );
  XNOR2_X1 U16759 ( .A(n13363), .B(n13362), .ZN(n13382) );
  XNOR2_X1 U16760 ( .A(n13364), .B(n14239), .ZN(n13365) );
  NAND2_X1 U16761 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n13365), .ZN(
        n13381) );
  XOR2_X1 U16762 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B(n13365), .Z(
        n19225) );
  INV_X1 U16763 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n21791) );
  XNOR2_X1 U16764 ( .A(n13367), .B(n13366), .ZN(n13375) );
  XNOR2_X1 U16765 ( .A(n13375), .B(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n19252) );
  XNOR2_X1 U16766 ( .A(n13369), .B(n13368), .ZN(n13370) );
  INV_X1 U16767 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n19550) );
  OR2_X1 U16768 ( .A1(n13370), .A2(n19550), .ZN(n13374) );
  XNOR2_X1 U16769 ( .A(n13370), .B(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n19266) );
  INV_X1 U16770 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n17962) );
  AOI21_X1 U16771 ( .B1(n14167), .B2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13371) );
  MUX2_X1 U16772 ( .A(n13371), .B(n14167), .S(n14161), .Z(n13373) );
  NOR2_X1 U16773 ( .A1(n14167), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13372) );
  NOR2_X1 U16774 ( .A1(n13373), .A2(n13372), .ZN(n19265) );
  NAND2_X1 U16775 ( .A1(n19266), .A2(n19265), .ZN(n19264) );
  NAND2_X1 U16776 ( .A1(n13374), .A2(n19264), .ZN(n19251) );
  NAND2_X1 U16777 ( .A1(n19252), .A2(n19251), .ZN(n19250) );
  OAI21_X1 U16778 ( .B1(n21791), .B2(n13375), .A(n19250), .ZN(n13379) );
  XNOR2_X1 U16779 ( .A(n13376), .B(n14235), .ZN(n13378) );
  INV_X1 U16780 ( .A(n13378), .ZN(n13377) );
  NAND2_X1 U16781 ( .A1(n13379), .A2(n13377), .ZN(n13380) );
  XNOR2_X1 U16782 ( .A(n13379), .B(n13378), .ZN(n19241) );
  NAND2_X1 U16783 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n19241), .ZN(
        n19240) );
  NAND2_X1 U16784 ( .A1(n13382), .A2(n13383), .ZN(n13384) );
  NAND2_X1 U16785 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n19216), .ZN(
        n19215) );
  INV_X1 U16786 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n19485) );
  NAND2_X1 U16787 ( .A1(n13388), .A2(n13385), .ZN(n13389) );
  NAND2_X1 U16788 ( .A1(n13388), .A2(n13387), .ZN(n13386) );
  NAND2_X1 U16789 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n19188), .ZN(
        n19187) );
  NAND2_X2 U16790 ( .A1(n13389), .A2(n19187), .ZN(n19426) );
  AND2_X2 U16791 ( .A1(n17914), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n17883) );
  INV_X1 U16792 ( .A(n17883), .ZN(n13397) );
  NAND2_X1 U16793 ( .A1(n19275), .A2(n13397), .ZN(n13390) );
  NAND2_X1 U16794 ( .A1(n13391), .A2(n13390), .ZN(n17773) );
  INV_X1 U16795 ( .A(n17910), .ZN(n13392) );
  NAND2_X1 U16796 ( .A1(n19141), .A2(n13392), .ZN(n13408) );
  NOR2_X1 U16797 ( .A1(n20049), .A2(n18189), .ZN(n19239) );
  INV_X1 U16798 ( .A(n19239), .ZN(n19145) );
  NOR2_X1 U16799 ( .A1(n20049), .A2(n20151), .ZN(n13393) );
  INV_X1 U16800 ( .A(n13393), .ZN(n19552) );
  NAND2_X1 U16801 ( .A1(n20134), .A2(n19552), .ZN(n20158) );
  NAND2_X1 U16802 ( .A1(n20156), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n19098) );
  INV_X1 U16803 ( .A(n19082), .ZN(n19053) );
  NOR2_X1 U16804 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n19053), .ZN(
        n17756) );
  OAI21_X1 U16805 ( .B1(n19067), .B2(n17756), .A(n18219), .ZN(n13407) );
  INV_X1 U16806 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n17981) );
  NAND2_X1 U16807 ( .A1(n17981), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n14744) );
  OAI21_X1 U16808 ( .B1(n13393), .B2(n20154), .A(n14744), .ZN(n19563) );
  NAND2_X1 U16809 ( .A1(n17753), .A2(n19945), .ZN(n13398) );
  INV_X1 U16810 ( .A(n19098), .ZN(n19143) );
  NAND2_X1 U16811 ( .A1(n19143), .A2(n13394), .ZN(n13395) );
  AND2_X1 U16812 ( .A1(n13398), .A2(n13395), .ZN(n13396) );
  AND2_X1 U16813 ( .A1(n19271), .A2(n13396), .ZN(n17758) );
  INV_X1 U16814 ( .A(n17758), .ZN(n13405) );
  NAND3_X1 U16815 ( .A1(n19275), .A2(n17914), .A3(n13397), .ZN(n13403) );
  INV_X1 U16816 ( .A(n13398), .ZN(n13401) );
  INV_X1 U16817 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n13399) );
  NOR2_X1 U16818 ( .A1(n19442), .A2(n13399), .ZN(n17897) );
  AOI21_X1 U16819 ( .B1(n13401), .B2(n13400), .A(n17897), .ZN(n13402) );
  NAND2_X1 U16820 ( .A1(n13403), .A2(n13402), .ZN(n13404) );
  AOI21_X1 U16821 ( .B1(n13405), .B2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n13404), .ZN(n13406) );
  OAI211_X1 U16822 ( .C1(n17884), .C2(n13408), .A(n13407), .B(n13406), .ZN(
        n13409) );
  NOR2_X1 U16823 ( .A1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15531) );
  NAND2_X1 U16824 ( .A1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15530) );
  INV_X1 U16825 ( .A(n15530), .ZN(n13412) );
  AND2_X1 U16826 ( .A1(n10056), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13413) );
  NAND2_X1 U16827 ( .A1(n15302), .A2(n13413), .ZN(n13414) );
  INV_X1 U16828 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14808) );
  NAND2_X1 U16829 ( .A1(n13415), .A2(n14808), .ZN(n13416) );
  INV_X1 U16830 ( .A(n14793), .ZN(n13477) );
  NOR2_X1 U16831 ( .A1(n11896), .A2(n13450), .ZN(n13443) );
  INV_X1 U16832 ( .A(n13443), .ZN(n13422) );
  INV_X1 U16833 ( .A(n13866), .ZN(n13420) );
  NAND2_X1 U16834 ( .A1(n11895), .A2(n13417), .ZN(n13457) );
  NAND2_X1 U16835 ( .A1(n13418), .A2(n13457), .ZN(n13419) );
  NAND2_X1 U16836 ( .A1(n13420), .A2(n13419), .ZN(n13938) );
  INV_X1 U16837 ( .A(n13990), .ZN(n18008) );
  NOR2_X1 U16838 ( .A1(n21533), .A2(n13865), .ZN(n13936) );
  OAI211_X1 U16839 ( .C1(n13450), .C2(n18008), .A(n13936), .B(n14381), .ZN(
        n13421) );
  OAI211_X1 U16840 ( .C1(n15971), .C2(n13422), .A(n13938), .B(n13421), .ZN(
        n13423) );
  NAND2_X1 U16841 ( .A1(n13423), .A2(n20935), .ZN(n13430) );
  NAND2_X1 U16842 ( .A1(n13425), .A2(n21532), .ZN(n13426) );
  OAI211_X1 U16843 ( .C1(n13424), .C2(n13426), .A(n10358), .B(n14136), .ZN(
        n13427) );
  NAND2_X1 U16844 ( .A1(n13427), .A2(n11871), .ZN(n13428) );
  NAND2_X1 U16845 ( .A1(n13432), .A2(n15147), .ZN(n14433) );
  AND2_X1 U16846 ( .A1(n15950), .A2(n14433), .ZN(n13863) );
  INV_X1 U16847 ( .A(n13433), .ZN(n13434) );
  OAI211_X1 U16848 ( .C1(n13435), .C2(n13431), .A(n13863), .B(n13434), .ZN(
        n13436) );
  INV_X1 U16849 ( .A(n13424), .ZN(n15960) );
  NAND2_X1 U16850 ( .A1(n15960), .A2(n15959), .ZN(n13988) );
  OAI21_X1 U16851 ( .B1(n13431), .B2(n11874), .A(n13988), .ZN(n13438) );
  NAND2_X1 U16852 ( .A1(n15496), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n14789) );
  OR2_X1 U16853 ( .A1(n13440), .A2(n13439), .ZN(n13442) );
  AND2_X1 U16854 ( .A1(n13442), .A2(n13441), .ZN(n13453) );
  NAND2_X1 U16855 ( .A1(n13453), .A2(n13443), .ZN(n14434) );
  INV_X1 U16856 ( .A(n14434), .ZN(n13444) );
  AND2_X1 U16857 ( .A1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n15748) );
  AND2_X1 U16858 ( .A1(n15748), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n15722) );
  AND2_X1 U16859 ( .A1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15723) );
  NAND2_X1 U16860 ( .A1(n15722), .A2(n15723), .ZN(n15705) );
  NOR2_X1 U16861 ( .A1(n15705), .A2(n15694), .ZN(n15689) );
  INV_X1 U16862 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n21118) );
  INV_X1 U16863 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n21144) );
  OAI21_X1 U16864 ( .B1(n21118), .B2(n21144), .A(n21131), .ZN(n21100) );
  AND2_X1 U16865 ( .A1(n21104), .A2(n21100), .ZN(n13445) );
  NAND2_X1 U16866 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n13445), .ZN(
        n15738) );
  NOR2_X1 U16867 ( .A1(n15738), .A2(n21804), .ZN(n13446) );
  AND2_X1 U16868 ( .A1(n15689), .A2(n13446), .ZN(n15587) );
  AND2_X1 U16869 ( .A1(n15587), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n13468) );
  INV_X1 U16870 ( .A(n13468), .ZN(n13447) );
  OR2_X1 U16871 ( .A1(n21117), .A2(n13447), .ZN(n13462) );
  OAI21_X1 U16872 ( .B1(n14136), .B2(n10358), .A(n14381), .ZN(n13449) );
  OAI21_X1 U16873 ( .B1(n11907), .B2(n13450), .A(n13449), .ZN(n13451) );
  INV_X1 U16874 ( .A(n13451), .ZN(n13452) );
  OAI211_X1 U16875 ( .C1(n13454), .C2(n14821), .A(n13453), .B(n13452), .ZN(
        n13455) );
  INV_X1 U16876 ( .A(n13455), .ZN(n13458) );
  NAND2_X1 U16877 ( .A1(n12623), .A2(n15147), .ZN(n13456) );
  OAI211_X1 U16878 ( .C1(n13448), .C2(n10358), .A(n13948), .B(n13459), .ZN(
        n13460) );
  AND2_X1 U16879 ( .A1(n13866), .A2(n10514), .ZN(n15937) );
  NAND2_X1 U16880 ( .A1(n15611), .A2(n21118), .ZN(n21136) );
  NAND2_X1 U16881 ( .A1(n21121), .A2(n21136), .ZN(n21116) );
  INV_X1 U16882 ( .A(n21116), .ZN(n15693) );
  INV_X1 U16883 ( .A(n21104), .ZN(n13461) );
  NAND2_X1 U16884 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n21101) );
  NOR2_X1 U16885 ( .A1(n13461), .A2(n21101), .ZN(n15741) );
  NAND2_X1 U16886 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n15741), .ZN(
        n15717) );
  NOR2_X1 U16887 ( .A1(n15705), .A2(n15717), .ZN(n15692) );
  NAND3_X1 U16888 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(n15692), .ZN(n15592) );
  NOR2_X1 U16889 ( .A1(n15683), .A2(n15592), .ZN(n13467) );
  NAND2_X1 U16890 ( .A1(n15693), .A2(n13467), .ZN(n15566) );
  NAND2_X1 U16891 ( .A1(n13462), .A2(n15566), .ZN(n15676) );
  INV_X1 U16892 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15637) );
  NAND4_X1 U16893 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A4(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15635) );
  NOR2_X1 U16894 ( .A1(n15637), .A2(n15635), .ZN(n13466) );
  NAND2_X1 U16895 ( .A1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n13466), .ZN(
        n13463) );
  NOR2_X1 U16896 ( .A1(n13464), .A2(n13463), .ZN(n13465) );
  NAND2_X1 U16897 ( .A1(n15676), .A2(n13465), .ZN(n15569) );
  INV_X1 U16898 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15547) );
  INV_X1 U16899 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15303) );
  NOR3_X1 U16900 ( .A1(n15540), .A2(n15530), .A3(n15303), .ZN(n15515) );
  INV_X1 U16901 ( .A(n21137), .ZN(n13476) );
  NAND2_X1 U16902 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n13475) );
  INV_X1 U16903 ( .A(n13466), .ZN(n15594) );
  NAND2_X1 U16904 ( .A1(n15614), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n13474) );
  NOR2_X1 U16905 ( .A1(n15742), .A2(n13467), .ZN(n13473) );
  NOR2_X1 U16906 ( .A1(n21117), .A2(n13468), .ZN(n13472) );
  OR2_X1 U16907 ( .A1(n15589), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13471) );
  NOR2_X1 U16908 ( .A1(n21137), .A2(n21119), .ZN(n15718) );
  AOI21_X1 U16909 ( .B1(n15627), .B2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n15718), .ZN(n15603) );
  OAI21_X1 U16910 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n21117), .A(
        n15579), .ZN(n15567) );
  AOI21_X1 U16911 ( .B1(n15548), .B2(n21137), .A(n15567), .ZN(n15557) );
  NAND2_X1 U16912 ( .A1(n15557), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15554) );
  NAND2_X1 U16913 ( .A1(n15579), .A2(n13476), .ZN(n15528) );
  OAI211_X1 U16914 ( .C1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n13476), .A(
        n15521), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15513) );
  NAND2_X1 U16915 ( .A1(n13478), .A2(n16884), .ZN(n13483) );
  INV_X1 U16916 ( .A(n13479), .ZN(n13480) );
  NOR2_X1 U16917 ( .A1(n13481), .A2(n13480), .ZN(n13482) );
  XNOR2_X1 U16918 ( .A(n13483), .B(n13482), .ZN(n16883) );
  OR2_X1 U16919 ( .A1(n16883), .A2(n17443), .ZN(n13495) );
  INV_X1 U16920 ( .A(n17163), .ZN(n13484) );
  NOR2_X1 U16921 ( .A1(n13484), .A2(n17162), .ZN(n13486) );
  OAI21_X1 U16922 ( .B1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n13486), .A(
        n13485), .ZN(n13487) );
  INV_X1 U16923 ( .A(n13487), .ZN(n13489) );
  NAND2_X1 U16924 ( .A1(n11487), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n16874) );
  INV_X1 U16925 ( .A(n16874), .ZN(n13488) );
  OAI21_X1 U16926 ( .B1(n16752), .B2(n18091), .A(n13490), .ZN(n13491) );
  INV_X1 U16927 ( .A(n13491), .ZN(n13494) );
  NOR2_X1 U16928 ( .A1(n16879), .A2(n20259), .ZN(n13492) );
  NAND3_X1 U16929 ( .A1(n13495), .A2(n13494), .A3(n13493), .ZN(P2_U3016) );
  NAND2_X1 U16930 ( .A1(n13496), .A2(n16974), .ZN(n13500) );
  NAND2_X1 U16931 ( .A1(n13498), .A2(n13497), .ZN(n13499) );
  INV_X1 U16932 ( .A(n16102), .ZN(n13502) );
  AOI21_X1 U16933 ( .B1(n13503), .B2(n13501), .A(n13502), .ZN(n14770) );
  NAND2_X1 U16934 ( .A1(n16117), .A2(n18063), .ZN(n13504) );
  NAND2_X1 U16935 ( .A1(n11487), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n14776) );
  OAI211_X1 U16936 ( .C1(n16114), .C2(n18060), .A(n13504), .B(n14776), .ZN(
        n13505) );
  NAND2_X1 U16937 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n17285) );
  INV_X1 U16938 ( .A(n17285), .ZN(n13507) );
  NOR4_X1 U16939 ( .A1(P1_ADDRESS_REG_16__SCAN_IN), .A2(
        P1_ADDRESS_REG_14__SCAN_IN), .A3(P1_ADDRESS_REG_13__SCAN_IN), .A4(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n13511) );
  NOR4_X1 U16940 ( .A1(P1_ADDRESS_REG_20__SCAN_IN), .A2(
        P1_ADDRESS_REG_19__SCAN_IN), .A3(P1_ADDRESS_REG_15__SCAN_IN), .A4(
        P1_ADDRESS_REG_17__SCAN_IN), .ZN(n13510) );
  NOR4_X1 U16941 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n13509) );
  NOR4_X1 U16942 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_7__SCAN_IN), .A3(P1_ADDRESS_REG_9__SCAN_IN), .A4(
        P1_ADDRESS_REG_8__SCAN_IN), .ZN(n13508) );
  AND4_X1 U16943 ( .A1(n13511), .A2(n13510), .A3(n13509), .A4(n13508), .ZN(
        n13516) );
  NOR4_X1 U16944 ( .A1(P1_ADDRESS_REG_2__SCAN_IN), .A2(
        P1_ADDRESS_REG_1__SCAN_IN), .A3(P1_ADDRESS_REG_28__SCAN_IN), .A4(
        P1_ADDRESS_REG_18__SCAN_IN), .ZN(n13514) );
  NOR4_X1 U16945 ( .A1(P1_ADDRESS_REG_24__SCAN_IN), .A2(
        P1_ADDRESS_REG_23__SCAN_IN), .A3(P1_ADDRESS_REG_22__SCAN_IN), .A4(
        P1_ADDRESS_REG_21__SCAN_IN), .ZN(n13513) );
  NOR4_X1 U16946 ( .A1(P1_ADDRESS_REG_12__SCAN_IN), .A2(
        P1_ADDRESS_REG_25__SCAN_IN), .A3(P1_ADDRESS_REG_27__SCAN_IN), .A4(
        P1_ADDRESS_REG_26__SCAN_IN), .ZN(n13512) );
  INV_X1 U16947 ( .A(P1_ADDRESS_REG_0__SCAN_IN), .ZN(n21542) );
  AND4_X1 U16948 ( .A1(n13514), .A2(n13513), .A3(n13512), .A4(n21542), .ZN(
        n13515) );
  NAND2_X1 U16949 ( .A1(n13516), .A2(n13515), .ZN(n13517) );
  INV_X1 U16950 ( .A(P1_M_IO_N_REG_SCAN_IN), .ZN(n21689) );
  INV_X1 U16951 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n21884) );
  NOR4_X1 U16952 ( .A1(P1_BE_N_REG_0__SCAN_IN), .A2(P1_BE_N_REG_1__SCAN_IN), 
        .A3(n21689), .A4(n21884), .ZN(n13519) );
  NOR4_X1 U16953 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_3__SCAN_IN), 
        .A3(P1_D_C_N_REG_SCAN_IN), .A4(P1_ADS_N_REG_SCAN_IN), .ZN(n13518) );
  NAND3_X1 U16954 ( .A1(n15223), .A2(n13519), .A3(n13518), .ZN(U214) );
  NOR2_X1 U16955 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(P2_BE_N_REG_1__SCAN_IN), 
        .ZN(n13521) );
  NOR4_X1 U16956 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n13520) );
  NAND4_X1 U16957 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(P2_W_R_N_REG_SCAN_IN), 
        .A3(n13521), .A4(n13520), .ZN(n13522) );
  NOR2_X1 U16958 ( .A1(n12798), .A2(n13522), .ZN(n18099) );
  NAND2_X1 U16959 ( .A1(n18099), .A2(U214), .ZN(U212) );
  NAND2_X1 U16960 ( .A1(n16322), .A2(n16218), .ZN(n16221) );
  AOI21_X1 U16961 ( .B1(n17050), .B2(n13523), .A(n16221), .ZN(n13538) );
  NOR2_X1 U16962 ( .A1(n16351), .A2(n11424), .ZN(n13524) );
  AOI211_X1 U16963 ( .C1(P2_EBX_REG_11__SCAN_IN), .C2(n20188), .A(n11487), .B(
        n13524), .ZN(n13525) );
  OAI21_X1 U16964 ( .B1(n17048), .B2(n16178), .A(n13525), .ZN(n13537) );
  OAI21_X1 U16965 ( .B1(n9782), .B2(n13527), .A(n13526), .ZN(n17366) );
  INV_X1 U16966 ( .A(n13528), .ZN(n13529) );
  OAI22_X1 U16967 ( .A1(n17366), .A2(n17991), .B1(n13529), .B2(n20192), .ZN(
        n13536) );
  INV_X1 U16968 ( .A(n17050), .ZN(n13534) );
  NAND2_X1 U16969 ( .A1(n13531), .A2(n13532), .ZN(n13533) );
  NAND2_X1 U16970 ( .A1(n13530), .A2(n13533), .ZN(n17370) );
  OAI22_X1 U16971 ( .A1(n16210), .A2(n13534), .B1(n17370), .B2(n20196), .ZN(
        n13535) );
  INV_X1 U16972 ( .A(n14051), .ZN(n20273) );
  MUX2_X1 U16973 ( .A(n14774), .B(n20273), .S(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .Z(n13547) );
  OAI21_X1 U16974 ( .B1(n13541), .B2(n13540), .A(n13539), .ZN(n16344) );
  OAI21_X1 U16975 ( .B1(n16349), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13924), .ZN(n20250) );
  OAI22_X1 U16976 ( .A1(n18091), .A2(n16344), .B1(n17443), .B2(n20250), .ZN(
        n13546) );
  OAI21_X1 U16977 ( .B1(n13543), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13542), .ZN(n20255) );
  NAND2_X1 U16978 ( .A1(n20280), .A2(n10091), .ZN(n13544) );
  NAND2_X1 U16979 ( .A1(n18058), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n20253) );
  OAI211_X1 U16980 ( .C1(n20255), .C2(n20290), .A(n13544), .B(n20253), .ZN(
        n13545) );
  OR3_X1 U16981 ( .A1(n13547), .A2(n13546), .A3(n13545), .ZN(P2_U3046) );
  NOR2_X1 U16982 ( .A1(n17920), .A2(n17917), .ZN(n13551) );
  INV_X1 U16983 ( .A(n13548), .ZN(n17775) );
  NAND2_X1 U16984 ( .A1(n17775), .A2(n19184), .ZN(n13550) );
  INV_X1 U16985 ( .A(n17917), .ZN(n13549) );
  AOI21_X1 U16986 ( .B1(n13550), .B2(n10490), .A(n13549), .ZN(n17909) );
  AOI211_X1 U16987 ( .C1(n13551), .C2(n13550), .A(n19109), .B(n17909), .ZN(
        n13573) );
  INV_X1 U16988 ( .A(n19043), .ZN(n13552) );
  NAND2_X1 U16989 ( .A1(n19141), .A2(n13552), .ZN(n13555) );
  NAND2_X1 U16990 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n19032), .ZN(
        n17943) );
  INV_X1 U16991 ( .A(n17943), .ZN(n13553) );
  NAND2_X1 U16992 ( .A1(n19275), .A2(n13553), .ZN(n13554) );
  NAND2_X1 U16993 ( .A1(n13555), .A2(n13554), .ZN(n17794) );
  AND2_X1 U16994 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n13556) );
  NAND2_X1 U16995 ( .A1(n17794), .A2(n13556), .ZN(n19010) );
  OR2_X1 U16996 ( .A1(n19010), .A2(n19289), .ZN(n17785) );
  NOR3_X1 U16997 ( .A1(n17785), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        n17937), .ZN(n13572) );
  NAND2_X1 U16998 ( .A1(n19141), .A2(n17925), .ZN(n13558) );
  NAND2_X1 U16999 ( .A1(n19275), .A2(n17929), .ZN(n13557) );
  AND2_X1 U17000 ( .A1(n13558), .A2(n13557), .ZN(n19009) );
  AND2_X1 U17001 ( .A1(n19009), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17784) );
  NOR2_X1 U17002 ( .A1(n19141), .A2(n19275), .ZN(n19087) );
  NOR3_X1 U17003 ( .A1(n17784), .A2(n19087), .A3(n17893), .ZN(n13571) );
  NAND2_X1 U17004 ( .A1(n19082), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13559) );
  OAI211_X1 U17005 ( .C1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A(n17778), .B(n13560), .ZN(n13569) );
  INV_X1 U17006 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n13561) );
  NAND2_X1 U17007 ( .A1(n19082), .A2(n13561), .ZN(n19000) );
  OAI21_X1 U17008 ( .B1(n13562), .B2(n19098), .A(n19271), .ZN(n13564) );
  NOR2_X1 U17009 ( .A1(n17778), .A2(n19145), .ZN(n13563) );
  NOR2_X1 U17010 ( .A1(n13564), .A2(n13563), .ZN(n19004) );
  NAND2_X1 U17011 ( .A1(n19000), .A2(n19004), .ZN(n17780) );
  INV_X1 U17012 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n13565) );
  NOR2_X1 U17013 ( .A1(n19442), .A2(n13565), .ZN(n17918) );
  NOR2_X1 U17014 ( .A1(n19159), .A2(n13566), .ZN(n13567) );
  AOI211_X1 U17015 ( .C1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .C2(n17780), .A(
        n17918), .B(n13567), .ZN(n13568) );
  OAI21_X1 U17016 ( .B1(n19148), .B2(n13569), .A(n13568), .ZN(n13570) );
  OR4_X1 U17017 ( .A1(n13573), .A2(n13572), .A3(n13571), .A4(n13570), .ZN(
        P3_U2802) );
  AND2_X1 U17018 ( .A1(n20742), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n17695) );
  NAND2_X1 U17019 ( .A1(n20819), .A2(n17695), .ZN(n17690) );
  NAND2_X1 U17020 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n20911) );
  INV_X1 U17021 ( .A(n20911), .ZN(n17515) );
  AND2_X1 U17022 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n17515), .ZN(n17688) );
  NOR2_X1 U17023 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n13575) );
  NOR3_X1 U17024 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(P2_STATEBS16_REG_SCAN_IN), .ZN(n13574) );
  NOR3_X1 U17025 ( .A1(n17688), .A2(n13575), .A3(n13574), .ZN(n13576) );
  AND2_X1 U17026 ( .A1(n17690), .A2(n13576), .ZN(P2_U3178) );
  NOR2_X1 U17027 ( .A1(n20939), .A2(n18052), .ZN(n13579) );
  NOR4_X1 U17028 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n21533), .A3(n20939), 
        .A4(n18052), .ZN(n13577) );
  AOI21_X1 U17029 ( .B1(n13578), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n13577), 
        .ZN(n18048) );
  OAI21_X1 U17030 ( .B1(n13579), .B2(n21349), .A(n18048), .ZN(P1_U3163) );
  NOR4_X1 U17031 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_11__SCAN_IN), .A3(P2_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_14__SCAN_IN), .ZN(n13589) );
  NOR4_X1 U17032 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_7__SCAN_IN), .A3(P2_DATAWIDTH_REG_8__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_9__SCAN_IN), .ZN(n13588) );
  AOI211_X1 U17033 ( .C1(P2_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_0__SCAN_IN), .A(P2_DATAWIDTH_REG_3__SCAN_IN), .B(
        P2_DATAWIDTH_REG_5__SCAN_IN), .ZN(n13580) );
  INV_X1 U17034 ( .A(P2_DATAWIDTH_REG_12__SCAN_IN), .ZN(n21883) );
  INV_X1 U17035 ( .A(P2_DATAWIDTH_REG_4__SCAN_IN), .ZN(n21766) );
  NAND3_X1 U17036 ( .A1(n13580), .A2(n21883), .A3(n21766), .ZN(n13586) );
  NOR4_X1 U17037 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_20__SCAN_IN), .A3(P2_DATAWIDTH_REG_21__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_22__SCAN_IN), .ZN(n13584) );
  NOR4_X1 U17038 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_16__SCAN_IN), .A3(P2_DATAWIDTH_REG_17__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_18__SCAN_IN), .ZN(n13583) );
  NOR4_X1 U17039 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n13582) );
  NOR4_X1 U17040 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_24__SCAN_IN), .A3(P2_DATAWIDTH_REG_25__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_26__SCAN_IN), .ZN(n13581) );
  NAND4_X1 U17041 ( .A1(n13584), .A2(n13583), .A3(n13582), .A4(n13581), .ZN(
        n13585) );
  NOR4_X1 U17042 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_2__SCAN_IN), .A3(n13586), .A4(n13585), .ZN(n13587) );
  NAND3_X1 U17043 ( .A1(n13589), .A2(n13588), .A3(n13587), .ZN(n13593) );
  INV_X1 U17044 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n13590) );
  NOR2_X1 U17045 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n13593), .ZN(n13594) );
  AOI22_X1 U17046 ( .A1(n13593), .A2(n13590), .B1(n13594), .B2(n20183), .ZN(
        P2_U2820) );
  INV_X1 U17047 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n13591) );
  INV_X1 U17048 ( .A(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n21711) );
  INV_X1 U17049 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20883) );
  NAND3_X1 U17050 ( .A1(n21711), .A2(n20883), .A3(n20183), .ZN(n13592) );
  AOI22_X1 U17051 ( .A1(n13593), .A2(n13591), .B1(n13594), .B2(n13592), .ZN(
        P2_U2821) );
  INV_X1 U17052 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n13596) );
  INV_X1 U17053 ( .A(n13593), .ZN(n20185) );
  OR2_X1 U17054 ( .A1(n13593), .A2(n13592), .ZN(n13595) );
  NAND2_X1 U17055 ( .A1(n13594), .A2(n20883), .ZN(n20187) );
  OAI211_X1 U17056 ( .C1(n13596), .C2(n20185), .A(n13595), .B(n20187), .ZN(
        P2_U2823) );
  NOR2_X1 U17057 ( .A1(n17986), .A2(n17696), .ZN(n13851) );
  NAND2_X1 U17058 ( .A1(n13851), .A2(n17654), .ZN(n20197) );
  INV_X1 U17059 ( .A(n20197), .ZN(n13599) );
  INV_X1 U17060 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n13598) );
  AND2_X1 U17061 ( .A1(n20888), .A2(n11386), .ZN(n13597) );
  NOR2_X1 U17062 ( .A1(n13603), .A2(n13597), .ZN(n13621) );
  OAI21_X1 U17063 ( .B1(n13599), .B2(n13598), .A(n13621), .ZN(P2_U2814) );
  INV_X1 U17064 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n13922) );
  AND2_X1 U17065 ( .A1(n17984), .A2(n17687), .ZN(n13600) );
  INV_X1 U17066 ( .A(BUF2_REG_8__SCAN_IN), .ZN(n18884) );
  NAND2_X1 U17067 ( .A1(n13676), .A2(BUF1_REG_8__SCAN_IN), .ZN(n13601) );
  OAI21_X1 U17068 ( .B1(n13676), .B2(n18884), .A(n13601), .ZN(n16792) );
  NAND2_X1 U17069 ( .A1(n13677), .A2(n16792), .ZN(n13609) );
  NAND2_X1 U17070 ( .A1(n17984), .A2(n20819), .ZN(n13602) );
  NAND2_X2 U17071 ( .A1(n13603), .A2(n13602), .ZN(n13685) );
  NAND2_X1 U17072 ( .A1(n13685), .A2(P2_UWORD_REG_8__SCAN_IN), .ZN(n13604) );
  OAI211_X1 U17073 ( .C1(n13852), .C2(n13922), .A(n13609), .B(n13604), .ZN(
        P2_U2960) );
  INV_X1 U17074 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n13917) );
  INV_X1 U17075 ( .A(BUF2_REG_14__SCAN_IN), .ZN(n13606) );
  NAND2_X1 U17076 ( .A1(n13676), .A2(BUF1_REG_14__SCAN_IN), .ZN(n13605) );
  OAI21_X1 U17077 ( .B1(n13676), .B2(n13606), .A(n13605), .ZN(n16745) );
  NAND2_X1 U17078 ( .A1(n13677), .A2(n16745), .ZN(n13613) );
  NAND2_X1 U17079 ( .A1(n13685), .A2(P2_UWORD_REG_14__SCAN_IN), .ZN(n13607) );
  OAI211_X1 U17080 ( .C1(n13852), .C2(n13917), .A(n13613), .B(n13607), .ZN(
        P2_U2966) );
  INV_X1 U17081 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n20229) );
  NAND2_X1 U17082 ( .A1(n13685), .A2(P2_LWORD_REG_8__SCAN_IN), .ZN(n13608) );
  OAI211_X1 U17083 ( .C1(n13852), .C2(n20229), .A(n13609), .B(n13608), .ZN(
        P2_U2975) );
  INV_X1 U17084 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n13919) );
  INV_X1 U17085 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n18807) );
  NAND2_X1 U17086 ( .A1(n13676), .A2(BUF1_REG_12__SCAN_IN), .ZN(n13610) );
  OAI21_X1 U17087 ( .B1(n13676), .B2(n18807), .A(n13610), .ZN(n16764) );
  NAND2_X1 U17088 ( .A1(n13677), .A2(n16764), .ZN(n13615) );
  NAND2_X1 U17089 ( .A1(n13685), .A2(P2_UWORD_REG_12__SCAN_IN), .ZN(n13611) );
  OAI211_X1 U17090 ( .C1(n13852), .C2(n13919), .A(n13615), .B(n13611), .ZN(
        P2_U2964) );
  INV_X1 U17091 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n20217) );
  NAND2_X1 U17092 ( .A1(n13685), .A2(P2_LWORD_REG_14__SCAN_IN), .ZN(n13612) );
  OAI211_X1 U17093 ( .C1(n13852), .C2(n20217), .A(n13613), .B(n13612), .ZN(
        P2_U2981) );
  INV_X1 U17094 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n20221) );
  NAND2_X1 U17095 ( .A1(n13685), .A2(P2_LWORD_REG_12__SCAN_IN), .ZN(n13614) );
  OAI211_X1 U17096 ( .C1(n13852), .C2(n20221), .A(n13615), .B(n13614), .ZN(
        P2_U2979) );
  INV_X1 U17097 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n20225) );
  INV_X1 U17098 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n18816) );
  NAND2_X1 U17099 ( .A1(n17525), .A2(BUF1_REG_10__SCAN_IN), .ZN(n13616) );
  OAI21_X1 U17100 ( .B1(n13676), .B2(n18816), .A(n13616), .ZN(n16778) );
  NAND2_X1 U17101 ( .A1(n13677), .A2(n16778), .ZN(n13619) );
  NAND2_X1 U17102 ( .A1(n13685), .A2(P2_LWORD_REG_10__SCAN_IN), .ZN(n13617) );
  OAI211_X1 U17103 ( .C1(n13852), .C2(n20225), .A(n13619), .B(n13617), .ZN(
        P2_U2977) );
  INV_X1 U17104 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n13915) );
  NAND2_X1 U17105 ( .A1(n13685), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n13618) );
  OAI211_X1 U17106 ( .C1(n13852), .C2(n13915), .A(n13619), .B(n13618), .ZN(
        P2_U2962) );
  INV_X1 U17107 ( .A(P2_READREQUEST_REG_SCAN_IN), .ZN(n13620) );
  NAND3_X1 U17108 ( .A1(n13621), .A2(n20197), .A3(n13620), .ZN(n13622) );
  OAI21_X1 U17109 ( .B1(n13623), .B2(n11471), .A(n13622), .ZN(n13624) );
  INV_X1 U17110 ( .A(n13624), .ZN(P2_U3612) );
  INV_X1 U17111 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n13629) );
  INV_X1 U17112 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n13628) );
  INV_X1 U17113 ( .A(n13685), .ZN(n13627) );
  INV_X1 U17114 ( .A(n13677), .ZN(n13626) );
  INV_X1 U17115 ( .A(BUF2_REG_15__SCAN_IN), .ZN(n13625) );
  INV_X1 U17116 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n14046) );
  MUX2_X1 U17117 ( .A(n13625), .B(n14046), .S(n17525), .Z(n14762) );
  OAI222_X1 U17118 ( .A1(n13852), .A2(n13629), .B1(n13628), .B2(n13627), .C1(
        n13626), .C2(n14762), .ZN(P2_U2982) );
  INV_X1 U17119 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n20178) );
  INV_X1 U17120 ( .A(n17491), .ZN(n17983) );
  INV_X1 U17121 ( .A(n17695), .ZN(n13630) );
  OAI22_X1 U17122 ( .A1(n15982), .A2(n20178), .B1(n17983), .B2(n13630), .ZN(
        P2_U2816) );
  AOI22_X1 U17123 ( .A1(n9676), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n13685), .B2(
        P2_UWORD_REG_1__SCAN_IN), .ZN(n13633) );
  INV_X1 U17124 ( .A(BUF2_REG_1__SCAN_IN), .ZN(n13632) );
  NAND2_X1 U17125 ( .A1(n13676), .A2(BUF1_REG_1__SCAN_IN), .ZN(n13631) );
  OAI21_X1 U17126 ( .B1(n13676), .B2(n13632), .A(n13631), .ZN(n17558) );
  NAND2_X1 U17127 ( .A1(n13677), .A2(n17558), .ZN(n13661) );
  NAND2_X1 U17128 ( .A1(n13633), .A2(n13661), .ZN(P2_U2953) );
  AOI22_X1 U17129 ( .A1(n9676), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n13685), .B2(
        P2_UWORD_REG_6__SCAN_IN), .ZN(n13636) );
  INV_X1 U17130 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n13635) );
  NAND2_X1 U17131 ( .A1(n17525), .A2(BUF1_REG_6__SCAN_IN), .ZN(n13634) );
  OAI21_X1 U17132 ( .B1(n17525), .B2(n13635), .A(n13634), .ZN(n17536) );
  NAND2_X1 U17133 ( .A1(n13677), .A2(n17536), .ZN(n13672) );
  NAND2_X1 U17134 ( .A1(n13636), .A2(n13672), .ZN(P2_U2958) );
  AOI22_X1 U17135 ( .A1(n9676), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n13685), .B2(
        P2_UWORD_REG_0__SCAN_IN), .ZN(n13638) );
  INV_X1 U17136 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n14163) );
  NAND2_X1 U17137 ( .A1(n13676), .A2(BUF1_REG_0__SCAN_IN), .ZN(n13637) );
  OAI21_X1 U17138 ( .B1(n17525), .B2(n14163), .A(n13637), .ZN(n17524) );
  NAND2_X1 U17139 ( .A1(n13677), .A2(n17524), .ZN(n13668) );
  NAND2_X1 U17140 ( .A1(n13638), .A2(n13668), .ZN(P2_U2952) );
  AOI22_X1 U17141 ( .A1(n9676), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n13685), .B2(
        P2_LWORD_REG_7__SCAN_IN), .ZN(n13641) );
  INV_X1 U17142 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n13640) );
  NAND2_X1 U17143 ( .A1(n13676), .A2(BUF1_REG_7__SCAN_IN), .ZN(n13639) );
  OAI21_X1 U17144 ( .B1(n17525), .B2(n13640), .A(n13639), .ZN(n17587) );
  NAND2_X1 U17145 ( .A1(n13677), .A2(n17587), .ZN(n13681) );
  NAND2_X1 U17146 ( .A1(n13641), .A2(n13681), .ZN(P2_U2974) );
  AOI22_X1 U17147 ( .A1(n9676), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n13685), .B2(
        P2_LWORD_REG_5__SCAN_IN), .ZN(n13644) );
  INV_X1 U17148 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n13643) );
  NAND2_X1 U17149 ( .A1(n17525), .A2(BUF1_REG_5__SCAN_IN), .ZN(n13642) );
  OAI21_X1 U17150 ( .B1(n13676), .B2(n13643), .A(n13642), .ZN(n17531) );
  NAND2_X1 U17151 ( .A1(n13677), .A2(n17531), .ZN(n13657) );
  NAND2_X1 U17152 ( .A1(n13644), .A2(n13657), .ZN(P2_U2972) );
  AOI22_X1 U17153 ( .A1(n9676), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n13685), .B2(
        P2_UWORD_REG_9__SCAN_IN), .ZN(n13647) );
  INV_X1 U17154 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n13646) );
  NAND2_X1 U17155 ( .A1(n17525), .A2(BUF1_REG_9__SCAN_IN), .ZN(n13645) );
  OAI21_X1 U17156 ( .B1(n13676), .B2(n13646), .A(n13645), .ZN(n16785) );
  NAND2_X1 U17157 ( .A1(n13677), .A2(n16785), .ZN(n13666) );
  NAND2_X1 U17158 ( .A1(n13647), .A2(n13666), .ZN(P2_U2961) );
  AOI22_X1 U17159 ( .A1(n9676), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n13685), .B2(
        P2_LWORD_REG_4__SCAN_IN), .ZN(n13650) );
  INV_X1 U17160 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n13649) );
  NAND2_X1 U17161 ( .A1(n13676), .A2(BUF1_REG_4__SCAN_IN), .ZN(n13648) );
  OAI21_X1 U17162 ( .B1(n17525), .B2(n13649), .A(n13648), .ZN(n17574) );
  NAND2_X1 U17163 ( .A1(n13677), .A2(n17574), .ZN(n13683) );
  NAND2_X1 U17164 ( .A1(n13650), .A2(n13683), .ZN(P2_U2971) );
  AOI22_X1 U17165 ( .A1(n9676), .A2(P2_EAX_REG_3__SCAN_IN), .B1(n13685), .B2(
        P2_LWORD_REG_3__SCAN_IN), .ZN(n13653) );
  INV_X1 U17166 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n13652) );
  NAND2_X1 U17167 ( .A1(n13676), .A2(BUF1_REG_3__SCAN_IN), .ZN(n13651) );
  OAI21_X1 U17168 ( .B1(n17525), .B2(n13652), .A(n13651), .ZN(n17569) );
  NAND2_X1 U17169 ( .A1(n13677), .A2(n17569), .ZN(n13687) );
  NAND2_X1 U17170 ( .A1(n13653), .A2(n13687), .ZN(P2_U2970) );
  AOI22_X1 U17171 ( .A1(n9676), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n13685), .B2(
        P2_LWORD_REG_2__SCAN_IN), .ZN(n13656) );
  INV_X1 U17172 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n13655) );
  NAND2_X1 U17173 ( .A1(n17525), .A2(BUF1_REG_2__SCAN_IN), .ZN(n13654) );
  OAI21_X1 U17174 ( .B1(n17525), .B2(n13655), .A(n13654), .ZN(n17563) );
  NAND2_X1 U17175 ( .A1(n13677), .A2(n17563), .ZN(n13659) );
  NAND2_X1 U17176 ( .A1(n13656), .A2(n13659), .ZN(P2_U2969) );
  AOI22_X1 U17177 ( .A1(n9676), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n13685), .B2(
        P2_UWORD_REG_5__SCAN_IN), .ZN(n13658) );
  NAND2_X1 U17178 ( .A1(n13658), .A2(n13657), .ZN(P2_U2957) );
  AOI22_X1 U17179 ( .A1(n9676), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n13685), .B2(
        P2_UWORD_REG_2__SCAN_IN), .ZN(n13660) );
  NAND2_X1 U17180 ( .A1(n13660), .A2(n13659), .ZN(P2_U2954) );
  AOI22_X1 U17181 ( .A1(n9676), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n13685), .B2(
        P2_LWORD_REG_1__SCAN_IN), .ZN(n13662) );
  NAND2_X1 U17182 ( .A1(n13662), .A2(n13661), .ZN(P2_U2968) );
  AOI22_X1 U17183 ( .A1(n9676), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n13685), .B2(
        P2_LWORD_REG_11__SCAN_IN), .ZN(n13665) );
  INV_X1 U17184 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n13664) );
  NAND2_X1 U17185 ( .A1(n13676), .A2(BUF1_REG_11__SCAN_IN), .ZN(n13663) );
  OAI21_X1 U17186 ( .B1(n13676), .B2(n13664), .A(n13663), .ZN(n16772) );
  NAND2_X1 U17187 ( .A1(n13677), .A2(n16772), .ZN(n13670) );
  NAND2_X1 U17188 ( .A1(n13665), .A2(n13670), .ZN(P2_U2978) );
  AOI22_X1 U17189 ( .A1(n9676), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n13685), .B2(
        P2_LWORD_REG_9__SCAN_IN), .ZN(n13667) );
  NAND2_X1 U17190 ( .A1(n13667), .A2(n13666), .ZN(P2_U2976) );
  AOI22_X1 U17191 ( .A1(n9676), .A2(P2_EAX_REG_0__SCAN_IN), .B1(n13685), .B2(
        P2_LWORD_REG_0__SCAN_IN), .ZN(n13669) );
  NAND2_X1 U17192 ( .A1(n13669), .A2(n13668), .ZN(P2_U2967) );
  AOI22_X1 U17193 ( .A1(n9676), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n13685), .B2(
        P2_UWORD_REG_11__SCAN_IN), .ZN(n13671) );
  NAND2_X1 U17194 ( .A1(n13671), .A2(n13670), .ZN(P2_U2963) );
  AOI22_X1 U17195 ( .A1(n9676), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n13685), .B2(
        P2_LWORD_REG_6__SCAN_IN), .ZN(n13673) );
  NAND2_X1 U17196 ( .A1(n13673), .A2(n13672), .ZN(P2_U2973) );
  AOI22_X1 U17197 ( .A1(n9676), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n13685), .B2(
        P2_LWORD_REG_13__SCAN_IN), .ZN(n13678) );
  INV_X1 U17198 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n13675) );
  NAND2_X1 U17199 ( .A1(n13676), .A2(BUF1_REG_13__SCAN_IN), .ZN(n13674) );
  OAI21_X1 U17200 ( .B1(n13676), .B2(n13675), .A(n13674), .ZN(n16757) );
  NAND2_X1 U17201 ( .A1(n13677), .A2(n16757), .ZN(n13679) );
  NAND2_X1 U17202 ( .A1(n13678), .A2(n13679), .ZN(P2_U2980) );
  AOI22_X1 U17203 ( .A1(n9676), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n13685), .B2(
        P2_UWORD_REG_13__SCAN_IN), .ZN(n13680) );
  NAND2_X1 U17204 ( .A1(n13680), .A2(n13679), .ZN(P2_U2965) );
  AOI22_X1 U17205 ( .A1(n9676), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n13685), .B2(
        P2_UWORD_REG_7__SCAN_IN), .ZN(n13682) );
  NAND2_X1 U17206 ( .A1(n13682), .A2(n13681), .ZN(P2_U2959) );
  AOI22_X1 U17207 ( .A1(n9676), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n13685), .B2(
        P2_UWORD_REG_4__SCAN_IN), .ZN(n13684) );
  NAND2_X1 U17208 ( .A1(n13684), .A2(n13683), .ZN(P2_U2956) );
  AOI22_X1 U17209 ( .A1(n9676), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n13685), .B2(
        P2_UWORD_REG_3__SCAN_IN), .ZN(n13688) );
  NAND2_X1 U17210 ( .A1(n13688), .A2(n13687), .ZN(P2_U2955) );
  INV_X1 U17211 ( .A(P3_EBX_REG_4__SCAN_IN), .ZN(n18764) );
  NAND3_X1 U17212 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n18763) );
  NOR3_X1 U17213 ( .A1(n18764), .A2(n18544), .A3(n18763), .ZN(n18762) );
  INV_X1 U17214 ( .A(P3_EBX_REG_8__SCAN_IN), .ZN(n18465) );
  NAND2_X1 U17215 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(P3_EBX_REG_6__SCAN_IN), 
        .ZN(n13750) );
  NOR4_X1 U17216 ( .A1(n18459), .A2(n18465), .A3(n18510), .A4(n13750), .ZN(
        n13725) );
  INV_X1 U17217 ( .A(P3_EBX_REG_10__SCAN_IN), .ZN(n18752) );
  NOR2_X1 U17218 ( .A1(n18717), .A2(n18752), .ZN(n13726) );
  NAND4_X1 U17219 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n18762), .A3(n13725), 
        .A4(n13726), .ZN(n13806) );
  NOR2_X1 U17220 ( .A1(n18410), .A2(n13806), .ZN(n18693) );
  NAND2_X1 U17221 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n18693), .ZN(n13771) );
  NOR2_X1 U17222 ( .A1(n18384), .A2(n13771), .ZN(n13774) );
  NAND2_X1 U17223 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n13774), .ZN(n13831) );
  NAND2_X1 U17224 ( .A1(n19577), .A2(n19588), .ZN(n13689) );
  NOR2_X1 U17225 ( .A1(n13691), .A2(n20047), .ZN(n13692) );
  AOI211_X1 U17226 ( .C1(n19588), .C2(n13831), .A(n18364), .B(n13832), .ZN(
        n13710) );
  AND2_X1 U17227 ( .A1(n18785), .A2(n19588), .ZN(n18782) );
  NOR2_X1 U17228 ( .A1(n18780), .A2(n13831), .ZN(n13834) );
  NOR2_X1 U17229 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n13834), .ZN(n13709) );
  INV_X1 U17230 ( .A(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13695) );
  NAND2_X1 U17231 ( .A1(n13185), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n13694) );
  NAND2_X1 U17232 ( .A1(n18699), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n13693) );
  OAI211_X1 U17233 ( .C1(n18735), .C2(n13695), .A(n13694), .B(n13693), .ZN(
        n13696) );
  INV_X1 U17234 ( .A(n13696), .ZN(n13700) );
  AOI22_X1 U17235 ( .A1(n18704), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n9683), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13699) );
  AOI22_X1 U17236 ( .A1(n18706), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n18705), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13698) );
  NAND2_X1 U17237 ( .A1(n18731), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n13697) );
  NAND4_X1 U17238 ( .A1(n13700), .A2(n13699), .A3(n13698), .A4(n13697), .ZN(
        n13707) );
  AOI22_X1 U17239 ( .A1(n18736), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n13878), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13705) );
  AOI22_X1 U17240 ( .A1(n13279), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n18596), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n13704) );
  AOI22_X1 U17241 ( .A1(n18740), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n18739), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13703) );
  AOI22_X1 U17242 ( .A1(n18738), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n18737), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13702) );
  NAND4_X1 U17243 ( .A1(n13705), .A2(n13704), .A3(n13703), .A4(n13702), .ZN(
        n13706) );
  OR2_X1 U17244 ( .A1(n13707), .A2(n13706), .ZN(n18851) );
  INV_X1 U17245 ( .A(n18851), .ZN(n13708) );
  OAI22_X1 U17246 ( .A1(n13710), .A2(n13709), .B1(n13708), .B2(n18770), .ZN(
        P3_U2686) );
  INV_X1 U17247 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n18768) );
  NAND2_X1 U17248 ( .A1(n9703), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n13712) );
  NAND2_X1 U17249 ( .A1(n18699), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n13711) );
  OAI211_X1 U17250 ( .C1(n18735), .C2(n18768), .A(n13712), .B(n13711), .ZN(
        n13713) );
  INV_X1 U17251 ( .A(n13713), .ZN(n13717) );
  AOI22_X1 U17252 ( .A1(n18704), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n18703), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13716) );
  AOI22_X1 U17253 ( .A1(n18706), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n18705), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13715) );
  NAND2_X1 U17254 ( .A1(n13795), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n13714) );
  NAND4_X1 U17255 ( .A1(n13717), .A2(n13716), .A3(n13715), .A4(n13714), .ZN(
        n13724) );
  AOI22_X1 U17256 ( .A1(n18736), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n13878), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n13722) );
  AOI22_X1 U17257 ( .A1(n13279), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n18596), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n13721) );
  AOI22_X1 U17258 ( .A1(n18740), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n18739), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n13720) );
  AOI22_X1 U17259 ( .A1(n13718), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n18737), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13719) );
  NAND4_X1 U17260 ( .A1(n13722), .A2(n13721), .A3(n13720), .A4(n13719), .ZN(
        n13723) );
  NOR2_X1 U17261 ( .A1(n13724), .A2(n13723), .ZN(n17738) );
  NAND3_X1 U17262 ( .A1(n18785), .A2(n18762), .A3(n13725), .ZN(n18747) );
  INV_X1 U17263 ( .A(n18747), .ZN(n13727) );
  NAND3_X1 U17264 ( .A1(n13727), .A2(n19588), .A3(n13726), .ZN(n18718) );
  INV_X1 U17265 ( .A(n18718), .ZN(n13729) );
  INV_X1 U17266 ( .A(P3_EBX_REG_12__SCAN_IN), .ZN(n13728) );
  NAND2_X1 U17267 ( .A1(n13729), .A2(n13728), .ZN(n13731) );
  NAND3_X1 U17268 ( .A1(n18718), .A2(P3_EBX_REG_12__SCAN_IN), .A3(n18770), 
        .ZN(n13730) );
  OAI211_X1 U17269 ( .C1(n17738), .C2(n18770), .A(n13731), .B(n13730), .ZN(
        P3_U2691) );
  INV_X1 U17270 ( .A(n13732), .ZN(n13733) );
  INV_X1 U17271 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .ZN(n21624) );
  NAND2_X1 U17272 ( .A1(n18052), .A2(n21376), .ZN(n20940) );
  OAI211_X1 U17273 ( .C1(n13733), .C2(n21624), .A(n14044), .B(n20940), .ZN(
        P1_U2801) );
  INV_X1 U17274 ( .A(n18706), .ZN(n18724) );
  INV_X1 U17275 ( .A(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n13762) );
  INV_X1 U17276 ( .A(n18705), .ZN(n18722) );
  INV_X1 U17277 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13759) );
  OAI22_X1 U17278 ( .A1(n18724), .A2(n13762), .B1(n18722), .B2(n13759), .ZN(
        n13737) );
  INV_X1 U17279 ( .A(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13735) );
  INV_X1 U17280 ( .A(n13734), .ZN(n18726) );
  INV_X1 U17281 ( .A(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13753) );
  OAI22_X1 U17282 ( .A1(n18728), .A2(n13735), .B1(n18726), .B2(n13753), .ZN(
        n13736) );
  AOI211_X1 U17283 ( .C1(n18731), .C2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A(
        n13737), .B(n13736), .ZN(n13739) );
  AOI22_X1 U17284 ( .A1(n9704), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n18732), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13738) );
  OAI211_X1 U17285 ( .C1(n9681), .C2(n21742), .A(n13739), .B(n13738), .ZN(
        n13745) );
  AOI22_X1 U17286 ( .A1(n18736), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n13878), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n13743) );
  AOI22_X1 U17287 ( .A1(n13279), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n18596), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13742) );
  AOI22_X1 U17288 ( .A1(n18738), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n18737), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13741) );
  AOI22_X1 U17289 ( .A1(n18740), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n18739), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n13740) );
  NAND4_X1 U17290 ( .A1(n13743), .A2(n13742), .A3(n13741), .A4(n13740), .ZN(
        n13744) );
  OR2_X1 U17291 ( .A1(n13745), .A2(n13744), .ZN(n18857) );
  INV_X1 U17292 ( .A(n18857), .ZN(n13749) );
  INV_X1 U17293 ( .A(n13834), .ZN(n13746) );
  NAND3_X1 U17294 ( .A1(n13746), .A2(P3_EBX_REG_16__SCAN_IN), .A3(n18770), 
        .ZN(n13748) );
  NAND3_X1 U17295 ( .A1(n18782), .A2(n13831), .A3(n13774), .ZN(n13747) );
  OAI211_X1 U17296 ( .C1(n13749), .C2(n18770), .A(n13748), .B(n13747), .ZN(
        P3_U2687) );
  NAND3_X1 U17297 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n18785), .A3(n18762), .ZN(
        n18756) );
  NOR3_X1 U17298 ( .A1(n18465), .A2(n13750), .A3(n18756), .ZN(n13829) );
  NOR2_X1 U17299 ( .A1(n13750), .A2(n18756), .ZN(n13751) );
  AOI22_X1 U17300 ( .A1(n13751), .A2(n19588), .B1(P3_EBX_REG_8__SCAN_IN), .B2(
        n18770), .ZN(n13770) );
  OAI22_X1 U17301 ( .A1(n18724), .A2(n13753), .B1(n18722), .B2(n13752), .ZN(
        n13756) );
  INV_X1 U17302 ( .A(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13754) );
  OAI22_X1 U17303 ( .A1(n18728), .A2(n21699), .B1(n18726), .B2(n13754), .ZN(
        n13755) );
  AOI211_X1 U17304 ( .C1(n18731), .C2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A(
        n13756), .B(n13755), .ZN(n13758) );
  AOI22_X1 U17305 ( .A1(n9703), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n18732), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13757) );
  OAI211_X1 U17306 ( .C1(n18735), .C2(n13759), .A(n13758), .B(n13757), .ZN(
        n13768) );
  INV_X1 U17307 ( .A(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n19647) );
  INV_X1 U17308 ( .A(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n13760) );
  OAI22_X1 U17309 ( .A1(n19647), .A2(n13761), .B1(n13819), .B2(n13760), .ZN(
        n13767) );
  INV_X1 U17310 ( .A(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n19621) );
  OAI22_X1 U17311 ( .A1(n11593), .A2(n19621), .B1(n14603), .B2(n13762), .ZN(
        n13766) );
  AOI22_X1 U17312 ( .A1(n18736), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n13878), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n13764) );
  AOI22_X1 U17313 ( .A1(n18738), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n18737), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13763) );
  NAND2_X1 U17314 ( .A1(n13764), .A2(n13763), .ZN(n13765) );
  OR4_X1 U17315 ( .A1(n13768), .A2(n13767), .A3(n13766), .A4(n13765), .ZN(
        n18881) );
  INV_X1 U17316 ( .A(n18881), .ZN(n13769) );
  OAI22_X1 U17317 ( .A1(n13829), .A2(n13770), .B1(n13769), .B2(n18770), .ZN(
        P3_U2695) );
  INV_X1 U17318 ( .A(n13771), .ZN(n13772) );
  NAND2_X1 U17319 ( .A1(n18785), .A2(n13772), .ZN(n13773) );
  NAND2_X1 U17320 ( .A1(n18770), .A2(n13773), .ZN(n18697) );
  NAND2_X1 U17321 ( .A1(n13774), .A2(n18782), .ZN(n13790) );
  INV_X1 U17322 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n18754) );
  NAND2_X1 U17323 ( .A1(n9704), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n13776) );
  NAND2_X1 U17324 ( .A1(n18699), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n13775) );
  OAI211_X1 U17325 ( .C1(n18735), .C2(n18754), .A(n13776), .B(n13775), .ZN(
        n13777) );
  INV_X1 U17326 ( .A(n13777), .ZN(n13781) );
  AOI22_X1 U17327 ( .A1(n18704), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n18703), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13780) );
  AOI22_X1 U17328 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n18706), .B1(
        n18705), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13779) );
  NAND2_X1 U17329 ( .A1(n18731), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n13778) );
  NAND4_X1 U17330 ( .A1(n13781), .A2(n13780), .A3(n13779), .A4(n13778), .ZN(
        n13787) );
  AOI22_X1 U17331 ( .A1(n18736), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13878), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n13785) );
  INV_X1 U17332 ( .A(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n19669) );
  AOI22_X1 U17333 ( .A1(n13279), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n18596), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n13784) );
  AOI22_X1 U17334 ( .A1(n18738), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n18737), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13783) );
  AOI22_X1 U17335 ( .A1(n18740), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n18739), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n13782) );
  NAND4_X1 U17336 ( .A1(n13785), .A2(n13784), .A3(n13783), .A4(n13782), .ZN(
        n13786) );
  NOR2_X1 U17337 ( .A1(n13787), .A2(n13786), .ZN(n14302) );
  INV_X1 U17338 ( .A(n14302), .ZN(n13788) );
  OR2_X1 U17339 ( .A1(n18770), .A2(n13788), .ZN(n13789) );
  OAI211_X1 U17340 ( .C1(n18697), .C2(P3_EBX_REG_15__SCAN_IN), .A(n13790), .B(
        n13789), .ZN(n13791) );
  INV_X1 U17341 ( .A(n13791), .ZN(P3_U2688) );
  INV_X1 U17342 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17707) );
  NAND2_X1 U17343 ( .A1(n9703), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n13793) );
  NAND2_X1 U17344 ( .A1(n18699), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n13792) );
  OAI211_X1 U17345 ( .C1(n9681), .C2(n17707), .A(n13793), .B(n13792), .ZN(
        n13794) );
  INV_X1 U17346 ( .A(n13794), .ZN(n13799) );
  AOI22_X1 U17347 ( .A1(n18704), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n9683), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13798) );
  AOI22_X1 U17348 ( .A1(n18706), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n18705), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13797) );
  NAND2_X1 U17349 ( .A1(n13795), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n13796) );
  NAND4_X1 U17350 ( .A1(n13799), .A2(n13798), .A3(n13797), .A4(n13796), .ZN(
        n13805) );
  AOI22_X1 U17351 ( .A1(n18736), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13878), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13803) );
  AOI22_X1 U17352 ( .A1(n13279), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n18596), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13802) );
  AOI22_X1 U17353 ( .A1(n18740), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n18739), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13801) );
  AOI22_X1 U17354 ( .A1(n18738), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n18737), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13800) );
  NAND4_X1 U17355 ( .A1(n13803), .A2(n13802), .A3(n13801), .A4(n13800), .ZN(
        n13804) );
  NOR2_X1 U17356 ( .A1(n13805), .A2(n13804), .ZN(n17736) );
  AOI211_X1 U17357 ( .C1(n18410), .C2(n13806), .A(n18693), .B(n18780), .ZN(
        n13807) );
  AOI21_X1 U17358 ( .B1(P3_EBX_REG_13__SCAN_IN), .B2(n13832), .A(n13807), .ZN(
        n13808) );
  OAI21_X1 U17359 ( .B1(n17736), .B2(n18770), .A(n13808), .ZN(P3_U2690) );
  INV_X1 U17360 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n18778) );
  INV_X1 U17361 ( .A(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13810) );
  OAI22_X1 U17362 ( .A1(n18724), .A2(n13810), .B1(n18722), .B2(n13809), .ZN(
        n13814) );
  INV_X1 U17363 ( .A(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13812) );
  INV_X1 U17364 ( .A(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13811) );
  OAI22_X1 U17365 ( .A1(n18728), .A2(n13812), .B1(n18726), .B2(n13811), .ZN(
        n13813) );
  AOI211_X1 U17366 ( .C1(n18731), .C2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A(
        n13814), .B(n13813), .ZN(n13816) );
  AOI22_X1 U17367 ( .A1(n13185), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n18732), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13815) );
  OAI211_X1 U17368 ( .C1(n18778), .C2(n18735), .A(n13816), .B(n13815), .ZN(
        n13828) );
  INV_X1 U17369 ( .A(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n13820) );
  AOI22_X1 U17370 ( .A1(n18740), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n18739), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13818) );
  NAND2_X1 U17371 ( .A1(n13279), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n13817) );
  OAI211_X1 U17372 ( .C1(n13820), .C2(n13819), .A(n13818), .B(n13817), .ZN(
        n13827) );
  INV_X1 U17373 ( .A(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13822) );
  INV_X1 U17374 ( .A(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13821) );
  OAI22_X1 U17375 ( .A1(n14593), .A2(n13822), .B1(n14591), .B2(n13821), .ZN(
        n13826) );
  INV_X1 U17376 ( .A(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13824) );
  OAI22_X1 U17377 ( .A1(n14596), .A2(n13824), .B1(n14594), .B2(n13823), .ZN(
        n13825) );
  NOR4_X1 U17378 ( .A1(n13828), .A2(n13827), .A3(n13826), .A4(n13825), .ZN(
        n14159) );
  OAI211_X1 U17379 ( .C1(n13829), .C2(P3_EBX_REG_9__SCAN_IN), .A(n18747), .B(
        n18770), .ZN(n13830) );
  OAI21_X1 U17380 ( .B1(n14159), .B2(n18770), .A(n13830), .ZN(P3_U2694) );
  INV_X1 U17381 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n13833) );
  OR2_X1 U17382 ( .A1(n13833), .A2(n13885), .ZN(n13850) );
  NAND3_X1 U17383 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n13834), .A3(n13833), 
        .ZN(n13849) );
  INV_X1 U17384 ( .A(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n19601) );
  INV_X1 U17385 ( .A(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n13836) );
  INV_X1 U17386 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13835) );
  OAI22_X1 U17387 ( .A1(n18724), .A2(n13836), .B1(n18722), .B2(n13835), .ZN(
        n13839) );
  INV_X1 U17388 ( .A(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13837) );
  INV_X1 U17389 ( .A(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n18723) );
  OAI22_X1 U17390 ( .A1(n18728), .A2(n13837), .B1(n18726), .B2(n18723), .ZN(
        n13838) );
  AOI211_X1 U17391 ( .C1(n18731), .C2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A(
        n13839), .B(n13838), .ZN(n13841) );
  AOI22_X1 U17392 ( .A1(n13185), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n18732), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13840) );
  OAI211_X1 U17393 ( .C1(n19601), .C2(n18735), .A(n13841), .B(n13840), .ZN(
        n13847) );
  AOI22_X1 U17394 ( .A1(n18736), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n13878), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13845) );
  AOI22_X1 U17395 ( .A1(n13279), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n18596), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n13844) );
  AOI22_X1 U17396 ( .A1(n18738), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n18737), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13843) );
  AOI22_X1 U17397 ( .A1(n18740), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n18739), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n13842) );
  NAND4_X1 U17398 ( .A1(n13845), .A2(n13844), .A3(n13843), .A4(n13842), .ZN(
        n13846) );
  OR2_X1 U17399 ( .A1(n13847), .A2(n13846), .ZN(n18846) );
  NAND2_X1 U17400 ( .A1(n18749), .A2(n18846), .ZN(n13848) );
  OAI211_X1 U17401 ( .C1(n13850), .C2(n18749), .A(n13849), .B(n13848), .ZN(
        P3_U2685) );
  INV_X1 U17402 ( .A(n13851), .ZN(n13853) );
  OAI21_X1 U17403 ( .B1(n17453), .B2(n13853), .A(n13852), .ZN(n13854) );
  INV_X1 U17404 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n13856) );
  INV_X1 U17405 ( .A(P2_UWORD_REG_3__SCAN_IN), .ZN(n21773) );
  INV_X2 U17406 ( .A(n20240), .ZN(n20243) );
  INV_X1 U17407 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n18164) );
  OAI222_X1 U17408 ( .A1(n20211), .A2(n13856), .B1(n20240), .B2(n21773), .C1(
        n20241), .C2(n18164), .ZN(P2_U2932) );
  INV_X1 U17409 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n13857) );
  INV_X1 U17410 ( .A(P2_UWORD_REG_11__SCAN_IN), .ZN(n21757) );
  INV_X1 U17411 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n18173) );
  OAI222_X1 U17412 ( .A1(n20211), .A2(n13857), .B1(n20240), .B2(n21757), .C1(
        n20241), .C2(n18173), .ZN(P2_U2924) );
  INV_X1 U17413 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n21882) );
  OR2_X1 U17414 ( .A1(n15971), .A2(n15147), .ZN(n13861) );
  NAND2_X1 U17415 ( .A1(n13866), .A2(n13858), .ZN(n13859) );
  NAND2_X1 U17416 ( .A1(n13859), .A2(n12622), .ZN(n13860) );
  NAND2_X1 U17417 ( .A1(n13861), .A2(n13860), .ZN(n20937) );
  INV_X1 U17418 ( .A(n15147), .ZN(n14822) );
  NAND3_X1 U17419 ( .A1(n14822), .A2(n13990), .A3(n14098), .ZN(n13862) );
  AND2_X1 U17420 ( .A1(n13862), .A2(n21532), .ZN(n21616) );
  OR2_X1 U17421 ( .A1(n20937), .A2(n21616), .ZN(n15952) );
  AND2_X1 U17422 ( .A1(n15952), .A2(n20935), .ZN(n20945) );
  AND2_X1 U17423 ( .A1(n13863), .A2(n12622), .ZN(n13864) );
  MUX2_X1 U17424 ( .A(n13864), .B(n14434), .S(n15971), .Z(n13868) );
  NAND2_X1 U17425 ( .A1(n13866), .A2(n13865), .ZN(n13867) );
  AND2_X1 U17426 ( .A1(n13868), .A2(n13867), .ZN(n15951) );
  INV_X1 U17427 ( .A(n15951), .ZN(n13869) );
  NAND2_X1 U17428 ( .A1(n13869), .A2(n20945), .ZN(n13870) );
  OAI21_X1 U17429 ( .B1(n21882), .B2(n20945), .A(n13870), .ZN(P1_U3484) );
  INV_X1 U17430 ( .A(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n19604) );
  INV_X1 U17431 ( .A(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13871) );
  INV_X1 U17432 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n18772) );
  OAI22_X1 U17433 ( .A1(n18724), .A2(n13871), .B1(n18722), .B2(n18772), .ZN(
        n13875) );
  INV_X1 U17434 ( .A(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13873) );
  INV_X1 U17435 ( .A(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13872) );
  OAI22_X1 U17436 ( .A1(n18728), .A2(n13873), .B1(n18726), .B2(n13872), .ZN(
        n13874) );
  AOI211_X1 U17437 ( .C1(n18731), .C2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A(
        n13875), .B(n13874), .ZN(n13877) );
  AOI22_X1 U17438 ( .A1(n9704), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n18732), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13876) );
  OAI211_X1 U17439 ( .C1(n18735), .C2(n19604), .A(n13877), .B(n13876), .ZN(
        n13884) );
  AOI22_X1 U17440 ( .A1(n18736), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n13878), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13882) );
  AOI22_X1 U17441 ( .A1(n13279), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n18596), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n13881) );
  AOI22_X1 U17442 ( .A1(n18738), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n18737), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13880) );
  AOI22_X1 U17443 ( .A1(n18740), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n18739), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13879) );
  NAND4_X1 U17444 ( .A1(n13882), .A2(n13881), .A3(n13880), .A4(n13879), .ZN(
        n13883) );
  NOR2_X1 U17445 ( .A1(n13884), .A2(n13883), .ZN(n17728) );
  NAND2_X1 U17446 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n13885), .ZN(n18584) );
  OAI21_X1 U17447 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n13885), .A(n18584), .ZN(
        n13886) );
  OR2_X1 U17448 ( .A1(n13886), .A2(n18749), .ZN(n13887) );
  OAI21_X1 U17449 ( .B1(n17728), .B2(n18770), .A(n13887), .ZN(P3_U2684) );
  INV_X1 U17450 ( .A(P3_EBX_REG_20__SCAN_IN), .ZN(n18585) );
  OAI21_X1 U17451 ( .B1(n18584), .B2(n18585), .A(n18770), .ZN(n18675) );
  INV_X1 U17452 ( .A(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n14670) );
  INV_X1 U17453 ( .A(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n14672) );
  OAI22_X1 U17454 ( .A1(n18724), .A2(n14672), .B1(n18722), .B2(n18768), .ZN(
        n13891) );
  INV_X1 U17455 ( .A(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13889) );
  INV_X1 U17456 ( .A(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13888) );
  OAI22_X1 U17457 ( .A1(n18728), .A2(n13889), .B1(n18726), .B2(n13888), .ZN(
        n13890) );
  AOI211_X1 U17458 ( .C1(n18731), .C2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A(
        n13891), .B(n13890), .ZN(n13893) );
  AOI22_X1 U17459 ( .A1(n13185), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n18732), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13892) );
  OAI211_X1 U17460 ( .C1(n9681), .C2(n14670), .A(n13893), .B(n13892), .ZN(
        n13899) );
  AOI22_X1 U17461 ( .A1(n18736), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n13878), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n13897) );
  AOI22_X1 U17462 ( .A1(n13279), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n18596), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n13896) );
  AOI22_X1 U17463 ( .A1(n18738), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n18737), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13895) );
  AOI22_X1 U17464 ( .A1(n18740), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n18739), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n13894) );
  NAND4_X1 U17465 ( .A1(n13897), .A2(n13896), .A3(n13895), .A4(n13894), .ZN(
        n13898) );
  OR2_X1 U17466 ( .A1(n13899), .A2(n13898), .ZN(n18840) );
  NAND2_X1 U17467 ( .A1(n18749), .A2(n18840), .ZN(n13901) );
  NOR2_X1 U17468 ( .A1(n18584), .A2(n18787), .ZN(n14579) );
  NAND2_X1 U17469 ( .A1(n18585), .A2(n14579), .ZN(n13900) );
  OAI211_X1 U17470 ( .C1(n18675), .C2(n18585), .A(n13901), .B(n13900), .ZN(
        P3_U2683) );
  INV_X1 U17471 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n13903) );
  AOI22_X1 U17472 ( .A1(n20243), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n20242), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n13902) );
  OAI21_X1 U17473 ( .B1(n13903), .B2(n20211), .A(n13902), .ZN(P2_U2928) );
  INV_X1 U17474 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n13905) );
  AOI22_X1 U17475 ( .A1(n20243), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n20242), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n13904) );
  OAI21_X1 U17476 ( .B1(n13905), .B2(n20211), .A(n13904), .ZN(P2_U2929) );
  INV_X1 U17477 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n13907) );
  AOI22_X1 U17478 ( .A1(n20243), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n20242), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n13906) );
  OAI21_X1 U17479 ( .B1(n13907), .B2(n20211), .A(n13906), .ZN(P2_U2934) );
  INV_X1 U17480 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n13909) );
  AOI22_X1 U17481 ( .A1(n20243), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n20242), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n13908) );
  OAI21_X1 U17482 ( .B1(n13909), .B2(n20211), .A(n13908), .ZN(P2_U2931) );
  INV_X1 U17483 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n13911) );
  AOI22_X1 U17484 ( .A1(n20243), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n20242), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n13910) );
  OAI21_X1 U17485 ( .B1(n13911), .B2(n20211), .A(n13910), .ZN(P2_U2930) );
  INV_X1 U17486 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n13913) );
  AOI22_X1 U17487 ( .A1(n20243), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n20242), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n13912) );
  OAI21_X1 U17488 ( .B1(n13913), .B2(n20211), .A(n13912), .ZN(P2_U2926) );
  AOI22_X1 U17489 ( .A1(n20243), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n20242), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n13914) );
  OAI21_X1 U17490 ( .B1(n13915), .B2(n20211), .A(n13914), .ZN(P2_U2925) );
  AOI22_X1 U17491 ( .A1(n20243), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(n20242), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .ZN(n13916) );
  OAI21_X1 U17492 ( .B1(n13917), .B2(n20211), .A(n13916), .ZN(P2_U2921) );
  AOI22_X1 U17493 ( .A1(n20243), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n20242), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n13918) );
  OAI21_X1 U17494 ( .B1(n13919), .B2(n20211), .A(n13918), .ZN(P2_U2923) );
  AOI22_X1 U17495 ( .A1(n20243), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n20242), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n13920) );
  OAI21_X1 U17496 ( .B1(n21700), .B2(n20211), .A(n13920), .ZN(P2_U2922) );
  AOI22_X1 U17497 ( .A1(n20243), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n20242), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n13921) );
  OAI21_X1 U17498 ( .B1(n13922), .B2(n20211), .A(n13921), .ZN(P2_U2927) );
  INV_X1 U17499 ( .A(n20249), .ZN(n18070) );
  XNOR2_X1 U17500 ( .A(n13924), .B(n13923), .ZN(n13925) );
  XOR2_X1 U17501 ( .A(n13925), .B(n14054), .Z(n14065) );
  NOR2_X1 U17502 ( .A1(n17136), .A2(n20829), .ZN(n14064) );
  AOI21_X1 U17503 ( .B1(n18070), .B2(n14065), .A(n14064), .ZN(n13929) );
  AOI21_X1 U17504 ( .B1(n14054), .B2(n13927), .A(n13926), .ZN(n14057) );
  NAND2_X1 U17505 ( .A1(n14057), .A2(n17155), .ZN(n13928) );
  OAI211_X1 U17506 ( .C1(n18060), .C2(n21776), .A(n13929), .B(n13928), .ZN(
        n13930) );
  AOI21_X1 U17507 ( .B1(n18063), .B2(n21776), .A(n13930), .ZN(n13931) );
  OAI21_X1 U17508 ( .B1(n14040), .B2(n17126), .A(n13931), .ZN(P2_U3013) );
  OAI21_X1 U17509 ( .B1(n15937), .B2(n15960), .A(n18008), .ZN(n13932) );
  OAI21_X1 U17510 ( .B1(n14098), .B2(n13424), .A(n13932), .ZN(n13934) );
  INV_X1 U17511 ( .A(n14433), .ZN(n13933) );
  AOI21_X1 U17512 ( .B1(n13934), .B2(n21532), .A(n13933), .ZN(n13935) );
  MUX2_X1 U17513 ( .A(n14434), .B(n13935), .S(n15971), .Z(n13941) );
  INV_X1 U17514 ( .A(n13936), .ZN(n13937) );
  OR2_X1 U17515 ( .A1(n14459), .A2(n13937), .ZN(n14130) );
  OAI211_X1 U17516 ( .C1(n13439), .C2(n14381), .A(n13938), .B(n14130), .ZN(
        n13939) );
  INV_X1 U17517 ( .A(n13939), .ZN(n13940) );
  NAND2_X1 U17518 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n18047) );
  NAND2_X1 U17519 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n15763), .ZN(n18053) );
  INV_X1 U17520 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n20944) );
  NOR2_X1 U17521 ( .A1(n18053), .A2(n20944), .ZN(n13942) );
  AOI21_X1 U17522 ( .B1(n15939), .B2(n20935), .A(n13942), .ZN(n18043) );
  NAND2_X1 U17523 ( .A1(n20939), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n13943) );
  INV_X1 U17524 ( .A(n13944), .ZN(n21471) );
  INV_X1 U17525 ( .A(n13945), .ZN(n13946) );
  AND4_X1 U17526 ( .A1(n13946), .A2(n14459), .A3(n13424), .A4(n13448), .ZN(
        n13947) );
  NAND2_X1 U17527 ( .A1(n13948), .A2(n13947), .ZN(n15935) );
  INV_X1 U17528 ( .A(n15937), .ZN(n14432) );
  INV_X1 U17529 ( .A(n13949), .ZN(n14456) );
  INV_X1 U17530 ( .A(n13950), .ZN(n13951) );
  NAND2_X1 U17531 ( .A1(n14456), .A2(n13951), .ZN(n13954) );
  OAI22_X1 U17532 ( .A1(n14432), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B1(
        n13954), .B2(n11896), .ZN(n13952) );
  AOI21_X1 U17533 ( .B1(n21471), .B2(n15935), .A(n13952), .ZN(n15938) );
  INV_X1 U17534 ( .A(n13953), .ZN(n21602) );
  NOR2_X1 U17535 ( .A1(n15938), .A2(n21602), .ZN(n13956) );
  INV_X1 U17536 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n15514) );
  AOI22_X1 U17537 ( .A1(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n21144), .B2(n15514), .ZN(
        n15777) );
  NAND2_X1 U17538 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n15776) );
  OAI22_X1 U17539 ( .A1(n21594), .A2(n13954), .B1(n15777), .B2(n15776), .ZN(
        n13955) );
  OAI21_X1 U17540 ( .B1(n13956), .B2(n13955), .A(n21597), .ZN(n13957) );
  OAI21_X1 U17541 ( .B1(n21597), .B2(n13958), .A(n13957), .ZN(P1_U3473) );
  INV_X1 U17542 ( .A(n14014), .ZN(n13960) );
  INV_X1 U17543 ( .A(n14161), .ZN(n13959) );
  NAND2_X1 U17544 ( .A1(n13959), .A2(n17962), .ZN(n14009) );
  NAND2_X1 U17545 ( .A1(n13960), .A2(n14009), .ZN(n14425) );
  INV_X1 U17546 ( .A(n14425), .ZN(n13987) );
  AND2_X1 U17547 ( .A1(n19571), .A2(n20150), .ZN(n13962) );
  INV_X1 U17548 ( .A(n20022), .ZN(n13961) );
  AOI22_X1 U17549 ( .A1(n20017), .A2(n13962), .B1(n13966), .B2(n13961), .ZN(
        n13974) );
  XNOR2_X1 U17550 ( .A(n19568), .B(n13963), .ZN(n13964) );
  OAI21_X1 U17551 ( .B1(n20149), .B2(n13964), .A(n20161), .ZN(n18190) );
  OR3_X1 U17552 ( .A1(n13966), .A2(n13965), .A3(n18190), .ZN(n13973) );
  OAI21_X1 U17553 ( .B1(n13968), .B2(n13967), .A(n18185), .ZN(n13970) );
  AND2_X1 U17554 ( .A1(n13970), .A2(n13969), .ZN(n14323) );
  OAI21_X1 U17555 ( .B1(n19577), .B2(n20022), .A(n14323), .ZN(n13971) );
  INV_X1 U17556 ( .A(n13971), .ZN(n13972) );
  OAI211_X1 U17557 ( .C1(n13974), .C2(n19583), .A(n13973), .B(n13972), .ZN(
        n13975) );
  NAND2_X1 U17558 ( .A1(n19546), .A2(n20021), .ZN(n19530) );
  INV_X1 U17559 ( .A(n13976), .ZN(n13977) );
  NAND2_X1 U17560 ( .A1(n13981), .A2(n13977), .ZN(n13978) );
  NAND2_X1 U17561 ( .A1(n13978), .A2(n14312), .ZN(n19428) );
  NOR2_X1 U17562 ( .A1(n19428), .A2(n20023), .ZN(n19355) );
  NOR3_X1 U17563 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n19355), .A3(
        n19522), .ZN(n14010) );
  NAND2_X1 U17564 ( .A1(n14312), .A2(n13979), .ZN(n13980) );
  NAND2_X1 U17565 ( .A1(n13981), .A2(n13980), .ZN(n19454) );
  AOI21_X1 U17566 ( .B1(n19546), .B2(n19314), .A(n17962), .ZN(n13982) );
  OAI21_X1 U17567 ( .B1(n14010), .B2(n13982), .A(n19442), .ZN(n13986) );
  INV_X1 U17568 ( .A(n20016), .ZN(n13983) );
  INV_X1 U17569 ( .A(P3_REIP_REG_0__SCAN_IN), .ZN(n13984) );
  NOR2_X1 U17570 ( .A1(n19442), .A2(n13984), .ZN(n14421) );
  AOI21_X1 U17571 ( .B1(n19545), .B2(n13987), .A(n14421), .ZN(n13985) );
  OAI211_X1 U17572 ( .C1(n13987), .C2(n19530), .A(n13986), .B(n13985), .ZN(
        P3_U2862) );
  INV_X1 U17573 ( .A(n13988), .ZN(n13989) );
  INV_X1 U17574 ( .A(n21060), .ZN(n21035) );
  NAND2_X1 U17575 ( .A1(n21035), .A2(n12634), .ZN(n14124) );
  NAND2_X1 U17576 ( .A1(n20939), .A2(n15763), .ZN(n21615) );
  INV_X2 U17577 ( .A(n21615), .ZN(n21054) );
  AOI22_X1 U17578 ( .A1(P1_UWORD_REG_14__SCAN_IN), .A2(n21054), .B1(n21053), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n13992) );
  OAI21_X1 U17579 ( .B1(n14799), .B2(n14124), .A(n13992), .ZN(P1_U2906) );
  AOI22_X1 U17580 ( .A1(P1_UWORD_REG_10__SCAN_IN), .A2(n21054), .B1(n21053), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n13993) );
  OAI21_X1 U17581 ( .B1(n15225), .B2(n14124), .A(n13993), .ZN(P1_U2910) );
  INV_X1 U17582 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n15229) );
  AOI22_X1 U17583 ( .A1(P1_UWORD_REG_9__SCAN_IN), .A2(n21054), .B1(n21053), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n13994) );
  OAI21_X1 U17584 ( .B1(n15229), .B2(n14124), .A(n13994), .ZN(P1_U2911) );
  INV_X1 U17585 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n21811) );
  AOI22_X1 U17586 ( .A1(P1_UWORD_REG_5__SCAN_IN), .A2(n21054), .B1(n21053), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n13995) );
  OAI21_X1 U17587 ( .B1(n21811), .B2(n14124), .A(n13995), .ZN(P1_U2915) );
  INV_X1 U17588 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n13997) );
  AOI22_X1 U17589 ( .A1(P1_UWORD_REG_4__SCAN_IN), .A2(n21054), .B1(n21053), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n13996) );
  OAI21_X1 U17590 ( .B1(n13997), .B2(n14124), .A(n13996), .ZN(P1_U2916) );
  AOI22_X1 U17591 ( .A1(P1_UWORD_REG_3__SCAN_IN), .A2(n21054), .B1(n21053), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n13998) );
  OAI21_X1 U17592 ( .B1(n12329), .B2(n14124), .A(n13998), .ZN(P1_U2917) );
  INV_X1 U17593 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n14000) );
  AOI22_X1 U17594 ( .A1(P1_UWORD_REG_7__SCAN_IN), .A2(n21054), .B1(n21053), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n13999) );
  OAI21_X1 U17595 ( .B1(n14000), .B2(n14124), .A(n13999), .ZN(P1_U2913) );
  INV_X1 U17596 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n14002) );
  AOI22_X1 U17597 ( .A1(P1_UWORD_REG_13__SCAN_IN), .A2(n21054), .B1(n21053), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n14001) );
  OAI21_X1 U17598 ( .B1(n14002), .B2(n14124), .A(n14001), .ZN(P1_U2907) );
  AOI22_X1 U17599 ( .A1(P1_UWORD_REG_12__SCAN_IN), .A2(n21054), .B1(n21053), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n14003) );
  OAI21_X1 U17600 ( .B1(n15212), .B2(n14124), .A(n14003), .ZN(P1_U2908) );
  INV_X1 U17601 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n14005) );
  AOI22_X1 U17602 ( .A1(P1_UWORD_REG_11__SCAN_IN), .A2(n21054), .B1(n21053), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n14004) );
  OAI21_X1 U17603 ( .B1(n14005), .B2(n14124), .A(n14004), .ZN(P1_U2909) );
  INV_X1 U17604 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n14007) );
  AOI22_X1 U17605 ( .A1(P1_UWORD_REG_6__SCAN_IN), .A2(n21054), .B1(n21053), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n14006) );
  OAI21_X1 U17606 ( .B1(n14007), .B2(n14124), .A(n14006), .ZN(P1_U2914) );
  AOI22_X1 U17607 ( .A1(P1_UWORD_REG_8__SCAN_IN), .A2(n21054), .B1(n21053), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n14008) );
  OAI21_X1 U17608 ( .B1(n15234), .B2(n14124), .A(n14008), .ZN(P1_U2912) );
  XNOR2_X1 U17609 ( .A(n14015), .B(n14009), .ZN(n19274) );
  INV_X1 U17610 ( .A(n19274), .ZN(n14019) );
  AND2_X1 U17611 ( .A1(n19546), .A2(n19467), .ZN(n19470) );
  OAI21_X1 U17612 ( .B1(n19454), .B2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n19470), .ZN(n14012) );
  NOR2_X1 U17613 ( .A1(n14010), .A2(n19527), .ZN(n14011) );
  MUX2_X1 U17614 ( .A(n14012), .B(n14011), .S(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .Z(n14018) );
  OAI21_X1 U17615 ( .B1(n14015), .B2(n14014), .A(n14013), .ZN(n14016) );
  INV_X1 U17616 ( .A(n14016), .ZN(n19276) );
  INV_X1 U17617 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n20136) );
  NOR2_X1 U17618 ( .A1(n19442), .A2(n20136), .ZN(n19273) );
  AOI21_X1 U17619 ( .B1(n19545), .B2(n19276), .A(n19273), .ZN(n14017) );
  OAI211_X1 U17620 ( .C1(n19530), .C2(n14019), .A(n14018), .B(n14017), .ZN(
        P3_U2861) );
  INV_X1 U17621 ( .A(n17524), .ZN(n14032) );
  INV_X1 U17622 ( .A(n14020), .ZN(n14021) );
  NAND2_X1 U17623 ( .A1(n14021), .A2(n11227), .ZN(n14763) );
  NAND2_X1 U17624 ( .A1(n17537), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n14022) );
  AOI22_X1 U17625 ( .A1(n14221), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n20888), .B2(n20919), .ZN(n14024) );
  NOR2_X1 U17626 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n14025) );
  NOR2_X1 U17627 ( .A1(n17537), .A2(n17703), .ZN(n14035) );
  OAI21_X1 U17628 ( .B1(n14026), .B2(n14025), .A(n14035), .ZN(n14027) );
  INV_X1 U17629 ( .A(n16344), .ZN(n14029) );
  NOR2_X1 U17630 ( .A1(n20914), .A2(n16344), .ZN(n14248) );
  INV_X1 U17631 ( .A(n14248), .ZN(n14028) );
  OAI211_X1 U17632 ( .C1(n17543), .C2(n14029), .A(n14028), .B(n16852), .ZN(
        n14031) );
  AOI22_X1 U17633 ( .A1(n16868), .A2(n14029), .B1(P2_EAX_REG_0__SCAN_IN), .B2(
        n16867), .ZN(n14030) );
  OAI211_X1 U17634 ( .C1(n14032), .C2(n14763), .A(n14031), .B(n14030), .ZN(
        P2_U2919) );
  INV_X1 U17635 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n16345) );
  MUX2_X1 U17636 ( .A(n14033), .B(n16345), .S(n16723), .Z(n14034) );
  OAI21_X1 U17637 ( .B1(n20914), .B2(n16733), .A(n14034), .ZN(P2_U2887) );
  INV_X1 U17638 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n20299) );
  NAND2_X1 U17639 ( .A1(n14221), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n14038) );
  NAND2_X1 U17640 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n17642) );
  NAND2_X1 U17641 ( .A1(n20909), .A2(n20919), .ZN(n20498) );
  AND2_X1 U17642 ( .A1(n17642), .A2(n20498), .ZN(n20695) );
  NAND2_X1 U17643 ( .A1(n20695), .A2(n20888), .ZN(n17618) );
  NAND2_X1 U17644 ( .A1(n14038), .A2(n17618), .ZN(n14039) );
  MUX2_X1 U17645 ( .A(n14041), .B(n14040), .S(n16728), .Z(n14042) );
  OAI21_X1 U17646 ( .B1(n17513), .B2(n16733), .A(n14042), .ZN(P2_U2886) );
  AND2_X1 U17647 ( .A1(n21617), .A2(n21533), .ZN(n14043) );
  OR2_X1 U17648 ( .A1(n14112), .A2(n10514), .ZN(n14169) );
  INV_X1 U17649 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n15279) );
  INV_X1 U17650 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n21032) );
  OR2_X1 U17651 ( .A1(n14112), .A2(n13450), .ZN(n14102) );
  NOR2_X1 U17652 ( .A1(n14801), .A2(n14046), .ZN(n14047) );
  AOI21_X1 U17653 ( .B1(DATAI_15_), .B2(n14801), .A(n14047), .ZN(n15280) );
  OAI222_X1 U17654 ( .A1(n14169), .A2(n15279), .B1(n14170), .B2(n21032), .C1(
        n14102), .C2(n15280), .ZN(P1_U2967) );
  INV_X1 U17655 ( .A(n17536), .ZN(n14050) );
  XNOR2_X1 U17656 ( .A(n14048), .B(n14049), .ZN(n17426) );
  INV_X1 U17657 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n20233) );
  OAI222_X1 U17658 ( .A1(n14763), .A2(n14050), .B1(n17426), .B2(n16864), .C1(
        n20233), .C2(n16744), .ZN(P2_U2913) );
  NOR2_X1 U17659 ( .A1(n14051), .A2(n14054), .ZN(n14056) );
  INV_X1 U17660 ( .A(n14052), .ZN(n20274) );
  AOI211_X1 U17661 ( .C1(n14054), .C2(n14053), .A(n20274), .B(n17419), .ZN(
        n14055) );
  AOI211_X1 U17662 ( .C1(n20267), .C2(n14057), .A(n14056), .B(n14055), .ZN(
        n14067) );
  OR2_X1 U17663 ( .A1(n14059), .A2(n14058), .ZN(n14060) );
  NAND2_X1 U17664 ( .A1(n14061), .A2(n14060), .ZN(n20907) );
  INV_X1 U17665 ( .A(n20907), .ZN(n14249) );
  OAI22_X1 U17666 ( .A1(n18091), .A2(n14249), .B1(n14062), .B2(n20259), .ZN(
        n14063) );
  AOI211_X1 U17667 ( .C1(n20279), .C2(n14065), .A(n14064), .B(n14063), .ZN(
        n14066) );
  NAND2_X1 U17668 ( .A1(n14067), .A2(n14066), .ZN(P2_U3045) );
  XNOR2_X1 U17669 ( .A(n17642), .B(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n20382) );
  AOI22_X1 U17670 ( .A1(n14221), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n20888), .B2(n20382), .ZN(n14069) );
  NAND2_X1 U17671 ( .A1(n14075), .A2(n14074), .ZN(n14078) );
  NAND2_X1 U17672 ( .A1(n17451), .A2(n14076), .ZN(n14077) );
  NAND2_X1 U17673 ( .A1(n14078), .A2(n14077), .ZN(n14216) );
  MUX2_X1 U17674 ( .A(n11013), .B(n14079), .S(n16728), .Z(n14080) );
  OAI21_X1 U17675 ( .B1(n20896), .B2(n16733), .A(n14080), .ZN(P2_U2885) );
  INV_X1 U17676 ( .A(n17587), .ZN(n14084) );
  OAI21_X1 U17677 ( .B1(n14081), .B2(n14083), .A(n14082), .ZN(n18073) );
  INV_X1 U17678 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n20231) );
  OAI222_X1 U17679 ( .A1(n14763), .A2(n14084), .B1(n18073), .B2(n16864), .C1(
        n20231), .C2(n16744), .ZN(P2_U2912) );
  INV_X1 U17680 ( .A(n14085), .ZN(n14088) );
  OAI21_X1 U17681 ( .B1(n14088), .B2(n14087), .A(n14086), .ZN(n15171) );
  OAI21_X1 U17682 ( .B1(n14089), .B2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13093), .ZN(n14152) );
  NAND2_X1 U17683 ( .A1(n15496), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n14146) );
  OAI21_X1 U17684 ( .B1(n21088), .B2(n14090), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n14091) );
  OAI211_X1 U17685 ( .C1(n14152), .C2(n20943), .A(n14146), .B(n14091), .ZN(
        n14092) );
  INV_X1 U17686 ( .A(n14092), .ZN(n14093) );
  OAI21_X1 U17687 ( .B1(n15511), .B2(n15171), .A(n14093), .ZN(P1_U2999) );
  OAI21_X1 U17688 ( .B1(n14095), .B2(n14094), .A(n14262), .ZN(n15164) );
  INV_X1 U17689 ( .A(n14385), .ZN(n14815) );
  NOR2_X1 U17690 ( .A1(n11872), .A2(n14381), .ZN(n14096) );
  NAND4_X1 U17691 ( .A1(n14097), .A2(n14815), .A3(n14096), .A4(n11861), .ZN(
        n14131) );
  INV_X1 U17692 ( .A(n15159), .ZN(n21134) );
  AOI22_X1 U17693 ( .A1(n15196), .A2(n21134), .B1(P1_EBX_REG_1__SCAN_IN), .B2(
        n15195), .ZN(n14101) );
  OAI21_X1 U17694 ( .B1(n15164), .B2(n15206), .A(n14101), .ZN(P1_U2871) );
  INV_X1 U17695 ( .A(DATAI_12_), .ZN(n14103) );
  INV_X1 U17696 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n18130) );
  MUX2_X1 U17697 ( .A(n14103), .B(n18130), .S(n15223), .Z(n15285) );
  INV_X1 U17698 ( .A(n15285), .ZN(n14104) );
  NAND2_X1 U17699 ( .A1(n21071), .A2(n14104), .ZN(n21080) );
  NAND2_X1 U17700 ( .A1(n14112), .A2(P1_UWORD_REG_12__SCAN_IN), .ZN(n14105) );
  OAI211_X1 U17701 ( .C1(n15212), .C2(n14169), .A(n21080), .B(n14105), .ZN(
        P1_U2949) );
  INV_X1 U17702 ( .A(DATAI_9_), .ZN(n14107) );
  INV_X1 U17703 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n14106) );
  MUX2_X1 U17704 ( .A(n14107), .B(n14106), .S(n15223), .Z(n15292) );
  INV_X1 U17705 ( .A(n15292), .ZN(n14108) );
  NAND2_X1 U17706 ( .A1(n21071), .A2(n14108), .ZN(n21073) );
  NAND2_X1 U17707 ( .A1(n14112), .A2(P1_UWORD_REG_9__SCAN_IN), .ZN(n14109) );
  OAI211_X1 U17708 ( .C1(n14169), .C2(n15229), .A(n21073), .B(n14109), .ZN(
        P1_U2946) );
  INV_X1 U17709 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n21043) );
  INV_X1 U17710 ( .A(DATAI_8_), .ZN(n14110) );
  INV_X1 U17711 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n21684) );
  MUX2_X1 U17712 ( .A(n14110), .B(n21684), .S(n15223), .Z(n15294) );
  INV_X1 U17713 ( .A(n15294), .ZN(n14111) );
  NAND2_X1 U17714 ( .A1(n21071), .A2(n14111), .ZN(n14115) );
  NAND2_X1 U17715 ( .A1(n14112), .A2(P1_LWORD_REG_8__SCAN_IN), .ZN(n14113) );
  OAI211_X1 U17716 ( .C1(n21043), .C2(n14169), .A(n14115), .B(n14113), .ZN(
        P1_U2960) );
  NAND2_X1 U17717 ( .A1(n21077), .A2(P1_UWORD_REG_8__SCAN_IN), .ZN(n14114) );
  OAI211_X1 U17718 ( .C1(n15234), .C2(n14169), .A(n14115), .B(n14114), .ZN(
        P1_U2945) );
  INV_X1 U17719 ( .A(n14082), .ZN(n14117) );
  OAI21_X1 U17720 ( .B1(n14117), .B2(n10639), .A(n14116), .ZN(n17412) );
  AOI22_X1 U17721 ( .A1(n16869), .A2(n16792), .B1(P2_EAX_REG_8__SCAN_IN), .B2(
        n16867), .ZN(n14118) );
  OAI21_X1 U17722 ( .B1(n17412), .B2(n16864), .A(n14118), .ZN(P2_U2911) );
  INV_X1 U17723 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n14120) );
  AOI22_X1 U17724 ( .A1(P1_UWORD_REG_1__SCAN_IN), .A2(n21054), .B1(n21053), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n14119) );
  OAI21_X1 U17725 ( .B1(n14120), .B2(n14124), .A(n14119), .ZN(P1_U2919) );
  INV_X1 U17726 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n14122) );
  AOI22_X1 U17727 ( .A1(P1_UWORD_REG_2__SCAN_IN), .A2(n21054), .B1(n21053), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n14121) );
  OAI21_X1 U17728 ( .B1(n14122), .B2(n14124), .A(n14121), .ZN(P1_U2918) );
  INV_X1 U17729 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n14125) );
  AOI22_X1 U17730 ( .A1(P1_UWORD_REG_0__SCAN_IN), .A2(n21054), .B1(n21053), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n14123) );
  OAI21_X1 U17731 ( .B1(n14125), .B2(n14124), .A(n14123), .ZN(P1_U2920) );
  NAND2_X1 U17732 ( .A1(n10514), .A2(n21532), .ZN(n14126) );
  OAI21_X1 U17733 ( .B1(n12622), .B2(n14126), .A(n14433), .ZN(n14127) );
  INV_X1 U17734 ( .A(n14127), .ZN(n14128) );
  OAI21_X1 U17735 ( .B1(n14822), .B2(n14131), .A(n14130), .ZN(n14132) );
  NAND2_X1 U17736 ( .A1(n14132), .A2(n20935), .ZN(n14133) );
  AND2_X1 U17737 ( .A1(n12571), .A2(n14385), .ZN(n14139) );
  INV_X1 U17738 ( .A(n14139), .ZN(n14135) );
  AND2_X1 U17739 ( .A1(n14136), .A2(n14135), .ZN(n14137) );
  NAND2_X1 U17740 ( .A1(n14801), .A2(DATAI_0_), .ZN(n14141) );
  NAND2_X1 U17741 ( .A1(n15223), .A2(BUF1_REG_0__SCAN_IN), .ZN(n14140) );
  AND2_X1 U17742 ( .A1(n14141), .A2(n14140), .ZN(n15271) );
  INV_X1 U17743 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n21059) );
  OAI222_X1 U17744 ( .A1(n15171), .A2(n15298), .B1(n15296), .B2(n15271), .C1(
        n14816), .C2(n21059), .ZN(P1_U2904) );
  NAND2_X1 U17745 ( .A1(n14801), .A2(DATAI_1_), .ZN(n14143) );
  NAND2_X1 U17746 ( .A1(n15223), .A2(BUF1_REG_1__SCAN_IN), .ZN(n14142) );
  AND2_X1 U17747 ( .A1(n14143), .A2(n14142), .ZN(n15266) );
  INV_X1 U17748 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n21056) );
  OAI222_X1 U17749 ( .A1(n15164), .A2(n15298), .B1(n15296), .B2(n15266), .C1(
        n14816), .C2(n21056), .ZN(P1_U2903) );
  INV_X1 U17750 ( .A(n14144), .ZN(n14145) );
  OAI21_X1 U17751 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n12674), .A(
        n14145), .ZN(n15166) );
  INV_X1 U17752 ( .A(n15166), .ZN(n14150) );
  INV_X1 U17753 ( .A(n14146), .ZN(n14149) );
  INV_X1 U17754 ( .A(n21117), .ZN(n15739) );
  NOR2_X1 U17755 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n15739), .ZN(
        n14147) );
  AOI21_X1 U17756 ( .B1(n15739), .B2(n21118), .A(n21119), .ZN(n21145) );
  AOI22_X1 U17757 ( .A1(n14147), .A2(n15589), .B1(n15611), .B2(n21145), .ZN(
        n14148) );
  AOI211_X1 U17758 ( .C1(n14150), .C2(n21135), .A(n14149), .B(n14148), .ZN(
        n14151) );
  OAI21_X1 U17759 ( .B1(n21139), .B2(n14152), .A(n14151), .ZN(P1_U3031) );
  NAND3_X1 U17760 ( .A1(n20018), .A2(n20161), .A3(n14153), .ZN(n14322) );
  NAND2_X1 U17761 ( .A1(n14155), .A2(n14154), .ZN(n14156) );
  INV_X1 U17762 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n18980) );
  INV_X1 U17763 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n18978) );
  INV_X1 U17764 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n18976) );
  INV_X1 U17765 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n14256) );
  NAND2_X1 U17766 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(P3_EAX_REG_0__SCAN_IN), 
        .ZN(n14255) );
  NOR2_X1 U17767 ( .A1(n14256), .A2(n14255), .ZN(n14232) );
  NAND4_X1 U17768 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n14232), .A3(
        P3_EAX_REG_4__SCAN_IN), .A4(P3_EAX_REG_3__SCAN_IN), .ZN(n14237) );
  NOR3_X1 U17769 ( .A1(n18978), .A2(n18976), .A3(n14237), .ZN(n18892) );
  AOI22_X1 U17770 ( .A1(n18886), .A2(P3_EAX_REG_9__SCAN_IN), .B1(n19588), .B2(
        n18878), .ZN(n14158) );
  AND2_X1 U17771 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n18878), .ZN(n14157) );
  NAND2_X1 U17772 ( .A1(n19588), .A2(n14157), .ZN(n18875) );
  INV_X1 U17773 ( .A(n18875), .ZN(n17733) );
  OAI222_X1 U17774 ( .A1(n18883), .A2(n13646), .B1(n18832), .B2(n14159), .C1(
        n14158), .C2(n17733), .ZN(P3_U2726) );
  AND2_X1 U17775 ( .A1(n9682), .A2(n19588), .ZN(n18891) );
  INV_X1 U17776 ( .A(n18891), .ZN(n18789) );
  INV_X1 U17777 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n18966) );
  OAI22_X1 U17778 ( .A1(n18789), .A2(P3_EAX_REG_0__SCAN_IN), .B1(n9682), .B2(
        n18966), .ZN(n14160) );
  AOI21_X1 U17779 ( .B1(n18888), .B2(n14161), .A(n14160), .ZN(n14162) );
  OAI21_X1 U17780 ( .B1(n14163), .B2(n18883), .A(n14162), .ZN(P3_U2735) );
  INV_X1 U17781 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n14165) );
  OAI211_X1 U17782 ( .C1(P3_EAX_REG_1__SCAN_IN), .C2(P3_EAX_REG_0__SCAN_IN), 
        .A(n18891), .B(n14255), .ZN(n14164) );
  OAI21_X1 U17783 ( .B1(n9682), .B2(n14165), .A(n14164), .ZN(n14166) );
  AOI21_X1 U17784 ( .B1(n18888), .B2(n14167), .A(n14166), .ZN(n14168) );
  OAI21_X1 U17785 ( .B1(n13632), .B2(n18883), .A(n14168), .ZN(P3_U2734) );
  AOI22_X1 U17786 ( .A1(n21084), .A2(P1_EAX_REG_21__SCAN_IN), .B1(
        P1_UWORD_REG_5__SCAN_IN), .B2(n14112), .ZN(n14174) );
  NAND2_X1 U17787 ( .A1(n14801), .A2(DATAI_5_), .ZN(n14172) );
  NAND2_X1 U17788 ( .A1(n15223), .A2(BUF1_REG_5__SCAN_IN), .ZN(n14171) );
  AND2_X1 U17789 ( .A1(n14172), .A2(n14171), .ZN(n15246) );
  INV_X1 U17790 ( .A(n15246), .ZN(n14173) );
  NAND2_X1 U17791 ( .A1(n21071), .A2(n14173), .ZN(n14194) );
  NAND2_X1 U17792 ( .A1(n14174), .A2(n14194), .ZN(P1_U2942) );
  AOI22_X1 U17793 ( .A1(n21084), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_UWORD_REG_0__SCAN_IN), .B2(n14112), .ZN(n14176) );
  INV_X1 U17794 ( .A(n15271), .ZN(n14175) );
  NAND2_X1 U17795 ( .A1(n21071), .A2(n14175), .ZN(n14181) );
  NAND2_X1 U17796 ( .A1(n14176), .A2(n14181), .ZN(P1_U2937) );
  AOI22_X1 U17797 ( .A1(n21084), .A2(P1_EAX_REG_20__SCAN_IN), .B1(
        P1_UWORD_REG_4__SCAN_IN), .B2(n14112), .ZN(n14180) );
  NAND2_X1 U17798 ( .A1(n14801), .A2(DATAI_4_), .ZN(n14178) );
  NAND2_X1 U17799 ( .A1(n15223), .A2(BUF1_REG_4__SCAN_IN), .ZN(n14177) );
  AND2_X1 U17800 ( .A1(n14178), .A2(n14177), .ZN(n15251) );
  INV_X1 U17801 ( .A(n15251), .ZN(n14179) );
  NAND2_X1 U17802 ( .A1(n21071), .A2(n14179), .ZN(n14202) );
  NAND2_X1 U17803 ( .A1(n14180), .A2(n14202), .ZN(P1_U2941) );
  AOI22_X1 U17804 ( .A1(n21084), .A2(P1_EAX_REG_0__SCAN_IN), .B1(
        P1_LWORD_REG_0__SCAN_IN), .B2(n21077), .ZN(n14182) );
  NAND2_X1 U17805 ( .A1(n14182), .A2(n14181), .ZN(P1_U2952) );
  AOI22_X1 U17806 ( .A1(n21084), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_UWORD_REG_2__SCAN_IN), .B2(n21077), .ZN(n14186) );
  NAND2_X1 U17807 ( .A1(n14801), .A2(DATAI_2_), .ZN(n14184) );
  NAND2_X1 U17808 ( .A1(n15223), .A2(BUF1_REG_2__SCAN_IN), .ZN(n14183) );
  AND2_X1 U17809 ( .A1(n14184), .A2(n14183), .ZN(n15261) );
  INV_X1 U17810 ( .A(n15261), .ZN(n14185) );
  NAND2_X1 U17811 ( .A1(n21071), .A2(n14185), .ZN(n14196) );
  NAND2_X1 U17812 ( .A1(n14186), .A2(n14196), .ZN(P1_U2939) );
  AOI22_X1 U17813 ( .A1(n21084), .A2(P1_EAX_REG_17__SCAN_IN), .B1(
        P1_UWORD_REG_1__SCAN_IN), .B2(n21077), .ZN(n14188) );
  INV_X1 U17814 ( .A(n15266), .ZN(n14187) );
  NAND2_X1 U17815 ( .A1(n21071), .A2(n14187), .ZN(n14212) );
  NAND2_X1 U17816 ( .A1(n14188), .A2(n14212), .ZN(P1_U2938) );
  AOI22_X1 U17817 ( .A1(n21084), .A2(P1_EAX_REG_19__SCAN_IN), .B1(
        P1_UWORD_REG_3__SCAN_IN), .B2(n21077), .ZN(n14191) );
  INV_X1 U17818 ( .A(DATAI_3_), .ZN(n14190) );
  NAND2_X1 U17819 ( .A1(n15223), .A2(BUF1_REG_3__SCAN_IN), .ZN(n14189) );
  OAI21_X1 U17820 ( .B1(n15223), .B2(n14190), .A(n14189), .ZN(n15255) );
  NAND2_X1 U17821 ( .A1(n21071), .A2(n15255), .ZN(n14192) );
  NAND2_X1 U17822 ( .A1(n14191), .A2(n14192), .ZN(P1_U2940) );
  AOI22_X1 U17823 ( .A1(n21084), .A2(P1_EAX_REG_3__SCAN_IN), .B1(
        P1_LWORD_REG_3__SCAN_IN), .B2(n21077), .ZN(n14193) );
  NAND2_X1 U17824 ( .A1(n14193), .A2(n14192), .ZN(P1_U2955) );
  AOI22_X1 U17825 ( .A1(n21084), .A2(P1_EAX_REG_5__SCAN_IN), .B1(
        P1_LWORD_REG_5__SCAN_IN), .B2(n21077), .ZN(n14195) );
  NAND2_X1 U17826 ( .A1(n14195), .A2(n14194), .ZN(P1_U2957) );
  AOI22_X1 U17827 ( .A1(n21084), .A2(P1_EAX_REG_2__SCAN_IN), .B1(
        P1_LWORD_REG_2__SCAN_IN), .B2(n21077), .ZN(n14197) );
  NAND2_X1 U17828 ( .A1(n14197), .A2(n14196), .ZN(P1_U2954) );
  AOI22_X1 U17829 ( .A1(n21084), .A2(P1_EAX_REG_23__SCAN_IN), .B1(
        P1_UWORD_REG_7__SCAN_IN), .B2(n21077), .ZN(n14201) );
  NAND2_X1 U17830 ( .A1(n14801), .A2(DATAI_7_), .ZN(n14199) );
  NAND2_X1 U17831 ( .A1(n15223), .A2(BUF1_REG_7__SCAN_IN), .ZN(n14198) );
  AND2_X1 U17832 ( .A1(n14199), .A2(n14198), .ZN(n15297) );
  INV_X1 U17833 ( .A(n15297), .ZN(n14200) );
  NAND2_X1 U17834 ( .A1(n21071), .A2(n14200), .ZN(n14204) );
  NAND2_X1 U17835 ( .A1(n14201), .A2(n14204), .ZN(P1_U2944) );
  AOI22_X1 U17836 ( .A1(n21084), .A2(P1_EAX_REG_4__SCAN_IN), .B1(
        P1_LWORD_REG_4__SCAN_IN), .B2(n21077), .ZN(n14203) );
  NAND2_X1 U17837 ( .A1(n14203), .A2(n14202), .ZN(P1_U2956) );
  AOI22_X1 U17838 ( .A1(n21084), .A2(P1_EAX_REG_7__SCAN_IN), .B1(
        P1_LWORD_REG_7__SCAN_IN), .B2(n21077), .ZN(n14205) );
  NAND2_X1 U17839 ( .A1(n14205), .A2(n14204), .ZN(P1_U2959) );
  AOI22_X1 U17840 ( .A1(n21084), .A2(P1_EAX_REG_6__SCAN_IN), .B1(
        P1_LWORD_REG_6__SCAN_IN), .B2(n21077), .ZN(n14209) );
  NAND2_X1 U17841 ( .A1(n14801), .A2(DATAI_6_), .ZN(n14207) );
  NAND2_X1 U17842 ( .A1(n15223), .A2(BUF1_REG_6__SCAN_IN), .ZN(n14206) );
  AND2_X1 U17843 ( .A1(n14207), .A2(n14206), .ZN(n15242) );
  INV_X1 U17844 ( .A(n15242), .ZN(n14208) );
  NAND2_X1 U17845 ( .A1(n21071), .A2(n14208), .ZN(n14210) );
  NAND2_X1 U17846 ( .A1(n14209), .A2(n14210), .ZN(P1_U2958) );
  AOI22_X1 U17847 ( .A1(n21084), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_UWORD_REG_6__SCAN_IN), .B2(n21077), .ZN(n14211) );
  NAND2_X1 U17848 ( .A1(n14211), .A2(n14210), .ZN(P1_U2943) );
  AOI22_X1 U17849 ( .A1(n21084), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_LWORD_REG_1__SCAN_IN), .B2(n21077), .ZN(n14213) );
  NAND2_X1 U17850 ( .A1(n14213), .A2(n14212), .ZN(P1_U2953) );
  OAI21_X1 U17851 ( .B1(n17642), .B2(n20900), .A(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n14219) );
  INV_X1 U17852 ( .A(n17642), .ZN(n20604) );
  NAND2_X1 U17853 ( .A1(n21853), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n20384) );
  INV_X1 U17854 ( .A(n20384), .ZN(n20437) );
  NAND2_X1 U17855 ( .A1(n20604), .A2(n20437), .ZN(n20469) );
  NAND2_X1 U17856 ( .A1(n14219), .A2(n20469), .ZN(n14220) );
  AOI22_X1 U17857 ( .A1(n14221), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n20888), .B2(n14220), .ZN(n14222) );
  NAND2_X1 U17858 ( .A1(n14223), .A2(n14222), .ZN(n14225) );
  OAI21_X1 U17859 ( .B1(n14225), .B2(n14224), .A(n14284), .ZN(n14226) );
  MUX2_X1 U17860 ( .A(n11004), .B(n14230), .S(n16728), .Z(n14231) );
  OAI21_X1 U17861 ( .B1(n20535), .B2(n16733), .A(n14231), .ZN(P2_U2884) );
  AND2_X1 U17862 ( .A1(n18891), .A2(n14232), .ZN(n14254) );
  AOI22_X1 U17863 ( .A1(n14254), .A2(P3_EAX_REG_3__SCAN_IN), .B1(
        P3_EAX_REG_4__SCAN_IN), .B2(n18886), .ZN(n14234) );
  NAND2_X1 U17864 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(P3_EAX_REG_3__SCAN_IN), 
        .ZN(n14233) );
  INV_X1 U17865 ( .A(n14254), .ZN(n14298) );
  NOR2_X1 U17866 ( .A1(n14233), .A2(n14298), .ZN(n14236) );
  OAI222_X1 U17867 ( .A1(n18832), .A2(n14235), .B1(n18883), .B2(n13649), .C1(
        n14234), .C2(n14236), .ZN(P3_U2731) );
  AOI21_X1 U17868 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n18886), .A(n14236), .ZN(
        n14238) );
  NOR2_X1 U17869 ( .A1(n18789), .A2(n14237), .ZN(n14240) );
  OAI222_X1 U17870 ( .A1(n18832), .A2(n14239), .B1(n18883), .B2(n13643), .C1(
        n14238), .C2(n14240), .ZN(P3_U2730) );
  AOI21_X1 U17871 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n18886), .A(n14240), .ZN(
        n14242) );
  INV_X1 U17872 ( .A(n14240), .ZN(n14241) );
  NOR2_X1 U17873 ( .A1(n14241), .A2(n18976), .ZN(n18885) );
  OAI222_X1 U17874 ( .A1(n18832), .A2(n14243), .B1(n18883), .B2(n13635), .C1(
        n14242), .C2(n18885), .ZN(P3_U2729) );
  OAI222_X1 U17875 ( .A1(n15166), .A2(n15203), .B1(n12635), .B2(n15204), .C1(
        n15171), .C2(n15206), .ZN(P1_U2872) );
  INV_X1 U17876 ( .A(n16785), .ZN(n14246) );
  NAND2_X1 U17877 ( .A1(n14116), .A2(n14244), .ZN(n14245) );
  NAND2_X1 U17878 ( .A1(n14359), .A2(n14245), .ZN(n17393) );
  INV_X1 U17879 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n20227) );
  OAI222_X1 U17880 ( .A1(n14763), .A2(n14246), .B1(n17393), .B2(n16864), .C1(
        n20227), .C2(n16744), .ZN(P2_U2910) );
  NAND2_X1 U17881 ( .A1(n17513), .A2(n14249), .ZN(n14346) );
  OAI21_X1 U17882 ( .B1(n17513), .B2(n14249), .A(n14346), .ZN(n14247) );
  NOR2_X1 U17883 ( .A1(n14247), .A2(n14248), .ZN(n14348) );
  AOI21_X1 U17884 ( .B1(n14248), .B2(n14247), .A(n14348), .ZN(n14252) );
  OAI22_X1 U17885 ( .A1(n14249), .A2(n16855), .B1(n16744), .B2(n11224), .ZN(
        n14250) );
  AOI21_X1 U17886 ( .B1(n16869), .B2(n17558), .A(n14250), .ZN(n14251) );
  OAI21_X1 U17887 ( .B1(n14252), .B2(n16872), .A(n14251), .ZN(P2_U2918) );
  INV_X1 U17888 ( .A(n9682), .ZN(n14257) );
  AOI221_X1 U17889 ( .B1(n14257), .B2(n14256), .C1(n14255), .C2(n14256), .A(
        n14254), .ZN(n14258) );
  INV_X1 U17890 ( .A(n14258), .ZN(n14259) );
  OAI222_X1 U17891 ( .A1(n18832), .A2(n14260), .B1(n14259), .B2(n18877), .C1(
        n18883), .C2(n13655), .ZN(P3_U2733) );
  NAND2_X1 U17892 ( .A1(n14263), .A2(n14262), .ZN(n14264) );
  AND2_X1 U17893 ( .A1(n14261), .A2(n14264), .ZN(n21017) );
  INV_X1 U17894 ( .A(n21017), .ZN(n14282) );
  NAND2_X1 U17895 ( .A1(n14266), .A2(n14265), .ZN(n14267) );
  NAND2_X1 U17896 ( .A1(n14270), .A2(n14267), .ZN(n21124) );
  INV_X1 U17897 ( .A(n21124), .ZN(n14268) );
  AOI22_X1 U17898 ( .A1(n15196), .A2(n14268), .B1(P1_EBX_REG_2__SCAN_IN), .B2(
        n15195), .ZN(n14269) );
  OAI21_X1 U17899 ( .B1(n14282), .B2(n15206), .A(n14269), .ZN(P1_U2870) );
  INV_X1 U17900 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n21052) );
  OAI222_X1 U17901 ( .A1(n14282), .A2(n15298), .B1(n15261), .B2(n15296), .C1(
        n14816), .C2(n21052), .ZN(P1_U2902) );
  XNOR2_X1 U17902 ( .A(n14411), .B(n14412), .ZN(n15510) );
  AOI21_X1 U17903 ( .B1(n14271), .B2(n14270), .A(n14417), .ZN(n21111) );
  AOI22_X1 U17904 ( .A1(n15196), .A2(n21111), .B1(P1_EBX_REG_3__SCAN_IN), .B2(
        n15195), .ZN(n14272) );
  OAI21_X1 U17905 ( .B1(n15510), .B2(n15206), .A(n14272), .ZN(P1_U2869) );
  NOR2_X1 U17906 ( .A1(n14274), .A2(n14273), .ZN(n21122) );
  INV_X1 U17907 ( .A(n21122), .ZN(n14276) );
  NAND3_X1 U17908 ( .A1(n14276), .A2(n21095), .A3(n14275), .ZN(n14281) );
  INV_X1 U17909 ( .A(n15496), .ZN(n21123) );
  INV_X1 U17910 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n14277) );
  OAI22_X1 U17911 ( .A1(n15504), .A2(n14278), .B1(n21123), .B2(n14277), .ZN(
        n14279) );
  AOI21_X1 U17912 ( .B1(n15507), .B2(n21028), .A(n14279), .ZN(n14280) );
  OAI211_X1 U17913 ( .C1(n15511), .C2(n14282), .A(n14281), .B(n14280), .ZN(
        P1_U2997) );
  NAND2_X1 U17914 ( .A1(n17537), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n14283) );
  AND2_X1 U17915 ( .A1(n16536), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n14286) );
  OR2_X1 U17916 ( .A1(n16367), .A2(n14286), .ZN(n14287) );
  NAND2_X1 U17917 ( .A1(n14506), .A2(n14287), .ZN(n20198) );
  AND2_X1 U17918 ( .A1(n14290), .A2(n14289), .ZN(n14291) );
  OR2_X1 U17919 ( .A1(n14288), .A2(n14291), .ZN(n20258) );
  MUX2_X1 U17920 ( .A(n20258), .B(n14292), .S(n16723), .Z(n14293) );
  OAI21_X1 U17921 ( .B1(n20198), .B2(n16733), .A(n14293), .ZN(P2_U2883) );
  NAND2_X1 U17922 ( .A1(n14298), .A2(P3_EAX_REG_3__SCAN_IN), .ZN(n14294) );
  OAI22_X1 U17923 ( .A1(n18832), .A2(n14295), .B1(n18877), .B2(n14294), .ZN(
        n14296) );
  AOI21_X1 U17924 ( .B1(n18889), .B2(BUF2_REG_3__SCAN_IN), .A(n14296), .ZN(
        n14297) );
  OAI21_X1 U17925 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n14298), .A(n14297), .ZN(
        P3_U2732) );
  INV_X1 U17926 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n18997) );
  INV_X1 U17927 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n18917) );
  INV_X1 U17928 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n18986) );
  INV_X1 U17929 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n18984) );
  INV_X1 U17930 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n18982) );
  NOR4_X1 U17931 ( .A1(n18917), .A2(n18986), .A3(n18984), .A4(n18982), .ZN(
        n14299) );
  AOI211_X1 U17932 ( .C1(n18997), .C2(n18865), .A(n18877), .B(n18860), .ZN(
        n14300) );
  AOI21_X1 U17933 ( .B1(n18889), .B2(BUF2_REG_15__SCAN_IN), .A(n14300), .ZN(
        n14301) );
  OAI21_X1 U17934 ( .B1(n14302), .B2(n18832), .A(n14301), .ZN(P3_U2720) );
  OAI21_X1 U17935 ( .B1(n14304), .B2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n14303), .ZN(n21140) );
  INV_X1 U17936 ( .A(n21140), .ZN(n14306) );
  MUX2_X1 U17937 ( .A(n15507), .B(n21088), .S(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .Z(n14305) );
  AND2_X1 U17938 ( .A1(n15496), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n21133) );
  AOI211_X1 U17939 ( .C1(n14306), .C2(n21095), .A(n14305), .B(n21133), .ZN(
        n14307) );
  OAI21_X1 U17940 ( .B1(n15511), .B2(n15164), .A(n14307), .ZN(P1_U2998) );
  INV_X1 U17941 ( .A(n15255), .ZN(n14308) );
  INV_X1 U17942 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n21050) );
  OAI222_X1 U17943 ( .A1(n15510), .A2(n15298), .B1(n15296), .B2(n14308), .C1(
        n14816), .C2(n21050), .ZN(P1_U2901) );
  INV_X1 U17944 ( .A(n14309), .ZN(n14315) );
  NAND2_X1 U17945 ( .A1(n14311), .A2(n14310), .ZN(n14314) );
  OAI211_X1 U17946 ( .C1(n14313), .C2(n14315), .A(n14312), .B(n14314), .ZN(
        n14736) );
  NAND3_X1 U17947 ( .A1(n14316), .A2(n14315), .A3(n14314), .ZN(n14317) );
  NOR2_X1 U17948 ( .A1(n14720), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n14329) );
  AOI21_X1 U17949 ( .B1(n14317), .B2(n14732), .A(n14329), .ZN(n14318) );
  NAND2_X1 U17950 ( .A1(n14319), .A2(n14318), .ZN(n20009) );
  NOR2_X1 U17951 ( .A1(n20022), .A2(n14320), .ZN(n14326) );
  NAND2_X1 U17952 ( .A1(n20018), .A2(n20161), .ZN(n14324) );
  OAI21_X1 U17953 ( .B1(n14321), .B2(n20041), .A(n20149), .ZN(n18894) );
  OAI211_X1 U17954 ( .C1(n14324), .C2(n18894), .A(n14323), .B(n14322), .ZN(
        n14325) );
  INV_X1 U17955 ( .A(n20026), .ZN(n19999) );
  INV_X1 U17956 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n19553) );
  NAND2_X1 U17957 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n20159), .ZN(n20133) );
  NOR2_X1 U17958 ( .A1(n19553), .A2(n20133), .ZN(n14327) );
  NOR2_X1 U17959 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n20134), .ZN(n19564) );
  AOI21_X1 U17960 ( .B1(n17979), .B2(n20009), .A(n14748), .ZN(n14339) );
  NAND2_X1 U17961 ( .A1(n19428), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n14328) );
  NAND2_X1 U17962 ( .A1(n14328), .A2(n19314), .ZN(n14734) );
  NAND2_X1 U17963 ( .A1(n14734), .A2(n14333), .ZN(n14331) );
  INV_X1 U17964 ( .A(n14329), .ZN(n14730) );
  NAND2_X1 U17965 ( .A1(n20023), .A2(n14730), .ZN(n14330) );
  NAND2_X1 U17966 ( .A1(n14331), .A2(n14330), .ZN(n14332) );
  NAND2_X1 U17967 ( .A1(n14332), .A2(n14338), .ZN(n20010) );
  INV_X1 U17968 ( .A(n17979), .ZN(n18577) );
  NAND2_X1 U17969 ( .A1(n14333), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n14729) );
  NAND2_X1 U17970 ( .A1(n14729), .A2(n14338), .ZN(n14334) );
  NAND2_X1 U17971 ( .A1(n14335), .A2(n14334), .ZN(n18535) );
  OAI22_X1 U17972 ( .A1(n20010), .A2(n18577), .B1(n14744), .B2(n18535), .ZN(
        n14336) );
  INV_X1 U17973 ( .A(n14336), .ZN(n14337) );
  OAI22_X1 U17974 ( .A1(n14339), .A2(n14338), .B1(n14748), .B2(n14337), .ZN(
        P3_U3285) );
  XOR2_X1 U17975 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B(n14506), .Z(n14345)
         );
  OR2_X1 U17976 ( .A1(n14288), .A2(n14341), .ZN(n14342) );
  NAND2_X1 U17977 ( .A1(n14340), .A2(n14342), .ZN(n17434) );
  INV_X1 U17978 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n14343) );
  MUX2_X1 U17979 ( .A(n17434), .B(n14343), .S(n16723), .Z(n14344) );
  OAI21_X1 U17980 ( .B1(n14345), .B2(n16733), .A(n14344), .ZN(P2_U2882) );
  INV_X1 U17981 ( .A(n14346), .ZN(n14347) );
  NOR2_X1 U17982 ( .A1(n14348), .A2(n14347), .ZN(n14354) );
  OR2_X1 U17983 ( .A1(n14350), .A2(n14349), .ZN(n14351) );
  NAND2_X1 U17984 ( .A1(n14352), .A2(n14351), .ZN(n20276) );
  INV_X1 U17985 ( .A(n20276), .ZN(n20894) );
  NAND2_X1 U17986 ( .A1(n20896), .A2(n20894), .ZN(n14558) );
  OAI21_X1 U17987 ( .B1(n20896), .B2(n20894), .A(n14558), .ZN(n14353) );
  NOR2_X1 U17988 ( .A1(n14354), .A2(n14353), .ZN(n14560) );
  AOI21_X1 U17989 ( .B1(n14354), .B2(n14353), .A(n14560), .ZN(n14357) );
  OAI22_X1 U17990 ( .A1(n20894), .A2(n16855), .B1(n16744), .B2(n21726), .ZN(
        n14355) );
  AOI21_X1 U17991 ( .B1(n16869), .B2(n17563), .A(n14355), .ZN(n14356) );
  OAI21_X1 U17992 ( .B1(n14357), .B2(n16872), .A(n14356), .ZN(P2_U2917) );
  AND2_X1 U17993 ( .A1(n14359), .A2(n14358), .ZN(n14360) );
  NOR2_X1 U17994 ( .A1(n9782), .A2(n14360), .ZN(n17389) );
  INV_X1 U17995 ( .A(n17389), .ZN(n16248) );
  AOI22_X1 U17996 ( .A1(n16869), .A2(n16778), .B1(P2_EAX_REG_10__SCAN_IN), 
        .B2(n16867), .ZN(n14361) );
  OAI21_X1 U17997 ( .B1(n16248), .B2(n16864), .A(n14361), .ZN(P2_U2909) );
  NOR2_X2 U17998 ( .A1(n15511), .A2(n15223), .ZN(n14400) );
  AOI22_X1 U17999 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n14401), .B1(DATAI_27_), 
        .B2(n14400), .ZN(n21496) );
  NAND3_X1 U18000 ( .A1(n9709), .A2(n14362), .A3(n14363), .ZN(n14373) );
  AOI22_X1 U18001 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n14401), .B1(DATAI_19_), 
        .B2(n14400), .ZN(n21439) );
  OR2_X1 U18002 ( .A1(n14367), .A2(n14366), .ZN(n14368) );
  NAND2_X1 U18003 ( .A1(n15792), .A2(n14457), .ZN(n21467) );
  NOR2_X1 U18004 ( .A1(n21467), .A2(n21417), .ZN(n21415) );
  OR2_X1 U18005 ( .A1(n15165), .A2(n11944), .ZN(n21236) );
  INV_X1 U18006 ( .A(n21236), .ZN(n14526) );
  NOR2_X1 U18007 ( .A1(n21681), .A2(n21464), .ZN(n14374) );
  INV_X1 U18008 ( .A(n14374), .ZN(n14369) );
  OAI22_X1 U18009 ( .A1(n14404), .A2(n21417), .B1(n14369), .B2(n21349), .ZN(
        n14370) );
  AOI21_X1 U18010 ( .B1(n21415), .B2(n14526), .A(n14370), .ZN(n14405) );
  OAI21_X1 U18011 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(
        P1_STATE2_REG_1__SCAN_IN), .A(n20939), .ZN(n21619) );
  AND2_X1 U18012 ( .A1(n15255), .A2(n15818), .ZN(n21492) );
  NAND2_X1 U18013 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n15818), .ZN(n14389) );
  OAI22_X1 U18014 ( .A1(n14405), .A2(n21400), .B1(n14404), .B2(n21321), .ZN(
        n14371) );
  AOI21_X1 U18015 ( .B1(n15790), .B2(n21493), .A(n14371), .ZN(n14377) );
  INV_X1 U18016 ( .A(n14372), .ZN(n21420) );
  NOR2_X1 U18017 ( .A1(n14373), .A2(n21420), .ZN(n14375) );
  NAND2_X1 U18018 ( .A1(n14407), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n14376) );
  OAI211_X1 U18019 ( .C1(n21496), .C2(n21476), .A(n14377), .B(n14376), .ZN(
        P1_U3156) );
  AOI22_X1 U18020 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n14401), .B1(DATAI_24_), 
        .B2(n14400), .ZN(n21480) );
  AOI22_X1 U18021 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n14401), .B1(DATAI_16_), 
        .B2(n14400), .ZN(n21428) );
  INV_X1 U18022 ( .A(n21428), .ZN(n21477) );
  NAND2_X1 U18023 ( .A1(n12634), .A2(n14402), .ZN(n21303) );
  OAI22_X1 U18024 ( .A1(n14405), .A2(n21394), .B1(n14404), .B2(n21303), .ZN(
        n14378) );
  AOI21_X1 U18025 ( .B1(n15790), .B2(n21477), .A(n14378), .ZN(n14380) );
  NAND2_X1 U18026 ( .A1(n14407), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n14379) );
  OAI211_X1 U18027 ( .C1(n21480), .C2(n21476), .A(n14380), .B(n14379), .ZN(
        P1_U3153) );
  AOI22_X1 U18028 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n14401), .B1(DATAI_26_), 
        .B2(n14400), .ZN(n21490) );
  AOI22_X1 U18029 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n14401), .B1(DATAI_18_), 
        .B2(n14400), .ZN(n21435) );
  INV_X1 U18030 ( .A(n21435), .ZN(n21931) );
  INV_X1 U18031 ( .A(n21928), .ZN(n21317) );
  OAI22_X1 U18032 ( .A1(n14405), .A2(n21936), .B1(n14404), .B2(n21317), .ZN(
        n14382) );
  AOI21_X1 U18033 ( .B1(n15790), .B2(n21931), .A(n14382), .ZN(n14384) );
  NAND2_X1 U18034 ( .A1(n14407), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n14383) );
  OAI211_X1 U18035 ( .C1(n21490), .C2(n21476), .A(n14384), .B(n14383), .ZN(
        P1_U3155) );
  AOI22_X1 U18036 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n14401), .B1(DATAI_31_), 
        .B2(n14400), .ZN(n21525) );
  AOI22_X1 U18037 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n14401), .B1(DATAI_23_), 
        .B2(n14400), .ZN(n21459) );
  INV_X1 U18038 ( .A(n21459), .ZN(n21519) );
  OAI22_X1 U18039 ( .A1(n14405), .A2(n21412), .B1(n14404), .B2(n21337), .ZN(
        n14386) );
  AOI21_X1 U18040 ( .B1(n15790), .B2(n21519), .A(n14386), .ZN(n14388) );
  NAND2_X1 U18041 ( .A1(n14407), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n14387) );
  OAI211_X1 U18042 ( .C1(n21525), .C2(n21476), .A(n14388), .B(n14387), .ZN(
        P1_U3160) );
  AOI22_X1 U18043 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n14401), .B1(DATAI_25_), 
        .B2(n14400), .ZN(n21486) );
  AOI22_X1 U18044 ( .A1(DATAI_17_), .A2(n14400), .B1(BUF1_REG_17__SCAN_IN), 
        .B2(n14401), .ZN(n21432) );
  INV_X1 U18045 ( .A(n21432), .ZN(n21483) );
  OR2_X1 U18046 ( .A1(n13450), .A2(n14389), .ZN(n21313) );
  OAI22_X1 U18047 ( .A1(n14405), .A2(n21397), .B1(n14404), .B2(n21313), .ZN(
        n14391) );
  AOI21_X1 U18048 ( .B1(n15790), .B2(n21483), .A(n14391), .ZN(n14393) );
  NAND2_X1 U18049 ( .A1(n14407), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n14392) );
  OAI211_X1 U18050 ( .C1(n21486), .C2(n21476), .A(n14393), .B(n14392), .ZN(
        P1_U3154) );
  AOI22_X1 U18051 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n14401), .B1(DATAI_30_), 
        .B2(n14400), .ZN(n21514) );
  AOI22_X1 U18052 ( .A1(DATAI_22_), .A2(n14400), .B1(BUF1_REG_22__SCAN_IN), 
        .B2(n14401), .ZN(n21451) );
  NAND2_X1 U18053 ( .A1(n11861), .A2(n14402), .ZN(n21333) );
  OAI22_X1 U18054 ( .A1(n14405), .A2(n21409), .B1(n14404), .B2(n21333), .ZN(
        n14394) );
  AOI21_X1 U18055 ( .B1(n15790), .B2(n21511), .A(n14394), .ZN(n14396) );
  NAND2_X1 U18056 ( .A1(n14407), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n14395) );
  OAI211_X1 U18057 ( .C1(n21514), .C2(n21476), .A(n14396), .B(n14395), .ZN(
        P1_U3159) );
  AOI22_X1 U18058 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n14401), .B1(DATAI_28_), 
        .B2(n14400), .ZN(n21502) );
  AOI22_X1 U18059 ( .A1(DATAI_20_), .A2(n14400), .B1(BUF1_REG_20__SCAN_IN), 
        .B2(n14401), .ZN(n21443) );
  INV_X1 U18060 ( .A(n21443), .ZN(n21499) );
  INV_X1 U18061 ( .A(n21497), .ZN(n21325) );
  OAI22_X1 U18062 ( .A1(n14405), .A2(n21403), .B1(n14404), .B2(n21325), .ZN(
        n14397) );
  AOI21_X1 U18063 ( .B1(n15790), .B2(n21499), .A(n14397), .ZN(n14399) );
  NAND2_X1 U18064 ( .A1(n14407), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n14398) );
  OAI211_X1 U18065 ( .C1(n21502), .C2(n21476), .A(n14399), .B(n14398), .ZN(
        P1_U3157) );
  AOI22_X1 U18066 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n14401), .B1(DATAI_29_), 
        .B2(n14400), .ZN(n21508) );
  AOI22_X1 U18067 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n14401), .B1(DATAI_21_), 
        .B2(n14400), .ZN(n21447) );
  INV_X1 U18068 ( .A(n21447), .ZN(n21505) );
  OAI22_X1 U18069 ( .A1(n14405), .A2(n21406), .B1(n14404), .B2(n21329), .ZN(
        n14406) );
  AOI21_X1 U18070 ( .B1(n15790), .B2(n21505), .A(n14406), .ZN(n14409) );
  NAND2_X1 U18071 ( .A1(n14407), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n14408) );
  OAI211_X1 U18072 ( .C1(n21508), .C2(n21476), .A(n14409), .B(n14408), .ZN(
        P1_U3158) );
  NAND2_X1 U18073 ( .A1(n14412), .A2(n14411), .ZN(n14414) );
  NAND2_X1 U18074 ( .A1(n14414), .A2(n14413), .ZN(n14415) );
  AND2_X1 U18075 ( .A1(n14410), .A2(n14415), .ZN(n21093) );
  INV_X1 U18076 ( .A(n21093), .ZN(n14419) );
  OAI21_X1 U18077 ( .B1(n14417), .B2(n14416), .A(n14576), .ZN(n21005) );
  INV_X1 U18078 ( .A(n21005), .ZN(n21103) );
  AOI22_X1 U18079 ( .A1(n15196), .A2(n21103), .B1(P1_EBX_REG_4__SCAN_IN), .B2(
        n15195), .ZN(n14418) );
  OAI21_X1 U18080 ( .B1(n14419), .B2(n15206), .A(n14418), .ZN(P1_U2868) );
  INV_X1 U18081 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n21048) );
  OAI222_X1 U18082 ( .A1(n14419), .A2(n15298), .B1(n15251), .B2(n15296), .C1(
        n14816), .C2(n21048), .ZN(P1_U2900) );
  INV_X1 U18083 ( .A(n16772), .ZN(n14420) );
  INV_X1 U18084 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n20223) );
  OAI222_X1 U18085 ( .A1(n14763), .A2(n14420), .B1(n17366), .B2(n16864), .C1(
        n20223), .C2(n16744), .ZN(P2_U2908) );
  INV_X1 U18086 ( .A(n19277), .ZN(n14426) );
  NAND3_X1 U18087 ( .A1(n20049), .A2(n19271), .A3(n19098), .ZN(n14422) );
  AOI21_X1 U18088 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n14422), .A(
        n14421), .ZN(n14424) );
  NAND2_X1 U18089 ( .A1(n19275), .A2(n14425), .ZN(n14423) );
  OAI211_X1 U18090 ( .C1(n14426), .C2(n14425), .A(n14424), .B(n14423), .ZN(
        P3_U2830) );
  AND2_X1 U18091 ( .A1(n14427), .A2(n14410), .ZN(n14429) );
  OR2_X1 U18092 ( .A1(n14429), .A2(n14428), .ZN(n20988) );
  XOR2_X1 U18093 ( .A(n14575), .B(n14576), .Z(n20991) );
  AOI22_X1 U18094 ( .A1(n20991), .A2(n15196), .B1(P1_EBX_REG_5__SCAN_IN), .B2(
        n15195), .ZN(n14430) );
  OAI21_X1 U18095 ( .B1(n20988), .B2(n15206), .A(n14430), .ZN(P1_U2867) );
  NOR2_X1 U18096 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n18052), .ZN(n14462) );
  XNOR2_X1 U18097 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n15783), .ZN(
        n14431) );
  NOR2_X1 U18098 ( .A1(n14432), .A2(n14431), .ZN(n14437) );
  NAND2_X1 U18099 ( .A1(n14434), .A2(n14433), .ZN(n14449) );
  NOR2_X1 U18100 ( .A1(n14435), .A2(n11896), .ZN(n14447) );
  XNOR2_X1 U18101 ( .A(n12589), .B(n13950), .ZN(n15778) );
  MUX2_X1 U18102 ( .A(n14449), .B(n14447), .S(n15778), .Z(n14436) );
  AOI211_X1 U18103 ( .C1(n15792), .C2(n15935), .A(n14437), .B(n14436), .ZN(
        n15781) );
  INV_X1 U18104 ( .A(n15781), .ZN(n14438) );
  MUX2_X1 U18105 ( .A(n15783), .B(n14438), .S(n15939), .Z(n15944) );
  AOI22_X1 U18106 ( .A1(n14462), .A2(n15783), .B1(n18052), .B2(n15944), .ZN(
        n14455) );
  NAND2_X1 U18107 ( .A1(n15783), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n14440) );
  XNOR2_X1 U18108 ( .A(n15788), .B(n14440), .ZN(n14441) );
  NAND2_X1 U18109 ( .A1(n15937), .A2(n14441), .ZN(n14451) );
  MUX2_X1 U18110 ( .A(n14442), .B(n15788), .S(n13950), .Z(n14444) );
  NOR2_X1 U18111 ( .A1(n14444), .A2(n14443), .ZN(n14448) );
  NAND2_X1 U18112 ( .A1(n13950), .A2(n15783), .ZN(n14445) );
  NAND2_X1 U18113 ( .A1(n14445), .A2(n15788), .ZN(n14446) );
  NAND2_X1 U18114 ( .A1(n9714), .A2(n14446), .ZN(n15784) );
  AOI22_X1 U18115 ( .A1(n14449), .A2(n14448), .B1(n14447), .B2(n15784), .ZN(
        n14450) );
  NAND2_X1 U18116 ( .A1(n14451), .A2(n14450), .ZN(n14452) );
  AOI21_X1 U18117 ( .B1(n14439), .B2(n15935), .A(n14452), .ZN(n15786) );
  NOR2_X1 U18118 ( .A1(n15939), .A2(n15788), .ZN(n14453) );
  AOI21_X1 U18119 ( .B1(n15786), .B2(n15939), .A(n14453), .ZN(n15933) );
  AOI22_X1 U18120 ( .A1(n14462), .A2(n15788), .B1(n15933), .B2(n18052), .ZN(
        n14454) );
  NOR2_X1 U18121 ( .A1(n14455), .A2(n14454), .ZN(n15956) );
  NAND2_X1 U18122 ( .A1(n15956), .A2(n14456), .ZN(n15766) );
  INV_X1 U18123 ( .A(n14457), .ZN(n14472) );
  OR2_X1 U18124 ( .A1(n14365), .A2(n14472), .ZN(n14458) );
  XNOR2_X1 U18125 ( .A(n14458), .B(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n21000) );
  INV_X1 U18126 ( .A(n14459), .ZN(n14460) );
  NAND2_X1 U18127 ( .A1(n21000), .A2(n14460), .ZN(n18044) );
  NAND2_X1 U18128 ( .A1(n18044), .A2(n15939), .ZN(n14461) );
  NAND2_X1 U18129 ( .A1(n14461), .A2(n18052), .ZN(n14465) );
  INV_X1 U18130 ( .A(n14462), .ZN(n14464) );
  AOI21_X1 U18131 ( .B1(n15939), .B2(n18052), .A(
        P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n14463) );
  AOI21_X1 U18132 ( .B1(n14465), .B2(n14464), .A(n14463), .ZN(n15955) );
  INV_X1 U18133 ( .A(n15955), .ZN(n15764) );
  AND3_X1 U18134 ( .A1(n15766), .A2(n20944), .A3(n15764), .ZN(n14466) );
  INV_X1 U18135 ( .A(n21146), .ZN(n14470) );
  NAND2_X1 U18136 ( .A1(n14363), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n21231) );
  XNOR2_X1 U18137 ( .A(n9709), .B(n21231), .ZN(n14467) );
  NAND2_X1 U18138 ( .A1(n21719), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n15769) );
  AOI22_X1 U18139 ( .A1(n14467), .A2(n21376), .B1(n15792), .B2(n15769), .ZN(
        n14469) );
  NAND2_X1 U18140 ( .A1(n14470), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n14468) );
  OAI21_X1 U18141 ( .B1(n14470), .B2(n14469), .A(n14468), .ZN(P1_U3476) );
  OAI222_X1 U18142 ( .A1(n20988), .A2(n15298), .B1(n15246), .B2(n15296), .C1(
        n14816), .C2(n12116), .ZN(P1_U2899) );
  INV_X1 U18143 ( .A(n14362), .ZN(n14471) );
  NOR2_X1 U18144 ( .A1(n21681), .A2(n21269), .ZN(n21301) );
  INV_X1 U18145 ( .A(n21268), .ZN(n21273) );
  NAND2_X1 U18146 ( .A1(n15792), .A2(n14472), .ZN(n21298) );
  INV_X1 U18147 ( .A(n21298), .ZN(n21270) );
  INV_X1 U18148 ( .A(n14500), .ZN(n14473) );
  AOI21_X1 U18149 ( .B1(n21270), .B2(n14526), .A(n14473), .ZN(n14476) );
  OAI211_X1 U18150 ( .C1(n21273), .C2(n21231), .A(n21376), .B(n14476), .ZN(
        n14474) );
  NAND2_X1 U18151 ( .A1(n14499), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n14480) );
  INV_X1 U18152 ( .A(n21508), .ZN(n21444) );
  INV_X1 U18153 ( .A(n14476), .ZN(n14477) );
  AOI22_X1 U18154 ( .A1(n14477), .A2(n21376), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n21301), .ZN(n14501) );
  OAI22_X1 U18155 ( .A1(n14501), .A2(n21406), .B1(n14500), .B2(n21329), .ZN(
        n14478) );
  AOI21_X1 U18156 ( .B1(n21341), .B2(n21444), .A(n14478), .ZN(n14479) );
  OAI211_X1 U18157 ( .C1(n21447), .C2(n14505), .A(n14480), .B(n14479), .ZN(
        P1_U3094) );
  NAND2_X1 U18158 ( .A1(n14499), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n14483) );
  INV_X1 U18159 ( .A(n21486), .ZN(n21429) );
  OAI22_X1 U18160 ( .A1(n14501), .A2(n21397), .B1(n14500), .B2(n21313), .ZN(
        n14481) );
  AOI21_X1 U18161 ( .B1(n21341), .B2(n21429), .A(n14481), .ZN(n14482) );
  OAI211_X1 U18162 ( .C1(n21432), .C2(n14505), .A(n14483), .B(n14482), .ZN(
        P1_U3090) );
  NAND2_X1 U18163 ( .A1(n14499), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n14486) );
  INV_X1 U18164 ( .A(n21502), .ZN(n21440) );
  OAI22_X1 U18165 ( .A1(n14501), .A2(n21403), .B1(n14500), .B2(n21325), .ZN(
        n14484) );
  AOI21_X1 U18166 ( .B1(n21341), .B2(n21440), .A(n14484), .ZN(n14485) );
  OAI211_X1 U18167 ( .C1(n21443), .C2(n14505), .A(n14486), .B(n14485), .ZN(
        P1_U3093) );
  NAND2_X1 U18168 ( .A1(n14499), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n14489) );
  INV_X1 U18169 ( .A(n21496), .ZN(n21436) );
  OAI22_X1 U18170 ( .A1(n14501), .A2(n21400), .B1(n14500), .B2(n21321), .ZN(
        n14487) );
  AOI21_X1 U18171 ( .B1(n21341), .B2(n21436), .A(n14487), .ZN(n14488) );
  OAI211_X1 U18172 ( .C1(n21439), .C2(n14505), .A(n14489), .B(n14488), .ZN(
        P1_U3092) );
  NAND2_X1 U18173 ( .A1(n14499), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n14492) );
  INV_X1 U18174 ( .A(n21490), .ZN(n21929) );
  OAI22_X1 U18175 ( .A1(n14501), .A2(n21936), .B1(n14500), .B2(n21317), .ZN(
        n14490) );
  AOI21_X1 U18176 ( .B1(n21341), .B2(n21929), .A(n14490), .ZN(n14491) );
  OAI211_X1 U18177 ( .C1(n21435), .C2(n14505), .A(n14492), .B(n14491), .ZN(
        P1_U3091) );
  NAND2_X1 U18178 ( .A1(n14499), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n14495) );
  INV_X1 U18179 ( .A(n21514), .ZN(n21448) );
  OAI22_X1 U18180 ( .A1(n14501), .A2(n21409), .B1(n14500), .B2(n21333), .ZN(
        n14493) );
  AOI21_X1 U18181 ( .B1(n21341), .B2(n21448), .A(n14493), .ZN(n14494) );
  OAI211_X1 U18182 ( .C1(n21451), .C2(n14505), .A(n14495), .B(n14494), .ZN(
        P1_U3095) );
  NAND2_X1 U18183 ( .A1(n14499), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n14498) );
  INV_X1 U18184 ( .A(n21525), .ZN(n21454) );
  OAI22_X1 U18185 ( .A1(n14501), .A2(n21412), .B1(n14500), .B2(n21337), .ZN(
        n14496) );
  AOI21_X1 U18186 ( .B1(n21341), .B2(n21454), .A(n14496), .ZN(n14497) );
  OAI211_X1 U18187 ( .C1(n21459), .C2(n14505), .A(n14498), .B(n14497), .ZN(
        P1_U3096) );
  NAND2_X1 U18188 ( .A1(n14499), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n14504) );
  INV_X1 U18189 ( .A(n21480), .ZN(n21425) );
  OAI22_X1 U18190 ( .A1(n14501), .A2(n21394), .B1(n14500), .B2(n21303), .ZN(
        n14502) );
  AOI21_X1 U18191 ( .B1(n21341), .B2(n21425), .A(n14502), .ZN(n14503) );
  OAI211_X1 U18192 ( .C1(n21428), .C2(n14505), .A(n14504), .B(n14503), .ZN(
        P1_U3089) );
  INV_X1 U18193 ( .A(n14506), .ZN(n14507) );
  AOI21_X1 U18194 ( .B1(n14507), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A(
        P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n14508) );
  NOR3_X1 U18195 ( .A1(n16698), .A2(n14508), .A3(n16733), .ZN(n14513) );
  NAND2_X1 U18196 ( .A1(n14340), .A2(n14510), .ZN(n14511) );
  AND2_X1 U18197 ( .A1(n14509), .A2(n14511), .ZN(n17423) );
  MUX2_X1 U18198 ( .A(P2_EBX_REG_6__SCAN_IN), .B(n17423), .S(n16728), .Z(
        n14512) );
  OR2_X1 U18199 ( .A1(n14513), .A2(n14512), .ZN(P2_U2881) );
  NAND2_X1 U18200 ( .A1(n13526), .A2(n14515), .ZN(n14516) );
  NAND2_X1 U18201 ( .A1(n14514), .A2(n14516), .ZN(n17354) );
  AOI22_X1 U18202 ( .A1(n16869), .A2(n16764), .B1(P2_EAX_REG_12__SCAN_IN), 
        .B2(n16867), .ZN(n14517) );
  OAI21_X1 U18203 ( .B1(n17354), .B2(n16864), .A(n14517), .ZN(P2_U2907) );
  XNOR2_X1 U18204 ( .A(n16698), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n14523) );
  NAND2_X1 U18205 ( .A1(n14509), .A2(n14519), .ZN(n14520) );
  AND2_X1 U18206 ( .A1(n14518), .A2(n14520), .ZN(n18080) );
  NAND2_X1 U18207 ( .A1(n18080), .A2(n16728), .ZN(n14522) );
  NAND2_X1 U18208 ( .A1(n16723), .A2(P2_EBX_REG_7__SCAN_IN), .ZN(n14521) );
  OAI211_X1 U18209 ( .C1(n14523), .C2(n16733), .A(n14522), .B(n14521), .ZN(
        P2_U2880) );
  NAND2_X1 U18210 ( .A1(n15945), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n21346) );
  NOR2_X1 U18211 ( .A1(n21681), .A2(n21346), .ZN(n21384) );
  INV_X1 U18212 ( .A(n15792), .ZN(n21022) );
  NAND2_X1 U18213 ( .A1(n14439), .A2(n21022), .ZN(n21379) );
  INV_X1 U18214 ( .A(n21379), .ZN(n21348) );
  NOR2_X1 U18215 ( .A1(n14525), .A2(n21346), .ZN(n14530) );
  AOI21_X1 U18216 ( .B1(n21348), .B2(n14526), .A(n14530), .ZN(n14528) );
  OAI211_X1 U18217 ( .C1(n21355), .C2(n21231), .A(n21376), .B(n14528), .ZN(
        n14527) );
  NAND2_X1 U18218 ( .A1(n14552), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n14533) );
  NAND2_X1 U18219 ( .A1(n15848), .A2(n15812), .ZN(n15896) );
  INV_X1 U18220 ( .A(n14528), .ZN(n14529) );
  AOI22_X1 U18221 ( .A1(n14529), .A2(n21376), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n21384), .ZN(n14554) );
  INV_X1 U18222 ( .A(n14530), .ZN(n14553) );
  OAI22_X1 U18223 ( .A1(n14554), .A2(n21406), .B1(n21329), .B2(n14553), .ZN(
        n14531) );
  AOI21_X1 U18224 ( .B1(n15930), .B2(n21505), .A(n14531), .ZN(n14532) );
  OAI211_X1 U18225 ( .C1(n21508), .C2(n21391), .A(n14533), .B(n14532), .ZN(
        P1_U3126) );
  NAND2_X1 U18226 ( .A1(n14552), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n14536) );
  OAI22_X1 U18227 ( .A1(n14554), .A2(n21394), .B1(n21303), .B2(n14553), .ZN(
        n14534) );
  AOI21_X1 U18228 ( .B1(n15930), .B2(n21477), .A(n14534), .ZN(n14535) );
  OAI211_X1 U18229 ( .C1(n21480), .C2(n21391), .A(n14536), .B(n14535), .ZN(
        P1_U3121) );
  NAND2_X1 U18230 ( .A1(n14552), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n14539) );
  OAI22_X1 U18231 ( .A1(n14554), .A2(n21403), .B1(n21325), .B2(n14553), .ZN(
        n14537) );
  AOI21_X1 U18232 ( .B1(n15930), .B2(n21499), .A(n14537), .ZN(n14538) );
  OAI211_X1 U18233 ( .C1(n21502), .C2(n21391), .A(n14539), .B(n14538), .ZN(
        P1_U3125) );
  NAND2_X1 U18234 ( .A1(n14552), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n14542) );
  OAI22_X1 U18235 ( .A1(n14554), .A2(n21409), .B1(n21333), .B2(n14553), .ZN(
        n14540) );
  AOI21_X1 U18236 ( .B1(n15930), .B2(n21511), .A(n14540), .ZN(n14541) );
  OAI211_X1 U18237 ( .C1(n21514), .C2(n21391), .A(n14542), .B(n14541), .ZN(
        P1_U3127) );
  NAND2_X1 U18238 ( .A1(n14552), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n14545) );
  OAI22_X1 U18239 ( .A1(n14554), .A2(n21400), .B1(n21321), .B2(n14553), .ZN(
        n14543) );
  AOI21_X1 U18240 ( .B1(n15930), .B2(n21493), .A(n14543), .ZN(n14544) );
  OAI211_X1 U18241 ( .C1(n21496), .C2(n21391), .A(n14545), .B(n14544), .ZN(
        P1_U3124) );
  NAND2_X1 U18242 ( .A1(n14552), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n14548) );
  OAI22_X1 U18243 ( .A1(n14554), .A2(n21397), .B1(n21313), .B2(n14553), .ZN(
        n14546) );
  AOI21_X1 U18244 ( .B1(n15930), .B2(n21483), .A(n14546), .ZN(n14547) );
  OAI211_X1 U18245 ( .C1(n21486), .C2(n21391), .A(n14548), .B(n14547), .ZN(
        P1_U3122) );
  NAND2_X1 U18246 ( .A1(n14552), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n14551) );
  OAI22_X1 U18247 ( .A1(n14554), .A2(n21412), .B1(n21337), .B2(n14553), .ZN(
        n14549) );
  AOI21_X1 U18248 ( .B1(n15930), .B2(n21519), .A(n14549), .ZN(n14550) );
  OAI211_X1 U18249 ( .C1(n21525), .C2(n21391), .A(n14551), .B(n14550), .ZN(
        P1_U3128) );
  NAND2_X1 U18250 ( .A1(n14552), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n14557) );
  OAI22_X1 U18251 ( .A1(n14554), .A2(n21936), .B1(n21317), .B2(n14553), .ZN(
        n14555) );
  AOI21_X1 U18252 ( .B1(n15930), .B2(n21931), .A(n14555), .ZN(n14556) );
  OAI211_X1 U18253 ( .C1(n21490), .C2(n21391), .A(n14557), .B(n14556), .ZN(
        P1_U3123) );
  INV_X1 U18254 ( .A(n14558), .ZN(n14559) );
  NOR2_X1 U18255 ( .A1(n14560), .A2(n14559), .ZN(n14566) );
  NAND2_X1 U18256 ( .A1(n14563), .A2(n14562), .ZN(n14564) );
  NAND2_X1 U18257 ( .A1(n14561), .A2(n14564), .ZN(n18090) );
  XNOR2_X1 U18258 ( .A(n20535), .B(n18090), .ZN(n14565) );
  NOR2_X1 U18259 ( .A1(n14566), .A2(n14565), .ZN(n16857) );
  AOI21_X1 U18260 ( .B1(n14566), .B2(n14565), .A(n16857), .ZN(n14569) );
  INV_X1 U18261 ( .A(n18090), .ZN(n20889) );
  AOI22_X1 U18262 ( .A1(n20889), .A2(n16868), .B1(P2_EAX_REG_3__SCAN_IN), .B2(
        n16867), .ZN(n14568) );
  NAND2_X1 U18263 ( .A1(n16869), .A2(n17569), .ZN(n14567) );
  OAI211_X1 U18264 ( .C1(n14569), .C2(n16872), .A(n14568), .B(n14567), .ZN(
        P2_U2916) );
  OR2_X1 U18265 ( .A1(n14428), .A2(n14572), .ZN(n14573) );
  AND2_X1 U18266 ( .A1(n14571), .A2(n14573), .ZN(n20983) );
  INV_X1 U18267 ( .A(n20983), .ZN(n14693) );
  OAI21_X1 U18268 ( .B1(n14576), .B2(n14575), .A(n14574), .ZN(n14577) );
  AND2_X1 U18269 ( .A1(n14577), .A2(n15132), .ZN(n20976) );
  AOI22_X1 U18270 ( .A1(n20976), .A2(n15196), .B1(P1_EBX_REG_6__SCAN_IN), .B2(
        n15195), .ZN(n14578) );
  OAI21_X1 U18271 ( .B1(n14693), .B2(n15206), .A(n14578), .ZN(P1_U2866) );
  NAND2_X1 U18272 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .ZN(n18626) );
  INV_X1 U18273 ( .A(n18626), .ZN(n14581) );
  NAND2_X1 U18274 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n14579), .ZN(n18677) );
  NAND2_X1 U18275 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n18656), .ZN(n18650) );
  NAND2_X1 U18276 ( .A1(P3_EBX_REG_25__SCAN_IN), .A2(n18649), .ZN(n18633) );
  NAND2_X1 U18277 ( .A1(n18777), .A2(n18638), .ZN(n14580) );
  OAI21_X1 U18278 ( .B1(n14581), .B2(n18780), .A(n14580), .ZN(n18628) );
  INV_X1 U18279 ( .A(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n14588) );
  INV_X1 U18280 ( .A(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n14582) );
  INV_X1 U18281 ( .A(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n21818) );
  OAI22_X1 U18282 ( .A1(n18724), .A2(n14582), .B1(n18722), .B2(n21818), .ZN(
        n14585) );
  INV_X1 U18283 ( .A(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n14583) );
  OAI22_X1 U18284 ( .A1(n18728), .A2(n14583), .B1(n18726), .B2(n17708), .ZN(
        n14584) );
  AOI211_X1 U18285 ( .C1(n18731), .C2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A(
        n14585), .B(n14584), .ZN(n14587) );
  AOI22_X1 U18286 ( .A1(n9704), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n18732), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n14586) );
  OAI211_X1 U18287 ( .C1(n18735), .C2(n14588), .A(n14587), .B(n14586), .ZN(
        n14600) );
  AOI22_X1 U18288 ( .A1(n13279), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n18596), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n14590) );
  AOI22_X1 U18289 ( .A1(n18740), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n18739), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n14589) );
  NAND2_X1 U18290 ( .A1(n14590), .A2(n14589), .ZN(n14599) );
  INV_X1 U18291 ( .A(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n14592) );
  INV_X1 U18292 ( .A(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n17709) );
  OAI22_X1 U18293 ( .A1(n14593), .A2(n14592), .B1(n14591), .B2(n17709), .ZN(
        n14598) );
  INV_X1 U18294 ( .A(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n21805) );
  OAI22_X1 U18295 ( .A1(n14596), .A2(n14595), .B1(n14594), .B2(n21805), .ZN(
        n14597) );
  NOR4_X1 U18296 ( .A1(n14600), .A2(n14599), .A3(n14598), .A4(n14597), .ZN(
        n14688) );
  INV_X1 U18297 ( .A(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n14609) );
  OAI22_X1 U18298 ( .A1(n14601), .A2(n18724), .B1(n18722), .B2(n19604), .ZN(
        n14606) );
  INV_X1 U18299 ( .A(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n14604) );
  INV_X1 U18300 ( .A(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n14602) );
  OAI22_X1 U18301 ( .A1(n18728), .A2(n14604), .B1(n14603), .B2(n14602), .ZN(
        n14605) );
  AOI211_X1 U18302 ( .C1(n18731), .C2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A(
        n14606), .B(n14605), .ZN(n14608) );
  AOI22_X1 U18303 ( .A1(n18736), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n18732), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n14607) );
  OAI211_X1 U18304 ( .C1(n18735), .C2(n14609), .A(n14608), .B(n14607), .ZN(
        n14615) );
  AOI22_X1 U18305 ( .A1(n18703), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n14680), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n14613) );
  AOI22_X1 U18306 ( .A1(n18738), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n14679), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n14612) );
  AOI22_X1 U18307 ( .A1(n18740), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n9703), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n14611) );
  AOI22_X1 U18308 ( .A1(n13279), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n18596), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n14610) );
  NAND4_X1 U18309 ( .A1(n14613), .A2(n14612), .A3(n14611), .A4(n14610), .ZN(
        n14614) );
  NOR2_X1 U18310 ( .A1(n14615), .A2(n14614), .ZN(n18636) );
  NAND2_X1 U18311 ( .A1(n9704), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n14617) );
  NAND2_X1 U18312 ( .A1(n18699), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n14616) );
  OAI211_X1 U18313 ( .C1(n18735), .C2(n19621), .A(n14617), .B(n14616), .ZN(
        n14618) );
  INV_X1 U18314 ( .A(n14618), .ZN(n14622) );
  AOI22_X1 U18315 ( .A1(n18704), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n18703), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n14621) );
  AOI22_X1 U18316 ( .A1(n18706), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n18705), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n14620) );
  NAND2_X1 U18317 ( .A1(n18731), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n14619) );
  NAND4_X1 U18318 ( .A1(n14622), .A2(n14621), .A3(n14620), .A4(n14619), .ZN(
        n14628) );
  AOI22_X1 U18319 ( .A1(n18736), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n14679), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n14626) );
  AOI22_X1 U18320 ( .A1(n13279), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n18596), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n14625) );
  AOI22_X1 U18321 ( .A1(n18740), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n18739), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n14624) );
  AOI22_X1 U18322 ( .A1(n18738), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n18737), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n14623) );
  NAND4_X1 U18323 ( .A1(n14626), .A2(n14625), .A3(n14624), .A4(n14623), .ZN(
        n14627) );
  OR2_X1 U18324 ( .A1(n14628), .A2(n14627), .ZN(n18652) );
  INV_X1 U18325 ( .A(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n18603) );
  NAND2_X1 U18326 ( .A1(n9704), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n14630) );
  NAND2_X1 U18327 ( .A1(n18699), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n14629) );
  OAI211_X1 U18328 ( .C1(n18735), .C2(n18603), .A(n14630), .B(n14629), .ZN(
        n14631) );
  INV_X1 U18329 ( .A(n14631), .ZN(n14635) );
  AOI22_X1 U18330 ( .A1(n18704), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n9683), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n14634) );
  AOI22_X1 U18331 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18706), .B1(
        n18705), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n14633) );
  NAND2_X1 U18332 ( .A1(n18731), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n14632) );
  NAND4_X1 U18333 ( .A1(n14635), .A2(n14634), .A3(n14633), .A4(n14632), .ZN(
        n14641) );
  AOI22_X1 U18334 ( .A1(n18736), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n14679), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n14639) );
  AOI22_X1 U18335 ( .A1(n13279), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n18596), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n14638) );
  AOI22_X1 U18336 ( .A1(n18740), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n18739), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n14637) );
  AOI22_X1 U18337 ( .A1(n18738), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n18737), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n14636) );
  NAND4_X1 U18338 ( .A1(n14639), .A2(n14638), .A3(n14637), .A4(n14636), .ZN(
        n14640) );
  OR2_X1 U18339 ( .A1(n14641), .A2(n14640), .ZN(n18653) );
  NAND2_X1 U18340 ( .A1(n18652), .A2(n18653), .ZN(n18651) );
  NAND2_X1 U18341 ( .A1(n9703), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n14643) );
  NAND2_X1 U18342 ( .A1(n18699), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n14642) );
  OAI211_X1 U18343 ( .C1(n18735), .C2(n19624), .A(n14643), .B(n14642), .ZN(
        n14644) );
  INV_X1 U18344 ( .A(n14644), .ZN(n14648) );
  AOI22_X1 U18345 ( .A1(n18704), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n18736), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n14647) );
  AOI22_X1 U18346 ( .A1(n18706), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n18705), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n14646) );
  NAND2_X1 U18347 ( .A1(n18731), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n14645) );
  NAND4_X1 U18348 ( .A1(n14648), .A2(n14647), .A3(n14646), .A4(n14645), .ZN(
        n14655) );
  AOI22_X1 U18349 ( .A1(n18738), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n14679), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n14653) );
  AOI22_X1 U18350 ( .A1(n9683), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n14649), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n14652) );
  AOI22_X1 U18351 ( .A1(n13279), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n18596), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n14651) );
  AOI22_X1 U18352 ( .A1(n18737), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n18739), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n14650) );
  NAND4_X1 U18353 ( .A1(n14653), .A2(n14652), .A3(n14651), .A4(n14650), .ZN(
        n14654) );
  NOR2_X1 U18354 ( .A1(n14655), .A2(n14654), .ZN(n18644) );
  NOR2_X1 U18355 ( .A1(n18651), .A2(n18644), .ZN(n18646) );
  INV_X1 U18356 ( .A(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n14658) );
  NAND2_X1 U18357 ( .A1(n9704), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n14657) );
  NAND2_X1 U18358 ( .A1(n18699), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n14656) );
  OAI211_X1 U18359 ( .C1(n18735), .C2(n14658), .A(n14657), .B(n14656), .ZN(
        n14659) );
  INV_X1 U18360 ( .A(n14659), .ZN(n14663) );
  AOI22_X1 U18361 ( .A1(n18704), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n9683), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n14662) );
  AOI22_X1 U18362 ( .A1(n18706), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n18705), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n14661) );
  NAND2_X1 U18363 ( .A1(n18731), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n14660) );
  NAND4_X1 U18364 ( .A1(n14663), .A2(n14662), .A3(n14661), .A4(n14660), .ZN(
        n14669) );
  AOI22_X1 U18365 ( .A1(n18736), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n13878), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n14667) );
  AOI22_X1 U18366 ( .A1(n13279), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n18596), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n14666) );
  AOI22_X1 U18367 ( .A1(n18740), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n18739), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n14665) );
  AOI22_X1 U18368 ( .A1(n18738), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n18737), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n14664) );
  NAND4_X1 U18369 ( .A1(n14667), .A2(n14666), .A3(n14665), .A4(n14664), .ZN(
        n14668) );
  OR2_X1 U18370 ( .A1(n14669), .A2(n14668), .ZN(n18641) );
  NAND2_X1 U18371 ( .A1(n18646), .A2(n18641), .ZN(n18640) );
  NOR2_X1 U18372 ( .A1(n18636), .A2(n18640), .ZN(n18635) );
  INV_X1 U18373 ( .A(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n14678) );
  OAI22_X1 U18374 ( .A1(n14671), .A2(n18724), .B1(n18722), .B2(n14670), .ZN(
        n14675) );
  INV_X1 U18375 ( .A(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n14673) );
  OAI22_X1 U18376 ( .A1(n18728), .A2(n14673), .B1(n18726), .B2(n14672), .ZN(
        n14674) );
  AOI211_X1 U18377 ( .C1(n18731), .C2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A(
        n14675), .B(n14674), .ZN(n14677) );
  AOI22_X1 U18378 ( .A1(n9703), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n18732), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n14676) );
  OAI211_X1 U18379 ( .C1(n18735), .C2(n14678), .A(n14677), .B(n14676), .ZN(
        n14686) );
  AOI22_X1 U18380 ( .A1(n18736), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n14679), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n14684) );
  AOI22_X1 U18381 ( .A1(n18738), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n14680), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n14683) );
  AOI22_X1 U18382 ( .A1(n13279), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n18596), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n14682) );
  AOI22_X1 U18383 ( .A1(n18740), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n18739), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n14681) );
  NAND4_X1 U18384 ( .A1(n14684), .A2(n14683), .A3(n14682), .A4(n14681), .ZN(
        n14685) );
  OR2_X1 U18385 ( .A1(n14686), .A2(n14685), .ZN(n18631) );
  NAND2_X1 U18386 ( .A1(n18635), .A2(n18631), .ZN(n18630) );
  OR2_X1 U18387 ( .A1(n18630), .A2(n14688), .ZN(n18625) );
  INV_X1 U18388 ( .A(n18625), .ZN(n14687) );
  AOI21_X1 U18389 ( .B1(n14688), .B2(n18630), .A(n14687), .ZN(n18802) );
  AOI22_X1 U18390 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n18628), .B1(n18802), 
        .B2(n18749), .ZN(n14692) );
  INV_X1 U18391 ( .A(P3_EBX_REG_28__SCAN_IN), .ZN(n14690) );
  INV_X1 U18392 ( .A(n18638), .ZN(n14689) );
  NAND3_X1 U18393 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n14690), .A3(n14689), 
        .ZN(n14691) );
  NAND2_X1 U18394 ( .A1(n14692), .A2(n14691), .ZN(P3_U2675) );
  OAI222_X1 U18395 ( .A1(n14693), .A2(n15298), .B1(n15242), .B2(n15296), .C1(
        n21045), .C2(n14816), .ZN(P1_U2898) );
  INV_X1 U18396 ( .A(n19164), .ZN(n19154) );
  INV_X1 U18397 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n14694) );
  AND2_X1 U18398 ( .A1(n19423), .A2(n19184), .ZN(n19130) );
  AOI22_X1 U18399 ( .A1(n19154), .A2(n14694), .B1(n19139), .B2(n19130), .ZN(
        n14695) );
  NOR2_X1 U18400 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n19165), .ZN(
        n19409) );
  NOR2_X1 U18401 ( .A1(n14695), .A2(n19409), .ZN(n14696) );
  XNOR2_X1 U18402 ( .A(n14696), .B(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n17828) );
  NOR2_X1 U18403 ( .A1(n20016), .A2(n18887), .ZN(n17964) );
  NAND2_X1 U18404 ( .A1(n19546), .A2(n17964), .ZN(n19324) );
  INV_X1 U18405 ( .A(n19324), .ZN(n17954) );
  INV_X1 U18406 ( .A(n19423), .ZN(n19185) );
  INV_X1 U18407 ( .A(n19139), .ZN(n19414) );
  NOR2_X1 U18408 ( .A1(n19185), .A2(n19414), .ZN(n19402) );
  AOI21_X1 U18409 ( .B1(n19402), .B2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n14697) );
  AND2_X1 U18410 ( .A1(n19423), .A2(n19387), .ZN(n19134) );
  NOR2_X1 U18411 ( .A1(n14697), .A2(n19134), .ZN(n17826) );
  INV_X1 U18412 ( .A(n19426), .ZN(n14698) );
  OR2_X1 U18413 ( .A1(n14708), .A2(n14698), .ZN(n14699) );
  NOR3_X1 U18414 ( .A1(n14698), .A2(n14707), .A3(n14708), .ZN(n19124) );
  AOI21_X1 U18415 ( .B1(n14707), .B2(n14699), .A(n19124), .ZN(n14700) );
  INV_X1 U18416 ( .A(n14700), .ZN(n17824) );
  NOR2_X1 U18417 ( .A1(n19442), .A2(n20093), .ZN(n14701) );
  AOI21_X1 U18418 ( .B1(n19527), .B2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n14701), .ZN(n14711) );
  INV_X1 U18419 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n19533) );
  OAI21_X1 U18420 ( .B1(n19533), .B2(n17962), .A(n19550), .ZN(n19462) );
  NOR2_X1 U18421 ( .A1(n19550), .A2(n19533), .ZN(n19464) );
  INV_X1 U18422 ( .A(n19532), .ZN(n19465) );
  AOI21_X1 U18423 ( .B1(n19314), .B2(n17962), .A(n19465), .ZN(n19539) );
  AOI22_X1 U18424 ( .A1(n20023), .A2(n19462), .B1(n19464), .B2(n19539), .ZN(
        n19523) );
  INV_X1 U18425 ( .A(n19523), .ZN(n14702) );
  INV_X1 U18426 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n19496) );
  NAND3_X1 U18427 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n19466) );
  NOR3_X1 U18428 ( .A1(n19496), .A2(n19485), .A3(n19466), .ZN(n14703) );
  NAND2_X1 U18429 ( .A1(n14702), .A2(n14703), .ZN(n19471) );
  OR2_X1 U18430 ( .A1(n13316), .A2(n19471), .ZN(n17955) );
  NAND3_X1 U18431 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n14703), .A3(
        n19462), .ZN(n19401) );
  NAND2_X1 U18432 ( .A1(n14703), .A2(n19464), .ZN(n19453) );
  NOR2_X1 U18433 ( .A1(n13316), .A2(n19453), .ZN(n17855) );
  NOR2_X1 U18434 ( .A1(n19314), .A2(n17855), .ZN(n19440) );
  AOI21_X1 U18435 ( .B1(n20023), .B2(n19401), .A(n19440), .ZN(n19379) );
  NAND2_X1 U18436 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n17855), .ZN(
        n19429) );
  INV_X1 U18437 ( .A(n19429), .ZN(n19450) );
  INV_X1 U18438 ( .A(n19428), .ZN(n19451) );
  AOI21_X1 U18439 ( .B1(n19139), .B2(n19450), .A(n19451), .ZN(n19407) );
  AOI211_X1 U18440 ( .C1(n20023), .C2(n19414), .A(n19407), .B(n14707), .ZN(
        n14704) );
  OAI211_X1 U18441 ( .C1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .C2(n19355), .A(
        n19379), .B(n14704), .ZN(n14705) );
  OAI221_X1 U18442 ( .B1(n14705), .B2(n14708), .C1(n14705), .C2(n19454), .A(
        n19546), .ZN(n14706) );
  AOI221_X1 U18443 ( .B1(n14708), .B2(n14707), .C1(n17955), .C2(n14707), .A(
        n14706), .ZN(n14709) );
  INV_X1 U18444 ( .A(n14709), .ZN(n14710) );
  OAI211_X1 U18445 ( .C1(n17824), .C2(n19530), .A(n14711), .B(n14710), .ZN(
        n14712) );
  AOI21_X1 U18446 ( .B1(n17954), .B2(n17826), .A(n14712), .ZN(n14713) );
  OAI21_X1 U18447 ( .B1(n19364), .B2(n17828), .A(n14713), .ZN(P3_U2848) );
  INV_X1 U18448 ( .A(n14744), .ZN(n20037) );
  INV_X1 U18449 ( .A(n14748), .ZN(n17982) );
  NOR2_X1 U18450 ( .A1(n19428), .A2(n14714), .ZN(n14722) );
  NAND2_X1 U18451 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n17962), .ZN(n14715) );
  OAI211_X1 U18452 ( .C1(n20001), .C2(n18577), .A(n17982), .B(n14715), .ZN(
        n14716) );
  OAI21_X1 U18453 ( .B1(n17982), .B2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n14716), .ZN(n14717) );
  OAI21_X1 U18454 ( .B1(n14748), .B2(n14718), .A(n14717), .ZN(P3_U3290) );
  INV_X1 U18455 ( .A(n14719), .ZN(n14721) );
  INV_X1 U18456 ( .A(n14720), .ZN(n14735) );
  NAND2_X1 U18457 ( .A1(n14721), .A2(n14735), .ZN(n18563) );
  OR2_X1 U18458 ( .A1(n14722), .A2(n18563), .ZN(n14724) );
  NAND2_X1 U18459 ( .A1(n14734), .A2(n14728), .ZN(n14723) );
  NAND2_X1 U18460 ( .A1(n14724), .A2(n14723), .ZN(n20003) );
  NOR2_X1 U18461 ( .A1(n20049), .A2(n17962), .ZN(n14742) );
  INV_X1 U18462 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n17871) );
  OAI22_X1 U18463 ( .A1(n17871), .A2(n19533), .B1(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14740) );
  NAND2_X1 U18464 ( .A1(n14742), .A2(n14740), .ZN(n14725) );
  OAI211_X1 U18465 ( .C1(n18563), .C2(n14744), .A(n17982), .B(n14725), .ZN(
        n14726) );
  AOI21_X1 U18466 ( .B1(n20003), .B2(n17979), .A(n14726), .ZN(n14727) );
  AOI21_X1 U18467 ( .B1(n14748), .B2(n14728), .A(n14727), .ZN(P3_U3289) );
  AND2_X1 U18468 ( .A1(n14730), .A2(n14729), .ZN(n14739) );
  INV_X1 U18469 ( .A(n20023), .ZN(n19536) );
  INV_X1 U18470 ( .A(n14731), .ZN(n14733) );
  NAND3_X1 U18471 ( .A1(n14734), .A2(n14733), .A3(n14732), .ZN(n14738) );
  NAND3_X1 U18472 ( .A1(n14736), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        n14735), .ZN(n14737) );
  OAI211_X1 U18473 ( .C1(n14739), .C2(n19536), .A(n14738), .B(n14737), .ZN(
        n20000) );
  INV_X1 U18474 ( .A(n14739), .ZN(n18554) );
  INV_X1 U18475 ( .A(n14740), .ZN(n14741) );
  NAND2_X1 U18476 ( .A1(n14742), .A2(n14741), .ZN(n14743) );
  OAI211_X1 U18477 ( .C1(n18554), .C2(n14744), .A(n17982), .B(n14743), .ZN(
        n14745) );
  AOI21_X1 U18478 ( .B1(n20000), .B2(n17979), .A(n14745), .ZN(n14746) );
  AOI21_X1 U18479 ( .B1(n14748), .B2(n14747), .A(n14746), .ZN(P3_U3288) );
  OR2_X1 U18480 ( .A1(n14751), .A2(n14752), .ZN(n14753) );
  NAND2_X1 U18481 ( .A1(n14750), .A2(n14753), .ZN(n17335) );
  AOI22_X1 U18482 ( .A1(n16869), .A2(n16745), .B1(P2_EAX_REG_14__SCAN_IN), 
        .B2(n16867), .ZN(n14754) );
  OAI21_X1 U18483 ( .B1(n17335), .B2(n16864), .A(n14754), .ZN(P2_U2905) );
  INV_X1 U18484 ( .A(n16757), .ZN(n14758) );
  AND2_X1 U18485 ( .A1(n14514), .A2(n14755), .ZN(n14756) );
  NOR2_X1 U18486 ( .A1(n14751), .A2(n14756), .ZN(n17346) );
  INV_X1 U18487 ( .A(n17346), .ZN(n14757) );
  INV_X1 U18488 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n20219) );
  OAI222_X1 U18489 ( .A1(n14763), .A2(n14758), .B1(n14757), .B2(n16864), .C1(
        n20219), .C2(n16744), .ZN(P2_U2906) );
  AOI21_X1 U18490 ( .B1(n14760), .B2(n14750), .A(n14759), .ZN(n17320) );
  INV_X1 U18491 ( .A(n17320), .ZN(n14761) );
  OAI222_X1 U18492 ( .A1(n14763), .A2(n14762), .B1(n14761), .B2(n16864), .C1(
        n13629), .C2(n16744), .ZN(P2_U2904) );
  NOR2_X1 U18493 ( .A1(n14764), .A2(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n17977) );
  NAND2_X1 U18494 ( .A1(n17977), .A2(n18722), .ZN(n19554) );
  NOR2_X1 U18495 ( .A1(n19554), .A2(P3_FLUSH_REG_SCAN_IN), .ZN(n14765) );
  OAI21_X1 U18496 ( .B1(n14765), .B2(n20133), .A(n19592), .ZN(n19559) );
  INV_X1 U18497 ( .A(n19559), .ZN(n14766) );
  NOR2_X1 U18498 ( .A1(n19239), .A2(n20158), .ZN(n17974) );
  AOI21_X1 U18499 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n17974), .ZN(n17975) );
  NOR2_X1 U18500 ( .A1(n14766), .A2(n17975), .ZN(n14768) );
  INV_X1 U18501 ( .A(n19905), .ZN(n19642) );
  NOR2_X1 U18502 ( .A1(n20134), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19593) );
  OR2_X1 U18503 ( .A1(n19593), .A2(n14766), .ZN(n17973) );
  OR2_X1 U18504 ( .A1(n19642), .A2(n17973), .ZN(n14767) );
  MUX2_X1 U18505 ( .A(n14768), .B(n14767), .S(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .Z(P3_U2864) );
  INV_X1 U18506 ( .A(n14770), .ZN(n16685) );
  NAND3_X1 U18507 ( .A1(n17326), .A2(n14771), .A3(n17325), .ZN(n14772) );
  NAND2_X1 U18508 ( .A1(n14772), .A2(n20257), .ZN(n17316) );
  OAI21_X1 U18509 ( .B1(n17419), .B2(n14773), .A(n17316), .ZN(n17277) );
  AOI21_X1 U18510 ( .B1(n14775), .B2(n14774), .A(n17277), .ZN(n17260) );
  INV_X1 U18511 ( .A(n17260), .ZN(n14778) );
  OAI21_X1 U18512 ( .B1(n17263), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n14776), .ZN(n14777) );
  AOI21_X1 U18513 ( .B1(n14778), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n14777), .ZN(n14779) );
  OAI21_X1 U18514 ( .B1(n16685), .B2(n20259), .A(n14779), .ZN(n14780) );
  INV_X1 U18515 ( .A(n14780), .ZN(n14785) );
  AOI21_X1 U18516 ( .B1(n14782), .B2(n14781), .A(n9755), .ZN(n16827) );
  INV_X1 U18517 ( .A(n16827), .ZN(n14783) );
  OR2_X1 U18518 ( .A1(n14783), .A2(n18091), .ZN(n14784) );
  OAI21_X1 U18519 ( .B1(n14788), .B2(n17443), .A(n14787), .ZN(P2_U3027) );
  OAI21_X1 U18520 ( .B1(n15504), .B2(n14790), .A(n14789), .ZN(n14791) );
  AOI21_X1 U18521 ( .B1(n14792), .B2(n15507), .A(n14791), .ZN(n14795) );
  OAI211_X1 U18522 ( .C1(n14806), .C2(n15511), .A(n14795), .B(n14794), .ZN(
        P1_U2969) );
  INV_X1 U18523 ( .A(DATAI_14_), .ZN(n14798) );
  INV_X1 U18524 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n14797) );
  MUX2_X1 U18525 ( .A(n14798), .B(n14797), .S(n15223), .Z(n21069) );
  OAI22_X1 U18526 ( .A1(n15272), .A2(n21069), .B1(n14799), .B2(n14816), .ZN(
        n14800) );
  AOI21_X1 U18527 ( .B1(BUF1_REG_30__SCAN_IN), .B2(n15274), .A(n14800), .ZN(
        n14804) );
  NAND2_X1 U18528 ( .A1(n15275), .A2(DATAI_30_), .ZN(n14803) );
  OAI211_X1 U18529 ( .C1(n14806), .C2(n15298), .A(n14804), .B(n14803), .ZN(
        P1_U2874) );
  OAI222_X1 U18530 ( .A1(n15203), .A2(n14807), .B1(n15206), .B2(n14806), .C1(
        n14805), .C2(n15204), .ZN(P1_U2842) );
  NAND2_X1 U18531 ( .A1(n15303), .A2(n14808), .ZN(n14810) );
  NAND4_X1 U18532 ( .A1(n15302), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A4(n10056), .ZN(n14809) );
  NAND2_X1 U18533 ( .A1(n15496), .A2(P1_REIP_REG_31__SCAN_IN), .ZN(n15517) );
  NAND2_X1 U18534 ( .A1(n21088), .A2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14811) );
  OAI211_X1 U18535 ( .C1(n14812), .C2(n21098), .A(n15517), .B(n14811), .ZN(
        n14813) );
  AOI21_X1 U18536 ( .B1(n14818), .B2(n21094), .A(n14813), .ZN(n14814) );
  OAI21_X1 U18537 ( .B1(n15519), .B2(n20943), .A(n14814), .ZN(P1_U2968) );
  AOI22_X1 U18538 ( .A1(n15275), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n15286), .ZN(n14819) );
  OAI211_X1 U18539 ( .C1(n15258), .C2(n18100), .A(n14820), .B(n14819), .ZN(
        P1_U2873) );
  INV_X1 U18540 ( .A(n20940), .ZN(n14962) );
  OR2_X1 U18541 ( .A1(P1_READREQUEST_REG_SCAN_IN), .A2(n14962), .ZN(n14824) );
  NAND2_X1 U18542 ( .A1(n14822), .A2(n14821), .ZN(n14823) );
  MUX2_X1 U18543 ( .A(n14824), .B(n14823), .S(n21611), .Z(P1_U3487) );
  OAI21_X1 U18544 ( .B1(n14844), .B2(n14829), .A(n14828), .ZN(n15527) );
  INV_X1 U18545 ( .A(n15527), .ZN(n14836) );
  NOR2_X1 U18546 ( .A1(n21015), .A2(n15300), .ZN(n14835) );
  AOI22_X1 U18547 ( .A1(n21024), .A2(P1_EBX_REG_29__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n21019), .ZN(n14832) );
  INV_X1 U18548 ( .A(n14842), .ZN(n14830) );
  NAND2_X1 U18549 ( .A1(n14830), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n14831) );
  OAI211_X1 U18550 ( .C1(n14833), .C2(P1_REIP_REG_29__SCAN_IN), .A(n14832), 
        .B(n14831), .ZN(n14834) );
  AOI211_X1 U18551 ( .C1(n14836), .C2(n20992), .A(n14835), .B(n14834), .ZN(
        n14837) );
  OAI21_X1 U18552 ( .B1(n15306), .B2(n15112), .A(n14837), .ZN(P1_U2811) );
  AOI21_X1 U18553 ( .B1(n14838), .B2(n13151), .A(n14825), .ZN(n15315) );
  INV_X1 U18554 ( .A(n15315), .ZN(n15216) );
  INV_X1 U18555 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n14841) );
  NAND3_X1 U18556 ( .A1(n14858), .A2(P1_REIP_REG_27__SCAN_IN), .A3(n14841), 
        .ZN(n14840) );
  AOI22_X1 U18557 ( .A1(n21024), .A2(P1_EBX_REG_28__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n21019), .ZN(n14839) );
  OAI211_X1 U18558 ( .C1(n14842), .C2(n14841), .A(n14840), .B(n14839), .ZN(
        n14847) );
  INV_X1 U18559 ( .A(n14862), .ZN(n14850) );
  AOI21_X1 U18560 ( .B1(n14850), .B2(n14849), .A(n14843), .ZN(n14845) );
  OR2_X1 U18561 ( .A1(n14845), .A2(n14844), .ZN(n15534) );
  NOR2_X1 U18562 ( .A1(n15534), .A2(n21026), .ZN(n14846) );
  AOI211_X1 U18563 ( .C1(n21027), .C2(n15312), .A(n14847), .B(n14846), .ZN(
        n14848) );
  OAI21_X1 U18564 ( .B1(n15216), .B2(n15112), .A(n14848), .ZN(P1_U2812) );
  XNOR2_X1 U18565 ( .A(n14850), .B(n14849), .ZN(n15541) );
  NAND2_X1 U18566 ( .A1(n14851), .A2(n20982), .ZN(n14860) );
  INV_X1 U18567 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n14857) );
  NAND2_X1 U18568 ( .A1(n20970), .A2(n14852), .ZN(n14869) );
  AOI22_X1 U18569 ( .A1(n21024), .A2(P1_EBX_REG_27__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n21019), .ZN(n14853) );
  OAI21_X1 U18570 ( .B1(n14869), .B2(n14857), .A(n14853), .ZN(n14856) );
  NOR2_X1 U18571 ( .A1(n21015), .A2(n14854), .ZN(n14855) );
  AOI211_X1 U18572 ( .C1(n14858), .C2(n14857), .A(n14856), .B(n14855), .ZN(
        n14859) );
  OAI211_X1 U18573 ( .C1(n15541), .C2(n21026), .A(n14860), .B(n14859), .ZN(
        P1_U2813) );
  OAI21_X1 U18574 ( .B1(n14896), .B2(n14877), .A(n14861), .ZN(n14863) );
  NAND2_X1 U18575 ( .A1(n14863), .A2(n14862), .ZN(n15550) );
  INV_X1 U18577 ( .A(n15322), .ZN(n14866) );
  NAND2_X1 U18578 ( .A1(n14866), .A2(n20982), .ZN(n14873) );
  INV_X1 U18579 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n21835) );
  NOR3_X1 U18580 ( .A1(n14878), .A2(P1_REIP_REG_26__SCAN_IN), .A3(n21835), 
        .ZN(n14871) );
  INV_X1 U18581 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n14868) );
  AOI22_X1 U18582 ( .A1(n21024), .A2(P1_EBX_REG_26__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n21019), .ZN(n14867) );
  OAI21_X1 U18583 ( .B1(n14869), .B2(n14868), .A(n14867), .ZN(n14870) );
  AOI211_X1 U18584 ( .C1(n21027), .C2(n15324), .A(n14871), .B(n14870), .ZN(
        n14872) );
  OAI211_X1 U18585 ( .C1(n21026), .C2(n15550), .A(n14873), .B(n14872), .ZN(
        P1_U2814) );
  AOI21_X1 U18586 ( .B1(n14876), .B2(n14874), .A(n14875), .ZN(n15333) );
  INV_X1 U18587 ( .A(n15333), .ZN(n15233) );
  XOR2_X1 U18588 ( .A(n14877), .B(n14896), .Z(n15563) );
  INV_X1 U18589 ( .A(n14878), .ZN(n14883) );
  OAI22_X1 U18590 ( .A1(n21003), .A2(n21702), .B1(n14879), .B2(n21001), .ZN(
        n14882) );
  NOR3_X1 U18591 ( .A1(n20968), .A2(n14880), .A3(n21835), .ZN(n14881) );
  AOI211_X1 U18592 ( .C1(n14883), .C2(n21835), .A(n14882), .B(n14881), .ZN(
        n14884) );
  OAI21_X1 U18593 ( .B1(n21015), .B2(n15331), .A(n14884), .ZN(n14885) );
  AOI21_X1 U18594 ( .B1(n15563), .B2(n20992), .A(n14885), .ZN(n14886) );
  OAI21_X1 U18595 ( .B1(n15233), .B2(n15112), .A(n14886), .ZN(P1_U2815) );
  INV_X1 U18596 ( .A(n14874), .ZN(n14888) );
  AOI21_X1 U18597 ( .B1(n14889), .B2(n14887), .A(n14888), .ZN(n15341) );
  INV_X1 U18598 ( .A(n15341), .ZN(n15238) );
  NAND2_X1 U18599 ( .A1(n20970), .A2(n14890), .ZN(n14907) );
  NAND2_X1 U18600 ( .A1(n14891), .A2(n14894), .ZN(n14893) );
  AOI22_X1 U18601 ( .A1(n21024), .A2(P1_EBX_REG_24__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n21019), .ZN(n14892) );
  OAI211_X1 U18602 ( .C1(n14907), .C2(n14894), .A(n14893), .B(n14892), .ZN(
        n14895) );
  AOI21_X1 U18603 ( .B1(n21027), .B2(n15337), .A(n14895), .ZN(n14900) );
  NAND2_X1 U18604 ( .A1(n14925), .A2(n14904), .ZN(n14897) );
  AOI21_X1 U18605 ( .B1(n14898), .B2(n14897), .A(n10528), .ZN(n15575) );
  NAND2_X1 U18606 ( .A1(n15575), .A2(n20992), .ZN(n14899) );
  OAI211_X1 U18607 ( .C1(n15238), .C2(n15112), .A(n14900), .B(n14899), .ZN(
        P1_U2816) );
  OAI21_X1 U18609 ( .B1(n14902), .B2(n14903), .A(n14887), .ZN(n15349) );
  XNOR2_X1 U18610 ( .A(n14925), .B(n14904), .ZN(n15586) );
  INV_X1 U18611 ( .A(n15586), .ZN(n14911) );
  NOR2_X1 U18612 ( .A1(n21015), .A2(n15343), .ZN(n14910) );
  INV_X1 U18613 ( .A(n14905), .ZN(n14919) );
  AOI21_X1 U18614 ( .B1(n14919), .B2(P1_REIP_REG_22__SCAN_IN), .A(
        P1_REIP_REG_23__SCAN_IN), .ZN(n14908) );
  AOI22_X1 U18615 ( .A1(n21024), .A2(P1_EBX_REG_23__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n21019), .ZN(n14906) );
  OAI21_X1 U18616 ( .B1(n14908), .B2(n14907), .A(n14906), .ZN(n14909) );
  AOI211_X1 U18617 ( .C1(n14911), .C2(n20992), .A(n14910), .B(n14909), .ZN(
        n14912) );
  OAI21_X1 U18618 ( .B1(n15349), .B2(n15112), .A(n14912), .ZN(P1_U2817) );
  INV_X1 U18619 ( .A(n14902), .ZN(n14914) );
  OAI21_X1 U18620 ( .B1(n14915), .B2(n14913), .A(n14914), .ZN(n15354) );
  INV_X1 U18621 ( .A(n14916), .ZN(n14936) );
  NAND2_X1 U18622 ( .A1(n15158), .A2(n14936), .ZN(n14917) );
  AND2_X1 U18623 ( .A1(n20970), .A2(n14917), .ZN(n14935) );
  AOI21_X1 U18624 ( .B1(n21016), .B2(n14939), .A(n14935), .ZN(n14922) );
  INV_X1 U18625 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n14921) );
  INV_X1 U18626 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n15353) );
  OAI22_X1 U18627 ( .A1(n21003), .A2(n15180), .B1(n15353), .B2(n21001), .ZN(
        n14918) );
  AOI21_X1 U18628 ( .B1(n14919), .B2(n14921), .A(n14918), .ZN(n14920) );
  OAI21_X1 U18629 ( .B1(n14922), .B2(n14921), .A(n14920), .ZN(n14927) );
  NOR2_X1 U18630 ( .A1(n14934), .A2(n14923), .ZN(n14924) );
  OR2_X1 U18631 ( .A1(n14925), .A2(n14924), .ZN(n15598) );
  NOR2_X1 U18632 ( .A1(n15598), .A2(n21026), .ZN(n14926) );
  AOI211_X1 U18633 ( .C1(n21027), .C2(n15357), .A(n14927), .B(n14926), .ZN(
        n14928) );
  OAI21_X1 U18634 ( .B1(n15354), .B2(n15112), .A(n14928), .ZN(P1_U2818) );
  INV_X1 U18635 ( .A(n14930), .ZN(n14931) );
  AOI21_X1 U18636 ( .B1(n10273), .B2(n14931), .A(n14913), .ZN(n15365) );
  INV_X1 U18637 ( .A(n15365), .ZN(n15250) );
  AND2_X1 U18638 ( .A1(n14954), .A2(n14932), .ZN(n14933) );
  NOR2_X1 U18639 ( .A1(n14934), .A2(n14933), .ZN(n15608) );
  INV_X1 U18640 ( .A(n14935), .ZN(n14948) );
  AOI22_X1 U18641 ( .A1(n21024), .A2(P1_EBX_REG_21__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n21019), .ZN(n14938) );
  NAND3_X1 U18642 ( .A1(n21016), .A2(n14939), .A3(n14936), .ZN(n14937) );
  OAI211_X1 U18643 ( .C1(n14948), .C2(n14939), .A(n14938), .B(n14937), .ZN(
        n14941) );
  NOR2_X1 U18644 ( .A1(n21015), .A2(n15363), .ZN(n14940) );
  AOI211_X1 U18645 ( .C1(n15608), .C2(n20992), .A(n14941), .B(n14940), .ZN(
        n14942) );
  OAI21_X1 U18646 ( .B1(n15250), .B2(n15112), .A(n14942), .ZN(P1_U2819) );
  AND2_X1 U18647 ( .A1(n14943), .A2(n14944), .ZN(n14945) );
  OR2_X1 U18648 ( .A1(n14945), .A2(n14930), .ZN(n15371) );
  AOI21_X1 U18649 ( .B1(n21016), .B2(n14946), .A(P1_REIP_REG_20__SCAN_IN), 
        .ZN(n14947) );
  NOR2_X1 U18650 ( .A1(n14948), .A2(n14947), .ZN(n14951) );
  INV_X1 U18651 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n14949) );
  INV_X1 U18652 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n15370) );
  OAI22_X1 U18653 ( .A1(n21003), .A2(n14949), .B1(n15370), .B2(n21001), .ZN(
        n14950) );
  AOI211_X1 U18654 ( .C1(n21027), .C2(n15374), .A(n14951), .B(n14950), .ZN(
        n14956) );
  NAND2_X1 U18655 ( .A1(n14960), .A2(n14952), .ZN(n14953) );
  AND2_X1 U18656 ( .A1(n14954), .A2(n14953), .ZN(n15621) );
  NAND2_X1 U18657 ( .A1(n15621), .A2(n20992), .ZN(n14955) );
  OAI211_X1 U18658 ( .C1(n15371), .C2(n15112), .A(n14956), .B(n14955), .ZN(
        P1_U2820) );
  NAND2_X1 U18659 ( .A1(n14957), .A2(n14958), .ZN(n14959) );
  NAND2_X1 U18660 ( .A1(n14943), .A2(n14959), .ZN(n15379) );
  OAI21_X1 U18661 ( .B1(n14984), .B2(n14961), .A(n14960), .ZN(n15625) );
  NAND2_X1 U18662 ( .A1(n15158), .A2(n14962), .ZN(n20986) );
  OAI21_X1 U18663 ( .B1(n21001), .B2(n15378), .A(n20986), .ZN(n14965) );
  INV_X1 U18664 ( .A(n21016), .ZN(n20999) );
  NOR3_X1 U18665 ( .A1(n20999), .A2(P1_REIP_REG_19__SCAN_IN), .A3(n14963), 
        .ZN(n14964) );
  AOI211_X1 U18666 ( .C1(P1_EBX_REG_19__SCAN_IN), .C2(n21024), .A(n14965), .B(
        n14964), .ZN(n14977) );
  NAND2_X1 U18667 ( .A1(n21016), .A2(n14966), .ZN(n15125) );
  INV_X1 U18668 ( .A(n14967), .ZN(n14972) );
  OR2_X1 U18669 ( .A1(n15125), .A2(n14972), .ZN(n15015) );
  INV_X1 U18670 ( .A(n14968), .ZN(n14974) );
  NOR3_X1 U18671 ( .A1(n15015), .A2(P1_REIP_REG_18__SCAN_IN), .A3(n14974), 
        .ZN(n14987) );
  INV_X1 U18672 ( .A(n20961), .ZN(n14969) );
  AND2_X1 U18673 ( .A1(n15158), .A2(n14969), .ZN(n20967) );
  INV_X1 U18674 ( .A(n14970), .ZN(n14971) );
  NAND2_X1 U18675 ( .A1(n20967), .A2(n14971), .ZN(n15061) );
  NAND2_X1 U18676 ( .A1(n20970), .A2(n15061), .ZN(n15116) );
  NAND2_X1 U18677 ( .A1(n20970), .A2(n14972), .ZN(n14973) );
  NAND2_X1 U18678 ( .A1(n15116), .A2(n14973), .ZN(n15044) );
  AND2_X1 U18679 ( .A1(n20970), .A2(n14974), .ZN(n14975) );
  OR2_X1 U18680 ( .A1(n15044), .A2(n14975), .ZN(n15000) );
  OAI21_X1 U18681 ( .B1(n14987), .B2(n15000), .A(P1_REIP_REG_19__SCAN_IN), 
        .ZN(n14976) );
  OAI211_X1 U18682 ( .C1(n15625), .C2(n21026), .A(n14977), .B(n14976), .ZN(
        n14978) );
  AOI21_X1 U18683 ( .B1(n15382), .B2(n21027), .A(n14978), .ZN(n14979) );
  OAI21_X1 U18684 ( .B1(n15379), .B2(n15112), .A(n14979), .ZN(P1_U2821) );
  XOR2_X1 U18685 ( .A(n14981), .B(n14980), .Z(n15390) );
  INV_X1 U18686 ( .A(n15390), .ZN(n15265) );
  INV_X1 U18687 ( .A(n15011), .ZN(n14983) );
  AOI21_X1 U18688 ( .B1(n14983), .B2(n15001), .A(n14982), .ZN(n14985) );
  OR2_X1 U18689 ( .A1(n14985), .A2(n14984), .ZN(n15641) );
  INV_X1 U18690 ( .A(n20986), .ZN(n21009) );
  AOI21_X1 U18691 ( .B1(n21019), .B2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n21009), .ZN(n14986) );
  OAI21_X1 U18692 ( .B1(n21003), .B2(n15184), .A(n14986), .ZN(n14988) );
  AOI211_X1 U18693 ( .C1(P1_REIP_REG_18__SCAN_IN), .C2(n15000), .A(n14988), 
        .B(n14987), .ZN(n14989) );
  OAI21_X1 U18694 ( .B1(n21026), .B2(n15641), .A(n14989), .ZN(n14990) );
  AOI21_X1 U18695 ( .B1(n15386), .B2(n21027), .A(n14990), .ZN(n14991) );
  OAI21_X1 U18696 ( .B1(n15265), .B2(n15112), .A(n14991), .ZN(P1_U2822) );
  AOI21_X1 U18697 ( .B1(n14994), .B2(n14993), .A(n14980), .ZN(n15401) );
  NAND2_X1 U18698 ( .A1(n15401), .A2(n20982), .ZN(n15006) );
  NAND2_X1 U18699 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(P1_REIP_REG_15__SCAN_IN), 
        .ZN(n14995) );
  INV_X1 U18700 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n21564) );
  OAI21_X1 U18701 ( .B1(n15015), .B2(n14995), .A(n21564), .ZN(n14999) );
  INV_X1 U18702 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n14997) );
  NAND2_X1 U18703 ( .A1(n21019), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n14996) );
  OAI211_X1 U18704 ( .C1(n21003), .C2(n14997), .A(n20986), .B(n14996), .ZN(
        n14998) );
  AOI21_X1 U18705 ( .B1(n15000), .B2(n14999), .A(n14998), .ZN(n15005) );
  XNOR2_X1 U18706 ( .A(n15011), .B(n15001), .ZN(n15652) );
  NAND2_X1 U18707 ( .A1(n15652), .A2(n20992), .ZN(n15004) );
  INV_X1 U18708 ( .A(n15399), .ZN(n15002) );
  NAND2_X1 U18709 ( .A1(n21027), .A2(n15002), .ZN(n15003) );
  NAND4_X1 U18710 ( .A1(n15006), .A2(n15005), .A3(n15004), .A4(n15003), .ZN(
        P1_U2823) );
  AOI21_X1 U18711 ( .B1(n15009), .B2(n15008), .A(n10274), .ZN(n15410) );
  INV_X1 U18712 ( .A(n15410), .ZN(n15278) );
  OAI21_X1 U18713 ( .B1(n15039), .B2(n15024), .A(n15010), .ZN(n15012) );
  AND2_X1 U18714 ( .A1(n15012), .A2(n15011), .ZN(n15663) );
  INV_X1 U18715 ( .A(n15663), .ZN(n15018) );
  OAI21_X1 U18716 ( .B1(n21001), .B2(n10151), .A(n20986), .ZN(n15014) );
  INV_X1 U18717 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n21561) );
  NOR3_X1 U18718 ( .A1(n15015), .A2(P1_REIP_REG_16__SCAN_IN), .A3(n21561), 
        .ZN(n15013) );
  AOI211_X1 U18719 ( .C1(P1_EBX_REG_16__SCAN_IN), .C2(n21024), .A(n15014), .B(
        n15013), .ZN(n15017) );
  NOR2_X1 U18720 ( .A1(n15015), .A2(P1_REIP_REG_15__SCAN_IN), .ZN(n15026) );
  OAI21_X1 U18721 ( .B1(n15026), .B2(n15044), .A(P1_REIP_REG_16__SCAN_IN), 
        .ZN(n15016) );
  OAI211_X1 U18722 ( .C1(n15018), .C2(n21026), .A(n15017), .B(n15016), .ZN(
        n15019) );
  AOI21_X1 U18723 ( .B1(n15407), .B2(n21027), .A(n15019), .ZN(n15020) );
  OAI21_X1 U18724 ( .B1(n15278), .B2(n15112), .A(n15020), .ZN(P1_U2824) );
  INV_X1 U18725 ( .A(n15087), .ZN(n15052) );
  INV_X1 U18726 ( .A(n15021), .ZN(n15050) );
  NAND2_X1 U18727 ( .A1(n15050), .A2(n15049), .ZN(n15051) );
  OAI21_X1 U18728 ( .B1(n15052), .B2(n15021), .A(n15051), .ZN(n15022) );
  OAI21_X1 U18729 ( .B1(n15034), .B2(n15023), .A(n15008), .ZN(n15419) );
  XOR2_X1 U18730 ( .A(n15024), .B(n15039), .Z(n15671) );
  INV_X1 U18731 ( .A(n15044), .ZN(n15029) );
  OAI21_X1 U18732 ( .B1(n21001), .B2(n15025), .A(n20986), .ZN(n15027) );
  AOI211_X1 U18733 ( .C1(P1_EBX_REG_15__SCAN_IN), .C2(n21024), .A(n15027), .B(
        n15026), .ZN(n15028) );
  OAI21_X1 U18734 ( .B1(n15029), .B2(n21561), .A(n15028), .ZN(n15031) );
  NOR2_X1 U18735 ( .A1(n21015), .A2(n15421), .ZN(n15030) );
  AOI211_X1 U18736 ( .C1(n20992), .C2(n15671), .A(n15031), .B(n15030), .ZN(
        n15032) );
  OAI21_X1 U18737 ( .B1(n15419), .B2(n15112), .A(n15032), .ZN(P1_U2825) );
  INV_X1 U18738 ( .A(n15033), .ZN(n15036) );
  INV_X1 U18739 ( .A(n15054), .ZN(n15035) );
  AOI21_X1 U18740 ( .B1(n15036), .B2(n15035), .A(n15034), .ZN(n15434) );
  NAND2_X1 U18741 ( .A1(n15434), .A2(n20982), .ZN(n15048) );
  OR2_X1 U18742 ( .A1(n15057), .A2(n15037), .ZN(n15038) );
  AND2_X1 U18743 ( .A1(n15039), .A2(n15038), .ZN(n15675) );
  NAND2_X1 U18744 ( .A1(n21019), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15040) );
  OAI211_X1 U18745 ( .C1(n21003), .C2(n15041), .A(n20986), .B(n15040), .ZN(
        n15046) );
  OR3_X1 U18746 ( .A1(n15125), .A2(n15060), .A3(n21558), .ZN(n15042) );
  NAND2_X1 U18747 ( .A1(n15042), .A2(n21557), .ZN(n15043) );
  AND2_X1 U18748 ( .A1(n15044), .A2(n15043), .ZN(n15045) );
  AOI211_X1 U18749 ( .C1(n15675), .C2(n20992), .A(n15046), .B(n15045), .ZN(
        n15047) );
  OAI211_X1 U18750 ( .C1(n21015), .C2(n15432), .A(n15048), .B(n15047), .ZN(
        P1_U2826) );
  OAI21_X1 U18751 ( .B1(n15050), .B2(n15049), .A(n15051), .ZN(n15088) );
  OAI21_X1 U18752 ( .B1(n15088), .B2(n15052), .A(n15051), .ZN(n15070) );
  NAND2_X1 U18753 ( .A1(n15070), .A2(n15069), .ZN(n15068) );
  INV_X1 U18754 ( .A(n15053), .ZN(n15055) );
  AOI21_X1 U18755 ( .B1(n15068), .B2(n15055), .A(n15054), .ZN(n15446) );
  NAND2_X1 U18756 ( .A1(n15446), .A2(n20982), .ZN(n15067) );
  INV_X1 U18757 ( .A(n15056), .ZN(n15059) );
  INV_X1 U18758 ( .A(n15074), .ZN(n15058) );
  AOI21_X1 U18759 ( .B1(n15059), .B2(n15058), .A(n15057), .ZN(n15682) );
  NOR3_X1 U18760 ( .A1(n15125), .A2(P1_REIP_REG_13__SCAN_IN), .A3(n15060), 
        .ZN(n15065) );
  OR2_X1 U18761 ( .A1(n15061), .A2(n15060), .ZN(n15081) );
  NAND3_X1 U18762 ( .A1(n20970), .A2(P1_REIP_REG_13__SCAN_IN), .A3(n15081), 
        .ZN(n15063) );
  AOI21_X1 U18763 ( .B1(n21019), .B2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n21009), .ZN(n15062) );
  OAI211_X1 U18764 ( .C1(n15190), .C2(n21003), .A(n15063), .B(n15062), .ZN(
        n15064) );
  AOI211_X1 U18765 ( .C1(n15682), .C2(n20992), .A(n15065), .B(n15064), .ZN(
        n15066) );
  OAI211_X1 U18766 ( .C1(n21015), .C2(n15444), .A(n15067), .B(n15066), .ZN(
        P1_U2827) );
  OAI21_X1 U18767 ( .B1(n15070), .B2(n15069), .A(n15068), .ZN(n15456) );
  INV_X1 U18768 ( .A(n15456), .ZN(n15071) );
  NAND2_X1 U18769 ( .A1(n15071), .A2(n20982), .ZN(n15086) );
  AND2_X1 U18770 ( .A1(n15092), .A2(n15072), .ZN(n15073) );
  NOR2_X1 U18771 ( .A1(n15074), .A2(n15073), .ZN(n15701) );
  INV_X1 U18772 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n15076) );
  NAND2_X1 U18773 ( .A1(n21019), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15075) );
  OAI211_X1 U18774 ( .C1(n21003), .C2(n15076), .A(n20986), .B(n15075), .ZN(
        n15077) );
  AOI21_X1 U18775 ( .B1(n15701), .B2(n20992), .A(n15077), .ZN(n15085) );
  INV_X1 U18776 ( .A(n15078), .ZN(n15453) );
  NAND2_X1 U18777 ( .A1(n21027), .A2(n15453), .ZN(n15084) );
  INV_X1 U18778 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n21554) );
  NAND2_X1 U18779 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(P1_REIP_REG_9__SCAN_IN), 
        .ZN(n15093) );
  OR3_X1 U18780 ( .A1(n15125), .A2(n21554), .A3(n15093), .ZN(n15080) );
  INV_X1 U18781 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n15079) );
  NAND2_X1 U18782 ( .A1(n15080), .A2(n15079), .ZN(n15082) );
  NAND3_X1 U18783 ( .A1(n15082), .A2(n20970), .A3(n15081), .ZN(n15083) );
  NAND4_X1 U18784 ( .A1(n15086), .A2(n15085), .A3(n15084), .A4(n15083), .ZN(
        P1_U2828) );
  XNOR2_X1 U18785 ( .A(n15088), .B(n15087), .ZN(n15462) );
  NAND2_X1 U18786 ( .A1(n15462), .A2(n20982), .ZN(n15099) );
  INV_X1 U18787 ( .A(n15093), .ZN(n15089) );
  OAI21_X1 U18788 ( .B1(n20968), .B2(n15089), .A(n15116), .ZN(n15105) );
  NAND2_X1 U18789 ( .A1(n15103), .A2(n15090), .ZN(n15091) );
  NAND2_X1 U18790 ( .A1(n15092), .A2(n15091), .ZN(n15708) );
  NOR3_X1 U18791 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(n15093), .A3(n15125), 
        .ZN(n15094) );
  AOI211_X1 U18792 ( .C1(n21019), .C2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n15094), .B(n21009), .ZN(n15096) );
  NAND2_X1 U18793 ( .A1(n21024), .A2(P1_EBX_REG_11__SCAN_IN), .ZN(n15095) );
  OAI211_X1 U18794 ( .C1(n21026), .C2(n15708), .A(n15096), .B(n15095), .ZN(
        n15097) );
  AOI21_X1 U18795 ( .B1(n15105), .B2(P1_REIP_REG_11__SCAN_IN), .A(n15097), 
        .ZN(n15098) );
  OAI211_X1 U18796 ( .C1(n21015), .C2(n15460), .A(n15099), .B(n15098), .ZN(
        P1_U2829) );
  OAI21_X1 U18797 ( .B1(n9719), .B2(n15100), .A(n15021), .ZN(n15473) );
  OR2_X1 U18798 ( .A1(n15121), .A2(n15101), .ZN(n15102) );
  NAND2_X1 U18799 ( .A1(n15103), .A2(n15102), .ZN(n15721) );
  INV_X1 U18800 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n15104) );
  NOR2_X1 U18801 ( .A1(n15125), .A2(n15104), .ZN(n15106) );
  OAI21_X1 U18802 ( .B1(P1_REIP_REG_10__SCAN_IN), .B2(n15106), .A(n15105), 
        .ZN(n15109) );
  OAI21_X1 U18803 ( .B1(n21001), .B2(n10156), .A(n20986), .ZN(n15107) );
  AOI21_X1 U18804 ( .B1(n21024), .B2(P1_EBX_REG_10__SCAN_IN), .A(n15107), .ZN(
        n15108) );
  OAI211_X1 U18805 ( .C1(n15721), .C2(n21026), .A(n15109), .B(n15108), .ZN(
        n15110) );
  AOI21_X1 U18806 ( .B1(n21027), .B2(n15470), .A(n15110), .ZN(n15111) );
  OAI21_X1 U18807 ( .B1(n15473), .B2(n15112), .A(n15111), .ZN(P1_U2830) );
  NOR2_X1 U18808 ( .A1(n15113), .A2(n15114), .ZN(n15115) );
  OR2_X1 U18809 ( .A1(n9719), .A2(n15115), .ZN(n15293) );
  INV_X1 U18810 ( .A(n15293), .ZN(n15482) );
  NAND2_X1 U18811 ( .A1(n15482), .A2(n20982), .ZN(n15128) );
  INV_X1 U18812 ( .A(n15116), .ZN(n15136) );
  INV_X1 U18813 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n15194) );
  NAND2_X1 U18814 ( .A1(n21019), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15117) );
  OAI211_X1 U18815 ( .C1(n21003), .C2(n15194), .A(n20986), .B(n15117), .ZN(
        n15118) );
  INV_X1 U18816 ( .A(n15118), .ZN(n15124) );
  NOR2_X1 U18817 ( .A1(n15134), .A2(n15119), .ZN(n15120) );
  OR2_X1 U18818 ( .A1(n15121), .A2(n15120), .ZN(n15731) );
  INV_X1 U18819 ( .A(n15731), .ZN(n15122) );
  NAND2_X1 U18820 ( .A1(n20992), .A2(n15122), .ZN(n15123) );
  OAI211_X1 U18821 ( .C1(n15125), .C2(P1_REIP_REG_9__SCAN_IN), .A(n15124), .B(
        n15123), .ZN(n15126) );
  AOI21_X1 U18822 ( .B1(P1_REIP_REG_9__SCAN_IN), .B2(n15136), .A(n15126), .ZN(
        n15127) );
  OAI211_X1 U18823 ( .C1(n21015), .C2(n15480), .A(n15128), .B(n15127), .ZN(
        P1_U2831) );
  AOI21_X1 U18824 ( .B1(n15130), .B2(n15129), .A(n15113), .ZN(n15490) );
  INV_X1 U18825 ( .A(n15488), .ZN(n15131) );
  NAND2_X1 U18826 ( .A1(n21027), .A2(n15131), .ZN(n15141) );
  INV_X1 U18827 ( .A(n15132), .ZN(n15202) );
  AOI21_X1 U18828 ( .B1(n15202), .B2(n15201), .A(n15133), .ZN(n15135) );
  OR2_X1 U18829 ( .A1(n15135), .A2(n15134), .ZN(n15751) );
  INV_X1 U18830 ( .A(n15751), .ZN(n15197) );
  AOI22_X1 U18831 ( .A1(n21024), .A2(P1_EBX_REG_8__SCAN_IN), .B1(
        P1_REIP_REG_8__SCAN_IN), .B2(n15136), .ZN(n15137) );
  OAI211_X1 U18832 ( .C1(n21001), .C2(n15138), .A(n15137), .B(n20986), .ZN(
        n15139) );
  AOI21_X1 U18833 ( .B1(n20992), .B2(n15197), .A(n15139), .ZN(n15140) );
  NAND2_X1 U18834 ( .A1(n15141), .A2(n15140), .ZN(n15144) );
  NAND3_X1 U18835 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(P1_REIP_REG_6__SCAN_IN), 
        .A3(P1_REIP_REG_5__SCAN_IN), .ZN(n15142) );
  NOR4_X1 U18836 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n20961), .A3(n20999), .A4(
        n15142), .ZN(n15143) );
  AOI211_X1 U18837 ( .C1(n15490), .C2(n20982), .A(n15144), .B(n15143), .ZN(
        n15145) );
  INV_X1 U18838 ( .A(n15145), .ZN(P1_U2832) );
  INV_X1 U18839 ( .A(n15149), .ZN(n15146) );
  AOI21_X1 U18840 ( .B1(n15147), .B2(n15146), .A(n20982), .ZN(n21010) );
  INV_X1 U18841 ( .A(n15148), .ZN(n15506) );
  INV_X1 U18842 ( .A(n14439), .ZN(n15774) );
  OR2_X1 U18843 ( .A1(n15149), .A2(n13439), .ZN(n21021) );
  INV_X1 U18844 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n21603) );
  NOR4_X1 U18845 ( .A1(n20999), .A2(n14277), .A3(P1_REIP_REG_3__SCAN_IN), .A4(
        n21603), .ZN(n15150) );
  AOI21_X1 U18846 ( .B1(n21111), .B2(n20992), .A(n15150), .ZN(n15152) );
  AOI22_X1 U18847 ( .A1(n21024), .A2(P1_EBX_REG_3__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n21019), .ZN(n15151) );
  OAI211_X1 U18848 ( .C1(n15774), .C2(n21021), .A(n15152), .B(n15151), .ZN(
        n15156) );
  NAND2_X1 U18849 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_2__SCAN_IN), 
        .ZN(n15154) );
  AOI21_X1 U18850 ( .B1(n21016), .B2(n15154), .A(n15153), .ZN(n21030) );
  INV_X1 U18851 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n21545) );
  NOR2_X1 U18852 ( .A1(n21030), .A2(n21545), .ZN(n15155) );
  AOI211_X1 U18853 ( .C1(n21027), .C2(n15506), .A(n15156), .B(n15155), .ZN(
        n15157) );
  OAI21_X1 U18854 ( .B1(n21010), .B2(n15510), .A(n15157), .ZN(P1_U2837) );
  OAI22_X1 U18855 ( .A1(n21021), .A2(n13944), .B1(n21603), .B2(n15158), .ZN(
        n15161) );
  OAI22_X1 U18856 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(n20999), .B1(n21026), 
        .B2(n15159), .ZN(n15160) );
  AOI211_X1 U18857 ( .C1(n21024), .C2(P1_EBX_REG_1__SCAN_IN), .A(n15161), .B(
        n15160), .ZN(n15163) );
  MUX2_X1 U18858 ( .A(n21015), .B(n21001), .S(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .Z(n15162) );
  OAI211_X1 U18859 ( .C1(n21010), .C2(n15164), .A(n15163), .B(n15162), .ZN(
        P1_U2839) );
  OAI22_X1 U18860 ( .A1(n21003), .A2(n12635), .B1(n15165), .B2(n21021), .ZN(
        n15168) );
  NOR2_X1 U18861 ( .A1(n21026), .A2(n15166), .ZN(n15167) );
  AOI211_X1 U18862 ( .C1(P1_REIP_REG_0__SCAN_IN), .C2(n20970), .A(n15168), .B(
        n15167), .ZN(n15170) );
  OAI21_X1 U18863 ( .B1(n21027), .B2(n21019), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n15169) );
  OAI211_X1 U18864 ( .C1(n21010), .C2(n15171), .A(n15170), .B(n15169), .ZN(
        P1_U2840) );
  OAI22_X1 U18865 ( .A1(n15512), .A2(n15203), .B1(n15204), .B2(n15172), .ZN(
        P1_U2841) );
  OAI222_X1 U18866 ( .A1(n15206), .A2(n15306), .B1(n15173), .B2(n15204), .C1(
        n15527), .C2(n15203), .ZN(P1_U2843) );
  INV_X1 U18867 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n15174) );
  OAI222_X1 U18868 ( .A1(n15206), .A2(n15216), .B1(n15174), .B2(n15204), .C1(
        n15534), .C2(n15203), .ZN(P1_U2844) );
  OAI222_X1 U18869 ( .A1(n15222), .A2(n15206), .B1(n15175), .B2(n15204), .C1(
        n15203), .C2(n15541), .ZN(P1_U2845) );
  INV_X1 U18870 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n15176) );
  OAI222_X1 U18871 ( .A1(n15206), .A2(n15322), .B1(n15176), .B2(n15204), .C1(
        n15550), .C2(n15203), .ZN(P1_U2846) );
  INV_X1 U18872 ( .A(n15563), .ZN(n15177) );
  OAI222_X1 U18873 ( .A1(n15233), .A2(n15206), .B1(n21702), .B2(n15204), .C1(
        n15203), .C2(n15177), .ZN(P1_U2847) );
  AOI22_X1 U18874 ( .A1(n15575), .A2(n15196), .B1(P1_EBX_REG_24__SCAN_IN), 
        .B2(n15195), .ZN(n15178) );
  OAI21_X1 U18875 ( .B1(n15238), .B2(n15206), .A(n15178), .ZN(P1_U2848) );
  INV_X1 U18876 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n15179) );
  OAI222_X1 U18877 ( .A1(n15349), .A2(n15206), .B1(n15179), .B2(n15204), .C1(
        n15203), .C2(n15586), .ZN(P1_U2849) );
  OAI222_X1 U18878 ( .A1(n15354), .A2(n15206), .B1(n15180), .B2(n15204), .C1(
        n15598), .C2(n15203), .ZN(P1_U2850) );
  AOI22_X1 U18879 ( .A1(n15608), .A2(n15196), .B1(P1_EBX_REG_21__SCAN_IN), 
        .B2(n15195), .ZN(n15181) );
  OAI21_X1 U18880 ( .B1(n15250), .B2(n15206), .A(n15181), .ZN(P1_U2851) );
  AOI22_X1 U18881 ( .A1(n15621), .A2(n15196), .B1(P1_EBX_REG_20__SCAN_IN), 
        .B2(n15195), .ZN(n15182) );
  OAI21_X1 U18882 ( .B1(n15371), .B2(n15206), .A(n15182), .ZN(P1_U2852) );
  INV_X1 U18883 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n15183) );
  OAI222_X1 U18884 ( .A1(n15206), .A2(n15379), .B1(n15183), .B2(n15204), .C1(
        n15625), .C2(n15203), .ZN(P1_U2853) );
  OAI222_X1 U18885 ( .A1(n15265), .A2(n15206), .B1(n15184), .B2(n15204), .C1(
        n15641), .C2(n15203), .ZN(P1_U2854) );
  INV_X1 U18886 ( .A(n15401), .ZN(n15270) );
  AOI22_X1 U18887 ( .A1(n15652), .A2(n15196), .B1(P1_EBX_REG_17__SCAN_IN), 
        .B2(n15195), .ZN(n15185) );
  OAI21_X1 U18888 ( .B1(n15270), .B2(n15206), .A(n15185), .ZN(P1_U2855) );
  AOI22_X1 U18889 ( .A1(n15663), .A2(n15196), .B1(P1_EBX_REG_16__SCAN_IN), 
        .B2(n15195), .ZN(n15186) );
  OAI21_X1 U18890 ( .B1(n15278), .B2(n15206), .A(n15186), .ZN(P1_U2856) );
  AOI22_X1 U18891 ( .A1(n15671), .A2(n15196), .B1(P1_EBX_REG_15__SCAN_IN), 
        .B2(n15195), .ZN(n15187) );
  OAI21_X1 U18892 ( .B1(n15419), .B2(n15206), .A(n15187), .ZN(P1_U2857) );
  INV_X1 U18893 ( .A(n15434), .ZN(n15281) );
  AOI22_X1 U18894 ( .A1(n15675), .A2(n15196), .B1(P1_EBX_REG_14__SCAN_IN), 
        .B2(n15195), .ZN(n15188) );
  OAI21_X1 U18895 ( .B1(n15281), .B2(n15206), .A(n15188), .ZN(P1_U2858) );
  INV_X1 U18896 ( .A(n15446), .ZN(n15283) );
  INV_X1 U18897 ( .A(n15682), .ZN(n15189) );
  OAI222_X1 U18898 ( .A1(n15283), .A2(n15206), .B1(n15190), .B2(n15204), .C1(
        n15189), .C2(n15203), .ZN(P1_U2859) );
  AOI22_X1 U18899 ( .A1(n15701), .A2(n15196), .B1(P1_EBX_REG_12__SCAN_IN), 
        .B2(n15195), .ZN(n15191) );
  OAI21_X1 U18900 ( .B1(n15456), .B2(n15206), .A(n15191), .ZN(P1_U2860) );
  INV_X1 U18901 ( .A(n15462), .ZN(n15289) );
  OAI222_X1 U18902 ( .A1(n15289), .A2(n15206), .B1(n15192), .B2(n15204), .C1(
        n15708), .C2(n15203), .ZN(P1_U2861) );
  INV_X1 U18903 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n15193) );
  OAI222_X1 U18904 ( .A1(n15473), .A2(n15206), .B1(n15193), .B2(n15204), .C1(
        n15721), .C2(n15203), .ZN(P1_U2862) );
  OAI222_X1 U18905 ( .A1(n15293), .A2(n15206), .B1(n15194), .B2(n15204), .C1(
        n15731), .C2(n15203), .ZN(P1_U2863) );
  INV_X1 U18906 ( .A(n15490), .ZN(n15295) );
  AOI22_X1 U18907 ( .A1(n15197), .A2(n15196), .B1(P1_EBX_REG_8__SCAN_IN), .B2(
        n15195), .ZN(n15198) );
  OAI21_X1 U18908 ( .B1(n15295), .B2(n15206), .A(n15198), .ZN(P1_U2864) );
  INV_X1 U18909 ( .A(n15129), .ZN(n15199) );
  AOI21_X1 U18910 ( .B1(n15200), .B2(n14571), .A(n15199), .ZN(n20971) );
  INV_X1 U18911 ( .A(n20971), .ZN(n15299) );
  INV_X1 U18912 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n15205) );
  XNOR2_X1 U18913 ( .A(n15202), .B(n15201), .ZN(n20962) );
  OAI222_X1 U18914 ( .A1(n15299), .A2(n15206), .B1(n15205), .B2(n15204), .C1(
        n15203), .C2(n20962), .ZN(P1_U2865) );
  INV_X1 U18915 ( .A(DATAI_13_), .ZN(n15208) );
  INV_X1 U18916 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n15207) );
  MUX2_X1 U18917 ( .A(n15208), .B(n15207), .S(n15223), .Z(n21066) );
  OAI22_X1 U18918 ( .A1(n15272), .A2(n21066), .B1(n14002), .B2(n14816), .ZN(
        n15209) );
  AOI21_X1 U18919 ( .B1(BUF1_REG_29__SCAN_IN), .B2(n15274), .A(n15209), .ZN(
        n15211) );
  NAND2_X1 U18920 ( .A1(n15275), .A2(DATAI_29_), .ZN(n15210) );
  OAI211_X1 U18921 ( .C1(n15306), .C2(n15298), .A(n15211), .B(n15210), .ZN(
        P1_U2875) );
  OAI22_X1 U18922 ( .A1(n15272), .A2(n15285), .B1(n15212), .B2(n14816), .ZN(
        n15213) );
  AOI21_X1 U18923 ( .B1(BUF1_REG_28__SCAN_IN), .B2(n15274), .A(n15213), .ZN(
        n15215) );
  NAND2_X1 U18924 ( .A1(n15275), .A2(DATAI_28_), .ZN(n15214) );
  OAI211_X1 U18925 ( .C1(n15216), .C2(n15298), .A(n15215), .B(n15214), .ZN(
        P1_U2876) );
  INV_X1 U18926 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n21718) );
  INV_X1 U18927 ( .A(n15272), .ZN(n15256) );
  INV_X1 U18928 ( .A(DATAI_11_), .ZN(n15218) );
  NAND2_X1 U18929 ( .A1(n15223), .A2(BUF1_REG_11__SCAN_IN), .ZN(n15217) );
  OAI21_X1 U18930 ( .B1(n15223), .B2(n15218), .A(n15217), .ZN(n21064) );
  AOI22_X1 U18931 ( .A1(n15256), .A2(n21064), .B1(P1_EAX_REG_27__SCAN_IN), 
        .B2(n15286), .ZN(n15219) );
  OAI21_X1 U18932 ( .B1(n15258), .B2(n21718), .A(n15219), .ZN(n15220) );
  AOI21_X1 U18933 ( .B1(n15275), .B2(DATAI_27_), .A(n15220), .ZN(n15221) );
  OAI21_X1 U18934 ( .B1(n15222), .B2(n15298), .A(n15221), .ZN(P1_U2877) );
  INV_X1 U18935 ( .A(DATAI_10_), .ZN(n15224) );
  INV_X1 U18936 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n18133) );
  MUX2_X1 U18937 ( .A(n15224), .B(n18133), .S(n15223), .Z(n21061) );
  OAI22_X1 U18938 ( .A1(n15272), .A2(n21061), .B1(n15225), .B2(n14816), .ZN(
        n15226) );
  AOI21_X1 U18939 ( .B1(n15274), .B2(BUF1_REG_26__SCAN_IN), .A(n15226), .ZN(
        n15228) );
  NAND2_X1 U18940 ( .A1(n15275), .A2(DATAI_26_), .ZN(n15227) );
  OAI211_X1 U18941 ( .C1(n15322), .C2(n15298), .A(n15228), .B(n15227), .ZN(
        P1_U2878) );
  OAI22_X1 U18942 ( .A1(n15272), .A2(n15292), .B1(n15229), .B2(n14816), .ZN(
        n15230) );
  AOI21_X1 U18943 ( .B1(n15274), .B2(BUF1_REG_25__SCAN_IN), .A(n15230), .ZN(
        n15232) );
  NAND2_X1 U18944 ( .A1(n15275), .A2(DATAI_25_), .ZN(n15231) );
  OAI211_X1 U18945 ( .C1(n15233), .C2(n15298), .A(n15232), .B(n15231), .ZN(
        P1_U2879) );
  OAI22_X1 U18946 ( .A1(n15272), .A2(n15294), .B1(n15234), .B2(n14816), .ZN(
        n15235) );
  AOI21_X1 U18947 ( .B1(n15274), .B2(BUF1_REG_24__SCAN_IN), .A(n15235), .ZN(
        n15237) );
  NAND2_X1 U18948 ( .A1(n15275), .A2(DATAI_24_), .ZN(n15236) );
  OAI211_X1 U18949 ( .C1(n15238), .C2(n15298), .A(n15237), .B(n15236), .ZN(
        P1_U2880) );
  OAI22_X1 U18950 ( .A1(n15272), .A2(n15297), .B1(n14000), .B2(n14816), .ZN(
        n15239) );
  AOI21_X1 U18951 ( .B1(n15274), .B2(BUF1_REG_23__SCAN_IN), .A(n15239), .ZN(
        n15241) );
  NAND2_X1 U18952 ( .A1(n15275), .A2(DATAI_23_), .ZN(n15240) );
  OAI211_X1 U18953 ( .C1(n15349), .C2(n15298), .A(n15241), .B(n15240), .ZN(
        P1_U2881) );
  OAI22_X1 U18954 ( .A1(n15272), .A2(n15242), .B1(n14007), .B2(n14816), .ZN(
        n15243) );
  AOI21_X1 U18955 ( .B1(n15274), .B2(BUF1_REG_22__SCAN_IN), .A(n15243), .ZN(
        n15245) );
  NAND2_X1 U18956 ( .A1(n15275), .A2(DATAI_22_), .ZN(n15244) );
  OAI211_X1 U18957 ( .C1(n15354), .C2(n15298), .A(n15245), .B(n15244), .ZN(
        P1_U2882) );
  OAI22_X1 U18958 ( .A1(n15272), .A2(n15246), .B1(n21811), .B2(n14816), .ZN(
        n15247) );
  AOI21_X1 U18959 ( .B1(n15274), .B2(BUF1_REG_21__SCAN_IN), .A(n15247), .ZN(
        n15249) );
  NAND2_X1 U18960 ( .A1(n15275), .A2(DATAI_21_), .ZN(n15248) );
  OAI211_X1 U18961 ( .C1(n15250), .C2(n15298), .A(n15249), .B(n15248), .ZN(
        P1_U2883) );
  OAI22_X1 U18962 ( .A1(n15272), .A2(n15251), .B1(n13997), .B2(n14816), .ZN(
        n15252) );
  AOI21_X1 U18963 ( .B1(n15274), .B2(BUF1_REG_20__SCAN_IN), .A(n15252), .ZN(
        n15254) );
  NAND2_X1 U18964 ( .A1(n15275), .A2(DATAI_20_), .ZN(n15253) );
  OAI211_X1 U18965 ( .C1(n15371), .C2(n15298), .A(n15254), .B(n15253), .ZN(
        P1_U2884) );
  INV_X1 U18966 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n17570) );
  AOI22_X1 U18967 ( .A1(n15256), .A2(n15255), .B1(P1_EAX_REG_19__SCAN_IN), 
        .B2(n15286), .ZN(n15257) );
  OAI21_X1 U18968 ( .B1(n15258), .B2(n17570), .A(n15257), .ZN(n15259) );
  AOI21_X1 U18969 ( .B1(n15275), .B2(DATAI_19_), .A(n15259), .ZN(n15260) );
  OAI21_X1 U18970 ( .B1(n15379), .B2(n15298), .A(n15260), .ZN(P1_U2885) );
  OAI22_X1 U18971 ( .A1(n15272), .A2(n15261), .B1(n14122), .B2(n14816), .ZN(
        n15262) );
  AOI21_X1 U18972 ( .B1(n15274), .B2(BUF1_REG_18__SCAN_IN), .A(n15262), .ZN(
        n15264) );
  NAND2_X1 U18973 ( .A1(n15275), .A2(DATAI_18_), .ZN(n15263) );
  OAI211_X1 U18974 ( .C1(n15265), .C2(n15298), .A(n15264), .B(n15263), .ZN(
        P1_U2886) );
  OAI22_X1 U18975 ( .A1(n15272), .A2(n15266), .B1(n14120), .B2(n14816), .ZN(
        n15267) );
  AOI21_X1 U18976 ( .B1(n15274), .B2(BUF1_REG_17__SCAN_IN), .A(n15267), .ZN(
        n15269) );
  NAND2_X1 U18977 ( .A1(n15275), .A2(DATAI_17_), .ZN(n15268) );
  OAI211_X1 U18978 ( .C1(n15270), .C2(n15298), .A(n15269), .B(n15268), .ZN(
        P1_U2887) );
  OAI22_X1 U18979 ( .A1(n15272), .A2(n15271), .B1(n14125), .B2(n14816), .ZN(
        n15273) );
  AOI21_X1 U18980 ( .B1(n15274), .B2(BUF1_REG_16__SCAN_IN), .A(n15273), .ZN(
        n15277) );
  NAND2_X1 U18981 ( .A1(n15275), .A2(DATAI_16_), .ZN(n15276) );
  OAI211_X1 U18982 ( .C1(n15278), .C2(n15298), .A(n15277), .B(n15276), .ZN(
        P1_U2888) );
  OAI222_X1 U18983 ( .A1(n15419), .A2(n15298), .B1(n15296), .B2(n15280), .C1(
        n15279), .C2(n14816), .ZN(P1_U2889) );
  OAI222_X1 U18984 ( .A1(n15281), .A2(n15298), .B1(n21069), .B2(n15296), .C1(
        n21034), .C2(n14816), .ZN(P1_U2890) );
  INV_X1 U18985 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n15282) );
  OAI222_X1 U18986 ( .A1(n15283), .A2(n15298), .B1(n21066), .B2(n15296), .C1(
        n15282), .C2(n14816), .ZN(P1_U2891) );
  INV_X1 U18987 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n15284) );
  OAI222_X1 U18988 ( .A1(n15456), .A2(n15298), .B1(n15285), .B2(n15296), .C1(
        n15284), .C2(n14816), .ZN(P1_U2892) );
  INV_X1 U18989 ( .A(n15296), .ZN(n15287) );
  AOI22_X1 U18990 ( .A1(n15287), .A2(n21064), .B1(P1_EAX_REG_11__SCAN_IN), 
        .B2(n15286), .ZN(n15288) );
  OAI21_X1 U18991 ( .B1(n15289), .B2(n15298), .A(n15288), .ZN(P1_U2893) );
  INV_X1 U18992 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n15290) );
  OAI222_X1 U18993 ( .A1(n15473), .A2(n15298), .B1(n21061), .B2(n15296), .C1(
        n15290), .C2(n14816), .ZN(P1_U2894) );
  INV_X1 U18994 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n15291) );
  OAI222_X1 U18995 ( .A1(n15293), .A2(n15298), .B1(n15292), .B2(n15296), .C1(
        n15291), .C2(n14816), .ZN(P1_U2895) );
  OAI222_X1 U18996 ( .A1(n15295), .A2(n15298), .B1(n15294), .B2(n15296), .C1(
        n21043), .C2(n14816), .ZN(P1_U2896) );
  OAI222_X1 U18997 ( .A1(n15299), .A2(n15298), .B1(n15297), .B2(n15296), .C1(
        n14816), .C2(n12052), .ZN(P1_U2897) );
  NOR2_X1 U18998 ( .A1(n21123), .A2(n21580), .ZN(n15523) );
  NOR2_X1 U18999 ( .A1(n15300), .A2(n21098), .ZN(n15301) );
  AOI211_X1 U19000 ( .C1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .C2(n21088), .A(
        n15523), .B(n15301), .ZN(n15305) );
  NAND2_X1 U19001 ( .A1(n15520), .A2(n21095), .ZN(n15304) );
  OAI211_X1 U19002 ( .C1(n15306), .C2(n15511), .A(n15305), .B(n15304), .ZN(
        P1_U2970) );
  NAND2_X1 U19003 ( .A1(n10056), .A2(n15548), .ZN(n15318) );
  NAND3_X1 U19004 ( .A1(n15346), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        n15318), .ZN(n15307) );
  OAI21_X1 U19005 ( .B1(n15317), .B2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n15307), .ZN(n15310) );
  MUX2_X1 U19006 ( .A(n15308), .B(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .S(
        n10056), .Z(n15309) );
  NAND2_X1 U19007 ( .A1(n15310), .A2(n15309), .ZN(n15311) );
  XOR2_X1 U19008 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n15311), .Z(
        n15538) );
  NAND2_X1 U19009 ( .A1(n15312), .A2(n15507), .ZN(n15313) );
  NAND2_X1 U19010 ( .A1(n15496), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n15529) );
  OAI211_X1 U19011 ( .C1(n15504), .C2(n21683), .A(n15313), .B(n15529), .ZN(
        n15314) );
  AOI21_X1 U19012 ( .B1(n15315), .B2(n21094), .A(n15314), .ZN(n15316) );
  OAI21_X1 U19013 ( .B1(n20943), .B2(n15538), .A(n15316), .ZN(P1_U2971) );
  OAI21_X1 U19014 ( .B1(n15335), .B2(n15394), .A(n15317), .ZN(n15319) );
  NAND2_X1 U19015 ( .A1(n15319), .A2(n15318), .ZN(n15320) );
  XOR2_X1 U19016 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B(n15320), .Z(
        n15556) );
  NAND2_X1 U19017 ( .A1(n15496), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n15549) );
  OAI21_X1 U19018 ( .B1(n15504), .B2(n15321), .A(n15549), .ZN(n15323) );
  OAI21_X1 U19019 ( .B1(n20943), .B2(n15556), .A(n15325), .ZN(P1_U2973) );
  NOR3_X1 U19020 ( .A1(n9693), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15328) );
  NAND2_X1 U19021 ( .A1(n15326), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15336) );
  NOR2_X1 U19022 ( .A1(n15336), .A2(n15572), .ZN(n15327) );
  MUX2_X1 U19023 ( .A(n15328), .B(n15327), .S(n10056), .Z(n15329) );
  XNOR2_X1 U19024 ( .A(n15329), .B(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15565) );
  NAND2_X1 U19025 ( .A1(n15496), .A2(P1_REIP_REG_25__SCAN_IN), .ZN(n15559) );
  NAND2_X1 U19026 ( .A1(n21088), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15330) );
  OAI211_X1 U19027 ( .C1(n15331), .C2(n21098), .A(n15559), .B(n15330), .ZN(
        n15332) );
  AOI21_X1 U19028 ( .B1(n15333), .B2(n21094), .A(n15332), .ZN(n15334) );
  OAI21_X1 U19029 ( .B1(n20943), .B2(n15565), .A(n15334), .ZN(P1_U2974) );
  NAND2_X1 U19030 ( .A1(n15337), .A2(n15507), .ZN(n15338) );
  NAND2_X1 U19031 ( .A1(n15496), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n15571) );
  OAI211_X1 U19032 ( .C1(n15504), .C2(n15339), .A(n15338), .B(n15571), .ZN(
        n15340) );
  AOI21_X1 U19033 ( .B1(n15341), .B2(n21094), .A(n15340), .ZN(n15342) );
  OAI21_X1 U19034 ( .B1(n20943), .B2(n15577), .A(n15342), .ZN(P1_U2975) );
  AND2_X1 U19035 ( .A1(n15496), .A2(P1_REIP_REG_23__SCAN_IN), .ZN(n15581) );
  NOR2_X1 U19036 ( .A1(n15343), .A2(n21098), .ZN(n15344) );
  AOI211_X1 U19037 ( .C1(n21088), .C2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n15581), .B(n15344), .ZN(n15348) );
  XNOR2_X1 U19038 ( .A(n15394), .B(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15345) );
  XNOR2_X1 U19039 ( .A(n9693), .B(n15345), .ZN(n15578) );
  NAND2_X1 U19040 ( .A1(n15578), .A2(n21095), .ZN(n15347) );
  OAI211_X1 U19041 ( .C1(n15349), .C2(n15511), .A(n15348), .B(n15347), .ZN(
        P1_U2976) );
  NAND2_X1 U19042 ( .A1(n15351), .A2(n15350), .ZN(n15352) );
  XOR2_X1 U19043 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n15352), .Z(
        n15602) );
  NAND2_X1 U19044 ( .A1(n15496), .A2(P1_REIP_REG_22__SCAN_IN), .ZN(n15596) );
  OAI21_X1 U19045 ( .B1(n15504), .B2(n15353), .A(n15596), .ZN(n15356) );
  NOR2_X1 U19046 ( .A1(n15354), .A2(n15511), .ZN(n15355) );
  AOI211_X1 U19047 ( .C1(n15507), .C2(n15357), .A(n15356), .B(n15355), .ZN(
        n15358) );
  OAI21_X1 U19048 ( .B1(n20943), .B2(n15602), .A(n15358), .ZN(P1_U2977) );
  NOR2_X1 U19049 ( .A1(n15359), .A2(n10056), .ZN(n15367) );
  INV_X1 U19050 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n21743) );
  NOR3_X1 U19051 ( .A1(n15360), .A2(n15394), .A3(n21743), .ZN(n15368) );
  MUX2_X1 U19052 ( .A(n15367), .B(n15368), .S(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .Z(n15361) );
  XNOR2_X1 U19053 ( .A(n15361), .B(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15610) );
  NAND2_X1 U19054 ( .A1(n15496), .A2(P1_REIP_REG_21__SCAN_IN), .ZN(n15604) );
  NAND2_X1 U19055 ( .A1(n21088), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15362) );
  OAI211_X1 U19056 ( .C1(n15363), .C2(n21098), .A(n15604), .B(n15362), .ZN(
        n15364) );
  AOI21_X1 U19057 ( .B1(n15365), .B2(n21094), .A(n15364), .ZN(n15366) );
  OAI21_X1 U19058 ( .B1(n15610), .B2(n20943), .A(n15366), .ZN(P1_U2978) );
  NOR2_X1 U19059 ( .A1(n15368), .A2(n15367), .ZN(n15369) );
  XOR2_X1 U19060 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .B(n15369), .Z(
        n15624) );
  NAND2_X1 U19061 ( .A1(n15496), .A2(P1_REIP_REG_20__SCAN_IN), .ZN(n15616) );
  OAI21_X1 U19062 ( .B1(n15504), .B2(n15370), .A(n15616), .ZN(n15373) );
  NOR2_X1 U19063 ( .A1(n15371), .A2(n15511), .ZN(n15372) );
  AOI211_X1 U19064 ( .C1(n15507), .C2(n15374), .A(n15373), .B(n15372), .ZN(
        n15375) );
  OAI21_X1 U19065 ( .B1(n15624), .B2(n20943), .A(n15375), .ZN(P1_U2979) );
  NAND2_X1 U19066 ( .A1(n15360), .A2(n15637), .ZN(n15376) );
  MUX2_X1 U19067 ( .A(n15360), .B(n15376), .S(n15394), .Z(n15377) );
  XOR2_X1 U19068 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B(n15377), .Z(
        n15633) );
  NAND2_X1 U19069 ( .A1(n15496), .A2(P1_REIP_REG_19__SCAN_IN), .ZN(n15626) );
  OAI21_X1 U19070 ( .B1(n15504), .B2(n15378), .A(n15626), .ZN(n15381) );
  NOR2_X1 U19071 ( .A1(n15379), .A2(n15511), .ZN(n15380) );
  AOI211_X1 U19072 ( .C1(n15507), .C2(n15382), .A(n15381), .B(n15380), .ZN(
        n15383) );
  OAI21_X1 U19073 ( .B1(n15633), .B2(n20943), .A(n15383), .ZN(P1_U2980) );
  OAI21_X1 U19074 ( .B1(n15385), .B2(n15384), .A(n15360), .ZN(n15645) );
  NAND2_X1 U19075 ( .A1(n15507), .A2(n15386), .ZN(n15387) );
  NAND2_X1 U19076 ( .A1(n15496), .A2(P1_REIP_REG_18__SCAN_IN), .ZN(n15638) );
  OAI211_X1 U19077 ( .C1(n15504), .C2(n15388), .A(n15387), .B(n15638), .ZN(
        n15389) );
  AOI21_X1 U19078 ( .B1(n15390), .B2(n21094), .A(n15389), .ZN(n15391) );
  OAI21_X1 U19079 ( .B1(n20943), .B2(n15645), .A(n15391), .ZN(P1_U2981) );
  NAND2_X1 U19080 ( .A1(n15392), .A2(n10637), .ZN(n15425) );
  AOI21_X1 U19081 ( .B1(n15425), .B2(n15404), .A(n15393), .ZN(n15396) );
  NOR2_X1 U19082 ( .A1(n15396), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15395) );
  MUX2_X1 U19083 ( .A(n15396), .B(n15395), .S(n15394), .Z(n15397) );
  XNOR2_X1 U19084 ( .A(n15397), .B(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15655) );
  AND2_X1 U19085 ( .A1(n15496), .A2(P1_REIP_REG_17__SCAN_IN), .ZN(n15649) );
  AOI21_X1 U19086 ( .B1(n21088), .B2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n15649), .ZN(n15398) );
  OAI21_X1 U19087 ( .B1(n15399), .B2(n21098), .A(n15398), .ZN(n15400) );
  AOI21_X1 U19088 ( .B1(n15401), .B2(n21094), .A(n15400), .ZN(n15402) );
  OAI21_X1 U19089 ( .B1(n15655), .B2(n20943), .A(n15402), .ZN(P1_U2982) );
  NOR2_X1 U19090 ( .A1(n15425), .A2(n15403), .ZN(n15416) );
  OAI21_X1 U19091 ( .B1(n15416), .B2(n10049), .A(n15412), .ZN(n15405) );
  XOR2_X1 U19092 ( .A(n15406), .B(n15405), .Z(n15665) );
  NAND2_X1 U19093 ( .A1(n15507), .A2(n15407), .ZN(n15408) );
  NAND2_X1 U19094 ( .A1(n15496), .A2(P1_REIP_REG_16__SCAN_IN), .ZN(n15659) );
  OAI211_X1 U19095 ( .C1(n15504), .C2(n10151), .A(n15408), .B(n15659), .ZN(
        n15409) );
  AOI21_X1 U19096 ( .B1(n15410), .B2(n21094), .A(n15409), .ZN(n15411) );
  OAI21_X1 U19097 ( .B1(n15665), .B2(n20943), .A(n15411), .ZN(P1_U2983) );
  INV_X1 U19098 ( .A(n15412), .ZN(n15413) );
  NOR2_X1 U19099 ( .A1(n15414), .A2(n15413), .ZN(n15418) );
  NOR2_X1 U19100 ( .A1(n15416), .A2(n15415), .ZN(n15417) );
  XOR2_X1 U19101 ( .A(n15418), .B(n15417), .Z(n15673) );
  INV_X1 U19102 ( .A(n15419), .ZN(n15423) );
  NAND2_X1 U19103 ( .A1(n15496), .A2(P1_REIP_REG_15__SCAN_IN), .ZN(n15666) );
  NAND2_X1 U19104 ( .A1(n21088), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15420) );
  OAI211_X1 U19105 ( .C1(n21098), .C2(n15421), .A(n15666), .B(n15420), .ZN(
        n15422) );
  AOI21_X1 U19106 ( .B1(n15423), .B2(n21094), .A(n15422), .ZN(n15424) );
  OAI21_X1 U19107 ( .B1(n15673), .B2(n20943), .A(n15424), .ZN(P1_U2984) );
  OAI21_X1 U19108 ( .B1(n15464), .B2(n15427), .A(n15426), .ZN(n15428) );
  NAND2_X1 U19109 ( .A1(n15428), .A2(n13076), .ZN(n15430) );
  XNOR2_X1 U19110 ( .A(n10056), .B(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15429) );
  XNOR2_X1 U19111 ( .A(n15430), .B(n15429), .ZN(n15680) );
  AND2_X1 U19112 ( .A1(n15496), .A2(P1_REIP_REG_14__SCAN_IN), .ZN(n15674) );
  AOI21_X1 U19113 ( .B1(n21088), .B2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n15674), .ZN(n15431) );
  OAI21_X1 U19114 ( .B1(n15432), .B2(n21098), .A(n15431), .ZN(n15433) );
  AOI21_X1 U19115 ( .B1(n15434), .B2(n21094), .A(n15433), .ZN(n15435) );
  OAI21_X1 U19116 ( .B1(n15680), .B2(n20943), .A(n15435), .ZN(P1_U2985) );
  INV_X1 U19117 ( .A(n15436), .ZN(n15437) );
  AOI21_X1 U19118 ( .B1(n15464), .B2(n15438), .A(n15437), .ZN(n15450) );
  AND2_X1 U19119 ( .A1(n15439), .A2(n15440), .ZN(n15449) );
  NAND2_X1 U19120 ( .A1(n15450), .A2(n15449), .ZN(n15448) );
  NAND2_X1 U19121 ( .A1(n15448), .A2(n15440), .ZN(n15441) );
  XNOR2_X1 U19122 ( .A(n15442), .B(n15441), .ZN(n15688) );
  AND2_X1 U19123 ( .A1(n15496), .A2(P1_REIP_REG_13__SCAN_IN), .ZN(n15681) );
  AOI21_X1 U19124 ( .B1(n21088), .B2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n15681), .ZN(n15443) );
  OAI21_X1 U19125 ( .B1(n15444), .B2(n21098), .A(n15443), .ZN(n15445) );
  AOI21_X1 U19126 ( .B1(n15446), .B2(n21094), .A(n15445), .ZN(n15447) );
  OAI21_X1 U19127 ( .B1(n15688), .B2(n20943), .A(n15447), .ZN(P1_U2986) );
  OAI21_X1 U19128 ( .B1(n15450), .B2(n15449), .A(n15448), .ZN(n15695) );
  NAND2_X1 U19129 ( .A1(n15695), .A2(n21095), .ZN(n15455) );
  NAND2_X1 U19130 ( .A1(n15496), .A2(P1_REIP_REG_12__SCAN_IN), .ZN(n15696) );
  OAI21_X1 U19131 ( .B1(n15504), .B2(n15451), .A(n15696), .ZN(n15452) );
  AOI21_X1 U19132 ( .B1(n15507), .B2(n15453), .A(n15452), .ZN(n15454) );
  OAI211_X1 U19133 ( .C1(n15511), .C2(n15456), .A(n15455), .B(n15454), .ZN(
        P1_U2987) );
  NAND3_X1 U19134 ( .A1(n15464), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        n10056), .ZN(n15457) );
  OR3_X1 U19135 ( .A1(n15392), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        n10056), .ZN(n15467) );
  NAND2_X1 U19136 ( .A1(n15457), .A2(n15467), .ZN(n15458) );
  XNOR2_X1 U19137 ( .A(n15458), .B(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n15712) );
  NAND2_X1 U19138 ( .A1(n15496), .A2(P1_REIP_REG_11__SCAN_IN), .ZN(n15707) );
  NAND2_X1 U19139 ( .A1(n21088), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n15459) );
  OAI211_X1 U19140 ( .C1(n21098), .C2(n15460), .A(n15707), .B(n15459), .ZN(
        n15461) );
  AOI21_X1 U19141 ( .B1(n15462), .B2(n21094), .A(n15461), .ZN(n15463) );
  OAI21_X1 U19142 ( .B1(n15712), .B2(n20943), .A(n15463), .ZN(P1_U2988) );
  NAND2_X1 U19143 ( .A1(n15392), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15466) );
  XNOR2_X1 U19144 ( .A(n15464), .B(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15465) );
  MUX2_X1 U19145 ( .A(n15466), .B(n15465), .S(n10056), .Z(n15468) );
  NAND2_X1 U19146 ( .A1(n15468), .A2(n15467), .ZN(n15713) );
  NAND2_X1 U19147 ( .A1(n15713), .A2(n21095), .ZN(n15472) );
  NAND2_X1 U19148 ( .A1(n15496), .A2(P1_REIP_REG_10__SCAN_IN), .ZN(n15720) );
  OAI21_X1 U19149 ( .B1(n15504), .B2(n10156), .A(n15720), .ZN(n15469) );
  AOI21_X1 U19150 ( .B1(n15507), .B2(n15470), .A(n15469), .ZN(n15471) );
  OAI211_X1 U19151 ( .C1(n15511), .C2(n15473), .A(n15472), .B(n15471), .ZN(
        P1_U2989) );
  AND2_X1 U19152 ( .A1(n15475), .A2(n15474), .ZN(n15478) );
  NAND2_X1 U19153 ( .A1(n10637), .A2(n15476), .ZN(n15477) );
  XNOR2_X1 U19154 ( .A(n15478), .B(n15477), .ZN(n15736) );
  NAND2_X1 U19155 ( .A1(n15496), .A2(P1_REIP_REG_9__SCAN_IN), .ZN(n15730) );
  OR2_X1 U19156 ( .A1(n15504), .A2(n10155), .ZN(n15479) );
  OAI211_X1 U19157 ( .C1(n21098), .C2(n15480), .A(n15730), .B(n15479), .ZN(
        n15481) );
  AOI21_X1 U19158 ( .B1(n15482), .B2(n21094), .A(n15481), .ZN(n15483) );
  OAI21_X1 U19159 ( .B1(n15736), .B2(n20943), .A(n15483), .ZN(P1_U2990) );
  XOR2_X1 U19160 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B(n15485), .Z(
        n15486) );
  XNOR2_X1 U19161 ( .A(n15484), .B(n15486), .ZN(n15755) );
  NAND2_X1 U19162 ( .A1(n15496), .A2(P1_REIP_REG_8__SCAN_IN), .ZN(n15749) );
  NAND2_X1 U19163 ( .A1(n21088), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n15487) );
  OAI211_X1 U19164 ( .C1(n21098), .C2(n15488), .A(n15749), .B(n15487), .ZN(
        n15489) );
  AOI21_X1 U19165 ( .B1(n15490), .B2(n21094), .A(n15489), .ZN(n15491) );
  OAI21_X1 U19166 ( .B1(n15755), .B2(n20943), .A(n15491), .ZN(P1_U2991) );
  NAND2_X1 U19167 ( .A1(n15493), .A2(n15492), .ZN(n15495) );
  XOR2_X1 U19168 ( .A(n15495), .B(n15494), .Z(n15762) );
  NAND2_X1 U19169 ( .A1(n15496), .A2(P1_REIP_REG_7__SCAN_IN), .ZN(n15757) );
  NAND2_X1 U19170 ( .A1(n21088), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15497) );
  OAI211_X1 U19171 ( .C1(n21098), .C2(n20974), .A(n15757), .B(n15497), .ZN(
        n15498) );
  AOI21_X1 U19172 ( .B1(n20971), .B2(n21094), .A(n15498), .ZN(n15499) );
  OAI21_X1 U19173 ( .B1(n15762), .B2(n20943), .A(n15499), .ZN(P1_U2992) );
  XNOR2_X1 U19174 ( .A(n15500), .B(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n15502) );
  NOR2_X1 U19175 ( .A1(n15502), .A2(n9692), .ZN(n21089) );
  AOI21_X1 U19176 ( .B1(n15502), .B2(n9692), .A(n21089), .ZN(n21109) );
  NAND2_X1 U19177 ( .A1(n21109), .A2(n21095), .ZN(n15509) );
  OAI22_X1 U19178 ( .A1(n15504), .A2(n15503), .B1(n21123), .B2(n21545), .ZN(
        n15505) );
  AOI21_X1 U19179 ( .B1(n15507), .B2(n15506), .A(n15505), .ZN(n15508) );
  OAI211_X1 U19180 ( .C1(n15511), .C2(n15510), .A(n15509), .B(n15508), .ZN(
        P1_U2996) );
  NAND3_X1 U19181 ( .A1(n15513), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n15528), .ZN(n15518) );
  NAND3_X1 U19182 ( .A1(n15515), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n15514), .ZN(n15516) );
  NAND2_X1 U19183 ( .A1(n15520), .A2(n21110), .ZN(n15526) );
  INV_X1 U19184 ( .A(n15521), .ZN(n15524) );
  NOR3_X1 U19185 ( .A1(n15540), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n15530), .ZN(n15522) );
  AOI211_X1 U19186 ( .C1(n15524), .C2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n15523), .B(n15522), .ZN(n15525) );
  OAI211_X1 U19187 ( .C1(n15527), .C2(n21125), .A(n15526), .B(n15525), .ZN(
        P1_U3002) );
  AND2_X1 U19188 ( .A1(n15554), .A2(n15528), .ZN(n15544) );
  INV_X1 U19189 ( .A(n15529), .ZN(n15533) );
  NOR3_X1 U19190 ( .A1(n15540), .A2(n13412), .A3(n15531), .ZN(n15532) );
  AOI211_X1 U19191 ( .C1(n15544), .C2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n15533), .B(n15532), .ZN(n15537) );
  INV_X1 U19192 ( .A(n15534), .ZN(n15535) );
  NAND2_X1 U19193 ( .A1(n15535), .A2(n21135), .ZN(n15536) );
  OAI211_X1 U19194 ( .C1(n15538), .C2(n21139), .A(n15537), .B(n15536), .ZN(
        P1_U3003) );
  OAI21_X1 U19195 ( .B1(n15540), .B2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n15539), .ZN(n15543) );
  NOR2_X1 U19196 ( .A1(n15541), .A2(n21125), .ZN(n15542) );
  AOI211_X1 U19197 ( .C1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n15544), .A(
        n15543), .B(n15542), .ZN(n15545) );
  OAI21_X1 U19198 ( .B1(n15569), .B2(n15548), .A(n15547), .ZN(n15553) );
  INV_X1 U19199 ( .A(n15549), .ZN(n15552) );
  NOR2_X1 U19200 ( .A1(n15550), .A2(n21125), .ZN(n15551) );
  AOI211_X1 U19201 ( .C1(n15554), .C2(n15553), .A(n15552), .B(n15551), .ZN(
        n15555) );
  OAI21_X1 U19202 ( .B1(n15556), .B2(n21139), .A(n15555), .ZN(P1_U3005) );
  NOR2_X1 U19203 ( .A1(n15557), .A2(n15558), .ZN(n15562) );
  NAND3_X1 U19204 ( .A1(n15558), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15560) );
  OAI21_X1 U19205 ( .B1(n15569), .B2(n15560), .A(n15559), .ZN(n15561) );
  AOI211_X1 U19206 ( .C1(n15563), .C2(n21135), .A(n15562), .B(n15561), .ZN(
        n15564) );
  OAI21_X1 U19207 ( .B1(n15565), .B2(n21139), .A(n15564), .ZN(P1_U3006) );
  NOR2_X1 U19208 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n15566), .ZN(
        n15568) );
  NOR2_X1 U19209 ( .A1(n15568), .A2(n15567), .ZN(n15573) );
  INV_X1 U19210 ( .A(n15569), .ZN(n15583) );
  NAND3_X1 U19211 ( .A1(n15583), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        n15572), .ZN(n15570) );
  OAI211_X1 U19212 ( .C1(n15573), .C2(n15572), .A(n15571), .B(n15570), .ZN(
        n15574) );
  AOI21_X1 U19213 ( .B1(n15575), .B2(n21135), .A(n15574), .ZN(n15576) );
  OAI21_X1 U19214 ( .B1(n15577), .B2(n21139), .A(n15576), .ZN(P1_U3007) );
  NAND2_X1 U19215 ( .A1(n15578), .A2(n21110), .ZN(n15585) );
  INV_X1 U19216 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15582) );
  NOR2_X1 U19217 ( .A1(n15579), .A2(n15582), .ZN(n15580) );
  AOI211_X1 U19218 ( .C1(n15583), .C2(n15582), .A(n15581), .B(n15580), .ZN(
        n15584) );
  OAI211_X1 U19219 ( .C1(n15586), .C2(n21125), .A(n15585), .B(n15584), .ZN(
        P1_U3008) );
  INV_X1 U19220 ( .A(n15587), .ZN(n15588) );
  OR2_X1 U19221 ( .A1(n21117), .A2(n15588), .ZN(n15591) );
  OR3_X1 U19222 ( .A1(n21118), .A2(n15589), .A3(n15592), .ZN(n15590) );
  NAND2_X1 U19223 ( .A1(n15591), .A2(n15590), .ZN(n15613) );
  NOR2_X1 U19224 ( .A1(n15611), .A2(n15592), .ZN(n15593) );
  NOR2_X1 U19225 ( .A1(n15613), .A2(n15593), .ZN(n15684) );
  NOR3_X1 U19226 ( .A1(n15684), .A2(n15594), .A3(n15683), .ZN(n15617) );
  NAND2_X1 U19227 ( .A1(n15617), .A2(n15595), .ZN(n15606) );
  XNOR2_X1 U19228 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .B(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15597) );
  OAI21_X1 U19229 ( .B1(n15606), .B2(n15597), .A(n15596), .ZN(n15600) );
  NOR2_X1 U19230 ( .A1(n15598), .A2(n21125), .ZN(n15599) );
  AOI211_X1 U19231 ( .C1(n15603), .C2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n15600), .B(n15599), .ZN(n15601) );
  OAI21_X1 U19232 ( .B1(n15602), .B2(n21139), .A(n15601), .ZN(P1_U3009) );
  NAND2_X1 U19233 ( .A1(n15603), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15605) );
  OAI211_X1 U19234 ( .C1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n15606), .A(
        n15605), .B(n15604), .ZN(n15607) );
  AOI21_X1 U19235 ( .B1(n15608), .B2(n21135), .A(n15607), .ZN(n15609) );
  OAI21_X1 U19236 ( .B1(n15610), .B2(n21139), .A(n15609), .ZN(P1_U3010) );
  INV_X1 U19237 ( .A(n15656), .ZN(n15685) );
  INV_X1 U19238 ( .A(n15611), .ZN(n15612) );
  OAI21_X1 U19239 ( .B1(n15613), .B2(n15612), .A(n21743), .ZN(n15615) );
  NAND3_X1 U19240 ( .A1(n15685), .A2(n15615), .A3(n15614), .ZN(n15620) );
  INV_X1 U19241 ( .A(n15616), .ZN(n15619) );
  INV_X1 U19242 ( .A(n15617), .ZN(n15628) );
  NOR3_X1 U19243 ( .A1(n15628), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A3(
        n21743), .ZN(n15618) );
  AOI211_X1 U19244 ( .C1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .C2(n15620), .A(
        n15619), .B(n15618), .ZN(n15623) );
  NAND2_X1 U19245 ( .A1(n15621), .A2(n21135), .ZN(n15622) );
  OAI211_X1 U19246 ( .C1(n15624), .C2(n21139), .A(n15623), .B(n15622), .ZN(
        P1_U3011) );
  INV_X1 U19247 ( .A(n15625), .ZN(n15631) );
  INV_X1 U19248 ( .A(n15626), .ZN(n15630) );
  AOI21_X1 U19249 ( .B1(n15628), .B2(n21743), .A(n15627), .ZN(n15629) );
  AOI211_X1 U19250 ( .C1(n15631), .C2(n21135), .A(n15630), .B(n15629), .ZN(
        n15632) );
  OAI21_X1 U19251 ( .B1(n15633), .B2(n21139), .A(n15632), .ZN(P1_U3012) );
  NAND2_X1 U19252 ( .A1(n21137), .A2(n15635), .ZN(n15634) );
  NAND2_X1 U19253 ( .A1(n15685), .A2(n15634), .ZN(n15651) );
  INV_X1 U19254 ( .A(n15635), .ZN(n15636) );
  NAND3_X1 U19255 ( .A1(n15676), .A2(n15637), .A3(n15636), .ZN(n15639) );
  NAND2_X1 U19256 ( .A1(n15639), .A2(n15638), .ZN(n15640) );
  AOI21_X1 U19257 ( .B1(n15651), .B2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n15640), .ZN(n15644) );
  INV_X1 U19258 ( .A(n15641), .ZN(n15642) );
  NAND2_X1 U19259 ( .A1(n15642), .A2(n21135), .ZN(n15643) );
  OAI211_X1 U19260 ( .C1(n15645), .C2(n21139), .A(n15644), .B(n15643), .ZN(
        P1_U3013) );
  INV_X1 U19261 ( .A(n15676), .ZN(n15648) );
  NAND3_X1 U19262 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15647) );
  OAI21_X1 U19263 ( .B1(n15648), .B2(n15647), .A(n15646), .ZN(n15650) );
  AOI21_X1 U19264 ( .B1(n15651), .B2(n15650), .A(n15649), .ZN(n15654) );
  NAND2_X1 U19265 ( .A1(n15652), .A2(n21135), .ZN(n15653) );
  OAI211_X1 U19266 ( .C1(n15655), .C2(n21139), .A(n15654), .B(n15653), .ZN(
        P1_U3014) );
  AOI21_X1 U19267 ( .B1(n15677), .B2(n21137), .A(n15656), .ZN(n15669) );
  NOR2_X1 U19268 ( .A1(n15677), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15657) );
  NAND2_X1 U19269 ( .A1(n15676), .A2(n15657), .ZN(n15667) );
  AOI21_X1 U19270 ( .B1(n15669), .B2(n15667), .A(n15658), .ZN(n15662) );
  NAND4_X1 U19271 ( .A1(n15676), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A4(n15658), .ZN(n15660) );
  NAND2_X1 U19272 ( .A1(n15660), .A2(n15659), .ZN(n15661) );
  AOI211_X1 U19273 ( .C1(n15663), .C2(n21135), .A(n15662), .B(n15661), .ZN(
        n15664) );
  OAI21_X1 U19274 ( .B1(n15665), .B2(n21139), .A(n15664), .ZN(P1_U3015) );
  OAI211_X1 U19275 ( .C1(n15669), .C2(n15668), .A(n15667), .B(n15666), .ZN(
        n15670) );
  AOI21_X1 U19276 ( .B1(n15671), .B2(n21135), .A(n15670), .ZN(n15672) );
  OAI21_X1 U19277 ( .B1(n15673), .B2(n21139), .A(n15672), .ZN(P1_U3016) );
  AOI21_X1 U19278 ( .B1(n15675), .B2(n21135), .A(n15674), .ZN(n15679) );
  MUX2_X1 U19279 ( .A(n15685), .B(n15648), .S(n15677), .Z(n15678) );
  OAI211_X1 U19280 ( .C1(n15680), .C2(n21139), .A(n15679), .B(n15678), .ZN(
        P1_U3017) );
  AOI21_X1 U19281 ( .B1(n15682), .B2(n21135), .A(n15681), .ZN(n15687) );
  MUX2_X1 U19282 ( .A(n15685), .B(n15684), .S(n15683), .Z(n15686) );
  OAI211_X1 U19283 ( .C1(n15688), .C2(n21139), .A(n15687), .B(n15686), .ZN(
        P1_U3018) );
  INV_X1 U19284 ( .A(n21119), .ZN(n15691) );
  INV_X1 U19285 ( .A(n15689), .ZN(n15698) );
  OAI21_X1 U19286 ( .B1(n15698), .B2(n15738), .A(n15739), .ZN(n15690) );
  OAI211_X1 U19287 ( .C1(n15742), .C2(n15692), .A(n15691), .B(n15690), .ZN(
        n15710) );
  AOI21_X1 U19288 ( .B1(n15694), .B2(n15693), .A(n15710), .ZN(n15704) );
  NAND2_X1 U19289 ( .A1(n15695), .A2(n21110), .ZN(n15703) );
  INV_X1 U19290 ( .A(n15696), .ZN(n15700) );
  NOR2_X1 U19291 ( .A1(n21101), .A2(n21116), .ZN(n15744) );
  INV_X1 U19292 ( .A(n15744), .ZN(n15697) );
  NAND2_X1 U19293 ( .A1(n21117), .A2(n15697), .ZN(n18036) );
  INV_X1 U19294 ( .A(n15738), .ZN(n15714) );
  NAND2_X1 U19295 ( .A1(n18036), .A2(n15714), .ZN(n15746) );
  NOR3_X1 U19296 ( .A1(n15746), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A3(
        n15698), .ZN(n15699) );
  AOI211_X1 U19297 ( .C1(n15701), .C2(n21135), .A(n15700), .B(n15699), .ZN(
        n15702) );
  OAI211_X1 U19298 ( .C1(n15704), .C2(n21804), .A(n15703), .B(n15702), .ZN(
        P1_U3019) );
  OR3_X1 U19299 ( .A1(n15746), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(
        n15705), .ZN(n15706) );
  OAI211_X1 U19300 ( .C1(n15708), .C2(n21125), .A(n15707), .B(n15706), .ZN(
        n15709) );
  AOI21_X1 U19301 ( .B1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n15710), .A(
        n15709), .ZN(n15711) );
  OAI21_X1 U19302 ( .B1(n15712), .B2(n21139), .A(n15711), .ZN(P1_U3020) );
  INV_X1 U19303 ( .A(n15713), .ZN(n15728) );
  NAND2_X1 U19304 ( .A1(n15742), .A2(n15714), .ZN(n15716) );
  INV_X1 U19305 ( .A(n15722), .ZN(n15715) );
  AOI211_X1 U19306 ( .C1(n15717), .C2(n15716), .A(n15715), .B(n21119), .ZN(
        n15719) );
  NOR2_X1 U19307 ( .A1(n15719), .A2(n15718), .ZN(n15734) );
  OAI21_X1 U19308 ( .B1(n15721), .B2(n21125), .A(n15720), .ZN(n15726) );
  INV_X1 U19309 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15724) );
  INV_X1 U19310 ( .A(n15746), .ZN(n18030) );
  NAND2_X1 U19311 ( .A1(n18030), .A2(n15722), .ZN(n15729) );
  AOI211_X1 U19312 ( .C1(n21728), .C2(n15724), .A(n15723), .B(n15729), .ZN(
        n15725) );
  AOI211_X1 U19313 ( .C1(n15734), .C2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n15726), .B(n15725), .ZN(n15727) );
  OAI21_X1 U19314 ( .B1(n15728), .B2(n21139), .A(n15727), .ZN(P1_U3021) );
  NOR2_X1 U19315 ( .A1(n15729), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15733) );
  OAI21_X1 U19316 ( .B1(n15731), .B2(n21125), .A(n15730), .ZN(n15732) );
  AOI211_X1 U19317 ( .C1(n15734), .C2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n15733), .B(n15732), .ZN(n15735) );
  OAI21_X1 U19318 ( .B1(n15736), .B2(n21139), .A(n15735), .ZN(P1_U3022) );
  NAND2_X1 U19319 ( .A1(n15737), .A2(n21104), .ZN(n18042) );
  INV_X1 U19320 ( .A(n18042), .ZN(n15743) );
  AOI21_X1 U19321 ( .B1(n15739), .B2(n15738), .A(n21119), .ZN(n15740) );
  OAI21_X1 U19322 ( .B1(n15742), .B2(n15741), .A(n15740), .ZN(n18038) );
  AOI21_X1 U19323 ( .B1(n15744), .B2(n15743), .A(n18038), .ZN(n18035) );
  INV_X1 U19324 ( .A(n18035), .ZN(n15745) );
  AOI21_X1 U19325 ( .B1(n18034), .B2(n21137), .A(n15745), .ZN(n15756) );
  OR3_X1 U19326 ( .A1(n15746), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(
        n18034), .ZN(n15758) );
  NAND2_X1 U19327 ( .A1(n15756), .A2(n15758), .ZN(n15753) );
  INV_X1 U19328 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n15747) );
  NAND3_X1 U19329 ( .A1(n18030), .A2(n15748), .A3(n15747), .ZN(n15750) );
  OAI211_X1 U19330 ( .C1(n21125), .C2(n15751), .A(n15750), .B(n15749), .ZN(
        n15752) );
  AOI21_X1 U19331 ( .B1(n15753), .B2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A(
        n15752), .ZN(n15754) );
  OAI21_X1 U19332 ( .B1(n21139), .B2(n15755), .A(n15754), .ZN(P1_U3023) );
  INV_X1 U19333 ( .A(n15756), .ZN(n15760) );
  OAI211_X1 U19334 ( .C1(n20962), .C2(n21125), .A(n15758), .B(n15757), .ZN(
        n15759) );
  AOI21_X1 U19335 ( .B1(n15760), .B2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n15759), .ZN(n15761) );
  OAI21_X1 U19336 ( .B1(n15762), .B2(n21139), .A(n15761), .ZN(P1_U3024) );
  AND2_X1 U19337 ( .A1(n15764), .A2(n15763), .ZN(n15765) );
  NAND2_X1 U19338 ( .A1(n15766), .A2(n15765), .ZN(n15968) );
  NAND2_X1 U19339 ( .A1(n15936), .A2(n15769), .ZN(n15767) );
  OAI211_X1 U19340 ( .C1(n21417), .C2(n14364), .A(n15968), .B(n15767), .ZN(
        n15768) );
  MUX2_X1 U19341 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n15768), .S(
        n21146), .Z(P1_U3478) );
  INV_X1 U19342 ( .A(n15769), .ZN(n15773) );
  NAND2_X1 U19343 ( .A1(n21468), .A2(n21376), .ZN(n21377) );
  MUX2_X1 U19344 ( .A(n21420), .B(n21377), .S(n14363), .Z(n15770) );
  OAI21_X1 U19345 ( .B1(n15773), .B2(n13944), .A(n15770), .ZN(n15771) );
  MUX2_X1 U19346 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n15771), .S(
        n21146), .Z(P1_U3477) );
  AOI211_X1 U19347 ( .C1(n14363), .C2(n21268), .A(n21419), .B(n15848), .ZN(
        n15772) );
  OAI222_X1 U19348 ( .A1(n14524), .A2(n21377), .B1(n15774), .B2(n15773), .C1(
        n21420), .C2(n15772), .ZN(n15775) );
  MUX2_X1 U19349 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n15775), .S(
        n21146), .Z(P1_U3475) );
  INV_X1 U19350 ( .A(n21594), .ZN(n15779) );
  INV_X1 U19351 ( .A(n15776), .ZN(n21596) );
  AOI22_X1 U19352 ( .A1(n15779), .A2(n15778), .B1(n15777), .B2(n21596), .ZN(
        n15780) );
  OAI21_X1 U19353 ( .B1(n15781), .B2(n21602), .A(n15780), .ZN(n15782) );
  MUX2_X1 U19354 ( .A(n15783), .B(n15782), .S(n21597), .Z(P1_U3472) );
  INV_X1 U19355 ( .A(n15784), .ZN(n15785) );
  OAI22_X1 U19356 ( .A1(n15786), .A2(n21602), .B1(n15785), .B2(n21594), .ZN(
        n15787) );
  MUX2_X1 U19357 ( .A(n15788), .B(n15787), .S(n21597), .Z(P1_U3469) );
  INV_X1 U19358 ( .A(n9709), .ZN(n15789) );
  OAI21_X1 U19359 ( .B1(n21169), .B2(n15790), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n15791) );
  NAND2_X1 U19360 ( .A1(n15791), .A2(n21376), .ZN(n15804) );
  INV_X1 U19361 ( .A(n15804), .ZN(n15799) );
  OR2_X1 U19362 ( .A1(n14439), .A2(n15792), .ZN(n21237) );
  INV_X1 U19363 ( .A(n21237), .ZN(n21175) );
  NAND2_X1 U19364 ( .A1(n21175), .A2(n13944), .ZN(n15803) );
  NAND2_X1 U19365 ( .A1(n15945), .A2(n15793), .ZN(n21240) );
  NOR2_X1 U19366 ( .A1(n15898), .A2(n21240), .ZN(n15800) );
  INV_X1 U19367 ( .A(n15852), .ZN(n15794) );
  INV_X1 U19368 ( .A(n21380), .ZN(n15851) );
  NAND2_X1 U19369 ( .A1(n15794), .A2(n15851), .ZN(n15813) );
  NAND2_X1 U19370 ( .A1(n15813), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15797) );
  INV_X1 U19371 ( .A(n15802), .ZN(n15795) );
  NOR2_X1 U19372 ( .A1(n15795), .A2(n21349), .ZN(n21460) );
  OAI211_X1 U19373 ( .C1(n15800), .C2(n21719), .A(n15797), .B(n21386), .ZN(
        n15798) );
  INV_X1 U19374 ( .A(n15800), .ZN(n21166) );
  OAI22_X1 U19375 ( .A1(n21167), .A2(n21480), .B1(n21166), .B2(n21303), .ZN(
        n15801) );
  AOI21_X1 U19376 ( .B1(n21169), .B2(n21477), .A(n15801), .ZN(n15806) );
  OR2_X1 U19377 ( .A1(n15802), .A2(n21349), .ZN(n15853) );
  INV_X1 U19378 ( .A(n21394), .ZN(n21466) );
  NAND2_X1 U19379 ( .A1(n21170), .A2(n21466), .ZN(n15805) );
  OAI211_X1 U19380 ( .C1(n21173), .C2(n15807), .A(n15806), .B(n15805), .ZN(
        P1_U3033) );
  INV_X1 U19381 ( .A(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n15811) );
  OAI22_X1 U19382 ( .A1(n21167), .A2(n21514), .B1(n21166), .B2(n21333), .ZN(
        n15808) );
  AOI21_X1 U19383 ( .B1(n21169), .B2(n21511), .A(n15808), .ZN(n15810) );
  INV_X1 U19384 ( .A(n21409), .ZN(n21510) );
  NAND2_X1 U19385 ( .A1(n21170), .A2(n21510), .ZN(n15809) );
  OAI211_X1 U19386 ( .C1(n21173), .C2(n15811), .A(n15810), .B(n15809), .ZN(
        P1_U3039) );
  INV_X1 U19387 ( .A(n15813), .ZN(n15815) );
  NOR3_X1 U19388 ( .A1(n21298), .A2(n21471), .A3(n21417), .ZN(n15814) );
  AOI21_X1 U19389 ( .B1(n21460), .B2(n15815), .A(n15814), .ZN(n15843) );
  OAI21_X1 U19390 ( .B1(n21261), .B2(n21292), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n15817) );
  NAND2_X1 U19391 ( .A1(n21270), .A2(n13944), .ZN(n15816) );
  AOI21_X1 U19392 ( .B1(n15817), .B2(n15816), .A(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n15819) );
  AND2_X1 U19393 ( .A1(n15853), .A2(n15818), .ZN(n21473) );
  AOI22_X1 U19394 ( .A1(n21465), .A2(n9850), .B1(
        P1_INSTQUEUE_REG_4__0__SCAN_IN), .B2(n15841), .ZN(n15820) );
  OAI21_X1 U19395 ( .B1(n15843), .B2(n21394), .A(n15820), .ZN(n15821) );
  AOI21_X1 U19396 ( .B1(n21292), .B2(n21477), .A(n15821), .ZN(n15822) );
  OAI21_X1 U19397 ( .B1(n21480), .B2(n15846), .A(n15822), .ZN(P1_U3065) );
  AOI22_X1 U19398 ( .A1(n21481), .A2(n9850), .B1(
        P1_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n15841), .ZN(n15823) );
  OAI21_X1 U19399 ( .B1(n15843), .B2(n21397), .A(n15823), .ZN(n15824) );
  AOI21_X1 U19400 ( .B1(n21292), .B2(n21483), .A(n15824), .ZN(n15825) );
  OAI21_X1 U19401 ( .B1(n21486), .B2(n15846), .A(n15825), .ZN(P1_U3066) );
  AOI22_X1 U19402 ( .A1(n21928), .A2(n9850), .B1(
        P1_INSTQUEUE_REG_4__2__SCAN_IN), .B2(n15841), .ZN(n15826) );
  OAI21_X1 U19403 ( .B1(n15843), .B2(n21936), .A(n15826), .ZN(n15827) );
  AOI21_X1 U19404 ( .B1(n21292), .B2(n21931), .A(n15827), .ZN(n15828) );
  OAI21_X1 U19405 ( .B1(n21490), .B2(n15846), .A(n15828), .ZN(P1_U3067) );
  AOI22_X1 U19406 ( .A1(n21491), .A2(n9850), .B1(
        P1_INSTQUEUE_REG_4__3__SCAN_IN), .B2(n15841), .ZN(n15829) );
  OAI21_X1 U19407 ( .B1(n15843), .B2(n21400), .A(n15829), .ZN(n15830) );
  AOI21_X1 U19408 ( .B1(n21292), .B2(n21493), .A(n15830), .ZN(n15831) );
  OAI21_X1 U19409 ( .B1(n21496), .B2(n15846), .A(n15831), .ZN(P1_U3068) );
  AOI22_X1 U19410 ( .A1(n21497), .A2(n9850), .B1(
        P1_INSTQUEUE_REG_4__4__SCAN_IN), .B2(n15841), .ZN(n15832) );
  OAI21_X1 U19411 ( .B1(n15843), .B2(n21403), .A(n15832), .ZN(n15833) );
  AOI21_X1 U19412 ( .B1(n21292), .B2(n21499), .A(n15833), .ZN(n15834) );
  OAI21_X1 U19413 ( .B1(n21502), .B2(n15846), .A(n15834), .ZN(P1_U3069) );
  AOI22_X1 U19414 ( .A1(n21503), .A2(n9850), .B1(
        P1_INSTQUEUE_REG_4__5__SCAN_IN), .B2(n15841), .ZN(n15835) );
  OAI21_X1 U19415 ( .B1(n15843), .B2(n21406), .A(n15835), .ZN(n15836) );
  AOI21_X1 U19416 ( .B1(n21292), .B2(n21505), .A(n15836), .ZN(n15837) );
  OAI21_X1 U19417 ( .B1(n21508), .B2(n15846), .A(n15837), .ZN(P1_U3070) );
  AOI22_X1 U19418 ( .A1(n21509), .A2(n9850), .B1(
        P1_INSTQUEUE_REG_4__6__SCAN_IN), .B2(n15841), .ZN(n15838) );
  OAI21_X1 U19419 ( .B1(n15843), .B2(n21409), .A(n15838), .ZN(n15839) );
  AOI21_X1 U19420 ( .B1(n21292), .B2(n21511), .A(n15839), .ZN(n15840) );
  OAI21_X1 U19421 ( .B1(n21514), .B2(n15846), .A(n15840), .ZN(P1_U3071) );
  AOI22_X1 U19422 ( .A1(n21516), .A2(n9850), .B1(
        P1_INSTQUEUE_REG_4__7__SCAN_IN), .B2(n15841), .ZN(n15842) );
  OAI21_X1 U19423 ( .B1(n15843), .B2(n21412), .A(n15842), .ZN(n15844) );
  AOI21_X1 U19424 ( .B1(n21292), .B2(n21519), .A(n15844), .ZN(n15845) );
  OAI21_X1 U19425 ( .B1(n21525), .B2(n15846), .A(n15845), .ZN(P1_U3072) );
  OR2_X1 U19426 ( .A1(n21379), .A2(n21471), .ZN(n15849) );
  OR2_X1 U19427 ( .A1(n15898), .A2(n21346), .ZN(n15863) );
  INV_X1 U19428 ( .A(n15857), .ZN(n15850) );
  NAND2_X1 U19429 ( .A1(n15850), .A2(n21376), .ZN(n15855) );
  AND2_X1 U19430 ( .A1(n15852), .A2(n15851), .ZN(n15899) );
  INV_X1 U19431 ( .A(n15853), .ZN(n21382) );
  NAND2_X1 U19432 ( .A1(n15899), .A2(n21382), .ZN(n15854) );
  INV_X1 U19433 ( .A(n15863), .ZN(n15888) );
  OAI21_X1 U19434 ( .B1(n15889), .B2(n15894), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n15856) );
  NAND2_X1 U19435 ( .A1(n15857), .A2(n15856), .ZN(n15858) );
  OAI211_X1 U19436 ( .C1(n15888), .C2(n21719), .A(n21386), .B(n15858), .ZN(
        n15887) );
  AOI22_X1 U19437 ( .A1(n21465), .A2(n15888), .B1(
        P1_INSTQUEUE_REG_8__0__SCAN_IN), .B2(n15887), .ZN(n15859) );
  OAI21_X1 U19438 ( .B1(n15892), .B2(n21394), .A(n15859), .ZN(n15860) );
  AOI21_X1 U19439 ( .B1(n15889), .B2(n21425), .A(n15860), .ZN(n15861) );
  OAI21_X1 U19440 ( .B1(n21428), .B2(n21375), .A(n15861), .ZN(P1_U3097) );
  INV_X1 U19441 ( .A(n15892), .ZN(n15865) );
  INV_X1 U19442 ( .A(n15887), .ZN(n15862) );
  OAI22_X1 U19443 ( .A1(n21313), .A2(n15863), .B1(n21759), .B2(n15862), .ZN(
        n15864) );
  AOI21_X1 U19444 ( .B1(n15865), .B2(n21482), .A(n15864), .ZN(n15867) );
  NAND2_X1 U19445 ( .A1(n15889), .A2(n21429), .ZN(n15866) );
  OAI211_X1 U19446 ( .C1(n21432), .C2(n21375), .A(n15867), .B(n15866), .ZN(
        P1_U3098) );
  AOI22_X1 U19447 ( .A1(n21928), .A2(n15888), .B1(
        P1_INSTQUEUE_REG_8__2__SCAN_IN), .B2(n15887), .ZN(n15869) );
  NAND2_X1 U19448 ( .A1(n15889), .A2(n21929), .ZN(n15868) );
  OAI211_X1 U19449 ( .C1(n15892), .C2(n21936), .A(n15869), .B(n15868), .ZN(
        n15870) );
  AOI21_X1 U19450 ( .B1(n15894), .B2(n21931), .A(n15870), .ZN(n15871) );
  INV_X1 U19451 ( .A(n15871), .ZN(P1_U3099) );
  AOI22_X1 U19452 ( .A1(n21491), .A2(n15888), .B1(
        P1_INSTQUEUE_REG_8__3__SCAN_IN), .B2(n15887), .ZN(n15873) );
  NAND2_X1 U19453 ( .A1(n15889), .A2(n21436), .ZN(n15872) );
  OAI211_X1 U19454 ( .C1(n15892), .C2(n21400), .A(n15873), .B(n15872), .ZN(
        n15874) );
  AOI21_X1 U19455 ( .B1(n15894), .B2(n21493), .A(n15874), .ZN(n15875) );
  INV_X1 U19456 ( .A(n15875), .ZN(P1_U3100) );
  AOI22_X1 U19457 ( .A1(n21497), .A2(n15888), .B1(
        P1_INSTQUEUE_REG_8__4__SCAN_IN), .B2(n15887), .ZN(n15877) );
  NAND2_X1 U19458 ( .A1(n15889), .A2(n21440), .ZN(n15876) );
  OAI211_X1 U19459 ( .C1(n15892), .C2(n21403), .A(n15877), .B(n15876), .ZN(
        n15878) );
  AOI21_X1 U19460 ( .B1(n15894), .B2(n21499), .A(n15878), .ZN(n15879) );
  INV_X1 U19461 ( .A(n15879), .ZN(P1_U3101) );
  AOI22_X1 U19462 ( .A1(n21503), .A2(n15888), .B1(
        P1_INSTQUEUE_REG_8__5__SCAN_IN), .B2(n15887), .ZN(n15881) );
  NAND2_X1 U19463 ( .A1(n15889), .A2(n21444), .ZN(n15880) );
  OAI211_X1 U19464 ( .C1(n15892), .C2(n21406), .A(n15881), .B(n15880), .ZN(
        n15882) );
  AOI21_X1 U19465 ( .B1(n15894), .B2(n21505), .A(n15882), .ZN(n15883) );
  INV_X1 U19466 ( .A(n15883), .ZN(P1_U3102) );
  AOI22_X1 U19467 ( .A1(n21509), .A2(n15888), .B1(
        P1_INSTQUEUE_REG_8__6__SCAN_IN), .B2(n15887), .ZN(n15884) );
  OAI21_X1 U19468 ( .B1(n15892), .B2(n21409), .A(n15884), .ZN(n15885) );
  AOI21_X1 U19469 ( .B1(n15889), .B2(n21448), .A(n15885), .ZN(n15886) );
  OAI21_X1 U19470 ( .B1(n21451), .B2(n21375), .A(n15886), .ZN(P1_U3103) );
  AOI22_X1 U19471 ( .A1(n21516), .A2(n15888), .B1(
        P1_INSTQUEUE_REG_8__7__SCAN_IN), .B2(n15887), .ZN(n15891) );
  NAND2_X1 U19472 ( .A1(n15889), .A2(n21454), .ZN(n15890) );
  OAI211_X1 U19473 ( .C1(n15892), .C2(n21412), .A(n15891), .B(n15890), .ZN(
        n15893) );
  AOI21_X1 U19474 ( .B1(n15894), .B2(n21519), .A(n15893), .ZN(n15895) );
  INV_X1 U19475 ( .A(n15895), .ZN(P1_U3104) );
  NAND3_X1 U19476 ( .A1(n15896), .A2(n21376), .A3(n15928), .ZN(n15897) );
  NAND2_X1 U19477 ( .A1(n15897), .A2(n21377), .ZN(n15902) );
  NOR2_X1 U19478 ( .A1(n21467), .A2(n21471), .ZN(n15900) );
  INV_X1 U19479 ( .A(n15899), .ZN(n15903) );
  INV_X1 U19480 ( .A(n15900), .ZN(n15901) );
  AOI22_X1 U19481 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n15903), .B1(n15902), 
        .B2(n15901), .ZN(n15904) );
  OAI211_X1 U19482 ( .C1(n9851), .C2(n21719), .A(n21473), .B(n15904), .ZN(
        n15926) );
  AOI22_X1 U19483 ( .A1(n21465), .A2(n9851), .B1(
        P1_INSTQUEUE_REG_12__0__SCAN_IN), .B2(n15926), .ZN(n15905) );
  OAI21_X1 U19484 ( .B1(n15928), .B2(n21428), .A(n15905), .ZN(n15906) );
  AOI21_X1 U19485 ( .B1(n15930), .B2(n21425), .A(n15906), .ZN(n15907) );
  OAI21_X1 U19486 ( .B1(n15932), .B2(n21394), .A(n15907), .ZN(P1_U3129) );
  AOI22_X1 U19487 ( .A1(n21481), .A2(n9851), .B1(
        P1_INSTQUEUE_REG_12__1__SCAN_IN), .B2(n15926), .ZN(n15908) );
  OAI21_X1 U19488 ( .B1(n15928), .B2(n21432), .A(n15908), .ZN(n15909) );
  AOI21_X1 U19489 ( .B1(n15930), .B2(n21429), .A(n15909), .ZN(n15910) );
  OAI21_X1 U19490 ( .B1(n15932), .B2(n21397), .A(n15910), .ZN(P1_U3130) );
  AOI22_X1 U19491 ( .A1(n21928), .A2(n9851), .B1(
        P1_INSTQUEUE_REG_12__2__SCAN_IN), .B2(n15926), .ZN(n15911) );
  OAI21_X1 U19492 ( .B1(n15928), .B2(n21435), .A(n15911), .ZN(n15912) );
  AOI21_X1 U19493 ( .B1(n15930), .B2(n21929), .A(n15912), .ZN(n15913) );
  OAI21_X1 U19494 ( .B1(n15932), .B2(n21936), .A(n15913), .ZN(P1_U3131) );
  AOI22_X1 U19495 ( .A1(n21491), .A2(n9851), .B1(
        P1_INSTQUEUE_REG_12__3__SCAN_IN), .B2(n15926), .ZN(n15914) );
  OAI21_X1 U19496 ( .B1(n15928), .B2(n21439), .A(n15914), .ZN(n15915) );
  AOI21_X1 U19497 ( .B1(n15930), .B2(n21436), .A(n15915), .ZN(n15916) );
  OAI21_X1 U19498 ( .B1(n15932), .B2(n21400), .A(n15916), .ZN(P1_U3132) );
  AOI22_X1 U19499 ( .A1(n21497), .A2(n9851), .B1(
        P1_INSTQUEUE_REG_12__4__SCAN_IN), .B2(n15926), .ZN(n15917) );
  OAI21_X1 U19500 ( .B1(n15928), .B2(n21443), .A(n15917), .ZN(n15918) );
  AOI21_X1 U19501 ( .B1(n15930), .B2(n21440), .A(n15918), .ZN(n15919) );
  OAI21_X1 U19502 ( .B1(n15932), .B2(n21403), .A(n15919), .ZN(P1_U3133) );
  AOI22_X1 U19503 ( .A1(n21503), .A2(n9851), .B1(
        P1_INSTQUEUE_REG_12__5__SCAN_IN), .B2(n15926), .ZN(n15920) );
  OAI21_X1 U19504 ( .B1(n15928), .B2(n21447), .A(n15920), .ZN(n15921) );
  AOI21_X1 U19505 ( .B1(n15930), .B2(n21444), .A(n15921), .ZN(n15922) );
  OAI21_X1 U19506 ( .B1(n15932), .B2(n21406), .A(n15922), .ZN(P1_U3134) );
  AOI22_X1 U19507 ( .A1(n21509), .A2(n9851), .B1(
        P1_INSTQUEUE_REG_12__6__SCAN_IN), .B2(n15926), .ZN(n15923) );
  OAI21_X1 U19508 ( .B1(n15928), .B2(n21451), .A(n15923), .ZN(n15924) );
  AOI21_X1 U19509 ( .B1(n15930), .B2(n21448), .A(n15924), .ZN(n15925) );
  OAI21_X1 U19510 ( .B1(n15932), .B2(n21409), .A(n15925), .ZN(P1_U3135) );
  AOI22_X1 U19511 ( .A1(n21516), .A2(n9851), .B1(
        P1_INSTQUEUE_REG_12__7__SCAN_IN), .B2(n15926), .ZN(n15927) );
  OAI21_X1 U19512 ( .B1(n15928), .B2(n21459), .A(n15927), .ZN(n15929) );
  AOI21_X1 U19513 ( .B1(n15930), .B2(n21454), .A(n15929), .ZN(n15931) );
  OAI21_X1 U19514 ( .B1(n15932), .B2(n21412), .A(n15931), .ZN(P1_U3136) );
  INV_X1 U19515 ( .A(n15933), .ZN(n15948) );
  AOI22_X1 U19516 ( .A1(n15936), .A2(n15935), .B1(n15934), .B2(n11736), .ZN(
        n21592) );
  NAND2_X1 U19517 ( .A1(n15937), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n21601) );
  AND3_X1 U19518 ( .A1(n21592), .A2(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(
        n21601), .ZN(n15943) );
  INV_X1 U19519 ( .A(n15943), .ZN(n15941) );
  INV_X1 U19520 ( .A(n15938), .ZN(n15940) );
  OAI211_X1 U19521 ( .C1(n15941), .C2(n21681), .A(n15940), .B(n15939), .ZN(
        n15942) );
  OAI21_X1 U19522 ( .B1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n15943), .A(
        n15942), .ZN(n15946) );
  AOI222_X1 U19523 ( .A1(n15946), .A2(n15945), .B1(n15946), .B2(n15944), .C1(
        n15945), .C2(n15944), .ZN(n15947) );
  AOI222_X1 U19524 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n15948), 
        .B1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n15947), .C1(n15948), 
        .C2(n15947), .ZN(n15949) );
  AND2_X1 U19525 ( .A1(n15949), .A2(n21147), .ZN(n15957) );
  NOR2_X1 U19526 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(P1_MORE_REG_SCAN_IN), .ZN(
        n15953) );
  OAI211_X1 U19527 ( .C1(n15953), .C2(n15952), .A(n15951), .B(n15950), .ZN(
        n15954) );
  OAI21_X1 U19528 ( .B1(n15967), .B2(n20939), .A(n18052), .ZN(n15965) );
  NAND4_X1 U19529 ( .A1(n15960), .A2(n15959), .A3(n18008), .A4(n15958), .ZN(
        n15964) );
  OAI21_X1 U19530 ( .B1(n21532), .B2(n15962), .A(n15961), .ZN(n15963) );
  AND2_X1 U19531 ( .A1(n15964), .A2(n15963), .ZN(n18046) );
  NOR2_X1 U19532 ( .A1(n15973), .A2(n20939), .ZN(n18054) );
  OAI21_X1 U19533 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n21532), .A(n18054), 
        .ZN(n18051) );
  NAND2_X1 U19534 ( .A1(n15967), .A2(n15966), .ZN(n15970) );
  INV_X1 U19535 ( .A(n18049), .ZN(n15969) );
  NAND3_X1 U19536 ( .A1(n15970), .A2(n15969), .A3(n15968), .ZN(n15975) );
  AND2_X1 U19537 ( .A1(n15971), .A2(n18049), .ZN(n15972) );
  OAI21_X1 U19538 ( .B1(n15973), .B2(n15972), .A(n20939), .ZN(n15974) );
  OAI21_X1 U19539 ( .B1(n18051), .B2(n15975), .A(n15974), .ZN(n15976) );
  INV_X1 U19540 ( .A(n15976), .ZN(P1_U3161) );
  OAI21_X1 U19541 ( .B1(n17984), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n20812), 
        .ZN(n15977) );
  NAND3_X1 U19542 ( .A1(n15978), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n15977), 
        .ZN(n15980) );
  OAI21_X1 U19543 ( .B1(P2_STATE2_REG_1__SCAN_IN), .B2(
        P2_STATE2_REG_2__SCAN_IN), .A(n17703), .ZN(n17684) );
  OAI21_X1 U19544 ( .B1(n20819), .B2(n20742), .A(n17684), .ZN(n15979) );
  NAND2_X1 U19545 ( .A1(n15980), .A2(n15979), .ZN(n15986) );
  NOR2_X1 U19546 ( .A1(n15981), .A2(n20742), .ZN(n17680) );
  INV_X1 U19547 ( .A(n17680), .ZN(n15984) );
  NOR2_X1 U19548 ( .A1(n20819), .A2(n20240), .ZN(n15983) );
  AOI211_X1 U19549 ( .C1(n20750), .C2(n15984), .A(n15983), .B(n15982), .ZN(
        n15985) );
  MUX2_X1 U19550 ( .A(n15986), .B(P2_REQUESTPENDING_REG_SCAN_IN), .S(n15985), 
        .Z(P2_U3610) );
  OAI21_X1 U19551 ( .B1(n13062), .B2(n15988), .A(n15987), .ZN(n17160) );
  OAI21_X1 U19552 ( .B1(n16009), .B2(n16887), .A(n20204), .ZN(n15990) );
  NAND2_X1 U19553 ( .A1(n15992), .A2(n16348), .ZN(n15997) );
  INV_X1 U19554 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n15994) );
  AOI22_X1 U19555 ( .A1(n20190), .A2(P2_REIP_REG_29__SCAN_IN), .B1(n20188), 
        .B2(P2_EBX_REG_29__SCAN_IN), .ZN(n15993) );
  OAI21_X1 U19556 ( .B1(n16178), .B2(n15994), .A(n15993), .ZN(n15995) );
  INV_X1 U19557 ( .A(n15995), .ZN(n15996) );
  AOI21_X1 U19558 ( .B1(n16001), .B2(n9754), .A(n16000), .ZN(n17169) );
  NAND2_X1 U19559 ( .A1(n17169), .A2(n20195), .ZN(n16002) );
  OAI211_X1 U19560 ( .C1(n20196), .C2(n17160), .A(n16003), .B(n16002), .ZN(
        P2_U2826) );
  NAND2_X1 U19561 ( .A1(n16004), .A2(n16005), .ZN(n16006) );
  INV_X1 U19562 ( .A(n16007), .ZN(n16024) );
  OAI21_X1 U19563 ( .B1(n16024), .B2(n16008), .A(n20204), .ZN(n16010) );
  AOI21_X1 U19564 ( .B1(n16210), .B2(n16010), .A(n16009), .ZN(n16016) );
  INV_X1 U19565 ( .A(n16011), .ZN(n16012) );
  NAND2_X1 U19566 ( .A1(n16012), .A2(n16348), .ZN(n16014) );
  AOI22_X1 U19567 ( .A1(n20190), .A2(P2_REIP_REG_28__SCAN_IN), .B1(n20188), 
        .B2(P2_EBX_REG_28__SCAN_IN), .ZN(n16013) );
  OAI211_X1 U19568 ( .C1(n16178), .C2(n10440), .A(n16014), .B(n16013), .ZN(
        n16015) );
  OAI21_X1 U19569 ( .B1(n9925), .B2(n17991), .A(n16017), .ZN(P2_U2827) );
  OAI21_X1 U19570 ( .B1(n16018), .B2(n16019), .A(n16004), .ZN(n17193) );
  AND2_X1 U19571 ( .A1(n16021), .A2(n16036), .ZN(n16038) );
  OAI21_X1 U19572 ( .B1(n16038), .B2(n16023), .A(n16022), .ZN(n16899) );
  INV_X1 U19573 ( .A(n16899), .ZN(n17191) );
  OAI21_X1 U19574 ( .B1(n9756), .B2(n16898), .A(n20204), .ZN(n16025) );
  AOI21_X1 U19575 ( .B1(n16210), .B2(n16025), .A(n16024), .ZN(n16031) );
  NAND2_X1 U19576 ( .A1(n16026), .A2(n16348), .ZN(n16028) );
  AOI22_X1 U19577 ( .A1(n20190), .A2(P2_REIP_REG_27__SCAN_IN), .B1(n20188), 
        .B2(P2_EBX_REG_27__SCAN_IN), .ZN(n16027) );
  OAI211_X1 U19578 ( .C1(n16178), .C2(n16029), .A(n16028), .B(n16027), .ZN(
        n16030) );
  AOI211_X1 U19579 ( .C1(n17191), .C2(n16354), .A(n16031), .B(n16030), .ZN(
        n16032) );
  OAI21_X1 U19580 ( .B1(n17193), .B2(n17991), .A(n16032), .ZN(P2_U2828) );
  INV_X1 U19581 ( .A(n16018), .ZN(n16034) );
  OAI21_X1 U19582 ( .B1(n16033), .B2(n16035), .A(n16034), .ZN(n17198) );
  NOR2_X1 U19583 ( .A1(n16021), .A2(n16036), .ZN(n16037) );
  INV_X1 U19584 ( .A(n17205), .ZN(n16046) );
  INV_X1 U19585 ( .A(n16039), .ZN(n16054) );
  OAI21_X1 U19586 ( .B1(n16054), .B2(n16907), .A(n20204), .ZN(n16040) );
  AOI21_X1 U19587 ( .B1(n16210), .B2(n16040), .A(n9756), .ZN(n16045) );
  AOI22_X1 U19588 ( .A1(n20190), .A2(P2_REIP_REG_26__SCAN_IN), .B1(n20188), 
        .B2(P2_EBX_REG_26__SCAN_IN), .ZN(n16042) );
  NAND2_X1 U19589 ( .A1(n20189), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n16041) );
  OAI211_X1 U19590 ( .C1(n16043), .C2(n20192), .A(n16042), .B(n16041), .ZN(
        n16044) );
  AOI211_X1 U19591 ( .C1(n16046), .C2(n16354), .A(n16045), .B(n16044), .ZN(
        n16047) );
  OAI21_X1 U19592 ( .B1(n17198), .B2(n17991), .A(n16047), .ZN(P2_U2829) );
  INV_X1 U19593 ( .A(n16033), .ZN(n16050) );
  OAI21_X1 U19594 ( .B1(n16049), .B2(n16051), .A(n16050), .ZN(n17211) );
  AOI21_X1 U19595 ( .B1(n16053), .B2(n16052), .A(n16021), .ZN(n17218) );
  OAI21_X1 U19596 ( .B1(n9757), .B2(n16919), .A(n20204), .ZN(n16055) );
  AOI21_X1 U19597 ( .B1(n16210), .B2(n16055), .A(n16054), .ZN(n16060) );
  XNOR2_X1 U19598 ( .A(n9678), .B(P2_EBX_REG_25__SCAN_IN), .ZN(n16058) );
  AOI22_X1 U19599 ( .A1(n20190), .A2(P2_REIP_REG_25__SCAN_IN), .B1(n20188), 
        .B2(P2_EBX_REG_25__SCAN_IN), .ZN(n16057) );
  NAND2_X1 U19600 ( .A1(n20189), .A2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n16056) );
  OAI211_X1 U19601 ( .C1(n16058), .C2(n20192), .A(n16057), .B(n16056), .ZN(
        n16059) );
  AOI211_X1 U19602 ( .C1(n17218), .C2(n16354), .A(n16060), .B(n16059), .ZN(
        n16061) );
  OAI21_X1 U19603 ( .B1(n17211), .B2(n17991), .A(n16061), .ZN(P2_U2830) );
  NAND2_X1 U19604 ( .A1(n16084), .A2(n16063), .ZN(n16064) );
  NAND2_X1 U19605 ( .A1(n16052), .A2(n16064), .ZN(n17229) );
  XOR2_X1 U19606 ( .A(P2_EBX_REG_24__SCAN_IN), .B(n16065), .Z(n16073) );
  AOI22_X1 U19607 ( .A1(n20190), .A2(P2_REIP_REG_24__SCAN_IN), .B1(n20188), 
        .B2(P2_EBX_REG_24__SCAN_IN), .ZN(n16066) );
  OAI21_X1 U19608 ( .B1(n16178), .B2(n16067), .A(n16066), .ZN(n16072) );
  INV_X1 U19609 ( .A(n16068), .ZN(n16069) );
  OAI21_X1 U19610 ( .B1(n16069), .B2(n16925), .A(n20204), .ZN(n16070) );
  AOI21_X1 U19611 ( .B1(n16210), .B2(n16070), .A(n9757), .ZN(n16071) );
  AOI211_X1 U19612 ( .C1(n16348), .C2(n16073), .A(n16072), .B(n16071), .ZN(
        n16078) );
  AND2_X1 U19613 ( .A1(n16074), .A2(n16075), .ZN(n16076) );
  NOR2_X1 U19614 ( .A1(n16049), .A2(n16076), .ZN(n17233) );
  NAND2_X1 U19615 ( .A1(n17233), .A2(n20195), .ZN(n16077) );
  OAI211_X1 U19616 ( .C1(n20196), .C2(n17229), .A(n16078), .B(n16077), .ZN(
        P2_U2831) );
  NAND2_X1 U19617 ( .A1(n16079), .A2(n16080), .ZN(n16081) );
  NAND2_X1 U19618 ( .A1(n16074), .A2(n16081), .ZN(n17236) );
  NAND2_X1 U19619 ( .A1(n9766), .A2(n16082), .ZN(n16083) );
  AND2_X1 U19620 ( .A1(n16084), .A2(n16083), .ZN(n17246) );
  AOI21_X1 U19621 ( .B1(n16085), .B2(n10190), .A(n17996), .ZN(n16086) );
  OAI21_X1 U19622 ( .B1(n16086), .B2(n17999), .A(n16068), .ZN(n16090) );
  INV_X1 U19623 ( .A(n20188), .ZN(n16346) );
  OAI22_X1 U19624 ( .A1(n16346), .A2(n16087), .B1(n20862), .B2(n16351), .ZN(
        n16088) );
  AOI21_X1 U19625 ( .B1(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n20189), .A(
        n16088), .ZN(n16089) );
  OAI211_X1 U19626 ( .C1(n20192), .C2(n13000), .A(n16090), .B(n16089), .ZN(
        n16091) );
  AOI21_X1 U19627 ( .B1(n17246), .B2(n16354), .A(n16091), .ZN(n16092) );
  OAI21_X1 U19628 ( .B1(n17236), .B2(n17991), .A(n16092), .ZN(P2_U2832) );
  OAI211_X1 U19629 ( .C1(n16093), .C2(n16956), .A(n17998), .B(n20204), .ZN(
        n16095) );
  AOI22_X1 U19630 ( .A1(n20190), .A2(P2_REIP_REG_21__SCAN_IN), .B1(n20188), 
        .B2(P2_EBX_REG_21__SCAN_IN), .ZN(n16094) );
  OAI211_X1 U19631 ( .C1(n16178), .C2(n10448), .A(n16095), .B(n16094), .ZN(
        n16096) );
  AOI21_X1 U19632 ( .B1(n16097), .B2(n16348), .A(n16096), .ZN(n16099) );
  NAND2_X1 U19633 ( .A1(n16813), .A2(n20195), .ZN(n16098) );
  OAI211_X1 U19634 ( .C1(n16675), .C2(n20196), .A(n16099), .B(n16098), .ZN(
        P2_U2834) );
  OAI21_X1 U19635 ( .B1(n9755), .B2(n10634), .A(n16100), .ZN(n17268) );
  AOI21_X1 U19636 ( .B1(n16103), .B2(n16102), .A(n16101), .ZN(n17266) );
  NOR2_X1 U19637 ( .A1(n16104), .A2(n20192), .ZN(n16110) );
  XNOR2_X1 U19638 ( .A(n16105), .B(n16966), .ZN(n16108) );
  AOI22_X1 U19639 ( .A1(n20190), .A2(P2_REIP_REG_20__SCAN_IN), .B1(n20188), 
        .B2(P2_EBX_REG_20__SCAN_IN), .ZN(n16107) );
  NAND2_X1 U19640 ( .A1(n20189), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n16106) );
  OAI211_X1 U19641 ( .C1(n16108), .C2(n17996), .A(n16107), .B(n16106), .ZN(
        n16109) );
  AOI211_X1 U19642 ( .C1(n17266), .C2(n16354), .A(n16110), .B(n16109), .ZN(
        n16111) );
  OAI21_X1 U19643 ( .B1(n17268), .B2(n17991), .A(n16111), .ZN(P2_U2835) );
  NOR2_X1 U19644 ( .A1(n16351), .A2(n21778), .ZN(n16112) );
  AOI211_X1 U19645 ( .C1(P2_EBX_REG_19__SCAN_IN), .C2(n20188), .A(n11487), .B(
        n16112), .ZN(n16113) );
  OAI21_X1 U19646 ( .B1(n16114), .B2(n16178), .A(n16113), .ZN(n16121) );
  INV_X1 U19647 ( .A(n16322), .ZN(n16358) );
  INV_X1 U19648 ( .A(n16116), .ZN(n16115) );
  NOR2_X1 U19649 ( .A1(n16358), .A2(n16115), .ZN(n16119) );
  OAI21_X1 U19650 ( .B1(n16116), .B2(n17996), .A(n16210), .ZN(n16118) );
  MUX2_X1 U19651 ( .A(n16119), .B(n16118), .S(n16117), .Z(n16120) );
  AOI211_X1 U19652 ( .C1(n16348), .C2(n16122), .A(n16121), .B(n16120), .ZN(
        n16124) );
  NAND2_X1 U19653 ( .A1(n16827), .A2(n20195), .ZN(n16123) );
  OAI211_X1 U19654 ( .C1(n16685), .C2(n20196), .A(n16124), .B(n16123), .ZN(
        P2_U2836) );
  OAI21_X1 U19655 ( .B1(n16125), .B2(n16126), .A(n14781), .ZN(n17273) );
  AOI21_X1 U19656 ( .B1(n16127), .B2(n20204), .A(n17999), .ZN(n16129) );
  INV_X1 U19657 ( .A(n16127), .ZN(n16128) );
  NAND2_X1 U19658 ( .A1(n16322), .A2(n16128), .ZN(n16150) );
  MUX2_X1 U19659 ( .A(n16129), .B(n16150), .S(n16977), .Z(n16132) );
  NOR2_X1 U19660 ( .A1(n16351), .A2(n20855), .ZN(n16130) );
  AOI211_X1 U19661 ( .C1(P2_EBX_REG_18__SCAN_IN), .C2(n20188), .A(n11487), .B(
        n16130), .ZN(n16131) );
  OAI211_X1 U19662 ( .C1(n16178), .C2(n16133), .A(n16132), .B(n16131), .ZN(
        n16137) );
  OAI21_X1 U19663 ( .B1(n16134), .B2(n16135), .A(n13501), .ZN(n17279) );
  NOR2_X1 U19664 ( .A1(n17279), .A2(n20196), .ZN(n16136) );
  AOI211_X1 U19665 ( .C1(n16348), .C2(n16138), .A(n16137), .B(n16136), .ZN(
        n16139) );
  OAI21_X1 U19666 ( .B1(n17273), .B2(n17991), .A(n16139), .ZN(P2_U2837) );
  INV_X1 U19667 ( .A(n16125), .ZN(n16141) );
  OAI21_X1 U19668 ( .B1(n16140), .B2(n16142), .A(n16141), .ZN(n17287) );
  NOR2_X1 U19669 ( .A1(n16143), .A2(n16983), .ZN(n16149) );
  NAND2_X1 U19670 ( .A1(n20188), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n16144) );
  OAI211_X1 U19671 ( .C1(n16351), .C2(n20853), .A(n16144), .B(n17136), .ZN(
        n16145) );
  AOI21_X1 U19672 ( .B1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n20189), .A(
        n16145), .ZN(n16148) );
  INV_X1 U19673 ( .A(n16983), .ZN(n16146) );
  NAND2_X1 U19674 ( .A1(n17999), .A2(n16146), .ZN(n16147) );
  OAI211_X1 U19675 ( .C1(n16150), .C2(n16149), .A(n16148), .B(n16147), .ZN(
        n16155) );
  INV_X1 U19676 ( .A(n16134), .ZN(n16152) );
  OAI21_X1 U19677 ( .B1(n16151), .B2(n16153), .A(n16152), .ZN(n17289) );
  NOR2_X1 U19678 ( .A1(n17289), .A2(n20196), .ZN(n16154) );
  AOI211_X1 U19679 ( .C1(n16348), .C2(n16156), .A(n16155), .B(n16154), .ZN(
        n16157) );
  OAI21_X1 U19680 ( .B1(n17287), .B2(n17991), .A(n16157), .ZN(P2_U2838) );
  AOI21_X1 U19681 ( .B1(n16159), .B2(n16158), .A(n16140), .ZN(n17305) );
  INV_X1 U19682 ( .A(n17305), .ZN(n16856) );
  AND2_X1 U19683 ( .A1(n16160), .A2(n16161), .ZN(n16162) );
  OR2_X1 U19684 ( .A1(n16162), .A2(n16151), .ZN(n17300) );
  INV_X1 U19685 ( .A(n17300), .ZN(n16995) );
  INV_X1 U19686 ( .A(n16164), .ZN(n16163) );
  AOI21_X1 U19687 ( .B1(n16163), .B2(n20204), .A(n17999), .ZN(n16166) );
  NAND2_X1 U19688 ( .A1(n16322), .A2(n16164), .ZN(n16165) );
  MUX2_X1 U19689 ( .A(n16166), .B(n16165), .S(n16992), .Z(n16170) );
  NAND2_X1 U19690 ( .A1(n20188), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n16167) );
  OAI211_X1 U19691 ( .C1(n16351), .C2(n20851), .A(n16167), .B(n17136), .ZN(
        n16168) );
  AOI21_X1 U19692 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n20189), .A(
        n16168), .ZN(n16169) );
  OAI211_X1 U19693 ( .C1(n20192), .C2(n16171), .A(n16170), .B(n16169), .ZN(
        n16172) );
  AOI21_X1 U19694 ( .B1(n16995), .B2(n16354), .A(n16172), .ZN(n16173) );
  OAI21_X1 U19695 ( .B1(n16856), .B2(n17991), .A(n16173), .ZN(P2_U2839) );
  NAND2_X1 U19696 ( .A1(n16336), .A2(n16174), .ZN(n16175) );
  XOR2_X1 U19697 ( .A(n17004), .B(n16175), .Z(n16186) );
  NOR2_X1 U19698 ( .A1(n16351), .A2(n20849), .ZN(n16176) );
  AOI211_X1 U19699 ( .C1(P2_EBX_REG_15__SCAN_IN), .C2(n20188), .A(n18058), .B(
        n16176), .ZN(n16177) );
  OAI21_X1 U19700 ( .B1(n17002), .B2(n16178), .A(n16177), .ZN(n16179) );
  AOI21_X1 U19701 ( .B1(n16180), .B2(n16348), .A(n16179), .ZN(n16185) );
  NAND2_X1 U19702 ( .A1(n16181), .A2(n16182), .ZN(n16183) );
  NAND2_X1 U19703 ( .A1(n16160), .A2(n16183), .ZN(n17317) );
  INV_X1 U19704 ( .A(n17317), .ZN(n16702) );
  AOI22_X1 U19705 ( .A1(n16702), .A2(n16354), .B1(n17320), .B2(n20195), .ZN(
        n16184) );
  OAI211_X1 U19706 ( .C1(n16186), .C2(n17996), .A(n16185), .B(n16184), .ZN(
        P2_U2840) );
  AOI21_X1 U19707 ( .B1(n16187), .B2(n20204), .A(n17999), .ZN(n16190) );
  INV_X1 U19708 ( .A(n16187), .ZN(n16188) );
  NAND2_X1 U19709 ( .A1(n16322), .A2(n16188), .ZN(n16189) );
  MUX2_X1 U19710 ( .A(n16190), .B(n16189), .S(n17017), .Z(n16201) );
  NAND2_X1 U19711 ( .A1(n16191), .A2(n16192), .ZN(n16193) );
  AND2_X1 U19712 ( .A1(n16181), .A2(n16193), .ZN(n17333) );
  NAND2_X1 U19713 ( .A1(n16194), .A2(n16348), .ZN(n16198) );
  NAND2_X1 U19714 ( .A1(n20188), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n16195) );
  OAI211_X1 U19715 ( .C1(n16351), .C2(n20848), .A(n16195), .B(n17136), .ZN(
        n16196) );
  AOI21_X1 U19716 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n20189), .A(
        n16196), .ZN(n16197) );
  NAND2_X1 U19717 ( .A1(n16198), .A2(n16197), .ZN(n16199) );
  AOI21_X1 U19718 ( .B1(n17333), .B2(n16354), .A(n16199), .ZN(n16200) );
  OAI211_X1 U19719 ( .C1(n17991), .C2(n17335), .A(n16201), .B(n16200), .ZN(
        P2_U2841) );
  OR2_X1 U19720 ( .A1(n16202), .A2(n16203), .ZN(n16204) );
  NAND2_X1 U19721 ( .A1(n16191), .A2(n16204), .ZN(n17344) );
  NAND2_X1 U19722 ( .A1(n20189), .A2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n16206) );
  AOI21_X1 U19723 ( .B1(n20188), .B2(P2_EBX_REG_13__SCAN_IN), .A(n11487), .ZN(
        n16205) );
  OAI211_X1 U19724 ( .C1(n16351), .C2(n20846), .A(n16206), .B(n16205), .ZN(
        n16207) );
  AOI21_X1 U19725 ( .B1(n16208), .B2(n16348), .A(n16207), .ZN(n16209) );
  OAI21_X1 U19726 ( .B1(n17344), .B2(n20196), .A(n16209), .ZN(n16216) );
  INV_X1 U19727 ( .A(n16212), .ZN(n16211) );
  OAI21_X1 U19728 ( .B1(n16211), .B2(n17996), .A(n16210), .ZN(n16214) );
  NOR2_X1 U19729 ( .A1(n16358), .A2(n16212), .ZN(n16213) );
  MUX2_X1 U19730 ( .A(n16214), .B(n16213), .S(n17029), .Z(n16215) );
  AOI211_X1 U19731 ( .C1(n20195), .C2(n17346), .A(n16216), .B(n16215), .ZN(
        n16217) );
  INV_X1 U19732 ( .A(n16217), .ZN(P2_U2842) );
  INV_X1 U19733 ( .A(n16218), .ZN(n16219) );
  AOI21_X1 U19734 ( .B1(n16219), .B2(n20204), .A(n17999), .ZN(n16220) );
  MUX2_X1 U19735 ( .A(n16221), .B(n16220), .S(n17039), .Z(n16233) );
  AND2_X1 U19736 ( .A1(n13530), .A2(n16222), .ZN(n16223) );
  OR2_X1 U19737 ( .A1(n16202), .A2(n16223), .ZN(n17358) );
  AOI21_X1 U19738 ( .B1(n16224), .B2(P2_EBX_REG_12__SCAN_IN), .A(n20192), .ZN(
        n16229) );
  NAND2_X1 U19739 ( .A1(n20189), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n16226) );
  AOI21_X1 U19740 ( .B1(n20188), .B2(P2_EBX_REG_12__SCAN_IN), .A(n11487), .ZN(
        n16225) );
  OAI211_X1 U19741 ( .C1(n16351), .C2(n16227), .A(n16226), .B(n16225), .ZN(
        n16228) );
  AOI21_X1 U19742 ( .B1(n11091), .B2(n16229), .A(n16228), .ZN(n16230) );
  OAI21_X1 U19743 ( .B1(n17358), .B2(n20196), .A(n16230), .ZN(n16231) );
  INV_X1 U19744 ( .A(n16231), .ZN(n16232) );
  OAI211_X1 U19745 ( .C1(n17991), .C2(n17354), .A(n16233), .B(n16232), .ZN(
        P2_U2843) );
  AOI21_X1 U19746 ( .B1(n16234), .B2(n20204), .A(n17999), .ZN(n16237) );
  INV_X1 U19747 ( .A(n16234), .ZN(n16235) );
  NAND2_X1 U19748 ( .A1(n16322), .A2(n16235), .ZN(n16236) );
  MUX2_X1 U19749 ( .A(n16237), .B(n16236), .S(n17062), .Z(n16247) );
  OR2_X1 U19750 ( .A1(n16238), .A2(n16239), .ZN(n16240) );
  AND2_X1 U19751 ( .A1(n13531), .A2(n16240), .ZN(n17381) );
  INV_X1 U19752 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n20843) );
  NAND2_X1 U19753 ( .A1(n20188), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n16241) );
  OAI211_X1 U19754 ( .C1(n16351), .C2(n20843), .A(n16241), .B(n17136), .ZN(
        n16242) );
  AOI21_X1 U19755 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n20189), .A(
        n16242), .ZN(n16243) );
  OAI21_X1 U19756 ( .B1(n16244), .B2(n20192), .A(n16243), .ZN(n16245) );
  AOI21_X1 U19757 ( .B1(n17381), .B2(n16354), .A(n16245), .ZN(n16246) );
  OAI211_X1 U19758 ( .C1(n17991), .C2(n16248), .A(n16247), .B(n16246), .ZN(
        P2_U2845) );
  NOR2_X1 U19759 ( .A1(n12943), .A2(n16249), .ZN(n16250) );
  XNOR2_X1 U19760 ( .A(n16250), .B(n17074), .ZN(n16261) );
  NOR2_X1 U19761 ( .A1(n17393), .A2(n17991), .ZN(n16260) );
  NOR2_X1 U19762 ( .A1(n16251), .A2(n16252), .ZN(n16253) );
  OR2_X1 U19763 ( .A1(n16238), .A2(n16253), .ZN(n17397) );
  NAND2_X1 U19764 ( .A1(n20189), .A2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16255) );
  AOI21_X1 U19765 ( .B1(n20188), .B2(P2_EBX_REG_9__SCAN_IN), .A(n11487), .ZN(
        n16254) );
  OAI211_X1 U19766 ( .C1(n16351), .C2(n20841), .A(n16255), .B(n16254), .ZN(
        n16256) );
  AOI21_X1 U19767 ( .B1(n16257), .B2(n16348), .A(n16256), .ZN(n16258) );
  OAI21_X1 U19768 ( .B1(n17397), .B2(n20196), .A(n16258), .ZN(n16259) );
  AOI211_X1 U19769 ( .C1(n16261), .C2(n20204), .A(n16260), .B(n16259), .ZN(
        n16262) );
  INV_X1 U19770 ( .A(n16262), .ZN(P2_U2846) );
  INV_X1 U19771 ( .A(n16264), .ZN(n16263) );
  AOI21_X1 U19772 ( .B1(n16263), .B2(n20204), .A(n17999), .ZN(n16266) );
  NAND2_X1 U19773 ( .A1(n16322), .A2(n16264), .ZN(n16265) );
  MUX2_X1 U19774 ( .A(n16266), .B(n16265), .S(n17092), .Z(n16275) );
  AND2_X1 U19775 ( .A1(n14518), .A2(n16267), .ZN(n16268) );
  OR2_X1 U19776 ( .A1(n16268), .A2(n16251), .ZN(n17090) );
  INV_X1 U19777 ( .A(n17090), .ZN(n17409) );
  AOI21_X1 U19778 ( .B1(n20188), .B2(P2_EBX_REG_8__SCAN_IN), .A(n11487), .ZN(
        n16269) );
  OAI21_X1 U19779 ( .B1(n20839), .B2(n16351), .A(n16269), .ZN(n16270) );
  AOI21_X1 U19780 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n20189), .A(
        n16270), .ZN(n16271) );
  OAI21_X1 U19781 ( .B1(n16272), .B2(n20192), .A(n16271), .ZN(n16273) );
  AOI21_X1 U19782 ( .B1(n17409), .B2(n16354), .A(n16273), .ZN(n16274) );
  OAI211_X1 U19783 ( .C1(n17991), .C2(n17412), .A(n16275), .B(n16274), .ZN(
        P2_U2847) );
  NAND2_X1 U19784 ( .A1(n16322), .A2(n16276), .ZN(n16278) );
  AOI21_X1 U19785 ( .B1(n10195), .B2(n20204), .A(n17999), .ZN(n16277) );
  MUX2_X1 U19786 ( .A(n16278), .B(n16277), .S(n18062), .Z(n16286) );
  NAND2_X1 U19787 ( .A1(n16279), .A2(n16348), .ZN(n16283) );
  NAND2_X1 U19788 ( .A1(n20188), .A2(P2_EBX_REG_7__SCAN_IN), .ZN(n16280) );
  OAI211_X1 U19789 ( .C1(n16351), .C2(n20837), .A(n16280), .B(n17136), .ZN(
        n16281) );
  AOI21_X1 U19790 ( .B1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n20189), .A(
        n16281), .ZN(n16282) );
  NAND2_X1 U19791 ( .A1(n16283), .A2(n16282), .ZN(n16284) );
  AOI21_X1 U19792 ( .B1(n18080), .B2(n16354), .A(n16284), .ZN(n16285) );
  OAI211_X1 U19793 ( .C1(n17991), .C2(n18073), .A(n16286), .B(n16285), .ZN(
        P2_U2848) );
  AOI21_X1 U19794 ( .B1(n16287), .B2(n20204), .A(n17999), .ZN(n16289) );
  NAND2_X1 U19795 ( .A1(n16322), .A2(n10196), .ZN(n16288) );
  MUX2_X1 U19796 ( .A(n16289), .B(n16288), .S(n17101), .Z(n16296) );
  NAND2_X1 U19797 ( .A1(n20188), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n16290) );
  OAI211_X1 U19798 ( .C1(n16351), .C2(n20835), .A(n16290), .B(n17136), .ZN(
        n16291) );
  AOI21_X1 U19799 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n20189), .A(
        n16291), .ZN(n16292) );
  OAI21_X1 U19800 ( .B1(n16293), .B2(n20192), .A(n16292), .ZN(n16294) );
  AOI21_X1 U19801 ( .B1(n17423), .B2(n16354), .A(n16294), .ZN(n16295) );
  OAI211_X1 U19802 ( .C1(n17426), .C2(n17991), .A(n16296), .B(n16295), .ZN(
        P2_U2849) );
  NAND2_X1 U19803 ( .A1(n16336), .A2(n20203), .ZN(n16297) );
  XOR2_X1 U19804 ( .A(n17113), .B(n16297), .Z(n16308) );
  XOR2_X1 U19805 ( .A(n16860), .B(n16298), .Z(n17440) );
  NAND2_X1 U19806 ( .A1(n20188), .A2(P2_EBX_REG_5__SCAN_IN), .ZN(n16299) );
  OAI211_X1 U19807 ( .C1(n16351), .C2(n16300), .A(n16299), .B(n17136), .ZN(
        n16301) );
  AOI21_X1 U19808 ( .B1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n20189), .A(
        n16301), .ZN(n16305) );
  INV_X1 U19809 ( .A(n16302), .ZN(n16303) );
  NAND2_X1 U19810 ( .A1(n16303), .A2(n16348), .ZN(n16304) );
  OAI211_X1 U19811 ( .C1(n17434), .C2(n20196), .A(n16305), .B(n16304), .ZN(
        n16306) );
  AOI21_X1 U19812 ( .B1(n20195), .B2(n17440), .A(n16306), .ZN(n16307) );
  OAI21_X1 U19813 ( .B1(n16308), .B2(n17996), .A(n16307), .ZN(P2_U2850) );
  AOI21_X1 U19814 ( .B1(n16309), .B2(n20204), .A(n17999), .ZN(n16312) );
  INV_X1 U19815 ( .A(n16309), .ZN(n16310) );
  NAND2_X1 U19816 ( .A1(n16322), .A2(n16310), .ZN(n16311) );
  MUX2_X1 U19817 ( .A(n16312), .B(n16311), .S(n17138), .Z(n16320) );
  NOR2_X1 U19818 ( .A1(n20192), .A2(n16314), .ZN(n16316) );
  OAI22_X1 U19819 ( .A1(n16346), .A2(n11004), .B1(n17135), .B2(n16351), .ZN(
        n16315) );
  AOI211_X1 U19820 ( .C1(n20189), .C2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n16316), .B(n16315), .ZN(n16317) );
  OAI21_X1 U19821 ( .B1(n17991), .B2(n18090), .A(n16317), .ZN(n16318) );
  AOI21_X1 U19822 ( .B1(n10798), .B2(n16354), .A(n16318), .ZN(n16319) );
  OAI211_X1 U19823 ( .C1(n20535), .C2(n20197), .A(n16320), .B(n16319), .ZN(
        P2_U2852) );
  AOI21_X1 U19824 ( .B1(n16334), .B2(n20204), .A(n17999), .ZN(n16324) );
  INV_X1 U19825 ( .A(n16334), .ZN(n16321) );
  NAND2_X1 U19826 ( .A1(n16322), .A2(n16321), .ZN(n16323) );
  MUX2_X1 U19827 ( .A(n16324), .B(n16323), .S(n17145), .Z(n16331) );
  NAND2_X1 U19828 ( .A1(n20276), .A2(n20195), .ZN(n16327) );
  OAI22_X1 U19829 ( .A1(n16346), .A2(n11013), .B1(n20830), .B2(n16351), .ZN(
        n16325) );
  AOI21_X1 U19830 ( .B1(n20189), .B2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n16325), .ZN(n16326) );
  OAI211_X1 U19831 ( .C1(n20192), .C2(n16328), .A(n16327), .B(n16326), .ZN(
        n16329) );
  AOI21_X1 U19832 ( .B1(n20281), .B2(n16354), .A(n16329), .ZN(n16330) );
  OAI211_X1 U19833 ( .C1(n20197), .C2(n20896), .A(n16331), .B(n16330), .ZN(
        P2_U2853) );
  AND2_X1 U19834 ( .A1(n16332), .A2(n17445), .ZN(n16333) );
  NOR2_X1 U19835 ( .A1(n16334), .A2(n16333), .ZN(n16335) );
  NAND2_X1 U19836 ( .A1(n16336), .A2(n16335), .ZN(n17466) );
  NAND2_X1 U19837 ( .A1(n17999), .A2(n21776), .ZN(n16343) );
  AOI22_X1 U19838 ( .A1(n20189), .A2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B1(
        n20195), .B2(n20907), .ZN(n16339) );
  AOI22_X1 U19839 ( .A1(n16348), .A2(n16337), .B1(P2_EBX_REG_1__SCAN_IN), .B2(
        n20188), .ZN(n16338) );
  OAI211_X1 U19840 ( .C1(n20829), .C2(n16351), .A(n16339), .B(n16338), .ZN(
        n16341) );
  NOR2_X1 U19841 ( .A1(n17513), .A2(n20197), .ZN(n16340) );
  AOI211_X1 U19842 ( .C1(n16354), .C2(n17467), .A(n16341), .B(n16340), .ZN(
        n16342) );
  OAI211_X1 U19843 ( .C1(n17466), .C2(n17996), .A(n16343), .B(n16342), .ZN(
        P2_U2854) );
  INV_X1 U19844 ( .A(n17445), .ZN(n16357) );
  OAI22_X1 U19845 ( .A1(n16346), .A2(n16345), .B1(n17991), .B2(n16344), .ZN(
        n16347) );
  AOI21_X1 U19846 ( .B1(n16349), .B2(n16348), .A(n16347), .ZN(n16350) );
  OAI21_X1 U19847 ( .B1(n20183), .B2(n16351), .A(n16350), .ZN(n16353) );
  NOR2_X1 U19848 ( .A1(n20914), .A2(n20197), .ZN(n16352) );
  AOI211_X1 U19849 ( .C1(n16354), .C2(n10091), .A(n16353), .B(n16352), .ZN(
        n16356) );
  OAI21_X1 U19850 ( .B1(n17999), .B2(n20189), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n16355) );
  OAI211_X1 U19851 ( .C1(n16358), .C2(n16357), .A(n16356), .B(n16355), .ZN(
        P2_U2855) );
  AND4_X1 U19852 ( .A1(n16360), .A2(n16711), .A3(n16359), .A4(n16719), .ZN(
        n16364) );
  AND4_X1 U19853 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__5__SCAN_IN), .A3(P2_INSTQUEUE_REG_0__7__SCAN_IN), 
        .A4(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n16361) );
  AND3_X1 U19854 ( .A1(n16739), .A2(n16700), .A3(n16361), .ZN(n16363) );
  NAND4_X1 U19855 ( .A1(n16364), .A2(n16363), .A3(n16362), .A4(n16731), .ZN(
        n16365) );
  NOR2_X1 U19856 ( .A1(n16365), .A2(n16563), .ZN(n16366) );
  AOI22_X1 U19857 ( .A1(n11190), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n16411), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n16371) );
  AOI22_X1 U19858 ( .A1(n10841), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n16464), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n16370) );
  AOI22_X1 U19859 ( .A1(n16466), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n16465), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n16369) );
  AOI22_X1 U19860 ( .A1(n10842), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10891), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n16368) );
  NAND4_X1 U19861 ( .A1(n16371), .A2(n16370), .A3(n16369), .A4(n16368), .ZN(
        n16377) );
  AOI22_X1 U19862 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n16472), .B1(
        n16471), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n16375) );
  AOI22_X1 U19863 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n16473), .B1(
        n17505), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n16374) );
  AOI22_X1 U19864 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n10848), .B1(
        n16437), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n16373) );
  AOI22_X1 U19865 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n10847), .B1(
        n16438), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n16372) );
  NAND4_X1 U19866 ( .A1(n16375), .A2(n16374), .A3(n16373), .A4(n16372), .ZN(
        n16376) );
  NOR2_X1 U19867 ( .A1(n16377), .A2(n16376), .ZN(n16695) );
  INV_X1 U19868 ( .A(n16695), .ZN(n16378) );
  AOI22_X1 U19869 ( .A1(n11190), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n16411), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n16382) );
  AOI22_X1 U19870 ( .A1(n10841), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n16464), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n16381) );
  AOI22_X1 U19871 ( .A1(n16466), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n16465), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n16380) );
  AOI22_X1 U19872 ( .A1(n10842), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n10891), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n16379) );
  NAND4_X1 U19873 ( .A1(n16382), .A2(n16381), .A3(n16380), .A4(n16379), .ZN(
        n16388) );
  AOI22_X1 U19874 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n16472), .B1(
        n16471), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n16386) );
  AOI22_X1 U19875 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n17505), .B1(
        n16473), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n16385) );
  AOI22_X1 U19876 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n10848), .B1(
        n16437), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n16384) );
  AOI22_X1 U19877 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n10847), .B1(
        n16438), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n16383) );
  NAND4_X1 U19878 ( .A1(n16386), .A2(n16385), .A3(n16384), .A4(n16383), .ZN(
        n16387) );
  NOR2_X1 U19879 ( .A1(n16388), .A2(n16387), .ZN(n16691) );
  AOI22_X1 U19880 ( .A1(n11190), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n16411), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n16392) );
  AOI22_X1 U19881 ( .A1(n10841), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n16464), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n16391) );
  AOI22_X1 U19882 ( .A1(n16466), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n16465), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n16390) );
  AOI22_X1 U19883 ( .A1(n10842), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10891), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n16389) );
  NAND4_X1 U19884 ( .A1(n16392), .A2(n16391), .A3(n16390), .A4(n16389), .ZN(
        n16398) );
  AOI22_X1 U19885 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n16472), .B1(
        n16471), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n16396) );
  AOI22_X1 U19886 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n17505), .B1(
        n16473), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n16395) );
  AOI22_X1 U19887 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n10848), .B1(
        n16437), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n16394) );
  AOI22_X1 U19888 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n10847), .B1(
        n16438), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n16393) );
  NAND4_X1 U19889 ( .A1(n16396), .A2(n16395), .A3(n16394), .A4(n16393), .ZN(
        n16397) );
  NAND2_X1 U19890 ( .A1(n16686), .A2(n16687), .ZN(n16681) );
  AOI22_X1 U19891 ( .A1(n11190), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n16411), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n16402) );
  AOI22_X1 U19892 ( .A1(n10841), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n16464), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n16401) );
  AOI22_X1 U19893 ( .A1(n16466), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n16465), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n16400) );
  AOI22_X1 U19894 ( .A1(n10842), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10891), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n16399) );
  NAND4_X1 U19895 ( .A1(n16402), .A2(n16401), .A3(n16400), .A4(n16399), .ZN(
        n16408) );
  AOI22_X1 U19896 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n16472), .B1(
        n16471), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n16406) );
  AOI22_X1 U19897 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n17505), .B1(
        n16473), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n16405) );
  AOI22_X1 U19898 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n10848), .B1(
        n16437), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n16404) );
  AOI22_X1 U19899 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n10847), .B1(
        n16438), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n16403) );
  NAND4_X1 U19900 ( .A1(n16406), .A2(n16405), .A3(n16404), .A4(n16403), .ZN(
        n16407) );
  NOR2_X1 U19901 ( .A1(n16408), .A2(n16407), .ZN(n16682) );
  AOI22_X1 U19902 ( .A1(n11190), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n16411), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n16415) );
  AOI22_X1 U19903 ( .A1(n10841), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n16464), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n16414) );
  AOI22_X1 U19904 ( .A1(n16466), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n16465), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n16413) );
  AOI22_X1 U19905 ( .A1(n10842), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n10891), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n16412) );
  NAND4_X1 U19906 ( .A1(n16415), .A2(n16414), .A3(n16413), .A4(n16412), .ZN(
        n16421) );
  AOI22_X1 U19907 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n16472), .B1(
        n16471), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n16419) );
  AOI22_X1 U19908 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n17505), .B1(
        n16473), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n16418) );
  AOI22_X1 U19909 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n10848), .B1(
        n16437), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n16417) );
  AOI22_X1 U19910 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n10847), .B1(
        n16438), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n16416) );
  NAND4_X1 U19911 ( .A1(n16419), .A2(n16418), .A3(n16417), .A4(n16416), .ZN(
        n16420) );
  NOR2_X1 U19912 ( .A1(n16421), .A2(n16420), .ZN(n16677) );
  INV_X1 U19913 ( .A(n16677), .ZN(n16422) );
  AOI22_X1 U19914 ( .A1(n11190), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n16411), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n16426) );
  AOI22_X1 U19915 ( .A1(n10841), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n16464), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n16425) );
  AOI22_X1 U19916 ( .A1(n16466), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n16465), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n16424) );
  AOI22_X1 U19917 ( .A1(n10842), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10891), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n16423) );
  NAND4_X1 U19918 ( .A1(n16426), .A2(n16425), .A3(n16424), .A4(n16423), .ZN(
        n16432) );
  AOI22_X1 U19919 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n16472), .B1(
        n16471), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n16430) );
  AOI22_X1 U19920 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n16473), .B1(
        n17505), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n16429) );
  AOI22_X1 U19921 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n10848), .B1(
        n16437), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n16428) );
  AOI22_X1 U19922 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n10847), .B1(
        n16438), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n16427) );
  NAND4_X1 U19923 ( .A1(n16430), .A2(n16429), .A3(n16428), .A4(n16427), .ZN(
        n16431) );
  NOR2_X1 U19924 ( .A1(n16432), .A2(n16431), .ZN(n16673) );
  AOI22_X1 U19925 ( .A1(n11190), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n16411), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n16436) );
  AOI22_X1 U19926 ( .A1(n10841), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n16464), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n16435) );
  AOI22_X1 U19927 ( .A1(n16466), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n16465), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n16434) );
  AOI22_X1 U19928 ( .A1(n10842), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n10891), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n16433) );
  NAND4_X1 U19929 ( .A1(n16436), .A2(n16435), .A3(n16434), .A4(n16433), .ZN(
        n16444) );
  AOI22_X1 U19930 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n16472), .B1(
        n16471), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n16442) );
  AOI22_X1 U19931 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n17505), .B1(
        n16473), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n16441) );
  AOI22_X1 U19932 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n10848), .B1(
        n16437), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n16440) );
  AOI22_X1 U19933 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n10847), .B1(
        n16438), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n16439) );
  NAND4_X1 U19934 ( .A1(n16442), .A2(n16441), .A3(n16440), .A4(n16439), .ZN(
        n16443) );
  AOI22_X1 U19935 ( .A1(n16612), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n9705), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n16455) );
  AOI22_X1 U19936 ( .A1(n9708), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n16613), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n16454) );
  AOI22_X1 U19937 ( .A1(n16489), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17500), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n16453) );
  AND2_X1 U19938 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n16449) );
  OR2_X1 U19939 ( .A1(n16449), .A2(n16448), .ZN(n16611) );
  INV_X1 U19940 ( .A(n16611), .ZN(n16588) );
  NAND2_X1 U19941 ( .A1(n9699), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n16450) );
  AND3_X1 U19942 ( .A1(n16588), .A2(n16451), .A3(n16450), .ZN(n16452) );
  NAND4_X1 U19943 ( .A1(n16455), .A2(n16454), .A3(n16453), .A4(n16452), .ZN(
        n16463) );
  AOI22_X1 U19944 ( .A1(n16612), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n9708), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n16461) );
  NAND2_X1 U19945 ( .A1(n16614), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n16456) );
  AND3_X1 U19946 ( .A1(n16457), .A2(n16611), .A3(n16456), .ZN(n16460) );
  AOI22_X1 U19947 ( .A1(n9680), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(n9684), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n16459) );
  AOI22_X1 U19948 ( .A1(n16489), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17500), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n16458) );
  NAND4_X1 U19949 ( .A1(n16461), .A2(n16460), .A3(n16459), .A4(n16458), .ZN(
        n16462) );
  NAND2_X1 U19950 ( .A1(n16463), .A2(n16462), .ZN(n16502) );
  NOR2_X1 U19951 ( .A1(n9710), .A2(n16502), .ZN(n16481) );
  AOI22_X1 U19952 ( .A1(n11190), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n16411), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n16470) );
  AOI22_X1 U19953 ( .A1(n10841), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n16464), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n16469) );
  AOI22_X1 U19954 ( .A1(n16466), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n16465), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n16468) );
  AOI22_X1 U19955 ( .A1(n10842), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n10891), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n16467) );
  NAND4_X1 U19956 ( .A1(n16470), .A2(n16469), .A3(n16468), .A4(n16467), .ZN(
        n16480) );
  AOI22_X1 U19957 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n16472), .B1(
        n16471), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n16478) );
  AOI22_X1 U19958 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n17505), .B1(
        n16473), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n16477) );
  AOI22_X1 U19959 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n10848), .B1(
        n16437), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n16476) );
  AOI22_X1 U19960 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n10847), .B1(
        n16438), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n16475) );
  NAND4_X1 U19961 ( .A1(n16478), .A2(n16477), .A3(n16476), .A4(n16475), .ZN(
        n16479) );
  XNOR2_X1 U19962 ( .A(n16481), .B(n16499), .ZN(n16503) );
  INV_X1 U19963 ( .A(n16502), .ZN(n16498) );
  NAND2_X1 U19964 ( .A1(n9710), .A2(n16498), .ZN(n16660) );
  AOI22_X1 U19965 ( .A1(n16612), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n16445), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n16488) );
  AOI22_X1 U19966 ( .A1(n9708), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n16613), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n16487) );
  NAND2_X1 U19967 ( .A1(n17500), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n16482) );
  AND3_X1 U19968 ( .A1(n16588), .A2(n16483), .A3(n16482), .ZN(n16486) );
  AOI22_X1 U19969 ( .A1(n16489), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n9699), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n16485) );
  NAND4_X1 U19970 ( .A1(n16488), .A2(n16487), .A3(n16486), .A4(n16485), .ZN(
        n16497) );
  AOI22_X1 U19971 ( .A1(n16612), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n9679), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n16495) );
  AOI22_X1 U19972 ( .A1(n9708), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n16613), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n16494) );
  AOI22_X1 U19973 ( .A1(n16489), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n16614), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n16493) );
  NAND2_X1 U19974 ( .A1(n17500), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n16490) );
  AND3_X1 U19975 ( .A1(n16491), .A2(n16611), .A3(n16490), .ZN(n16492) );
  NAND4_X1 U19976 ( .A1(n16495), .A2(n16494), .A3(n16493), .A4(n16492), .ZN(
        n16496) );
  AND2_X1 U19977 ( .A1(n16497), .A2(n16496), .ZN(n16501) );
  AND2_X1 U19978 ( .A1(n16499), .A2(n16498), .ZN(n16500) );
  NAND2_X1 U19979 ( .A1(n16500), .A2(n16501), .ZN(n16505) );
  OAI211_X1 U19980 ( .C1(n16501), .C2(n16500), .A(n16536), .B(n16505), .ZN(
        n16654) );
  NAND2_X1 U19981 ( .A1(n9710), .A2(n16501), .ZN(n16656) );
  NOR3_X1 U19982 ( .A1(n16503), .A2(n16502), .A3(n16656), .ZN(n16504) );
  INV_X1 U19983 ( .A(n16505), .ZN(n16520) );
  AOI22_X1 U19984 ( .A1(n16612), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n9708), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n16511) );
  NAND2_X1 U19985 ( .A1(n17500), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n16506) );
  AND3_X1 U19986 ( .A1(n16588), .A2(n16507), .A3(n16506), .ZN(n16510) );
  AOI22_X1 U19987 ( .A1(n9680), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9684), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n16509) );
  AOI22_X1 U19988 ( .A1(n16489), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9699), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n16508) );
  NAND4_X1 U19989 ( .A1(n16511), .A2(n16510), .A3(n16509), .A4(n16508), .ZN(
        n16519) );
  AOI22_X1 U19990 ( .A1(n16612), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n9708), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n16517) );
  INV_X1 U19991 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n20303) );
  NAND2_X1 U19992 ( .A1(n17500), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n16512) );
  AND3_X1 U19993 ( .A1(n16513), .A2(n16611), .A3(n16512), .ZN(n16516) );
  AOI22_X1 U19994 ( .A1(n9680), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n16613), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n16515) );
  AOI22_X1 U19995 ( .A1(n16489), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n9698), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n16514) );
  NAND4_X1 U19996 ( .A1(n16517), .A2(n16516), .A3(n16515), .A4(n16514), .ZN(
        n16518) );
  AND2_X1 U19997 ( .A1(n16519), .A2(n16518), .ZN(n16543) );
  NAND2_X1 U19998 ( .A1(n16520), .A2(n16543), .ZN(n16535) );
  OAI211_X1 U19999 ( .C1(n16520), .C2(n16543), .A(n16535), .B(n16536), .ZN(
        n16540) );
  INV_X1 U20000 ( .A(n16641), .ZN(n16539) );
  AOI22_X1 U20001 ( .A1(n16612), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n9679), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n16526) );
  AOI22_X1 U20002 ( .A1(n9708), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n9685), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n16525) );
  NAND2_X1 U20003 ( .A1(n17500), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n16521) );
  AND3_X1 U20004 ( .A1(n16588), .A2(n16522), .A3(n16521), .ZN(n16524) );
  AOI22_X1 U20005 ( .A1(n16489), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9698), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n16523) );
  NAND4_X1 U20006 ( .A1(n16526), .A2(n16525), .A3(n16524), .A4(n16523), .ZN(
        n16534) );
  AOI22_X1 U20007 ( .A1(n16612), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n9705), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n16532) );
  AOI22_X1 U20008 ( .A1(n9708), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(n9685), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n16531) );
  AOI22_X1 U20009 ( .A1(n16489), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n9699), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n16530) );
  NAND2_X1 U20010 ( .A1(n17500), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n16527) );
  AND3_X1 U20011 ( .A1(n16528), .A2(n16611), .A3(n16527), .ZN(n16529) );
  NAND4_X1 U20012 ( .A1(n16532), .A2(n16531), .A3(n16530), .A4(n16529), .ZN(
        n16533) );
  AND2_X1 U20013 ( .A1(n16534), .A2(n16533), .ZN(n16545) );
  INV_X1 U20014 ( .A(n16535), .ZN(n16537) );
  INV_X1 U20015 ( .A(n16545), .ZN(n16642) );
  OAI211_X1 U20016 ( .C1(n16545), .C2(n16537), .A(n16564), .B(n16536), .ZN(
        n16644) );
  NAND2_X1 U20017 ( .A1(n16539), .A2(n16538), .ZN(n16548) );
  INV_X1 U20018 ( .A(n16540), .ZN(n16541) );
  INV_X1 U20019 ( .A(n16543), .ZN(n16544) );
  NOR2_X1 U20020 ( .A1(n17984), .A2(n16544), .ZN(n16650) );
  AND2_X1 U20021 ( .A1(n16650), .A2(n16545), .ZN(n16546) );
  AOI22_X1 U20022 ( .A1(n16612), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n16445), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n16554) );
  AOI22_X1 U20023 ( .A1(n9708), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n9685), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n16553) );
  NAND2_X1 U20024 ( .A1(n17500), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n16549) );
  AND3_X1 U20025 ( .A1(n16588), .A2(n16550), .A3(n16549), .ZN(n16552) );
  AOI22_X1 U20026 ( .A1(n16489), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n9699), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n16551) );
  NAND4_X1 U20027 ( .A1(n16554), .A2(n16553), .A3(n16552), .A4(n16551), .ZN(
        n16562) );
  AOI22_X1 U20028 ( .A1(n16612), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n9679), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n16560) );
  AOI22_X1 U20029 ( .A1(n9708), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(n9685), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n16559) );
  AOI22_X1 U20030 ( .A1(n16489), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n9699), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n16558) );
  NAND2_X1 U20031 ( .A1(n17500), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n16555) );
  AND3_X1 U20032 ( .A1(n16556), .A2(n16611), .A3(n16555), .ZN(n16557) );
  NAND4_X1 U20033 ( .A1(n16560), .A2(n16559), .A3(n16558), .A4(n16557), .ZN(
        n16561) );
  NAND2_X1 U20034 ( .A1(n16562), .A2(n16561), .ZN(n16567) );
  NOR2_X1 U20035 ( .A1(n16564), .A2(n16567), .ZN(n16584) );
  AOI211_X1 U20036 ( .C1(n16567), .C2(n16564), .A(n16563), .B(n16584), .ZN(
        n16565) );
  OAI21_X1 U20037 ( .B1(n16566), .B2(n16565), .A(n16569), .ZN(n16637) );
  INV_X1 U20038 ( .A(n16567), .ZN(n16568) );
  NAND2_X1 U20039 ( .A1(n9710), .A2(n16568), .ZN(n16636) );
  AOI22_X1 U20040 ( .A1(n16612), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n16445), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n16575) );
  AOI22_X1 U20041 ( .A1(n9708), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n16613), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n16574) );
  NAND2_X1 U20042 ( .A1(n17500), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n16570) );
  AND3_X1 U20043 ( .A1(n16588), .A2(n16571), .A3(n16570), .ZN(n16573) );
  AOI22_X1 U20044 ( .A1(n16489), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n16614), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n16572) );
  NAND4_X1 U20045 ( .A1(n16575), .A2(n16574), .A3(n16573), .A4(n16572), .ZN(
        n16583) );
  AOI22_X1 U20046 ( .A1(n16612), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n9705), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n16581) );
  AOI22_X1 U20047 ( .A1(n9708), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(n9684), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n16580) );
  AOI22_X1 U20048 ( .A1(n16489), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n9698), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n16579) );
  NAND2_X1 U20049 ( .A1(n17500), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n16576) );
  AND3_X1 U20050 ( .A1(n16577), .A2(n16611), .A3(n16576), .ZN(n16578) );
  NAND4_X1 U20051 ( .A1(n16581), .A2(n16580), .A3(n16579), .A4(n16578), .ZN(
        n16582) );
  AND2_X1 U20052 ( .A1(n16583), .A2(n16582), .ZN(n16631) );
  INV_X1 U20053 ( .A(n16584), .ZN(n16630) );
  NAND2_X1 U20054 ( .A1(n17984), .A2(n16631), .ZN(n16585) );
  NOR2_X1 U20055 ( .A1(n16630), .A2(n16585), .ZN(n16603) );
  AOI22_X1 U20056 ( .A1(n16612), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n9708), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n16592) );
  NAND2_X1 U20057 ( .A1(n9698), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n16586) );
  AND3_X1 U20058 ( .A1(n16588), .A2(n16587), .A3(n16586), .ZN(n16591) );
  AOI22_X1 U20059 ( .A1(n16445), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n16613), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n16590) );
  AOI22_X1 U20060 ( .A1(n16489), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17500), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n16589) );
  NAND4_X1 U20061 ( .A1(n16592), .A2(n16591), .A3(n16590), .A4(n16589), .ZN(
        n16601) );
  AOI22_X1 U20062 ( .A1(n16445), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n16593), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n16599) );
  NAND2_X1 U20063 ( .A1(n9699), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n16594) );
  AND3_X1 U20064 ( .A1(n16595), .A2(n16611), .A3(n16594), .ZN(n16598) );
  AOI22_X1 U20065 ( .A1(n16612), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n9685), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n16597) );
  AOI22_X1 U20066 ( .A1(n9708), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17500), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n16596) );
  NAND4_X1 U20067 ( .A1(n16599), .A2(n16598), .A3(n16597), .A4(n16596), .ZN(
        n16600) );
  AND2_X1 U20068 ( .A1(n16601), .A2(n16600), .ZN(n16602) );
  NAND2_X1 U20069 ( .A1(n16603), .A2(n16602), .ZN(n16604) );
  OAI21_X1 U20070 ( .B1(n16603), .B2(n16602), .A(n16604), .ZN(n16626) );
  AOI22_X1 U20071 ( .A1(n16612), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17500), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n16607) );
  NAND2_X1 U20072 ( .A1(n16614), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n16605) );
  NAND4_X1 U20073 ( .A1(n16607), .A2(n16606), .A3(n16605), .A4(n16611), .ZN(
        n16621) );
  AOI22_X1 U20074 ( .A1(n9705), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(n9708), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n16609) );
  AOI22_X1 U20075 ( .A1(n16489), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n9684), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n16608) );
  NAND2_X1 U20076 ( .A1(n16609), .A2(n16608), .ZN(n16620) );
  AOI211_X1 U20077 ( .C1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .C2(n17500), .A(
        n16611), .B(n16610), .ZN(n16618) );
  AOI22_X1 U20078 ( .A1(n16612), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n9705), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n16617) );
  AOI22_X1 U20079 ( .A1(n9708), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9685), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n16616) );
  AOI22_X1 U20080 ( .A1(n16489), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9699), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n16615) );
  NAND4_X1 U20081 ( .A1(n16618), .A2(n16617), .A3(n16616), .A4(n16615), .ZN(
        n16619) );
  OAI21_X1 U20082 ( .B1(n16621), .B2(n16620), .A(n16619), .ZN(n16622) );
  XNOR2_X1 U20083 ( .A(n16623), .B(n16622), .ZN(n16755) );
  NOR2_X1 U20084 ( .A1(n16879), .A2(n16723), .ZN(n16624) );
  AOI21_X1 U20085 ( .B1(P2_EBX_REG_30__SCAN_IN), .B2(n16723), .A(n16624), .ZN(
        n16625) );
  OAI21_X1 U20086 ( .B1(n16755), .B2(n16733), .A(n16625), .ZN(P2_U2857) );
  NAND2_X1 U20087 ( .A1(n16627), .A2(n16626), .ZN(n16756) );
  NAND3_X1 U20088 ( .A1(n9724), .A2(n16737), .A3(n16756), .ZN(n16629) );
  NAND2_X1 U20089 ( .A1(n16723), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n16628) );
  OAI211_X1 U20090 ( .C1(n17160), .C2(n16723), .A(n16629), .B(n16628), .ZN(
        P2_U2858) );
  NAND2_X1 U20091 ( .A1(n16569), .A2(n16630), .ZN(n16632) );
  XNOR2_X1 U20092 ( .A(n16632), .B(n16631), .ZN(n16770) );
  NOR2_X1 U20093 ( .A1(n17183), .A2(n16723), .ZN(n16634) );
  AOI21_X1 U20094 ( .B1(P2_EBX_REG_28__SCAN_IN), .B2(n16723), .A(n16634), .ZN(
        n16635) );
  OAI21_X1 U20095 ( .B1(n16770), .B2(n16733), .A(n16635), .ZN(P2_U2859) );
  NAND2_X1 U20096 ( .A1(n16771), .A2(n16737), .ZN(n16639) );
  NAND2_X1 U20097 ( .A1(n16723), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n16638) );
  OAI211_X1 U20098 ( .C1(n16899), .C2(n16723), .A(n16639), .B(n16638), .ZN(
        P2_U2860) );
  NAND2_X1 U20099 ( .A1(n16640), .A2(n16650), .ZN(n16649) );
  NAND2_X1 U20100 ( .A1(n16641), .A2(n16649), .ZN(n16646) );
  NOR2_X1 U20101 ( .A1(n16642), .A2(n17984), .ZN(n16643) );
  XNOR2_X1 U20102 ( .A(n16644), .B(n16643), .ZN(n16645) );
  XNOR2_X1 U20103 ( .A(n16646), .B(n16645), .ZN(n16784) );
  NOR2_X1 U20104 ( .A1(n17205), .A2(n16723), .ZN(n16647) );
  AOI21_X1 U20105 ( .B1(P2_EBX_REG_26__SCAN_IN), .B2(n16723), .A(n16647), .ZN(
        n16648) );
  OAI21_X1 U20106 ( .B1(n16784), .B2(n16733), .A(n16648), .ZN(P2_U2861) );
  OAI21_X1 U20107 ( .B1(n16640), .B2(n16650), .A(n16649), .ZN(n16791) );
  NAND2_X1 U20108 ( .A1(n17218), .A2(n16728), .ZN(n16652) );
  NAND2_X1 U20109 ( .A1(n16723), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n16651) );
  OAI211_X1 U20110 ( .C1(n16791), .C2(n16733), .A(n16652), .B(n16651), .ZN(
        P2_U2862) );
  AOI21_X1 U20111 ( .B1(n9779), .B2(n16654), .A(n16653), .ZN(n16655) );
  XOR2_X1 U20112 ( .A(n16656), .B(n16655), .Z(n16798) );
  NOR2_X1 U20113 ( .A1(n17229), .A2(n16723), .ZN(n16657) );
  AOI21_X1 U20114 ( .B1(P2_EBX_REG_24__SCAN_IN), .B2(n16723), .A(n16657), .ZN(
        n16658) );
  OAI21_X1 U20115 ( .B1(n16798), .B2(n16733), .A(n16658), .ZN(P2_U2863) );
  INV_X1 U20116 ( .A(n17246), .ZN(n16664) );
  AOI21_X1 U20117 ( .B1(n16661), .B2(n16660), .A(n16659), .ZN(n16802) );
  NAND2_X1 U20118 ( .A1(n16802), .A2(n16737), .ZN(n16663) );
  NAND2_X1 U20119 ( .A1(n16723), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n16662) );
  OAI211_X1 U20120 ( .C1(n16664), .C2(n16723), .A(n16663), .B(n16662), .ZN(
        P2_U2864) );
  OR2_X1 U20121 ( .A1(n12811), .A2(n16665), .ZN(n16666) );
  NAND2_X1 U20122 ( .A1(n9766), .A2(n16666), .ZN(n17993) );
  OR2_X1 U20123 ( .A1(n16667), .A2(n16668), .ZN(n16670) );
  AND2_X1 U20124 ( .A1(n16670), .A2(n16669), .ZN(n16811) );
  AOI22_X1 U20125 ( .A1(n16811), .A2(n16737), .B1(P2_EBX_REG_22__SCAN_IN), 
        .B2(n16723), .ZN(n16671) );
  OAI21_X1 U20126 ( .B1(n17993), .B2(n16723), .A(n16671), .ZN(P2_U2865) );
  AOI21_X1 U20127 ( .B1(n16673), .B2(n16672), .A(n16667), .ZN(n16817) );
  AOI22_X1 U20128 ( .A1(n16817), .A2(n16737), .B1(P2_EBX_REG_21__SCAN_IN), 
        .B2(n16723), .ZN(n16674) );
  OAI21_X1 U20129 ( .B1(n16675), .B2(n16723), .A(n16674), .ZN(P2_U2866) );
  NAND2_X1 U20130 ( .A1(n16676), .A2(n16677), .ZN(n16678) );
  NAND2_X1 U20131 ( .A1(n16672), .A2(n16678), .ZN(n16820) );
  NAND2_X1 U20132 ( .A1(n17266), .A2(n16728), .ZN(n16680) );
  NAND2_X1 U20133 ( .A1(n16723), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n16679) );
  OAI211_X1 U20134 ( .C1(n16820), .C2(n16733), .A(n16680), .B(n16679), .ZN(
        P2_U2867) );
  NAND2_X1 U20135 ( .A1(n16681), .A2(n16682), .ZN(n16683) );
  AND2_X1 U20136 ( .A1(n16676), .A2(n16683), .ZN(n16831) );
  AOI22_X1 U20137 ( .A1(n16831), .A2(n16737), .B1(P2_EBX_REG_19__SCAN_IN), 
        .B2(n16723), .ZN(n16684) );
  OAI21_X1 U20138 ( .B1(n16685), .B2(n16723), .A(n16684), .ZN(P2_U2868) );
  OR2_X1 U20139 ( .A1(n16686), .A2(n16687), .ZN(n16688) );
  AND2_X1 U20140 ( .A1(n16681), .A2(n16688), .ZN(n16837) );
  AOI22_X1 U20141 ( .A1(n16837), .A2(n16737), .B1(P2_EBX_REG_18__SCAN_IN), 
        .B2(n16723), .ZN(n16689) );
  OAI21_X1 U20142 ( .B1(n17279), .B2(n16723), .A(n16689), .ZN(P2_U2869) );
  AND2_X1 U20143 ( .A1(n16690), .A2(n16691), .ZN(n16692) );
  NOR2_X1 U20144 ( .A1(n16686), .A2(n16692), .ZN(n16843) );
  AOI22_X1 U20145 ( .A1(n16843), .A2(n16737), .B1(P2_EBX_REG_17__SCAN_IN), 
        .B2(n16723), .ZN(n16693) );
  OAI21_X1 U20146 ( .B1(n17289), .B2(n16723), .A(n16693), .ZN(P2_U2870) );
  NAND2_X1 U20147 ( .A1(n16694), .A2(n16695), .ZN(n16696) );
  AND2_X1 U20148 ( .A1(n16690), .A2(n16696), .ZN(n16853) );
  AOI22_X1 U20149 ( .A1(n16853), .A2(n16737), .B1(P2_EBX_REG_16__SCAN_IN), 
        .B2(n16723), .ZN(n16697) );
  OAI21_X1 U20150 ( .B1(n17300), .B2(n16723), .A(n16697), .ZN(P2_U2871) );
  INV_X1 U20151 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n16705) );
  NAND2_X1 U20152 ( .A1(n16698), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n16735) );
  NAND2_X1 U20153 ( .A1(n16736), .A2(n16731), .ZN(n16725) );
  NOR2_X1 U20154 ( .A1(n16725), .A2(n16724), .ZN(n16720) );
  NAND2_X1 U20155 ( .A1(n16720), .A2(n16719), .ZN(n16718) );
  NOR2_X1 U20156 ( .A1(n16718), .A2(n16715), .ZN(n16712) );
  NAND2_X1 U20157 ( .A1(n16712), .A2(n16711), .ZN(n16710) );
  NOR2_X1 U20158 ( .A1(n16710), .A2(n16706), .ZN(n16701) );
  OAI211_X1 U20159 ( .C1(n16701), .C2(n16700), .A(n16737), .B(n16694), .ZN(
        n16704) );
  NAND2_X1 U20160 ( .A1(n16702), .A2(n16728), .ZN(n16703) );
  OAI211_X1 U20161 ( .C1(n16728), .C2(n16705), .A(n16704), .B(n16703), .ZN(
        P2_U2872) );
  XNOR2_X1 U20162 ( .A(n16710), .B(n16706), .ZN(n16709) );
  NOR2_X1 U20163 ( .A1(n16728), .A2(n11096), .ZN(n16707) );
  AOI21_X1 U20164 ( .B1(n17333), .B2(n16728), .A(n16707), .ZN(n16708) );
  OAI21_X1 U20165 ( .B1(n16709), .B2(n16733), .A(n16708), .ZN(P2_U2873) );
  OAI211_X1 U20166 ( .C1(n16712), .C2(n16711), .A(n16710), .B(n16737), .ZN(
        n16714) );
  NAND2_X1 U20167 ( .A1(n16723), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n16713) );
  OAI211_X1 U20168 ( .C1(n17344), .C2(n16723), .A(n16714), .B(n16713), .ZN(
        P2_U2874) );
  XNOR2_X1 U20169 ( .A(n16718), .B(n16715), .ZN(n16717) );
  INV_X1 U20170 ( .A(P2_EBX_REG_12__SCAN_IN), .ZN(n21819) );
  MUX2_X1 U20171 ( .A(n17358), .B(n21819), .S(n16723), .Z(n16716) );
  OAI21_X1 U20172 ( .B1(n16717), .B2(n16733), .A(n16716), .ZN(P2_U2875) );
  OAI211_X1 U20173 ( .C1(n16720), .C2(n16719), .A(n16718), .B(n16737), .ZN(
        n16722) );
  NAND2_X1 U20174 ( .A1(n16723), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n16721) );
  OAI211_X1 U20175 ( .C1(n17370), .C2(n16723), .A(n16722), .B(n16721), .ZN(
        P2_U2876) );
  XNOR2_X1 U20176 ( .A(n16725), .B(n16724), .ZN(n16730) );
  NOR2_X1 U20177 ( .A1(n16728), .A2(n16726), .ZN(n16727) );
  AOI21_X1 U20178 ( .B1(n17381), .B2(n16728), .A(n16727), .ZN(n16729) );
  OAI21_X1 U20179 ( .B1(n16730), .B2(n16733), .A(n16729), .ZN(P2_U2877) );
  XNOR2_X1 U20180 ( .A(n16736), .B(n16731), .ZN(n16734) );
  INV_X1 U20181 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n21847) );
  MUX2_X1 U20182 ( .A(n17397), .B(n21847), .S(n16723), .Z(n16732) );
  OAI21_X1 U20183 ( .B1(n16734), .B2(n16733), .A(n16732), .ZN(P2_U2878) );
  INV_X1 U20184 ( .A(n16735), .ZN(n16740) );
  INV_X1 U20185 ( .A(n16736), .ZN(n16738) );
  OAI211_X1 U20186 ( .C1(n16740), .C2(n16739), .A(n16738), .B(n16737), .ZN(
        n16742) );
  NAND2_X1 U20187 ( .A1(n16723), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n16741) );
  OAI211_X1 U20188 ( .C1(n17090), .C2(n16723), .A(n16742), .B(n16741), .ZN(
        P2_U2879) );
  INV_X1 U20189 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n16747) );
  AND2_X1 U20190 ( .A1(n16744), .A2(n16743), .ZN(n16846) );
  AOI22_X1 U20191 ( .A1(n16846), .A2(n16745), .B1(P2_EAX_REG_30__SCAN_IN), 
        .B2(n16867), .ZN(n16746) );
  OAI21_X1 U20192 ( .B1(n16850), .B2(n16747), .A(n16746), .ZN(n16748) );
  INV_X1 U20193 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n16749) );
  NOR2_X1 U20194 ( .A1(n12797), .A2(n16749), .ZN(n16750) );
  OAI21_X1 U20195 ( .B1(n16752), .B2(n16855), .A(n16751), .ZN(n16753) );
  INV_X1 U20196 ( .A(n16753), .ZN(n16754) );
  OAI21_X1 U20197 ( .B1(n16755), .B2(n16872), .A(n16754), .ZN(P2_U2889) );
  INV_X1 U20198 ( .A(n17169), .ZN(n16763) );
  NAND3_X1 U20199 ( .A1(n9724), .A2(n16852), .A3(n16756), .ZN(n16762) );
  INV_X1 U20200 ( .A(BUF2_REG_29__SCAN_IN), .ZN(n16759) );
  AOI22_X1 U20201 ( .A1(n16846), .A2(n16757), .B1(P2_EAX_REG_29__SCAN_IN), 
        .B2(n16867), .ZN(n16758) );
  OAI21_X1 U20202 ( .B1(n16850), .B2(n16759), .A(n16758), .ZN(n16760) );
  AOI21_X1 U20203 ( .B1(n16845), .B2(BUF1_REG_29__SCAN_IN), .A(n16760), .ZN(
        n16761) );
  OAI211_X1 U20204 ( .C1(n16763), .C2(n16855), .A(n16762), .B(n16761), .ZN(
        P2_U2890) );
  INV_X1 U20205 ( .A(BUF2_REG_28__SCAN_IN), .ZN(n16767) );
  NAND2_X1 U20206 ( .A1(n16845), .A2(BUF1_REG_28__SCAN_IN), .ZN(n16766) );
  AOI22_X1 U20207 ( .A1(n16846), .A2(n16764), .B1(P2_EAX_REG_28__SCAN_IN), 
        .B2(n16867), .ZN(n16765) );
  OAI211_X1 U20208 ( .C1(n16850), .C2(n16767), .A(n16766), .B(n16765), .ZN(
        n16768) );
  AOI21_X1 U20209 ( .B1(n17176), .B2(n16868), .A(n16768), .ZN(n16769) );
  OAI21_X1 U20210 ( .B1(n16770), .B2(n16872), .A(n16769), .ZN(P2_U2891) );
  INV_X1 U20211 ( .A(BUF2_REG_27__SCAN_IN), .ZN(n16774) );
  AOI22_X1 U20212 ( .A1(n16846), .A2(n16772), .B1(P2_EAX_REG_27__SCAN_IN), 
        .B2(n16867), .ZN(n16773) );
  OAI21_X1 U20213 ( .B1(n16850), .B2(n16774), .A(n16773), .ZN(n16775) );
  AOI21_X1 U20214 ( .B1(n16845), .B2(BUF1_REG_27__SCAN_IN), .A(n16775), .ZN(
        n16776) );
  OAI211_X1 U20215 ( .C1(n17193), .C2(n16855), .A(n16777), .B(n16776), .ZN(
        P2_U2892) );
  INV_X1 U20216 ( .A(BUF2_REG_26__SCAN_IN), .ZN(n16780) );
  AOI22_X1 U20217 ( .A1(n16846), .A2(n16778), .B1(P2_EAX_REG_26__SCAN_IN), 
        .B2(n16867), .ZN(n16779) );
  OAI21_X1 U20218 ( .B1(n16850), .B2(n16780), .A(n16779), .ZN(n16782) );
  NOR2_X1 U20219 ( .A1(n17198), .A2(n16855), .ZN(n16781) );
  AOI211_X1 U20220 ( .C1(n16845), .C2(BUF1_REG_26__SCAN_IN), .A(n16782), .B(
        n16781), .ZN(n16783) );
  OAI21_X1 U20221 ( .B1(n16784), .B2(n16872), .A(n16783), .ZN(P2_U2893) );
  INV_X1 U20222 ( .A(BUF2_REG_25__SCAN_IN), .ZN(n16787) );
  AOI22_X1 U20223 ( .A1(n16846), .A2(n16785), .B1(P2_EAX_REG_25__SCAN_IN), 
        .B2(n16867), .ZN(n16786) );
  OAI21_X1 U20224 ( .B1(n16850), .B2(n16787), .A(n16786), .ZN(n16789) );
  NOR2_X1 U20225 ( .A1(n17211), .A2(n16855), .ZN(n16788) );
  AOI211_X1 U20226 ( .C1(n16845), .C2(BUF1_REG_25__SCAN_IN), .A(n16789), .B(
        n16788), .ZN(n16790) );
  OAI21_X1 U20227 ( .B1(n16872), .B2(n16791), .A(n16790), .ZN(P2_U2894) );
  INV_X1 U20228 ( .A(BUF2_REG_24__SCAN_IN), .ZN(n16795) );
  NAND2_X1 U20229 ( .A1(n16845), .A2(BUF1_REG_24__SCAN_IN), .ZN(n16794) );
  AOI22_X1 U20230 ( .A1(n16846), .A2(n16792), .B1(P2_EAX_REG_24__SCAN_IN), 
        .B2(n16867), .ZN(n16793) );
  OAI211_X1 U20231 ( .C1(n16850), .C2(n16795), .A(n16794), .B(n16793), .ZN(
        n16796) );
  AOI21_X1 U20232 ( .B1(n17233), .B2(n16868), .A(n16796), .ZN(n16797) );
  OAI21_X1 U20233 ( .B1(n16798), .B2(n16872), .A(n16797), .ZN(P2_U2895) );
  INV_X1 U20234 ( .A(BUF2_REG_23__SCAN_IN), .ZN(n16800) );
  AOI22_X1 U20235 ( .A1(n16846), .A2(n17587), .B1(P2_EAX_REG_23__SCAN_IN), 
        .B2(n16867), .ZN(n16799) );
  OAI21_X1 U20236 ( .B1(n16850), .B2(n16800), .A(n16799), .ZN(n16801) );
  AOI21_X1 U20237 ( .B1(n16845), .B2(BUF1_REG_23__SCAN_IN), .A(n16801), .ZN(
        n16804) );
  NAND2_X1 U20238 ( .A1(n16802), .A2(n16852), .ZN(n16803) );
  OAI211_X1 U20239 ( .C1(n17236), .C2(n16855), .A(n16804), .B(n16803), .ZN(
        P2_U2896) );
  OR2_X1 U20240 ( .A1(n12763), .A2(n16805), .ZN(n16806) );
  NAND2_X1 U20241 ( .A1(n16079), .A2(n16806), .ZN(n17992) );
  INV_X1 U20242 ( .A(BUF2_REG_22__SCAN_IN), .ZN(n16809) );
  NAND2_X1 U20243 ( .A1(n16845), .A2(BUF1_REG_22__SCAN_IN), .ZN(n16808) );
  AOI22_X1 U20244 ( .A1(n16846), .A2(n17536), .B1(P2_EAX_REG_22__SCAN_IN), 
        .B2(n16867), .ZN(n16807) );
  OAI211_X1 U20245 ( .C1(n16850), .C2(n16809), .A(n16808), .B(n16807), .ZN(
        n16810) );
  AOI21_X1 U20246 ( .B1(n16811), .B2(n16852), .A(n16810), .ZN(n16812) );
  OAI21_X1 U20247 ( .B1(n17992), .B2(n16855), .A(n16812), .ZN(P2_U2897) );
  INV_X1 U20248 ( .A(n16813), .ZN(n16819) );
  INV_X1 U20249 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n17721) );
  NAND2_X1 U20250 ( .A1(n16845), .A2(BUF1_REG_21__SCAN_IN), .ZN(n16815) );
  AOI22_X1 U20251 ( .A1(n16846), .A2(n17531), .B1(P2_EAX_REG_21__SCAN_IN), 
        .B2(n16867), .ZN(n16814) );
  OAI211_X1 U20252 ( .C1(n16850), .C2(n17721), .A(n16815), .B(n16814), .ZN(
        n16816) );
  AOI21_X1 U20253 ( .B1(n16817), .B2(n16852), .A(n16816), .ZN(n16818) );
  OAI21_X1 U20254 ( .B1(n16819), .B2(n16855), .A(n16818), .ZN(P2_U2898) );
  INV_X1 U20255 ( .A(n16820), .ZN(n16825) );
  INV_X1 U20256 ( .A(BUF2_REG_20__SCAN_IN), .ZN(n16823) );
  NAND2_X1 U20257 ( .A1(n16845), .A2(BUF1_REG_20__SCAN_IN), .ZN(n16822) );
  AOI22_X1 U20258 ( .A1(n16846), .A2(n17574), .B1(P2_EAX_REG_20__SCAN_IN), 
        .B2(n16867), .ZN(n16821) );
  OAI211_X1 U20259 ( .C1(n16850), .C2(n16823), .A(n16822), .B(n16821), .ZN(
        n16824) );
  AOI21_X1 U20260 ( .B1(n16825), .B2(n16852), .A(n16824), .ZN(n16826) );
  OAI21_X1 U20261 ( .B1(n17268), .B2(n16855), .A(n16826), .ZN(P2_U2899) );
  INV_X1 U20262 ( .A(BUF2_REG_19__SCAN_IN), .ZN(n17727) );
  NAND2_X1 U20263 ( .A1(n16845), .A2(BUF1_REG_19__SCAN_IN), .ZN(n16829) );
  AOI22_X1 U20264 ( .A1(n16846), .A2(n17569), .B1(P2_EAX_REG_19__SCAN_IN), 
        .B2(n16867), .ZN(n16828) );
  OAI211_X1 U20265 ( .C1(n16850), .C2(n17727), .A(n16829), .B(n16828), .ZN(
        n16830) );
  AOI21_X1 U20266 ( .B1(n16831), .B2(n16852), .A(n16830), .ZN(n16832) );
  OAI21_X1 U20267 ( .B1(n14783), .B2(n16855), .A(n16832), .ZN(P2_U2900) );
  INV_X1 U20268 ( .A(BUF2_REG_18__SCAN_IN), .ZN(n16835) );
  NAND2_X1 U20269 ( .A1(n16845), .A2(BUF1_REG_18__SCAN_IN), .ZN(n16834) );
  AOI22_X1 U20270 ( .A1(n16846), .A2(n17563), .B1(P2_EAX_REG_18__SCAN_IN), 
        .B2(n16867), .ZN(n16833) );
  OAI211_X1 U20271 ( .C1(n16850), .C2(n16835), .A(n16834), .B(n16833), .ZN(
        n16836) );
  AOI21_X1 U20272 ( .B1(n16837), .B2(n16852), .A(n16836), .ZN(n16838) );
  OAI21_X1 U20273 ( .B1(n17273), .B2(n16855), .A(n16838), .ZN(P2_U2901) );
  INV_X1 U20274 ( .A(BUF2_REG_17__SCAN_IN), .ZN(n16841) );
  NAND2_X1 U20275 ( .A1(n16845), .A2(BUF1_REG_17__SCAN_IN), .ZN(n16840) );
  AOI22_X1 U20276 ( .A1(n16846), .A2(n17558), .B1(P2_EAX_REG_17__SCAN_IN), 
        .B2(n16867), .ZN(n16839) );
  OAI211_X1 U20277 ( .C1(n16850), .C2(n16841), .A(n16840), .B(n16839), .ZN(
        n16842) );
  AOI21_X1 U20278 ( .B1(n16843), .B2(n16852), .A(n16842), .ZN(n16844) );
  OAI21_X1 U20279 ( .B1(n17287), .B2(n16855), .A(n16844), .ZN(P2_U2902) );
  INV_X1 U20280 ( .A(BUF2_REG_16__SCAN_IN), .ZN(n16849) );
  NAND2_X1 U20281 ( .A1(n16845), .A2(BUF1_REG_16__SCAN_IN), .ZN(n16848) );
  AOI22_X1 U20282 ( .A1(n16846), .A2(n17524), .B1(P2_EAX_REG_16__SCAN_IN), 
        .B2(n16867), .ZN(n16847) );
  OAI211_X1 U20283 ( .C1(n16850), .C2(n16849), .A(n16848), .B(n16847), .ZN(
        n16851) );
  AOI21_X1 U20284 ( .B1(n16853), .B2(n16852), .A(n16851), .ZN(n16854) );
  OAI21_X1 U20285 ( .B1(n16856), .B2(n16855), .A(n16854), .ZN(P2_U2903) );
  INV_X1 U20286 ( .A(n17440), .ZN(n16865) );
  AOI21_X1 U20287 ( .B1(n18090), .B2(n20535), .A(n16857), .ZN(n16861) );
  NAND2_X1 U20288 ( .A1(n14561), .A2(n16858), .ZN(n16859) );
  AND2_X1 U20289 ( .A1(n16860), .A2(n16859), .ZN(n20263) );
  NOR2_X1 U20290 ( .A1(n16861), .A2(n20263), .ZN(n16866) );
  OR3_X1 U20291 ( .A1(n16866), .A2(n20198), .A3(n16872), .ZN(n16863) );
  AOI22_X1 U20292 ( .A1(n16869), .A2(n17531), .B1(P2_EAX_REG_5__SCAN_IN), .B2(
        n16867), .ZN(n16862) );
  OAI211_X1 U20293 ( .C1(n16865), .C2(n16864), .A(n16863), .B(n16862), .ZN(
        P2_U2914) );
  XNOR2_X1 U20294 ( .A(n16866), .B(n20198), .ZN(n16873) );
  AOI22_X1 U20295 ( .A1(n20263), .A2(n16868), .B1(P2_EAX_REG_4__SCAN_IN), .B2(
        n16867), .ZN(n16871) );
  NAND2_X1 U20296 ( .A1(n16869), .A2(n17574), .ZN(n16870) );
  OAI211_X1 U20297 ( .C1(n16873), .C2(n16872), .A(n16871), .B(n16870), .ZN(
        P2_U2915) );
  OAI21_X1 U20298 ( .B1(n18060), .B2(n16875), .A(n16874), .ZN(n16876) );
  AOI21_X1 U20299 ( .B1(n16877), .B2(n18063), .A(n16876), .ZN(n16878) );
  OAI21_X1 U20300 ( .B1(n16879), .B2(n17126), .A(n16878), .ZN(n16880) );
  OAI21_X1 U20301 ( .B1(n16883), .B2(n20249), .A(n16882), .ZN(P2_U2984) );
  INV_X1 U20302 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n20871) );
  NOR2_X1 U20303 ( .A1(n17136), .A2(n20871), .ZN(n17161) );
  NOR2_X1 U20304 ( .A1(n16887), .A2(n17146), .ZN(n16888) );
  AOI211_X1 U20305 ( .C1(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .C2(n20247), .A(
        n17161), .B(n16888), .ZN(n16889) );
  OAI21_X1 U20306 ( .B1(n17160), .B2(n17126), .A(n16889), .ZN(n16890) );
  AOI21_X1 U20307 ( .B1(n17155), .B2(n17172), .A(n16890), .ZN(n16891) );
  OAI21_X1 U20308 ( .B1(n17175), .B2(n20249), .A(n16891), .ZN(P2_U2985) );
  INV_X1 U20309 ( .A(n16892), .ZN(n16893) );
  XNOR2_X1 U20310 ( .A(n16894), .B(n17188), .ZN(n16895) );
  NAND2_X1 U20311 ( .A1(n11487), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n17186) );
  NAND2_X1 U20312 ( .A1(n20247), .A2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16897) );
  OAI211_X1 U20313 ( .C1(n16898), .C2(n17146), .A(n17186), .B(n16897), .ZN(
        n16901) );
  NOR2_X1 U20314 ( .A1(n16899), .A2(n17126), .ZN(n16900) );
  INV_X1 U20315 ( .A(n16916), .ZN(n16914) );
  NAND2_X1 U20316 ( .A1(n16917), .A2(n16914), .ZN(n16903) );
  XOR2_X1 U20317 ( .A(n16904), .B(n16903), .Z(n17210) );
  NOR2_X1 U20318 ( .A1(n17136), .A2(n16906), .ZN(n17201) );
  NOR2_X1 U20319 ( .A1(n16907), .A2(n17146), .ZN(n16908) );
  AOI211_X1 U20320 ( .C1(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .C2(n20247), .A(
        n17201), .B(n16908), .ZN(n16909) );
  OAI21_X1 U20321 ( .B1(n17205), .B2(n17126), .A(n16909), .ZN(n16910) );
  AOI21_X1 U20322 ( .B1(n17155), .B2(n17208), .A(n16910), .ZN(n16911) );
  OAI21_X1 U20323 ( .B1(n17210), .B2(n20249), .A(n16911), .ZN(P2_U2988) );
  AND2_X1 U20324 ( .A1(n16914), .A2(n16913), .ZN(n16915) );
  OAI22_X1 U20325 ( .A1(n16917), .A2(n16916), .B1(n16912), .B2(n16915), .ZN(
        n17222) );
  NAND2_X1 U20326 ( .A1(n11487), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n17212) );
  NAND2_X1 U20327 ( .A1(n20247), .A2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n16918) );
  OAI211_X1 U20328 ( .C1(n16919), .C2(n17146), .A(n17212), .B(n16918), .ZN(
        n16920) );
  AOI21_X1 U20329 ( .B1(n17218), .B2(n20252), .A(n16920), .ZN(n16922) );
  NAND2_X1 U20330 ( .A1(n16923), .A2(n17214), .ZN(n17219) );
  OAI211_X1 U20331 ( .C1(n17222), .C2(n20249), .A(n16922), .B(n16921), .ZN(
        P2_U2989) );
  OAI21_X1 U20332 ( .B1(n16940), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n16923), .ZN(n17235) );
  INV_X1 U20333 ( .A(n17229), .ZN(n16930) );
  NAND2_X1 U20334 ( .A1(n18058), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n17228) );
  NAND2_X1 U20335 ( .A1(n20247), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n16924) );
  OAI211_X1 U20336 ( .C1(n16925), .C2(n17146), .A(n17228), .B(n16924), .ZN(
        n16929) );
  XNOR2_X1 U20337 ( .A(n16927), .B(n10602), .ZN(n16928) );
  OAI21_X1 U20338 ( .B1(n20256), .B2(n17235), .A(n9809), .ZN(P2_U2990) );
  NOR2_X1 U20339 ( .A1(n16932), .A2(n16933), .ZN(n16948) );
  OAI21_X1 U20340 ( .B1(n16948), .B2(n16946), .A(n16934), .ZN(n16935) );
  XOR2_X1 U20341 ( .A(n16936), .B(n16935), .Z(n17249) );
  NAND2_X1 U20342 ( .A1(n11487), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n17242) );
  NAND2_X1 U20343 ( .A1(n20247), .A2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n16937) );
  OAI211_X1 U20344 ( .C1(n16938), .C2(n17146), .A(n17242), .B(n16937), .ZN(
        n16939) );
  AOI21_X1 U20345 ( .B1(n17246), .B2(n20252), .A(n16939), .ZN(n16942) );
  OAI211_X1 U20346 ( .C1(n17249), .C2(n20249), .A(n16942), .B(n16941), .ZN(
        P2_U2991) );
  OAI21_X1 U20347 ( .B1(n16944), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n16943), .ZN(n17258) );
  NOR2_X1 U20348 ( .A1(n16946), .A2(n16945), .ZN(n16947) );
  XNOR2_X1 U20349 ( .A(n16948), .B(n16947), .ZN(n17256) );
  NOR2_X1 U20350 ( .A1(n17136), .A2(n16949), .ZN(n17251) );
  NOR2_X1 U20351 ( .A1(n17995), .A2(n17146), .ZN(n16950) );
  AOI211_X1 U20352 ( .C1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .C2(n20247), .A(
        n17251), .B(n16950), .ZN(n16951) );
  OAI21_X1 U20353 ( .B1(n17993), .B2(n17126), .A(n16951), .ZN(n16952) );
  AOI21_X1 U20354 ( .B1(n17256), .B2(n18070), .A(n16952), .ZN(n16953) );
  OAI21_X1 U20355 ( .B1(n20256), .B2(n17258), .A(n16953), .ZN(P2_U2992) );
  AOI21_X1 U20356 ( .B1(n20247), .B2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n16954), .ZN(n16955) );
  OAI21_X1 U20357 ( .B1(n16956), .B2(n17146), .A(n16955), .ZN(n16957) );
  NAND2_X1 U20358 ( .A1(n16962), .A2(n16961), .ZN(n16963) );
  XNOR2_X1 U20359 ( .A(n16964), .B(n16963), .ZN(n17272) );
  NAND2_X1 U20360 ( .A1(n11487), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n17261) );
  NAND2_X1 U20361 ( .A1(n20247), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n16965) );
  OAI211_X1 U20362 ( .C1(n16966), .C2(n17146), .A(n17261), .B(n16965), .ZN(
        n16967) );
  AOI21_X1 U20363 ( .B1(n17266), .B2(n20252), .A(n16967), .ZN(n16971) );
  NAND2_X1 U20364 ( .A1(n17270), .A2(n17155), .ZN(n16970) );
  OAI211_X1 U20365 ( .C1(n17272), .C2(n20249), .A(n16971), .B(n16970), .ZN(
        P2_U2994) );
  NAND2_X1 U20366 ( .A1(n16974), .A2(n16973), .ZN(n16975) );
  XNOR2_X1 U20367 ( .A(n16972), .B(n16975), .ZN(n17284) );
  NOR2_X1 U20368 ( .A1(n17136), .A2(n20855), .ZN(n17276) );
  NOR2_X1 U20369 ( .A1(n16977), .A2(n17146), .ZN(n16978) );
  AOI211_X1 U20370 ( .C1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(n20247), .A(
        n17276), .B(n16978), .ZN(n16979) );
  OAI21_X1 U20371 ( .B1(n17279), .B2(n17126), .A(n16979), .ZN(n16980) );
  AOI21_X1 U20372 ( .B1(n17282), .B2(n17155), .A(n16980), .ZN(n16981) );
  OAI21_X1 U20373 ( .B1(n17284), .B2(n20249), .A(n16981), .ZN(P2_U2996) );
  XNOR2_X1 U20374 ( .A(n17295), .B(n17292), .ZN(n16988) );
  INV_X1 U20375 ( .A(n17289), .ZN(n16987) );
  NAND2_X1 U20376 ( .A1(n11487), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n17288) );
  NAND2_X1 U20377 ( .A1(n20247), .A2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n16982) );
  OAI211_X1 U20378 ( .C1(n17146), .C2(n16983), .A(n17288), .B(n16982), .ZN(
        n16986) );
  XNOR2_X1 U20379 ( .A(n16989), .B(n16990), .ZN(n17309) );
  NAND2_X1 U20380 ( .A1(n18058), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n17299) );
  NAND2_X1 U20381 ( .A1(n20247), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n16991) );
  OAI211_X1 U20382 ( .C1(n17146), .C2(n16992), .A(n17299), .B(n16991), .ZN(
        n16994) );
  AOI21_X1 U20383 ( .B1(n17301), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16993) );
  OAI21_X1 U20384 ( .B1(n20249), .B2(n17309), .A(n16996), .ZN(P2_U2998) );
  XNOR2_X1 U20385 ( .A(n16997), .B(n17315), .ZN(n17323) );
  NAND2_X1 U20386 ( .A1(n16999), .A2(n16998), .ZN(n17000) );
  XNOR2_X1 U20387 ( .A(n17001), .B(n17000), .ZN(n17310) );
  NAND2_X1 U20388 ( .A1(n11487), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n17311) );
  OAI21_X1 U20389 ( .B1(n18060), .B2(n17002), .A(n17311), .ZN(n17003) );
  AOI21_X1 U20390 ( .B1(n18063), .B2(n17004), .A(n17003), .ZN(n17005) );
  OAI21_X1 U20391 ( .B1(n17317), .B2(n17126), .A(n17005), .ZN(n17006) );
  AOI21_X1 U20392 ( .B1(n17310), .B2(n18070), .A(n17006), .ZN(n17007) );
  OAI21_X1 U20393 ( .B1(n20256), .B2(n17323), .A(n17007), .ZN(P2_U2999) );
  NAND2_X1 U20394 ( .A1(n17009), .A2(n17008), .ZN(n17027) );
  INV_X1 U20395 ( .A(n17025), .ZN(n17010) );
  AOI21_X1 U20396 ( .B1(n17027), .B2(n17024), .A(n17010), .ZN(n17014) );
  NAND2_X1 U20397 ( .A1(n17012), .A2(n17011), .ZN(n17013) );
  XNOR2_X1 U20398 ( .A(n17014), .B(n17013), .ZN(n17340) );
  NAND2_X1 U20399 ( .A1(n17324), .A2(n17155), .ZN(n17020) );
  NOR2_X1 U20400 ( .A1(n17136), .A2(n20848), .ZN(n17332) );
  AOI21_X1 U20401 ( .B1(n20247), .B2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n17332), .ZN(n17016) );
  OAI21_X1 U20402 ( .B1(n17146), .B2(n17017), .A(n17016), .ZN(n17018) );
  AOI21_X1 U20403 ( .B1(n17333), .B2(n20252), .A(n17018), .ZN(n17019) );
  OAI211_X1 U20404 ( .C1(n17340), .C2(n20249), .A(n17020), .B(n17019), .ZN(
        P2_U3000) );
  NAND2_X1 U20405 ( .A1(n17023), .A2(n17022), .ZN(n17353) );
  NAND2_X1 U20406 ( .A1(n17025), .A2(n17024), .ZN(n17026) );
  XNOR2_X1 U20407 ( .A(n17027), .B(n17026), .ZN(n17351) );
  NOR2_X1 U20408 ( .A1(n17344), .A2(n17126), .ZN(n17031) );
  NAND2_X1 U20409 ( .A1(n11487), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n17343) );
  NAND2_X1 U20410 ( .A1(n20247), .A2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n17028) );
  OAI211_X1 U20411 ( .C1(n17146), .C2(n17029), .A(n17343), .B(n17028), .ZN(
        n17030) );
  AOI211_X1 U20412 ( .C1(n17351), .C2(n18070), .A(n17031), .B(n17030), .ZN(
        n17032) );
  OAI21_X1 U20413 ( .B1(n17353), .B2(n20256), .A(n17032), .ZN(P2_U3001) );
  XNOR2_X1 U20414 ( .A(n9771), .B(n17327), .ZN(n17365) );
  NAND2_X1 U20415 ( .A1(n17033), .A2(n17043), .ZN(n17036) );
  XNOR2_X1 U20416 ( .A(n17034), .B(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n17035) );
  XNOR2_X1 U20417 ( .A(n17036), .B(n17035), .ZN(n17362) );
  NAND2_X1 U20418 ( .A1(n11487), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n17357) );
  OAI21_X1 U20419 ( .B1(n18060), .B2(n17037), .A(n17357), .ZN(n17038) );
  AOI21_X1 U20420 ( .B1(n18063), .B2(n17039), .A(n17038), .ZN(n17040) );
  OAI21_X1 U20421 ( .B1(n17358), .B2(n17126), .A(n17040), .ZN(n17041) );
  AOI21_X1 U20422 ( .B1(n17362), .B2(n18070), .A(n17041), .ZN(n17042) );
  OAI21_X1 U20423 ( .B1(n17365), .B2(n20256), .A(n17042), .ZN(P2_U3002) );
  OAI21_X1 U20424 ( .B1(n17060), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n9771), .ZN(n17379) );
  INV_X1 U20425 ( .A(n17043), .ZN(n17044) );
  NOR2_X1 U20426 ( .A1(n17045), .A2(n17044), .ZN(n17047) );
  XOR2_X1 U20427 ( .A(n17047), .B(n17046), .Z(n17376) );
  NAND2_X1 U20428 ( .A1(n11487), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n17369) );
  OAI21_X1 U20429 ( .B1(n18060), .B2(n17048), .A(n17369), .ZN(n17049) );
  AOI21_X1 U20430 ( .B1(n18063), .B2(n17050), .A(n17049), .ZN(n17051) );
  OAI21_X1 U20431 ( .B1(n17370), .B2(n17126), .A(n17051), .ZN(n17052) );
  AOI21_X1 U20432 ( .B1(n17376), .B2(n18070), .A(n17052), .ZN(n17053) );
  OAI21_X1 U20433 ( .B1(n17379), .B2(n20256), .A(n17053), .ZN(P2_U3003) );
  NAND2_X1 U20434 ( .A1(n17055), .A2(n17054), .ZN(n17059) );
  AND2_X1 U20435 ( .A1(n17057), .A2(n17056), .ZN(n17068) );
  NAND2_X1 U20436 ( .A1(n17068), .A2(n17069), .ZN(n17067) );
  NAND2_X1 U20437 ( .A1(n17067), .A2(n17071), .ZN(n17058) );
  XOR2_X1 U20438 ( .A(n17059), .B(n17058), .Z(n17392) );
  NAND2_X1 U20439 ( .A1(n17380), .A2(n17155), .ZN(n17065) );
  NAND2_X1 U20440 ( .A1(n11487), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n17382) );
  NAND2_X1 U20441 ( .A1(n20247), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n17061) );
  OAI211_X1 U20442 ( .C1(n17146), .C2(n17062), .A(n17382), .B(n17061), .ZN(
        n17063) );
  AOI21_X1 U20443 ( .B1(n17381), .B2(n20252), .A(n17063), .ZN(n17064) );
  OAI211_X1 U20444 ( .C1(n17392), .C2(n20249), .A(n17065), .B(n17064), .ZN(
        P2_U3004) );
  INV_X1 U20445 ( .A(n17067), .ZN(n17072) );
  AOI21_X1 U20446 ( .B1(n17069), .B2(n17071), .A(n17068), .ZN(n17070) );
  AOI21_X1 U20447 ( .B1(n17072), .B2(n17071), .A(n17070), .ZN(n17401) );
  NOR2_X1 U20448 ( .A1(n17397), .A2(n17126), .ZN(n17076) );
  NAND2_X1 U20449 ( .A1(n18058), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n17396) );
  NAND2_X1 U20450 ( .A1(n20247), .A2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n17073) );
  OAI211_X1 U20451 ( .C1(n17146), .C2(n17074), .A(n17396), .B(n17073), .ZN(
        n17075) );
  AOI211_X1 U20452 ( .C1(n17401), .C2(n18070), .A(n17076), .B(n17075), .ZN(
        n17077) );
  OAI21_X1 U20453 ( .B1(n17404), .B2(n20256), .A(n17077), .ZN(P2_U3005) );
  XNOR2_X1 U20454 ( .A(n17078), .B(n17079), .ZN(n17416) );
  XNOR2_X1 U20455 ( .A(n17080), .B(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n17098) );
  INV_X1 U20456 ( .A(n17081), .ZN(n17083) );
  OAI21_X1 U20457 ( .B1(n17098), .B2(n17083), .A(n17082), .ZN(n18065) );
  INV_X1 U20458 ( .A(n17084), .ZN(n18066) );
  NOR2_X1 U20459 ( .A1(n18065), .A2(n18066), .ZN(n18064) );
  NOR2_X1 U20460 ( .A1(n18064), .A2(n18068), .ZN(n17089) );
  INV_X1 U20461 ( .A(n17085), .ZN(n17087) );
  NAND2_X1 U20462 ( .A1(n17087), .A2(n17086), .ZN(n17088) );
  XNOR2_X1 U20463 ( .A(n17089), .B(n17088), .ZN(n17414) );
  NOR2_X1 U20464 ( .A1(n17090), .A2(n17126), .ZN(n17094) );
  NAND2_X1 U20465 ( .A1(n11487), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n17406) );
  NAND2_X1 U20466 ( .A1(n20247), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n17091) );
  OAI211_X1 U20467 ( .C1(n17146), .C2(n17092), .A(n17406), .B(n17091), .ZN(
        n17093) );
  AOI211_X1 U20468 ( .C1(n17414), .C2(n18070), .A(n17094), .B(n17093), .ZN(
        n17095) );
  OAI21_X1 U20469 ( .B1(n17416), .B2(n20256), .A(n17095), .ZN(P2_U3006) );
  XNOR2_X1 U20470 ( .A(n17097), .B(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n17430) );
  XNOR2_X1 U20471 ( .A(n17081), .B(n17098), .ZN(n17428) );
  NAND2_X1 U20472 ( .A1(n17423), .A2(n20252), .ZN(n17100) );
  NOR2_X1 U20473 ( .A1(n17136), .A2(n20835), .ZN(n17422) );
  AOI21_X1 U20474 ( .B1(n20247), .B2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n17422), .ZN(n17099) );
  OAI211_X1 U20475 ( .C1(n17101), .C2(n17146), .A(n17100), .B(n17099), .ZN(
        n17102) );
  AOI21_X1 U20476 ( .B1(n17428), .B2(n18070), .A(n17102), .ZN(n17103) );
  OAI21_X1 U20477 ( .B1(n17430), .B2(n20256), .A(n17103), .ZN(P2_U3008) );
  XNOR2_X1 U20478 ( .A(n17104), .B(n17105), .ZN(n17444) );
  AOI21_X1 U20479 ( .B1(n17109), .B2(n17107), .A(n10267), .ZN(n17108) );
  AOI21_X1 U20480 ( .B1(n17106), .B2(n17109), .A(n17108), .ZN(n17431) );
  NAND2_X1 U20481 ( .A1(n17431), .A2(n17155), .ZN(n17115) );
  INV_X1 U20482 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17110) );
  NAND2_X1 U20483 ( .A1(n18058), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n17432) );
  OAI21_X1 U20484 ( .B1(n18060), .B2(n17110), .A(n17432), .ZN(n17112) );
  NOR2_X1 U20485 ( .A1(n17434), .A2(n17126), .ZN(n17111) );
  AOI211_X1 U20486 ( .C1(n17113), .C2(n18063), .A(n17112), .B(n17111), .ZN(
        n17114) );
  OAI211_X1 U20487 ( .C1(n17444), .C2(n20249), .A(n17115), .B(n17114), .ZN(
        P2_U3009) );
  NAND2_X1 U20488 ( .A1(n17116), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n17131) );
  NOR2_X1 U20489 ( .A1(n17116), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n17130) );
  AOI21_X1 U20490 ( .B1(n17117), .B2(n17131), .A(n17130), .ZN(n17119) );
  XNOR2_X1 U20491 ( .A(n20193), .B(n20264), .ZN(n17118) );
  XNOR2_X1 U20492 ( .A(n17119), .B(n17118), .ZN(n20268) );
  INV_X1 U20493 ( .A(n20268), .ZN(n17129) );
  XNOR2_X1 U20494 ( .A(n17121), .B(n20264), .ZN(n17122) );
  XNOR2_X1 U20495 ( .A(n17120), .B(n17122), .ZN(n20266) );
  NAND2_X1 U20496 ( .A1(n11487), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n20269) );
  OAI21_X1 U20497 ( .B1(n18060), .B2(n17123), .A(n20269), .ZN(n17124) );
  AOI21_X1 U20498 ( .B1(n18063), .B2(n20201), .A(n17124), .ZN(n17125) );
  OAI21_X1 U20499 ( .B1(n20258), .B2(n17126), .A(n17125), .ZN(n17127) );
  AOI21_X1 U20500 ( .B1(n20266), .B2(n17155), .A(n17127), .ZN(n17128) );
  OAI21_X1 U20501 ( .B1(n17129), .B2(n20249), .A(n17128), .ZN(P2_U3010) );
  INV_X1 U20502 ( .A(n17130), .ZN(n17132) );
  NAND2_X1 U20503 ( .A1(n17132), .A2(n17131), .ZN(n17134) );
  XNOR2_X1 U20504 ( .A(n17134), .B(n17133), .ZN(n18093) );
  INV_X1 U20505 ( .A(n18093), .ZN(n17143) );
  NOR2_X1 U20506 ( .A1(n17136), .A2(n17135), .ZN(n18087) );
  AOI21_X1 U20507 ( .B1(n20247), .B2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n18087), .ZN(n17137) );
  OAI21_X1 U20508 ( .B1(n17146), .B2(n17138), .A(n17137), .ZN(n17139) );
  AOI21_X1 U20509 ( .B1(n10798), .B2(n20252), .A(n17139), .ZN(n17142) );
  NAND3_X1 U20510 ( .A1(n18086), .A2(n17155), .A3(n18085), .ZN(n17141) );
  OAI211_X1 U20511 ( .C1(n17143), .C2(n20249), .A(n17142), .B(n17141), .ZN(
        P2_U3011) );
  NAND2_X1 U20512 ( .A1(n20281), .A2(n20252), .ZN(n17159) );
  NAND2_X1 U20513 ( .A1(n11487), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n20282) );
  NAND2_X1 U20514 ( .A1(n20247), .A2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n17144) );
  OAI211_X1 U20515 ( .C1(n17146), .C2(n17145), .A(n20282), .B(n17144), .ZN(
        n17147) );
  INV_X1 U20516 ( .A(n17147), .ZN(n17158) );
  OAI21_X1 U20517 ( .B1(n17150), .B2(n17149), .A(n17148), .ZN(n17151) );
  INV_X1 U20518 ( .A(n17151), .ZN(n20278) );
  NAND2_X1 U20519 ( .A1(n20278), .A2(n18070), .ZN(n17157) );
  INV_X1 U20520 ( .A(n17152), .ZN(n17153) );
  NAND2_X1 U20521 ( .A1(n17154), .A2(n17153), .ZN(n20286) );
  NAND3_X1 U20522 ( .A1(n20287), .A2(n17155), .A3(n20286), .ZN(n17156) );
  NAND4_X1 U20523 ( .A1(n17159), .A2(n17158), .A3(n17157), .A4(n17156), .ZN(
        P2_U3012) );
  AOI21_X1 U20524 ( .B1(n17163), .B2(n17162), .A(n17161), .ZN(n17167) );
  INV_X1 U20525 ( .A(n17178), .ZN(n17164) );
  NAND2_X1 U20526 ( .A1(n17164), .A2(n17188), .ZN(n17187) );
  NAND2_X1 U20527 ( .A1(n17189), .A2(n17187), .ZN(n17181) );
  NOR2_X1 U20528 ( .A1(n17178), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n17165) );
  OAI21_X1 U20529 ( .B1(n17181), .B2(n17165), .A(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n17166) );
  NAND2_X1 U20530 ( .A1(n17167), .A2(n17166), .ZN(n17168) );
  AOI21_X1 U20531 ( .B1(n17169), .B2(n20277), .A(n17168), .ZN(n17170) );
  NAND2_X1 U20532 ( .A1(n17172), .A2(n20267), .ZN(n17173) );
  OAI211_X1 U20533 ( .C1(n17175), .C2(n17443), .A(n17174), .B(n17173), .ZN(
        P2_U3017) );
  INV_X1 U20534 ( .A(n17177), .ZN(n17180) );
  NOR3_X1 U20535 ( .A1(n17178), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        n17188), .ZN(n17179) );
  AOI211_X1 U20536 ( .C1(n17181), .C2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n17180), .B(n17179), .ZN(n17182) );
  OAI21_X1 U20537 ( .B1(n17183), .B2(n20259), .A(n17182), .ZN(n17184) );
  OAI211_X1 U20538 ( .C1(n17189), .C2(n17188), .A(n17187), .B(n17186), .ZN(
        n17190) );
  AOI21_X1 U20539 ( .B1(n17191), .B2(n20280), .A(n17190), .ZN(n17192) );
  OAI21_X1 U20540 ( .B1(n18091), .B2(n17193), .A(n17192), .ZN(n17194) );
  OAI21_X1 U20541 ( .B1(n17197), .B2(n17443), .A(n17196), .ZN(P2_U3019) );
  NOR2_X1 U20542 ( .A1(n17198), .A2(n18091), .ZN(n17207) );
  NAND2_X1 U20543 ( .A1(n17225), .A2(n20257), .ZN(n17215) );
  NAND3_X1 U20544 ( .A1(n17199), .A2(n17394), .A3(n17214), .ZN(n17213) );
  AOI21_X1 U20545 ( .B1(n17215), .B2(n17213), .A(n17202), .ZN(n17200) );
  AOI211_X1 U20546 ( .C1(n17203), .C2(n17202), .A(n17201), .B(n17200), .ZN(
        n17204) );
  OAI21_X1 U20547 ( .B1(n17205), .B2(n20259), .A(n17204), .ZN(n17206) );
  AOI211_X1 U20548 ( .C1(n17208), .C2(n20267), .A(n17207), .B(n17206), .ZN(
        n17209) );
  OAI21_X1 U20549 ( .B1(n17210), .B2(n17443), .A(n17209), .ZN(P2_U3020) );
  NOR2_X1 U20550 ( .A1(n17211), .A2(n18091), .ZN(n17217) );
  OAI211_X1 U20551 ( .C1(n17215), .C2(n17214), .A(n17213), .B(n17212), .ZN(
        n17216) );
  AOI211_X1 U20552 ( .C1(n17218), .C2(n20280), .A(n17217), .B(n17216), .ZN(
        n17221) );
  OAI211_X1 U20553 ( .C1(n17222), .C2(n17443), .A(n17221), .B(n17220), .ZN(
        P2_U3021) );
  NAND2_X1 U20554 ( .A1(n17394), .A2(n17223), .ZN(n17224) );
  NAND2_X1 U20555 ( .A1(n10602), .A2(n17224), .ZN(n17226) );
  NAND3_X1 U20556 ( .A1(n20257), .A2(n17226), .A3(n17225), .ZN(n17227) );
  OAI211_X1 U20557 ( .C1(n17229), .C2(n20259), .A(n17228), .B(n17227), .ZN(
        n17232) );
  NOR2_X1 U20558 ( .A1(n17230), .A2(n17443), .ZN(n17231) );
  AOI211_X1 U20559 ( .C1(n20277), .C2(n17233), .A(n17232), .B(n17231), .ZN(
        n17234) );
  OAI21_X1 U20560 ( .B1(n20290), .B2(n17235), .A(n17234), .ZN(P2_U3022) );
  NOR2_X1 U20561 ( .A1(n17236), .A2(n18091), .ZN(n17245) );
  NOR3_X1 U20562 ( .A1(n17238), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        n17237), .ZN(n17250) );
  OAI21_X1 U20563 ( .B1(n17252), .B2(n17250), .A(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17243) );
  NAND4_X1 U20564 ( .A1(n17240), .A2(n17394), .A3(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A4(n17239), .ZN(n17241) );
  NAND3_X1 U20565 ( .A1(n17243), .A2(n17242), .A3(n17241), .ZN(n17244) );
  AOI211_X1 U20566 ( .C1(n17246), .C2(n20280), .A(n17245), .B(n17244), .ZN(
        n17248) );
  OAI211_X1 U20567 ( .C1(n17249), .C2(n17443), .A(n17248), .B(n17247), .ZN(
        P2_U3023) );
  NOR2_X1 U20568 ( .A1(n17992), .A2(n18091), .ZN(n17255) );
  AOI211_X1 U20569 ( .C1(n17252), .C2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n17251), .B(n17250), .ZN(n17253) );
  OAI21_X1 U20570 ( .B1(n17993), .B2(n20259), .A(n17253), .ZN(n17254) );
  AOI211_X1 U20571 ( .C1(n17256), .C2(n20279), .A(n17255), .B(n17254), .ZN(
        n17257) );
  OAI21_X1 U20572 ( .B1(n20290), .B2(n17258), .A(n17257), .ZN(P2_U3024) );
  NOR2_X1 U20573 ( .A1(n17260), .A2(n17259), .ZN(n17265) );
  XNOR2_X1 U20574 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n17262) );
  OAI21_X1 U20575 ( .B1(n17263), .B2(n17262), .A(n17261), .ZN(n17264) );
  AOI211_X1 U20576 ( .C1(n17266), .C2(n20280), .A(n17265), .B(n17264), .ZN(
        n17267) );
  OAI21_X1 U20577 ( .B1(n18091), .B2(n17268), .A(n17267), .ZN(n17269) );
  AOI21_X1 U20578 ( .B1(n17270), .B2(n20267), .A(n17269), .ZN(n17271) );
  OAI21_X1 U20579 ( .B1(n17272), .B2(n17443), .A(n17271), .ZN(P2_U3026) );
  NOR2_X1 U20580 ( .A1(n17273), .A2(n18091), .ZN(n17281) );
  INV_X1 U20581 ( .A(n17313), .ZN(n17286) );
  NOR3_X1 U20582 ( .A1(n17286), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n17274), .ZN(n17275) );
  AOI211_X1 U20583 ( .C1(n17277), .C2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n17276), .B(n17275), .ZN(n17278) );
  OAI21_X1 U20584 ( .B1(n17279), .B2(n20259), .A(n17278), .ZN(n17280) );
  AOI211_X1 U20585 ( .C1(n17282), .C2(n20267), .A(n17281), .B(n17280), .ZN(
        n17283) );
  OAI21_X1 U20586 ( .B1(n17284), .B2(n17443), .A(n17283), .ZN(P2_U3028) );
  OAI22_X1 U20587 ( .A1(n17295), .A2(n20290), .B1(n17286), .B2(n17285), .ZN(
        n17293) );
  NOR2_X1 U20588 ( .A1(n17287), .A2(n18091), .ZN(n17291) );
  OAI21_X1 U20589 ( .B1(n17289), .B2(n20259), .A(n17288), .ZN(n17290) );
  AOI211_X1 U20590 ( .C1(n17293), .C2(n17292), .A(n17291), .B(n17290), .ZN(
        n17298) );
  INV_X1 U20591 ( .A(n17294), .ZN(n17296) );
  NOR2_X1 U20592 ( .A1(n17419), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n17297) );
  OAI21_X1 U20593 ( .B1(n17300), .B2(n20259), .A(n17299), .ZN(n17304) );
  AOI21_X1 U20594 ( .B1(n17301), .B2(n20267), .A(n17313), .ZN(n17302) );
  NOR3_X1 U20595 ( .A1(n17302), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        n17315), .ZN(n17303) );
  NAND2_X1 U20596 ( .A1(n17306), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n17307) );
  OAI211_X1 U20597 ( .C1(n17443), .C2(n17309), .A(n17308), .B(n17307), .ZN(
        P2_U3030) );
  NAND2_X1 U20598 ( .A1(n17310), .A2(n20279), .ZN(n17322) );
  INV_X1 U20599 ( .A(n17311), .ZN(n17312) );
  AOI21_X1 U20600 ( .B1(n17313), .B2(n17315), .A(n17312), .ZN(n17314) );
  OAI21_X1 U20601 ( .B1(n17316), .B2(n17315), .A(n17314), .ZN(n17319) );
  NOR2_X1 U20602 ( .A1(n17317), .A2(n20259), .ZN(n17318) );
  AOI211_X1 U20603 ( .C1(n17320), .C2(n20277), .A(n17319), .B(n17318), .ZN(
        n17321) );
  OAI211_X1 U20604 ( .C1(n17323), .C2(n20290), .A(n17322), .B(n17321), .ZN(
        P2_U3031) );
  INV_X1 U20605 ( .A(n20257), .ZN(n17437) );
  AOI21_X1 U20606 ( .B1(n17326), .B2(n17325), .A(n17437), .ZN(n17361) );
  AND2_X1 U20607 ( .A1(n17341), .A2(n17327), .ZN(n17355) );
  NOR2_X1 U20608 ( .A1(n17361), .A2(n17355), .ZN(n17349) );
  INV_X1 U20609 ( .A(n17349), .ZN(n17337) );
  NOR2_X1 U20610 ( .A1(n17328), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n17330) );
  INV_X1 U20611 ( .A(n17341), .ZN(n17329) );
  AOI211_X1 U20612 ( .C1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(n17330), .B(n17329), .ZN(
        n17331) );
  AOI211_X1 U20613 ( .C1(n17333), .C2(n20280), .A(n17332), .B(n17331), .ZN(
        n17334) );
  OAI21_X1 U20614 ( .B1(n18091), .B2(n17335), .A(n17334), .ZN(n17336) );
  AOI21_X1 U20615 ( .B1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n17337), .A(
        n17336), .ZN(n17338) );
  OAI211_X1 U20616 ( .C1(n17340), .C2(n17443), .A(n17339), .B(n17338), .ZN(
        P2_U3032) );
  NAND3_X1 U20617 ( .A1(n17341), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A3(
        n17348), .ZN(n17342) );
  OAI211_X1 U20618 ( .C1(n17344), .C2(n20259), .A(n17343), .B(n17342), .ZN(
        n17345) );
  AOI21_X1 U20619 ( .B1(n20277), .B2(n17346), .A(n17345), .ZN(n17347) );
  OAI21_X1 U20620 ( .B1(n17349), .B2(n17348), .A(n17347), .ZN(n17350) );
  AOI21_X1 U20621 ( .B1(n17351), .B2(n20279), .A(n17350), .ZN(n17352) );
  OAI21_X1 U20622 ( .B1(n17353), .B2(n20290), .A(n17352), .ZN(P2_U3033) );
  NOR2_X1 U20623 ( .A1(n17354), .A2(n18091), .ZN(n17360) );
  INV_X1 U20624 ( .A(n17355), .ZN(n17356) );
  OAI211_X1 U20625 ( .C1(n17358), .C2(n20259), .A(n17357), .B(n17356), .ZN(
        n17359) );
  AOI211_X1 U20626 ( .C1(n17361), .C2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n17360), .B(n17359), .ZN(n17364) );
  NAND2_X1 U20627 ( .A1(n17362), .A2(n20279), .ZN(n17363) );
  OAI211_X1 U20628 ( .C1(n17365), .C2(n20290), .A(n17364), .B(n17363), .ZN(
        P2_U3034) );
  INV_X1 U20629 ( .A(n17366), .ZN(n17375) );
  AND2_X1 U20630 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17367) );
  NAND3_X1 U20631 ( .A1(n17367), .A2(n17394), .A3(n17372), .ZN(n17368) );
  OAI211_X1 U20632 ( .C1(n17370), .C2(n20259), .A(n17369), .B(n17368), .ZN(
        n17374) );
  INV_X1 U20633 ( .A(n17371), .ZN(n17400) );
  AOI21_X1 U20634 ( .B1(n10240), .B2(n20257), .A(n17400), .ZN(n17386) );
  NAND3_X1 U20635 ( .A1(n17385), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(
        n17394), .ZN(n17383) );
  AOI21_X1 U20636 ( .B1(n17386), .B2(n17383), .A(n17372), .ZN(n17373) );
  AOI211_X1 U20637 ( .C1(n20277), .C2(n17375), .A(n17374), .B(n17373), .ZN(
        n17378) );
  NAND2_X1 U20638 ( .A1(n17376), .A2(n20279), .ZN(n17377) );
  OAI211_X1 U20639 ( .C1(n17379), .C2(n20290), .A(n17378), .B(n17377), .ZN(
        P2_U3035) );
  NAND2_X1 U20640 ( .A1(n17381), .A2(n20280), .ZN(n17384) );
  NAND3_X1 U20641 ( .A1(n17384), .A2(n17383), .A3(n17382), .ZN(n17388) );
  NOR2_X1 U20642 ( .A1(n17386), .A2(n17385), .ZN(n17387) );
  AOI211_X1 U20643 ( .C1(n20277), .C2(n17389), .A(n17388), .B(n17387), .ZN(
        n17390) );
  OAI211_X1 U20644 ( .C1(n17392), .C2(n17443), .A(n17391), .B(n17390), .ZN(
        P2_U3036) );
  NOR2_X1 U20645 ( .A1(n17393), .A2(n18091), .ZN(n17399) );
  NAND2_X1 U20646 ( .A1(n10240), .A2(n17394), .ZN(n17395) );
  OAI211_X1 U20647 ( .C1(n17397), .C2(n20259), .A(n17396), .B(n17395), .ZN(
        n17398) );
  AOI211_X1 U20648 ( .C1(n17400), .C2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n17399), .B(n17398), .ZN(n17403) );
  NAND2_X1 U20649 ( .A1(n17401), .A2(n20279), .ZN(n17402) );
  OAI211_X1 U20650 ( .C1(n17404), .C2(n20290), .A(n17403), .B(n17402), .ZN(
        P2_U3037) );
  NAND3_X1 U20651 ( .A1(n18076), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A3(
        n20257), .ZN(n17411) );
  OAI21_X1 U20652 ( .B1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n17405), .ZN(n17407) );
  OAI21_X1 U20653 ( .B1(n18075), .B2(n17407), .A(n17406), .ZN(n17408) );
  AOI21_X1 U20654 ( .B1(n17409), .B2(n20280), .A(n17408), .ZN(n17410) );
  OAI211_X1 U20655 ( .C1(n18091), .C2(n17412), .A(n17411), .B(n17410), .ZN(
        n17413) );
  AOI21_X1 U20656 ( .B1(n17414), .B2(n20279), .A(n17413), .ZN(n17415) );
  OAI21_X1 U20657 ( .B1(n17416), .B2(n20290), .A(n17415), .ZN(P2_U3038) );
  OAI21_X1 U20658 ( .B1(n17419), .B2(n17418), .A(n17417), .ZN(n17420) );
  OAI21_X1 U20659 ( .B1(n17421), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n17420), .ZN(n17425) );
  AOI21_X1 U20660 ( .B1(n17423), .B2(n20280), .A(n17422), .ZN(n17424) );
  OAI211_X1 U20661 ( .C1(n18091), .C2(n17426), .A(n17425), .B(n17424), .ZN(
        n17427) );
  AOI21_X1 U20662 ( .B1(n17428), .B2(n20279), .A(n17427), .ZN(n17429) );
  OAI21_X1 U20663 ( .B1(n17430), .B2(n20290), .A(n17429), .ZN(P2_U3040) );
  NAND2_X1 U20664 ( .A1(n17431), .A2(n20267), .ZN(n17442) );
  NOR2_X1 U20665 ( .A1(n18096), .A2(n18095), .ZN(n20265) );
  OAI221_X1 U20666 ( .B1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .C1(n17436), .C2(n20264), .A(
        n20265), .ZN(n17433) );
  OAI211_X1 U20667 ( .C1(n17434), .C2(n20259), .A(n17433), .B(n17432), .ZN(
        n17439) );
  NOR2_X1 U20668 ( .A1(n18096), .A2(n17435), .ZN(n20261) );
  NOR3_X1 U20669 ( .A1(n20261), .A2(n17437), .A3(n17436), .ZN(n17438) );
  AOI211_X1 U20670 ( .C1(n20277), .C2(n17440), .A(n17439), .B(n17438), .ZN(
        n17441) );
  OAI211_X1 U20671 ( .C1(n17444), .C2(n17443), .A(n17442), .B(n17441), .ZN(
        P2_U3041) );
  MUX2_X1 U20672 ( .A(n17445), .B(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .S(
        n12943), .Z(n17446) );
  NAND2_X1 U20673 ( .A1(n17446), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n17487) );
  INV_X1 U20674 ( .A(n17447), .ZN(n17509) );
  INV_X1 U20675 ( .A(n11209), .ZN(n17448) );
  NAND2_X1 U20676 ( .A1(n17449), .A2(n17448), .ZN(n17473) );
  MUX2_X1 U20677 ( .A(n17473), .B(n17498), .S(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n17450) );
  AOI21_X1 U20678 ( .B1(n10091), .B2(n17509), .A(n17450), .ZN(n17646) );
  OAI21_X1 U20679 ( .B1(n17646), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n11386), 
        .ZN(n17452) );
  AOI22_X1 U20680 ( .A1(n17487), .A2(n17452), .B1(n17451), .B2(n17685), .ZN(
        n17464) );
  INV_X1 U20681 ( .A(n17453), .ZN(n17456) );
  NOR2_X1 U20682 ( .A1(n17986), .A2(n17454), .ZN(n17455) );
  NAND2_X1 U20683 ( .A1(n17456), .A2(n17455), .ZN(n17460) );
  NAND4_X1 U20684 ( .A1(n17460), .A2(n17459), .A3(n17458), .A4(n17457), .ZN(
        n17657) );
  NAND2_X1 U20685 ( .A1(n17657), .A2(n20180), .ZN(n17462) );
  AOI22_X1 U20686 ( .A1(n17688), .A2(P2_FLUSH_REG_SCAN_IN), .B1(n17703), .B2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n17461) );
  NAND2_X1 U20687 ( .A1(n17462), .A2(n17461), .ZN(n17990) );
  NAND2_X1 U20688 ( .A1(n17511), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n17463) );
  OAI21_X1 U20689 ( .B1(n17464), .B2(n17511), .A(n17463), .ZN(P2_U3601) );
  NAND2_X1 U20690 ( .A1(n12943), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17465) );
  NAND2_X1 U20691 ( .A1(n17466), .A2(n17465), .ZN(n17489) );
  NAND2_X1 U20692 ( .A1(n17467), .A2(n17509), .ZN(n17475) );
  INV_X1 U20693 ( .A(n17468), .ZN(n17471) );
  INV_X1 U20694 ( .A(n17469), .ZN(n17470) );
  NAND2_X1 U20695 ( .A1(n17471), .A2(n17470), .ZN(n17472) );
  AOI22_X1 U20696 ( .A1(n17498), .A2(n10580), .B1(n17473), .B2(n17472), .ZN(
        n17474) );
  NAND2_X1 U20697 ( .A1(n17475), .A2(n17474), .ZN(n17643) );
  AOI22_X1 U20698 ( .A1(n20903), .A2(n17685), .B1(n17491), .B2(n17643), .ZN(
        n17476) );
  OAI21_X1 U20699 ( .B1(n17487), .B2(n17489), .A(n17476), .ZN(n17477) );
  MUX2_X1 U20700 ( .A(n17477), .B(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .S(
        n17511), .Z(P2_U3600) );
  AND2_X1 U20701 ( .A1(n11465), .A2(n17478), .ZN(n17501) );
  NAND2_X1 U20702 ( .A1(n17479), .A2(n11000), .ZN(n17495) );
  NAND2_X1 U20703 ( .A1(n17480), .A2(n17495), .ZN(n17486) );
  NAND2_X1 U20704 ( .A1(n20281), .A2(n17509), .ZN(n17485) );
  OR2_X1 U20705 ( .A1(n17653), .A2(n17652), .ZN(n17494) );
  NOR2_X1 U20706 ( .A1(n17481), .A2(n17482), .ZN(n17483) );
  AOI22_X1 U20707 ( .A1(n17494), .A2(n17486), .B1(n17483), .B2(n17498), .ZN(
        n17484) );
  OAI211_X1 U20708 ( .C1(n17501), .C2(n17486), .A(n17485), .B(n17484), .ZN(
        n17641) );
  INV_X1 U20709 ( .A(n20896), .ZN(n17490) );
  INV_X1 U20710 ( .A(n17487), .ZN(n17488) );
  AOI222_X1 U20711 ( .A1(n17641), .A2(n17491), .B1(n17685), .B2(n17490), .C1(
        n17489), .C2(n17488), .ZN(n17493) );
  NAND2_X1 U20712 ( .A1(n17511), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n17492) );
  OAI21_X1 U20713 ( .B1(n17493), .B2(n17511), .A(n17492), .ZN(P2_U3599) );
  INV_X1 U20714 ( .A(n17685), .ZN(n17510) );
  AOI22_X1 U20715 ( .A1(n17494), .A2(n17495), .B1(n17482), .B2(n17498), .ZN(
        n17504) );
  INV_X1 U20716 ( .A(n17495), .ZN(n17496) );
  AOI21_X1 U20717 ( .B1(n17498), .B2(n17497), .A(n17496), .ZN(n17499) );
  OAI21_X1 U20718 ( .B1(n17501), .B2(n17500), .A(n17499), .ZN(n17502) );
  INV_X1 U20719 ( .A(n17502), .ZN(n17503) );
  MUX2_X1 U20720 ( .A(n17504), .B(n17503), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n17507) );
  INV_X1 U20721 ( .A(n17505), .ZN(n17506) );
  NAND2_X1 U20722 ( .A1(n17507), .A2(n17506), .ZN(n17508) );
  AOI21_X1 U20723 ( .B1(n10798), .B2(n17509), .A(n17508), .ZN(n17649) );
  OAI22_X1 U20724 ( .A1(n20535), .A2(n17510), .B1(n17649), .B2(n17983), .ZN(
        n17512) );
  MUX2_X1 U20725 ( .A(n17512), .B(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n17511), .Z(P2_U3596) );
  INV_X1 U20726 ( .A(n20497), .ZN(n20536) );
  AOI21_X1 U20727 ( .B1(n20348), .B2(n20310), .A(n20691), .ZN(n17514) );
  INV_X1 U20728 ( .A(n20888), .ZN(n20692) );
  NAND2_X1 U20729 ( .A1(n21853), .A2(n20900), .ZN(n20351) );
  NOR2_X1 U20730 ( .A1(n20498), .A2(n20351), .ZN(n20315) );
  NOR2_X1 U20731 ( .A1(n21853), .A2(n20900), .ZN(n20694) );
  INV_X1 U20732 ( .A(n20694), .ZN(n20741) );
  NOR2_X1 U20733 ( .A1(n17642), .A2(n20741), .ZN(n20796) );
  NOR2_X1 U20734 ( .A1(n20315), .A2(n20796), .ZN(n17522) );
  OAI21_X1 U20735 ( .B1(n9836), .B2(n20315), .A(n20748), .ZN(n17518) );
  INV_X1 U20736 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17530) );
  INV_X1 U20737 ( .A(n17519), .ZN(n17523) );
  OAI21_X1 U20738 ( .B1(n17520), .B2(n20315), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n17521) );
  AOI22_X2 U20739 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n17590), .B1(
        BUF1_REG_24__SCAN_IN), .B2(n17589), .ZN(n20759) );
  INV_X1 U20740 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n18125) );
  OAI22_X2 U20741 ( .A1(n18125), .A2(n17592), .B1(n16849), .B2(n17591), .ZN(
        n20756) );
  AND2_X1 U20742 ( .A1(n17588), .A2(n17526), .ZN(n20745) );
  AOI22_X1 U20743 ( .A1(n20756), .A2(n20316), .B1(n20745), .B2(n20315), .ZN(
        n17527) );
  OAI21_X1 U20744 ( .B1(n20759), .B2(n20310), .A(n17527), .ZN(n17528) );
  AOI21_X1 U20745 ( .B1(n20317), .B2(n20746), .A(n17528), .ZN(n17529) );
  OAI21_X1 U20746 ( .B1(n20321), .B2(n17530), .A(n17529), .ZN(P2_U3048) );
  AOI22_X1 U20747 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n17589), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n17590), .ZN(n20789) );
  AOI22_X1 U20748 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n17589), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n17590), .ZN(n20720) );
  AOI22_X1 U20749 ( .A1(n20316), .A2(n20786), .B1(n20315), .B2(n20784), .ZN(
        n17532) );
  OAI21_X1 U20750 ( .B1(n20789), .B2(n20310), .A(n17532), .ZN(n17533) );
  AOI21_X1 U20751 ( .B1(n20317), .B2(n20785), .A(n17533), .ZN(n17534) );
  OAI21_X1 U20752 ( .B1(n20321), .B2(n17535), .A(n17534), .ZN(P2_U3053) );
  AOI22_X1 U20753 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n17590), .B1(
        BUF1_REG_30__SCAN_IN), .B2(n17589), .ZN(n20795) );
  NOR2_X1 U20754 ( .A1(n20310), .A2(n20795), .ZN(n17539) );
  AOI22_X1 U20755 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n17589), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n17590), .ZN(n20726) );
  INV_X1 U20756 ( .A(n20315), .ZN(n20309) );
  NAND2_X1 U20757 ( .A1(n17588), .A2(n17537), .ZN(n20724) );
  OAI22_X1 U20758 ( .A1(n20348), .A2(n20726), .B1(n20309), .B2(n20724), .ZN(
        n17538) );
  AOI211_X1 U20759 ( .C1(n20317), .C2(n20791), .A(n17539), .B(n17538), .ZN(
        n17540) );
  OAI21_X1 U20760 ( .B1(n20321), .B2(n17541), .A(n17540), .ZN(P2_U3054) );
  NOR2_X2 U20761 ( .A1(n20497), .A2(n20476), .ZN(n20344) );
  NOR2_X1 U20762 ( .A1(n20377), .A2(n20344), .ZN(n17548) );
  INV_X1 U20763 ( .A(n20748), .ZN(n20661) );
  NOR3_X1 U20764 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20909), .A3(
        n20351), .ZN(n17549) );
  INV_X1 U20765 ( .A(n17549), .ZN(n17594) );
  OAI21_X1 U20766 ( .B1(n17544), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n17594), 
        .ZN(n17545) );
  NOR2_X1 U20767 ( .A1(n17618), .A2(n20351), .ZN(n17551) );
  AOI21_X1 U20768 ( .B1(n17545), .B2(n20692), .A(n17551), .ZN(n17546) );
  INV_X1 U20769 ( .A(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17557) );
  OAI21_X1 U20770 ( .B1(n17550), .B2(n17549), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n17553) );
  INV_X1 U20771 ( .A(n17551), .ZN(n17552) );
  NAND2_X1 U20772 ( .A1(n17553), .A2(n17552), .ZN(n17596) );
  INV_X1 U20773 ( .A(n20745), .ZN(n20538) );
  INV_X1 U20774 ( .A(n20759), .ZN(n17629) );
  AOI22_X1 U20775 ( .A1(n20377), .A2(n20756), .B1(n20344), .B2(n17629), .ZN(
        n17554) );
  OAI21_X1 U20776 ( .B1(n20538), .B2(n17594), .A(n17554), .ZN(n17555) );
  AOI21_X1 U20777 ( .B1(n17596), .B2(n20746), .A(n17555), .ZN(n17556) );
  OAI21_X1 U20778 ( .B1(n17599), .B2(n17557), .A(n17556), .ZN(P2_U3064) );
  INV_X1 U20779 ( .A(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n17562) );
  INV_X1 U20780 ( .A(n20760), .ZN(n20510) );
  AOI22_X1 U20781 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n17589), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n17590), .ZN(n20708) );
  INV_X1 U20782 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n18110) );
  AOI22_X1 U20783 ( .A1(n20377), .A2(n20762), .B1(n20344), .B2(n20705), .ZN(
        n17559) );
  OAI21_X1 U20784 ( .B1(n20510), .B2(n17594), .A(n17559), .ZN(n17560) );
  AOI21_X1 U20785 ( .B1(n17596), .B2(n20761), .A(n17560), .ZN(n17561) );
  OAI21_X1 U20786 ( .B1(n17599), .B2(n17562), .A(n17561), .ZN(P2_U3065) );
  INV_X1 U20787 ( .A(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17568) );
  NAND2_X1 U20788 ( .A1(n17588), .A2(n17564), .ZN(n20709) );
  AOI22_X1 U20789 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n17589), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n17590), .ZN(n20713) );
  AOI22_X2 U20790 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n17590), .B1(
        BUF1_REG_26__SCAN_IN), .B2(n17589), .ZN(n20771) );
  INV_X1 U20791 ( .A(n20771), .ZN(n20634) );
  AOI22_X1 U20792 ( .A1(n20377), .A2(n20768), .B1(n20344), .B2(n20634), .ZN(
        n17565) );
  OAI21_X1 U20793 ( .B1(n20709), .B2(n17594), .A(n17565), .ZN(n17566) );
  AOI21_X1 U20794 ( .B1(n17596), .B2(n20767), .A(n17566), .ZN(n17567) );
  OAI21_X1 U20795 ( .B1(n17599), .B2(n17568), .A(n17567), .ZN(P2_U3066) );
  INV_X1 U20796 ( .A(n20772), .ZN(n20555) );
  OAI22_X2 U20797 ( .A1(n17570), .A2(n17592), .B1(n17727), .B2(n17591), .ZN(
        n20774) );
  AOI22_X2 U20798 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n17589), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n17590), .ZN(n20777) );
  INV_X1 U20799 ( .A(n20777), .ZN(n20638) );
  AOI22_X1 U20800 ( .A1(n20377), .A2(n20774), .B1(n20344), .B2(n20638), .ZN(
        n17571) );
  OAI21_X1 U20801 ( .B1(n20555), .B2(n17594), .A(n17571), .ZN(n17572) );
  AOI21_X1 U20802 ( .B1(n17596), .B2(n20773), .A(n17572), .ZN(n17573) );
  OAI21_X1 U20803 ( .B1(n17599), .B2(n10871), .A(n17573), .ZN(P2_U3067) );
  INV_X1 U20804 ( .A(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17579) );
  AND2_X1 U20805 ( .A1(n17588), .A2(n17575), .ZN(n20778) );
  INV_X1 U20806 ( .A(n20778), .ZN(n20308) );
  INV_X1 U20807 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n21772) );
  OAI22_X2 U20808 ( .A1(n21772), .A2(n17592), .B1(n16823), .B2(n17591), .ZN(
        n20780) );
  AOI22_X2 U20809 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n17590), .B1(
        BUF1_REG_28__SCAN_IN), .B2(n17589), .ZN(n20783) );
  INV_X1 U20810 ( .A(n20783), .ZN(n20641) );
  AOI22_X1 U20811 ( .A1(n20377), .A2(n20780), .B1(n20344), .B2(n20641), .ZN(
        n17576) );
  OAI21_X1 U20812 ( .B1(n20308), .B2(n17594), .A(n17576), .ZN(n17577) );
  AOI21_X1 U20813 ( .B1(n17596), .B2(n20779), .A(n17577), .ZN(n17578) );
  OAI21_X1 U20814 ( .B1(n17599), .B2(n17579), .A(n17578), .ZN(P2_U3068) );
  INV_X1 U20815 ( .A(n20784), .ZN(n20719) );
  INV_X1 U20816 ( .A(n20789), .ZN(n20678) );
  AOI22_X1 U20817 ( .A1(n20377), .A2(n20786), .B1(n20344), .B2(n20678), .ZN(
        n17580) );
  OAI21_X1 U20818 ( .B1(n20719), .B2(n17594), .A(n17580), .ZN(n17581) );
  AOI21_X1 U20819 ( .B1(n17596), .B2(n20785), .A(n17581), .ZN(n17582) );
  OAI21_X1 U20820 ( .B1(n17599), .B2(n17583), .A(n17582), .ZN(P2_U3069) );
  INV_X1 U20821 ( .A(n20795), .ZN(n20647) );
  AOI22_X1 U20822 ( .A1(n20377), .A2(n20792), .B1(n20344), .B2(n20647), .ZN(
        n17584) );
  OAI21_X1 U20823 ( .B1(n20724), .B2(n17594), .A(n17584), .ZN(n17585) );
  AOI21_X1 U20824 ( .B1(n17596), .B2(n20791), .A(n17585), .ZN(n17586) );
  OAI21_X1 U20825 ( .B1(n17599), .B2(n10969), .A(n17586), .ZN(P2_U3070) );
  INV_X1 U20826 ( .A(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n17598) );
  AND2_X1 U20827 ( .A1(n17588), .A2(n10734), .ZN(n20797) );
  INV_X1 U20828 ( .A(n20797), .ZN(n20574) );
  AOI22_X1 U20829 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n17590), .B1(
        BUF1_REG_23__SCAN_IN), .B2(n17589), .ZN(n20738) );
  INV_X1 U20830 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n18178) );
  AOI22_X1 U20831 ( .A1(n20377), .A2(n20800), .B1(n20344), .B2(n20733), .ZN(
        n17593) );
  OAI21_X1 U20832 ( .B1(n20574), .B2(n17594), .A(n17593), .ZN(n17595) );
  AOI21_X1 U20833 ( .B1(n17596), .B2(n20798), .A(n17595), .ZN(n17597) );
  OAI21_X1 U20834 ( .B1(n17599), .B2(n17598), .A(n17597), .ZN(P2_U3071) );
  NAND2_X1 U20835 ( .A1(n20535), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20470) );
  OAI21_X1 U20836 ( .B1(n20470), .B2(n20666), .A(n20888), .ZN(n17607) );
  NAND2_X1 U20837 ( .A1(n20437), .A2(n20909), .ZN(n17606) );
  INV_X1 U20838 ( .A(n17606), .ZN(n17600) );
  OR2_X1 U20839 ( .A1(n17607), .A2(n17600), .ZN(n17604) );
  NAND2_X1 U20840 ( .A1(n10929), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n17601) );
  NAND2_X1 U20841 ( .A1(n17601), .A2(n20750), .ZN(n17602) );
  NOR2_X1 U20842 ( .A1(n20919), .A2(n17606), .ZN(n20429) );
  AOI21_X1 U20843 ( .B1(n17602), .B2(n10616), .A(n20661), .ZN(n17603) );
  INV_X1 U20844 ( .A(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17612) );
  INV_X1 U20845 ( .A(n20430), .ZN(n17609) );
  AOI22_X1 U20846 ( .A1(n20756), .A2(n20440), .B1(n20745), .B2(n20429), .ZN(
        n17608) );
  OAI21_X1 U20847 ( .B1(n20759), .B2(n17609), .A(n17608), .ZN(n17610) );
  AOI21_X1 U20848 ( .B1(n20746), .B2(n20431), .A(n17610), .ZN(n17611) );
  OAI21_X1 U20849 ( .B1(n20435), .B2(n17612), .A(n17611), .ZN(P2_U3088) );
  NAND2_X1 U20850 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n20900), .ZN(
        n20602) );
  NOR2_X1 U20851 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20602), .ZN(
        n20543) );
  NAND2_X1 U20852 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20543), .ZN(
        n20575) );
  OAI221_X1 U20853 ( .B1(n20691), .B2(n20633), .C1(n20691), .C2(n20601), .A(
        n20575), .ZN(n17613) );
  NAND2_X1 U20854 ( .A1(n20750), .A2(n17613), .ZN(n17614) );
  NOR2_X1 U20855 ( .A1(n20909), .A2(n20602), .ZN(n20613) );
  INV_X1 U20856 ( .A(n20613), .ZN(n20607) );
  NOR2_X1 U20857 ( .A1(n20607), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n20595) );
  INV_X1 U20858 ( .A(n20598), .ZN(n17624) );
  INV_X1 U20859 ( .A(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17623) );
  OAI21_X1 U20860 ( .B1(n17616), .B2(n20595), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n17617) );
  INV_X1 U20861 ( .A(n20595), .ZN(n17620) );
  AOI22_X1 U20862 ( .A1(n20597), .A2(n20756), .B1(n20562), .B2(n17629), .ZN(
        n17619) );
  OAI21_X1 U20863 ( .B1(n20538), .B2(n17620), .A(n17619), .ZN(n17621) );
  AOI21_X1 U20864 ( .B1(n20596), .B2(n20746), .A(n17621), .ZN(n17622) );
  OAI21_X1 U20865 ( .B1(n17624), .B2(n17623), .A(n17622), .ZN(P2_U3128) );
  OAI21_X1 U20866 ( .B1(n20686), .B2(n20652), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n17628) );
  INV_X1 U20867 ( .A(n20382), .ZN(n17625) );
  NOR2_X1 U20868 ( .A1(n17625), .A2(n21853), .ZN(n17630) );
  INV_X1 U20869 ( .A(n20695), .ZN(n20383) );
  NAND2_X1 U20870 ( .A1(n17630), .A2(n20383), .ZN(n17627) );
  NOR2_X1 U20871 ( .A1(n20498), .A2(n20741), .ZN(n20650) );
  OAI211_X1 U20872 ( .C1(n20650), .C2(n20750), .A(n17631), .B(n20748), .ZN(
        n17626) );
  INV_X1 U20873 ( .A(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17636) );
  AOI22_X1 U20874 ( .A1(n20686), .A2(n20756), .B1(n20652), .B2(n17629), .ZN(
        n17635) );
  NAND3_X1 U20875 ( .A1(n17630), .A2(n20750), .A3(n20383), .ZN(n17633) );
  INV_X1 U20876 ( .A(n17631), .ZN(n17632) );
  AOI22_X1 U20877 ( .A1(n20651), .A2(n20746), .B1(n20745), .B2(n20650), .ZN(
        n17634) );
  OAI211_X1 U20878 ( .C1(n20656), .C2(n17636), .A(n17635), .B(n17634), .ZN(
        P2_U3144) );
  AOI22_X1 U20879 ( .A1(n20686), .A2(n20762), .B1(n20652), .B2(n20705), .ZN(
        n17638) );
  AOI22_X1 U20880 ( .A1(n20651), .A2(n20761), .B1(n20650), .B2(n20760), .ZN(
        n17637) );
  OAI211_X1 U20881 ( .C1(n20656), .C2(n17639), .A(n17638), .B(n17637), .ZN(
        P2_U3145) );
  INV_X1 U20882 ( .A(n17640), .ZN(n17683) );
  MUX2_X1 U20883 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n17641), .S(
        n17657), .Z(n17662) );
  OAI21_X1 U20884 ( .B1(n17643), .B2(n20919), .A(n17642), .ZN(n17645) );
  OAI21_X1 U20885 ( .B1(n17643), .B2(n20909), .A(n17657), .ZN(n17644) );
  AOI21_X1 U20886 ( .B1(n17646), .B2(n17645), .A(n17644), .ZN(n17647) );
  OAI21_X1 U20887 ( .B1(n17662), .B2(n20900), .A(n17647), .ZN(n17663) );
  INV_X1 U20888 ( .A(n17663), .ZN(n17648) );
  INV_X1 U20889 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18015) );
  AOI21_X1 U20890 ( .B1(n17648), .B2(n18015), .A(n17662), .ZN(n17679) );
  MUX2_X1 U20891 ( .A(n17650), .B(n17649), .S(n17657), .Z(n17678) );
  MUX2_X1 U20892 ( .A(n17653), .B(n17652), .S(n17651), .Z(n17656) );
  NOR2_X1 U20893 ( .A1(n17656), .A2(n17655), .ZN(n20925) );
  INV_X1 U20894 ( .A(n17657), .ZN(n17676) );
  NOR2_X1 U20895 ( .A1(n17659), .A2(n17658), .ZN(n17660) );
  NAND2_X1 U20896 ( .A1(n17661), .A2(n17660), .ZN(n20181) );
  NOR2_X1 U20897 ( .A1(P2_FLUSH_REG_SCAN_IN), .A2(P2_MORE_REG_SCAN_IN), .ZN(
        n17674) );
  NAND2_X1 U20898 ( .A1(n20900), .A2(n17662), .ZN(n17664) );
  NAND3_X1 U20899 ( .A1(n17678), .A2(n17664), .A3(n17663), .ZN(n17665) );
  NAND3_X1 U20900 ( .A1(n21853), .A2(n18015), .A3(n17665), .ZN(n17666) );
  OAI21_X1 U20901 ( .B1(n17668), .B2(n17667), .A(n17666), .ZN(n17669) );
  INV_X1 U20902 ( .A(n17669), .ZN(n17673) );
  INV_X1 U20903 ( .A(n17986), .ZN(n17671) );
  INV_X1 U20904 ( .A(n17985), .ZN(n17670) );
  NAND3_X1 U20905 ( .A1(n17671), .A2(n9710), .A3(n17670), .ZN(n17672) );
  OAI211_X1 U20906 ( .C1(n20181), .C2(n17674), .A(n17673), .B(n17672), .ZN(
        n17675) );
  AOI21_X1 U20907 ( .B1(n17676), .B2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n17675), .ZN(n17677) );
  OAI211_X1 U20908 ( .C1(n17679), .C2(n17678), .A(n20925), .B(n17677), .ZN(
        n17692) );
  OAI21_X1 U20909 ( .B1(n17692), .B2(P2_STATE2_REG_1__SCAN_IN), .A(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n17681) );
  OAI211_X1 U20910 ( .C1(n17683), .C2(n17682), .A(n17681), .B(n17680), .ZN(
        n17700) );
  OAI21_X1 U20911 ( .B1(n17685), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n17684), 
        .ZN(n17686) );
  OAI21_X1 U20912 ( .B1(n17700), .B2(n17687), .A(n17686), .ZN(n17694) );
  INV_X1 U20913 ( .A(n18013), .ZN(n20922) );
  INV_X1 U20914 ( .A(n17688), .ZN(n18011) );
  OAI211_X1 U20915 ( .C1(n20922), .C2(n18011), .A(n17690), .B(n17689), .ZN(
        n17691) );
  AOI21_X1 U20916 ( .B1(n17692), .B2(n20180), .A(n17691), .ZN(n17693) );
  OAI211_X1 U20917 ( .C1(n17700), .C2(n17703), .A(n17694), .B(n17693), .ZN(
        P2_U3176) );
  INV_X1 U20918 ( .A(n17700), .ZN(n17704) );
  OAI211_X1 U20919 ( .C1(n17704), .C2(n17695), .A(P2_STATE2_REG_1__SCAN_IN), 
        .B(n20819), .ZN(n17702) );
  INV_X1 U20920 ( .A(n20658), .ZN(n17699) );
  OAI21_X1 U20921 ( .B1(n17697), .B2(n20819), .A(n17696), .ZN(n17698) );
  NAND3_X1 U20922 ( .A1(n17700), .A2(n17699), .A3(n17698), .ZN(n17701) );
  NAND3_X1 U20923 ( .A1(n17702), .A2(n17996), .A3(n17701), .ZN(P2_U3177) );
  OAI21_X1 U20924 ( .B1(n17704), .B2(n17703), .A(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n17705) );
  NAND2_X1 U20925 ( .A1(n17705), .A2(n18011), .ZN(P2_U3593) );
  NAND4_X1 U20926 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(P3_EAX_REG_19__SCAN_IN), 
        .A3(P3_EAX_REG_18__SCAN_IN), .A4(P3_EAX_REG_17__SCAN_IN), .ZN(n18786)
         );
  INV_X1 U20927 ( .A(n18854), .ZN(n18847) );
  NOR2_X1 U20928 ( .A1(n18786), .A2(n18847), .ZN(n18841) );
  AOI21_X1 U20929 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n18886), .A(n18841), .ZN(
        n17725) );
  NAND2_X1 U20930 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n18841), .ZN(n18837) );
  INV_X1 U20931 ( .A(n18837), .ZN(n17724) );
  OAI22_X1 U20932 ( .A1(n17708), .A2(n18724), .B1(n18722), .B2(n17707), .ZN(
        n17712) );
  OAI22_X1 U20933 ( .A1(n18728), .A2(n17710), .B1(n18726), .B2(n17709), .ZN(
        n17711) );
  AOI211_X1 U20934 ( .C1(n18731), .C2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A(
        n17712), .B(n17711), .ZN(n17714) );
  AOI22_X1 U20935 ( .A1(n9704), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n18732), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n17713) );
  OAI211_X1 U20936 ( .C1(n9681), .C2(n21818), .A(n17714), .B(n17713), .ZN(
        n17720) );
  AOI22_X1 U20937 ( .A1(n18736), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n13878), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n17718) );
  AOI22_X1 U20938 ( .A1(n13279), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n18596), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n17717) );
  AOI22_X1 U20939 ( .A1(n18738), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n18737), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n17716) );
  AOI22_X1 U20940 ( .A1(n18740), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n18739), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n17715) );
  NAND4_X1 U20941 ( .A1(n17718), .A2(n17717), .A3(n17716), .A4(n17715), .ZN(
        n17719) );
  NOR2_X1 U20942 ( .A1(n17720), .A2(n17719), .ZN(n18673) );
  OAI22_X1 U20943 ( .A1(n18832), .A2(n18673), .B1(n18788), .B2(n17721), .ZN(
        n17722) );
  AOI21_X1 U20944 ( .B1(BUF2_REG_5__SCAN_IN), .B2(n18827), .A(n17722), .ZN(
        n17723) );
  OAI21_X1 U20945 ( .B1(n17725), .B2(n17724), .A(n17723), .ZN(P3_U2714) );
  NAND3_X1 U20946 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(P3_EAX_REG_17__SCAN_IN), 
        .A3(n18854), .ZN(n18848) );
  INV_X1 U20947 ( .A(n18848), .ZN(n17726) );
  AOI21_X1 U20948 ( .B1(P3_EAX_REG_19__SCAN_IN), .B2(n18886), .A(n17726), .ZN(
        n17732) );
  NAND2_X1 U20949 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n17726), .ZN(n18842) );
  INV_X1 U20950 ( .A(n18842), .ZN(n17731) );
  OAI22_X1 U20951 ( .A1(n18832), .A2(n17728), .B1(n18788), .B2(n17727), .ZN(
        n17729) );
  AOI21_X1 U20952 ( .B1(BUF2_REG_3__SCAN_IN), .B2(n18827), .A(n17729), .ZN(
        n17730) );
  OAI21_X1 U20953 ( .B1(n17732), .B2(n17731), .A(n17730), .ZN(P3_U2716) );
  NAND2_X1 U20954 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17733), .ZN(n18872) );
  NOR2_X1 U20955 ( .A1(n18986), .A2(n18872), .ZN(n17737) );
  AOI21_X1 U20956 ( .B1(n18886), .B2(P3_EAX_REG_13__SCAN_IN), .A(n17740), .ZN(
        n17735) );
  NAND2_X1 U20957 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n17740), .ZN(n18868) );
  INV_X1 U20958 ( .A(n18868), .ZN(n17734) );
  OAI222_X1 U20959 ( .A1(n18883), .A2(n13675), .B1(n18832), .B2(n17736), .C1(
        n17735), .C2(n17734), .ZN(P3_U2722) );
  AOI21_X1 U20960 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n18886), .A(n17737), .ZN(
        n17739) );
  OAI222_X1 U20961 ( .A1(n18883), .A2(n18807), .B1(n17740), .B2(n17739), .C1(
        n18832), .C2(n17738), .ZN(P3_U2723) );
  INV_X1 U20962 ( .A(n18998), .ZN(n17741) );
  NOR2_X1 U20963 ( .A1(n17743), .A2(n19184), .ZN(n17751) );
  NAND3_X1 U20964 ( .A1(n17907), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n17762) );
  INV_X1 U20965 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n17881) );
  AND2_X1 U20966 ( .A1(n19030), .A2(n17871), .ZN(n17746) );
  INV_X1 U20967 ( .A(n17746), .ZN(n17745) );
  OAI21_X1 U20968 ( .B1(n19184), .B2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n17744) );
  OAI211_X1 U20969 ( .C1(n17762), .C2(n17881), .A(n17745), .B(n17744), .ZN(
        n17750) );
  NAND2_X1 U20970 ( .A1(n17871), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n17754) );
  NAND2_X1 U20971 ( .A1(n17762), .A2(n17754), .ZN(n17747) );
  OAI21_X1 U20972 ( .B1(n17763), .B2(n17747), .A(n17746), .ZN(n17749) );
  NAND3_X1 U20973 ( .A1(n17747), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n17748) );
  OAI211_X1 U20974 ( .C1(n17751), .C2(n17750), .A(n17749), .B(n17748), .ZN(
        n17876) );
  INV_X1 U20975 ( .A(n17884), .ZN(n17879) );
  NAND2_X1 U20976 ( .A1(n17879), .A2(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n17752) );
  NAND2_X1 U20977 ( .A1(n17881), .A2(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n17863) );
  OAI211_X1 U20978 ( .C1(n17879), .C2(n17754), .A(n17752), .B(n17863), .ZN(
        n17874) );
  OR2_X1 U20979 ( .A1(n19148), .A2(n17753), .ZN(n17770) );
  XNOR2_X1 U20980 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(
        P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n17759) );
  INV_X1 U20981 ( .A(n17754), .ZN(n17868) );
  NAND2_X1 U20982 ( .A1(n17883), .A2(n17868), .ZN(n17755) );
  OAI211_X1 U20983 ( .C1(n17883), .C2(n17871), .A(n17755), .B(n17863), .ZN(
        n17865) );
  INV_X1 U20984 ( .A(n17756), .ZN(n17757) );
  NAND2_X1 U20985 ( .A1(n17758), .A2(n17757), .ZN(n17767) );
  AOI21_X1 U20986 ( .B1(n19141), .B2(n17874), .A(n17760), .ZN(n17761) );
  OAI21_X1 U20987 ( .B1(n17876), .B2(n19109), .A(n17761), .ZN(P3_U2799) );
  NAND2_X1 U20988 ( .A1(n17763), .A2(n17762), .ZN(n17764) );
  XNOR2_X1 U20989 ( .A(n17764), .B(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n17888) );
  INV_X1 U20990 ( .A(n17765), .ZN(n17766) );
  NAND2_X1 U20991 ( .A1(n17766), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n17861) );
  NOR3_X1 U20992 ( .A1(n17785), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n17861), .ZN(n17772) );
  NOR2_X1 U20993 ( .A1(n19442), .A2(n20123), .ZN(n17880) );
  AOI21_X1 U20994 ( .B1(n19067), .B2(n18211), .A(n17880), .ZN(n17769) );
  NAND2_X1 U20995 ( .A1(n17767), .A2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n17768) );
  OAI211_X1 U20996 ( .C1(n17770), .C2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n17769), .B(n17768), .ZN(n17771) );
  AOI211_X1 U20997 ( .C1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .C2(n17773), .A(
        n17772), .B(n17771), .ZN(n17774) );
  OAI21_X1 U20998 ( .B1(n17888), .B2(n19109), .A(n17774), .ZN(P3_U2800) );
  NAND2_X1 U20999 ( .A1(n17775), .A2(n10490), .ZN(n17776) );
  MUX2_X1 U21000 ( .A(n17776), .B(n10490), .S(n19184), .Z(n17777) );
  NAND2_X1 U21001 ( .A1(n17777), .A2(n10023), .ZN(n17942) );
  NAND2_X1 U21002 ( .A1(n17778), .A2(n18243), .ZN(n17783) );
  INV_X1 U21003 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n17779) );
  NOR2_X1 U21004 ( .A1(n19442), .A2(n17779), .ZN(n17924) );
  AOI21_X1 U21005 ( .B1(n19067), .B2(n18242), .A(n17924), .ZN(n17782) );
  NAND2_X1 U21006 ( .A1(n17780), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17781) );
  OAI211_X1 U21007 ( .C1(n19148), .C2(n17783), .A(n17782), .B(n17781), .ZN(
        n17787) );
  AOI21_X1 U21008 ( .B1(n17937), .B2(n17785), .A(n17784), .ZN(n17786) );
  NOR2_X1 U21009 ( .A1(n17787), .A2(n17786), .ZN(n17788) );
  OAI21_X1 U21010 ( .B1(n17942), .B2(n19109), .A(n17788), .ZN(P3_U2803) );
  INV_X1 U21011 ( .A(n17789), .ZN(n17790) );
  AOI21_X1 U21012 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n17791), .A(
        n17790), .ZN(n17953) );
  NAND2_X1 U21013 ( .A1(n19275), .A2(n17943), .ZN(n19033) );
  NAND2_X1 U21014 ( .A1(n19141), .A2(n19043), .ZN(n17792) );
  NAND3_X1 U21015 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n19033), .A3(
        n17792), .ZN(n17793) );
  OAI21_X1 U21016 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n17794), .A(
        n17793), .ZN(n17799) );
  NOR2_X1 U21017 ( .A1(n19148), .A2(n11529), .ZN(n19022) );
  INV_X1 U21018 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n21690) );
  AND2_X1 U21019 ( .A1(n11529), .A2(n19945), .ZN(n19041) );
  AOI211_X1 U21020 ( .C1(n19143), .C2(n17795), .A(n19237), .B(n19041), .ZN(
        n19038) );
  OAI21_X1 U21021 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n19053), .A(
        n19038), .ZN(n19011) );
  OAI22_X1 U21022 ( .A1(n19442), .A2(n21849), .B1(n19159), .B2(n17796), .ZN(
        n17797) );
  AOI221_X1 U21023 ( .B1(n19022), .B2(n21690), .C1(n19011), .C2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(n17797), .ZN(n17798) );
  OAI211_X1 U21024 ( .C1(n17953), .C2(n19109), .A(n17799), .B(n17798), .ZN(
        P3_U2806) );
  XOR2_X1 U21025 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B(n17800), .Z(
        n17972) );
  NAND2_X1 U21026 ( .A1(n19426), .A2(n19275), .ZN(n17802) );
  NAND2_X1 U21027 ( .A1(n19141), .A2(n19423), .ZN(n17801) );
  NAND2_X1 U21028 ( .A1(n17802), .A2(n17801), .ZN(n17845) );
  NOR2_X1 U21029 ( .A1(n19189), .A2(n19325), .ZN(n19135) );
  AOI21_X1 U21030 ( .B1(n19275), .B2(n19385), .A(n19135), .ZN(n19086) );
  OAI21_X1 U21031 ( .B1(n19123), .B2(n19110), .A(n19086), .ZN(n19120) );
  NOR2_X1 U21032 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n10019), .ZN(
        n17970) );
  INV_X1 U21033 ( .A(n17970), .ZN(n17805) );
  NOR2_X1 U21034 ( .A1(n18353), .A2(n17808), .ZN(n19099) );
  AOI21_X1 U21035 ( .B1(n18353), .B2(n17808), .A(n19099), .ZN(n18356) );
  NOR2_X1 U21036 ( .A1(n19442), .A2(n20099), .ZN(n17969) );
  NAND2_X1 U21037 ( .A1(n11533), .A2(n19945), .ZN(n19079) );
  NAND2_X1 U21038 ( .A1(n11533), .A2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n19100) );
  AOI21_X1 U21039 ( .B1(n19239), .B2(n19100), .A(n19237), .ZN(n19097) );
  AOI21_X1 U21040 ( .B1(n18353), .B2(n19079), .A(n19097), .ZN(n17803) );
  AOI211_X1 U21041 ( .C1(n18356), .C2(n19243), .A(n17969), .B(n17803), .ZN(
        n17804) );
  OAI21_X1 U21042 ( .B1(n19123), .B2(n17805), .A(n17804), .ZN(n17806) );
  AOI21_X1 U21043 ( .B1(n19120), .B2(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n17806), .ZN(n17807) );
  OAI21_X1 U21044 ( .B1(n19109), .B2(n17972), .A(n17807), .ZN(P3_U2813) );
  INV_X1 U21045 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n19128) );
  NOR2_X1 U21046 ( .A1(n18562), .A2(n17810), .ZN(n18379) );
  INV_X1 U21047 ( .A(n18379), .ZN(n18380) );
  NOR2_X1 U21048 ( .A1(n19128), .A2(n18380), .ZN(n17809) );
  OAI21_X1 U21049 ( .B1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n17809), .A(
        n17808), .ZN(n18369) );
  AOI21_X1 U21050 ( .B1(n19239), .B2(n17810), .A(n19237), .ZN(n17820) );
  OAI21_X1 U21051 ( .B1(n18379), .B2(n19098), .A(n17820), .ZN(n19127) );
  AOI22_X1 U21052 ( .A1(n19494), .A2(P3_REIP_REG_16__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n19127), .ZN(n17813) );
  NOR2_X1 U21053 ( .A1(n19148), .A2(n17810), .ZN(n19129) );
  OAI211_X1 U21054 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n19129), .B(n17811), .ZN(n17812) );
  OAI211_X1 U21055 ( .C1(n19159), .C2(n18369), .A(n17813), .B(n17812), .ZN(
        n17814) );
  AOI21_X1 U21056 ( .B1(n19050), .B2(n10019), .A(n17814), .ZN(n17818) );
  OAI21_X1 U21057 ( .B1(n19325), .B2(n19030), .A(n17815), .ZN(n17816) );
  XNOR2_X1 U21058 ( .A(n17816), .B(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n19381) );
  NAND2_X1 U21059 ( .A1(n19381), .A2(n19191), .ZN(n17817) );
  OAI211_X1 U21060 ( .C1(n19086), .C2(n10019), .A(n17818), .B(n17817), .ZN(
        P3_U2814) );
  INV_X1 U21061 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n18401) );
  NAND2_X1 U21062 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17819), .ZN(
        n18402) );
  AOI21_X1 U21063 ( .B1(n18401), .B2(n18402), .A(n18379), .ZN(n18393) );
  AOI21_X1 U21064 ( .B1(n17819), .B2(n19945), .A(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17821) );
  OAI22_X1 U21065 ( .A1(n17821), .A2(n17820), .B1(n19442), .B2(n20093), .ZN(
        n17822) );
  AOI21_X1 U21066 ( .B1(n18393), .B2(n19243), .A(n17822), .ZN(n17823) );
  OAI21_X1 U21067 ( .B1(n17824), .B2(n19267), .A(n17823), .ZN(n17825) );
  AOI21_X1 U21068 ( .B1(n19141), .B2(n17826), .A(n17825), .ZN(n17827) );
  OAI21_X1 U21069 ( .B1(n19109), .B2(n17828), .A(n17827), .ZN(P3_U2816) );
  NAND2_X1 U21070 ( .A1(n19130), .A2(n19432), .ZN(n17830) );
  NAND3_X1 U21071 ( .A1(n9830), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(
        n17830), .ZN(n17829) );
  OAI211_X1 U21072 ( .C1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n17830), .A(
        n17829), .B(n19164), .ZN(n19421) );
  INV_X1 U21073 ( .A(n19421), .ZN(n17842) );
  INV_X1 U21074 ( .A(n17845), .ZN(n19175) );
  OAI22_X1 U21075 ( .A1(n19426), .A2(n19267), .B1(n19423), .B2(n19189), .ZN(
        n17844) );
  INV_X1 U21076 ( .A(n17844), .ZN(n17831) );
  OAI21_X1 U21077 ( .B1(n19175), .B2(n19432), .A(n17831), .ZN(n19177) );
  NAND2_X1 U21078 ( .A1(n19432), .A2(n17832), .ZN(n19437) );
  INV_X1 U21079 ( .A(n18426), .ZN(n17833) );
  NOR3_X1 U21080 ( .A1(n18562), .A2(n19217), .A3(n19218), .ZN(n18491) );
  NAND2_X1 U21081 ( .A1(n17833), .A2(n18491), .ZN(n18441) );
  NAND2_X1 U21082 ( .A1(n19146), .A2(n18491), .ZN(n19142) );
  INV_X1 U21083 ( .A(n19142), .ZN(n18418) );
  AOI21_X1 U21084 ( .B1(n17834), .B2(n18441), .A(n18418), .ZN(n18429) );
  INV_X1 U21085 ( .A(n19147), .ZN(n17836) );
  INV_X1 U21086 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n18462) );
  NOR3_X1 U21087 ( .A1(n19217), .A2(n19218), .A3(n19594), .ZN(n19199) );
  NAND2_X1 U21088 ( .A1(n17849), .A2(n19199), .ZN(n17846) );
  NOR2_X1 U21089 ( .A1(n18462), .A2(n17846), .ZN(n19179) );
  NAND2_X1 U21090 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n19179), .ZN(
        n19178) );
  NAND2_X1 U21091 ( .A1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n19278), .ZN(
        n17835) );
  AOI22_X1 U21092 ( .A1(n17836), .A2(n19945), .B1(n19178), .B2(n17835), .ZN(
        n17838) );
  NOR2_X1 U21093 ( .A1(n19442), .A2(n20087), .ZN(n17837) );
  AOI211_X1 U21094 ( .C1(n18429), .C2(n19243), .A(n17838), .B(n17837), .ZN(
        n17839) );
  OAI21_X1 U21095 ( .B1(n19175), .B2(n19437), .A(n17839), .ZN(n17840) );
  AOI21_X1 U21096 ( .B1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n19177), .A(
        n17840), .ZN(n17841) );
  OAI21_X1 U21097 ( .B1(n17842), .B2(n19109), .A(n17841), .ZN(P3_U2819) );
  INV_X1 U21098 ( .A(n19130), .ZN(n19173) );
  NAND3_X1 U21099 ( .A1(n19173), .A2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(
        n9752), .ZN(n17843) );
  OAI211_X1 U21100 ( .C1(n19173), .C2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n17843), .B(n19172), .ZN(n19459) );
  INV_X1 U21101 ( .A(n19459), .ZN(n17854) );
  MUX2_X1 U21102 ( .A(n17845), .B(n17844), .S(
        P3_INSTADDRPOINTER_REG_9__SCAN_IN), .Z(n17852) );
  INV_X1 U21103 ( .A(n17846), .ZN(n17847) );
  AOI21_X1 U21104 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n19278), .A(
        n17847), .ZN(n17850) );
  INV_X1 U21105 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n18470) );
  NAND3_X1 U21106 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17848), .A3(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n18478) );
  NOR2_X1 U21107 ( .A1(n18470), .A2(n18478), .ZN(n18466) );
  NAND3_X1 U21108 ( .A1(n17849), .A2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A3(
        n18491), .ZN(n18443) );
  OAI21_X1 U21109 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n18466), .A(
        n18443), .ZN(n18454) );
  OAI22_X1 U21110 ( .A1(n19179), .A2(n17850), .B1(n19281), .B2(n18454), .ZN(
        n17851) );
  NOR2_X1 U21111 ( .A1(n19442), .A2(n20084), .ZN(n19458) );
  NOR3_X1 U21112 ( .A1(n17852), .A2(n17851), .A3(n19458), .ZN(n17853) );
  OAI21_X1 U21113 ( .B1(n17854), .B2(n19109), .A(n17853), .ZN(P3_U2821) );
  NAND2_X1 U21114 ( .A1(n17856), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17905) );
  NAND2_X1 U21115 ( .A1(n19336), .A2(n17855), .ZN(n17963) );
  NOR2_X1 U21116 ( .A1(n19290), .A2(n17963), .ZN(n17857) );
  NAND2_X1 U21117 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n17857), .ZN(
        n17930) );
  INV_X1 U21118 ( .A(n19336), .ZN(n17959) );
  NOR2_X1 U21119 ( .A1(n17959), .A2(n19401), .ZN(n17866) );
  NAND2_X1 U21120 ( .A1(n19110), .A2(n17866), .ZN(n19311) );
  NOR2_X1 U21121 ( .A1(n19027), .A2(n19311), .ZN(n19295) );
  AOI21_X1 U21122 ( .B1(n17856), .B2(n19295), .A(n19536), .ZN(n17927) );
  AOI221_X1 U21123 ( .B1(n17905), .B2(n19428), .C1(n17930), .C2(n19428), .A(
        n17927), .ZN(n17860) );
  NAND2_X1 U21124 ( .A1(n17857), .A2(n17856), .ZN(n17858) );
  NAND2_X1 U21125 ( .A1(n19454), .A2(n17858), .ZN(n17859) );
  NAND2_X1 U21126 ( .A1(n17860), .A2(n17859), .ZN(n17892) );
  AOI211_X1 U21127 ( .C1(n19467), .C2(n17861), .A(n19522), .B(n17892), .ZN(
        n17862) );
  NOR2_X1 U21128 ( .A1(n17862), .A2(n19494), .ZN(n17885) );
  INV_X1 U21129 ( .A(n17885), .ZN(n17872) );
  INV_X1 U21130 ( .A(n19530), .ZN(n19322) );
  INV_X1 U21131 ( .A(n19470), .ZN(n19514) );
  NOR2_X1 U21132 ( .A1(n19514), .A2(n17863), .ZN(n17864) );
  AOI211_X1 U21133 ( .C1(n19322), .C2(n17865), .A(n9843), .B(n17864), .ZN(
        n17870) );
  INV_X1 U21134 ( .A(n17963), .ZN(n19313) );
  AND2_X1 U21135 ( .A1(n20023), .A2(n17866), .ZN(n17902) );
  AOI21_X1 U21136 ( .B1(n19313), .B2(n19454), .A(n17902), .ZN(n17867) );
  OAI22_X1 U21137 ( .A1(n19451), .A2(n17930), .B1(n17867), .B2(n19290), .ZN(
        n17877) );
  NOR3_X1 U21138 ( .A1(n19522), .A2(n17893), .A3(n17905), .ZN(n17878) );
  NAND4_X1 U21139 ( .A1(n17877), .A2(n17878), .A3(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A4(n17868), .ZN(n17869) );
  OAI211_X1 U21140 ( .C1(n17872), .C2(n17871), .A(n17870), .B(n17869), .ZN(
        n17873) );
  AOI21_X1 U21141 ( .B1(n17874), .B2(n17954), .A(n17873), .ZN(n17875) );
  OAI21_X1 U21142 ( .B1(n17876), .B2(n19364), .A(n17875), .ZN(P3_U2831) );
  AOI22_X1 U21143 ( .A1(n17878), .A2(n17877), .B1(n19322), .B2(n17914), .ZN(
        n17889) );
  OAI22_X1 U21144 ( .A1(n17879), .A2(n19324), .B1(n17889), .B2(n17899), .ZN(
        n17882) );
  AOI21_X1 U21145 ( .B1(n17882), .B2(n17881), .A(n17880), .ZN(n17887) );
  OAI22_X1 U21146 ( .A1(n17884), .A2(n19324), .B1(n17883), .B2(n19530), .ZN(
        n17890) );
  OAI21_X1 U21147 ( .B1(n17890), .B2(n17885), .A(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n17886) );
  OAI211_X1 U21148 ( .C1(n17888), .C2(n19364), .A(n17887), .B(n17886), .ZN(
        P3_U2832) );
  OAI21_X1 U21149 ( .B1(n17910), .B2(n19324), .A(n17889), .ZN(n17898) );
  INV_X1 U21150 ( .A(n17890), .ZN(n17895) );
  OR2_X1 U21151 ( .A1(n19454), .A2(n20023), .ZN(n19439) );
  AND2_X1 U21152 ( .A1(n19439), .A2(n17937), .ZN(n17891) );
  OR3_X1 U21153 ( .A1(n17892), .A2(n17891), .A3(n19527), .ZN(n17911) );
  AOI22_X1 U21154 ( .A1(n17911), .A2(n19442), .B1(n19470), .B2(n17893), .ZN(
        n17894) );
  AOI21_X1 U21155 ( .B1(n17895), .B2(n17894), .A(n17899), .ZN(n17896) );
  AOI211_X1 U21156 ( .C1(n17899), .C2(n17898), .A(n17897), .B(n17896), .ZN(
        n17900) );
  OAI21_X1 U21157 ( .B1(n17901), .B2(n19364), .A(n17900), .ZN(P3_U2833) );
  INV_X1 U21158 ( .A(n17964), .ZN(n19476) );
  NAND3_X1 U21159 ( .A1(n19426), .A2(n19336), .A3(n20021), .ZN(n17903) );
  AOI21_X1 U21160 ( .B1(n19313), .B2(n19539), .A(n17902), .ZN(n19292) );
  OAI211_X1 U21161 ( .C1(n19476), .C2(n17904), .A(n17903), .B(n19292), .ZN(
        n19327) );
  NAND2_X1 U21162 ( .A1(n19327), .A2(n19110), .ZN(n17936) );
  NOR3_X1 U21163 ( .A1(n19335), .A2(n19027), .A3(n17905), .ZN(n17906) );
  AOI21_X1 U21164 ( .B1(n17907), .B2(n19545), .A(n17906), .ZN(n17923) );
  NOR4_X1 U21165 ( .A1(n17909), .A2(n17908), .A3(n17907), .A4(n20016), .ZN(
        n17916) );
  NAND2_X1 U21166 ( .A1(n17910), .A2(n17964), .ZN(n17913) );
  INV_X1 U21167 ( .A(n17911), .ZN(n17912) );
  OAI211_X1 U21168 ( .C1(n17914), .C2(n19543), .A(n17913), .B(n17912), .ZN(
        n17915) );
  OAI211_X1 U21169 ( .C1(n17916), .C2(n17915), .A(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n19442), .ZN(n17922) );
  NOR2_X1 U21170 ( .A1(n19364), .A2(n17917), .ZN(n17919) );
  AOI21_X1 U21171 ( .B1(n17920), .B2(n17919), .A(n17918), .ZN(n17921) );
  OAI211_X1 U21172 ( .C1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .C2(n17923), .A(
        n17922), .B(n17921), .ZN(P3_U2834) );
  AOI21_X1 U21173 ( .B1(n19527), .B2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n17924), .ZN(n17941) );
  INV_X1 U21174 ( .A(n17925), .ZN(n17935) );
  OAI22_X1 U21175 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n19314), .B1(
        n17926), .B2(n19451), .ZN(n17928) );
  AOI211_X1 U21176 ( .C1(n20021), .C2(n17929), .A(n17928), .B(n17927), .ZN(
        n17934) );
  OAI21_X1 U21177 ( .B1(n19428), .B2(n19060), .A(n17930), .ZN(n19319) );
  INV_X1 U21178 ( .A(n19319), .ZN(n17932) );
  AOI21_X1 U21179 ( .B1(n19326), .B2(n19313), .A(n19314), .ZN(n17931) );
  AOI21_X1 U21180 ( .B1(n17932), .B2(n19532), .A(n17931), .ZN(n17945) );
  OAI21_X1 U21181 ( .B1(n19465), .B2(n19296), .A(n17945), .ZN(n19297) );
  INV_X1 U21182 ( .A(n19297), .ZN(n17933) );
  OAI211_X1 U21183 ( .C1(n17935), .C2(n19476), .A(n17934), .B(n17933), .ZN(
        n19282) );
  OAI21_X1 U21184 ( .B1(n19314), .B2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n17939) );
  NOR2_X1 U21185 ( .A1(n19027), .A2(n17936), .ZN(n19307) );
  NAND4_X1 U21186 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A4(n19307), .ZN(n19284) );
  OAI21_X1 U21187 ( .B1(n19284), .B2(n19289), .A(n17937), .ZN(n17938) );
  OAI211_X1 U21188 ( .C1(n19282), .C2(n17939), .A(n17938), .B(n19546), .ZN(
        n17940) );
  OAI211_X1 U21189 ( .C1(n17942), .C2(n19364), .A(n17941), .B(n17940), .ZN(
        P3_U2835) );
  AOI22_X1 U21190 ( .A1(n20021), .A2(n17943), .B1(n17964), .B2(n19043), .ZN(
        n17944) );
  NAND3_X1 U21191 ( .A1(n17945), .A2(n17944), .A3(n19551), .ZN(n17948) );
  INV_X1 U21192 ( .A(n19295), .ZN(n17946) );
  AOI211_X1 U21193 ( .C1(n20023), .C2(n17946), .A(n19035), .B(n17948), .ZN(
        n17947) );
  NOR2_X1 U21194 ( .A1(n19494), .A2(n17947), .ZN(n19306) );
  OAI211_X1 U21195 ( .C1(n17948), .C2(n19467), .A(n19306), .B(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17952) );
  NOR3_X1 U21196 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17949), .A3(
        n19335), .ZN(n17950) );
  AOI21_X1 U21197 ( .B1(n19494), .B2(P3_REIP_REG_24__SCAN_IN), .A(n17950), 
        .ZN(n17951) );
  OAI211_X1 U21198 ( .C1(n17953), .C2(n19364), .A(n17952), .B(n17951), .ZN(
        P3_U2838) );
  NAND2_X1 U21199 ( .A1(n19426), .A2(n19322), .ZN(n17958) );
  NAND2_X1 U21200 ( .A1(n19423), .A2(n17954), .ZN(n17957) );
  NAND2_X1 U21201 ( .A1(n19546), .A2(n19386), .ZN(n17956) );
  NOR2_X1 U21202 ( .A1(n17959), .A2(n19461), .ZN(n19366) );
  INV_X1 U21203 ( .A(n19385), .ZN(n17961) );
  NOR2_X1 U21204 ( .A1(n19325), .A2(n19476), .ZN(n19392) );
  INV_X1 U21205 ( .A(n19392), .ZN(n17960) );
  OAI211_X1 U21206 ( .C1(n19543), .C2(n17961), .A(n17960), .B(n19546), .ZN(
        n19380) );
  NAND2_X1 U21207 ( .A1(n17962), .A2(n19428), .ZN(n19463) );
  INV_X1 U21208 ( .A(n19463), .ZN(n19534) );
  NOR3_X1 U21209 ( .A1(n19534), .A2(n17963), .A3(n10019), .ZN(n17965) );
  OR2_X1 U21210 ( .A1(n20021), .A2(n17964), .ZN(n19351) );
  INV_X1 U21211 ( .A(n19351), .ZN(n19431) );
  OAI22_X1 U21212 ( .A1(n19465), .A2(n17965), .B1(n19110), .B2(n19431), .ZN(
        n17966) );
  AOI211_X1 U21213 ( .C1(n20023), .C2(n19311), .A(n19380), .B(n17966), .ZN(
        n19367) );
  INV_X1 U21214 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17967) );
  NOR3_X1 U21215 ( .A1(n19494), .A2(n19367), .A3(n17967), .ZN(n17968) );
  AOI211_X1 U21216 ( .C1(n17970), .C2(n19366), .A(n17969), .B(n17968), .ZN(
        n17971) );
  OAI21_X1 U21217 ( .B1(n19364), .B2(n17972), .A(n17971), .ZN(P3_U2845) );
  NAND2_X1 U21218 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19715) );
  AOI221_X1 U21219 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n19715), .C1(n17974), 
        .C2(n19715), .A(n17973), .ZN(n19558) );
  NOR2_X1 U21220 ( .A1(n17975), .A2(n11693), .ZN(n17976) );
  OAI21_X1 U21221 ( .B1(n17976), .B2(n19642), .A(n19559), .ZN(n19556) );
  AOI22_X1 U21222 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n19558), .B1(
        n19556), .B2(n11696), .ZN(P3_U2865) );
  NOR2_X1 U21223 ( .A1(n17978), .A2(n17977), .ZN(n20025) );
  NAND3_X1 U21224 ( .A1(n17982), .A2(n17979), .A3(n20025), .ZN(n17980) );
  OAI21_X1 U21225 ( .B1(n17982), .B2(n17981), .A(n17980), .ZN(P3_U3284) );
  NOR4_X1 U21226 ( .A1(n17986), .A2(n17985), .A3(n17984), .A4(n17983), .ZN(
        n17987) );
  NAND2_X1 U21227 ( .A1(n17990), .A2(n17987), .ZN(n17988) );
  OAI21_X1 U21228 ( .B1(n17990), .B2(n17989), .A(n17988), .ZN(P2_U3595) );
  OAI22_X1 U21229 ( .A1(n17993), .A2(n20196), .B1(n17992), .B2(n17991), .ZN(
        n17994) );
  INV_X1 U21230 ( .A(n17994), .ZN(n18007) );
  INV_X1 U21231 ( .A(n17995), .ZN(n17997) );
  AOI21_X1 U21232 ( .B1(n17998), .B2(n17997), .A(n17996), .ZN(n18000) );
  OAI21_X1 U21233 ( .B1(n18000), .B2(n17999), .A(n16085), .ZN(n18005) );
  AOI22_X1 U21234 ( .A1(n20190), .A2(P2_REIP_REG_22__SCAN_IN), .B1(n20188), 
        .B2(P2_EBX_REG_22__SCAN_IN), .ZN(n18004) );
  OR2_X1 U21235 ( .A1(n18001), .A2(n20192), .ZN(n18003) );
  NAND2_X1 U21236 ( .A1(n20189), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n18002) );
  AND4_X1 U21237 ( .A1(n18005), .A2(n18004), .A3(n18003), .A4(n18002), .ZN(
        n18006) );
  NAND2_X1 U21238 ( .A1(n18007), .A2(n18006), .ZN(P2_U2833) );
  INV_X1 U21239 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n21541) );
  NAND2_X1 U21240 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n21541), .ZN(n21531) );
  INV_X1 U21241 ( .A(HOLD), .ZN(n20817) );
  AOI21_X1 U21242 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n21533), .A(n18008), 
        .ZN(n18010) );
  OAI211_X1 U21243 ( .C1(n21541), .C2(n20817), .A(P1_STATE_REG_0__SCAN_IN), 
        .B(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n18009) );
  OAI211_X1 U21244 ( .C1(n21531), .C2(n20817), .A(n18010), .B(n18009), .ZN(
        P1_U3195) );
  INV_X1 U21245 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n18180) );
  NOR2_X1 U21246 ( .A1(n21058), .A2(n18180), .ZN(P1_U2905) );
  AOI21_X1 U21247 ( .B1(n18013), .B2(n18012), .A(n18011), .ZN(n18014) );
  NOR2_X1 U21248 ( .A1(n20748), .A2(n18014), .ZN(n20917) );
  INV_X1 U21249 ( .A(n20917), .ZN(n20918) );
  NOR2_X1 U21250 ( .A1(n18015), .A2(n20918), .ZN(P2_U3047) );
  INV_X1 U21251 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n18016) );
  NOR2_X1 U21252 ( .A1(n21123), .A2(n18016), .ZN(n18029) );
  AOI21_X1 U21253 ( .B1(n21088), .B2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n18029), .ZN(n18021) );
  XNOR2_X1 U21254 ( .A(n18018), .B(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n18019) );
  XNOR2_X1 U21255 ( .A(n18017), .B(n18019), .ZN(n18031) );
  AOI22_X1 U21256 ( .A1(n18031), .A2(n21095), .B1(n21094), .B2(n20983), .ZN(
        n18020) );
  OAI211_X1 U21257 ( .C1(n20985), .C2(n21098), .A(n18021), .B(n18020), .ZN(
        P1_U2993) );
  INV_X1 U21258 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n18022) );
  NOR2_X1 U21259 ( .A1(n21123), .A2(n18022), .ZN(n18037) );
  AOI21_X1 U21260 ( .B1(n21088), .B2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A(
        n18037), .ZN(n18028) );
  INV_X1 U21261 ( .A(n18025), .ZN(n18039) );
  INV_X1 U21262 ( .A(n20988), .ZN(n18026) );
  AOI22_X1 U21263 ( .A1(n18039), .A2(n21095), .B1(n21094), .B2(n18026), .ZN(
        n18027) );
  OAI211_X1 U21264 ( .C1(n20997), .C2(n21098), .A(n18028), .B(n18027), .ZN(
        P1_U2994) );
  AOI21_X1 U21265 ( .B1(n21135), .B2(n20976), .A(n18029), .ZN(n18033) );
  AOI22_X1 U21266 ( .A1(n18031), .A2(n21110), .B1(n18030), .B2(n18034), .ZN(
        n18032) );
  OAI211_X1 U21267 ( .C1(n18035), .C2(n18034), .A(n18033), .B(n18032), .ZN(
        P1_U3025) );
  NAND2_X1 U21268 ( .A1(n18036), .A2(n21100), .ZN(n21115) );
  AOI21_X1 U21269 ( .B1(n20991), .B2(n21135), .A(n18037), .ZN(n18041) );
  AOI22_X1 U21270 ( .A1(n18039), .A2(n21110), .B1(n18038), .B2(
        P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n18040) );
  OAI211_X1 U21271 ( .C1(n21115), .C2(n18042), .A(n18041), .B(n18040), .ZN(
        P1_U3026) );
  OR3_X1 U21272 ( .A1(n18044), .A2(n18043), .A3(n21602), .ZN(n18045) );
  OAI21_X1 U21273 ( .B1(n21597), .B2(n12613), .A(n18045), .ZN(P1_U3468) );
  AOI21_X1 U21274 ( .B1(n18048), .B2(n18047), .A(n18046), .ZN(n18050) );
  AOI211_X1 U21275 ( .C1(n18052), .C2(n18051), .A(n18050), .B(n18049), .ZN(
        P1_U3162) );
  OAI21_X1 U21276 ( .B1(n18054), .B2(n21719), .A(n18053), .ZN(P1_U3466) );
  XNOR2_X1 U21277 ( .A(n18056), .B(n18055), .ZN(n18057) );
  NAND2_X1 U21278 ( .A1(n18058), .A2(P2_REIP_REG_7__SCAN_IN), .ZN(n18074) );
  OAI21_X1 U21279 ( .B1(n18060), .B2(n18059), .A(n18074), .ZN(n18061) );
  AOI21_X1 U21280 ( .B1(n18063), .B2(n18062), .A(n18061), .ZN(n18072) );
  INV_X1 U21281 ( .A(n18064), .ZN(n18069) );
  OAI21_X1 U21282 ( .B1(n18066), .B2(n18068), .A(n18065), .ZN(n18067) );
  OAI21_X1 U21283 ( .B1(n18069), .B2(n18068), .A(n18067), .ZN(n18081) );
  AOI22_X1 U21284 ( .A1(n18081), .A2(n18070), .B1(n20252), .B2(n18080), .ZN(
        n18071) );
  OAI211_X1 U21285 ( .C1(n20256), .C2(n18084), .A(n18072), .B(n18071), .ZN(
        P2_U3007) );
  INV_X1 U21286 ( .A(n18073), .ZN(n18079) );
  OAI21_X1 U21287 ( .B1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n18075), .A(
        n18074), .ZN(n18078) );
  AND3_X1 U21288 ( .A1(n18076), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(
        n20257), .ZN(n18077) );
  AOI211_X1 U21289 ( .C1(n18079), .C2(n20277), .A(n18078), .B(n18077), .ZN(
        n18083) );
  AOI22_X1 U21290 ( .A1(n18081), .A2(n20279), .B1(n20280), .B2(n18080), .ZN(
        n18082) );
  OAI211_X1 U21291 ( .C1(n20290), .C2(n18084), .A(n18083), .B(n18082), .ZN(
        P2_U3039) );
  NAND3_X1 U21292 ( .A1(n18086), .A2(n10158), .A3(n20267), .ZN(n18089) );
  AOI21_X1 U21293 ( .B1(n10798), .B2(n20280), .A(n18087), .ZN(n18088) );
  OAI211_X1 U21294 ( .C1(n18091), .C2(n18090), .A(n18089), .B(n18088), .ZN(
        n18092) );
  AOI21_X1 U21295 ( .B1(n18093), .B2(n20279), .A(n18092), .ZN(n18094) );
  OAI221_X1 U21296 ( .B1(n20261), .B2(n18096), .C1(n20261), .C2(n18095), .A(
        n18094), .ZN(P2_U3043) );
  NOR3_X1 U21297 ( .A1(P3_BE_N_REG_3__SCAN_IN), .A2(P3_W_R_N_REG_SCAN_IN), 
        .A3(P3_BE_N_REG_0__SCAN_IN), .ZN(n18098) );
  NOR4_X1 U21298 ( .A1(P3_BE_N_REG_1__SCAN_IN), .A2(P3_BE_N_REG_2__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n18097) );
  INV_X2 U21299 ( .A(n18179), .ZN(U215) );
  NAND4_X1 U21300 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n18098), .A3(n18097), .A4(
        U215), .ZN(U213) );
  INV_X1 U21301 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n20210) );
  INV_X2 U21302 ( .A(U214), .ZN(n18144) );
  OAI222_X1 U21303 ( .A1(U212), .A2(n20210), .B1(n18148), .B2(n18100), .C1(
        U214), .C2(n18180), .ZN(U216) );
  AOI22_X1 U21304 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(n18142), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n18144), .ZN(n18101) );
  OAI21_X1 U21305 ( .B1(n16749), .B2(n18148), .A(n18101), .ZN(U217) );
  INV_X1 U21306 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n18103) );
  AOI22_X1 U21307 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(n18142), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n18144), .ZN(n18102) );
  OAI21_X1 U21308 ( .B1(n18103), .B2(n18148), .A(n18102), .ZN(U218) );
  INV_X1 U21309 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n18105) );
  AOI22_X1 U21310 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(n18142), .B1(
        P1_DATAO_REG_28__SCAN_IN), .B2(n18144), .ZN(n18104) );
  OAI21_X1 U21311 ( .B1(n18105), .B2(n18148), .A(n18104), .ZN(U219) );
  INV_X1 U21312 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n18106) );
  OAI222_X1 U21313 ( .A1(U214), .A2(n18106), .B1(n18148), .B2(n21718), .C1(
        U212), .C2(n18173), .ZN(U220) );
  INV_X1 U21314 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n18108) );
  AOI22_X1 U21315 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(n18142), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n18144), .ZN(n18107) );
  OAI21_X1 U21316 ( .B1(n18108), .B2(n18148), .A(n18107), .ZN(U221) );
  AOI22_X1 U21317 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(n18142), .B1(
        P1_DATAO_REG_25__SCAN_IN), .B2(n18144), .ZN(n18109) );
  OAI21_X1 U21318 ( .B1(n18110), .B2(n18148), .A(n18109), .ZN(U222) );
  INV_X1 U21319 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n18112) );
  AOI22_X1 U21320 ( .A1(P2_DATAO_REG_24__SCAN_IN), .A2(n18142), .B1(
        P1_DATAO_REG_24__SCAN_IN), .B2(n18144), .ZN(n18111) );
  OAI21_X1 U21321 ( .B1(n18112), .B2(n18148), .A(n18111), .ZN(U223) );
  INV_X1 U21322 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n18114) );
  AOI22_X1 U21323 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(n18142), .B1(
        P1_DATAO_REG_23__SCAN_IN), .B2(n18144), .ZN(n18113) );
  OAI21_X1 U21324 ( .B1(n18114), .B2(n18148), .A(n18113), .ZN(U224) );
  INV_X1 U21325 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n18116) );
  AOI22_X1 U21326 ( .A1(P2_DATAO_REG_22__SCAN_IN), .A2(n18142), .B1(
        P1_DATAO_REG_22__SCAN_IN), .B2(n18144), .ZN(n18115) );
  OAI21_X1 U21327 ( .B1(n18116), .B2(n18148), .A(n18115), .ZN(U225) );
  INV_X1 U21328 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n18118) );
  AOI22_X1 U21329 ( .A1(P2_DATAO_REG_21__SCAN_IN), .A2(n18142), .B1(
        P1_DATAO_REG_21__SCAN_IN), .B2(n18144), .ZN(n18117) );
  OAI21_X1 U21330 ( .B1(n18118), .B2(n18148), .A(n18117), .ZN(U226) );
  AOI22_X1 U21331 ( .A1(P2_DATAO_REG_20__SCAN_IN), .A2(n18142), .B1(
        P1_DATAO_REG_20__SCAN_IN), .B2(n18144), .ZN(n18119) );
  OAI21_X1 U21332 ( .B1(n21772), .B2(n18148), .A(n18119), .ZN(U227) );
  AOI222_X1 U21333 ( .A1(n18144), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n18145), 
        .B2(BUF1_REG_19__SCAN_IN), .C1(n18142), .C2(P2_DATAO_REG_19__SCAN_IN), 
        .ZN(n18120) );
  INV_X1 U21334 ( .A(n18120), .ZN(U228) );
  AOI222_X1 U21335 ( .A1(n18144), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n18145), 
        .B2(BUF1_REG_18__SCAN_IN), .C1(n18142), .C2(P2_DATAO_REG_18__SCAN_IN), 
        .ZN(n18121) );
  INV_X1 U21336 ( .A(n18121), .ZN(U229) );
  INV_X1 U21337 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n18123) );
  AOI22_X1 U21338 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(n18142), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n18144), .ZN(n18122) );
  OAI21_X1 U21339 ( .B1(n18123), .B2(n18148), .A(n18122), .ZN(U230) );
  AOI22_X1 U21340 ( .A1(P2_DATAO_REG_16__SCAN_IN), .A2(n18142), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n18144), .ZN(n18124) );
  OAI21_X1 U21341 ( .B1(n18125), .B2(n18148), .A(n18124), .ZN(U231) );
  AOI22_X1 U21342 ( .A1(P2_DATAO_REG_15__SCAN_IN), .A2(n18142), .B1(
        P1_DATAO_REG_15__SCAN_IN), .B2(n18144), .ZN(n18126) );
  OAI21_X1 U21343 ( .B1(n14046), .B2(n18148), .A(n18126), .ZN(U232) );
  AOI22_X1 U21344 ( .A1(P2_DATAO_REG_14__SCAN_IN), .A2(n18142), .B1(
        P1_DATAO_REG_14__SCAN_IN), .B2(n18144), .ZN(n18127) );
  OAI21_X1 U21345 ( .B1(n14797), .B2(n18148), .A(n18127), .ZN(U233) );
  AOI22_X1 U21346 ( .A1(P2_DATAO_REG_13__SCAN_IN), .A2(n18142), .B1(
        P1_DATAO_REG_13__SCAN_IN), .B2(n18144), .ZN(n18128) );
  OAI21_X1 U21347 ( .B1(n15207), .B2(n18148), .A(n18128), .ZN(U234) );
  AOI22_X1 U21348 ( .A1(P2_DATAO_REG_12__SCAN_IN), .A2(n18142), .B1(
        P1_DATAO_REG_12__SCAN_IN), .B2(n18144), .ZN(n18129) );
  OAI21_X1 U21349 ( .B1(n18130), .B2(n18148), .A(n18129), .ZN(U235) );
  INV_X1 U21350 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n20222) );
  AOI22_X1 U21351 ( .A1(BUF1_REG_11__SCAN_IN), .A2(n18145), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n18144), .ZN(n18131) );
  OAI21_X1 U21352 ( .B1(n20222), .B2(U212), .A(n18131), .ZN(U236) );
  AOI22_X1 U21353 ( .A1(P2_DATAO_REG_10__SCAN_IN), .A2(n18142), .B1(
        P1_DATAO_REG_10__SCAN_IN), .B2(n18144), .ZN(n18132) );
  OAI21_X1 U21354 ( .B1(n18133), .B2(n18148), .A(n18132), .ZN(U237) );
  INV_X1 U21355 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n18155) );
  AOI22_X1 U21356 ( .A1(BUF1_REG_9__SCAN_IN), .A2(n18145), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n18144), .ZN(n18134) );
  OAI21_X1 U21357 ( .B1(n18155), .B2(U212), .A(n18134), .ZN(U238) );
  AOI22_X1 U21358 ( .A1(P2_DATAO_REG_8__SCAN_IN), .A2(n18142), .B1(
        P1_DATAO_REG_8__SCAN_IN), .B2(n18144), .ZN(n18135) );
  OAI21_X1 U21359 ( .B1(n21684), .B2(n18148), .A(n18135), .ZN(U239) );
  INV_X1 U21360 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n18153) );
  INV_X1 U21361 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n21809) );
  INV_X1 U21362 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n21747) );
  OAI222_X1 U21363 ( .A1(U212), .A2(n18153), .B1(n18148), .B2(n21809), .C1(
        U214), .C2(n21747), .ZN(U240) );
  INV_X1 U21364 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n18137) );
  AOI22_X1 U21365 ( .A1(P2_DATAO_REG_6__SCAN_IN), .A2(n18142), .B1(
        P1_DATAO_REG_6__SCAN_IN), .B2(n18144), .ZN(n18136) );
  OAI21_X1 U21366 ( .B1(n18137), .B2(n18148), .A(n18136), .ZN(U241) );
  INV_X1 U21367 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n18151) );
  AOI22_X1 U21368 ( .A1(BUF1_REG_5__SCAN_IN), .A2(n18145), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(n18144), .ZN(n18138) );
  OAI21_X1 U21369 ( .B1(n18151), .B2(U212), .A(n18138), .ZN(U242) );
  INV_X1 U21370 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n18140) );
  AOI22_X1 U21371 ( .A1(P2_DATAO_REG_4__SCAN_IN), .A2(n18142), .B1(
        P1_DATAO_REG_4__SCAN_IN), .B2(n18144), .ZN(n18139) );
  OAI21_X1 U21372 ( .B1(n18140), .B2(n18148), .A(n18139), .ZN(U243) );
  INV_X1 U21373 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n21732) );
  AOI22_X1 U21374 ( .A1(BUF1_REG_3__SCAN_IN), .A2(n18145), .B1(
        P1_DATAO_REG_3__SCAN_IN), .B2(n18144), .ZN(n18141) );
  OAI21_X1 U21375 ( .B1(n21732), .B2(U212), .A(n18141), .ZN(U244) );
  AOI222_X1 U21376 ( .A1(n18144), .A2(P1_DATAO_REG_2__SCAN_IN), .B1(n18145), 
        .B2(BUF1_REG_2__SCAN_IN), .C1(n18142), .C2(P2_DATAO_REG_2__SCAN_IN), 
        .ZN(n18143) );
  INV_X1 U21377 ( .A(n18143), .ZN(U245) );
  INV_X1 U21378 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n21763) );
  AOI22_X1 U21379 ( .A1(BUF1_REG_1__SCAN_IN), .A2(n18145), .B1(
        P1_DATAO_REG_1__SCAN_IN), .B2(n18144), .ZN(n18146) );
  OAI21_X1 U21380 ( .B1(n21763), .B2(U212), .A(n18146), .ZN(U246) );
  INV_X1 U21381 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n21057) );
  INV_X1 U21382 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n18147) );
  INV_X1 U21383 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n18149) );
  OAI222_X1 U21384 ( .A1(U214), .A2(n21057), .B1(n18148), .B2(n18147), .C1(
        U212), .C2(n18149), .ZN(U247) );
  AOI22_X1 U21385 ( .A1(n18179), .A2(n18149), .B1(n14163), .B2(U215), .ZN(U251) );
  AOI22_X1 U21386 ( .A1(n18179), .A2(n21763), .B1(n13632), .B2(U215), .ZN(U252) );
  INV_X1 U21387 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n21825) );
  AOI22_X1 U21388 ( .A1(n18174), .A2(n21825), .B1(n13655), .B2(U215), .ZN(U253) );
  AOI22_X1 U21389 ( .A1(n18174), .A2(n21732), .B1(n13652), .B2(U215), .ZN(U254) );
  OAI22_X1 U21390 ( .A1(U215), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n18174), .ZN(n18150) );
  INV_X1 U21391 ( .A(n18150), .ZN(U255) );
  AOI22_X1 U21392 ( .A1(n18179), .A2(n18151), .B1(n13643), .B2(U215), .ZN(U256) );
  OAI22_X1 U21393 ( .A1(U215), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n18179), .ZN(n18152) );
  INV_X1 U21394 ( .A(n18152), .ZN(U257) );
  AOI22_X1 U21395 ( .A1(n18179), .A2(n18153), .B1(n13640), .B2(U215), .ZN(U258) );
  OAI22_X1 U21396 ( .A1(U215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n18179), .ZN(n18154) );
  INV_X1 U21397 ( .A(n18154), .ZN(U259) );
  AOI22_X1 U21398 ( .A1(n18179), .A2(n18155), .B1(n13646), .B2(U215), .ZN(U260) );
  OAI22_X1 U21399 ( .A1(U215), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n18179), .ZN(n18156) );
  INV_X1 U21400 ( .A(n18156), .ZN(U261) );
  OAI22_X1 U21401 ( .A1(U215), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n18174), .ZN(n18157) );
  INV_X1 U21402 ( .A(n18157), .ZN(U262) );
  OAI22_X1 U21403 ( .A1(U215), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n18179), .ZN(n18158) );
  INV_X1 U21404 ( .A(n18158), .ZN(U263) );
  OAI22_X1 U21405 ( .A1(U215), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n18174), .ZN(n18159) );
  INV_X1 U21406 ( .A(n18159), .ZN(U264) );
  OAI22_X1 U21407 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n18179), .ZN(n18160) );
  INV_X1 U21408 ( .A(n18160), .ZN(U265) );
  OAI22_X1 U21409 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n18174), .ZN(n18161) );
  INV_X1 U21410 ( .A(n18161), .ZN(U266) );
  OAI22_X1 U21411 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n18179), .ZN(n18162) );
  INV_X1 U21412 ( .A(n18162), .ZN(U267) );
  OAI22_X1 U21413 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n18174), .ZN(n18163) );
  INV_X1 U21414 ( .A(n18163), .ZN(U268) );
  INV_X1 U21415 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n21855) );
  AOI22_X1 U21416 ( .A1(n18179), .A2(n21855), .B1(n16835), .B2(U215), .ZN(U269) );
  AOI22_X1 U21417 ( .A1(n18179), .A2(n18164), .B1(n17727), .B2(U215), .ZN(U270) );
  OAI22_X1 U21418 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n18179), .ZN(n18165) );
  INV_X1 U21419 ( .A(n18165), .ZN(U271) );
  OAI22_X1 U21420 ( .A1(U215), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n18174), .ZN(n18166) );
  INV_X1 U21421 ( .A(n18166), .ZN(U272) );
  OAI22_X1 U21422 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n18174), .ZN(n18167) );
  INV_X1 U21423 ( .A(n18167), .ZN(U273) );
  OAI22_X1 U21424 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n18179), .ZN(n18168) );
  INV_X1 U21425 ( .A(n18168), .ZN(U274) );
  OAI22_X1 U21426 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n18179), .ZN(n18169) );
  INV_X1 U21427 ( .A(n18169), .ZN(U275) );
  OAI22_X1 U21428 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n18179), .ZN(n18170) );
  INV_X1 U21429 ( .A(n18170), .ZN(U276) );
  OAI22_X1 U21430 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n18179), .ZN(n18171) );
  INV_X1 U21431 ( .A(n18171), .ZN(U277) );
  AOI22_X1 U21432 ( .A1(n18174), .A2(n18173), .B1(n16774), .B2(U215), .ZN(U278) );
  OAI22_X1 U21433 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n18179), .ZN(n18175) );
  INV_X1 U21434 ( .A(n18175), .ZN(U279) );
  OAI22_X1 U21435 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n18179), .ZN(n18176) );
  INV_X1 U21436 ( .A(n18176), .ZN(U280) );
  OAI22_X1 U21437 ( .A1(U215), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n18179), .ZN(n18177) );
  INV_X1 U21438 ( .A(n18177), .ZN(U281) );
  AOI22_X1 U21439 ( .A1(n18179), .A2(n20210), .B1(n18178), .B2(U215), .ZN(U282) );
  INV_X1 U21440 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n21879) );
  AOI222_X1 U21441 ( .A1(n18180), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n20210), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .C1(n21879), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n18181) );
  INV_X2 U21442 ( .A(n18183), .ZN(n18182) );
  INV_X1 U21443 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n21823) );
  INV_X1 U21444 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n20844) );
  AOI22_X1 U21445 ( .A1(n18182), .A2(n21823), .B1(n20844), .B2(n18183), .ZN(
        U347) );
  INV_X1 U21446 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n20085) );
  INV_X1 U21447 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n20842) );
  AOI22_X1 U21448 ( .A1(n18182), .A2(n20085), .B1(n20842), .B2(n18183), .ZN(
        U348) );
  INV_X1 U21449 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n20083) );
  INV_X1 U21450 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n20840) );
  AOI22_X1 U21451 ( .A1(n18182), .A2(n20083), .B1(n20840), .B2(n18183), .ZN(
        U349) );
  INV_X1 U21452 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n21775) );
  INV_X1 U21453 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n20838) );
  AOI22_X1 U21454 ( .A1(n18182), .A2(n21775), .B1(n20838), .B2(n18183), .ZN(
        U350) );
  INV_X1 U21455 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n20080) );
  INV_X1 U21456 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n20836) );
  AOI22_X1 U21457 ( .A1(n18182), .A2(n20080), .B1(n20836), .B2(n18183), .ZN(
        U351) );
  INV_X1 U21458 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n20079) );
  INV_X1 U21459 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n20834) );
  AOI22_X1 U21460 ( .A1(n18182), .A2(n20079), .B1(n20834), .B2(n18183), .ZN(
        U352) );
  INV_X1 U21461 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n21865) );
  INV_X1 U21462 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n20833) );
  AOI22_X1 U21463 ( .A1(n18182), .A2(n21865), .B1(n20833), .B2(n18183), .ZN(
        U353) );
  INV_X1 U21464 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n20076) );
  INV_X1 U21465 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n20832) );
  AOI22_X1 U21466 ( .A1(n18182), .A2(n20076), .B1(n20832), .B2(n18183), .ZN(
        U354) );
  INV_X1 U21467 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n20122) );
  INV_X1 U21468 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n20874) );
  AOI22_X1 U21469 ( .A1(n18182), .A2(n20122), .B1(n20874), .B2(n18183), .ZN(
        U355) );
  INV_X1 U21470 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n20119) );
  INV_X1 U21471 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n20872) );
  AOI22_X1 U21472 ( .A1(n18182), .A2(n20119), .B1(n20872), .B2(n18183), .ZN(
        U356) );
  INV_X1 U21473 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n20118) );
  INV_X1 U21474 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n21840) );
  AOI22_X1 U21475 ( .A1(n18182), .A2(n20118), .B1(n21840), .B2(n18183), .ZN(
        U357) );
  INV_X1 U21476 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n20116) );
  INV_X1 U21477 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n20868) );
  AOI22_X1 U21478 ( .A1(n18182), .A2(n20116), .B1(n20868), .B2(n18183), .ZN(
        U358) );
  INV_X1 U21479 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n20115) );
  INV_X1 U21480 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n21748) );
  AOI22_X1 U21481 ( .A1(n18182), .A2(n20115), .B1(n21748), .B2(n18183), .ZN(
        U359) );
  INV_X1 U21482 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n21812) );
  INV_X1 U21483 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n20867) );
  AOI22_X1 U21484 ( .A1(n18182), .A2(n21812), .B1(n20867), .B2(n18183), .ZN(
        U360) );
  INV_X1 U21485 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n20112) );
  INV_X1 U21486 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n20865) );
  AOI22_X1 U21487 ( .A1(n18182), .A2(n20112), .B1(n20865), .B2(n18183), .ZN(
        U361) );
  INV_X1 U21488 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n20110) );
  INV_X1 U21489 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n20863) );
  AOI22_X1 U21490 ( .A1(n18182), .A2(n20110), .B1(n20863), .B2(n18183), .ZN(
        U362) );
  INV_X1 U21491 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n20109) );
  INV_X1 U21492 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n20861) );
  AOI22_X1 U21493 ( .A1(n18182), .A2(n20109), .B1(n20861), .B2(n18183), .ZN(
        U363) );
  INV_X1 U21494 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n20107) );
  INV_X1 U21495 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n20860) );
  AOI22_X1 U21496 ( .A1(n18182), .A2(n20107), .B1(n20860), .B2(n18183), .ZN(
        U364) );
  INV_X1 U21497 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n20075) );
  INV_X1 U21498 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n20831) );
  AOI22_X1 U21499 ( .A1(n18182), .A2(n20075), .B1(n20831), .B2(n18183), .ZN(
        U365) );
  INV_X1 U21500 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n20106) );
  INV_X1 U21501 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n20858) );
  AOI22_X1 U21502 ( .A1(n18182), .A2(n20106), .B1(n20858), .B2(n18183), .ZN(
        U366) );
  INV_X1 U21503 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n20103) );
  INV_X1 U21504 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n20857) );
  AOI22_X1 U21505 ( .A1(n18182), .A2(n20103), .B1(n20857), .B2(n18183), .ZN(
        U367) );
  INV_X1 U21506 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n20102) );
  INV_X1 U21507 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n20856) );
  AOI22_X1 U21508 ( .A1(n18182), .A2(n20102), .B1(n20856), .B2(n18183), .ZN(
        U368) );
  INV_X1 U21509 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n20100) );
  INV_X1 U21510 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n20854) );
  AOI22_X1 U21511 ( .A1(n18182), .A2(n20100), .B1(n20854), .B2(n18183), .ZN(
        U369) );
  INV_X1 U21512 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n20098) );
  INV_X1 U21513 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n20852) );
  AOI22_X1 U21514 ( .A1(n18182), .A2(n20098), .B1(n20852), .B2(n18183), .ZN(
        U370) );
  INV_X1 U21515 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n20096) );
  INV_X1 U21516 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n20850) );
  AOI22_X1 U21517 ( .A1(n18182), .A2(n20096), .B1(n20850), .B2(n18183), .ZN(
        U371) );
  INV_X1 U21518 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n20094) );
  INV_X1 U21519 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n21898) );
  AOI22_X1 U21520 ( .A1(n18182), .A2(n20094), .B1(n21898), .B2(n18183), .ZN(
        U372) );
  INV_X1 U21521 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n20092) );
  INV_X1 U21522 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n20847) );
  AOI22_X1 U21523 ( .A1(n18182), .A2(n20092), .B1(n20847), .B2(n18183), .ZN(
        U373) );
  INV_X1 U21524 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n20090) );
  INV_X1 U21525 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n21691) );
  AOI22_X1 U21526 ( .A1(n18182), .A2(n20090), .B1(n21691), .B2(n18183), .ZN(
        U374) );
  INV_X1 U21527 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n20088) );
  INV_X1 U21528 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n20845) );
  AOI22_X1 U21529 ( .A1(n18182), .A2(n20088), .B1(n20845), .B2(n18183), .ZN(
        U375) );
  INV_X1 U21530 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n20073) );
  INV_X1 U21531 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n20828) );
  AOI22_X1 U21532 ( .A1(n18182), .A2(n20073), .B1(n20828), .B2(n18183), .ZN(
        U376) );
  NOR2_X1 U21533 ( .A1(P3_STATE_REG_2__SCAN_IN), .A2(n20067), .ZN(n20064) );
  OAI22_X1 U21534 ( .A1(n20062), .A2(n20064), .B1(n20067), .B2(
        P3_STATE_REG_1__SCAN_IN), .ZN(n20056) );
  INV_X1 U21535 ( .A(n20056), .ZN(n20132) );
  AOI21_X1 U21536 ( .B1(P3_STATE_REG_0__SCAN_IN), .B2(P3_ADS_N_REG_SCAN_IN), 
        .A(n20132), .ZN(n18184) );
  INV_X1 U21537 ( .A(n18184), .ZN(P3_U2633) );
  INV_X1 U21538 ( .A(n18185), .ZN(n18191) );
  NOR2_X1 U21539 ( .A1(n18937), .A2(n18191), .ZN(n18186) );
  OAI21_X1 U21540 ( .B1(n18186), .B2(n18935), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n18187) );
  OAI21_X1 U21541 ( .B1(n20167), .B2(n20156), .A(n18187), .ZN(P3_U2634) );
  INV_X1 U21542 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n20072) );
  AOI21_X1 U21543 ( .B1(n20067), .B2(n20072), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n18188) );
  AOI22_X1 U21544 ( .A1(n20144), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n18188), 
        .B2(n20164), .ZN(P3_U2635) );
  OAI21_X1 U21545 ( .B1(n20058), .B2(BS16), .A(n20132), .ZN(n20130) );
  OAI21_X1 U21546 ( .B1(n20132), .B2(n18189), .A(n20130), .ZN(P3_U2636) );
  OAI211_X1 U21547 ( .C1(n18937), .C2(n18191), .A(n18190), .B(n20018), .ZN(
        n20028) );
  NAND2_X1 U21548 ( .A1(n18192), .A2(n20028), .ZN(n20148) );
  INV_X1 U21549 ( .A(n20148), .ZN(n18194) );
  OAI21_X1 U21550 ( .B1(n18194), .B2(n19553), .A(n18193), .ZN(P3_U2637) );
  NOR4_X1 U21551 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_21__SCAN_IN), .A3(P3_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_23__SCAN_IN), .ZN(n18198) );
  NOR4_X1 U21552 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_17__SCAN_IN), .A3(P3_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_19__SCAN_IN), .ZN(n18197) );
  NOR4_X1 U21553 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_29__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n18196) );
  NOR4_X1 U21554 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_25__SCAN_IN), .A3(P3_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_27__SCAN_IN), .ZN(n18195) );
  NAND4_X1 U21555 ( .A1(n18198), .A2(n18197), .A3(n18196), .A4(n18195), .ZN(
        n18204) );
  NOR4_X1 U21556 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_3__SCAN_IN), .A3(P3_DATAWIDTH_REG_4__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_6__SCAN_IN), .ZN(n18202) );
  AOI211_X1 U21557 ( .C1(P3_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_10__SCAN_IN), .B(
        P3_DATAWIDTH_REG_5__SCAN_IN), .ZN(n18201) );
  NOR4_X1 U21558 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_13__SCAN_IN), .A3(P3_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_15__SCAN_IN), .ZN(n18200) );
  NOR4_X1 U21559 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_8__SCAN_IN), .A3(P3_DATAWIDTH_REG_9__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_11__SCAN_IN), .ZN(n18199) );
  NAND4_X1 U21560 ( .A1(n18202), .A2(n18201), .A3(n18200), .A4(n18199), .ZN(
        n18203) );
  NOR2_X1 U21561 ( .A1(n18204), .A2(n18203), .ZN(n20143) );
  INV_X1 U21562 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n18206) );
  NOR3_X1 U21563 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n18207) );
  OAI21_X1 U21564 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n18207), .A(n20143), .ZN(
        n18205) );
  OAI21_X1 U21565 ( .B1(n20143), .B2(n18206), .A(n18205), .ZN(P3_U2638) );
  INV_X1 U21566 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20131) );
  AOI21_X1 U21567 ( .B1(n20136), .B2(n20131), .A(n18207), .ZN(n18208) );
  INV_X1 U21568 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20125) );
  INV_X1 U21569 ( .A(n20143), .ZN(n20138) );
  AOI22_X1 U21570 ( .A1(n20143), .A2(n18208), .B1(n20125), .B2(n20138), .ZN(
        P3_U2639) );
  NAND2_X1 U21571 ( .A1(n18580), .A2(n18209), .ZN(n18224) );
  OAI22_X1 U21572 ( .A1(n10506), .A2(n18558), .B1(n20123), .B2(n18228), .ZN(
        n18212) );
  OAI21_X1 U21573 ( .B1(n18581), .B2(n18214), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n18215) );
  OAI211_X1 U21574 ( .C1(P3_EBX_REG_30__SCAN_IN), .C2(n18224), .A(n18216), .B(
        n18215), .ZN(P3_U2641) );
  AOI211_X1 U21575 ( .C1(n18219), .C2(n18218), .A(n18217), .B(n18536), .ZN(
        n18223) );
  NAND3_X1 U21576 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .A3(n18246), .ZN(n18221) );
  OAI22_X1 U21577 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n18221), .B1(n18220), 
        .B2(n18558), .ZN(n18222) );
  AOI211_X1 U21578 ( .C1(P3_EBX_REG_29__SCAN_IN), .C2(n18581), .A(n18223), .B(
        n18222), .ZN(n18227) );
  INV_X1 U21579 ( .A(n18224), .ZN(n18225) );
  OAI21_X1 U21580 ( .B1(n18230), .B2(n21826), .A(n18225), .ZN(n18226) );
  OAI211_X1 U21581 ( .C1(n18228), .C2(n13399), .A(n18227), .B(n18226), .ZN(
        P3_U2642) );
  AOI22_X1 U21582 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n18540), .B1(
        n18581), .B2(P3_EBX_REG_28__SCAN_IN), .ZN(n18239) );
  NAND2_X1 U21583 ( .A1(n18579), .A2(n18229), .ZN(n18251) );
  INV_X1 U21584 ( .A(n18251), .ZN(n18260) );
  AOI211_X1 U21585 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n18247), .A(n18230), .B(
        n18567), .ZN(n18235) );
  AOI211_X1 U21586 ( .C1(n18233), .C2(n18232), .A(n18231), .B(n18536), .ZN(
        n18234) );
  NAND2_X1 U21587 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .ZN(n18236) );
  OAI211_X1 U21588 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(P3_REIP_REG_27__SCAN_IN), .A(n18246), .B(n18236), .ZN(n18237) );
  NAND3_X1 U21589 ( .A1(n18239), .A2(n18238), .A3(n18237), .ZN(P3_U2643) );
  AOI211_X1 U21590 ( .C1(n18242), .C2(n18241), .A(n18240), .B(n18536), .ZN(
        n18245) );
  OAI22_X1 U21591 ( .A1(n18243), .A2(n18558), .B1(n18568), .B2(n18248), .ZN(
        n18244) );
  AOI211_X1 U21592 ( .C1(n18246), .C2(n17779), .A(n18245), .B(n18244), .ZN(
        n18250) );
  OAI211_X1 U21593 ( .C1(n18253), .C2(n18248), .A(n18580), .B(n18247), .ZN(
        n18249) );
  OAI211_X1 U21594 ( .C1(n18251), .C2(n17779), .A(n18250), .B(n18249), .ZN(
        P3_U2644) );
  AOI22_X1 U21595 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n18540), .B1(
        n18581), .B2(P3_EBX_REG_26__SCAN_IN), .ZN(n18262) );
  INV_X1 U21596 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n20113) );
  NAND2_X1 U21597 ( .A1(n18551), .A2(n18252), .ZN(n18267) );
  INV_X1 U21598 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n20114) );
  OAI21_X1 U21599 ( .B1(n20113), .B2(n18267), .A(n20114), .ZN(n18259) );
  AOI211_X1 U21600 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n18270), .A(n18253), .B(
        n18567), .ZN(n18258) );
  AOI211_X1 U21601 ( .C1(n18256), .C2(n18255), .A(n18254), .B(n18536), .ZN(
        n18257) );
  AOI211_X1 U21602 ( .C1(n18260), .C2(n18259), .A(n18258), .B(n18257), .ZN(
        n18261) );
  NAND2_X1 U21603 ( .A1(n18262), .A2(n18261), .ZN(P3_U2645) );
  NAND2_X1 U21604 ( .A1(n18551), .A2(n18284), .ZN(n18298) );
  NAND2_X1 U21605 ( .A1(n18564), .A2(n18298), .ZN(n18292) );
  AOI21_X1 U21606 ( .B1(n18551), .B2(n21849), .A(n18292), .ZN(n18274) );
  INV_X1 U21607 ( .A(n18263), .ZN(n18266) );
  INV_X1 U21608 ( .A(n18264), .ZN(n18265) );
  AOI211_X1 U21609 ( .C1(n19012), .C2(n18266), .A(n18265), .B(n18536), .ZN(
        n18269) );
  OAI22_X1 U21610 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n18267), .B1(n18271), 
        .B2(n18568), .ZN(n18268) );
  AOI211_X1 U21611 ( .C1(n18540), .C2(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n18269), .B(n18268), .ZN(n18273) );
  OAI211_X1 U21612 ( .C1(n18275), .C2(n18271), .A(n18580), .B(n18270), .ZN(
        n18272) );
  OAI211_X1 U21613 ( .C1(n18274), .C2(n20113), .A(n18273), .B(n18272), .ZN(
        P3_U2646) );
  NAND2_X1 U21614 ( .A1(n18551), .A2(n21849), .ZN(n18283) );
  AOI22_X1 U21615 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n18540), .B1(
        n18581), .B2(P3_EBX_REG_24__SCAN_IN), .ZN(n18282) );
  AOI211_X1 U21616 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n18293), .A(n18275), .B(
        n18567), .ZN(n18280) );
  AOI211_X1 U21617 ( .C1(n18278), .C2(n18277), .A(n18276), .B(n18536), .ZN(
        n18279) );
  AOI211_X1 U21618 ( .C1(P3_REIP_REG_24__SCAN_IN), .C2(n18292), .A(n18280), 
        .B(n18279), .ZN(n18281) );
  OAI211_X1 U21619 ( .C1(n18284), .C2(n18283), .A(n18282), .B(n18281), .ZN(
        P3_U2647) );
  INV_X1 U21620 ( .A(n18285), .ZN(n18297) );
  INV_X1 U21621 ( .A(n18286), .ZN(n18289) );
  INV_X1 U21622 ( .A(n18287), .ZN(n18288) );
  AOI211_X1 U21623 ( .C1(n19036), .C2(n18289), .A(n18288), .B(n18536), .ZN(
        n18291) );
  OAI22_X1 U21624 ( .A1(n10497), .A2(n18558), .B1(n18568), .B2(n18294), .ZN(
        n18290) );
  AOI211_X1 U21625 ( .C1(P3_REIP_REG_23__SCAN_IN), .C2(n18292), .A(n18291), 
        .B(n18290), .ZN(n18296) );
  OAI211_X1 U21626 ( .C1(n18302), .C2(n18294), .A(n18580), .B(n18293), .ZN(
        n18295) );
  OAI211_X1 U21627 ( .C1(n18298), .C2(n18297), .A(n18296), .B(n18295), .ZN(
        P3_U2648) );
  AOI21_X1 U21628 ( .B1(n18551), .B2(n18299), .A(n18576), .ZN(n18328) );
  AOI211_X1 U21629 ( .C1(n18301), .C2(n9847), .A(n18300), .B(n18536), .ZN(
        n18306) );
  AOI211_X1 U21630 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n18316), .A(n18302), .B(
        n18567), .ZN(n18305) );
  AOI22_X1 U21631 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n18540), .B1(
        n18581), .B2(P3_EBX_REG_22__SCAN_IN), .ZN(n18303) );
  INV_X1 U21632 ( .A(n18303), .ZN(n18304) );
  NOR3_X1 U21633 ( .A1(n18306), .A2(n18305), .A3(n18304), .ZN(n18309) );
  NAND3_X1 U21634 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(P3_REIP_REG_20__SCAN_IN), 
        .A3(P3_REIP_REG_18__SCAN_IN), .ZN(n18307) );
  NAND2_X1 U21635 ( .A1(n18551), .A2(n18329), .ZN(n18346) );
  NOR2_X1 U21636 ( .A1(n18307), .A2(n18346), .ZN(n18314) );
  OAI221_X1 U21637 ( .B1(P3_REIP_REG_21__SCAN_IN), .B2(P3_REIP_REG_22__SCAN_IN), .C1(n21832), .C2(n20108), .A(n18314), .ZN(n18308) );
  OAI211_X1 U21638 ( .C1(n20108), .C2(n18328), .A(n18309), .B(n18308), .ZN(
        P3_U2649) );
  AOI22_X1 U21639 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n18540), .B1(
        n18581), .B2(P3_EBX_REG_21__SCAN_IN), .ZN(n18319) );
  INV_X1 U21640 ( .A(n18328), .ZN(n18315) );
  INV_X1 U21641 ( .A(n18310), .ZN(n18311) );
  AOI211_X1 U21642 ( .C1(n19066), .C2(n18312), .A(n18311), .B(n18536), .ZN(
        n18313) );
  AOI221_X1 U21643 ( .B1(n18315), .B2(P3_REIP_REG_21__SCAN_IN), .C1(n18314), 
        .C2(n21832), .A(n18313), .ZN(n18318) );
  OAI211_X1 U21644 ( .C1(n18323), .C2(n18676), .A(n18580), .B(n18316), .ZN(
        n18317) );
  NAND3_X1 U21645 ( .A1(n18319), .A2(n18318), .A3(n18317), .ZN(P3_U2650) );
  INV_X1 U21646 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n20105) );
  AOI211_X1 U21647 ( .C1(n18321), .C2(n18330), .A(n18320), .B(n18536), .ZN(
        n18322) );
  AOI21_X1 U21648 ( .B1(n18540), .B2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n18322), .ZN(n18327) );
  INV_X1 U21649 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n20104) );
  INV_X1 U21650 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n20101) );
  NOR4_X1 U21651 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n20104), .A3(n20101), 
        .A4(n18346), .ZN(n18325) );
  AOI211_X1 U21652 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n18337), .A(n18323), .B(
        n18567), .ZN(n18324) );
  AOI211_X1 U21653 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n18581), .A(n18325), .B(
        n18324), .ZN(n18326) );
  OAI211_X1 U21654 ( .C1(n20105), .C2(n18328), .A(n18327), .B(n18326), .ZN(
        P3_U2651) );
  NOR2_X1 U21655 ( .A1(n20101), .A2(n18346), .ZN(n18336) );
  OR2_X1 U21656 ( .A1(n18329), .A2(n18574), .ZN(n18357) );
  NAND2_X1 U21657 ( .A1(n18564), .A2(n18357), .ZN(n18362) );
  INV_X1 U21658 ( .A(n18362), .ZN(n18352) );
  OAI21_X1 U21659 ( .B1(P3_REIP_REG_18__SCAN_IN), .B2(n18346), .A(n18352), 
        .ZN(n18335) );
  INV_X1 U21660 ( .A(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n18333) );
  NAND2_X1 U21661 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n19099), .ZN(
        n18341) );
  AOI21_X1 U21662 ( .B1(n18333), .B2(n18341), .A(n19051), .ZN(n18331) );
  INV_X1 U21663 ( .A(n18331), .ZN(n19104) );
  OAI21_X1 U21664 ( .B1(n18341), .B2(n18342), .A(n10503), .ZN(n18344) );
  OAI221_X1 U21665 ( .B1(n18331), .B2(n18330), .C1(n19104), .C2(n18344), .A(
        n20050), .ZN(n18332) );
  OAI211_X1 U21666 ( .C1(n18333), .C2(n18558), .A(n19442), .B(n18332), .ZN(
        n18334) );
  AOI221_X1 U21667 ( .B1(n18336), .B2(n20104), .C1(n18335), .C2(
        P3_REIP_REG_19__SCAN_IN), .A(n18334), .ZN(n18339) );
  OAI211_X1 U21668 ( .C1(n18347), .C2(n18340), .A(n18580), .B(n18337), .ZN(
        n18338) );
  OAI211_X1 U21669 ( .C1(n18340), .C2(n18568), .A(n18339), .B(n18338), .ZN(
        P3_U2652) );
  OAI21_X1 U21670 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n19099), .A(
        n18341), .ZN(n19111) );
  NAND2_X1 U21671 ( .A1(n20050), .A2(n18518), .ZN(n18561) );
  INV_X1 U21672 ( .A(n18342), .ZN(n18354) );
  INV_X1 U21673 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n19114) );
  OAI221_X1 U21674 ( .B1(n19111), .B2(n18354), .C1(n19111), .C2(n19114), .A(
        n20050), .ZN(n18343) );
  AOI22_X1 U21675 ( .A1(n19111), .A2(n18344), .B1(n18561), .B2(n18343), .ZN(
        n18345) );
  AOI211_X1 U21676 ( .C1(n18581), .C2(P3_EBX_REG_18__SCAN_IN), .A(n19494), .B(
        n18345), .ZN(n18351) );
  NOR2_X1 U21677 ( .A1(P3_REIP_REG_18__SCAN_IN), .A2(n18346), .ZN(n18349) );
  AOI211_X1 U21678 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n18363), .A(n18347), .B(
        n18567), .ZN(n18348) );
  AOI211_X1 U21679 ( .C1(n18540), .C2(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n18349), .B(n18348), .ZN(n18350) );
  OAI211_X1 U21680 ( .C1(n18352), .C2(n20101), .A(n18351), .B(n18350), .ZN(
        P3_U2653) );
  OAI22_X1 U21681 ( .A1(n18353), .A2(n18558), .B1(n18568), .B2(n18364), .ZN(
        n18361) );
  AOI21_X1 U21682 ( .B1(n18354), .B2(n18369), .A(n18518), .ZN(n18355) );
  XNOR2_X1 U21683 ( .A(n18356), .B(n18355), .ZN(n18359) );
  OAI22_X1 U21684 ( .A1(n18536), .A2(n18359), .B1(n18358), .B2(n18357), .ZN(
        n18360) );
  AOI211_X1 U21685 ( .C1(P3_REIP_REG_17__SCAN_IN), .C2(n18362), .A(n18361), 
        .B(n18360), .ZN(n18366) );
  OAI211_X1 U21686 ( .C1(n18367), .C2(n18364), .A(n18580), .B(n18363), .ZN(
        n18365) );
  NAND3_X1 U21687 ( .A1(n18366), .A2(n19442), .A3(n18365), .ZN(P3_U2654) );
  NAND3_X1 U21688 ( .A1(n18551), .A2(P3_REIP_REG_15__SCAN_IN), .A3(n18377), 
        .ZN(n18376) );
  INV_X1 U21689 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n20097) );
  INV_X1 U21690 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n20095) );
  NAND2_X1 U21691 ( .A1(n18377), .A2(n18564), .ZN(n18397) );
  OAI21_X1 U21692 ( .B1(n20095), .B2(n18397), .A(n18579), .ZN(n18387) );
  AOI211_X1 U21693 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n18383), .A(n18367), .B(
        n18567), .ZN(n18374) );
  INV_X1 U21694 ( .A(P3_EBX_REG_16__SCAN_IN), .ZN(n18372) );
  NAND2_X1 U21695 ( .A1(n18370), .A2(n18369), .ZN(n18368) );
  OAI211_X1 U21696 ( .C1(n18370), .C2(n18369), .A(n20050), .B(n18368), .ZN(
        n18371) );
  OAI211_X1 U21697 ( .C1(n18568), .C2(n18372), .A(n19442), .B(n18371), .ZN(
        n18373) );
  AOI211_X1 U21698 ( .C1(n18540), .C2(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n18374), .B(n18373), .ZN(n18375) );
  OAI221_X1 U21699 ( .B1(P3_REIP_REG_16__SCAN_IN), .B2(n18376), .C1(n20097), 
        .C2(n18387), .A(n18375), .ZN(P3_U2655) );
  AOI21_X1 U21700 ( .B1(n18551), .B2(n18377), .A(P3_REIP_REG_15__SCAN_IN), 
        .ZN(n18388) );
  NOR2_X1 U21701 ( .A1(n18378), .A2(n18518), .ZN(n18392) );
  AOI22_X1 U21702 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n18380), .B1(
        n18379), .B2(n19128), .ZN(n19125) );
  XOR2_X1 U21703 ( .A(n18392), .B(n19125), .Z(n18381) );
  OAI22_X1 U21704 ( .A1(n18568), .A2(n18384), .B1(n18536), .B2(n18381), .ZN(
        n18382) );
  AOI211_X1 U21705 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(n18540), .A(
        n19494), .B(n18382), .ZN(n18386) );
  OAI211_X1 U21706 ( .C1(n18389), .C2(n18384), .A(n18580), .B(n18383), .ZN(
        n18385) );
  OAI211_X1 U21707 ( .C1(n18388), .C2(n18387), .A(n18386), .B(n18385), .ZN(
        P3_U2656) );
  AOI211_X1 U21708 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n18409), .A(n18389), .B(
        n18567), .ZN(n18396) );
  INV_X1 U21709 ( .A(n17819), .ZN(n18390) );
  OAI211_X1 U21710 ( .C1(n18390), .C2(n18522), .A(n10503), .B(n18393), .ZN(
        n18391) );
  OAI211_X1 U21711 ( .C1(n18393), .C2(n18392), .A(n20050), .B(n18391), .ZN(
        n18394) );
  NAND2_X1 U21712 ( .A1(n19442), .A2(n18394), .ZN(n18395) );
  AOI211_X1 U21713 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n18581), .A(n18396), .B(
        n18395), .ZN(n18400) );
  NOR3_X1 U21714 ( .A1(n18574), .A2(n20091), .A3(n18406), .ZN(n18398) );
  OAI211_X1 U21715 ( .C1(P3_REIP_REG_14__SCAN_IN), .C2(n18398), .A(n18397), 
        .B(n18579), .ZN(n18399) );
  OAI211_X1 U21716 ( .C1(n18558), .C2(n18401), .A(n18400), .B(n18399), .ZN(
        P3_U2657) );
  AOI22_X1 U21717 ( .A1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n18540), .B1(
        n18581), .B2(P3_EBX_REG_13__SCAN_IN), .ZN(n18414) );
  INV_X1 U21718 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n19162) );
  NOR2_X1 U21719 ( .A1(n19162), .A2(n19142), .ZN(n18403) );
  OAI21_X1 U21720 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n18403), .A(
        n18402), .ZN(n19152) );
  NOR2_X1 U21721 ( .A1(n19147), .A2(n18522), .ZN(n18417) );
  AOI21_X1 U21722 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n18417), .A(
        n18518), .ZN(n18404) );
  XNOR2_X1 U21723 ( .A(n19152), .B(n18404), .ZN(n18405) );
  AOI21_X1 U21724 ( .B1(n18405), .B2(n20050), .A(n19494), .ZN(n18413) );
  OR2_X1 U21725 ( .A1(n18574), .A2(n18406), .ZN(n18408) );
  OAI21_X1 U21726 ( .B1(n18422), .B2(n18574), .A(n18564), .ZN(n18433) );
  NOR2_X1 U21727 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n18574), .ZN(n18421) );
  NOR2_X1 U21728 ( .A1(n18433), .A2(n18421), .ZN(n18407) );
  MUX2_X1 U21729 ( .A(n18408), .B(n18407), .S(P3_REIP_REG_13__SCAN_IN), .Z(
        n18412) );
  OAI211_X1 U21730 ( .C1(n18415), .C2(n18410), .A(n18580), .B(n18409), .ZN(
        n18411) );
  NAND4_X1 U21731 ( .A1(n18414), .A2(n18413), .A3(n18412), .A4(n18411), .ZN(
        P3_U2658) );
  AOI211_X1 U21732 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n18434), .A(n18415), .B(
        n18567), .ZN(n18416) );
  AOI21_X1 U21733 ( .B1(n18540), .B2(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n18416), .ZN(n18425) );
  NOR2_X1 U21734 ( .A1(n18417), .A2(n18518), .ZN(n18419) );
  AOI22_X1 U21735 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n19142), .B1(
        n18418), .B2(n19162), .ZN(n19158) );
  XNOR2_X1 U21736 ( .A(n18419), .B(n19158), .ZN(n18420) );
  AOI22_X1 U21737 ( .A1(n18581), .A2(P3_EBX_REG_12__SCAN_IN), .B1(n20050), 
        .B2(n18420), .ZN(n18424) );
  AOI22_X1 U21738 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n18433), .B1(n18422), 
        .B2(n18421), .ZN(n18423) );
  NAND4_X1 U21739 ( .A1(n18425), .A2(n18424), .A3(n18423), .A4(n19442), .ZN(
        P3_U2659) );
  NAND2_X1 U21740 ( .A1(n17848), .A2(n18547), .ZN(n18477) );
  OAI21_X1 U21741 ( .B1(n18426), .B2(n18477), .A(n10503), .ZN(n18428) );
  AOI21_X1 U21742 ( .B1(n18429), .B2(n18428), .A(n19494), .ZN(n18427) );
  OAI21_X1 U21743 ( .B1(n18429), .B2(n18428), .A(n18427), .ZN(n18430) );
  AOI22_X1 U21744 ( .A1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n18540), .B1(
        n18523), .B2(n18430), .ZN(n18437) );
  OAI21_X1 U21745 ( .B1(n18574), .B2(n18431), .A(n20087), .ZN(n18432) );
  AOI22_X1 U21746 ( .A1(n18581), .A2(P3_EBX_REG_11__SCAN_IN), .B1(n18433), 
        .B2(n18432), .ZN(n18436) );
  OAI211_X1 U21747 ( .C1(n18440), .C2(n18717), .A(n18580), .B(n18434), .ZN(
        n18435) );
  NAND3_X1 U21748 ( .A1(n18437), .A2(n18436), .A3(n18435), .ZN(P3_U2660) );
  NAND2_X1 U21749 ( .A1(n18551), .A2(n18438), .ZN(n18450) );
  INV_X1 U21750 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n20086) );
  OAI21_X1 U21751 ( .B1(n18574), .B2(n18438), .A(n18564), .ZN(n18439) );
  INV_X1 U21752 ( .A(n18439), .ZN(n18451) );
  AOI211_X1 U21753 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n18458), .A(n18440), .B(
        n18567), .ZN(n18448) );
  INV_X1 U21754 ( .A(n18443), .ZN(n18442) );
  OAI21_X1 U21755 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n18442), .A(
        n18441), .ZN(n18444) );
  INV_X1 U21756 ( .A(n18444), .ZN(n19171) );
  OAI21_X1 U21757 ( .B1(n18443), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n10503), .ZN(n18445) );
  INV_X1 U21758 ( .A(n18445), .ZN(n18453) );
  AOI221_X1 U21759 ( .B1(n19171), .B2(n18445), .C1(n18444), .C2(n18453), .A(
        n19494), .ZN(n18446) );
  OAI22_X1 U21760 ( .A1(n18481), .A2(n18446), .B1(n18568), .B2(n18752), .ZN(
        n18447) );
  AOI211_X1 U21761 ( .C1(n18540), .C2(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n18448), .B(n18447), .ZN(n18449) );
  OAI221_X1 U21762 ( .B1(P3_REIP_REG_10__SCAN_IN), .B2(n18450), .C1(n20086), 
        .C2(n18451), .A(n18449), .ZN(P3_U2661) );
  INV_X1 U21763 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n21712) );
  NAND4_X1 U21764 ( .A1(n18551), .A2(n18511), .A3(P3_REIP_REG_5__SCAN_IN), 
        .A4(P3_REIP_REG_4__SCAN_IN), .ZN(n18499) );
  NOR2_X1 U21765 ( .A1(n21712), .A2(n18499), .ZN(n18483) );
  NAND2_X1 U21766 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(n18483), .ZN(n18475) );
  AOI221_X1 U21767 ( .B1(n20082), .B2(n20084), .C1(n18475), .C2(n20084), .A(
        n18451), .ZN(n18457) );
  INV_X1 U21768 ( .A(n17848), .ZN(n18467) );
  NOR4_X1 U21769 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n19192), .A3(
        n18467), .A4(n18522), .ZN(n18452) );
  AOI211_X1 U21770 ( .C1(n18453), .C2(n18454), .A(n19494), .B(n18452), .ZN(
        n18455) );
  OAI22_X1 U21771 ( .A1(n18481), .A2(n18455), .B1(n18561), .B2(n18454), .ZN(
        n18456) );
  AOI211_X1 U21772 ( .C1(P3_EBX_REG_9__SCAN_IN), .C2(n18581), .A(n18457), .B(
        n18456), .ZN(n18461) );
  OAI211_X1 U21773 ( .C1(n18464), .C2(n18459), .A(n18580), .B(n18458), .ZN(
        n18460) );
  OAI211_X1 U21774 ( .C1(n18558), .C2(n18462), .A(n18461), .B(n18460), .ZN(
        P3_U2662) );
  AOI221_X1 U21775 ( .B1(n18463), .B2(n18551), .C1(n18489), .C2(n18551), .A(
        n18576), .ZN(n18476) );
  INV_X1 U21776 ( .A(n18464), .ZN(n18473) );
  OAI222_X1 U21777 ( .A1(n18567), .A2(n18485), .B1(n18567), .B2(
        P3_EBX_REG_8__SCAN_IN), .C1(n18568), .C2(n18465), .ZN(n18472) );
  AOI21_X1 U21778 ( .B1(n18470), .B2(n18478), .A(n18466), .ZN(n19183) );
  INV_X1 U21779 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n19198) );
  NOR2_X1 U21780 ( .A1(n18467), .A2(n19198), .ZN(n19193) );
  AOI21_X1 U21781 ( .B1(n18547), .B2(n19193), .A(n18518), .ZN(n18468) );
  XNOR2_X1 U21782 ( .A(n19183), .B(n18468), .ZN(n18469) );
  OAI22_X1 U21783 ( .A1(n18470), .A2(n18558), .B1(n18536), .B2(n18469), .ZN(
        n18471) );
  AOI211_X1 U21784 ( .C1(n18473), .C2(n18472), .A(n19494), .B(n18471), .ZN(
        n18474) );
  OAI221_X1 U21785 ( .B1(P3_REIP_REG_8__SCAN_IN), .B2(n18475), .C1(n20082), 
        .C2(n18476), .A(n18474), .ZN(P3_U2663) );
  INV_X1 U21786 ( .A(n18476), .ZN(n18484) );
  INV_X1 U21787 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n20081) );
  AND2_X1 U21788 ( .A1(n18477), .A2(n10503), .ZN(n18492) );
  OAI21_X1 U21789 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n18491), .A(
        n18478), .ZN(n19209) );
  OAI21_X1 U21790 ( .B1(n18492), .B2(n19209), .A(n19442), .ZN(n18479) );
  AOI21_X1 U21791 ( .B1(n18492), .B2(n19209), .A(n18479), .ZN(n18480) );
  OAI22_X1 U21792 ( .A1(n18481), .A2(n18480), .B1(n19198), .B2(n18558), .ZN(
        n18482) );
  AOI221_X1 U21793 ( .B1(n18484), .B2(P3_REIP_REG_7__SCAN_IN), .C1(n18483), 
        .C2(n20081), .A(n18482), .ZN(n18487) );
  OAI211_X1 U21794 ( .C1(n18490), .C2(n18488), .A(n18580), .B(n18485), .ZN(
        n18486) );
  OAI211_X1 U21795 ( .C1(n18488), .C2(n18568), .A(n18487), .B(n18486), .ZN(
        P3_U2664) );
  AOI21_X1 U21796 ( .B1(n18551), .B2(n18489), .A(n18576), .ZN(n18502) );
  AOI211_X1 U21797 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n18507), .A(n18490), .B(
        n18567), .ZN(n18497) );
  OR2_X1 U21798 ( .A1(n18562), .A2(n19217), .ZN(n18500) );
  AOI21_X1 U21799 ( .B1(n19218), .B2(n18500), .A(n18491), .ZN(n19220) );
  NAND2_X1 U21800 ( .A1(n20050), .A2(n18492), .ZN(n18495) );
  INV_X1 U21801 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n18575) );
  NAND2_X1 U21802 ( .A1(n20050), .A2(n18575), .ZN(n18560) );
  OAI21_X1 U21803 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n18560), .A(
        n18561), .ZN(n18493) );
  AOI22_X1 U21804 ( .A1(n18581), .A2(P3_EBX_REG_6__SCAN_IN), .B1(n19220), .B2(
        n18493), .ZN(n18494) );
  OAI211_X1 U21805 ( .C1(n19220), .C2(n18495), .A(n18494), .B(n19442), .ZN(
        n18496) );
  AOI211_X1 U21806 ( .C1(n18540), .C2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n18497), .B(n18496), .ZN(n18498) );
  OAI221_X1 U21807 ( .B1(P3_REIP_REG_6__SCAN_IN), .B2(n18499), .C1(n21712), 
        .C2(n18502), .A(n18498), .ZN(P3_U2665) );
  AND2_X1 U21808 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n19227), .ZN(
        n18517) );
  AOI21_X1 U21809 ( .B1(n18517), .B2(n18575), .A(n18518), .ZN(n18520) );
  OAI21_X1 U21810 ( .B1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n18517), .A(
        n18500), .ZN(n19230) );
  XOR2_X1 U21811 ( .A(n18520), .B(n19230), .Z(n18501) );
  OAI21_X1 U21812 ( .B1(n18536), .B2(n18501), .A(n19442), .ZN(n18506) );
  INV_X1 U21813 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n20078) );
  NAND2_X1 U21814 ( .A1(n18551), .A2(n18511), .ZN(n18530) );
  NOR2_X1 U21815 ( .A1(n20078), .A2(n18530), .ZN(n18504) );
  INV_X1 U21816 ( .A(n18502), .ZN(n18503) );
  MUX2_X1 U21817 ( .A(n18504), .B(n18503), .S(P3_REIP_REG_5__SCAN_IN), .Z(
        n18505) );
  AOI211_X1 U21818 ( .C1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .C2(n18540), .A(
        n18506), .B(n18505), .ZN(n18509) );
  OAI211_X1 U21819 ( .C1(n18513), .C2(n18510), .A(n18580), .B(n18507), .ZN(
        n18508) );
  OAI211_X1 U21820 ( .C1(n18510), .C2(n18568), .A(n18509), .B(n18508), .ZN(
        P3_U2666) );
  OAI21_X1 U21821 ( .B1(n18574), .B2(n18511), .A(n18564), .ZN(n18512) );
  INV_X1 U21822 ( .A(n18512), .ZN(n18531) );
  AOI211_X1 U21823 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n18541), .A(n18513), .B(
        n18567), .ZN(n18528) );
  NOR2_X1 U21824 ( .A1(n18699), .A2(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n18514) );
  NAND2_X1 U21825 ( .A1(n20169), .A2(n19565), .ZN(n20172) );
  OAI22_X1 U21826 ( .A1(n18568), .A2(n18764), .B1(n18514), .B2(n20172), .ZN(
        n18515) );
  AOI21_X1 U21827 ( .B1(n18540), .B2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n18515), .ZN(n18526) );
  NAND2_X1 U21828 ( .A1(n18516), .A2(n21869), .ZN(n19247) );
  NAND2_X1 U21829 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18516), .ZN(
        n18532) );
  AOI21_X1 U21830 ( .B1(n21869), .B2(n18532), .A(n18517), .ZN(n19244) );
  INV_X1 U21831 ( .A(n19244), .ZN(n18519) );
  AOI221_X1 U21832 ( .B1(n18520), .B2(n18519), .C1(n18518), .C2(n19244), .A(
        n19494), .ZN(n18521) );
  OAI21_X1 U21833 ( .B1(n18522), .B2(n19247), .A(n18521), .ZN(n18524) );
  NAND2_X1 U21834 ( .A1(n18524), .A2(n18523), .ZN(n18525) );
  NAND2_X1 U21835 ( .A1(n18526), .A2(n18525), .ZN(n18527) );
  NOR2_X1 U21836 ( .A1(n18528), .A2(n18527), .ZN(n18529) );
  OAI221_X1 U21837 ( .B1(P3_REIP_REG_4__SCAN_IN), .B2(n18530), .C1(n20078), 
        .C2(n18531), .A(n18529), .ZN(P3_U2667) );
  AOI221_X1 U21838 ( .B1(n18574), .B2(n20077), .C1(n18550), .C2(n20077), .A(
        n18531), .ZN(n18539) );
  NAND2_X1 U21839 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n18546) );
  INV_X1 U21840 ( .A(n18546), .ZN(n18533) );
  OAI21_X1 U21841 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n18533), .A(
        n18532), .ZN(n19249) );
  OAI21_X1 U21842 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n18546), .A(
        n10503), .ZN(n18534) );
  XNOR2_X1 U21843 ( .A(n19249), .B(n18534), .ZN(n18537) );
  OAI22_X1 U21844 ( .A1(n18537), .A2(n18536), .B1(n20172), .B2(n18535), .ZN(
        n18538) );
  AOI211_X1 U21845 ( .C1(n18540), .C2(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n18539), .B(n18538), .ZN(n18543) );
  OAI211_X1 U21846 ( .C1(n18545), .C2(n18544), .A(n18580), .B(n18541), .ZN(
        n18542) );
  OAI211_X1 U21847 ( .C1(n18544), .C2(n18568), .A(n18543), .B(n18542), .ZN(
        P3_U2668) );
  INV_X1 U21848 ( .A(P3_EBX_REG_0__SCAN_IN), .ZN(n18784) );
  INV_X1 U21849 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n18779) );
  NAND2_X1 U21850 ( .A1(n18784), .A2(n18779), .ZN(n18566) );
  AOI211_X1 U21851 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n18566), .A(n18545), .B(
        n18567), .ZN(n18556) );
  OAI21_X1 U21852 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n18546), .ZN(n19263) );
  OAI22_X1 U21853 ( .A1(n18547), .A2(n19263), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n18546), .ZN(n18548) );
  OAI22_X1 U21854 ( .A1(n18559), .A2(n18548), .B1(n18561), .B2(n19263), .ZN(
        n18549) );
  AOI21_X1 U21855 ( .B1(P3_REIP_REG_2__SCAN_IN), .B2(n18576), .A(n18549), .ZN(
        n18553) );
  OAI211_X1 U21856 ( .C1(P3_REIP_REG_1__SCAN_IN), .C2(P3_REIP_REG_2__SCAN_IN), 
        .A(n18551), .B(n18550), .ZN(n18552) );
  OAI211_X1 U21857 ( .C1(n20172), .C2(n18554), .A(n18553), .B(n18552), .ZN(
        n18555) );
  AOI211_X1 U21858 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n18581), .A(n18556), .B(
        n18555), .ZN(n18557) );
  OAI21_X1 U21859 ( .B1(n19272), .B2(n18558), .A(n18557), .ZN(P3_U2669) );
  OAI211_X1 U21860 ( .C1(n18575), .C2(n18559), .A(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B(n18558), .ZN(n18572) );
  NAND3_X1 U21861 ( .A1(n18562), .A2(n18561), .A3(n18560), .ZN(n18571) );
  OAI22_X1 U21862 ( .A1(n18564), .A2(n20136), .B1(n20172), .B2(n18563), .ZN(
        n18570) );
  NOR2_X1 U21863 ( .A1(n18784), .A2(n18779), .ZN(n18773) );
  INV_X1 U21864 ( .A(n18773), .ZN(n18565) );
  NAND2_X1 U21865 ( .A1(n18566), .A2(n18565), .ZN(n18781) );
  OAI22_X1 U21866 ( .A1(n18568), .A2(n18779), .B1(n18567), .B2(n18781), .ZN(
        n18569) );
  AOI211_X1 U21867 ( .C1(n18572), .C2(n18571), .A(n18570), .B(n18569), .ZN(
        n18573) );
  OAI21_X1 U21868 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n18574), .A(n18573), .ZN(
        P3_U2670) );
  NOR2_X1 U21869 ( .A1(n18576), .A2(n18575), .ZN(n18578) );
  AOI22_X1 U21870 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(n18579), .B1(n18578), 
        .B2(n18577), .ZN(n18583) );
  OAI21_X1 U21871 ( .B1(n18581), .B2(n18580), .A(P3_EBX_REG_0__SCAN_IN), .ZN(
        n18582) );
  OAI211_X1 U21872 ( .C1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n20172), .A(
        n18583), .B(n18582), .ZN(P3_U2671) );
  AND4_X1 U21873 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(P3_EBX_REG_23__SCAN_IN), 
        .A3(P3_EBX_REG_22__SCAN_IN), .A4(P3_EBX_REG_21__SCAN_IN), .ZN(n18587)
         );
  INV_X1 U21874 ( .A(P3_EBX_REG_26__SCAN_IN), .ZN(n18634) );
  NOR4_X1 U21875 ( .A1(n18634), .A2(n18585), .A3(n18584), .A4(n18626), .ZN(
        n18586) );
  NAND4_X1 U21876 ( .A1(P3_EBX_REG_25__SCAN_IN), .A2(P3_EBX_REG_24__SCAN_IN), 
        .A3(n18587), .A4(n18586), .ZN(n18620) );
  NOR2_X1 U21877 ( .A1(n18621), .A2(n18620), .ZN(n18619) );
  NAND2_X1 U21878 ( .A1(n18777), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n18589) );
  NAND2_X1 U21879 ( .A1(n18619), .A2(n19588), .ZN(n18588) );
  OAI22_X1 U21880 ( .A1(n18619), .A2(n18589), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n18588), .ZN(P3_U2672) );
  INV_X1 U21881 ( .A(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n18595) );
  INV_X1 U21882 ( .A(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n18590) );
  INV_X1 U21883 ( .A(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n18659) );
  OAI22_X1 U21884 ( .A1(n18724), .A2(n18590), .B1(n18722), .B2(n18659), .ZN(
        n18592) );
  INV_X1 U21885 ( .A(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n18680) );
  OAI22_X1 U21886 ( .A1(n18728), .A2(n18680), .B1(n18726), .B2(n11586), .ZN(
        n18591) );
  AOI211_X1 U21887 ( .C1(n18731), .C2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A(
        n18592), .B(n18591), .ZN(n18594) );
  AOI22_X1 U21888 ( .A1(n13185), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n18732), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n18593) );
  OAI211_X1 U21889 ( .C1(n9681), .C2(n18595), .A(n18594), .B(n18593), .ZN(
        n18602) );
  AOI22_X1 U21890 ( .A1(n18736), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n13878), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n18600) );
  AOI22_X1 U21891 ( .A1(n13279), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n18596), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n18599) );
  AOI22_X1 U21892 ( .A1(n18738), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n18737), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n18598) );
  AOI22_X1 U21893 ( .A1(n18740), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n18739), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n18597) );
  NAND4_X1 U21894 ( .A1(n18600), .A2(n18599), .A3(n18598), .A4(n18597), .ZN(
        n18601) );
  NOR2_X1 U21895 ( .A1(n18602), .A2(n18601), .ZN(n18624) );
  NOR2_X1 U21896 ( .A1(n18625), .A2(n18624), .ZN(n18618) );
  INV_X1 U21897 ( .A(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n18604) );
  OAI22_X1 U21898 ( .A1(n18604), .A2(n18724), .B1(n18722), .B2(n18603), .ZN(
        n18608) );
  INV_X1 U21899 ( .A(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n18606) );
  INV_X1 U21900 ( .A(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n18605) );
  OAI22_X1 U21901 ( .A1(n18728), .A2(n18606), .B1(n18726), .B2(n18605), .ZN(
        n18607) );
  AOI211_X1 U21902 ( .C1(n18731), .C2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A(
        n18608), .B(n18607), .ZN(n18610) );
  AOI22_X1 U21903 ( .A1(n9703), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n18732), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n18609) );
  OAI211_X1 U21904 ( .C1(n19640), .C2(n18735), .A(n18610), .B(n18609), .ZN(
        n18616) );
  AOI22_X1 U21905 ( .A1(n18736), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n13878), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n18614) );
  AOI22_X1 U21906 ( .A1(n13279), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n18596), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n18613) );
  AOI22_X1 U21907 ( .A1(n18738), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n18737), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n18612) );
  AOI22_X1 U21908 ( .A1(n18740), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n18739), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n18611) );
  NAND4_X1 U21909 ( .A1(n18614), .A2(n18613), .A3(n18612), .A4(n18611), .ZN(
        n18615) );
  NOR2_X1 U21910 ( .A1(n18616), .A2(n18615), .ZN(n18617) );
  XNOR2_X1 U21911 ( .A(n18618), .B(n18617), .ZN(n18793) );
  AOI211_X1 U21912 ( .C1(n18621), .C2(n18620), .A(n18619), .B(n18749), .ZN(
        n18622) );
  AOI21_X1 U21913 ( .B1(n18749), .B2(n18793), .A(n18622), .ZN(n18623) );
  INV_X1 U21914 ( .A(n18623), .ZN(P3_U2673) );
  XNOR2_X1 U21915 ( .A(n18625), .B(n18624), .ZN(n18801) );
  OAI21_X1 U21916 ( .B1(n18638), .B2(n18626), .A(n21826), .ZN(n18627) );
  OAI21_X1 U21917 ( .B1(n21826), .B2(n18628), .A(n18627), .ZN(n18629) );
  OAI21_X1 U21918 ( .B1(n18801), .B2(n18770), .A(n18629), .ZN(P3_U2674) );
  OAI21_X1 U21919 ( .B1(n18635), .B2(n18631), .A(n18630), .ZN(n18811) );
  NAND3_X1 U21920 ( .A1(n18638), .A2(P3_EBX_REG_27__SCAN_IN), .A3(n18770), 
        .ZN(n18632) );
  OAI221_X1 U21921 ( .B1(n18638), .B2(P3_EBX_REG_27__SCAN_IN), .C1(n18777), 
        .C2(n18811), .A(n18632), .ZN(P3_U2676) );
  OAI21_X1 U21922 ( .B1(n18634), .B2(n18749), .A(n18633), .ZN(n18637) );
  AOI21_X1 U21923 ( .B1(n18636), .B2(n18640), .A(n18635), .ZN(n18812) );
  AOI22_X1 U21924 ( .A1(n18638), .A2(n18637), .B1(n18812), .B2(n18749), .ZN(
        n18639) );
  INV_X1 U21925 ( .A(n18639), .ZN(P3_U2677) );
  AOI21_X1 U21926 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n18777), .A(n18649), .ZN(
        n18642) );
  OAI21_X1 U21927 ( .B1(n18646), .B2(n18641), .A(n18640), .ZN(n18821) );
  OAI22_X1 U21928 ( .A1(n18643), .A2(n18642), .B1(n18821), .B2(n18770), .ZN(
        P3_U2678) );
  AOI21_X1 U21929 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n18777), .A(n18655), .ZN(
        n18648) );
  AND2_X1 U21930 ( .A1(n18651), .A2(n18644), .ZN(n18645) );
  NOR2_X1 U21931 ( .A1(n18646), .A2(n18645), .ZN(n18822) );
  INV_X1 U21932 ( .A(n18822), .ZN(n18647) );
  OAI22_X1 U21933 ( .A1(n18649), .A2(n18648), .B1(n18647), .B2(n18770), .ZN(
        P3_U2679) );
  INV_X1 U21934 ( .A(n18650), .ZN(n18672) );
  AOI21_X1 U21935 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n18777), .A(n18672), .ZN(
        n18654) );
  OAI21_X1 U21936 ( .B1(n18653), .B2(n18652), .A(n18651), .ZN(n18833) );
  OAI22_X1 U21937 ( .A1(n18655), .A2(n18654), .B1(n18777), .B2(n18833), .ZN(
        P3_U2680) );
  AOI21_X1 U21938 ( .B1(P3_EBX_REG_22__SCAN_IN), .B2(n18777), .A(n18656), .ZN(
        n18671) );
  NAND2_X1 U21939 ( .A1(n13185), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n18658) );
  NAND2_X1 U21940 ( .A1(n18699), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n18657) );
  OAI211_X1 U21941 ( .C1(n9681), .C2(n18659), .A(n18658), .B(n18657), .ZN(
        n18660) );
  INV_X1 U21942 ( .A(n18660), .ZN(n18664) );
  AOI22_X1 U21943 ( .A1(n18704), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n18703), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n18663) );
  AOI22_X1 U21944 ( .A1(n18706), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n18705), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n18662) );
  NAND2_X1 U21945 ( .A1(n18731), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n18661) );
  NAND4_X1 U21946 ( .A1(n18664), .A2(n18663), .A3(n18662), .A4(n18661), .ZN(
        n18670) );
  AOI22_X1 U21947 ( .A1(n18736), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n13878), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n18668) );
  AOI22_X1 U21948 ( .A1(n13279), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n18596), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n18667) );
  AOI22_X1 U21949 ( .A1(n18740), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n18739), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n18666) );
  AOI22_X1 U21950 ( .A1(n18738), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n18737), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n18665) );
  NAND4_X1 U21951 ( .A1(n18668), .A2(n18667), .A3(n18666), .A4(n18665), .ZN(
        n18669) );
  NOR2_X1 U21952 ( .A1(n18670), .A2(n18669), .ZN(n18834) );
  OAI22_X1 U21953 ( .A1(n18672), .A2(n18671), .B1(n18834), .B2(n18770), .ZN(
        P3_U2681) );
  OR2_X1 U21954 ( .A1(n18770), .A2(n18673), .ZN(n18674) );
  OAI221_X1 U21955 ( .B1(P3_EBX_REG_21__SCAN_IN), .B2(n18677), .C1(n18676), 
        .C2(n18675), .A(n18674), .ZN(P3_U2682) );
  INV_X1 U21956 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n18698) );
  INV_X1 U21957 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n18686) );
  INV_X1 U21958 ( .A(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n18679) );
  OAI22_X1 U21959 ( .A1(n18724), .A2(n18679), .B1(n18722), .B2(n18678), .ZN(
        n18683) );
  INV_X1 U21960 ( .A(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n18681) );
  OAI22_X1 U21961 ( .A1(n18728), .A2(n18681), .B1(n18726), .B2(n18680), .ZN(
        n18682) );
  AOI211_X1 U21962 ( .C1(n18731), .C2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A(
        n18683), .B(n18682), .ZN(n18685) );
  AOI22_X1 U21963 ( .A1(n9703), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n18732), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n18684) );
  OAI211_X1 U21964 ( .C1(n9681), .C2(n18686), .A(n18685), .B(n18684), .ZN(
        n18692) );
  AOI22_X1 U21965 ( .A1(n18736), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n13878), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n18690) );
  AOI22_X1 U21966 ( .A1(n13279), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n18596), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n18689) );
  AOI22_X1 U21967 ( .A1(n18738), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n18737), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n18688) );
  AOI22_X1 U21968 ( .A1(n18740), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n18739), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n18687) );
  NAND4_X1 U21969 ( .A1(n18690), .A2(n18689), .A3(n18688), .A4(n18687), .ZN(
        n18691) );
  OR2_X1 U21970 ( .A1(n18692), .A2(n18691), .ZN(n18864) );
  INV_X1 U21971 ( .A(n18693), .ZN(n18694) );
  NOR3_X1 U21972 ( .A1(n18780), .A2(P3_EBX_REG_14__SCAN_IN), .A3(n18694), .ZN(
        n18695) );
  AOI21_X1 U21973 ( .B1(n18749), .B2(n18864), .A(n18695), .ZN(n18696) );
  OAI21_X1 U21974 ( .B1(n18698), .B2(n18697), .A(n18696), .ZN(P3_U2689) );
  NAND2_X1 U21975 ( .A1(n9704), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n18701) );
  NAND2_X1 U21976 ( .A1(n18699), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n18700) );
  OAI211_X1 U21977 ( .C1(n9681), .C2(n18772), .A(n18701), .B(n18700), .ZN(
        n18702) );
  INV_X1 U21978 ( .A(n18702), .ZN(n18710) );
  AOI22_X1 U21979 ( .A1(n18704), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n9683), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n18709) );
  AOI22_X1 U21980 ( .A1(n18706), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n18705), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n18708) );
  NAND2_X1 U21981 ( .A1(n18731), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n18707) );
  NAND4_X1 U21982 ( .A1(n18710), .A2(n18709), .A3(n18708), .A4(n18707), .ZN(
        n18716) );
  AOI22_X1 U21983 ( .A1(n18736), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n13878), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n18714) );
  AOI22_X1 U21984 ( .A1(n13279), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n18596), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n18713) );
  AOI22_X1 U21985 ( .A1(n18740), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n18739), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n18712) );
  AOI22_X1 U21986 ( .A1(n18738), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n18737), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n18711) );
  NAND4_X1 U21987 ( .A1(n18714), .A2(n18713), .A3(n18712), .A4(n18711), .ZN(
        n18715) );
  NOR2_X1 U21988 ( .A1(n18716), .A2(n18715), .ZN(n18869) );
  OAI21_X1 U21989 ( .B1(n18752), .B2(n18747), .A(n18717), .ZN(n18719) );
  NAND3_X1 U21990 ( .A1(n18719), .A2(n18718), .A3(n18777), .ZN(n18720) );
  OAI21_X1 U21991 ( .B1(n18869), .B2(n18770), .A(n18720), .ZN(P3_U2692) );
  NAND2_X1 U21992 ( .A1(n18777), .A2(n18747), .ZN(n18751) );
  OAI22_X1 U21993 ( .A1(n18724), .A2(n18723), .B1(n18722), .B2(n18721), .ZN(
        n18730) );
  INV_X1 U21994 ( .A(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n18727) );
  OAI22_X1 U21995 ( .A1(n18728), .A2(n18727), .B1(n18726), .B2(n18725), .ZN(
        n18729) );
  AOI211_X1 U21996 ( .C1(n18731), .C2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A(
        n18730), .B(n18729), .ZN(n18734) );
  AOI22_X1 U21997 ( .A1(n9704), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n18732), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n18733) );
  OAI211_X1 U21998 ( .C1(n13835), .C2(n18735), .A(n18734), .B(n18733), .ZN(
        n18746) );
  AOI22_X1 U21999 ( .A1(n18736), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n13878), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n18744) );
  AOI22_X1 U22000 ( .A1(n13279), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n18596), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n18743) );
  AOI22_X1 U22001 ( .A1(n18738), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n18737), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n18742) );
  AOI22_X1 U22002 ( .A1(n18740), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n18739), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n18741) );
  NAND4_X1 U22003 ( .A1(n18744), .A2(n18743), .A3(n18742), .A4(n18741), .ZN(
        n18745) );
  OR2_X1 U22004 ( .A1(n18746), .A2(n18745), .ZN(n18873) );
  NOR3_X1 U22005 ( .A1(n18747), .A2(n18787), .A3(P3_EBX_REG_10__SCAN_IN), .ZN(
        n18748) );
  AOI21_X1 U22006 ( .B1(n18749), .B2(n18873), .A(n18748), .ZN(n18750) );
  OAI21_X1 U22007 ( .B1(n18752), .B2(n18751), .A(n18750), .ZN(P3_U2693) );
  NOR2_X1 U22008 ( .A1(n18756), .A2(n18787), .ZN(n18757) );
  NAND2_X1 U22009 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n18757), .ZN(n18755) );
  NAND3_X1 U22010 ( .A1(n18755), .A2(P3_EBX_REG_7__SCAN_IN), .A3(n18777), .ZN(
        n18753) );
  OAI221_X1 U22011 ( .B1(n18755), .B2(P3_EBX_REG_7__SCAN_IN), .C1(n18777), 
        .C2(n18754), .A(n18753), .ZN(P3_U2696) );
  INV_X1 U22012 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n18759) );
  NAND2_X1 U22013 ( .A1(n18777), .A2(n18756), .ZN(n18760) );
  AOI22_X1 U22014 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n18749), .B1(
        n18757), .B2(n18759), .ZN(n18758) );
  OAI21_X1 U22015 ( .B1(n18759), .B2(n18760), .A(n18758), .ZN(P3_U2697) );
  AOI21_X1 U22016 ( .B1(n18785), .B2(n18762), .A(P3_EBX_REG_5__SCAN_IN), .ZN(
        n18761) );
  OAI22_X1 U22017 ( .A1(n18761), .A2(n18760), .B1(n17707), .B2(n18770), .ZN(
        P3_U2698) );
  INV_X1 U22018 ( .A(n18762), .ZN(n18766) );
  NOR2_X1 U22019 ( .A1(n18763), .A2(n18780), .ZN(n18775) );
  NAND2_X1 U22020 ( .A1(P3_EBX_REG_3__SCAN_IN), .A2(n18775), .ZN(n18769) );
  OAI21_X1 U22021 ( .B1(n18749), .B2(n18764), .A(n18769), .ZN(n18765) );
  OAI21_X1 U22022 ( .B1(n18780), .B2(n18766), .A(n18765), .ZN(n18767) );
  OAI21_X1 U22023 ( .B1(n18777), .B2(n18768), .A(n18767), .ZN(P3_U2699) );
  OAI211_X1 U22024 ( .C1(n18775), .C2(P3_EBX_REG_3__SCAN_IN), .A(n18770), .B(
        n18769), .ZN(n18771) );
  OAI21_X1 U22025 ( .B1(n18777), .B2(n18772), .A(n18771), .ZN(P3_U2700) );
  OR2_X1 U22026 ( .A1(n18787), .A2(n18773), .ZN(n18774) );
  AOI21_X1 U22027 ( .B1(n18785), .B2(n18774), .A(P3_EBX_REG_2__SCAN_IN), .ZN(
        n18776) );
  AOI211_X1 U22028 ( .C1(n18749), .C2(n13835), .A(n18776), .B(n18775), .ZN(
        P3_U2701) );
  OAI222_X1 U22029 ( .A1(n18781), .A2(n18780), .B1(n18779), .B2(n18785), .C1(
        n18778), .C2(n18777), .ZN(P3_U2702) );
  AOI22_X1 U22030 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18749), .B1(
        n18782), .B2(n18784), .ZN(n18783) );
  OAI21_X1 U22031 ( .B1(n18785), .B2(n18784), .A(n18783), .ZN(P3_U2703) );
  INV_X1 U22032 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n18961) );
  INV_X1 U22033 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n18957) );
  INV_X1 U22034 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n18950) );
  INV_X1 U22035 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n18948) );
  NAND2_X1 U22036 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n18824), .ZN(n18823) );
  NAND2_X1 U22037 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n18803), .ZN(n18798) );
  INV_X1 U22038 ( .A(n18798), .ZN(n18794) );
  NAND2_X1 U22039 ( .A1(n18794), .A2(P3_EAX_REG_30__SCAN_IN), .ZN(n18792) );
  NAND2_X1 U22040 ( .A1(n18886), .A2(n18798), .ZN(n18797) );
  OAI21_X1 U22041 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(n18789), .A(n18797), .ZN(
        n18790) );
  AOI22_X1 U22042 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n18858), .B1(
        P3_EAX_REG_31__SCAN_IN), .B2(n18790), .ZN(n18791) );
  OAI21_X1 U22043 ( .B1(P3_EAX_REG_31__SCAN_IN), .B2(n18792), .A(n18791), .ZN(
        P3_U2704) );
  INV_X1 U22044 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n18896) );
  AOI22_X1 U22045 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n18858), .B1(n18888), .B2(
        n18793), .ZN(n18796) );
  AOI22_X1 U22046 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n18827), .B1(n18794), .B2(
        n18896), .ZN(n18795) );
  OAI211_X1 U22047 ( .C1(n18797), .C2(n18896), .A(n18796), .B(n18795), .ZN(
        P3_U2705) );
  AOI22_X1 U22048 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n18827), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n18858), .ZN(n18800) );
  OAI211_X1 U22049 ( .C1(n18803), .C2(P3_EAX_REG_29__SCAN_IN), .A(n18886), .B(
        n18798), .ZN(n18799) );
  OAI211_X1 U22050 ( .C1(n18801), .C2(n18832), .A(n18800), .B(n18799), .ZN(
        P3_U2706) );
  AOI22_X1 U22051 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n18858), .B1(n18888), .B2(
        n18802), .ZN(n18806) );
  AOI211_X1 U22052 ( .C1(n18961), .C2(n18808), .A(n18803), .B(n18877), .ZN(
        n18804) );
  INV_X1 U22053 ( .A(n18804), .ZN(n18805) );
  OAI211_X1 U22054 ( .C1(n18863), .C2(n18807), .A(n18806), .B(n18805), .ZN(
        P3_U2707) );
  AOI22_X1 U22055 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n18827), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n18858), .ZN(n18810) );
  OAI211_X1 U22056 ( .C1(n9759), .C2(P3_EAX_REG_27__SCAN_IN), .A(n18886), .B(
        n18808), .ZN(n18809) );
  OAI211_X1 U22057 ( .C1(n18811), .C2(n18832), .A(n18810), .B(n18809), .ZN(
        P3_U2708) );
  AOI22_X1 U22058 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n18858), .B1(n18888), .B2(
        n18812), .ZN(n18815) );
  AOI211_X1 U22059 ( .C1(n18957), .C2(n18817), .A(n9759), .B(n18877), .ZN(
        n18813) );
  INV_X1 U22060 ( .A(n18813), .ZN(n18814) );
  OAI211_X1 U22061 ( .C1(n18863), .C2(n18816), .A(n18815), .B(n18814), .ZN(
        P3_U2709) );
  AOI22_X1 U22062 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n18827), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n18858), .ZN(n18820) );
  OAI211_X1 U22063 ( .C1(n18818), .C2(P3_EAX_REG_25__SCAN_IN), .A(n18886), .B(
        n18817), .ZN(n18819) );
  OAI211_X1 U22064 ( .C1(n18821), .C2(n18832), .A(n18820), .B(n18819), .ZN(
        P3_U2710) );
  AOI22_X1 U22065 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n18858), .B1(n18888), .B2(
        n18822), .ZN(n18826) );
  OAI211_X1 U22066 ( .C1(n18824), .C2(P3_EAX_REG_24__SCAN_IN), .A(n18886), .B(
        n18823), .ZN(n18825) );
  OAI211_X1 U22067 ( .C1(n18863), .C2(n18884), .A(n18826), .B(n18825), .ZN(
        P3_U2711) );
  AOI22_X1 U22068 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n18827), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n18858), .ZN(n18831) );
  OAI211_X1 U22069 ( .C1(P3_EAX_REG_23__SCAN_IN), .C2(n18829), .A(n18886), .B(
        n18828), .ZN(n18830) );
  OAI211_X1 U22070 ( .C1(n18833), .C2(n18832), .A(n18831), .B(n18830), .ZN(
        P3_U2712) );
  INV_X1 U22071 ( .A(n18834), .ZN(n18835) );
  AOI22_X1 U22072 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n18858), .B1(n18888), .B2(
        n18835), .ZN(n18839) );
  OAI21_X1 U22073 ( .B1(n18950), .B2(n18877), .A(n18837), .ZN(n18836) );
  OAI21_X1 U22074 ( .B1(n18950), .B2(n18837), .A(n18836), .ZN(n18838) );
  OAI211_X1 U22075 ( .C1(n13635), .C2(n18863), .A(n18839), .B(n18838), .ZN(
        P3_U2713) );
  AOI22_X1 U22076 ( .A1(n18858), .A2(BUF2_REG_20__SCAN_IN), .B1(n18888), .B2(
        n18840), .ZN(n18845) );
  INV_X1 U22077 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n18946) );
  AOI211_X1 U22078 ( .C1(n18946), .C2(n18842), .A(n18841), .B(n18877), .ZN(
        n18843) );
  INV_X1 U22079 ( .A(n18843), .ZN(n18844) );
  OAI211_X1 U22080 ( .C1(n18863), .C2(n13649), .A(n18845), .B(n18844), .ZN(
        P3_U2715) );
  AOI22_X1 U22081 ( .A1(n18858), .A2(BUF2_REG_18__SCAN_IN), .B1(n18888), .B2(
        n18846), .ZN(n18850) );
  INV_X1 U22082 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n18941) );
  NOR2_X1 U22083 ( .A1(n18941), .A2(n18847), .ZN(n18852) );
  OAI211_X1 U22084 ( .C1(n18852), .C2(P3_EAX_REG_18__SCAN_IN), .A(n18886), .B(
        n18848), .ZN(n18849) );
  OAI211_X1 U22085 ( .C1(n18863), .C2(n13655), .A(n18850), .B(n18849), .ZN(
        P3_U2717) );
  AOI22_X1 U22086 ( .A1(n18858), .A2(BUF2_REG_17__SCAN_IN), .B1(n18888), .B2(
        n18851), .ZN(n18856) );
  INV_X1 U22087 ( .A(n18852), .ZN(n18853) );
  OAI211_X1 U22088 ( .C1(n18854), .C2(P3_EAX_REG_17__SCAN_IN), .A(n18886), .B(
        n18853), .ZN(n18855) );
  OAI211_X1 U22089 ( .C1(n18863), .C2(n13632), .A(n18856), .B(n18855), .ZN(
        P3_U2718) );
  AOI22_X1 U22090 ( .A1(n18858), .A2(BUF2_REG_16__SCAN_IN), .B1(n18888), .B2(
        n18857), .ZN(n18862) );
  OAI211_X1 U22091 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n18860), .A(n18886), .B(
        n18859), .ZN(n18861) );
  OAI211_X1 U22092 ( .C1(n18863), .C2(n14163), .A(n18862), .B(n18861), .ZN(
        P3_U2719) );
  AOI22_X1 U22093 ( .A1(n18889), .A2(BUF2_REG_14__SCAN_IN), .B1(n18888), .B2(
        n18864), .ZN(n18867) );
  NAND3_X1 U22094 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(n18886), .A3(n18865), 
        .ZN(n18866) );
  OAI211_X1 U22095 ( .C1(P3_EAX_REG_14__SCAN_IN), .C2(n18868), .A(n18867), .B(
        n18866), .ZN(P3_U2721) );
  NAND2_X1 U22096 ( .A1(n18886), .A2(n18872), .ZN(n18876) );
  INV_X1 U22097 ( .A(n18869), .ZN(n18870) );
  AOI22_X1 U22098 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n18889), .B1(n18888), .B2(
        n18870), .ZN(n18871) );
  OAI221_X1 U22099 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n18872), .C1(n18986), 
        .C2(n18876), .A(n18871), .ZN(P3_U2724) );
  AOI22_X1 U22100 ( .A1(n18889), .A2(BUF2_REG_10__SCAN_IN), .B1(n18888), .B2(
        n18873), .ZN(n18874) );
  OAI221_X1 U22101 ( .B1(n18876), .B2(n18984), .C1(n18876), .C2(n18875), .A(
        n18874), .ZN(P3_U2725) );
  AOI211_X1 U22102 ( .C1(n18879), .C2(n18980), .A(n18878), .B(n18877), .ZN(
        n18880) );
  AOI21_X1 U22103 ( .B1(n18888), .B2(n18881), .A(n18880), .ZN(n18882) );
  OAI21_X1 U22104 ( .B1(n18884), .B2(n18883), .A(n18882), .ZN(P3_U2727) );
  AOI21_X1 U22105 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n18886), .A(n18885), .ZN(
        n18893) );
  AOI22_X1 U22106 ( .A1(n18889), .A2(BUF2_REG_7__SCAN_IN), .B1(n18888), .B2(
        n18887), .ZN(n18890) );
  OAI221_X1 U22107 ( .B1(n18893), .B2(n18892), .C1(n18893), .C2(n18891), .A(
        n18890), .ZN(P3_U2728) );
  NAND2_X1 U22108 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n19143), .ZN(n18930) );
  NOR2_X1 U22109 ( .A1(n21879), .A2(n18916), .ZN(P3_U2736) );
  NOR2_X1 U22110 ( .A1(n18934), .A2(n19565), .ZN(n18908) );
  INV_X2 U22111 ( .A(n18930), .ZN(n18932) );
  AOI22_X1 U22112 ( .A1(P3_UWORD_REG_14__SCAN_IN), .A2(n18932), .B1(n18923), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n18895) );
  OAI21_X1 U22113 ( .B1(n18896), .B2(n18912), .A(n18895), .ZN(P3_U2737) );
  INV_X1 U22114 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n18963) );
  AOI22_X1 U22115 ( .A1(n18932), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n18923), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n18897) );
  OAI21_X1 U22116 ( .B1(n18963), .B2(n18912), .A(n18897), .ZN(P3_U2738) );
  AOI22_X1 U22117 ( .A1(n18932), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n18923), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n18898) );
  OAI21_X1 U22118 ( .B1(n18961), .B2(n18912), .A(n18898), .ZN(P3_U2739) );
  INV_X1 U22119 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n18959) );
  AOI22_X1 U22120 ( .A1(n18932), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n18923), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n18899) );
  OAI21_X1 U22121 ( .B1(n18959), .B2(n18912), .A(n18899), .ZN(P3_U2740) );
  AOI22_X1 U22122 ( .A1(n18932), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n18923), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n18900) );
  OAI21_X1 U22123 ( .B1(n18957), .B2(n18912), .A(n18900), .ZN(P3_U2741) );
  INV_X1 U22124 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n21680) );
  AOI22_X1 U22125 ( .A1(n18932), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n18923), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n18901) );
  OAI21_X1 U22126 ( .B1(n21680), .B2(n18912), .A(n18901), .ZN(P3_U2742) );
  INV_X1 U22127 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n18954) );
  AOI22_X1 U22128 ( .A1(n18932), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n18923), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n18902) );
  OAI21_X1 U22129 ( .B1(n18954), .B2(n18912), .A(n18902), .ZN(P3_U2743) );
  INV_X1 U22130 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n18952) );
  AOI22_X1 U22131 ( .A1(n18932), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n18923), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n18903) );
  OAI21_X1 U22132 ( .B1(n18952), .B2(n18912), .A(n18903), .ZN(P3_U2744) );
  AOI22_X1 U22133 ( .A1(n18932), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n18923), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n18904) );
  OAI21_X1 U22134 ( .B1(n18950), .B2(n18912), .A(n18904), .ZN(P3_U2745) );
  AOI22_X1 U22135 ( .A1(n18932), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n18923), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n18905) );
  OAI21_X1 U22136 ( .B1(n18948), .B2(n18912), .A(n18905), .ZN(P3_U2746) );
  AOI22_X1 U22137 ( .A1(n18932), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n18923), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n18906) );
  OAI21_X1 U22138 ( .B1(n18946), .B2(n18912), .A(n18906), .ZN(P3_U2747) );
  INV_X1 U22139 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n18944) );
  AOI22_X1 U22140 ( .A1(n18932), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n18923), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n18907) );
  OAI21_X1 U22141 ( .B1(n18944), .B2(n18912), .A(n18907), .ZN(P3_U2748) );
  INV_X1 U22142 ( .A(P3_UWORD_REG_2__SCAN_IN), .ZN(n21745) );
  AOI22_X1 U22143 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n18908), .B1(n18923), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n18909) );
  OAI21_X1 U22144 ( .B1(n21745), .B2(n18930), .A(n18909), .ZN(P3_U2749) );
  AOI22_X1 U22145 ( .A1(n18932), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n18923), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n18910) );
  OAI21_X1 U22146 ( .B1(n18941), .B2(n18912), .A(n18910), .ZN(P3_U2750) );
  INV_X1 U22147 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n18939) );
  AOI22_X1 U22148 ( .A1(n18932), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n18923), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n18911) );
  OAI21_X1 U22149 ( .B1(n18939), .B2(n18912), .A(n18911), .ZN(P3_U2751) );
  AOI22_X1 U22150 ( .A1(n18932), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n18923), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n18913) );
  OAI21_X1 U22151 ( .B1(n18997), .B2(n18934), .A(n18913), .ZN(P3_U2752) );
  INV_X1 U22152 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n18993) );
  AOI22_X1 U22153 ( .A1(n18932), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n18923), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n18914) );
  OAI21_X1 U22154 ( .B1(n18993), .B2(n18934), .A(n18914), .ZN(P3_U2753) );
  INV_X1 U22155 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n18991) );
  AOI22_X1 U22156 ( .A1(n18932), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n18923), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n18915) );
  OAI21_X1 U22157 ( .B1(n18991), .B2(n18934), .A(n18915), .ZN(P3_U2754) );
  INV_X1 U22158 ( .A(P3_DATAO_REG_12__SCAN_IN), .ZN(n21696) );
  INV_X1 U22159 ( .A(P3_LWORD_REG_12__SCAN_IN), .ZN(n21762) );
  OAI222_X1 U22160 ( .A1(n18934), .A2(n18917), .B1(n18916), .B2(n21696), .C1(
        n18930), .C2(n21762), .ZN(P3_U2755) );
  AOI22_X1 U22161 ( .A1(n18932), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n18923), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n18918) );
  OAI21_X1 U22162 ( .B1(n18986), .B2(n18934), .A(n18918), .ZN(P3_U2756) );
  AOI22_X1 U22163 ( .A1(n18932), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n18923), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n18919) );
  OAI21_X1 U22164 ( .B1(n18984), .B2(n18934), .A(n18919), .ZN(P3_U2757) );
  AOI22_X1 U22165 ( .A1(n18932), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n18923), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n18920) );
  OAI21_X1 U22166 ( .B1(n18982), .B2(n18934), .A(n18920), .ZN(P3_U2758) );
  AOI22_X1 U22167 ( .A1(n18932), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n18923), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n18921) );
  OAI21_X1 U22168 ( .B1(n18980), .B2(n18934), .A(n18921), .ZN(P3_U2759) );
  AOI22_X1 U22169 ( .A1(n18932), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n18923), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n18922) );
  OAI21_X1 U22170 ( .B1(n18978), .B2(n18934), .A(n18922), .ZN(P3_U2760) );
  AOI22_X1 U22171 ( .A1(n18932), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n18923), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n18924) );
  OAI21_X1 U22172 ( .B1(n18976), .B2(n18934), .A(n18924), .ZN(P3_U2761) );
  INV_X1 U22173 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n18974) );
  AOI22_X1 U22174 ( .A1(n18932), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n18923), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n18925) );
  OAI21_X1 U22175 ( .B1(n18974), .B2(n18934), .A(n18925), .ZN(P3_U2762) );
  INV_X1 U22176 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n18972) );
  AOI22_X1 U22177 ( .A1(n18932), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n18923), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n18926) );
  OAI21_X1 U22178 ( .B1(n18972), .B2(n18934), .A(n18926), .ZN(P3_U2763) );
  INV_X1 U22179 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n18970) );
  AOI22_X1 U22180 ( .A1(n18932), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n18923), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n18927) );
  OAI21_X1 U22181 ( .B1(n18970), .B2(n18934), .A(n18927), .ZN(P3_U2764) );
  INV_X1 U22182 ( .A(P3_LWORD_REG_2__SCAN_IN), .ZN(n21900) );
  AOI22_X1 U22183 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n18928), .B1(n18923), .B2(
        P3_DATAO_REG_2__SCAN_IN), .ZN(n18929) );
  OAI21_X1 U22184 ( .B1(n21900), .B2(n18930), .A(n18929), .ZN(P3_U2765) );
  AOI22_X1 U22185 ( .A1(n18932), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n18923), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n18931) );
  OAI21_X1 U22186 ( .B1(n14165), .B2(n18934), .A(n18931), .ZN(P3_U2766) );
  AOI22_X1 U22187 ( .A1(n18932), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n18923), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n18933) );
  OAI21_X1 U22188 ( .B1(n18966), .B2(n18934), .A(n18933), .ZN(P3_U2767) );
  INV_X1 U22189 ( .A(n20161), .ZN(n20152) );
  AOI21_X1 U22190 ( .B1(n20150), .B2(n20152), .A(n18935), .ZN(n18936) );
  NAND2_X2 U22191 ( .A1(n20041), .A2(n18936), .ZN(n18996) );
  NAND2_X2 U22192 ( .A1(n18937), .A2(n18936), .ZN(n18994) );
  AOI22_X1 U22193 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n9841), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n18994), .ZN(n18938) );
  OAI21_X1 U22194 ( .B1(n18939), .B2(n18996), .A(n18938), .ZN(P3_U2768) );
  AOI22_X1 U22195 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n9841), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n18994), .ZN(n18940) );
  OAI21_X1 U22196 ( .B1(n18941), .B2(n18996), .A(n18940), .ZN(P3_U2769) );
  INV_X1 U22197 ( .A(n18994), .ZN(n18989) );
  AOI22_X1 U22198 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n9841), .B1(
        P3_EAX_REG_18__SCAN_IN), .B2(n18987), .ZN(n18942) );
  OAI21_X1 U22199 ( .B1(n18989), .B2(n21745), .A(n18942), .ZN(P3_U2770) );
  AOI22_X1 U22200 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n9841), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n18994), .ZN(n18943) );
  OAI21_X1 U22201 ( .B1(n18944), .B2(n18996), .A(n18943), .ZN(P3_U2771) );
  AOI22_X1 U22202 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n9841), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n18994), .ZN(n18945) );
  OAI21_X1 U22203 ( .B1(n18946), .B2(n18996), .A(n18945), .ZN(P3_U2772) );
  AOI22_X1 U22204 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n9841), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n18994), .ZN(n18947) );
  OAI21_X1 U22205 ( .B1(n18948), .B2(n18996), .A(n18947), .ZN(P3_U2773) );
  AOI22_X1 U22206 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n9841), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n18994), .ZN(n18949) );
  OAI21_X1 U22207 ( .B1(n18950), .B2(n18996), .A(n18949), .ZN(P3_U2774) );
  AOI22_X1 U22208 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n9841), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n18994), .ZN(n18951) );
  OAI21_X1 U22209 ( .B1(n18952), .B2(n18996), .A(n18951), .ZN(P3_U2775) );
  AOI22_X1 U22210 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n9841), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n18994), .ZN(n18953) );
  OAI21_X1 U22211 ( .B1(n18954), .B2(n18996), .A(n18953), .ZN(P3_U2776) );
  AOI22_X1 U22212 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n9841), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n18994), .ZN(n18955) );
  OAI21_X1 U22213 ( .B1(n21680), .B2(n18996), .A(n18955), .ZN(P3_U2777) );
  AOI22_X1 U22214 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n9841), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n18994), .ZN(n18956) );
  OAI21_X1 U22215 ( .B1(n18957), .B2(n18996), .A(n18956), .ZN(P3_U2778) );
  AOI22_X1 U22216 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n9841), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n18994), .ZN(n18958) );
  OAI21_X1 U22217 ( .B1(n18959), .B2(n18996), .A(n18958), .ZN(P3_U2779) );
  AOI22_X1 U22218 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n9841), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n18994), .ZN(n18960) );
  OAI21_X1 U22219 ( .B1(n18961), .B2(n18996), .A(n18960), .ZN(P3_U2780) );
  AOI22_X1 U22220 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n9841), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n18994), .ZN(n18962) );
  OAI21_X1 U22221 ( .B1(n18963), .B2(n18996), .A(n18962), .ZN(P3_U2781) );
  INV_X1 U22222 ( .A(P3_UWORD_REG_14__SCAN_IN), .ZN(n21789) );
  AOI22_X1 U22223 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n9841), .B1(
        P3_EAX_REG_30__SCAN_IN), .B2(n18987), .ZN(n18964) );
  OAI21_X1 U22224 ( .B1(n18989), .B2(n21789), .A(n18964), .ZN(P3_U2782) );
  AOI22_X1 U22225 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n9841), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n18994), .ZN(n18965) );
  OAI21_X1 U22226 ( .B1(n18966), .B2(n18996), .A(n18965), .ZN(P3_U2783) );
  AOI22_X1 U22227 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n9841), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n18994), .ZN(n18967) );
  OAI21_X1 U22228 ( .B1(n14165), .B2(n18996), .A(n18967), .ZN(P3_U2784) );
  AOI22_X1 U22229 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n9841), .B1(
        P3_EAX_REG_2__SCAN_IN), .B2(n18987), .ZN(n18968) );
  OAI21_X1 U22230 ( .B1(n18989), .B2(n21900), .A(n18968), .ZN(P3_U2785) );
  AOI22_X1 U22231 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n9841), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n18994), .ZN(n18969) );
  OAI21_X1 U22232 ( .B1(n18970), .B2(n18996), .A(n18969), .ZN(P3_U2786) );
  AOI22_X1 U22233 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n9841), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n18994), .ZN(n18971) );
  OAI21_X1 U22234 ( .B1(n18972), .B2(n18996), .A(n18971), .ZN(P3_U2787) );
  AOI22_X1 U22235 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n9841), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n18994), .ZN(n18973) );
  OAI21_X1 U22236 ( .B1(n18974), .B2(n18996), .A(n18973), .ZN(P3_U2788) );
  AOI22_X1 U22237 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n9841), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n18994), .ZN(n18975) );
  OAI21_X1 U22238 ( .B1(n18976), .B2(n18996), .A(n18975), .ZN(P3_U2789) );
  AOI22_X1 U22239 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n9841), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n18994), .ZN(n18977) );
  OAI21_X1 U22240 ( .B1(n18978), .B2(n18996), .A(n18977), .ZN(P3_U2790) );
  AOI22_X1 U22241 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n9841), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n18994), .ZN(n18979) );
  OAI21_X1 U22242 ( .B1(n18980), .B2(n18996), .A(n18979), .ZN(P3_U2791) );
  AOI22_X1 U22243 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n9841), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n18994), .ZN(n18981) );
  OAI21_X1 U22244 ( .B1(n18982), .B2(n18996), .A(n18981), .ZN(P3_U2792) );
  AOI22_X1 U22245 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n9841), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n18994), .ZN(n18983) );
  OAI21_X1 U22246 ( .B1(n18984), .B2(n18996), .A(n18983), .ZN(P3_U2793) );
  AOI22_X1 U22247 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n9841), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n18994), .ZN(n18985) );
  OAI21_X1 U22248 ( .B1(n18986), .B2(n18996), .A(n18985), .ZN(P3_U2794) );
  AOI22_X1 U22249 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n9841), .B1(
        P3_EAX_REG_12__SCAN_IN), .B2(n18987), .ZN(n18988) );
  OAI21_X1 U22250 ( .B1(n18989), .B2(n21762), .A(n18988), .ZN(P3_U2795) );
  AOI22_X1 U22251 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n9841), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n18994), .ZN(n18990) );
  OAI21_X1 U22252 ( .B1(n18991), .B2(n18996), .A(n18990), .ZN(P3_U2796) );
  AOI22_X1 U22253 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n9841), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n18994), .ZN(n18992) );
  OAI21_X1 U22254 ( .B1(n18993), .B2(n18996), .A(n18992), .ZN(P3_U2797) );
  AOI22_X1 U22255 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n9841), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n18994), .ZN(n18995) );
  OAI21_X1 U22256 ( .B1(n18997), .B2(n18996), .A(n18995), .ZN(P3_U2798) );
  OAI21_X1 U22257 ( .B1(n18999), .B2(n19289), .A(n18998), .ZN(n19287) );
  NOR2_X1 U22258 ( .A1(n19442), .A2(n20114), .ZN(n19286) );
  INV_X1 U22259 ( .A(n19000), .ZN(n19001) );
  NOR2_X1 U22260 ( .A1(n19067), .A2(n19001), .ZN(n19006) );
  AOI21_X1 U22261 ( .B1(n19002), .B2(n19945), .A(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n19003) );
  OAI22_X1 U22262 ( .A1(n19006), .A2(n19005), .B1(n19004), .B2(n19003), .ZN(
        n19007) );
  AOI211_X1 U22263 ( .C1(n19287), .C2(n19191), .A(n19286), .B(n19007), .ZN(
        n19008) );
  OAI221_X1 U22264 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n19010), 
        .C1(n19289), .C2(n19009), .A(n19008), .ZN(P3_U2804) );
  AOI22_X1 U22265 ( .A1(n19067), .A2(n19012), .B1(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n19011), .ZN(n19025) );
  NAND2_X1 U22266 ( .A1(n19032), .A2(n19296), .ZN(n19014) );
  INV_X1 U22267 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n19013) );
  XOR2_X1 U22268 ( .A(n19014), .B(n19013), .Z(n19294) );
  NOR2_X1 U22269 ( .A1(n19042), .A2(n19291), .ZN(n19015) );
  XNOR2_X1 U22270 ( .A(n19015), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n19301) );
  INV_X1 U22271 ( .A(n19016), .ZN(n19018) );
  NOR2_X1 U22272 ( .A1(n19018), .A2(n19017), .ZN(n19019) );
  XNOR2_X1 U22273 ( .A(n19019), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n19305) );
  OAI22_X1 U22274 ( .A1(n19189), .A2(n19301), .B1(n19109), .B2(n19305), .ZN(
        n19020) );
  AOI21_X1 U22275 ( .B1(n19275), .B2(n19294), .A(n19020), .ZN(n19024) );
  NAND2_X1 U22276 ( .A1(n19494), .A2(P3_REIP_REG_25__SCAN_IN), .ZN(n19303) );
  OAI211_X1 U22277 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(n19022), .B(n19021), .ZN(n19023) );
  NAND4_X1 U22278 ( .A1(n19025), .A2(n19024), .A3(n19303), .A4(n19023), .ZN(
        P3_U2805) );
  INV_X1 U22279 ( .A(n19026), .ZN(n19076) );
  INV_X1 U22280 ( .A(n19027), .ZN(n19028) );
  AOI21_X1 U22281 ( .B1(n19118), .B2(n19028), .A(n19047), .ZN(n19029) );
  AOI211_X1 U22282 ( .C1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n19030), .A(
        n19076), .B(n19029), .ZN(n19031) );
  XNOR2_X1 U22283 ( .A(n19031), .B(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n19310) );
  INV_X1 U22284 ( .A(n19032), .ZN(n19034) );
  AOI21_X1 U22285 ( .B1(n19035), .B2(n19034), .A(n19033), .ZN(n19040) );
  NAND2_X1 U22286 ( .A1(n19494), .A2(P3_REIP_REG_23__SCAN_IN), .ZN(n19309) );
  OAI21_X1 U22287 ( .B1(n19067), .B2(n19082), .A(n19036), .ZN(n19037) );
  OAI211_X1 U22288 ( .C1(n19038), .C2(n10497), .A(n19309), .B(n19037), .ZN(
        n19039) );
  AOI211_X1 U22289 ( .C1(n19041), .C2(n9816), .A(n19040), .B(n19039), .ZN(
        n19046) );
  INV_X1 U22290 ( .A(n19042), .ZN(n19044) );
  OAI211_X1 U22291 ( .C1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n19044), .A(
        n19141), .B(n19043), .ZN(n19045) );
  OAI211_X1 U22292 ( .C1(n19109), .C2(n19310), .A(n19046), .B(n19045), .ZN(
        P3_U2807) );
  AOI21_X1 U22293 ( .B1(n19325), .B2(n19326), .A(n19047), .ZN(n19048) );
  NOR2_X1 U22294 ( .A1(n19076), .A2(n19048), .ZN(n19049) );
  XNOR2_X1 U22295 ( .A(n19049), .B(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n19334) );
  AND2_X1 U22296 ( .A1(n19326), .A2(n19050), .ZN(n19061) );
  OAI21_X1 U22297 ( .B1(n19087), .B2(n19326), .A(n19086), .ZN(n19073) );
  OAI21_X1 U22298 ( .B1(n19051), .B2(n19098), .A(n19271), .ZN(n19052) );
  AOI21_X1 U22299 ( .B1(n19239), .B2(n19054), .A(n19052), .ZN(n19078) );
  OAI21_X1 U22300 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n19053), .A(
        n19078), .ZN(n19070) );
  AOI22_X1 U22301 ( .A1(n19494), .A2(P3_REIP_REG_22__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n19070), .ZN(n19057) );
  NOR2_X1 U22302 ( .A1(n19148), .A2(n19054), .ZN(n19072) );
  OAI211_X1 U22303 ( .C1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A(n19072), .B(n19055), .ZN(n19056) );
  OAI211_X1 U22304 ( .C1(n19159), .C2(n19058), .A(n19057), .B(n19056), .ZN(
        n19059) );
  AOI221_X1 U22305 ( .B1(n19061), .B2(n19060), .C1(n19073), .C2(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n19059), .ZN(n19062) );
  OAI21_X1 U22306 ( .B1(n19109), .B2(n19334), .A(n19062), .ZN(P3_U2808) );
  NAND2_X1 U22307 ( .A1(n19184), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n19117) );
  OAI22_X1 U22308 ( .A1(n19118), .A2(n19064), .B1(n19340), .B2(n19090), .ZN(
        n19065) );
  XNOR2_X1 U22309 ( .A(n19065), .B(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n19347) );
  AOI22_X1 U22310 ( .A1(n19494), .A2(P3_REIP_REG_21__SCAN_IN), .B1(n19067), 
        .B2(n19066), .ZN(n19068) );
  INV_X1 U22311 ( .A(n19068), .ZN(n19069) );
  AOI221_X1 U22312 ( .B1(n19072), .B2(n19071), .C1(n19070), .C2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(n19069), .ZN(n19075) );
  NOR2_X1 U22313 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n19340), .ZN(
        n19344) );
  NOR2_X1 U22314 ( .A1(n19337), .A2(n19123), .ZN(n19107) );
  AOI22_X1 U22315 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n19073), .B1(
        n19344), .B2(n19107), .ZN(n19074) );
  OAI211_X1 U22316 ( .C1(n19347), .C2(n19109), .A(n19075), .B(n19074), .ZN(
        P3_U2809) );
  INV_X1 U22317 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n21705) );
  AND2_X1 U22318 ( .A1(n19116), .A2(n21705), .ZN(n19093) );
  AOI211_X1 U22319 ( .C1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n19090), .A(
        n19093), .B(n19076), .ZN(n19077) );
  XOR2_X1 U22320 ( .A(n19315), .B(n19077), .Z(n19359) );
  INV_X1 U22321 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n19080) );
  AOI221_X1 U22322 ( .B1(n19081), .B2(n19080), .C1(n19079), .C2(n19080), .A(
        n19078), .ZN(n19085) );
  AOI21_X1 U22323 ( .B1(n19159), .B2(n19053), .A(n19083), .ZN(n19084) );
  AOI211_X1 U22324 ( .C1(P3_REIP_REG_20__SCAN_IN), .C2(n19494), .A(n19085), 
        .B(n19084), .ZN(n19089) );
  NOR2_X1 U22325 ( .A1(n19337), .A2(n21705), .ZN(n19349) );
  OAI21_X1 U22326 ( .B1(n19087), .B2(n19349), .A(n19086), .ZN(n19106) );
  NOR2_X1 U22327 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n21705), .ZN(
        n19348) );
  AOI22_X1 U22328 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n19106), .B1(
        n19107), .B2(n19348), .ZN(n19088) );
  OAI211_X1 U22329 ( .C1(n19109), .C2(n19359), .A(n19089), .B(n19088), .ZN(
        P3_U2810) );
  INV_X1 U22330 ( .A(n19118), .ZN(n19092) );
  INV_X1 U22331 ( .A(n19116), .ZN(n19091) );
  INV_X1 U22332 ( .A(n19090), .ZN(n19094) );
  AOI21_X1 U22333 ( .B1(n19092), .B2(n19091), .A(n19094), .ZN(n19096) );
  AOI21_X1 U22334 ( .B1(n19118), .B2(n21705), .A(n19093), .ZN(n19095) );
  OAI22_X1 U22335 ( .A1(n19096), .A2(n21705), .B1(n19095), .B2(n19094), .ZN(
        n19365) );
  OAI21_X1 U22336 ( .B1(n19099), .B2(n19098), .A(n19097), .ZN(n19113) );
  AOI22_X1 U22337 ( .A1(n19494), .A2(P3_REIP_REG_19__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n19113), .ZN(n19103) );
  NOR2_X1 U22338 ( .A1(n19148), .A2(n19100), .ZN(n19115) );
  OAI211_X1 U22339 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n19115), .B(n19101), .ZN(n19102) );
  OAI211_X1 U22340 ( .C1(n19159), .C2(n19104), .A(n19103), .B(n19102), .ZN(
        n19105) );
  AOI221_X1 U22341 ( .B1(n19107), .B2(n21705), .C1(n19106), .C2(
        P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A(n19105), .ZN(n19108) );
  OAI21_X1 U22342 ( .B1(n19365), .B2(n19109), .A(n19108), .ZN(P3_U2811) );
  NAND2_X1 U22343 ( .A1(n19110), .A2(n19368), .ZN(n19374) );
  OAI22_X1 U22344 ( .A1(n19442), .A2(n20101), .B1(n19159), .B2(n19111), .ZN(
        n19112) );
  AOI221_X1 U22345 ( .B1(n19115), .B2(n19114), .C1(n19113), .C2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(n19112), .ZN(n19122) );
  NAND2_X1 U22346 ( .A1(n19117), .A2(n19116), .ZN(n19119) );
  XOR2_X1 U22347 ( .A(n19119), .B(n19118), .Z(n19369) );
  AOI22_X1 U22348 ( .A1(n19369), .A2(n19191), .B1(n19120), .B2(
        P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n19121) );
  OAI211_X1 U22349 ( .C1(n19123), .C2(n19374), .A(n19122), .B(n19121), .ZN(
        P3_U2812) );
  NOR2_X1 U22350 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n19124), .ZN(
        n19395) );
  NAND2_X1 U22351 ( .A1(n19275), .A2(n19385), .ZN(n19138) );
  OAI22_X1 U22352 ( .A1(n19442), .A2(n20095), .B1(n19159), .B2(n19125), .ZN(
        n19126) );
  AOI221_X1 U22353 ( .B1(n19129), .B2(n19128), .C1(n19127), .C2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(n19126), .ZN(n19137) );
  NAND3_X1 U22354 ( .A1(n19130), .A2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        n19139), .ZN(n19131) );
  AOI21_X1 U22355 ( .B1(n19132), .B2(n19131), .A(n19409), .ZN(n19133) );
  XNOR2_X1 U22356 ( .A(n19133), .B(n19400), .ZN(n19396) );
  OR2_X1 U22357 ( .A1(n19134), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n19391) );
  AOI22_X1 U22358 ( .A1(n19396), .A2(n19191), .B1(n19135), .B2(n19391), .ZN(
        n19136) );
  OAI211_X1 U22359 ( .C1(n19395), .C2(n19138), .A(n19137), .B(n19136), .ZN(
        P3_U2815) );
  INV_X1 U22360 ( .A(n19402), .ZN(n19140) );
  NAND2_X1 U22361 ( .A1(n19139), .A2(n19426), .ZN(n19404) );
  AOI22_X1 U22362 ( .A1(n19141), .A2(n19140), .B1(n19275), .B2(n19404), .ZN(
        n19170) );
  OAI21_X1 U22363 ( .B1(n17848), .B2(n19145), .A(n19271), .ZN(n19197) );
  AOI21_X1 U22364 ( .B1(n19143), .B2(n19142), .A(n19197), .ZN(n19144) );
  OAI21_X1 U22365 ( .B1(n19146), .B2(n19145), .A(n19144), .ZN(n19161) );
  NOR2_X1 U22366 ( .A1(n19148), .A2(n19147), .ZN(n19163) );
  OAI211_X1 U22367 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(n19163), .B(n19149), .ZN(n19151) );
  NAND2_X1 U22368 ( .A1(n19494), .A2(P3_REIP_REG_13__SCAN_IN), .ZN(n19150) );
  OAI211_X1 U22369 ( .C1(n19159), .C2(n19152), .A(n19151), .B(n19150), .ZN(
        n19153) );
  AOI21_X1 U22370 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n19161), .A(
        n19153), .ZN(n19157) );
  AOI22_X1 U22371 ( .A1(n19154), .A2(n19165), .B1(n19184), .B2(n19402), .ZN(
        n19155) );
  XOR2_X1 U22372 ( .A(n14694), .B(n19155), .Z(n19410) );
  NOR2_X1 U22373 ( .A1(n19175), .A2(n19408), .ZN(n19167) );
  AOI22_X1 U22374 ( .A1(n19191), .A2(n19410), .B1(n19409), .B2(n19167), .ZN(
        n19156) );
  OAI211_X1 U22375 ( .C1(n19170), .C2(n14694), .A(n19157), .B(n19156), .ZN(
        P3_U2817) );
  INV_X1 U22376 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n20089) );
  OAI22_X1 U22377 ( .A1(n19442), .A2(n20089), .B1(n19159), .B2(n19158), .ZN(
        n19160) );
  AOI221_X1 U22378 ( .B1(n19163), .B2(n19162), .C1(n19161), .C2(
        P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A(n19160), .ZN(n19169) );
  OAI21_X1 U22379 ( .B1(n19408), .B2(n19173), .A(n19164), .ZN(n19166) );
  XNOR2_X1 U22380 ( .A(n19166), .B(n19165), .ZN(n19413) );
  AOI22_X1 U22381 ( .A1(n19191), .A2(n19413), .B1(n19167), .B2(n19165), .ZN(
        n19168) );
  OAI211_X1 U22382 ( .C1(n19170), .C2(n19165), .A(n19169), .B(n19168), .ZN(
        P3_U2818) );
  AOI22_X1 U22383 ( .A1(n19494), .A2(P3_REIP_REG_10__SCAN_IN), .B1(n19171), 
        .B2(n19243), .ZN(n19182) );
  OAI21_X1 U22384 ( .B1(n19173), .B2(n10263), .A(n19172), .ZN(n19174) );
  XOR2_X1 U22385 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B(n19174), .Z(
        n19438) );
  OAI21_X1 U22386 ( .B1(n19175), .B2(n10263), .A(n19445), .ZN(n19176) );
  AOI22_X1 U22387 ( .A1(n19191), .A2(n19438), .B1(n19177), .B2(n19176), .ZN(
        n19181) );
  OAI211_X1 U22388 ( .C1(n19179), .C2(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n19278), .B(n19178), .ZN(n19180) );
  NAND3_X1 U22389 ( .A1(n19182), .A2(n19181), .A3(n19180), .ZN(P3_U2820) );
  AOI22_X1 U22390 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n19197), .B1(
        n19183), .B2(n19243), .ZN(n19196) );
  MUX2_X1 U22391 ( .A(n19185), .B(n19475), .S(n19184), .Z(n19186) );
  NAND2_X1 U22392 ( .A1(n19186), .A2(n9752), .ZN(n19477) );
  OAI21_X1 U22393 ( .B1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n19188), .A(
        n19187), .ZN(n19472) );
  OAI22_X1 U22394 ( .A1(n19472), .A2(n19267), .B1(n19189), .B2(n19475), .ZN(
        n19190) );
  AOI21_X1 U22395 ( .B1(n19191), .B2(n19477), .A(n19190), .ZN(n19195) );
  NAND2_X1 U22396 ( .A1(n19494), .A2(P3_REIP_REG_8__SCAN_IN), .ZN(n19480) );
  OAI211_X1 U22397 ( .C1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(n19193), .A(
        n19945), .B(n19192), .ZN(n19194) );
  NAND4_X1 U22398 ( .A1(n19196), .A2(n19195), .A3(n19480), .A4(n19194), .ZN(
        P3_U2822) );
  NOR2_X1 U22399 ( .A1(n19442), .A2(n20081), .ZN(n19484) );
  AOI221_X1 U22400 ( .B1(n19199), .B2(n19198), .C1(n19197), .C2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A(n19484), .ZN(n19208) );
  AOI21_X1 U22401 ( .B1(n19202), .B2(n19201), .A(n19200), .ZN(n19203) );
  XOR2_X1 U22402 ( .A(n19203), .B(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .Z(
        n19483) );
  OAI21_X1 U22403 ( .B1(n19205), .B2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n19204), .ZN(n19206) );
  INV_X1 U22404 ( .A(n19206), .ZN(n19486) );
  AOI22_X1 U22405 ( .A1(n19483), .A2(n19275), .B1(n19277), .B2(n19486), .ZN(
        n19207) );
  OAI211_X1 U22406 ( .C1(n19281), .C2(n19209), .A(n19208), .B(n19207), .ZN(
        P3_U2823) );
  OR2_X1 U22407 ( .A1(n19211), .A2(n19210), .ZN(n19212) );
  AND2_X1 U22408 ( .A1(n19213), .A2(n19212), .ZN(n19499) );
  NOR2_X1 U22409 ( .A1(n19217), .A2(n19594), .ZN(n19214) );
  AOI22_X1 U22410 ( .A1(n19277), .A2(n19499), .B1(n19218), .B2(n19214), .ZN(
        n19222) );
  OAI21_X1 U22411 ( .B1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n19216), .A(
        n19215), .ZN(n19501) );
  OAI21_X1 U22412 ( .B1(n19217), .B2(n19594), .A(n19278), .ZN(n19228) );
  OAI22_X1 U22413 ( .A1(n19267), .A2(n19501), .B1(n19218), .B2(n19228), .ZN(
        n19219) );
  AOI21_X1 U22414 ( .B1(n19220), .B2(n19243), .A(n19219), .ZN(n19221) );
  OAI211_X1 U22415 ( .C1(n19442), .C2(n21712), .A(n19222), .B(n19221), .ZN(
        P3_U2824) );
  OAI21_X1 U22416 ( .B1(n19225), .B2(n19224), .A(n19223), .ZN(n19506) );
  XNOR2_X1 U22417 ( .A(n19226), .B(n10259), .ZN(n19502) );
  INV_X1 U22418 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n21714) );
  NOR2_X1 U22419 ( .A1(n19442), .A2(n21714), .ZN(n19503) );
  AOI21_X1 U22420 ( .B1(n19227), .B2(n19271), .A(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n19229) );
  OAI22_X1 U22421 ( .A1(n19281), .A2(n19230), .B1(n19229), .B2(n19228), .ZN(
        n19231) );
  AOI211_X1 U22422 ( .C1(n19277), .C2(n19502), .A(n19503), .B(n19231), .ZN(
        n19232) );
  OAI21_X1 U22423 ( .B1(n19267), .B2(n19506), .A(n19232), .ZN(P3_U2825) );
  OAI21_X1 U22424 ( .B1(n19235), .B2(n19234), .A(n19233), .ZN(n19236) );
  INV_X1 U22425 ( .A(n19236), .ZN(n19512) );
  NOR2_X1 U22426 ( .A1(n19442), .A2(n20078), .ZN(n19511) );
  AOI21_X1 U22427 ( .B1(n19277), .B2(n19512), .A(n19511), .ZN(n19246) );
  AOI21_X1 U22428 ( .B1(n19239), .B2(n19238), .A(n19237), .ZN(n19258) );
  OAI21_X1 U22429 ( .B1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n19241), .A(
        n19240), .ZN(n19519) );
  OAI22_X1 U22430 ( .A1(n19258), .A2(n21869), .B1(n19267), .B2(n19519), .ZN(
        n19242) );
  AOI21_X1 U22431 ( .B1(n19244), .B2(n19243), .A(n19242), .ZN(n19245) );
  OAI211_X1 U22432 ( .C1(n19594), .C2(n19247), .A(n19246), .B(n19245), .ZN(
        P3_U2826) );
  NAND2_X1 U22433 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n19271), .ZN(
        n19256) );
  XOR2_X1 U22434 ( .A(n19248), .B(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .Z(
        n19526) );
  NAND2_X1 U22435 ( .A1(n19494), .A2(P3_REIP_REG_3__SCAN_IN), .ZN(n19520) );
  OAI21_X1 U22436 ( .B1(n19281), .B2(n19249), .A(n19520), .ZN(n19254) );
  OAI21_X1 U22437 ( .B1(n19252), .B2(n19251), .A(n19250), .ZN(n19531) );
  NOR2_X1 U22438 ( .A1(n19267), .A2(n19531), .ZN(n19253) );
  AOI211_X1 U22439 ( .C1(n19277), .C2(n19526), .A(n19254), .B(n19253), .ZN(
        n19255) );
  OAI221_X1 U22440 ( .B1(n19258), .B2(n19257), .C1(n19258), .C2(n19256), .A(
        n19255), .ZN(P3_U2827) );
  OAI21_X1 U22441 ( .B1(n19261), .B2(n19260), .A(n19259), .ZN(n19262) );
  INV_X1 U22442 ( .A(n19262), .ZN(n19544) );
  NAND2_X1 U22443 ( .A1(n19494), .A2(P3_REIP_REG_2__SCAN_IN), .ZN(n19548) );
  OAI21_X1 U22444 ( .B1(n19281), .B2(n19263), .A(n19548), .ZN(n19269) );
  OAI21_X1 U22445 ( .B1(n19266), .B2(n19265), .A(n19264), .ZN(n19542) );
  NOR2_X1 U22446 ( .A1(n19267), .A2(n19542), .ZN(n19268) );
  AOI211_X1 U22447 ( .C1(n19277), .C2(n19544), .A(n19269), .B(n19268), .ZN(
        n19270) );
  OAI221_X1 U22448 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n19594), .C1(
        n19272), .C2(n19271), .A(n19270), .ZN(P3_U2828) );
  AOI21_X1 U22449 ( .B1(n19275), .B2(n19274), .A(n19273), .ZN(n19280) );
  AOI22_X1 U22450 ( .A1(n19278), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B1(
        n19277), .B2(n19276), .ZN(n19279) );
  OAI211_X1 U22451 ( .C1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n19281), .A(
        n19280), .B(n19279), .ZN(P3_U2829) );
  OAI21_X1 U22452 ( .B1(n19282), .B2(n19289), .A(n19546), .ZN(n19283) );
  AOI21_X1 U22453 ( .B1(n19284), .B2(n19289), .A(n19283), .ZN(n19285) );
  AOI211_X1 U22454 ( .C1(n19287), .C2(n19478), .A(n19286), .B(n19285), .ZN(
        n19288) );
  OAI21_X1 U22455 ( .B1(n19289), .B2(n19551), .A(n19288), .ZN(P3_U2836) );
  NOR4_X1 U22456 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n19292), .A3(
        n19291), .A4(n19290), .ZN(n19293) );
  AOI21_X1 U22457 ( .B1(n19294), .B2(n20021), .A(n19293), .ZN(n19300) );
  AOI21_X1 U22458 ( .B1(n19296), .B2(n19295), .A(n19536), .ZN(n19298) );
  OAI21_X1 U22459 ( .B1(n19298), .B2(n19297), .A(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n19299) );
  OAI211_X1 U22460 ( .C1(n19301), .C2(n19476), .A(n19300), .B(n19299), .ZN(
        n19302) );
  AOI22_X1 U22461 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n19527), .B1(
        n19546), .B2(n19302), .ZN(n19304) );
  OAI211_X1 U22462 ( .C1(n19305), .C2(n19364), .A(n19304), .B(n19303), .ZN(
        P3_U2837) );
  OAI221_X1 U22463 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n19307), 
        .C1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n19551), .A(n19306), .ZN(
        n19308) );
  OAI211_X1 U22464 ( .C1(n19310), .C2(n19364), .A(n19309), .B(n19308), .ZN(
        P3_U2839) );
  OAI21_X1 U22465 ( .B1(n19368), .B2(n19311), .A(n20023), .ZN(n19312) );
  OAI221_X1 U22466 ( .B1(n19314), .B2(n19313), .C1(n19314), .C2(n19349), .A(
        n19312), .ZN(n19350) );
  AOI21_X1 U22467 ( .B1(n19315), .B2(n19454), .A(n19350), .ZN(n19316) );
  OAI21_X1 U22468 ( .B1(n19326), .B2(n19431), .A(n19316), .ZN(n19338) );
  INV_X1 U22469 ( .A(n19317), .ZN(n19318) );
  NAND2_X1 U22470 ( .A1(n19439), .A2(n19318), .ZN(n19320) );
  NAND2_X1 U22471 ( .A1(n19320), .A2(n19319), .ZN(n19321) );
  OR2_X1 U22472 ( .A1(n19338), .A2(n19321), .ZN(n19323) );
  AOI22_X1 U22473 ( .A1(n19323), .A2(n19546), .B1(n19322), .B2(n19385), .ZN(
        n19330) );
  OR2_X1 U22474 ( .A1(n19325), .A2(n19324), .ZN(n19329) );
  AOI21_X1 U22475 ( .B1(n19327), .B2(n19326), .A(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n19328) );
  AOI21_X1 U22476 ( .B1(n19330), .B2(n19329), .A(n19328), .ZN(n19331) );
  AOI21_X1 U22477 ( .B1(n19527), .B2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n19331), .ZN(n19333) );
  NAND2_X1 U22478 ( .A1(n19494), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n19332) );
  OAI211_X1 U22479 ( .C1(n19334), .C2(n19364), .A(n19333), .B(n19332), .ZN(
        P3_U2840) );
  NOR2_X1 U22480 ( .A1(n19368), .A2(n19335), .ZN(n19360) );
  NAND2_X1 U22481 ( .A1(n19336), .A2(n19450), .ZN(n19375) );
  AOI221_X1 U22482 ( .B1(n19337), .B2(n19428), .C1(n19375), .C2(n19428), .A(
        n19380), .ZN(n19354) );
  INV_X1 U22483 ( .A(n19355), .ZN(n19339) );
  AOI21_X1 U22484 ( .B1(n19340), .B2(n19339), .A(n19338), .ZN(n19342) );
  AOI211_X1 U22485 ( .C1(n19354), .C2(n19342), .A(n19494), .B(n19341), .ZN(
        n19343) );
  AOI21_X1 U22486 ( .B1(n19344), .B2(n19360), .A(n19343), .ZN(n19346) );
  NAND2_X1 U22487 ( .A1(n19494), .A2(P3_REIP_REG_21__SCAN_IN), .ZN(n19345) );
  OAI211_X1 U22488 ( .C1(n19347), .C2(n19364), .A(n19346), .B(n19345), .ZN(
        P3_U2841) );
  AOI22_X1 U22489 ( .A1(n19494), .A2(P3_REIP_REG_20__SCAN_IN), .B1(n19360), 
        .B2(n19348), .ZN(n19358) );
  INV_X1 U22490 ( .A(n19349), .ZN(n19352) );
  AOI21_X1 U22491 ( .B1(n19352), .B2(n19351), .A(n19350), .ZN(n19353) );
  AOI21_X1 U22492 ( .B1(n19354), .B2(n19353), .A(n19494), .ZN(n19361) );
  NOR3_X1 U22493 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n19355), .A3(
        n20151), .ZN(n19356) );
  OAI21_X1 U22494 ( .B1(n19361), .B2(n19356), .A(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n19357) );
  OAI211_X1 U22495 ( .C1(n19359), .C2(n19364), .A(n19358), .B(n19357), .ZN(
        P3_U2842) );
  AOI22_X1 U22496 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n19361), .B1(
        n19360), .B2(n21705), .ZN(n19363) );
  NAND2_X1 U22497 ( .A1(n19494), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n19362) );
  OAI211_X1 U22498 ( .C1(n19365), .C2(n19364), .A(n19363), .B(n19362), .ZN(
        P3_U2843) );
  INV_X1 U22499 ( .A(n19366), .ZN(n19384) );
  OAI21_X1 U22500 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n19465), .A(
        n19367), .ZN(n19371) );
  NOR2_X1 U22501 ( .A1(n19494), .A2(n19368), .ZN(n19370) );
  AOI22_X1 U22502 ( .A1(n19371), .A2(n19370), .B1(n19478), .B2(n19369), .ZN(
        n19373) );
  NAND2_X1 U22503 ( .A1(n19494), .A2(P3_REIP_REG_18__SCAN_IN), .ZN(n19372) );
  OAI211_X1 U22504 ( .C1(n19374), .C2(n19384), .A(n19373), .B(n19372), .ZN(
        P3_U2844) );
  OAI21_X1 U22505 ( .B1(n19428), .B2(n19400), .A(n19375), .ZN(n19378) );
  INV_X1 U22506 ( .A(n19387), .ZN(n19376) );
  NAND2_X1 U22507 ( .A1(n19439), .A2(n19376), .ZN(n19377) );
  NAND3_X1 U22508 ( .A1(n19379), .A2(n19378), .A3(n19377), .ZN(n19390) );
  OAI221_X1 U22509 ( .B1(n19380), .B2(n19467), .C1(n19380), .C2(n19390), .A(
        n19442), .ZN(n19383) );
  AOI22_X1 U22510 ( .A1(n19494), .A2(P3_REIP_REG_16__SCAN_IN), .B1(n19478), 
        .B2(n19381), .ZN(n19382) );
  OAI221_X1 U22511 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n19384), 
        .C1(n10019), .C2(n19383), .A(n19382), .ZN(P3_U2846) );
  NAND2_X1 U22512 ( .A1(n20021), .A2(n19385), .ZN(n19394) );
  NAND2_X1 U22513 ( .A1(n19387), .A2(n19386), .ZN(n19388) );
  NAND2_X1 U22514 ( .A1(n19388), .A2(n19400), .ZN(n19389) );
  AOI22_X1 U22515 ( .A1(n19392), .A2(n19391), .B1(n19390), .B2(n19389), .ZN(
        n19393) );
  OAI21_X1 U22516 ( .B1(n19395), .B2(n19394), .A(n19393), .ZN(n19397) );
  AOI22_X1 U22517 ( .A1(n19546), .A2(n19397), .B1(n19478), .B2(n19396), .ZN(
        n19399) );
  NAND2_X1 U22518 ( .A1(n19494), .A2(P3_REIP_REG_15__SCAN_IN), .ZN(n19398) );
  OAI211_X1 U22519 ( .C1(n19551), .C2(n19400), .A(n19399), .B(n19398), .ZN(
        P3_U2847) );
  INV_X1 U22520 ( .A(n19439), .ZN(n19405) );
  NAND2_X1 U22521 ( .A1(n20023), .A2(n19401), .ZN(n19422) );
  AOI21_X1 U22522 ( .B1(n19439), .B2(n19408), .A(n19440), .ZN(n19433) );
  OAI211_X1 U22523 ( .C1(n19402), .C2(n19476), .A(n19422), .B(n19433), .ZN(
        n19403) );
  AOI21_X1 U22524 ( .B1(n20021), .B2(n19404), .A(n19403), .ZN(n19415) );
  OAI211_X1 U22525 ( .C1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n19405), .A(
        n19546), .B(n19415), .ZN(n19406) );
  OAI21_X1 U22526 ( .B1(n19407), .B2(n19406), .A(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n19412) );
  NOR2_X1 U22527 ( .A1(n19408), .A2(n19461), .ZN(n19418) );
  AOI22_X1 U22528 ( .A1(n19478), .A2(n19410), .B1(n19409), .B2(n19418), .ZN(
        n19411) );
  OAI221_X1 U22529 ( .B1(n19494), .B2(n19412), .C1(n19442), .C2(n20091), .A(
        n19411), .ZN(P3_U2849) );
  AOI22_X1 U22530 ( .A1(n19494), .A2(P3_REIP_REG_12__SCAN_IN), .B1(n19478), 
        .B2(n19413), .ZN(n19420) );
  NOR2_X1 U22531 ( .A1(n19414), .A2(n19429), .ZN(n19416) );
  OAI211_X1 U22532 ( .C1(n19416), .C2(n19451), .A(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B(n19415), .ZN(n19417) );
  OAI211_X1 U22533 ( .C1(n19418), .C2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n19546), .B(n19417), .ZN(n19419) );
  OAI211_X1 U22534 ( .C1(n19551), .C2(n19165), .A(n19420), .B(n19419), .ZN(
        P3_U2850) );
  AOI22_X1 U22535 ( .A1(n19494), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n19478), 
        .B2(n19421), .ZN(n19436) );
  AND2_X1 U22536 ( .A1(n19546), .A2(n19422), .ZN(n19425) );
  OR2_X1 U22537 ( .A1(n19423), .A2(n19476), .ZN(n19424) );
  OAI211_X1 U22538 ( .C1(n19426), .C2(n19543), .A(n19425), .B(n19424), .ZN(
        n19427) );
  INV_X1 U22539 ( .A(n19427), .ZN(n19456) );
  OAI21_X1 U22540 ( .B1(n10263), .B2(n19429), .A(n19428), .ZN(n19430) );
  OAI211_X1 U22541 ( .C1(n19432), .C2(n19431), .A(n19456), .B(n19430), .ZN(
        n19443) );
  OAI21_X1 U22542 ( .B1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n19451), .A(
        n19433), .ZN(n19434) );
  OAI211_X1 U22543 ( .C1(n19443), .C2(n19434), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n19442), .ZN(n19435) );
  OAI211_X1 U22544 ( .C1(n19461), .C2(n19437), .A(n19436), .B(n19435), .ZN(
        P3_U2851) );
  AOI22_X1 U22545 ( .A1(n19494), .A2(P3_REIP_REG_10__SCAN_IN), .B1(n19478), 
        .B2(n19438), .ZN(n19449) );
  OAI21_X1 U22546 ( .B1(n10263), .B2(n19440), .A(n19439), .ZN(n19441) );
  INV_X1 U22547 ( .A(n19441), .ZN(n19444) );
  OAI211_X1 U22548 ( .C1(n19444), .C2(n19443), .A(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B(n19442), .ZN(n19448) );
  INV_X1 U22549 ( .A(n19461), .ZN(n19446) );
  NAND3_X1 U22550 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n19446), .A3(
        n19445), .ZN(n19447) );
  NAND3_X1 U22551 ( .A1(n19449), .A2(n19448), .A3(n19447), .ZN(P3_U2852) );
  AOI211_X1 U22552 ( .C1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .C2(n19451), .A(
        n19465), .B(n19450), .ZN(n19452) );
  AOI21_X1 U22553 ( .B1(n19454), .B2(n19453), .A(n19452), .ZN(n19455) );
  AOI211_X1 U22554 ( .C1(n19456), .C2(n19455), .A(n19494), .B(n10263), .ZN(
        n19457) );
  AOI211_X1 U22555 ( .C1(n19478), .C2(n19459), .A(n19458), .B(n19457), .ZN(
        n19460) );
  OAI21_X1 U22556 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n19461), .A(
        n19460), .ZN(P3_U2853) );
  INV_X1 U22557 ( .A(n19467), .ZN(n19469) );
  NOR2_X1 U22558 ( .A1(n19496), .A2(n19485), .ZN(n19468) );
  OR2_X1 U22559 ( .A1(n19536), .A2(n19462), .ZN(n19540) );
  OAI211_X1 U22560 ( .C1(n19465), .C2(n19464), .A(n19540), .B(n19463), .ZN(
        n19513) );
  AOI21_X1 U22561 ( .B1(n19467), .B2(n19466), .A(n19513), .ZN(n19492) );
  OAI21_X1 U22562 ( .B1(n19469), .B2(n19468), .A(n19492), .ZN(n19487) );
  AOI21_X1 U22563 ( .B1(n19470), .B2(n19487), .A(n19527), .ZN(n19482) );
  OAI22_X1 U22564 ( .A1(n19472), .A2(n19543), .B1(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n19471), .ZN(n19473) );
  INV_X1 U22565 ( .A(n19473), .ZN(n19474) );
  OAI21_X1 U22566 ( .B1(n19476), .B2(n19475), .A(n19474), .ZN(n19479) );
  AOI22_X1 U22567 ( .A1(n19546), .A2(n19479), .B1(n19478), .B2(n19477), .ZN(
        n19481) );
  OAI211_X1 U22568 ( .C1(n19482), .C2(n13316), .A(n19481), .B(n19480), .ZN(
        P3_U2854) );
  INV_X1 U22569 ( .A(n19483), .ZN(n19491) );
  AOI21_X1 U22570 ( .B1(n19527), .B2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n19484), .ZN(n19490) );
  NOR3_X1 U22571 ( .A1(n19523), .A2(n19522), .A3(n21791), .ZN(n19515) );
  NAND3_X1 U22572 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A3(n19515), .ZN(n19497) );
  OAI22_X1 U22573 ( .A1(n19497), .A2(n19496), .B1(n19522), .B2(n19485), .ZN(
        n19488) );
  AOI22_X1 U22574 ( .A1(n19488), .A2(n19487), .B1(n19545), .B2(n19486), .ZN(
        n19489) );
  OAI211_X1 U22575 ( .C1(n19530), .C2(n19491), .A(n19490), .B(n19489), .ZN(
        P3_U2855) );
  AOI21_X1 U22576 ( .B1(n19546), .B2(n19492), .A(n19494), .ZN(n19493) );
  INV_X1 U22577 ( .A(n19493), .ZN(n19509) );
  NAND2_X1 U22578 ( .A1(n19494), .A2(P3_REIP_REG_6__SCAN_IN), .ZN(n19495) );
  OAI221_X1 U22579 ( .B1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n19497), .C1(
        n19496), .C2(n19509), .A(n19495), .ZN(n19498) );
  AOI21_X1 U22580 ( .B1(n19545), .B2(n19499), .A(n19498), .ZN(n19500) );
  OAI21_X1 U22581 ( .B1(n19530), .B2(n19501), .A(n19500), .ZN(P3_U2856) );
  NAND2_X1 U22582 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n19515), .ZN(
        n19510) );
  NAND2_X1 U22583 ( .A1(n19545), .A2(n19502), .ZN(n19505) );
  INV_X1 U22584 ( .A(n19503), .ZN(n19504) );
  OAI211_X1 U22585 ( .C1(n19506), .C2(n19530), .A(n19505), .B(n19504), .ZN(
        n19507) );
  INV_X1 U22586 ( .A(n19507), .ZN(n19508) );
  OAI221_X1 U22587 ( .B1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n19510), .C1(
        n10259), .C2(n19509), .A(n19508), .ZN(P3_U2857) );
  AOI21_X1 U22588 ( .B1(n19545), .B2(n19512), .A(n19511), .ZN(n19518) );
  NOR2_X1 U22589 ( .A1(n21791), .A2(n19513), .ZN(n19521) );
  OAI21_X1 U22590 ( .B1(n19521), .B2(n19514), .A(n19551), .ZN(n19516) );
  INV_X1 U22591 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n21906) );
  AOI22_X1 U22592 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n19516), .B1(
        n19515), .B2(n21906), .ZN(n19517) );
  OAI211_X1 U22593 ( .C1(n19530), .C2(n19519), .A(n19518), .B(n19517), .ZN(
        P3_U2858) );
  INV_X1 U22594 ( .A(n19520), .ZN(n19525) );
  AOI211_X1 U22595 ( .C1(n19523), .C2(n21791), .A(n19522), .B(n19521), .ZN(
        n19524) );
  AOI211_X1 U22596 ( .C1(n19545), .C2(n19526), .A(n19525), .B(n19524), .ZN(
        n19529) );
  NAND2_X1 U22597 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n19527), .ZN(
        n19528) );
  OAI211_X1 U22598 ( .C1(n19531), .C2(n19530), .A(n19529), .B(n19528), .ZN(
        P3_U2859) );
  NAND2_X1 U22599 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n19537) );
  OAI21_X1 U22600 ( .B1(n19534), .B2(n19533), .A(n19532), .ZN(n19535) );
  OAI21_X1 U22601 ( .B1(n19537), .B2(n19536), .A(n19535), .ZN(n19538) );
  OAI222_X1 U22602 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n19539), .C1(n19550), .C2(
        n19538), .ZN(n19541) );
  OAI211_X1 U22603 ( .C1(n19543), .C2(n19542), .A(n19541), .B(n19540), .ZN(
        n19547) );
  AOI22_X1 U22604 ( .A1(n19547), .A2(n19546), .B1(n19545), .B2(n19544), .ZN(
        n19549) );
  OAI211_X1 U22605 ( .C1(n19551), .C2(n19550), .A(n19549), .B(n19548), .ZN(
        P3_U2860) );
  AOI21_X1 U22606 ( .B1(n19554), .B2(n19553), .A(n19552), .ZN(n20044) );
  OAI21_X1 U22607 ( .B1(n20044), .B2(n19593), .A(n19559), .ZN(n19555) );
  OAI221_X1 U22608 ( .B1(n11692), .B2(n20158), .C1(n11692), .C2(n19559), .A(
        n19555), .ZN(P3_U2863) );
  NAND2_X1 U22609 ( .A1(n11696), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19804) );
  INV_X1 U22610 ( .A(n19804), .ZN(n19782) );
  NAND2_X1 U22611 ( .A1(n20013), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n19739) );
  INV_X1 U22612 ( .A(n19739), .ZN(n19693) );
  NOR2_X1 U22613 ( .A1(n19782), .A2(n19693), .ZN(n19557) );
  OAI22_X1 U22614 ( .A1(n19558), .A2(n20013), .B1(n19557), .B2(n19556), .ZN(
        P3_U2866) );
  NOR2_X1 U22615 ( .A1(n19560), .A2(n19559), .ZN(P3_U2867) );
  NOR2_X1 U22616 ( .A1(n19594), .A2(n16849), .ZN(n19873) );
  NOR2_X1 U22617 ( .A1(n20013), .A2(n19715), .ZN(n19943) );
  INV_X1 U22618 ( .A(n19943), .ZN(n19938) );
  NOR2_X2 U22619 ( .A1(n19938), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19934) );
  INV_X1 U22620 ( .A(n19934), .ZN(n19607) );
  NOR2_X1 U22621 ( .A1(n11696), .A2(n20013), .ZN(n19875) );
  INV_X1 U22622 ( .A(n19875), .ZN(n19872) );
  NAND2_X1 U22623 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n11693), .ZN(
        n19784) );
  NOR2_X2 U22624 ( .A1(n19872), .A2(n19784), .ZN(n19976) );
  NAND2_X1 U22625 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n19945), .ZN(n19880) );
  INV_X1 U22626 ( .A(n19880), .ZN(n19940) );
  NOR2_X2 U22627 ( .A1(n19592), .A2(n14163), .ZN(n19941) );
  NAND2_X1 U22628 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19943), .ZN(
        n19631) );
  INV_X1 U22629 ( .A(n19631), .ZN(n19993) );
  NAND2_X1 U22630 ( .A1(n11693), .A2(n11692), .ZN(n20005) );
  NAND2_X1 U22631 ( .A1(n11696), .A2(n20013), .ZN(n19643) );
  NOR2_X2 U22632 ( .A1(n20005), .A2(n19643), .ZN(n19666) );
  NOR2_X1 U22633 ( .A1(n19993), .A2(n19666), .ZN(n19617) );
  NAND2_X1 U22634 ( .A1(n20151), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n19827) );
  INV_X1 U22635 ( .A(n19827), .ZN(n19939) );
  NOR2_X1 U22636 ( .A1(n19617), .A2(n19939), .ZN(n19586) );
  AOI22_X1 U22637 ( .A1(n19976), .A2(n19940), .B1(n19941), .B2(n19586), .ZN(
        n19567) );
  INV_X1 U22638 ( .A(n19592), .ZN(n19908) );
  NOR2_X1 U22639 ( .A1(n11692), .A2(n20134), .ZN(n19561) );
  NOR2_X1 U22640 ( .A1(n19934), .A2(n19976), .ZN(n19904) );
  OAI22_X1 U22641 ( .A1(n19561), .A2(n19617), .B1(n19904), .B2(n19905), .ZN(
        n19562) );
  NAND2_X1 U22642 ( .A1(n19908), .A2(n19562), .ZN(n19589) );
  NAND2_X1 U22643 ( .A1(n19564), .A2(n19563), .ZN(n19587) );
  NOR2_X2 U22644 ( .A1(n19565), .A2(n19587), .ZN(n19946) );
  AOI22_X1 U22645 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n19589), .B1(
        n19666), .B2(n19946), .ZN(n19566) );
  OAI211_X1 U22646 ( .C1(n19949), .C2(n19607), .A(n19567), .B(n19566), .ZN(
        P3_U2868) );
  INV_X1 U22647 ( .A(n19976), .ZN(n19998) );
  NOR2_X1 U22648 ( .A1(n16787), .A2(n19594), .ZN(n19911) );
  NAND2_X1 U22649 ( .A1(n19945), .A2(BUF2_REG_17__SCAN_IN), .ZN(n19914) );
  INV_X1 U22650 ( .A(n19914), .ZN(n19951) );
  NOR2_X2 U22651 ( .A1(n19592), .A2(n13632), .ZN(n19950) );
  AOI22_X1 U22652 ( .A1(n19934), .A2(n19951), .B1(n19586), .B2(n19950), .ZN(
        n19570) );
  NOR2_X2 U22653 ( .A1(n19568), .A2(n19587), .ZN(n19952) );
  AOI22_X1 U22654 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n19589), .B1(
        n19666), .B2(n19952), .ZN(n19569) );
  OAI211_X1 U22655 ( .C1(n19998), .C2(n19955), .A(n19570), .B(n19569), .ZN(
        P3_U2869) );
  NOR2_X1 U22656 ( .A1(n19594), .A2(n16835), .ZN(n19883) );
  INV_X1 U22657 ( .A(n19883), .ZN(n19961) );
  NAND2_X1 U22658 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n19945), .ZN(n19886) );
  INV_X1 U22659 ( .A(n19886), .ZN(n19956) );
  NOR2_X2 U22660 ( .A1(n19592), .A2(n13655), .ZN(n19957) );
  AOI22_X1 U22661 ( .A1(n19976), .A2(n19956), .B1(n19586), .B2(n19957), .ZN(
        n19573) );
  NOR2_X2 U22662 ( .A1(n19571), .A2(n19587), .ZN(n19958) );
  AOI22_X1 U22663 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n19589), .B1(
        n19666), .B2(n19958), .ZN(n19572) );
  OAI211_X1 U22664 ( .C1(n19607), .C2(n19961), .A(n19573), .B(n19572), .ZN(
        P3_U2870) );
  NAND2_X1 U22665 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n19877), .ZN(n19920) );
  NAND2_X1 U22666 ( .A1(n19945), .A2(BUF2_REG_19__SCAN_IN), .ZN(n19967) );
  INV_X1 U22667 ( .A(n19967), .ZN(n19917) );
  NOR2_X2 U22668 ( .A1(n19592), .A2(n13652), .ZN(n19962) );
  AOI22_X1 U22669 ( .A1(n19934), .A2(n19917), .B1(n19586), .B2(n19962), .ZN(
        n19576) );
  NOR2_X2 U22670 ( .A1(n19574), .A2(n19587), .ZN(n19964) );
  AOI22_X1 U22671 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19589), .B1(
        n19666), .B2(n19964), .ZN(n19575) );
  OAI211_X1 U22672 ( .C1(n19998), .C2(n19920), .A(n19576), .B(n19575), .ZN(
        P3_U2871) );
  NOR2_X1 U22673 ( .A1(n19594), .A2(n16823), .ZN(n19921) );
  INV_X1 U22674 ( .A(n19921), .ZN(n19973) );
  NAND2_X1 U22675 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n19945), .ZN(n19925) );
  INV_X1 U22676 ( .A(n19925), .ZN(n19968) );
  NOR2_X2 U22677 ( .A1(n19592), .A2(n13649), .ZN(n19969) );
  AOI22_X1 U22678 ( .A1(n19976), .A2(n19968), .B1(n19586), .B2(n19969), .ZN(
        n19579) );
  NOR2_X2 U22679 ( .A1(n19577), .A2(n19587), .ZN(n19970) );
  AOI22_X1 U22680 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n19589), .B1(
        n19666), .B2(n19970), .ZN(n19578) );
  OAI211_X1 U22681 ( .C1(n19607), .C2(n19973), .A(n19579), .B(n19578), .ZN(
        P3_U2872) );
  NAND2_X1 U22682 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n19945), .ZN(n19981) );
  NAND2_X1 U22683 ( .A1(n19945), .A2(BUF2_REG_21__SCAN_IN), .ZN(n19929) );
  INV_X1 U22684 ( .A(n19929), .ZN(n19975) );
  NOR2_X2 U22685 ( .A1(n19592), .A2(n13643), .ZN(n19974) );
  AOI22_X1 U22686 ( .A1(n19934), .A2(n19975), .B1(n19586), .B2(n19974), .ZN(
        n19582) );
  NOR2_X2 U22687 ( .A1(n19580), .A2(n19587), .ZN(n19977) );
  AOI22_X1 U22688 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19589), .B1(
        n19666), .B2(n19977), .ZN(n19581) );
  OAI211_X1 U22689 ( .C1(n19998), .C2(n19981), .A(n19582), .B(n19581), .ZN(
        P3_U2873) );
  NAND2_X1 U22690 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n19945), .ZN(n19897) );
  NAND2_X1 U22691 ( .A1(n19945), .A2(BUF2_REG_22__SCAN_IN), .ZN(n19987) );
  INV_X1 U22692 ( .A(n19987), .ZN(n19894) );
  NOR2_X2 U22693 ( .A1(n19592), .A2(n13635), .ZN(n19982) );
  AOI22_X1 U22694 ( .A1(n19934), .A2(n19894), .B1(n19586), .B2(n19982), .ZN(
        n19585) );
  NOR2_X2 U22695 ( .A1(n19583), .A2(n19587), .ZN(n19984) );
  AOI22_X1 U22696 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19589), .B1(
        n19666), .B2(n19984), .ZN(n19584) );
  OAI211_X1 U22697 ( .C1(n19998), .C2(n19897), .A(n19585), .B(n19584), .ZN(
        P3_U2874) );
  NOR2_X1 U22698 ( .A1(n19594), .A2(n16800), .ZN(n19898) );
  INV_X1 U22699 ( .A(n19898), .ZN(n19997) );
  NAND2_X1 U22700 ( .A1(n19945), .A2(BUF2_REG_31__SCAN_IN), .ZN(n19903) );
  INV_X1 U22701 ( .A(n19903), .ZN(n19991) );
  NOR2_X2 U22702 ( .A1(n19592), .A2(n13640), .ZN(n19989) );
  AOI22_X1 U22703 ( .A1(n19976), .A2(n19991), .B1(n19586), .B2(n19989), .ZN(
        n19591) );
  NOR2_X2 U22704 ( .A1(n19588), .A2(n19587), .ZN(n19992) );
  AOI22_X1 U22705 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19589), .B1(
        n19666), .B2(n19992), .ZN(n19590) );
  OAI211_X1 U22706 ( .C1(n19607), .C2(n19997), .A(n19591), .B(n19590), .ZN(
        P3_U2875) );
  NOR2_X1 U22707 ( .A1(n19593), .A2(n19592), .ZN(n19942) );
  NAND2_X1 U22708 ( .A1(n19942), .A2(n11693), .ZN(n19692) );
  OAI22_X1 U22709 ( .A1(n19594), .A2(n19938), .B1(n19643), .B2(n19692), .ZN(
        n19610) );
  NAND2_X1 U22710 ( .A1(n11693), .A2(n19827), .ZN(n19871) );
  NOR2_X1 U22711 ( .A1(n19643), .A2(n19871), .ZN(n19613) );
  AOI22_X1 U22712 ( .A1(n19873), .A2(n19993), .B1(n19941), .B2(n19613), .ZN(
        n19596) );
  NOR2_X1 U22713 ( .A1(n19643), .A2(n19784), .ZN(n19654) );
  AOI22_X1 U22714 ( .A1(n19934), .A2(n19940), .B1(n19946), .B2(n19688), .ZN(
        n19595) );
  OAI211_X1 U22715 ( .C1(n21742), .C2(n19610), .A(n19596), .B(n19595), .ZN(
        P3_U2876) );
  AOI22_X1 U22716 ( .A1(n19993), .A2(n19951), .B1(n19950), .B2(n19613), .ZN(
        n19598) );
  INV_X1 U22717 ( .A(n19610), .ZN(n19614) );
  AOI22_X1 U22718 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19614), .B1(
        n19952), .B2(n19688), .ZN(n19597) );
  OAI211_X1 U22719 ( .C1(n19607), .C2(n19955), .A(n19598), .B(n19597), .ZN(
        P3_U2877) );
  AOI22_X1 U22720 ( .A1(n19993), .A2(n19883), .B1(n19957), .B2(n19613), .ZN(
        n19600) );
  AOI22_X1 U22721 ( .A1(n19934), .A2(n19956), .B1(n19958), .B2(n19654), .ZN(
        n19599) );
  OAI211_X1 U22722 ( .C1(n19601), .C2(n19610), .A(n19600), .B(n19599), .ZN(
        P3_U2878) );
  INV_X1 U22723 ( .A(n19920), .ZN(n19963) );
  AOI22_X1 U22724 ( .A1(n19934), .A2(n19963), .B1(n19962), .B2(n19613), .ZN(
        n19603) );
  AOI22_X1 U22725 ( .A1(n19993), .A2(n19917), .B1(n19964), .B2(n19654), .ZN(
        n19602) );
  OAI211_X1 U22726 ( .C1(n19604), .C2(n19610), .A(n19603), .B(n19602), .ZN(
        P3_U2879) );
  AOI22_X1 U22727 ( .A1(n19993), .A2(n19921), .B1(n19969), .B2(n19613), .ZN(
        n19606) );
  AOI22_X1 U22728 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19614), .B1(
        n19970), .B2(n19654), .ZN(n19605) );
  OAI211_X1 U22729 ( .C1(n19607), .C2(n19925), .A(n19606), .B(n19605), .ZN(
        P3_U2880) );
  INV_X1 U22730 ( .A(n19981), .ZN(n19926) );
  AOI22_X1 U22731 ( .A1(n19934), .A2(n19926), .B1(n19974), .B2(n19613), .ZN(
        n19609) );
  AOI22_X1 U22732 ( .A1(n19993), .A2(n19975), .B1(n19977), .B2(n19654), .ZN(
        n19608) );
  OAI211_X1 U22733 ( .C1(n21818), .C2(n19610), .A(n19609), .B(n19608), .ZN(
        P3_U2881) );
  INV_X1 U22734 ( .A(n19897), .ZN(n19983) );
  AOI22_X1 U22735 ( .A1(n19934), .A2(n19983), .B1(n19982), .B2(n19613), .ZN(
        n19612) );
  AOI22_X1 U22736 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19614), .B1(
        n19984), .B2(n19654), .ZN(n19611) );
  OAI211_X1 U22737 ( .C1(n19631), .C2(n19987), .A(n19612), .B(n19611), .ZN(
        P3_U2882) );
  AOI22_X1 U22738 ( .A1(n19934), .A2(n19991), .B1(n19989), .B2(n19613), .ZN(
        n19616) );
  AOI22_X1 U22739 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19614), .B1(
        n19992), .B2(n19654), .ZN(n19615) );
  OAI211_X1 U22740 ( .C1(n19631), .C2(n19997), .A(n19616), .B(n19615), .ZN(
        P3_U2883) );
  NOR2_X1 U22741 ( .A1(n11693), .A2(n19643), .ZN(n19694) );
  INV_X1 U22742 ( .A(n19694), .ZN(n19644) );
  NOR2_X2 U22743 ( .A1(n19644), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19711) );
  NOR2_X1 U22744 ( .A1(n19688), .A2(n19711), .ZN(n19671) );
  OAI21_X1 U22745 ( .B1(n19905), .B2(n19617), .A(n19671), .ZN(n19618) );
  OAI211_X1 U22746 ( .C1(n20134), .C2(n19711), .A(n19618), .B(n19908), .ZN(
        n19634) );
  INV_X1 U22747 ( .A(n19634), .ZN(n19641) );
  NOR2_X1 U22748 ( .A1(n19939), .A2(n19671), .ZN(n19637) );
  AOI22_X1 U22749 ( .A1(n19993), .A2(n19940), .B1(n19941), .B2(n19637), .ZN(
        n19620) );
  AOI22_X1 U22750 ( .A1(n19873), .A2(n19666), .B1(n19946), .B2(n19711), .ZN(
        n19619) );
  OAI211_X1 U22751 ( .C1(n19641), .C2(n19621), .A(n19620), .B(n19619), .ZN(
        P3_U2884) );
  AOI22_X1 U22752 ( .A1(n19666), .A2(n19951), .B1(n19950), .B2(n19637), .ZN(
        n19623) );
  AOI22_X1 U22753 ( .A1(n19993), .A2(n19911), .B1(n19952), .B2(n19711), .ZN(
        n19622) );
  OAI211_X1 U22754 ( .C1(n19641), .C2(n19624), .A(n19623), .B(n19622), .ZN(
        P3_U2885) );
  INV_X1 U22755 ( .A(n19666), .ZN(n19664) );
  AOI22_X1 U22756 ( .A1(n19993), .A2(n19956), .B1(n19957), .B2(n19637), .ZN(
        n19626) );
  AOI22_X1 U22757 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19634), .B1(
        n19958), .B2(n19711), .ZN(n19625) );
  OAI211_X1 U22758 ( .C1(n19664), .C2(n19961), .A(n19626), .B(n19625), .ZN(
        P3_U2886) );
  AOI22_X1 U22759 ( .A1(n19666), .A2(n19917), .B1(n19962), .B2(n19637), .ZN(
        n19628) );
  AOI22_X1 U22760 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19634), .B1(
        n19964), .B2(n19711), .ZN(n19627) );
  OAI211_X1 U22761 ( .C1(n19631), .C2(n19920), .A(n19628), .B(n19627), .ZN(
        P3_U2887) );
  AOI22_X1 U22762 ( .A1(n19666), .A2(n19921), .B1(n19969), .B2(n19637), .ZN(
        n19630) );
  AOI22_X1 U22763 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19634), .B1(
        n19970), .B2(n19711), .ZN(n19629) );
  OAI211_X1 U22764 ( .C1(n19631), .C2(n19925), .A(n19630), .B(n19629), .ZN(
        P3_U2888) );
  AOI22_X1 U22765 ( .A1(n19993), .A2(n19926), .B1(n19974), .B2(n19637), .ZN(
        n19633) );
  AOI22_X1 U22766 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19634), .B1(
        n19977), .B2(n19711), .ZN(n19632) );
  OAI211_X1 U22767 ( .C1(n19664), .C2(n19929), .A(n19633), .B(n19632), .ZN(
        P3_U2889) );
  AOI22_X1 U22768 ( .A1(n19993), .A2(n19983), .B1(n19982), .B2(n19637), .ZN(
        n19636) );
  AOI22_X1 U22769 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19634), .B1(
        n19984), .B2(n19711), .ZN(n19635) );
  OAI211_X1 U22770 ( .C1(n19664), .C2(n19987), .A(n19636), .B(n19635), .ZN(
        P3_U2890) );
  AOI22_X1 U22771 ( .A1(n19666), .A2(n19898), .B1(n19989), .B2(n19637), .ZN(
        n19639) );
  AOI22_X1 U22772 ( .A1(n19993), .A2(n19991), .B1(n19992), .B2(n19711), .ZN(
        n19638) );
  OAI211_X1 U22773 ( .C1(n19641), .C2(n19640), .A(n19639), .B(n19638), .ZN(
        P3_U2891) );
  OAI21_X1 U22774 ( .B1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n19642), .A(
        n19942), .ZN(n19738) );
  NOR2_X1 U22775 ( .A1(n19643), .A2(n19738), .ZN(n19670) );
  NOR2_X1 U22776 ( .A1(n19939), .A2(n19644), .ZN(n19665) );
  AOI22_X1 U22777 ( .A1(n19666), .A2(n19940), .B1(n19941), .B2(n19665), .ZN(
        n19646) );
  NAND2_X1 U22778 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19694), .ZN(
        n19732) );
  AOI22_X1 U22779 ( .A1(n19873), .A2(n19688), .B1(n19946), .B2(n19734), .ZN(
        n19645) );
  OAI211_X1 U22780 ( .C1(n19670), .C2(n19647), .A(n19646), .B(n19645), .ZN(
        P3_U2892) );
  INV_X1 U22781 ( .A(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n19650) );
  AOI22_X1 U22782 ( .A1(n19666), .A2(n19911), .B1(n19950), .B2(n19665), .ZN(
        n19649) );
  AOI22_X1 U22783 ( .A1(n19952), .A2(n19734), .B1(n19951), .B2(n19654), .ZN(
        n19648) );
  OAI211_X1 U22784 ( .C1(n19670), .C2(n19650), .A(n19649), .B(n19648), .ZN(
        P3_U2893) );
  INV_X1 U22785 ( .A(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n19653) );
  AOI22_X1 U22786 ( .A1(n19883), .A2(n19688), .B1(n19957), .B2(n19665), .ZN(
        n19652) );
  AOI22_X1 U22787 ( .A1(n19666), .A2(n19956), .B1(n19958), .B2(n19734), .ZN(
        n19651) );
  OAI211_X1 U22788 ( .C1(n19670), .C2(n19653), .A(n19652), .B(n19651), .ZN(
        P3_U2894) );
  INV_X1 U22789 ( .A(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n21896) );
  AOI22_X1 U22790 ( .A1(n19666), .A2(n19963), .B1(n19962), .B2(n19665), .ZN(
        n19656) );
  AOI22_X1 U22791 ( .A1(n19964), .A2(n19734), .B1(n19917), .B2(n19654), .ZN(
        n19655) );
  OAI211_X1 U22792 ( .C1(n19670), .C2(n21896), .A(n19656), .B(n19655), .ZN(
        P3_U2895) );
  AOI22_X1 U22793 ( .A1(n19921), .A2(n19688), .B1(n19969), .B2(n19665), .ZN(
        n19658) );
  INV_X1 U22794 ( .A(n19670), .ZN(n19661) );
  AOI22_X1 U22795 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19661), .B1(
        n19970), .B2(n19734), .ZN(n19657) );
  OAI211_X1 U22796 ( .C1(n19664), .C2(n19925), .A(n19658), .B(n19657), .ZN(
        P3_U2896) );
  AOI22_X1 U22797 ( .A1(n19975), .A2(n19688), .B1(n19974), .B2(n19665), .ZN(
        n19660) );
  AOI22_X1 U22798 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19661), .B1(
        n19977), .B2(n19734), .ZN(n19659) );
  OAI211_X1 U22799 ( .C1(n19664), .C2(n19981), .A(n19660), .B(n19659), .ZN(
        P3_U2897) );
  AOI22_X1 U22800 ( .A1(n19894), .A2(n19688), .B1(n19982), .B2(n19665), .ZN(
        n19663) );
  AOI22_X1 U22801 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19661), .B1(
        n19984), .B2(n19734), .ZN(n19662) );
  OAI211_X1 U22802 ( .C1(n19664), .C2(n19897), .A(n19663), .B(n19662), .ZN(
        P3_U2898) );
  AOI22_X1 U22803 ( .A1(n19898), .A2(n19688), .B1(n19989), .B2(n19665), .ZN(
        n19668) );
  AOI22_X1 U22804 ( .A1(n19666), .A2(n19991), .B1(n19992), .B2(n19734), .ZN(
        n19667) );
  OAI211_X1 U22805 ( .C1(n19670), .C2(n19669), .A(n19668), .B(n19667), .ZN(
        P3_U2899) );
  NOR2_X2 U22806 ( .A1(n20005), .A2(n19739), .ZN(n19752) );
  NOR2_X1 U22807 ( .A1(n19734), .A2(n19752), .ZN(n19716) );
  NOR2_X1 U22808 ( .A1(n19939), .A2(n19716), .ZN(n19687) );
  AOI22_X1 U22809 ( .A1(n19941), .A2(n19687), .B1(n19940), .B2(n19688), .ZN(
        n19674) );
  OAI21_X1 U22810 ( .B1(n19671), .B2(n19905), .A(n19716), .ZN(n19672) );
  OAI211_X1 U22811 ( .C1(n19752), .C2(n20134), .A(n19908), .B(n19672), .ZN(
        n19689) );
  AOI22_X1 U22812 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19689), .B1(
        n19946), .B2(n19752), .ZN(n19673) );
  OAI211_X1 U22813 ( .C1(n19949), .C2(n19709), .A(n19674), .B(n19673), .ZN(
        P3_U2900) );
  AOI22_X1 U22814 ( .A1(n19911), .A2(n19688), .B1(n19950), .B2(n19687), .ZN(
        n19676) );
  AOI22_X1 U22815 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19689), .B1(
        n19952), .B2(n19752), .ZN(n19675) );
  OAI211_X1 U22816 ( .C1(n19914), .C2(n19709), .A(n19676), .B(n19675), .ZN(
        P3_U2901) );
  AOI22_X1 U22817 ( .A1(n19957), .A2(n19687), .B1(n19956), .B2(n19688), .ZN(
        n19678) );
  AOI22_X1 U22818 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19689), .B1(
        n19958), .B2(n19752), .ZN(n19677) );
  OAI211_X1 U22819 ( .C1(n19961), .C2(n19709), .A(n19678), .B(n19677), .ZN(
        P3_U2902) );
  AOI22_X1 U22820 ( .A1(n19963), .A2(n19688), .B1(n19962), .B2(n19687), .ZN(
        n19680) );
  AOI22_X1 U22821 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19689), .B1(
        n19964), .B2(n19752), .ZN(n19679) );
  OAI211_X1 U22822 ( .C1(n19967), .C2(n19709), .A(n19680), .B(n19679), .ZN(
        P3_U2903) );
  AOI22_X1 U22823 ( .A1(n19969), .A2(n19687), .B1(n19968), .B2(n19688), .ZN(
        n19682) );
  AOI22_X1 U22824 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19689), .B1(
        n19970), .B2(n19752), .ZN(n19681) );
  OAI211_X1 U22825 ( .C1(n19973), .C2(n19709), .A(n19682), .B(n19681), .ZN(
        P3_U2904) );
  AOI22_X1 U22826 ( .A1(n19926), .A2(n19688), .B1(n19974), .B2(n19687), .ZN(
        n19684) );
  AOI22_X1 U22827 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19689), .B1(
        n19977), .B2(n19752), .ZN(n19683) );
  OAI211_X1 U22828 ( .C1(n19929), .C2(n19709), .A(n19684), .B(n19683), .ZN(
        P3_U2905) );
  AOI22_X1 U22829 ( .A1(n19983), .A2(n19688), .B1(n19982), .B2(n19687), .ZN(
        n19686) );
  AOI22_X1 U22830 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19689), .B1(
        n19984), .B2(n19752), .ZN(n19685) );
  OAI211_X1 U22831 ( .C1(n19987), .C2(n19709), .A(n19686), .B(n19685), .ZN(
        P3_U2906) );
  AOI22_X1 U22832 ( .A1(n19991), .A2(n19688), .B1(n19989), .B2(n19687), .ZN(
        n19691) );
  AOI22_X1 U22833 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19689), .B1(
        n19992), .B2(n19752), .ZN(n19690) );
  OAI211_X1 U22834 ( .C1(n19997), .C2(n19709), .A(n19691), .B(n19690), .ZN(
        P3_U2907) );
  NOR2_X1 U22835 ( .A1(n19739), .A2(n19871), .ZN(n19710) );
  AOI22_X1 U22836 ( .A1(n19873), .A2(n19734), .B1(n19941), .B2(n19710), .ZN(
        n19696) );
  INV_X1 U22837 ( .A(n19692), .ZN(n19874) );
  AOI22_X1 U22838 ( .A1(n19877), .A2(n19694), .B1(n19693), .B2(n19874), .ZN(
        n19712) );
  NOR2_X2 U22839 ( .A1(n19739), .A2(n19784), .ZN(n19772) );
  AOI22_X1 U22840 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19712), .B1(
        n19946), .B2(n19772), .ZN(n19695) );
  OAI211_X1 U22841 ( .C1(n19880), .C2(n19709), .A(n19696), .B(n19695), .ZN(
        P3_U2908) );
  AOI22_X1 U22842 ( .A1(n19951), .A2(n19734), .B1(n19950), .B2(n19710), .ZN(
        n19698) );
  AOI22_X1 U22843 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19712), .B1(
        n19952), .B2(n19772), .ZN(n19697) );
  OAI211_X1 U22844 ( .C1(n19955), .C2(n19709), .A(n19698), .B(n19697), .ZN(
        P3_U2909) );
  AOI22_X1 U22845 ( .A1(n19957), .A2(n19710), .B1(n19956), .B2(n19711), .ZN(
        n19700) );
  AOI22_X1 U22846 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19712), .B1(
        n19958), .B2(n19772), .ZN(n19699) );
  OAI211_X1 U22847 ( .C1(n19961), .C2(n19732), .A(n19700), .B(n19699), .ZN(
        P3_U2910) );
  AOI22_X1 U22848 ( .A1(n19963), .A2(n19711), .B1(n19962), .B2(n19710), .ZN(
        n19702) );
  AOI22_X1 U22849 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19712), .B1(
        n19964), .B2(n19772), .ZN(n19701) );
  OAI211_X1 U22850 ( .C1(n19967), .C2(n19732), .A(n19702), .B(n19701), .ZN(
        P3_U2911) );
  AOI22_X1 U22851 ( .A1(n19921), .A2(n19734), .B1(n19969), .B2(n19710), .ZN(
        n19704) );
  AOI22_X1 U22852 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19712), .B1(
        n19970), .B2(n19772), .ZN(n19703) );
  OAI211_X1 U22853 ( .C1(n19925), .C2(n19709), .A(n19704), .B(n19703), .ZN(
        P3_U2912) );
  AOI22_X1 U22854 ( .A1(n19975), .A2(n19734), .B1(n19974), .B2(n19710), .ZN(
        n19706) );
  AOI22_X1 U22855 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19712), .B1(
        n19977), .B2(n19772), .ZN(n19705) );
  OAI211_X1 U22856 ( .C1(n19981), .C2(n19709), .A(n19706), .B(n19705), .ZN(
        P3_U2913) );
  AOI22_X1 U22857 ( .A1(n19894), .A2(n19734), .B1(n19982), .B2(n19710), .ZN(
        n19708) );
  AOI22_X1 U22858 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19712), .B1(
        n19984), .B2(n19772), .ZN(n19707) );
  OAI211_X1 U22859 ( .C1(n19897), .C2(n19709), .A(n19708), .B(n19707), .ZN(
        P3_U2914) );
  AOI22_X1 U22860 ( .A1(n19991), .A2(n19711), .B1(n19989), .B2(n19710), .ZN(
        n19714) );
  AOI22_X1 U22861 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19712), .B1(
        n19992), .B2(n19772), .ZN(n19713) );
  OAI211_X1 U22862 ( .C1(n19997), .C2(n19732), .A(n19714), .B(n19713), .ZN(
        P3_U2915) );
  INV_X1 U22863 ( .A(n19752), .ZN(n19759) );
  NOR2_X1 U22864 ( .A1(n19715), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19783) );
  NAND2_X1 U22865 ( .A1(n11692), .A2(n19783), .ZN(n19803) );
  INV_X1 U22866 ( .A(n19803), .ZN(n19795) );
  NOR2_X1 U22867 ( .A1(n19772), .A2(n19795), .ZN(n19760) );
  NOR2_X1 U22868 ( .A1(n19939), .A2(n19760), .ZN(n19733) );
  AOI22_X1 U22869 ( .A1(n19941), .A2(n19733), .B1(n19940), .B2(n19734), .ZN(
        n19719) );
  OAI21_X1 U22870 ( .B1(n19716), .B2(n19905), .A(n19760), .ZN(n19717) );
  OAI211_X1 U22871 ( .C1(n19795), .C2(n20134), .A(n19908), .B(n19717), .ZN(
        n19735) );
  AOI22_X1 U22872 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19735), .B1(
        n19946), .B2(n19795), .ZN(n19718) );
  OAI211_X1 U22873 ( .C1(n19949), .C2(n19759), .A(n19719), .B(n19718), .ZN(
        P3_U2916) );
  AOI22_X1 U22874 ( .A1(n19951), .A2(n19752), .B1(n19950), .B2(n19733), .ZN(
        n19721) );
  AOI22_X1 U22875 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19735), .B1(
        n19952), .B2(n19795), .ZN(n19720) );
  OAI211_X1 U22876 ( .C1(n19955), .C2(n19732), .A(n19721), .B(n19720), .ZN(
        P3_U2917) );
  AOI22_X1 U22877 ( .A1(n19957), .A2(n19733), .B1(n19956), .B2(n19734), .ZN(
        n19723) );
  AOI22_X1 U22878 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19735), .B1(
        n19958), .B2(n19795), .ZN(n19722) );
  OAI211_X1 U22879 ( .C1(n19961), .C2(n19759), .A(n19723), .B(n19722), .ZN(
        P3_U2918) );
  AOI22_X1 U22880 ( .A1(n19963), .A2(n19734), .B1(n19962), .B2(n19733), .ZN(
        n19725) );
  AOI22_X1 U22881 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19735), .B1(
        n19964), .B2(n19795), .ZN(n19724) );
  OAI211_X1 U22882 ( .C1(n19967), .C2(n19759), .A(n19725), .B(n19724), .ZN(
        P3_U2919) );
  AOI22_X1 U22883 ( .A1(n19921), .A2(n19752), .B1(n19969), .B2(n19733), .ZN(
        n19727) );
  AOI22_X1 U22884 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19735), .B1(
        n19970), .B2(n19795), .ZN(n19726) );
  OAI211_X1 U22885 ( .C1(n19925), .C2(n19732), .A(n19727), .B(n19726), .ZN(
        P3_U2920) );
  AOI22_X1 U22886 ( .A1(n19975), .A2(n19752), .B1(n19974), .B2(n19733), .ZN(
        n19729) );
  AOI22_X1 U22887 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19735), .B1(
        n19977), .B2(n19795), .ZN(n19728) );
  OAI211_X1 U22888 ( .C1(n19981), .C2(n19732), .A(n19729), .B(n19728), .ZN(
        P3_U2921) );
  AOI22_X1 U22889 ( .A1(n19894), .A2(n19752), .B1(n19982), .B2(n19733), .ZN(
        n19731) );
  AOI22_X1 U22890 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19735), .B1(
        n19984), .B2(n19795), .ZN(n19730) );
  OAI211_X1 U22891 ( .C1(n19897), .C2(n19732), .A(n19731), .B(n19730), .ZN(
        P3_U2922) );
  AOI22_X1 U22892 ( .A1(n19991), .A2(n19734), .B1(n19989), .B2(n19733), .ZN(
        n19737) );
  AOI22_X1 U22893 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19735), .B1(
        n19992), .B2(n19795), .ZN(n19736) );
  OAI211_X1 U22894 ( .C1(n19997), .C2(n19759), .A(n19737), .B(n19736), .ZN(
        P3_U2923) );
  AND2_X1 U22895 ( .A1(n19827), .A2(n19783), .ZN(n19755) );
  AOI22_X1 U22896 ( .A1(n19873), .A2(n19772), .B1(n19941), .B2(n19755), .ZN(
        n19741) );
  OR2_X1 U22897 ( .A1(n19739), .A2(n19738), .ZN(n19756) );
  NAND2_X1 U22898 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19783), .ZN(
        n19826) );
  AOI22_X1 U22899 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19756), .B1(
        n19946), .B2(n19819), .ZN(n19740) );
  OAI211_X1 U22900 ( .C1(n19880), .C2(n19759), .A(n19741), .B(n19740), .ZN(
        P3_U2924) );
  INV_X1 U22901 ( .A(n19772), .ZN(n19781) );
  AOI22_X1 U22902 ( .A1(n19911), .A2(n19752), .B1(n19950), .B2(n19755), .ZN(
        n19743) );
  AOI22_X1 U22903 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19756), .B1(
        n19952), .B2(n19819), .ZN(n19742) );
  OAI211_X1 U22904 ( .C1(n19914), .C2(n19781), .A(n19743), .B(n19742), .ZN(
        P3_U2925) );
  AOI22_X1 U22905 ( .A1(n19957), .A2(n19755), .B1(n19956), .B2(n19752), .ZN(
        n19745) );
  AOI22_X1 U22906 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19756), .B1(
        n19958), .B2(n19819), .ZN(n19744) );
  OAI211_X1 U22907 ( .C1(n19961), .C2(n19781), .A(n19745), .B(n19744), .ZN(
        P3_U2926) );
  AOI22_X1 U22908 ( .A1(n19963), .A2(n19752), .B1(n19962), .B2(n19755), .ZN(
        n19747) );
  AOI22_X1 U22909 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19756), .B1(
        n19964), .B2(n19819), .ZN(n19746) );
  OAI211_X1 U22910 ( .C1(n19967), .C2(n19781), .A(n19747), .B(n19746), .ZN(
        P3_U2927) );
  AOI22_X1 U22911 ( .A1(n19921), .A2(n19772), .B1(n19969), .B2(n19755), .ZN(
        n19749) );
  AOI22_X1 U22912 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19756), .B1(
        n19970), .B2(n19819), .ZN(n19748) );
  OAI211_X1 U22913 ( .C1(n19925), .C2(n19759), .A(n19749), .B(n19748), .ZN(
        P3_U2928) );
  AOI22_X1 U22914 ( .A1(n19926), .A2(n19752), .B1(n19974), .B2(n19755), .ZN(
        n19751) );
  AOI22_X1 U22915 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19756), .B1(
        n19977), .B2(n19819), .ZN(n19750) );
  OAI211_X1 U22916 ( .C1(n19929), .C2(n19781), .A(n19751), .B(n19750), .ZN(
        P3_U2929) );
  AOI22_X1 U22917 ( .A1(n19983), .A2(n19752), .B1(n19982), .B2(n19755), .ZN(
        n19754) );
  AOI22_X1 U22918 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19756), .B1(
        n19984), .B2(n19819), .ZN(n19753) );
  OAI211_X1 U22919 ( .C1(n19987), .C2(n19781), .A(n19754), .B(n19753), .ZN(
        P3_U2930) );
  AOI22_X1 U22920 ( .A1(n19898), .A2(n19772), .B1(n19989), .B2(n19755), .ZN(
        n19758) );
  AOI22_X1 U22921 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19756), .B1(
        n19992), .B2(n19819), .ZN(n19757) );
  OAI211_X1 U22922 ( .C1(n19903), .C2(n19759), .A(n19758), .B(n19757), .ZN(
        P3_U2931) );
  NOR2_X2 U22923 ( .A1(n20005), .A2(n19804), .ZN(n19845) );
  NOR2_X1 U22924 ( .A1(n19819), .A2(n19845), .ZN(n19805) );
  NOR2_X1 U22925 ( .A1(n19939), .A2(n19805), .ZN(n19777) );
  AOI22_X1 U22926 ( .A1(n19941), .A2(n19777), .B1(n19940), .B2(n19772), .ZN(
        n19763) );
  OAI21_X1 U22927 ( .B1(n19760), .B2(n19905), .A(n19805), .ZN(n19761) );
  OAI211_X1 U22928 ( .C1(n19845), .C2(n20134), .A(n19908), .B(n19761), .ZN(
        n19778) );
  AOI22_X1 U22929 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19778), .B1(
        n19946), .B2(n19845), .ZN(n19762) );
  OAI211_X1 U22930 ( .C1(n19949), .C2(n19803), .A(n19763), .B(n19762), .ZN(
        P3_U2932) );
  AOI22_X1 U22931 ( .A1(n19951), .A2(n19795), .B1(n19950), .B2(n19777), .ZN(
        n19765) );
  AOI22_X1 U22932 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19778), .B1(
        n19952), .B2(n19845), .ZN(n19764) );
  OAI211_X1 U22933 ( .C1(n19955), .C2(n19781), .A(n19765), .B(n19764), .ZN(
        P3_U2933) );
  AOI22_X1 U22934 ( .A1(n19957), .A2(n19777), .B1(n19956), .B2(n19772), .ZN(
        n19767) );
  AOI22_X1 U22935 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19778), .B1(
        n19958), .B2(n19845), .ZN(n19766) );
  OAI211_X1 U22936 ( .C1(n19961), .C2(n19803), .A(n19767), .B(n19766), .ZN(
        P3_U2934) );
  AOI22_X1 U22937 ( .A1(n19917), .A2(n19795), .B1(n19962), .B2(n19777), .ZN(
        n19769) );
  AOI22_X1 U22938 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19778), .B1(
        n19964), .B2(n19845), .ZN(n19768) );
  OAI211_X1 U22939 ( .C1(n19920), .C2(n19781), .A(n19769), .B(n19768), .ZN(
        P3_U2935) );
  AOI22_X1 U22940 ( .A1(n19969), .A2(n19777), .B1(n19968), .B2(n19772), .ZN(
        n19771) );
  AOI22_X1 U22941 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19778), .B1(
        n19970), .B2(n19845), .ZN(n19770) );
  OAI211_X1 U22942 ( .C1(n19973), .C2(n19803), .A(n19771), .B(n19770), .ZN(
        P3_U2936) );
  AOI22_X1 U22943 ( .A1(n19926), .A2(n19772), .B1(n19974), .B2(n19777), .ZN(
        n19774) );
  AOI22_X1 U22944 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19778), .B1(
        n19977), .B2(n19845), .ZN(n19773) );
  OAI211_X1 U22945 ( .C1(n19929), .C2(n19803), .A(n19774), .B(n19773), .ZN(
        P3_U2937) );
  AOI22_X1 U22946 ( .A1(n19894), .A2(n19795), .B1(n19982), .B2(n19777), .ZN(
        n19776) );
  AOI22_X1 U22947 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19778), .B1(
        n19984), .B2(n19845), .ZN(n19775) );
  OAI211_X1 U22948 ( .C1(n19897), .C2(n19781), .A(n19776), .B(n19775), .ZN(
        P3_U2938) );
  AOI22_X1 U22949 ( .A1(n19898), .A2(n19795), .B1(n19989), .B2(n19777), .ZN(
        n19780) );
  AOI22_X1 U22950 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19778), .B1(
        n19992), .B2(n19845), .ZN(n19779) );
  OAI211_X1 U22951 ( .C1(n19903), .C2(n19781), .A(n19780), .B(n19779), .ZN(
        P3_U2939) );
  NOR2_X1 U22952 ( .A1(n19804), .A2(n19871), .ZN(n19828) );
  AOI22_X1 U22953 ( .A1(n19941), .A2(n19828), .B1(n19940), .B2(n19795), .ZN(
        n19786) );
  AOI22_X1 U22954 ( .A1(n19877), .A2(n19783), .B1(n19782), .B2(n19874), .ZN(
        n19800) );
  NOR2_X2 U22955 ( .A1(n19804), .A2(n19784), .ZN(n19861) );
  AOI22_X1 U22956 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19800), .B1(
        n19946), .B2(n19861), .ZN(n19785) );
  OAI211_X1 U22957 ( .C1(n19949), .C2(n19826), .A(n19786), .B(n19785), .ZN(
        P3_U2940) );
  AOI22_X1 U22958 ( .A1(n19951), .A2(n19819), .B1(n19950), .B2(n19828), .ZN(
        n19788) );
  AOI22_X1 U22959 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19800), .B1(
        n19952), .B2(n19861), .ZN(n19787) );
  OAI211_X1 U22960 ( .C1(n19955), .C2(n19803), .A(n19788), .B(n19787), .ZN(
        P3_U2941) );
  AOI22_X1 U22961 ( .A1(n19883), .A2(n19819), .B1(n19957), .B2(n19828), .ZN(
        n19790) );
  AOI22_X1 U22962 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19800), .B1(
        n19958), .B2(n19861), .ZN(n19789) );
  OAI211_X1 U22963 ( .C1(n19886), .C2(n19803), .A(n19790), .B(n19789), .ZN(
        P3_U2942) );
  AOI22_X1 U22964 ( .A1(n19917), .A2(n19819), .B1(n19962), .B2(n19828), .ZN(
        n19792) );
  AOI22_X1 U22965 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19800), .B1(
        n19964), .B2(n19861), .ZN(n19791) );
  OAI211_X1 U22966 ( .C1(n19920), .C2(n19803), .A(n19792), .B(n19791), .ZN(
        P3_U2943) );
  AOI22_X1 U22967 ( .A1(n19969), .A2(n19828), .B1(n19968), .B2(n19795), .ZN(
        n19794) );
  AOI22_X1 U22968 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19800), .B1(
        n19970), .B2(n19861), .ZN(n19793) );
  OAI211_X1 U22969 ( .C1(n19973), .C2(n19826), .A(n19794), .B(n19793), .ZN(
        P3_U2944) );
  AOI22_X1 U22970 ( .A1(n19926), .A2(n19795), .B1(n19974), .B2(n19828), .ZN(
        n19797) );
  AOI22_X1 U22971 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19800), .B1(
        n19977), .B2(n19861), .ZN(n19796) );
  OAI211_X1 U22972 ( .C1(n19929), .C2(n19826), .A(n19797), .B(n19796), .ZN(
        P3_U2945) );
  AOI22_X1 U22973 ( .A1(n19894), .A2(n19819), .B1(n19982), .B2(n19828), .ZN(
        n19799) );
  AOI22_X1 U22974 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19800), .B1(
        n19984), .B2(n19861), .ZN(n19798) );
  OAI211_X1 U22975 ( .C1(n19897), .C2(n19803), .A(n19799), .B(n19798), .ZN(
        P3_U2946) );
  AOI22_X1 U22976 ( .A1(n19898), .A2(n19819), .B1(n19989), .B2(n19828), .ZN(
        n19802) );
  AOI22_X1 U22977 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19800), .B1(
        n19992), .B2(n19861), .ZN(n19801) );
  OAI211_X1 U22978 ( .C1(n19903), .C2(n19803), .A(n19802), .B(n19801), .ZN(
        P3_U2947) );
  INV_X1 U22979 ( .A(n19845), .ZN(n19835) );
  NOR2_X1 U22980 ( .A1(n11693), .A2(n19804), .ZN(n19876) );
  NAND2_X1 U22981 ( .A1(n11692), .A2(n19876), .ZN(n19902) );
  INV_X1 U22982 ( .A(n19902), .ZN(n19889) );
  NOR2_X1 U22983 ( .A1(n19861), .A2(n19889), .ZN(n19849) );
  NOR2_X1 U22984 ( .A1(n19939), .A2(n19849), .ZN(n19822) );
  AOI22_X1 U22985 ( .A1(n19941), .A2(n19822), .B1(n19940), .B2(n19819), .ZN(
        n19808) );
  OAI21_X1 U22986 ( .B1(n19805), .B2(n19905), .A(n19849), .ZN(n19806) );
  OAI211_X1 U22987 ( .C1(n19889), .C2(n20134), .A(n19908), .B(n19806), .ZN(
        n19823) );
  AOI22_X1 U22988 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19823), .B1(
        n19946), .B2(n19889), .ZN(n19807) );
  OAI211_X1 U22989 ( .C1(n19949), .C2(n19835), .A(n19808), .B(n19807), .ZN(
        P3_U2948) );
  AOI22_X1 U22990 ( .A1(n19911), .A2(n19819), .B1(n19950), .B2(n19822), .ZN(
        n19810) );
  AOI22_X1 U22991 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19823), .B1(
        n19952), .B2(n19889), .ZN(n19809) );
  OAI211_X1 U22992 ( .C1(n19914), .C2(n19835), .A(n19810), .B(n19809), .ZN(
        P3_U2949) );
  AOI22_X1 U22993 ( .A1(n19957), .A2(n19822), .B1(n19956), .B2(n19819), .ZN(
        n19812) );
  AOI22_X1 U22994 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19823), .B1(
        n19958), .B2(n19889), .ZN(n19811) );
  OAI211_X1 U22995 ( .C1(n19961), .C2(n19835), .A(n19812), .B(n19811), .ZN(
        P3_U2950) );
  AOI22_X1 U22996 ( .A1(n19963), .A2(n19819), .B1(n19962), .B2(n19822), .ZN(
        n19814) );
  AOI22_X1 U22997 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19823), .B1(
        n19964), .B2(n19889), .ZN(n19813) );
  OAI211_X1 U22998 ( .C1(n19967), .C2(n19835), .A(n19814), .B(n19813), .ZN(
        P3_U2951) );
  AOI22_X1 U22999 ( .A1(n19921), .A2(n19845), .B1(n19969), .B2(n19822), .ZN(
        n19816) );
  AOI22_X1 U23000 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19823), .B1(
        n19970), .B2(n19889), .ZN(n19815) );
  OAI211_X1 U23001 ( .C1(n19925), .C2(n19826), .A(n19816), .B(n19815), .ZN(
        P3_U2952) );
  AOI22_X1 U23002 ( .A1(n19926), .A2(n19819), .B1(n19974), .B2(n19822), .ZN(
        n19818) );
  AOI22_X1 U23003 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19823), .B1(
        n19977), .B2(n19889), .ZN(n19817) );
  OAI211_X1 U23004 ( .C1(n19929), .C2(n19835), .A(n19818), .B(n19817), .ZN(
        P3_U2953) );
  AOI22_X1 U23005 ( .A1(n19983), .A2(n19819), .B1(n19982), .B2(n19822), .ZN(
        n19821) );
  AOI22_X1 U23006 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19823), .B1(
        n19984), .B2(n19889), .ZN(n19820) );
  OAI211_X1 U23007 ( .C1(n19987), .C2(n19835), .A(n19821), .B(n19820), .ZN(
        P3_U2954) );
  AOI22_X1 U23008 ( .A1(n19898), .A2(n19845), .B1(n19989), .B2(n19822), .ZN(
        n19825) );
  AOI22_X1 U23009 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19823), .B1(
        n19992), .B2(n19889), .ZN(n19824) );
  OAI211_X1 U23010 ( .C1(n19903), .C2(n19826), .A(n19825), .B(n19824), .ZN(
        P3_U2955) );
  INV_X1 U23011 ( .A(n19861), .ZN(n19870) );
  AND2_X1 U23012 ( .A1(n19827), .A2(n19876), .ZN(n19844) );
  AOI22_X1 U23013 ( .A1(n19941), .A2(n19844), .B1(n19940), .B2(n19845), .ZN(
        n19830) );
  AOI22_X1 U23014 ( .A1(n19877), .A2(n19828), .B1(n19942), .B2(n19876), .ZN(
        n19846) );
  NAND2_X1 U23015 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19876), .ZN(
        n19924) );
  INV_X1 U23016 ( .A(n19924), .ZN(n19933) );
  AOI22_X1 U23017 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19846), .B1(
        n19946), .B2(n19933), .ZN(n19829) );
  OAI211_X1 U23018 ( .C1(n19949), .C2(n19870), .A(n19830), .B(n19829), .ZN(
        P3_U2956) );
  AOI22_X1 U23019 ( .A1(n19911), .A2(n19845), .B1(n19950), .B2(n19844), .ZN(
        n19832) );
  AOI22_X1 U23020 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19846), .B1(
        n19952), .B2(n19933), .ZN(n19831) );
  OAI211_X1 U23021 ( .C1(n19914), .C2(n19870), .A(n19832), .B(n19831), .ZN(
        P3_U2957) );
  AOI22_X1 U23022 ( .A1(n19883), .A2(n19861), .B1(n19957), .B2(n19844), .ZN(
        n19834) );
  AOI22_X1 U23023 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19846), .B1(
        n19958), .B2(n19933), .ZN(n19833) );
  OAI211_X1 U23024 ( .C1(n19886), .C2(n19835), .A(n19834), .B(n19833), .ZN(
        P3_U2958) );
  AOI22_X1 U23025 ( .A1(n19963), .A2(n19845), .B1(n19962), .B2(n19844), .ZN(
        n19837) );
  AOI22_X1 U23026 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19846), .B1(
        n19964), .B2(n19933), .ZN(n19836) );
  OAI211_X1 U23027 ( .C1(n19967), .C2(n19870), .A(n19837), .B(n19836), .ZN(
        P3_U2959) );
  AOI22_X1 U23028 ( .A1(n19969), .A2(n19844), .B1(n19968), .B2(n19845), .ZN(
        n19839) );
  AOI22_X1 U23029 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19846), .B1(
        n19970), .B2(n19933), .ZN(n19838) );
  OAI211_X1 U23030 ( .C1(n19973), .C2(n19870), .A(n19839), .B(n19838), .ZN(
        P3_U2960) );
  AOI22_X1 U23031 ( .A1(n19926), .A2(n19845), .B1(n19974), .B2(n19844), .ZN(
        n19841) );
  AOI22_X1 U23032 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19846), .B1(
        n19977), .B2(n19933), .ZN(n19840) );
  OAI211_X1 U23033 ( .C1(n19929), .C2(n19870), .A(n19841), .B(n19840), .ZN(
        P3_U2961) );
  AOI22_X1 U23034 ( .A1(n19983), .A2(n19845), .B1(n19982), .B2(n19844), .ZN(
        n19843) );
  AOI22_X1 U23035 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19846), .B1(
        n19984), .B2(n19933), .ZN(n19842) );
  OAI211_X1 U23036 ( .C1(n19987), .C2(n19870), .A(n19843), .B(n19842), .ZN(
        P3_U2962) );
  AOI22_X1 U23037 ( .A1(n19991), .A2(n19845), .B1(n19989), .B2(n19844), .ZN(
        n19848) );
  AOI22_X1 U23038 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19846), .B1(
        n19992), .B2(n19933), .ZN(n19847) );
  OAI211_X1 U23039 ( .C1(n19997), .C2(n19870), .A(n19848), .B(n19847), .ZN(
        P3_U2963) );
  NOR2_X2 U23040 ( .A1(n20005), .A2(n19872), .ZN(n19990) );
  NOR2_X1 U23041 ( .A1(n19933), .A2(n19990), .ZN(n19906) );
  NOR2_X1 U23042 ( .A1(n19939), .A2(n19906), .ZN(n19866) );
  AOI22_X1 U23043 ( .A1(n19941), .A2(n19866), .B1(n19940), .B2(n19861), .ZN(
        n19852) );
  OAI21_X1 U23044 ( .B1(n19849), .B2(n19905), .A(n19906), .ZN(n19850) );
  OAI211_X1 U23045 ( .C1(n19990), .C2(n20134), .A(n19908), .B(n19850), .ZN(
        n19867) );
  AOI22_X1 U23046 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19867), .B1(
        n19946), .B2(n19990), .ZN(n19851) );
  OAI211_X1 U23047 ( .C1(n19949), .C2(n19902), .A(n19852), .B(n19851), .ZN(
        P3_U2964) );
  AOI22_X1 U23048 ( .A1(n19951), .A2(n19889), .B1(n19950), .B2(n19866), .ZN(
        n19854) );
  AOI22_X1 U23049 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19867), .B1(
        n19952), .B2(n19990), .ZN(n19853) );
  OAI211_X1 U23050 ( .C1(n19955), .C2(n19870), .A(n19854), .B(n19853), .ZN(
        P3_U2965) );
  AOI22_X1 U23051 ( .A1(n19957), .A2(n19866), .B1(n19956), .B2(n19861), .ZN(
        n19856) );
  AOI22_X1 U23052 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19867), .B1(
        n19958), .B2(n19990), .ZN(n19855) );
  OAI211_X1 U23053 ( .C1(n19961), .C2(n19902), .A(n19856), .B(n19855), .ZN(
        P3_U2966) );
  AOI22_X1 U23054 ( .A1(n19917), .A2(n19889), .B1(n19962), .B2(n19866), .ZN(
        n19858) );
  AOI22_X1 U23055 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19867), .B1(
        n19964), .B2(n19990), .ZN(n19857) );
  OAI211_X1 U23056 ( .C1(n19920), .C2(n19870), .A(n19858), .B(n19857), .ZN(
        P3_U2967) );
  AOI22_X1 U23057 ( .A1(n19969), .A2(n19866), .B1(n19968), .B2(n19861), .ZN(
        n19860) );
  AOI22_X1 U23058 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19867), .B1(
        n19970), .B2(n19990), .ZN(n19859) );
  OAI211_X1 U23059 ( .C1(n19973), .C2(n19902), .A(n19860), .B(n19859), .ZN(
        P3_U2968) );
  AOI22_X1 U23060 ( .A1(n19926), .A2(n19861), .B1(n19974), .B2(n19866), .ZN(
        n19863) );
  AOI22_X1 U23061 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19867), .B1(
        n19977), .B2(n19990), .ZN(n19862) );
  OAI211_X1 U23062 ( .C1(n19929), .C2(n19902), .A(n19863), .B(n19862), .ZN(
        P3_U2969) );
  AOI22_X1 U23063 ( .A1(n19894), .A2(n19889), .B1(n19982), .B2(n19866), .ZN(
        n19865) );
  AOI22_X1 U23064 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19867), .B1(
        n19984), .B2(n19990), .ZN(n19864) );
  OAI211_X1 U23065 ( .C1(n19897), .C2(n19870), .A(n19865), .B(n19864), .ZN(
        P3_U2970) );
  AOI22_X1 U23066 ( .A1(n19898), .A2(n19889), .B1(n19989), .B2(n19866), .ZN(
        n19869) );
  AOI22_X1 U23067 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19867), .B1(
        n19992), .B2(n19990), .ZN(n19868) );
  OAI211_X1 U23068 ( .C1(n19903), .C2(n19870), .A(n19869), .B(n19868), .ZN(
        P3_U2971) );
  NOR2_X1 U23069 ( .A1(n19872), .A2(n19871), .ZN(n19944) );
  AOI22_X1 U23070 ( .A1(n19873), .A2(n19933), .B1(n19941), .B2(n19944), .ZN(
        n19879) );
  AOI22_X1 U23071 ( .A1(n19877), .A2(n19876), .B1(n19875), .B2(n19874), .ZN(
        n19899) );
  AOI22_X1 U23072 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19899), .B1(
        n19976), .B2(n19946), .ZN(n19878) );
  OAI211_X1 U23073 ( .C1(n19880), .C2(n19902), .A(n19879), .B(n19878), .ZN(
        P3_U2972) );
  AOI22_X1 U23074 ( .A1(n19951), .A2(n19933), .B1(n19950), .B2(n19944), .ZN(
        n19882) );
  AOI22_X1 U23075 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19899), .B1(
        n19976), .B2(n19952), .ZN(n19881) );
  OAI211_X1 U23076 ( .C1(n19955), .C2(n19902), .A(n19882), .B(n19881), .ZN(
        P3_U2973) );
  AOI22_X1 U23077 ( .A1(n19883), .A2(n19933), .B1(n19957), .B2(n19944), .ZN(
        n19885) );
  AOI22_X1 U23078 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19899), .B1(
        n19976), .B2(n19958), .ZN(n19884) );
  OAI211_X1 U23079 ( .C1(n19886), .C2(n19902), .A(n19885), .B(n19884), .ZN(
        P3_U2974) );
  AOI22_X1 U23080 ( .A1(n19963), .A2(n19889), .B1(n19962), .B2(n19944), .ZN(
        n19888) );
  AOI22_X1 U23081 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19899), .B1(
        n19976), .B2(n19964), .ZN(n19887) );
  OAI211_X1 U23082 ( .C1(n19967), .C2(n19924), .A(n19888), .B(n19887), .ZN(
        P3_U2975) );
  AOI22_X1 U23083 ( .A1(n19969), .A2(n19944), .B1(n19968), .B2(n19889), .ZN(
        n19891) );
  AOI22_X1 U23084 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19899), .B1(
        n19976), .B2(n19970), .ZN(n19890) );
  OAI211_X1 U23085 ( .C1(n19973), .C2(n19924), .A(n19891), .B(n19890), .ZN(
        P3_U2976) );
  AOI22_X1 U23086 ( .A1(n19975), .A2(n19933), .B1(n19974), .B2(n19944), .ZN(
        n19893) );
  AOI22_X1 U23087 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19899), .B1(
        n19976), .B2(n19977), .ZN(n19892) );
  OAI211_X1 U23088 ( .C1(n19981), .C2(n19902), .A(n19893), .B(n19892), .ZN(
        P3_U2977) );
  AOI22_X1 U23089 ( .A1(n19894), .A2(n19933), .B1(n19982), .B2(n19944), .ZN(
        n19896) );
  AOI22_X1 U23090 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19899), .B1(
        n19976), .B2(n19984), .ZN(n19895) );
  OAI211_X1 U23091 ( .C1(n19897), .C2(n19902), .A(n19896), .B(n19895), .ZN(
        P3_U2978) );
  AOI22_X1 U23092 ( .A1(n19898), .A2(n19933), .B1(n19989), .B2(n19944), .ZN(
        n19901) );
  AOI22_X1 U23093 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19899), .B1(
        n19976), .B2(n19992), .ZN(n19900) );
  OAI211_X1 U23094 ( .C1(n19903), .C2(n19902), .A(n19901), .B(n19900), .ZN(
        P3_U2979) );
  INV_X1 U23095 ( .A(n19990), .ZN(n19980) );
  NOR2_X1 U23096 ( .A1(n19904), .A2(n19939), .ZN(n19932) );
  AOI22_X1 U23097 ( .A1(n19941), .A2(n19932), .B1(n19940), .B2(n19933), .ZN(
        n19910) );
  OAI21_X1 U23098 ( .B1(n19906), .B2(n19905), .A(n19904), .ZN(n19907) );
  OAI211_X1 U23099 ( .C1(n19934), .C2(n20134), .A(n19908), .B(n19907), .ZN(
        n19935) );
  AOI22_X1 U23100 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19935), .B1(
        n19934), .B2(n19946), .ZN(n19909) );
  OAI211_X1 U23101 ( .C1(n19949), .C2(n19980), .A(n19910), .B(n19909), .ZN(
        P3_U2980) );
  AOI22_X1 U23102 ( .A1(n19911), .A2(n19933), .B1(n19950), .B2(n19932), .ZN(
        n19913) );
  AOI22_X1 U23103 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19935), .B1(
        n19934), .B2(n19952), .ZN(n19912) );
  OAI211_X1 U23104 ( .C1(n19914), .C2(n19980), .A(n19913), .B(n19912), .ZN(
        P3_U2981) );
  AOI22_X1 U23105 ( .A1(n19957), .A2(n19932), .B1(n19956), .B2(n19933), .ZN(
        n19916) );
  AOI22_X1 U23106 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19935), .B1(
        n19934), .B2(n19958), .ZN(n19915) );
  OAI211_X1 U23107 ( .C1(n19961), .C2(n19980), .A(n19916), .B(n19915), .ZN(
        P3_U2982) );
  AOI22_X1 U23108 ( .A1(n19917), .A2(n19990), .B1(n19962), .B2(n19932), .ZN(
        n19919) );
  AOI22_X1 U23109 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19935), .B1(
        n19934), .B2(n19964), .ZN(n19918) );
  OAI211_X1 U23110 ( .C1(n19920), .C2(n19924), .A(n19919), .B(n19918), .ZN(
        P3_U2983) );
  AOI22_X1 U23111 ( .A1(n19921), .A2(n19990), .B1(n19969), .B2(n19932), .ZN(
        n19923) );
  AOI22_X1 U23112 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19935), .B1(
        n19934), .B2(n19970), .ZN(n19922) );
  OAI211_X1 U23113 ( .C1(n19925), .C2(n19924), .A(n19923), .B(n19922), .ZN(
        P3_U2984) );
  AOI22_X1 U23114 ( .A1(n19926), .A2(n19933), .B1(n19974), .B2(n19932), .ZN(
        n19928) );
  AOI22_X1 U23115 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19935), .B1(
        n19934), .B2(n19977), .ZN(n19927) );
  OAI211_X1 U23116 ( .C1(n19929), .C2(n19980), .A(n19928), .B(n19927), .ZN(
        P3_U2985) );
  AOI22_X1 U23117 ( .A1(n19983), .A2(n19933), .B1(n19982), .B2(n19932), .ZN(
        n19931) );
  AOI22_X1 U23118 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19935), .B1(
        n19934), .B2(n19984), .ZN(n19930) );
  OAI211_X1 U23119 ( .C1(n19987), .C2(n19980), .A(n19931), .B(n19930), .ZN(
        P3_U2986) );
  AOI22_X1 U23120 ( .A1(n19991), .A2(n19933), .B1(n19989), .B2(n19932), .ZN(
        n19937) );
  AOI22_X1 U23121 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19935), .B1(
        n19934), .B2(n19992), .ZN(n19936) );
  OAI211_X1 U23122 ( .C1(n19997), .C2(n19980), .A(n19937), .B(n19936), .ZN(
        P3_U2987) );
  NOR2_X1 U23123 ( .A1(n19939), .A2(n19938), .ZN(n19988) );
  AOI22_X1 U23124 ( .A1(n19941), .A2(n19988), .B1(n19940), .B2(n19990), .ZN(
        n19948) );
  AOI22_X1 U23125 ( .A1(n19945), .A2(n19944), .B1(n19943), .B2(n19942), .ZN(
        n19994) );
  AOI22_X1 U23126 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19994), .B1(
        n19993), .B2(n19946), .ZN(n19947) );
  OAI211_X1 U23127 ( .C1(n19949), .C2(n19998), .A(n19948), .B(n19947), .ZN(
        P3_U2988) );
  AOI22_X1 U23128 ( .A1(n19976), .A2(n19951), .B1(n19950), .B2(n19988), .ZN(
        n19954) );
  AOI22_X1 U23129 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19994), .B1(
        n19993), .B2(n19952), .ZN(n19953) );
  OAI211_X1 U23130 ( .C1(n19955), .C2(n19980), .A(n19954), .B(n19953), .ZN(
        P3_U2989) );
  AOI22_X1 U23131 ( .A1(n19957), .A2(n19988), .B1(n19956), .B2(n19990), .ZN(
        n19960) );
  AOI22_X1 U23132 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19994), .B1(
        n19993), .B2(n19958), .ZN(n19959) );
  OAI211_X1 U23133 ( .C1(n19998), .C2(n19961), .A(n19960), .B(n19959), .ZN(
        P3_U2990) );
  AOI22_X1 U23134 ( .A1(n19963), .A2(n19990), .B1(n19962), .B2(n19988), .ZN(
        n19966) );
  AOI22_X1 U23135 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19994), .B1(
        n19993), .B2(n19964), .ZN(n19965) );
  OAI211_X1 U23136 ( .C1(n19998), .C2(n19967), .A(n19966), .B(n19965), .ZN(
        P3_U2991) );
  AOI22_X1 U23137 ( .A1(n19969), .A2(n19988), .B1(n19968), .B2(n19990), .ZN(
        n19972) );
  AOI22_X1 U23138 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19994), .B1(
        n19993), .B2(n19970), .ZN(n19971) );
  OAI211_X1 U23139 ( .C1(n19998), .C2(n19973), .A(n19972), .B(n19971), .ZN(
        P3_U2992) );
  AOI22_X1 U23140 ( .A1(n19976), .A2(n19975), .B1(n19974), .B2(n19988), .ZN(
        n19979) );
  AOI22_X1 U23141 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19994), .B1(
        n19993), .B2(n19977), .ZN(n19978) );
  OAI211_X1 U23142 ( .C1(n19981), .C2(n19980), .A(n19979), .B(n19978), .ZN(
        P3_U2993) );
  AOI22_X1 U23143 ( .A1(n19983), .A2(n19990), .B1(n19982), .B2(n19988), .ZN(
        n19986) );
  AOI22_X1 U23144 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19994), .B1(
        n19993), .B2(n19984), .ZN(n19985) );
  OAI211_X1 U23145 ( .C1(n19998), .C2(n19987), .A(n19986), .B(n19985), .ZN(
        P3_U2994) );
  AOI22_X1 U23146 ( .A1(n19991), .A2(n19990), .B1(n19989), .B2(n19988), .ZN(
        n19996) );
  AOI22_X1 U23147 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19994), .B1(
        n19993), .B2(n19992), .ZN(n19995) );
  OAI211_X1 U23148 ( .C1(n19998), .C2(n19997), .A(n19996), .B(n19995), .ZN(
        P3_U2995) );
  AOI22_X1 U23149 ( .A1(n20026), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n20000), .B2(n19999), .ZN(n20030) );
  INV_X1 U23150 ( .A(n20030), .ZN(n20008) );
  NOR2_X1 U23151 ( .A1(n20001), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20004) );
  NAND3_X1 U23152 ( .A1(n20001), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20002) );
  OAI21_X1 U23153 ( .B1(n20004), .B2(n20003), .A(n20002), .ZN(n20006) );
  OAI21_X1 U23154 ( .B1(n20026), .B2(n20006), .A(n20005), .ZN(n20007) );
  AOI222_X1 U23155 ( .A1(n11696), .A2(n20008), .B1(n11696), .B2(n20007), .C1(
        n20008), .C2(n20007), .ZN(n20015) );
  OAI21_X1 U23156 ( .B1(n20026), .B2(n20009), .A(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n20012) );
  OR2_X1 U23157 ( .A1(n20026), .A2(n20010), .ZN(n20011) );
  NAND2_X1 U23158 ( .A1(n20012), .A2(n20011), .ZN(n20032) );
  INV_X1 U23159 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20013) );
  OAI21_X1 U23160 ( .B1(n20032), .B2(n20013), .A(n19560), .ZN(n20014) );
  OR2_X1 U23161 ( .A1(n20015), .A2(n20014), .ZN(n20036) );
  NOR2_X1 U23162 ( .A1(P3_MORE_REG_SCAN_IN), .A2(P3_FLUSH_REG_SCAN_IN), .ZN(
        n20029) );
  OAI22_X1 U23163 ( .A1(n20019), .A2(n20018), .B1(n20017), .B2(n20016), .ZN(
        n20020) );
  AOI221_X1 U23164 ( .B1(n20023), .B2(n20022), .C1(n20021), .C2(n20022), .A(
        n20020), .ZN(n20147) );
  AOI211_X1 U23165 ( .C1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .C2(n20026), .A(
        n20025), .B(n20024), .ZN(n20027) );
  OAI211_X1 U23166 ( .C1(n20029), .C2(n20028), .A(n20147), .B(n20027), .ZN(
        n20034) );
  OAI21_X1 U23167 ( .B1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(n20030), .ZN(n20031) );
  AND2_X1 U23168 ( .A1(n20032), .A2(n20031), .ZN(n20033) );
  NOR2_X1 U23169 ( .A1(n20034), .A2(n20033), .ZN(n20035) );
  AOI22_X1 U23170 ( .A1(n20037), .A2(n20154), .B1(n20152), .B2(n18932), .ZN(
        n20045) );
  INV_X1 U23171 ( .A(n20038), .ZN(n20040) );
  INV_X1 U23172 ( .A(n20048), .ZN(n20039) );
  AOI211_X1 U23173 ( .C1(n20041), .C2(n20040), .A(n20047), .B(n20039), .ZN(
        n20042) );
  NOR2_X1 U23174 ( .A1(n20042), .A2(n20156), .ZN(n20135) );
  OAI211_X1 U23175 ( .C1(P3_STATE2_REG_2__SCAN_IN), .C2(n20161), .A(n20135), 
        .B(n20043), .ZN(n20052) );
  OAI22_X1 U23176 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n20045), .B1(n20044), 
        .B2(n20052), .ZN(n20046) );
  OAI21_X1 U23177 ( .B1(n20048), .B2(n20047), .A(n20046), .ZN(P3_U2996) );
  NOR4_X1 U23178 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n20156), .A3(n20049), 
        .A4(n20161), .ZN(n20054) );
  AOI211_X1 U23179 ( .C1(n20152), .C2(n18932), .A(n20050), .B(n20054), .ZN(
        n20051) );
  OAI21_X1 U23180 ( .B1(P3_STATE2_REG_1__SCAN_IN), .B2(n20052), .A(n20051), 
        .ZN(P3_U2997) );
  INV_X1 U23181 ( .A(n20133), .ZN(n20053) );
  NOR4_X1 U23182 ( .A1(n20154), .A2(n20055), .A3(n20054), .A4(n20053), .ZN(
        P3_U2998) );
  AND2_X1 U23183 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n20056), .ZN(
        P3_U2999) );
  AND2_X1 U23184 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n20056), .ZN(
        P3_U3000) );
  AND2_X1 U23185 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n20056), .ZN(
        P3_U3001) );
  AND2_X1 U23186 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n20056), .ZN(
        P3_U3002) );
  AND2_X1 U23187 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n20056), .ZN(
        P3_U3003) );
  AND2_X1 U23188 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n20056), .ZN(
        P3_U3004) );
  AND2_X1 U23189 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n20056), .ZN(
        P3_U3005) );
  AND2_X1 U23190 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n20056), .ZN(
        P3_U3006) );
  AND2_X1 U23191 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n20056), .ZN(
        P3_U3007) );
  AND2_X1 U23192 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n20056), .ZN(
        P3_U3008) );
  AND2_X1 U23193 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n20057), .ZN(
        P3_U3009) );
  AND2_X1 U23194 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n20057), .ZN(
        P3_U3010) );
  AND2_X1 U23195 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n20057), .ZN(
        P3_U3011) );
  AND2_X1 U23196 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n20057), .ZN(
        P3_U3012) );
  AND2_X1 U23197 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n20057), .ZN(
        P3_U3013) );
  AND2_X1 U23198 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n20057), .ZN(
        P3_U3014) );
  AND2_X1 U23199 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n20057), .ZN(
        P3_U3015) );
  AND2_X1 U23200 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n20057), .ZN(
        P3_U3016) );
  AND2_X1 U23201 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n20057), .ZN(
        P3_U3017) );
  AND2_X1 U23202 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n20057), .ZN(
        P3_U3018) );
  AND2_X1 U23203 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n20057), .ZN(
        P3_U3019) );
  INV_X1 U23204 ( .A(P3_DATAWIDTH_REG_10__SCAN_IN), .ZN(n21725) );
  NOR2_X1 U23205 ( .A1(n21725), .A2(n20132), .ZN(P3_U3020) );
  AND2_X1 U23206 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n20057), .ZN(P3_U3021) );
  AND2_X1 U23207 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n20056), .ZN(P3_U3022) );
  AND2_X1 U23208 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n20056), .ZN(P3_U3023) );
  AND2_X1 U23209 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n20056), .ZN(P3_U3024) );
  INV_X1 U23210 ( .A(P3_DATAWIDTH_REG_5__SCAN_IN), .ZN(n21765) );
  NOR2_X1 U23211 ( .A1(n21765), .A2(n20132), .ZN(P3_U3025) );
  AND2_X1 U23212 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n20057), .ZN(P3_U3026) );
  AND2_X1 U23213 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n20057), .ZN(P3_U3027) );
  AND2_X1 U23214 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n20057), .ZN(P3_U3028) );
  NAND2_X1 U23215 ( .A1(n20152), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n20071) );
  OAI21_X1 U23216 ( .B1(n20058), .B2(n20817), .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n20059) );
  AOI22_X1 U23217 ( .A1(n20067), .A2(n20072), .B1(n20164), .B2(n20059), .ZN(
        n20061) );
  NAND3_X1 U23218 ( .A1(NA), .A2(n20067), .A3(n20062), .ZN(n20060) );
  OAI211_X1 U23219 ( .C1(P3_STATE_REG_2__SCAN_IN), .C2(n20071), .A(n20061), 
        .B(n20060), .ZN(P3_U3029) );
  NOR3_X1 U23220 ( .A1(P3_STATE_REG_2__SCAN_IN), .A2(n20062), .A3(n20817), 
        .ZN(n20063) );
  AOI221_X1 U23221 ( .B1(n20064), .B2(P3_REQUESTPENDING_REG_SCAN_IN), .C1(
        n20817), .C2(P3_REQUESTPENDING_REG_SCAN_IN), .A(n20063), .ZN(n20066)
         );
  OAI211_X1 U23222 ( .C1(n20066), .C2(n20067), .A(n20071), .B(n20065), .ZN(
        P3_U3030) );
  INV_X1 U23223 ( .A(NA), .ZN(n21536) );
  OAI21_X1 U23224 ( .B1(P3_STATE_REG_1__SCAN_IN), .B2(n21536), .A(n20067), 
        .ZN(n20070) );
  OAI222_X1 U23225 ( .A1(n20072), .A2(n20817), .B1(P3_STATE_REG_1__SCAN_IN), 
        .B2(P3_REQUESTPENDING_REG_SCAN_IN), .C1(n20071), .C2(NA), .ZN(n20068)
         );
  OAI211_X1 U23226 ( .C1(P3_REQUESTPENDING_REG_SCAN_IN), .C2(HOLD), .A(
        P3_STATE_REG_0__SCAN_IN), .B(n20068), .ZN(n20069) );
  OAI221_X1 U23227 ( .B1(n20072), .B2(n20071), .C1(n20072), .C2(n20070), .A(
        n20069), .ZN(P3_U3031) );
  INV_X1 U23228 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n20074) );
  OAI222_X1 U23229 ( .A1(n20136), .A2(n20124), .B1(n20073), .B2(n20121), .C1(
        n20074), .C2(n20117), .ZN(P3_U3032) );
  OAI222_X1 U23230 ( .A1(n20117), .A2(n20077), .B1(n20075), .B2(n20121), .C1(
        n20074), .C2(n20124), .ZN(P3_U3033) );
  OAI222_X1 U23231 ( .A1(n20077), .A2(n20124), .B1(n20076), .B2(n20121), .C1(
        n20078), .C2(n20117), .ZN(P3_U3034) );
  OAI222_X1 U23232 ( .A1(n20117), .A2(n21714), .B1(n21865), .B2(n20121), .C1(
        n20078), .C2(n20124), .ZN(P3_U3035) );
  OAI222_X1 U23233 ( .A1(n21714), .A2(n20124), .B1(n20079), .B2(n20121), .C1(
        n21712), .C2(n20117), .ZN(P3_U3036) );
  OAI222_X1 U23234 ( .A1(n21712), .A2(n20124), .B1(n20080), .B2(n20121), .C1(
        n20081), .C2(n20117), .ZN(P3_U3037) );
  OAI222_X1 U23235 ( .A1(n20117), .A2(n20082), .B1(n21775), .B2(n20144), .C1(
        n20081), .C2(n20124), .ZN(P3_U3038) );
  OAI222_X1 U23236 ( .A1(n20117), .A2(n20084), .B1(n20083), .B2(n20121), .C1(
        n20082), .C2(n20124), .ZN(P3_U3039) );
  OAI222_X1 U23237 ( .A1(n20117), .A2(n20086), .B1(n20085), .B2(n20121), .C1(
        n20084), .C2(n20124), .ZN(P3_U3040) );
  OAI222_X1 U23238 ( .A1(n20117), .A2(n20087), .B1(n21823), .B2(n20121), .C1(
        n20086), .C2(n20124), .ZN(P3_U3041) );
  OAI222_X1 U23239 ( .A1(n20117), .A2(n20089), .B1(n20088), .B2(n20121), .C1(
        n20087), .C2(n20124), .ZN(P3_U3042) );
  OAI222_X1 U23240 ( .A1(n20117), .A2(n20091), .B1(n20090), .B2(n20144), .C1(
        n20089), .C2(n20124), .ZN(P3_U3043) );
  OAI222_X1 U23241 ( .A1(n20117), .A2(n20093), .B1(n20092), .B2(n20144), .C1(
        n20091), .C2(n20124), .ZN(P3_U3044) );
  OAI222_X1 U23242 ( .A1(n20117), .A2(n20095), .B1(n20094), .B2(n20144), .C1(
        n20093), .C2(n20124), .ZN(P3_U3045) );
  OAI222_X1 U23243 ( .A1(n20117), .A2(n20097), .B1(n20096), .B2(n20144), .C1(
        n20095), .C2(n20124), .ZN(P3_U3046) );
  OAI222_X1 U23244 ( .A1(n20117), .A2(n20099), .B1(n20098), .B2(n20144), .C1(
        n20097), .C2(n20124), .ZN(P3_U3047) );
  OAI222_X1 U23245 ( .A1(n20117), .A2(n20101), .B1(n20100), .B2(n20144), .C1(
        n20099), .C2(n20124), .ZN(P3_U3048) );
  OAI222_X1 U23246 ( .A1(n20117), .A2(n20104), .B1(n20102), .B2(n20144), .C1(
        n20101), .C2(n20124), .ZN(P3_U3049) );
  OAI222_X1 U23247 ( .A1(n20104), .A2(n20124), .B1(n20103), .B2(n20144), .C1(
        n20105), .C2(n20117), .ZN(P3_U3050) );
  OAI222_X1 U23248 ( .A1(n20117), .A2(n21832), .B1(n20106), .B2(n20144), .C1(
        n20105), .C2(n20124), .ZN(P3_U3051) );
  OAI222_X1 U23249 ( .A1(n21832), .A2(n20124), .B1(n20107), .B2(n20144), .C1(
        n20108), .C2(n20117), .ZN(P3_U3052) );
  INV_X1 U23250 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n20111) );
  OAI222_X1 U23251 ( .A1(n20117), .A2(n20111), .B1(n20109), .B2(n20144), .C1(
        n20108), .C2(n20124), .ZN(P3_U3053) );
  OAI222_X1 U23252 ( .A1(n20111), .A2(n20124), .B1(n20110), .B2(n20121), .C1(
        n21849), .C2(n20117), .ZN(P3_U3054) );
  OAI222_X1 U23253 ( .A1(n20117), .A2(n20113), .B1(n20112), .B2(n20121), .C1(
        n21849), .C2(n20124), .ZN(P3_U3055) );
  OAI222_X1 U23254 ( .A1(n20117), .A2(n20114), .B1(n21812), .B2(n20121), .C1(
        n20113), .C2(n20124), .ZN(P3_U3056) );
  OAI222_X1 U23255 ( .A1(n20117), .A2(n17779), .B1(n20115), .B2(n20121), .C1(
        n20114), .C2(n20124), .ZN(P3_U3057) );
  OAI222_X1 U23256 ( .A1(n20117), .A2(n13565), .B1(n20116), .B2(n20121), .C1(
        n17779), .C2(n20124), .ZN(P3_U3058) );
  OAI222_X1 U23257 ( .A1(n13565), .A2(n20124), .B1(n20118), .B2(n20121), .C1(
        n13399), .C2(n20117), .ZN(P3_U3059) );
  OAI222_X1 U23258 ( .A1(n20117), .A2(n20123), .B1(n20119), .B2(n20121), .C1(
        n13399), .C2(n20124), .ZN(P3_U3060) );
  OAI222_X1 U23259 ( .A1(n20124), .A2(n20123), .B1(n20122), .B2(n20121), .C1(
        n20120), .C2(n20117), .ZN(P3_U3061) );
  INV_X1 U23260 ( .A(P3_BE_N_REG_3__SCAN_IN), .ZN(n21716) );
  AOI22_X1 U23261 ( .A1(n20144), .A2(n20125), .B1(n21716), .B2(n20164), .ZN(
        P3_U3274) );
  OAI22_X1 U23262 ( .A1(n20164), .A2(P3_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P3_BE_N_REG_2__SCAN_IN), .B2(n20144), .ZN(n20126) );
  INV_X1 U23263 ( .A(n20126), .ZN(P3_U3275) );
  OAI22_X1 U23264 ( .A1(n20164), .A2(P3_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P3_BE_N_REG_1__SCAN_IN), .B2(n20144), .ZN(n20127) );
  INV_X1 U23265 ( .A(n20127), .ZN(P3_U3276) );
  OAI22_X1 U23266 ( .A1(n20164), .A2(P3_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P3_BE_N_REG_0__SCAN_IN), .B2(n20121), .ZN(n20128) );
  INV_X1 U23267 ( .A(n20128), .ZN(P3_U3277) );
  OAI21_X1 U23268 ( .B1(n20132), .B2(P3_DATAWIDTH_REG_0__SCAN_IN), .A(n20130), 
        .ZN(n20129) );
  INV_X1 U23269 ( .A(n20129), .ZN(P3_U3280) );
  OAI21_X1 U23270 ( .B1(n20132), .B2(n20131), .A(n20130), .ZN(P3_U3281) );
  OAI21_X1 U23271 ( .B1(n20135), .B2(n20134), .A(n20133), .ZN(P3_U3282) );
  AOI21_X1 U23272 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n20137) );
  AOI22_X1 U23273 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .B1(n20137), .B2(n20136), .ZN(n20140) );
  INV_X1 U23274 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n20139) );
  AOI22_X1 U23275 ( .A1(n20143), .A2(n20140), .B1(n20139), .B2(n20138), .ZN(
        P3_U3292) );
  INV_X1 U23276 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20142) );
  OAI21_X1 U23277 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(P3_REIP_REG_0__SCAN_IN), 
        .A(n20143), .ZN(n20141) );
  OAI21_X1 U23278 ( .B1(n20143), .B2(n20142), .A(n20141), .ZN(P3_U3293) );
  INV_X1 U23279 ( .A(P3_READREQUEST_REG_SCAN_IN), .ZN(n20170) );
  OAI22_X1 U23280 ( .A1(n20164), .A2(n20170), .B1(P3_W_R_N_REG_SCAN_IN), .B2(
        n20144), .ZN(n20145) );
  INV_X1 U23281 ( .A(n20145), .ZN(P3_U3294) );
  NAND2_X1 U23282 ( .A1(n20148), .A2(P3_MORE_REG_SCAN_IN), .ZN(n20146) );
  OAI21_X1 U23283 ( .B1(n20148), .B2(n20147), .A(n20146), .ZN(P3_U3295) );
  OAI21_X1 U23284 ( .B1(P3_STATEBS16_REG_SCAN_IN), .B2(n20150), .A(n20149), 
        .ZN(n20153) );
  AOI211_X1 U23285 ( .C1(n20168), .C2(n20153), .A(n20152), .B(n20151), .ZN(
        n20157) );
  INV_X1 U23286 ( .A(n20154), .ZN(n20155) );
  OAI21_X1 U23287 ( .B1(n20157), .B2(n20156), .A(n20155), .ZN(n20163) );
  OAI21_X1 U23288 ( .B1(n20159), .B2(n20158), .A(n20166), .ZN(n20160) );
  AOI21_X1 U23289 ( .B1(n18932), .B2(n20161), .A(n20160), .ZN(n20162) );
  MUX2_X1 U23290 ( .A(n20163), .B(P3_REQUESTPENDING_REG_SCAN_IN), .S(n20162), 
        .Z(P3_U3296) );
  OAI22_X1 U23291 ( .A1(n20164), .A2(P3_MEMORYFETCH_REG_SCAN_IN), .B1(
        P3_M_IO_N_REG_SCAN_IN), .B2(n20121), .ZN(n20165) );
  INV_X1 U23292 ( .A(n20165), .ZN(P3_U3297) );
  NAND2_X1 U23293 ( .A1(n20167), .A2(n20166), .ZN(n20173) );
  INV_X1 U23294 ( .A(n20173), .ZN(n20171) );
  AOI22_X1 U23295 ( .A1(n20171), .A2(n20170), .B1(n20169), .B2(n20168), .ZN(
        P3_U3298) );
  OAI21_X1 U23296 ( .B1(n20173), .B2(P3_MEMORYFETCH_REG_SCAN_IN), .A(n20172), 
        .ZN(n20174) );
  INV_X1 U23297 ( .A(n20174), .ZN(P3_U3299) );
  INV_X1 U23298 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n20177) );
  NAND2_X1 U23299 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n20827), .ZN(n20816) );
  NAND2_X1 U23300 ( .A1(n20177), .A2(n20175), .ZN(n20813) );
  OAI21_X1 U23301 ( .B1(n20177), .B2(n20816), .A(n20813), .ZN(n20884) );
  AOI21_X1 U23302 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(P2_ADS_N_REG_SCAN_IN), 
        .A(n20884), .ZN(n20176) );
  INV_X1 U23303 ( .A(n20176), .ZN(P2_U2815) );
  INV_X1 U23304 ( .A(n20807), .ZN(n20822) );
  NAND2_X1 U23305 ( .A1(n20177), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n20931) );
  INV_X2 U23306 ( .A(n20931), .ZN(n20930) );
  AOI22_X1 U23307 ( .A1(n20930), .A2(n20178), .B1(P2_D_C_N_REG_SCAN_IN), .B2(
        n20931), .ZN(n20179) );
  OAI21_X1 U23308 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n20822), .A(n20179), 
        .ZN(P2_U2817) );
  INV_X1 U23309 ( .A(BS16), .ZN(n21779) );
  AOI21_X1 U23310 ( .B1(n20822), .B2(n21779), .A(n20881), .ZN(n20880) );
  INV_X1 U23311 ( .A(n20880), .ZN(n20882) );
  OAI21_X1 U23312 ( .B1(n20884), .B2(n20691), .A(n20882), .ZN(P2_U2818) );
  AND2_X1 U23313 ( .A1(n20181), .A2(n20180), .ZN(n20928) );
  OAI21_X1 U23314 ( .B1(n20928), .B2(n18012), .A(n20182), .ZN(P2_U2819) );
  OAI21_X1 U23315 ( .B1(n20829), .B2(n20183), .A(n20185), .ZN(n20184) );
  OAI21_X1 U23316 ( .B1(n20185), .B2(P2_BYTEENABLE_REG_2__SCAN_IN), .A(n20184), 
        .ZN(n20186) );
  OAI221_X1 U23317 ( .B1(n20187), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n20187), .C2(P2_REIP_REG_0__SCAN_IN), .A(n20186), .ZN(P2_U2822) );
  AOI22_X1 U23318 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n20189), .B1(
        P2_EBX_REG_4__SCAN_IN), .B2(n20188), .ZN(n20209) );
  AOI21_X1 U23319 ( .B1(n20190), .B2(P2_REIP_REG_4__SCAN_IN), .A(n18058), .ZN(
        n20191) );
  OAI21_X1 U23320 ( .B1(n20193), .B2(n20192), .A(n20191), .ZN(n20194) );
  AOI21_X1 U23321 ( .B1(n20263), .B2(n20195), .A(n20194), .ZN(n20208) );
  OAI22_X1 U23322 ( .A1(n20198), .A2(n20197), .B1(n20196), .B2(n20258), .ZN(
        n20199) );
  INV_X1 U23323 ( .A(n20199), .ZN(n20207) );
  NAND2_X1 U23324 ( .A1(n20200), .A2(n20201), .ZN(n20202) );
  MUX2_X1 U23325 ( .A(n20202), .B(n20201), .S(n12943), .Z(n20205) );
  NAND3_X1 U23326 ( .A1(n20205), .A2(n20204), .A3(n20203), .ZN(n20206) );
  NAND4_X1 U23327 ( .A1(n20209), .A2(n20208), .A3(n20207), .A4(n20206), .ZN(
        P2_U2851) );
  NOR2_X1 U23328 ( .A1(n20241), .A2(n20210), .ZN(P2_U2920) );
  INV_X1 U23329 ( .A(n20211), .ZN(n20213) );
  AOI22_X1 U23330 ( .A1(n20213), .A2(P2_EAX_REG_18__SCAN_IN), .B1(
        P2_UWORD_REG_2__SCAN_IN), .B2(n20243), .ZN(n20212) );
  OAI21_X1 U23331 ( .B1(n21855), .B2(n20241), .A(n20212), .ZN(P2_U2933) );
  INV_X1 U23332 ( .A(P2_UWORD_REG_0__SCAN_IN), .ZN(n21792) );
  AOI22_X1 U23333 ( .A1(n20242), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n20213), 
        .B2(P2_EAX_REG_16__SCAN_IN), .ZN(n20214) );
  OAI21_X1 U23334 ( .B1(n21792), .B2(n20240), .A(n20214), .ZN(P2_U2935) );
  AOI22_X1 U23335 ( .A1(n20243), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n20242), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n20215) );
  OAI21_X1 U23336 ( .B1(n13629), .B2(n20245), .A(n20215), .ZN(P2_U2936) );
  AOI22_X1 U23337 ( .A1(n20243), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n20242), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n20216) );
  OAI21_X1 U23338 ( .B1(n20217), .B2(n20245), .A(n20216), .ZN(P2_U2937) );
  AOI22_X1 U23339 ( .A1(n20243), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n20242), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n20218) );
  OAI21_X1 U23340 ( .B1(n20219), .B2(n20245), .A(n20218), .ZN(P2_U2938) );
  AOI22_X1 U23341 ( .A1(n20243), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n20242), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n20220) );
  OAI21_X1 U23342 ( .B1(n20221), .B2(n20245), .A(n20220), .ZN(P2_U2939) );
  INV_X1 U23343 ( .A(P2_LWORD_REG_11__SCAN_IN), .ZN(n21697) );
  OAI222_X1 U23344 ( .A1(n20240), .A2(n21697), .B1(n20245), .B2(n20223), .C1(
        n20241), .C2(n20222), .ZN(P2_U2940) );
  AOI22_X1 U23345 ( .A1(n20243), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n20242), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n20224) );
  OAI21_X1 U23346 ( .B1(n20225), .B2(n20245), .A(n20224), .ZN(P2_U2941) );
  AOI22_X1 U23347 ( .A1(n20243), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n20242), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n20226) );
  OAI21_X1 U23348 ( .B1(n20227), .B2(n20245), .A(n20226), .ZN(P2_U2942) );
  AOI22_X1 U23349 ( .A1(n20243), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n20242), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n20228) );
  OAI21_X1 U23350 ( .B1(n20229), .B2(n20245), .A(n20228), .ZN(P2_U2943) );
  AOI22_X1 U23351 ( .A1(n20243), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n20242), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n20230) );
  OAI21_X1 U23352 ( .B1(n20231), .B2(n20245), .A(n20230), .ZN(P2_U2944) );
  AOI22_X1 U23353 ( .A1(n20243), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n20242), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n20232) );
  OAI21_X1 U23354 ( .B1(n20233), .B2(n20245), .A(n20232), .ZN(P2_U2945) );
  INV_X1 U23355 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n21868) );
  AOI22_X1 U23356 ( .A1(n20243), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n20242), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n20234) );
  OAI21_X1 U23357 ( .B1(n21868), .B2(n20245), .A(n20234), .ZN(P2_U2946) );
  INV_X1 U23358 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n20236) );
  AOI22_X1 U23359 ( .A1(n20243), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n20242), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n20235) );
  OAI21_X1 U23360 ( .B1(n20236), .B2(n20245), .A(n20235), .ZN(P2_U2947) );
  AOI22_X1 U23361 ( .A1(P2_EAX_REG_3__SCAN_IN), .A2(n20238), .B1(n20243), .B2(
        P2_LWORD_REG_3__SCAN_IN), .ZN(n20237) );
  OAI21_X1 U23362 ( .B1(n21732), .B2(n20241), .A(n20237), .ZN(P2_U2948) );
  AOI222_X1 U23363 ( .A1(n20242), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(n20238), 
        .B2(P2_EAX_REG_2__SCAN_IN), .C1(n20243), .C2(P2_LWORD_REG_2__SCAN_IN), 
        .ZN(n20239) );
  INV_X1 U23364 ( .A(n20239), .ZN(P2_U2949) );
  INV_X1 U23365 ( .A(P2_LWORD_REG_1__SCAN_IN), .ZN(n21749) );
  OAI222_X1 U23366 ( .A1(n20241), .A2(n21763), .B1(n20245), .B2(n11224), .C1(
        n20240), .C2(n21749), .ZN(P2_U2950) );
  AOI22_X1 U23367 ( .A1(n20243), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n20242), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n20244) );
  OAI21_X1 U23368 ( .B1(n11215), .B2(n20245), .A(n20244), .ZN(P2_U2951) );
  OAI21_X1 U23369 ( .B1(n20247), .B2(n20246), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n20248) );
  OAI21_X1 U23370 ( .B1(n20250), .B2(n20249), .A(n20248), .ZN(n20251) );
  AOI21_X1 U23371 ( .B1(n10091), .B2(n20252), .A(n20251), .ZN(n20254) );
  OAI211_X1 U23372 ( .C1(n20256), .C2(n20255), .A(n20254), .B(n20253), .ZN(
        P2_U3014) );
  NAND2_X1 U23373 ( .A1(n20257), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n20260) );
  OAI22_X1 U23374 ( .A1(n20261), .A2(n20260), .B1(n20259), .B2(n20258), .ZN(
        n20262) );
  INV_X1 U23375 ( .A(n20262), .ZN(n20272) );
  AOI22_X1 U23376 ( .A1(n20265), .A2(n20264), .B1(n20263), .B2(n20277), .ZN(
        n20271) );
  AOI22_X1 U23377 ( .A1(n20268), .A2(n20279), .B1(n20267), .B2(n20266), .ZN(
        n20270) );
  NAND4_X1 U23378 ( .A1(n20272), .A2(n20271), .A3(n20270), .A4(n20269), .ZN(
        P2_U3042) );
  AOI21_X1 U23379 ( .B1(n20275), .B2(n20274), .A(n20273), .ZN(n20296) );
  AOI22_X1 U23380 ( .A1(n20279), .A2(n20278), .B1(n20277), .B2(n20276), .ZN(
        n20294) );
  NAND2_X1 U23381 ( .A1(n20281), .A2(n20280), .ZN(n20283) );
  OAI211_X1 U23382 ( .C1(n20285), .C2(n20284), .A(n20283), .B(n20282), .ZN(
        n20292) );
  NAND2_X1 U23383 ( .A1(n20287), .A2(n20286), .ZN(n20289) );
  OAI21_X1 U23384 ( .B1(n20290), .B2(n20289), .A(n20288), .ZN(n20291) );
  NOR2_X1 U23385 ( .A1(n20292), .A2(n20291), .ZN(n20293) );
  OAI211_X1 U23386 ( .C1(n20296), .C2(n20295), .A(n20294), .B(n20293), .ZN(
        P2_U3044) );
  AOI22_X1 U23387 ( .A1(n20705), .A2(n20801), .B1(n20760), .B2(n20315), .ZN(
        n20298) );
  AOI22_X1 U23388 ( .A1(n20317), .A2(n20761), .B1(n20316), .B2(n20762), .ZN(
        n20297) );
  OAI211_X1 U23389 ( .C1(n20321), .C2(n20299), .A(n20298), .B(n20297), .ZN(
        P2_U3049) );
  OAI22_X1 U23390 ( .A1(n20310), .A2(n20771), .B1(n20309), .B2(n20709), .ZN(
        n20300) );
  INV_X1 U23391 ( .A(n20300), .ZN(n20302) );
  AOI22_X1 U23392 ( .A1(n20317), .A2(n20767), .B1(n20316), .B2(n20768), .ZN(
        n20301) );
  OAI211_X1 U23393 ( .C1(n20321), .C2(n20303), .A(n20302), .B(n20301), .ZN(
        P2_U3050) );
  OAI22_X1 U23394 ( .A1(n20310), .A2(n20777), .B1(n20309), .B2(n20555), .ZN(
        n20304) );
  INV_X1 U23395 ( .A(n20304), .ZN(n20306) );
  AOI22_X1 U23396 ( .A1(n20317), .A2(n20773), .B1(n20316), .B2(n20774), .ZN(
        n20305) );
  OAI211_X1 U23397 ( .C1(n20321), .C2(n20307), .A(n20306), .B(n20305), .ZN(
        P2_U3051) );
  INV_X1 U23398 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n20314) );
  OAI22_X1 U23399 ( .A1(n20310), .A2(n20783), .B1(n20309), .B2(n20308), .ZN(
        n20311) );
  INV_X1 U23400 ( .A(n20311), .ZN(n20313) );
  AOI22_X1 U23401 ( .A1(n20317), .A2(n20779), .B1(n20316), .B2(n20780), .ZN(
        n20312) );
  OAI211_X1 U23402 ( .C1(n20321), .C2(n20314), .A(n20313), .B(n20312), .ZN(
        P2_U3052) );
  INV_X1 U23403 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n20320) );
  AOI22_X1 U23404 ( .A1(n20733), .A2(n20801), .B1(n20315), .B2(n20797), .ZN(
        n20319) );
  AOI22_X1 U23405 ( .A1(n20317), .A2(n20798), .B1(n20316), .B2(n20800), .ZN(
        n20318) );
  OAI211_X1 U23406 ( .C1(n20321), .C2(n20320), .A(n20319), .B(n20318), .ZN(
        P2_U3055) );
  OR2_X1 U23407 ( .A1(n20351), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20324) );
  INV_X1 U23408 ( .A(n10926), .ZN(n20322) );
  NOR3_X2 U23409 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20919), .A3(
        n20351), .ZN(n20342) );
  OAI21_X1 U23410 ( .B1(n20322), .B2(n20342), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20323) );
  AOI22_X1 U23411 ( .A1(n20343), .A2(n20746), .B1(n20745), .B2(n20342), .ZN(
        n20329) );
  OAI22_X1 U23412 ( .A1(n20470), .A2(n20497), .B1(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n20351), .ZN(n20327) );
  INV_X1 U23413 ( .A(n20342), .ZN(n20325) );
  OAI211_X1 U23414 ( .C1(n10926), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n20692), 
        .B(n20325), .ZN(n20326) );
  NAND3_X1 U23415 ( .A1(n20327), .A2(n20748), .A3(n20326), .ZN(n20345) );
  AOI22_X1 U23416 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20345), .B1(
        n20344), .B2(n20756), .ZN(n20328) );
  OAI211_X1 U23417 ( .C1(n20759), .C2(n20348), .A(n20329), .B(n20328), .ZN(
        P2_U3056) );
  AOI22_X1 U23418 ( .A1(n20343), .A2(n20761), .B1(n20760), .B2(n20342), .ZN(
        n20331) );
  AOI22_X1 U23419 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20345), .B1(
        n20344), .B2(n20762), .ZN(n20330) );
  OAI211_X1 U23420 ( .C1(n20765), .C2(n20348), .A(n20331), .B(n20330), .ZN(
        P2_U3057) );
  AOI22_X1 U23421 ( .A1(n20343), .A2(n20767), .B1(n20766), .B2(n20342), .ZN(
        n20333) );
  AOI22_X1 U23422 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20345), .B1(
        n20344), .B2(n20768), .ZN(n20332) );
  OAI211_X1 U23423 ( .C1(n20771), .C2(n20348), .A(n20333), .B(n20332), .ZN(
        P2_U3058) );
  AOI22_X1 U23424 ( .A1(n20343), .A2(n20773), .B1(n20772), .B2(n20342), .ZN(
        n20335) );
  AOI22_X1 U23425 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20345), .B1(
        n20344), .B2(n20774), .ZN(n20334) );
  OAI211_X1 U23426 ( .C1(n20777), .C2(n20348), .A(n20335), .B(n20334), .ZN(
        P2_U3059) );
  AOI22_X1 U23427 ( .A1(n20343), .A2(n20779), .B1(n20778), .B2(n20342), .ZN(
        n20337) );
  AOI22_X1 U23428 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20345), .B1(
        n20344), .B2(n20780), .ZN(n20336) );
  OAI211_X1 U23429 ( .C1(n20783), .C2(n20348), .A(n20337), .B(n20336), .ZN(
        P2_U3060) );
  AOI22_X1 U23430 ( .A1(n20343), .A2(n20785), .B1(n20784), .B2(n20342), .ZN(
        n20339) );
  AOI22_X1 U23431 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20345), .B1(
        n20344), .B2(n20786), .ZN(n20338) );
  OAI211_X1 U23432 ( .C1(n20789), .C2(n20348), .A(n20339), .B(n20338), .ZN(
        P2_U3061) );
  AOI22_X1 U23433 ( .A1(n20343), .A2(n20791), .B1(n20790), .B2(n20342), .ZN(
        n20341) );
  AOI22_X1 U23434 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20345), .B1(
        n20344), .B2(n20792), .ZN(n20340) );
  OAI211_X1 U23435 ( .C1(n20795), .C2(n20348), .A(n20341), .B(n20340), .ZN(
        P2_U3062) );
  AOI22_X1 U23436 ( .A1(n20343), .A2(n20798), .B1(n20797), .B2(n20342), .ZN(
        n20347) );
  AOI22_X1 U23437 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20345), .B1(
        n20344), .B2(n20800), .ZN(n20346) );
  OAI211_X1 U23438 ( .C1(n20806), .C2(n20348), .A(n20347), .B(n20346), .ZN(
        P2_U3063) );
  INV_X1 U23439 ( .A(n20377), .ZN(n20371) );
  INV_X1 U23440 ( .A(n20351), .ZN(n20349) );
  NAND2_X1 U23441 ( .A1(n20604), .A2(n20349), .ZN(n20353) );
  INV_X1 U23442 ( .A(n20353), .ZN(n20376) );
  AOI22_X1 U23443 ( .A1(n20756), .A2(n20387), .B1(n20745), .B2(n20376), .ZN(
        n20362) );
  OAI21_X1 U23444 ( .B1(n20470), .B2(n20350), .A(n20888), .ZN(n20360) );
  NOR2_X1 U23445 ( .A1(n20909), .A2(n20351), .ZN(n20356) );
  INV_X1 U23446 ( .A(n20352), .ZN(n20357) );
  OAI21_X1 U23447 ( .B1(n20357), .B2(n20742), .A(n20750), .ZN(n20354) );
  AOI21_X1 U23448 ( .B1(n20354), .B2(n20353), .A(n20661), .ZN(n20355) );
  INV_X1 U23449 ( .A(n20356), .ZN(n20359) );
  OAI21_X1 U23450 ( .B1(n20357), .B2(n20376), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20358) );
  AOI22_X1 U23451 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20379), .B1(
        n20378), .B2(n20746), .ZN(n20361) );
  OAI211_X1 U23452 ( .C1(n20759), .C2(n20371), .A(n20362), .B(n20361), .ZN(
        P2_U3072) );
  AOI22_X1 U23453 ( .A1(n20705), .A2(n20377), .B1(n20760), .B2(n20376), .ZN(
        n20364) );
  AOI22_X1 U23454 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20379), .B1(
        n20378), .B2(n20761), .ZN(n20363) );
  OAI211_X1 U23455 ( .C1(n20708), .C2(n20412), .A(n20364), .B(n20363), .ZN(
        P2_U3073) );
  AOI22_X1 U23456 ( .A1(n20387), .A2(n20768), .B1(n20376), .B2(n20766), .ZN(
        n20366) );
  AOI22_X1 U23457 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20379), .B1(
        n20378), .B2(n20767), .ZN(n20365) );
  OAI211_X1 U23458 ( .C1(n20771), .C2(n20371), .A(n20366), .B(n20365), .ZN(
        P2_U3074) );
  AOI22_X1 U23459 ( .A1(n20774), .A2(n20387), .B1(n20772), .B2(n20376), .ZN(
        n20368) );
  AOI22_X1 U23460 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20379), .B1(
        n20378), .B2(n20773), .ZN(n20367) );
  OAI211_X1 U23461 ( .C1(n20777), .C2(n20371), .A(n20368), .B(n20367), .ZN(
        P2_U3075) );
  AOI22_X1 U23462 ( .A1(n20780), .A2(n20387), .B1(n20778), .B2(n20376), .ZN(
        n20370) );
  AOI22_X1 U23463 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20379), .B1(
        n20378), .B2(n20779), .ZN(n20369) );
  OAI211_X1 U23464 ( .C1(n20783), .C2(n20371), .A(n20370), .B(n20369), .ZN(
        P2_U3076) );
  AOI22_X1 U23465 ( .A1(n20377), .A2(n20678), .B1(n20376), .B2(n20784), .ZN(
        n20373) );
  AOI22_X1 U23466 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20379), .B1(
        n20378), .B2(n20785), .ZN(n20372) );
  OAI211_X1 U23467 ( .C1(n20720), .C2(n20412), .A(n20373), .B(n20372), .ZN(
        P2_U3077) );
  AOI22_X1 U23468 ( .A1(n20377), .A2(n20647), .B1(n20376), .B2(n20790), .ZN(
        n20375) );
  AOI22_X1 U23469 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20379), .B1(
        n20378), .B2(n20791), .ZN(n20374) );
  OAI211_X1 U23470 ( .C1(n20726), .C2(n20412), .A(n20375), .B(n20374), .ZN(
        P2_U3078) );
  AOI22_X1 U23471 ( .A1(n20733), .A2(n20377), .B1(n20797), .B2(n20376), .ZN(
        n20381) );
  AOI22_X1 U23472 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20379), .B1(
        n20378), .B2(n20798), .ZN(n20380) );
  OAI211_X1 U23473 ( .C1(n20738), .C2(n20412), .A(n20381), .B(n20380), .ZN(
        P2_U3079) );
  NAND3_X1 U23474 ( .A1(n20383), .A2(n20382), .A3(n21853), .ZN(n20390) );
  NOR2_X1 U23475 ( .A1(n20384), .A2(n20498), .ZN(n20407) );
  INV_X1 U23476 ( .A(n20407), .ZN(n20388) );
  NAND3_X1 U23477 ( .A1(n20385), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(n20388), 
        .ZN(n20392) );
  INV_X1 U23478 ( .A(n20392), .ZN(n20386) );
  AOI211_X2 U23479 ( .C1(n20742), .C2(n20390), .A(n20658), .B(n20386), .ZN(
        n20408) );
  AOI22_X1 U23480 ( .A1(n20408), .A2(n20746), .B1(n20745), .B2(n20407), .ZN(
        n20394) );
  OAI21_X1 U23481 ( .B1(n20387), .B2(n20430), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n20389) );
  AOI22_X1 U23482 ( .A1(n20390), .A2(n20389), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(n20388), .ZN(n20391) );
  NAND3_X1 U23483 ( .A1(n20392), .A2(n20391), .A3(n20748), .ZN(n20409) );
  AOI22_X1 U23484 ( .A1(n20756), .A2(n20430), .B1(
        P2_INSTQUEUE_REG_4__0__SCAN_IN), .B2(n20409), .ZN(n20393) );
  OAI211_X1 U23485 ( .C1(n20759), .C2(n20412), .A(n20394), .B(n20393), .ZN(
        P2_U3080) );
  AOI22_X1 U23486 ( .A1(n20408), .A2(n20761), .B1(n20760), .B2(n20407), .ZN(
        n20396) );
  AOI22_X1 U23487 ( .A1(n20430), .A2(n20762), .B1(
        P2_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n20409), .ZN(n20395) );
  OAI211_X1 U23488 ( .C1(n20765), .C2(n20412), .A(n20396), .B(n20395), .ZN(
        P2_U3081) );
  AOI22_X1 U23489 ( .A1(n20408), .A2(n20767), .B1(n20766), .B2(n20407), .ZN(
        n20398) );
  AOI22_X1 U23490 ( .A1(n20430), .A2(n20768), .B1(
        P2_INSTQUEUE_REG_4__2__SCAN_IN), .B2(n20409), .ZN(n20397) );
  OAI211_X1 U23491 ( .C1(n20771), .C2(n20412), .A(n20398), .B(n20397), .ZN(
        P2_U3082) );
  AOI22_X1 U23492 ( .A1(n20408), .A2(n20773), .B1(n20772), .B2(n20407), .ZN(
        n20400) );
  AOI22_X1 U23493 ( .A1(n20774), .A2(n20430), .B1(
        P2_INSTQUEUE_REG_4__3__SCAN_IN), .B2(n20409), .ZN(n20399) );
  OAI211_X1 U23494 ( .C1(n20777), .C2(n20412), .A(n20400), .B(n20399), .ZN(
        P2_U3083) );
  AOI22_X1 U23495 ( .A1(n20408), .A2(n20779), .B1(n20778), .B2(n20407), .ZN(
        n20402) );
  AOI22_X1 U23496 ( .A1(n20780), .A2(n20430), .B1(
        P2_INSTQUEUE_REG_4__4__SCAN_IN), .B2(n20409), .ZN(n20401) );
  OAI211_X1 U23497 ( .C1(n20783), .C2(n20412), .A(n20402), .B(n20401), .ZN(
        P2_U3084) );
  AOI22_X1 U23498 ( .A1(n20408), .A2(n20785), .B1(n20784), .B2(n20407), .ZN(
        n20404) );
  AOI22_X1 U23499 ( .A1(n20430), .A2(n20786), .B1(
        P2_INSTQUEUE_REG_4__5__SCAN_IN), .B2(n20409), .ZN(n20403) );
  OAI211_X1 U23500 ( .C1(n20789), .C2(n20412), .A(n20404), .B(n20403), .ZN(
        P2_U3085) );
  AOI22_X1 U23501 ( .A1(n20408), .A2(n20791), .B1(n20790), .B2(n20407), .ZN(
        n20406) );
  AOI22_X1 U23502 ( .A1(n20430), .A2(n20792), .B1(
        P2_INSTQUEUE_REG_4__6__SCAN_IN), .B2(n20409), .ZN(n20405) );
  OAI211_X1 U23503 ( .C1(n20795), .C2(n20412), .A(n20406), .B(n20405), .ZN(
        P2_U3086) );
  AOI22_X1 U23504 ( .A1(n20408), .A2(n20798), .B1(n20797), .B2(n20407), .ZN(
        n20411) );
  AOI22_X1 U23505 ( .A1(n20430), .A2(n20800), .B1(
        P2_INSTQUEUE_REG_4__7__SCAN_IN), .B2(n20409), .ZN(n20410) );
  OAI211_X1 U23506 ( .C1(n20806), .C2(n20412), .A(n20411), .B(n20410), .ZN(
        P2_U3087) );
  INV_X1 U23507 ( .A(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n20415) );
  AOI22_X1 U23508 ( .A1(n20440), .A2(n20762), .B1(n20760), .B2(n20429), .ZN(
        n20414) );
  AOI22_X1 U23509 ( .A1(n20761), .A2(n20431), .B1(n20705), .B2(n20430), .ZN(
        n20413) );
  OAI211_X1 U23510 ( .C1(n20435), .C2(n20415), .A(n20414), .B(n20413), .ZN(
        P2_U3089) );
  INV_X1 U23511 ( .A(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n20418) );
  AOI22_X1 U23512 ( .A1(n20440), .A2(n20768), .B1(n20766), .B2(n20429), .ZN(
        n20417) );
  AOI22_X1 U23513 ( .A1(n20431), .A2(n20767), .B1(n20430), .B2(n20634), .ZN(
        n20416) );
  OAI211_X1 U23514 ( .C1(n20435), .C2(n20418), .A(n20417), .B(n20416), .ZN(
        P2_U3090) );
  AOI22_X1 U23515 ( .A1(n20774), .A2(n20440), .B1(n20429), .B2(n20772), .ZN(
        n20420) );
  AOI22_X1 U23516 ( .A1(n20431), .A2(n20773), .B1(n20430), .B2(n20638), .ZN(
        n20419) );
  OAI211_X1 U23517 ( .C1(n20435), .C2(n20421), .A(n20420), .B(n20419), .ZN(
        P2_U3091) );
  INV_X1 U23518 ( .A(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n20424) );
  AOI22_X1 U23519 ( .A1(n20430), .A2(n20641), .B1(n20429), .B2(n20778), .ZN(
        n20423) );
  AOI22_X1 U23520 ( .A1(n20779), .A2(n20431), .B1(n20780), .B2(n20440), .ZN(
        n20422) );
  OAI211_X1 U23521 ( .C1(n20435), .C2(n20424), .A(n20423), .B(n20422), .ZN(
        P2_U3092) );
  AOI22_X1 U23522 ( .A1(n20430), .A2(n20678), .B1(n20429), .B2(n20784), .ZN(
        n20426) );
  AOI22_X1 U23523 ( .A1(n20431), .A2(n20785), .B1(n20440), .B2(n20786), .ZN(
        n20425) );
  OAI211_X1 U23524 ( .C1(n20435), .C2(n10930), .A(n20426), .B(n20425), .ZN(
        P2_U3093) );
  AOI22_X1 U23525 ( .A1(n20430), .A2(n20647), .B1(n20429), .B2(n20790), .ZN(
        n20428) );
  AOI22_X1 U23526 ( .A1(n20431), .A2(n20791), .B1(n20440), .B2(n20792), .ZN(
        n20427) );
  OAI211_X1 U23527 ( .C1(n20435), .C2(n10962), .A(n20428), .B(n20427), .ZN(
        P2_U3094) );
  INV_X1 U23528 ( .A(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n20434) );
  AOI22_X1 U23529 ( .A1(n20440), .A2(n20800), .B1(n20797), .B2(n20429), .ZN(
        n20433) );
  AOI22_X1 U23530 ( .A1(n20798), .A2(n20431), .B1(n20733), .B2(n20430), .ZN(
        n20432) );
  OAI211_X1 U23531 ( .C1(n20435), .C2(n20434), .A(n20433), .B(n20432), .ZN(
        P2_U3095) );
  NAND2_X1 U23532 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20437), .ZN(
        n20471) );
  NOR2_X1 U23533 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20471), .ZN(
        n20460) );
  INV_X1 U23534 ( .A(n20460), .ZN(n20441) );
  NAND3_X1 U23535 ( .A1(n20436), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(n20441), 
        .ZN(n20445) );
  NAND2_X1 U23536 ( .A1(n20695), .A2(n20437), .ZN(n20443) );
  OAI21_X1 U23537 ( .B1(n20443), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n20742), 
        .ZN(n20438) );
  AOI22_X1 U23538 ( .A1(n20461), .A2(n20746), .B1(n20745), .B2(n20460), .ZN(
        n20447) );
  OAI21_X1 U23539 ( .B1(n20440), .B2(n20493), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n20442) );
  AOI22_X1 U23540 ( .A1(n20443), .A2(n20442), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(n20441), .ZN(n20444) );
  NAND3_X1 U23541 ( .A1(n20445), .A2(n20444), .A3(n20748), .ZN(n20462) );
  AOI22_X1 U23542 ( .A1(n20756), .A2(n20493), .B1(
        P2_INSTQUEUE_REG_6__0__SCAN_IN), .B2(n20462), .ZN(n20446) );
  OAI211_X1 U23543 ( .C1(n20759), .C2(n20465), .A(n20447), .B(n20446), .ZN(
        P2_U3096) );
  AOI22_X1 U23544 ( .A1(n20461), .A2(n20761), .B1(n20760), .B2(n20460), .ZN(
        n20449) );
  AOI22_X1 U23545 ( .A1(n20493), .A2(n20762), .B1(
        P2_INSTQUEUE_REG_6__1__SCAN_IN), .B2(n20462), .ZN(n20448) );
  OAI211_X1 U23546 ( .C1(n20765), .C2(n20465), .A(n20449), .B(n20448), .ZN(
        P2_U3097) );
  AOI22_X1 U23547 ( .A1(n20461), .A2(n20767), .B1(n20766), .B2(n20460), .ZN(
        n20451) );
  AOI22_X1 U23548 ( .A1(n20493), .A2(n20768), .B1(
        P2_INSTQUEUE_REG_6__2__SCAN_IN), .B2(n20462), .ZN(n20450) );
  OAI211_X1 U23549 ( .C1(n20771), .C2(n20465), .A(n20451), .B(n20450), .ZN(
        P2_U3098) );
  AOI22_X1 U23550 ( .A1(n20461), .A2(n20773), .B1(n20772), .B2(n20460), .ZN(
        n20453) );
  AOI22_X1 U23551 ( .A1(n20774), .A2(n20493), .B1(
        P2_INSTQUEUE_REG_6__3__SCAN_IN), .B2(n20462), .ZN(n20452) );
  OAI211_X1 U23552 ( .C1(n20777), .C2(n20465), .A(n20453), .B(n20452), .ZN(
        P2_U3099) );
  AOI22_X1 U23553 ( .A1(n20461), .A2(n20779), .B1(n20778), .B2(n20460), .ZN(
        n20455) );
  AOI22_X1 U23554 ( .A1(n20780), .A2(n20493), .B1(
        P2_INSTQUEUE_REG_6__4__SCAN_IN), .B2(n20462), .ZN(n20454) );
  OAI211_X1 U23555 ( .C1(n20783), .C2(n20465), .A(n20455), .B(n20454), .ZN(
        P2_U3100) );
  AOI22_X1 U23556 ( .A1(n20461), .A2(n20785), .B1(n20784), .B2(n20460), .ZN(
        n20457) );
  AOI22_X1 U23557 ( .A1(n20493), .A2(n20786), .B1(
        P2_INSTQUEUE_REG_6__5__SCAN_IN), .B2(n20462), .ZN(n20456) );
  OAI211_X1 U23558 ( .C1(n20789), .C2(n20465), .A(n20457), .B(n20456), .ZN(
        P2_U3101) );
  AOI22_X1 U23559 ( .A1(n20461), .A2(n20791), .B1(n20790), .B2(n20460), .ZN(
        n20459) );
  AOI22_X1 U23560 ( .A1(n20493), .A2(n20792), .B1(
        P2_INSTQUEUE_REG_6__6__SCAN_IN), .B2(n20462), .ZN(n20458) );
  OAI211_X1 U23561 ( .C1(n20795), .C2(n20465), .A(n20459), .B(n20458), .ZN(
        P2_U3102) );
  AOI22_X1 U23562 ( .A1(n20461), .A2(n20798), .B1(n20797), .B2(n20460), .ZN(
        n20464) );
  AOI22_X1 U23563 ( .A1(n20493), .A2(n20800), .B1(
        P2_INSTQUEUE_REG_6__7__SCAN_IN), .B2(n20462), .ZN(n20463) );
  OAI211_X1 U23564 ( .C1(n20806), .C2(n20465), .A(n20464), .B(n20463), .ZN(
        P2_U3103) );
  INV_X1 U23565 ( .A(n20493), .ZN(n20487) );
  AND2_X1 U23566 ( .A1(n20469), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n20466) );
  NAND2_X1 U23567 ( .A1(n20467), .A2(n20466), .ZN(n20472) );
  OAI21_X1 U23568 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n20471), .A(n20742), 
        .ZN(n20468) );
  AND2_X1 U23569 ( .A1(n20472), .A2(n20468), .ZN(n20492) );
  INV_X1 U23570 ( .A(n20469), .ZN(n20503) );
  AOI22_X1 U23571 ( .A1(n20492), .A2(n20746), .B1(n20503), .B2(n20745), .ZN(
        n20478) );
  NOR2_X1 U23572 ( .A1(n20470), .A2(n20747), .ZN(n20887) );
  INV_X1 U23573 ( .A(n20471), .ZN(n20475) );
  OAI211_X1 U23574 ( .C1(n20503), .C2(n20750), .A(n20472), .B(n20748), .ZN(
        n20473) );
  INV_X1 U23575 ( .A(n20473), .ZN(n20474) );
  AOI22_X1 U23576 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20494), .B1(
        n20499), .B2(n20756), .ZN(n20477) );
  OAI211_X1 U23577 ( .C1(n20759), .C2(n20487), .A(n20478), .B(n20477), .ZN(
        P2_U3104) );
  AOI22_X1 U23578 ( .A1(n20492), .A2(n20761), .B1(n20503), .B2(n20760), .ZN(
        n20480) );
  AOI22_X1 U23579 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20494), .B1(
        n20493), .B2(n20705), .ZN(n20479) );
  OAI211_X1 U23580 ( .C1(n20708), .C2(n20534), .A(n20480), .B(n20479), .ZN(
        P2_U3105) );
  AOI22_X1 U23581 ( .A1(n20492), .A2(n20767), .B1(n20503), .B2(n20766), .ZN(
        n20482) );
  AOI22_X1 U23582 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20494), .B1(
        n20493), .B2(n20634), .ZN(n20481) );
  OAI211_X1 U23583 ( .C1(n20713), .C2(n20534), .A(n20482), .B(n20481), .ZN(
        P2_U3106) );
  AOI22_X1 U23584 ( .A1(n20492), .A2(n20773), .B1(n20503), .B2(n20772), .ZN(
        n20484) );
  AOI22_X1 U23585 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20494), .B1(
        n20499), .B2(n20774), .ZN(n20483) );
  OAI211_X1 U23586 ( .C1(n20777), .C2(n20487), .A(n20484), .B(n20483), .ZN(
        P2_U3107) );
  AOI22_X1 U23587 ( .A1(n20492), .A2(n20779), .B1(n20503), .B2(n20778), .ZN(
        n20486) );
  AOI22_X1 U23588 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20494), .B1(
        n20499), .B2(n20780), .ZN(n20485) );
  OAI211_X1 U23589 ( .C1(n20783), .C2(n20487), .A(n20486), .B(n20485), .ZN(
        P2_U3108) );
  AOI22_X1 U23590 ( .A1(n20492), .A2(n20785), .B1(n20503), .B2(n20784), .ZN(
        n20489) );
  AOI22_X1 U23591 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20494), .B1(
        n20493), .B2(n20678), .ZN(n20488) );
  OAI211_X1 U23592 ( .C1(n20720), .C2(n20534), .A(n20489), .B(n20488), .ZN(
        P2_U3109) );
  AOI22_X1 U23593 ( .A1(n20492), .A2(n20791), .B1(n20503), .B2(n20790), .ZN(
        n20491) );
  AOI22_X1 U23594 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20494), .B1(
        n20493), .B2(n20647), .ZN(n20490) );
  OAI211_X1 U23595 ( .C1(n20726), .C2(n20534), .A(n20491), .B(n20490), .ZN(
        P2_U3110) );
  AOI22_X1 U23596 ( .A1(n20492), .A2(n20798), .B1(n20503), .B2(n20797), .ZN(
        n20496) );
  AOI22_X1 U23597 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20494), .B1(
        n20493), .B2(n20733), .ZN(n20495) );
  OAI211_X1 U23598 ( .C1(n20738), .C2(n20534), .A(n20496), .B(n20495), .ZN(
        P2_U3111) );
  OR2_X2 U23599 ( .A1(n20690), .A2(n20497), .ZN(n20556) );
  NOR2_X1 U23600 ( .A1(n20498), .A2(n20602), .ZN(n20519) );
  AOI22_X1 U23601 ( .A1(n20756), .A2(n20577), .B1(n20745), .B2(n20519), .ZN(
        n20509) );
  OAI21_X1 U23602 ( .B1(n20577), .B2(n20499), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n20500) );
  NAND2_X1 U23603 ( .A1(n20500), .A2(n20888), .ZN(n20507) );
  NOR2_X1 U23604 ( .A1(n20507), .A2(n20503), .ZN(n20501) );
  OAI21_X2 U23605 ( .B1(n20502), .B2(n20519), .A(n20748), .ZN(n20531) );
  NOR2_X1 U23606 ( .A1(n20503), .A2(n20519), .ZN(n20506) );
  OAI21_X1 U23607 ( .B1(n20504), .B2(n20519), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20505) );
  AOI22_X1 U23608 ( .A1(n20531), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n20746), .B2(n20530), .ZN(n20508) );
  OAI211_X1 U23609 ( .C1(n20759), .C2(n20534), .A(n20509), .B(n20508), .ZN(
        P2_U3112) );
  INV_X1 U23610 ( .A(n20519), .ZN(n20528) );
  OAI22_X1 U23611 ( .A1(n20556), .A2(n20708), .B1(n20510), .B2(n20528), .ZN(
        n20511) );
  INV_X1 U23612 ( .A(n20511), .ZN(n20513) );
  AOI22_X1 U23613 ( .A1(n20531), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n20761), .B2(n20530), .ZN(n20512) );
  OAI211_X1 U23614 ( .C1(n20765), .C2(n20534), .A(n20513), .B(n20512), .ZN(
        P2_U3113) );
  OAI22_X1 U23615 ( .A1(n20556), .A2(n20713), .B1(n20709), .B2(n20528), .ZN(
        n20514) );
  INV_X1 U23616 ( .A(n20514), .ZN(n20516) );
  AOI22_X1 U23617 ( .A1(n20531), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n20767), .B2(n20530), .ZN(n20515) );
  OAI211_X1 U23618 ( .C1(n20771), .C2(n20534), .A(n20516), .B(n20515), .ZN(
        P2_U3114) );
  AOI22_X1 U23619 ( .A1(n20774), .A2(n20577), .B1(n20772), .B2(n20519), .ZN(
        n20518) );
  AOI22_X1 U23620 ( .A1(n20531), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n20773), .B2(n20530), .ZN(n20517) );
  OAI211_X1 U23621 ( .C1(n20777), .C2(n20534), .A(n20518), .B(n20517), .ZN(
        P2_U3115) );
  AOI22_X1 U23622 ( .A1(n20780), .A2(n20577), .B1(n20778), .B2(n20519), .ZN(
        n20521) );
  AOI22_X1 U23623 ( .A1(n20531), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n20779), .B2(n20530), .ZN(n20520) );
  OAI211_X1 U23624 ( .C1(n20783), .C2(n20534), .A(n20521), .B(n20520), .ZN(
        P2_U3116) );
  OAI22_X1 U23625 ( .A1(n20556), .A2(n20720), .B1(n20719), .B2(n20528), .ZN(
        n20522) );
  INV_X1 U23626 ( .A(n20522), .ZN(n20524) );
  AOI22_X1 U23627 ( .A1(n20531), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n20785), .B2(n20530), .ZN(n20523) );
  OAI211_X1 U23628 ( .C1(n20789), .C2(n20534), .A(n20524), .B(n20523), .ZN(
        P2_U3117) );
  OAI22_X1 U23629 ( .A1(n20556), .A2(n20726), .B1(n20724), .B2(n20528), .ZN(
        n20525) );
  INV_X1 U23630 ( .A(n20525), .ZN(n20527) );
  AOI22_X1 U23631 ( .A1(n20531), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n20791), .B2(n20530), .ZN(n20526) );
  OAI211_X1 U23632 ( .C1(n20795), .C2(n20534), .A(n20527), .B(n20526), .ZN(
        P2_U3118) );
  OAI22_X1 U23633 ( .A1(n20556), .A2(n20738), .B1(n20574), .B2(n20528), .ZN(
        n20529) );
  INV_X1 U23634 ( .A(n20529), .ZN(n20533) );
  AOI22_X1 U23635 ( .A1(n20531), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n20798), .B2(n20530), .ZN(n20532) );
  OAI211_X1 U23636 ( .C1(n20806), .C2(n20534), .A(n20533), .B(n20532), .ZN(
        P2_U3119) );
  AOI21_X1 U23637 ( .B1(n20753), .B2(n20536), .A(n20692), .ZN(n20540) );
  AOI21_X1 U23638 ( .B1(n20541), .B2(n20575), .A(n20742), .ZN(n20537) );
  INV_X1 U23639 ( .A(n20746), .ZN(n20547) );
  OAI22_X1 U23640 ( .A1(n20556), .A2(n20759), .B1(n20538), .B2(n20575), .ZN(
        n20539) );
  INV_X1 U23641 ( .A(n20539), .ZN(n20546) );
  INV_X1 U23642 ( .A(n20540), .ZN(n20544) );
  OAI211_X1 U23643 ( .C1(n20541), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n20575), 
        .B(n20692), .ZN(n20542) );
  OAI211_X1 U23644 ( .C1(n20544), .C2(n20543), .A(n20748), .B(n20542), .ZN(
        n20578) );
  AOI22_X1 U23645 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20578), .B1(
        n20562), .B2(n20756), .ZN(n20545) );
  OAI211_X1 U23646 ( .C1(n20582), .C2(n20547), .A(n20546), .B(n20545), .ZN(
        P2_U3120) );
  INV_X1 U23647 ( .A(n20761), .ZN(n20550) );
  INV_X1 U23648 ( .A(n20575), .ZN(n20561) );
  AOI22_X1 U23649 ( .A1(n20705), .A2(n20577), .B1(n20760), .B2(n20561), .ZN(
        n20549) );
  AOI22_X1 U23650 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20578), .B1(
        n20562), .B2(n20762), .ZN(n20548) );
  OAI211_X1 U23651 ( .C1(n20582), .C2(n20550), .A(n20549), .B(n20548), .ZN(
        P2_U3121) );
  INV_X1 U23652 ( .A(n20767), .ZN(n20554) );
  OAI22_X1 U23653 ( .A1(n20556), .A2(n20771), .B1(n20709), .B2(n20575), .ZN(
        n20551) );
  INV_X1 U23654 ( .A(n20551), .ZN(n20553) );
  AOI22_X1 U23655 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20578), .B1(
        n20562), .B2(n20768), .ZN(n20552) );
  OAI211_X1 U23656 ( .C1(n20582), .C2(n20554), .A(n20553), .B(n20552), .ZN(
        P2_U3122) );
  INV_X1 U23657 ( .A(n20773), .ZN(n20560) );
  OAI22_X1 U23658 ( .A1(n20556), .A2(n20777), .B1(n20555), .B2(n20575), .ZN(
        n20557) );
  INV_X1 U23659 ( .A(n20557), .ZN(n20559) );
  AOI22_X1 U23660 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20578), .B1(
        n20562), .B2(n20774), .ZN(n20558) );
  OAI211_X1 U23661 ( .C1(n20582), .C2(n20560), .A(n20559), .B(n20558), .ZN(
        P2_U3123) );
  INV_X1 U23662 ( .A(n20779), .ZN(n20565) );
  AOI22_X1 U23663 ( .A1(n20780), .A2(n20562), .B1(n20778), .B2(n20561), .ZN(
        n20564) );
  AOI22_X1 U23664 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20578), .B1(
        n20577), .B2(n20641), .ZN(n20563) );
  OAI211_X1 U23665 ( .C1(n20582), .C2(n20565), .A(n20564), .B(n20563), .ZN(
        P2_U3124) );
  INV_X1 U23666 ( .A(n20785), .ZN(n20569) );
  OAI22_X1 U23667 ( .A1(n20601), .A2(n20720), .B1(n20575), .B2(n20719), .ZN(
        n20566) );
  INV_X1 U23668 ( .A(n20566), .ZN(n20568) );
  AOI22_X1 U23669 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20578), .B1(
        n20577), .B2(n20678), .ZN(n20567) );
  OAI211_X1 U23670 ( .C1(n20582), .C2(n20569), .A(n20568), .B(n20567), .ZN(
        P2_U3125) );
  INV_X1 U23671 ( .A(n20791), .ZN(n20573) );
  OAI22_X1 U23672 ( .A1(n20601), .A2(n20726), .B1(n20575), .B2(n20724), .ZN(
        n20570) );
  INV_X1 U23673 ( .A(n20570), .ZN(n20572) );
  AOI22_X1 U23674 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20578), .B1(
        n20577), .B2(n20647), .ZN(n20571) );
  OAI211_X1 U23675 ( .C1(n20582), .C2(n20573), .A(n20572), .B(n20571), .ZN(
        P2_U3126) );
  INV_X1 U23676 ( .A(n20798), .ZN(n20581) );
  OAI22_X1 U23677 ( .A1(n20601), .A2(n20738), .B1(n20575), .B2(n20574), .ZN(
        n20576) );
  INV_X1 U23678 ( .A(n20576), .ZN(n20580) );
  AOI22_X1 U23679 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20578), .B1(
        n20577), .B2(n20733), .ZN(n20579) );
  OAI211_X1 U23680 ( .C1(n20582), .C2(n20581), .A(n20580), .B(n20579), .ZN(
        P2_U3127) );
  AOI22_X1 U23681 ( .A1(n20596), .A2(n20761), .B1(n20760), .B2(n20595), .ZN(
        n20584) );
  AOI22_X1 U23682 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20598), .B1(
        n20597), .B2(n20762), .ZN(n20583) );
  OAI211_X1 U23683 ( .C1(n20765), .C2(n20601), .A(n20584), .B(n20583), .ZN(
        P2_U3129) );
  AOI22_X1 U23684 ( .A1(n20596), .A2(n20767), .B1(n20766), .B2(n20595), .ZN(
        n20586) );
  AOI22_X1 U23685 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20598), .B1(
        n20597), .B2(n20768), .ZN(n20585) );
  OAI211_X1 U23686 ( .C1(n20771), .C2(n20601), .A(n20586), .B(n20585), .ZN(
        P2_U3130) );
  AOI22_X1 U23687 ( .A1(n20596), .A2(n20773), .B1(n20772), .B2(n20595), .ZN(
        n20588) );
  AOI22_X1 U23688 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20598), .B1(
        n20597), .B2(n20774), .ZN(n20587) );
  OAI211_X1 U23689 ( .C1(n20777), .C2(n20601), .A(n20588), .B(n20587), .ZN(
        P2_U3131) );
  AOI22_X1 U23690 ( .A1(n20596), .A2(n20779), .B1(n20778), .B2(n20595), .ZN(
        n20590) );
  AOI22_X1 U23691 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20598), .B1(
        n20597), .B2(n20780), .ZN(n20589) );
  OAI211_X1 U23692 ( .C1(n20783), .C2(n20601), .A(n20590), .B(n20589), .ZN(
        P2_U3132) );
  AOI22_X1 U23693 ( .A1(n20596), .A2(n20785), .B1(n20784), .B2(n20595), .ZN(
        n20592) );
  AOI22_X1 U23694 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20598), .B1(
        n20597), .B2(n20786), .ZN(n20591) );
  OAI211_X1 U23695 ( .C1(n20789), .C2(n20601), .A(n20592), .B(n20591), .ZN(
        P2_U3133) );
  AOI22_X1 U23696 ( .A1(n20596), .A2(n20791), .B1(n20790), .B2(n20595), .ZN(
        n20594) );
  AOI22_X1 U23697 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20598), .B1(
        n20597), .B2(n20792), .ZN(n20593) );
  OAI211_X1 U23698 ( .C1(n20795), .C2(n20601), .A(n20594), .B(n20593), .ZN(
        P2_U3134) );
  AOI22_X1 U23699 ( .A1(n20596), .A2(n20798), .B1(n20797), .B2(n20595), .ZN(
        n20600) );
  AOI22_X1 U23700 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20598), .B1(
        n20597), .B2(n20800), .ZN(n20599) );
  OAI211_X1 U23701 ( .C1(n20806), .C2(n20601), .A(n20600), .B(n20599), .ZN(
        P2_U3135) );
  INV_X1 U23702 ( .A(n20602), .ZN(n20603) );
  NAND2_X1 U23703 ( .A1(n20604), .A2(n20603), .ZN(n20609) );
  AND2_X1 U23704 ( .A1(n20609), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n20605) );
  NAND2_X1 U23705 ( .A1(n20606), .A2(n20605), .ZN(n20610) );
  OAI21_X1 U23706 ( .B1(n20607), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n20742), 
        .ZN(n20608) );
  AND2_X1 U23707 ( .A1(n20610), .A2(n20608), .ZN(n20629) );
  INV_X1 U23708 ( .A(n20609), .ZN(n20628) );
  AOI22_X1 U23709 ( .A1(n20629), .A2(n20746), .B1(n20745), .B2(n20628), .ZN(
        n20615) );
  OAI211_X1 U23710 ( .C1(n20628), .C2(n20750), .A(n20610), .B(n20748), .ZN(
        n20611) );
  INV_X1 U23711 ( .A(n20611), .ZN(n20612) );
  OAI221_X1 U23712 ( .B1(n20613), .B2(n20885), .C1(n20613), .C2(n20753), .A(
        n20612), .ZN(n20630) );
  AOI22_X1 U23713 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20630), .B1(
        n20652), .B2(n20756), .ZN(n20614) );
  OAI211_X1 U23714 ( .C1(n20759), .C2(n20633), .A(n20615), .B(n20614), .ZN(
        P2_U3136) );
  AOI22_X1 U23715 ( .A1(n20629), .A2(n20761), .B1(n20760), .B2(n20628), .ZN(
        n20617) );
  AOI22_X1 U23716 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20630), .B1(
        n20652), .B2(n20762), .ZN(n20616) );
  OAI211_X1 U23717 ( .C1(n20765), .C2(n20633), .A(n20617), .B(n20616), .ZN(
        P2_U3137) );
  AOI22_X1 U23718 ( .A1(n20629), .A2(n20767), .B1(n20766), .B2(n20628), .ZN(
        n20619) );
  AOI22_X1 U23719 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20630), .B1(
        n20652), .B2(n20768), .ZN(n20618) );
  OAI211_X1 U23720 ( .C1(n20771), .C2(n20633), .A(n20619), .B(n20618), .ZN(
        P2_U3138) );
  AOI22_X1 U23721 ( .A1(n20629), .A2(n20773), .B1(n20772), .B2(n20628), .ZN(
        n20621) );
  AOI22_X1 U23722 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20630), .B1(
        n20652), .B2(n20774), .ZN(n20620) );
  OAI211_X1 U23723 ( .C1(n20777), .C2(n20633), .A(n20621), .B(n20620), .ZN(
        P2_U3139) );
  AOI22_X1 U23724 ( .A1(n20629), .A2(n20779), .B1(n20778), .B2(n20628), .ZN(
        n20623) );
  AOI22_X1 U23725 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20630), .B1(
        n20652), .B2(n20780), .ZN(n20622) );
  OAI211_X1 U23726 ( .C1(n20783), .C2(n20633), .A(n20623), .B(n20622), .ZN(
        P2_U3140) );
  AOI22_X1 U23727 ( .A1(n20629), .A2(n20785), .B1(n20784), .B2(n20628), .ZN(
        n20625) );
  AOI22_X1 U23728 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20630), .B1(
        n20652), .B2(n20786), .ZN(n20624) );
  OAI211_X1 U23729 ( .C1(n20789), .C2(n20633), .A(n20625), .B(n20624), .ZN(
        P2_U3141) );
  AOI22_X1 U23730 ( .A1(n20629), .A2(n20791), .B1(n20790), .B2(n20628), .ZN(
        n20627) );
  AOI22_X1 U23731 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20630), .B1(
        n20652), .B2(n20792), .ZN(n20626) );
  OAI211_X1 U23732 ( .C1(n20795), .C2(n20633), .A(n20627), .B(n20626), .ZN(
        P2_U3142) );
  AOI22_X1 U23733 ( .A1(n20629), .A2(n20798), .B1(n20797), .B2(n20628), .ZN(
        n20632) );
  AOI22_X1 U23734 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20630), .B1(
        n20652), .B2(n20800), .ZN(n20631) );
  OAI211_X1 U23735 ( .C1(n20806), .C2(n20633), .A(n20632), .B(n20631), .ZN(
        P2_U3143) );
  INV_X1 U23736 ( .A(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n20637) );
  AOI22_X1 U23737 ( .A1(n20651), .A2(n20767), .B1(n20650), .B2(n20766), .ZN(
        n20636) );
  AOI22_X1 U23738 ( .A1(n20686), .A2(n20768), .B1(n20652), .B2(n20634), .ZN(
        n20635) );
  OAI211_X1 U23739 ( .C1(n20656), .C2(n20637), .A(n20636), .B(n20635), .ZN(
        P2_U3146) );
  AOI22_X1 U23740 ( .A1(n20651), .A2(n20773), .B1(n20650), .B2(n20772), .ZN(
        n20640) );
  AOI22_X1 U23741 ( .A1(n20686), .A2(n20774), .B1(n20652), .B2(n20638), .ZN(
        n20639) );
  OAI211_X1 U23742 ( .C1(n20656), .C2(n10865), .A(n20640), .B(n20639), .ZN(
        P2_U3147) );
  INV_X1 U23743 ( .A(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n20644) );
  AOI22_X1 U23744 ( .A1(n20651), .A2(n20779), .B1(n20650), .B2(n20778), .ZN(
        n20643) );
  AOI22_X1 U23745 ( .A1(n20686), .A2(n20780), .B1(n20652), .B2(n20641), .ZN(
        n20642) );
  OAI211_X1 U23746 ( .C1(n20656), .C2(n20644), .A(n20643), .B(n20642), .ZN(
        P2_U3148) );
  AOI22_X1 U23747 ( .A1(n20651), .A2(n20785), .B1(n20650), .B2(n20784), .ZN(
        n20646) );
  AOI22_X1 U23748 ( .A1(n20686), .A2(n20786), .B1(n20652), .B2(n20678), .ZN(
        n20645) );
  OAI211_X1 U23749 ( .C1(n20656), .C2(n10922), .A(n20646), .B(n20645), .ZN(
        P2_U3149) );
  AOI22_X1 U23750 ( .A1(n20651), .A2(n20791), .B1(n20650), .B2(n20790), .ZN(
        n20649) );
  AOI22_X1 U23751 ( .A1(n20686), .A2(n20792), .B1(n20652), .B2(n20647), .ZN(
        n20648) );
  OAI211_X1 U23752 ( .C1(n20656), .C2(n10958), .A(n20649), .B(n20648), .ZN(
        P2_U3150) );
  INV_X1 U23753 ( .A(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n20655) );
  AOI22_X1 U23754 ( .A1(n20651), .A2(n20798), .B1(n20650), .B2(n20797), .ZN(
        n20654) );
  AOI22_X1 U23755 ( .A1(n20686), .A2(n20800), .B1(n20652), .B2(n20733), .ZN(
        n20653) );
  OAI211_X1 U23756 ( .C1(n20656), .C2(n20655), .A(n20654), .B(n20653), .ZN(
        P2_U3151) );
  NOR2_X1 U23757 ( .A1(n20741), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20665) );
  INV_X1 U23758 ( .A(n20665), .ZN(n20659) );
  NAND3_X1 U23759 ( .A1(n20909), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(
        n20694), .ZN(n20662) );
  INV_X1 U23760 ( .A(n20662), .ZN(n20684) );
  AOI211_X2 U23761 ( .C1(n20659), .C2(n20742), .A(n20658), .B(n20660), .ZN(
        n20685) );
  AOI22_X1 U23762 ( .A1(n20685), .A2(n20746), .B1(n20745), .B2(n20684), .ZN(
        n20669) );
  INV_X1 U23763 ( .A(n20666), .ZN(n20664) );
  AOI211_X1 U23764 ( .C1(P2_STATE2_REG_3__SCAN_IN), .C2(n20662), .A(n20661), 
        .B(n20660), .ZN(n20663) );
  OAI221_X1 U23765 ( .B1(n20665), .B2(n20664), .C1(n20665), .C2(n20753), .A(
        n20663), .ZN(n20687) );
  AOI22_X1 U23766 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20687), .B1(
        n20732), .B2(n20756), .ZN(n20668) );
  OAI211_X1 U23767 ( .C1(n20759), .C2(n20683), .A(n20669), .B(n20668), .ZN(
        P2_U3152) );
  AOI22_X1 U23768 ( .A1(n20685), .A2(n20761), .B1(n20760), .B2(n20684), .ZN(
        n20671) );
  AOI22_X1 U23769 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20687), .B1(
        n20686), .B2(n20705), .ZN(n20670) );
  OAI211_X1 U23770 ( .C1(n20708), .C2(n20730), .A(n20671), .B(n20670), .ZN(
        P2_U3153) );
  AOI22_X1 U23771 ( .A1(n20685), .A2(n20767), .B1(n20766), .B2(n20684), .ZN(
        n20673) );
  AOI22_X1 U23772 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20687), .B1(
        n20732), .B2(n20768), .ZN(n20672) );
  OAI211_X1 U23773 ( .C1(n20771), .C2(n20683), .A(n20673), .B(n20672), .ZN(
        P2_U3154) );
  AOI22_X1 U23774 ( .A1(n20685), .A2(n20773), .B1(n20772), .B2(n20684), .ZN(
        n20675) );
  AOI22_X1 U23775 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20687), .B1(
        n20732), .B2(n20774), .ZN(n20674) );
  OAI211_X1 U23776 ( .C1(n20777), .C2(n20683), .A(n20675), .B(n20674), .ZN(
        P2_U3155) );
  AOI22_X1 U23777 ( .A1(n20685), .A2(n20779), .B1(n20778), .B2(n20684), .ZN(
        n20677) );
  AOI22_X1 U23778 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20687), .B1(
        n20732), .B2(n20780), .ZN(n20676) );
  OAI211_X1 U23779 ( .C1(n20783), .C2(n20683), .A(n20677), .B(n20676), .ZN(
        P2_U3156) );
  AOI22_X1 U23780 ( .A1(n20685), .A2(n20785), .B1(n20784), .B2(n20684), .ZN(
        n20680) );
  AOI22_X1 U23781 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20687), .B1(
        n20686), .B2(n20678), .ZN(n20679) );
  OAI211_X1 U23782 ( .C1(n20720), .C2(n20730), .A(n20680), .B(n20679), .ZN(
        P2_U3157) );
  AOI22_X1 U23783 ( .A1(n20685), .A2(n20791), .B1(n20790), .B2(n20684), .ZN(
        n20682) );
  AOI22_X1 U23784 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20687), .B1(
        n20732), .B2(n20792), .ZN(n20681) );
  OAI211_X1 U23785 ( .C1(n20795), .C2(n20683), .A(n20682), .B(n20681), .ZN(
        P2_U3158) );
  AOI22_X1 U23786 ( .A1(n20685), .A2(n20798), .B1(n20797), .B2(n20684), .ZN(
        n20689) );
  AOI22_X1 U23787 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20687), .B1(
        n20686), .B2(n20733), .ZN(n20688) );
  OAI211_X1 U23788 ( .C1(n20738), .C2(n20730), .A(n20689), .B(n20688), .ZN(
        P2_U3159) );
  INV_X1 U23789 ( .A(n20805), .ZN(n20716) );
  AOI22_X1 U23790 ( .A1(n20756), .A2(n20716), .B1(n20745), .B2(n20731), .ZN(
        n20704) );
  AOI21_X1 U23791 ( .B1(n10869), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n20697) );
  AOI21_X1 U23792 ( .B1(n20730), .B2(n20805), .A(n20691), .ZN(n20693) );
  NOR2_X1 U23793 ( .A1(n20693), .A2(n20692), .ZN(n20698) );
  NAND2_X1 U23794 ( .A1(n20695), .A2(n20694), .ZN(n20701) );
  NAND2_X1 U23795 ( .A1(n20698), .A2(n20701), .ZN(n20696) );
  OAI211_X1 U23796 ( .C1(n20731), .C2(n20697), .A(n20696), .B(n20748), .ZN(
        n20735) );
  INV_X1 U23797 ( .A(n20698), .ZN(n20702) );
  INV_X1 U23798 ( .A(n10869), .ZN(n20699) );
  OAI21_X1 U23799 ( .B1(n20699), .B2(n20731), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20700) );
  OAI21_X2 U23800 ( .B1(n20702), .B2(n20701), .A(n20700), .ZN(n20734) );
  AOI22_X1 U23801 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20735), .B1(
        n20746), .B2(n20734), .ZN(n20703) );
  OAI211_X1 U23802 ( .C1(n20759), .C2(n20730), .A(n20704), .B(n20703), .ZN(
        P2_U3160) );
  AOI22_X1 U23803 ( .A1(n20705), .A2(n20732), .B1(n20760), .B2(n20731), .ZN(
        n20707) );
  AOI22_X1 U23804 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20735), .B1(
        n20761), .B2(n20734), .ZN(n20706) );
  OAI211_X1 U23805 ( .C1(n20708), .C2(n20805), .A(n20707), .B(n20706), .ZN(
        P2_U3161) );
  INV_X1 U23806 ( .A(n20731), .ZN(n20725) );
  OAI22_X1 U23807 ( .A1(n20730), .A2(n20771), .B1(n20709), .B2(n20725), .ZN(
        n20710) );
  INV_X1 U23808 ( .A(n20710), .ZN(n20712) );
  AOI22_X1 U23809 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20735), .B1(
        n20767), .B2(n20734), .ZN(n20711) );
  OAI211_X1 U23810 ( .C1(n20713), .C2(n20805), .A(n20712), .B(n20711), .ZN(
        P2_U3162) );
  AOI22_X1 U23811 ( .A1(n20774), .A2(n20716), .B1(n20772), .B2(n20731), .ZN(
        n20715) );
  AOI22_X1 U23812 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20735), .B1(
        n20773), .B2(n20734), .ZN(n20714) );
  OAI211_X1 U23813 ( .C1(n20777), .C2(n20730), .A(n20715), .B(n20714), .ZN(
        P2_U3163) );
  AOI22_X1 U23814 ( .A1(n20780), .A2(n20716), .B1(n20778), .B2(n20731), .ZN(
        n20718) );
  AOI22_X1 U23815 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20735), .B1(
        n20779), .B2(n20734), .ZN(n20717) );
  OAI211_X1 U23816 ( .C1(n20783), .C2(n20730), .A(n20718), .B(n20717), .ZN(
        P2_U3164) );
  OAI22_X1 U23817 ( .A1(n20805), .A2(n20720), .B1(n20725), .B2(n20719), .ZN(
        n20721) );
  INV_X1 U23818 ( .A(n20721), .ZN(n20723) );
  AOI22_X1 U23819 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20735), .B1(
        n20785), .B2(n20734), .ZN(n20722) );
  OAI211_X1 U23820 ( .C1(n20789), .C2(n20730), .A(n20723), .B(n20722), .ZN(
        P2_U3165) );
  OAI22_X1 U23821 ( .A1(n20805), .A2(n20726), .B1(n20725), .B2(n20724), .ZN(
        n20727) );
  INV_X1 U23822 ( .A(n20727), .ZN(n20729) );
  AOI22_X1 U23823 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20735), .B1(
        n20791), .B2(n20734), .ZN(n20728) );
  OAI211_X1 U23824 ( .C1(n20795), .C2(n20730), .A(n20729), .B(n20728), .ZN(
        P2_U3166) );
  AOI22_X1 U23825 ( .A1(n20733), .A2(n20732), .B1(n20797), .B2(n20731), .ZN(
        n20737) );
  AOI22_X1 U23826 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20735), .B1(
        n20798), .B2(n20734), .ZN(n20736) );
  OAI211_X1 U23827 ( .C1(n20738), .C2(n20805), .A(n20737), .B(n20736), .ZN(
        P2_U3167) );
  NOR2_X1 U23828 ( .A1(n20796), .A2(n20742), .ZN(n20739) );
  NAND2_X1 U23829 ( .A1(n20740), .A2(n20739), .ZN(n20749) );
  NOR2_X1 U23830 ( .A1(n20909), .A2(n20741), .ZN(n20755) );
  INV_X1 U23831 ( .A(n20755), .ZN(n20743) );
  OAI21_X1 U23832 ( .B1(n20743), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n20742), 
        .ZN(n20744) );
  AND2_X1 U23833 ( .A1(n20749), .A2(n20744), .ZN(n20799) );
  AOI22_X1 U23834 ( .A1(n20799), .A2(n20746), .B1(n20745), .B2(n20796), .ZN(
        n20758) );
  INV_X1 U23835 ( .A(n20747), .ZN(n20754) );
  OAI211_X1 U23836 ( .C1(n20796), .C2(n20750), .A(n20749), .B(n20748), .ZN(
        n20751) );
  INV_X1 U23837 ( .A(n20751), .ZN(n20752) );
  OAI221_X1 U23838 ( .B1(n20755), .B2(n20754), .C1(n20755), .C2(n20753), .A(
        n20752), .ZN(n20802) );
  AOI22_X1 U23839 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20802), .B1(
        n20801), .B2(n20756), .ZN(n20757) );
  OAI211_X1 U23840 ( .C1(n20759), .C2(n20805), .A(n20758), .B(n20757), .ZN(
        P2_U3168) );
  AOI22_X1 U23841 ( .A1(n20799), .A2(n20761), .B1(n20760), .B2(n20796), .ZN(
        n20764) );
  AOI22_X1 U23842 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20802), .B1(
        n20801), .B2(n20762), .ZN(n20763) );
  OAI211_X1 U23843 ( .C1(n20765), .C2(n20805), .A(n20764), .B(n20763), .ZN(
        P2_U3169) );
  AOI22_X1 U23844 ( .A1(n20799), .A2(n20767), .B1(n20766), .B2(n20796), .ZN(
        n20770) );
  AOI22_X1 U23845 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20802), .B1(
        n20801), .B2(n20768), .ZN(n20769) );
  OAI211_X1 U23846 ( .C1(n20771), .C2(n20805), .A(n20770), .B(n20769), .ZN(
        P2_U3170) );
  AOI22_X1 U23847 ( .A1(n20799), .A2(n20773), .B1(n20772), .B2(n20796), .ZN(
        n20776) );
  AOI22_X1 U23848 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20802), .B1(
        n20801), .B2(n20774), .ZN(n20775) );
  OAI211_X1 U23849 ( .C1(n20777), .C2(n20805), .A(n20776), .B(n20775), .ZN(
        P2_U3171) );
  AOI22_X1 U23850 ( .A1(n20799), .A2(n20779), .B1(n20778), .B2(n20796), .ZN(
        n20782) );
  AOI22_X1 U23851 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20802), .B1(
        n20801), .B2(n20780), .ZN(n20781) );
  OAI211_X1 U23852 ( .C1(n20783), .C2(n20805), .A(n20782), .B(n20781), .ZN(
        P2_U3172) );
  AOI22_X1 U23853 ( .A1(n20799), .A2(n20785), .B1(n20784), .B2(n20796), .ZN(
        n20788) );
  AOI22_X1 U23854 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20802), .B1(
        n20801), .B2(n20786), .ZN(n20787) );
  OAI211_X1 U23855 ( .C1(n20789), .C2(n20805), .A(n20788), .B(n20787), .ZN(
        P2_U3173) );
  AOI22_X1 U23856 ( .A1(n20799), .A2(n20791), .B1(n20790), .B2(n20796), .ZN(
        n20794) );
  AOI22_X1 U23857 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20802), .B1(
        n20801), .B2(n20792), .ZN(n20793) );
  OAI211_X1 U23858 ( .C1(n20795), .C2(n20805), .A(n20794), .B(n20793), .ZN(
        P2_U3174) );
  AOI22_X1 U23859 ( .A1(n20799), .A2(n20798), .B1(n20797), .B2(n20796), .ZN(
        n20804) );
  AOI22_X1 U23860 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20802), .B1(
        n20801), .B2(n20800), .ZN(n20803) );
  OAI211_X1 U23861 ( .C1(n20806), .C2(n20805), .A(n20804), .B(n20803), .ZN(
        P2_U3175) );
  AND2_X1 U23862 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n20881), .ZN(
        P2_U3179) );
  AND2_X1 U23863 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n20881), .ZN(
        P2_U3180) );
  AND2_X1 U23864 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n20881), .ZN(
        P2_U3181) );
  AND2_X1 U23865 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n20881), .ZN(
        P2_U3182) );
  INV_X1 U23866 ( .A(P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n21894) );
  NOR2_X1 U23867 ( .A1(n21894), .A2(n20884), .ZN(P2_U3183) );
  AND2_X1 U23868 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n20881), .ZN(
        P2_U3184) );
  AND2_X1 U23869 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n20881), .ZN(
        P2_U3185) );
  AND2_X1 U23870 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n20881), .ZN(
        P2_U3186) );
  AND2_X1 U23871 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n20881), .ZN(
        P2_U3187) );
  AND2_X1 U23872 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n20881), .ZN(
        P2_U3188) );
  AND2_X1 U23873 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n20881), .ZN(
        P2_U3189) );
  AND2_X1 U23874 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n20881), .ZN(
        P2_U3190) );
  AND2_X1 U23875 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n20881), .ZN(
        P2_U3191) );
  AND2_X1 U23876 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n20881), .ZN(
        P2_U3192) );
  AND2_X1 U23877 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n20881), .ZN(
        P2_U3193) );
  AND2_X1 U23878 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n20881), .ZN(
        P2_U3194) );
  AND2_X1 U23879 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n20881), .ZN(
        P2_U3195) );
  AND2_X1 U23880 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n20881), .ZN(
        P2_U3196) );
  AND2_X1 U23881 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n20881), .ZN(
        P2_U3197) );
  NOR2_X1 U23882 ( .A1(n21883), .A2(n20884), .ZN(P2_U3198) );
  AND2_X1 U23883 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n20881), .ZN(
        P2_U3199) );
  AND2_X1 U23884 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n20881), .ZN(
        P2_U3200) );
  AND2_X1 U23885 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n20881), .ZN(P2_U3201) );
  AND2_X1 U23886 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n20881), .ZN(P2_U3202) );
  AND2_X1 U23887 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n20881), .ZN(P2_U3203) );
  AND2_X1 U23888 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n20881), .ZN(P2_U3204) );
  AND2_X1 U23889 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n20881), .ZN(P2_U3205) );
  NOR2_X1 U23890 ( .A1(n21766), .A2(n20884), .ZN(P2_U3206) );
  AND2_X1 U23891 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n20881), .ZN(P2_U3207) );
  AND2_X1 U23892 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n20881), .ZN(P2_U3208) );
  NAND2_X1 U23893 ( .A1(n20819), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n20821) );
  NAND3_X1 U23894 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(
        P2_STATE_REG_0__SCAN_IN), .A3(n20821), .ZN(n20809) );
  AOI211_X1 U23895 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(n20817), .A(
        n20807), .B(n20930), .ZN(n20808) );
  NOR2_X1 U23896 ( .A1(n21536), .A2(n20813), .ZN(n20826) );
  AOI211_X1 U23897 ( .C1(n20827), .C2(n20809), .A(n20808), .B(n20826), .ZN(
        n20810) );
  INV_X1 U23898 ( .A(n20810), .ZN(P2_U3209) );
  INV_X1 U23899 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n20811) );
  AOI21_X1 U23900 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n20817), .A(n20827), 
        .ZN(n20818) );
  NOR2_X1 U23901 ( .A1(n20811), .A2(n20818), .ZN(n20814) );
  AOI21_X1 U23902 ( .B1(n20814), .B2(n20813), .A(n20812), .ZN(n20815) );
  OAI211_X1 U23903 ( .C1(n20817), .C2(n20816), .A(n20815), .B(n20821), .ZN(
        P2_U3210) );
  AOI21_X1 U23904 ( .B1(n20820), .B2(n20819), .A(n20818), .ZN(n20825) );
  OAI22_X1 U23905 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(n20822), .B1(NA), 
        .B2(n20821), .ZN(n20823) );
  OAI211_X1 U23906 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .B(n20823), .ZN(n20824) );
  OAI21_X1 U23907 ( .B1(n20826), .B2(n20825), .A(n20824), .ZN(P2_U3211) );
  OAI222_X1 U23908 ( .A1(n20873), .A2(n20829), .B1(n20828), .B2(n20930), .C1(
        n20830), .C2(n20876), .ZN(P2_U3212) );
  OAI222_X1 U23909 ( .A1(n20876), .A2(n17135), .B1(n20831), .B2(n20930), .C1(
        n20830), .C2(n20873), .ZN(P2_U3213) );
  OAI222_X1 U23910 ( .A1(n20876), .A2(n11396), .B1(n20832), .B2(n20930), .C1(
        n17135), .C2(n20873), .ZN(P2_U3214) );
  OAI222_X1 U23911 ( .A1(n20876), .A2(n16300), .B1(n20833), .B2(n20930), .C1(
        n11396), .C2(n20873), .ZN(P2_U3215) );
  OAI222_X1 U23912 ( .A1(n20876), .A2(n20835), .B1(n20834), .B2(n20930), .C1(
        n16300), .C2(n20873), .ZN(P2_U3216) );
  OAI222_X1 U23913 ( .A1(n20876), .A2(n20837), .B1(n20836), .B2(n20930), .C1(
        n20835), .C2(n20873), .ZN(P2_U3217) );
  OAI222_X1 U23914 ( .A1(n20876), .A2(n20839), .B1(n20838), .B2(n20930), .C1(
        n20837), .C2(n20873), .ZN(P2_U3218) );
  OAI222_X1 U23915 ( .A1(n20876), .A2(n20841), .B1(n20840), .B2(n20930), .C1(
        n20839), .C2(n20873), .ZN(P2_U3219) );
  OAI222_X1 U23916 ( .A1(n20876), .A2(n20843), .B1(n20842), .B2(n20930), .C1(
        n20841), .C2(n20873), .ZN(P2_U3220) );
  OAI222_X1 U23917 ( .A1(n20876), .A2(n11424), .B1(n20844), .B2(n20930), .C1(
        n20843), .C2(n20873), .ZN(P2_U3221) );
  OAI222_X1 U23918 ( .A1(n20876), .A2(n16227), .B1(n20845), .B2(n20930), .C1(
        n11424), .C2(n20873), .ZN(P2_U3222) );
  OAI222_X1 U23919 ( .A1(n20876), .A2(n20846), .B1(n21691), .B2(n20930), .C1(
        n16227), .C2(n20873), .ZN(P2_U3223) );
  OAI222_X1 U23920 ( .A1(n20876), .A2(n20848), .B1(n20847), .B2(n20930), .C1(
        n20846), .C2(n20873), .ZN(P2_U3224) );
  OAI222_X1 U23921 ( .A1(n20876), .A2(n20849), .B1(n21898), .B2(n20930), .C1(
        n20848), .C2(n20873), .ZN(P2_U3225) );
  OAI222_X1 U23922 ( .A1(n20876), .A2(n20851), .B1(n20850), .B2(n20930), .C1(
        n20849), .C2(n20873), .ZN(P2_U3226) );
  OAI222_X1 U23923 ( .A1(n20876), .A2(n20853), .B1(n20852), .B2(n20930), .C1(
        n20851), .C2(n20873), .ZN(P2_U3227) );
  OAI222_X1 U23924 ( .A1(n20876), .A2(n20855), .B1(n20854), .B2(n20930), .C1(
        n20853), .C2(n20873), .ZN(P2_U3228) );
  OAI222_X1 U23925 ( .A1(n20876), .A2(n21778), .B1(n20856), .B2(n20930), .C1(
        n20855), .C2(n20873), .ZN(P2_U3229) );
  OAI222_X1 U23926 ( .A1(n20876), .A2(n11462), .B1(n20857), .B2(n20930), .C1(
        n21778), .C2(n20873), .ZN(P2_U3230) );
  OAI222_X1 U23927 ( .A1(n20876), .A2(n20859), .B1(n20858), .B2(n20930), .C1(
        n11462), .C2(n20873), .ZN(P2_U3231) );
  OAI222_X1 U23928 ( .A1(n20876), .A2(n16949), .B1(n20860), .B2(n20930), .C1(
        n20859), .C2(n20873), .ZN(P2_U3232) );
  OAI222_X1 U23929 ( .A1(n20876), .A2(n20862), .B1(n20861), .B2(n20930), .C1(
        n16949), .C2(n20873), .ZN(P2_U3233) );
  OAI222_X1 U23930 ( .A1(n20876), .A2(n20864), .B1(n20863), .B2(n20930), .C1(
        n20862), .C2(n20873), .ZN(P2_U3234) );
  OAI222_X1 U23931 ( .A1(n20876), .A2(n20866), .B1(n20865), .B2(n20930), .C1(
        n20864), .C2(n20873), .ZN(P2_U3235) );
  OAI222_X1 U23932 ( .A1(n20876), .A2(n16906), .B1(n20867), .B2(n20930), .C1(
        n20866), .C2(n20873), .ZN(P2_U3236) );
  OAI222_X1 U23933 ( .A1(n20876), .A2(n20869), .B1(n21748), .B2(n20930), .C1(
        n16906), .C2(n20873), .ZN(P2_U3237) );
  INV_X1 U23934 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n20870) );
  OAI222_X1 U23935 ( .A1(n20873), .A2(n20869), .B1(n20868), .B2(n20930), .C1(
        n20870), .C2(n20876), .ZN(P2_U3238) );
  OAI222_X1 U23936 ( .A1(n20876), .A2(n20871), .B1(n21840), .B2(n20930), .C1(
        n20870), .C2(n20873), .ZN(P2_U3239) );
  OAI222_X1 U23937 ( .A1(n20876), .A2(n12838), .B1(n20872), .B2(n20930), .C1(
        n20871), .C2(n20873), .ZN(P2_U3240) );
  OAI222_X1 U23938 ( .A1(n20876), .A2(n20875), .B1(n20874), .B2(n20930), .C1(
        n12838), .C2(n20873), .ZN(P2_U3241) );
  OAI22_X1 U23939 ( .A1(n20931), .A2(P2_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P2_BE_N_REG_3__SCAN_IN), .B2(n20930), .ZN(n20877) );
  INV_X1 U23940 ( .A(n20877), .ZN(P2_U3585) );
  MUX2_X1 U23941 ( .A(P2_BYTEENABLE_REG_2__SCAN_IN), .B(P2_BE_N_REG_2__SCAN_IN), .S(n20931), .Z(P2_U3586) );
  OAI22_X1 U23942 ( .A1(n20931), .A2(P2_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P2_BE_N_REG_1__SCAN_IN), .B2(n20930), .ZN(n20878) );
  INV_X1 U23943 ( .A(n20878), .ZN(P2_U3587) );
  OAI22_X1 U23944 ( .A1(n20931), .A2(P2_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P2_BE_N_REG_0__SCAN_IN), .B2(n20930), .ZN(n20879) );
  INV_X1 U23945 ( .A(n20879), .ZN(P2_U3588) );
  AOI21_X1 U23946 ( .B1(n20881), .B2(n21711), .A(n20880), .ZN(P2_U3591) );
  OAI21_X1 U23947 ( .B1(n20884), .B2(n20883), .A(n20882), .ZN(P2_U3592) );
  NAND2_X1 U23948 ( .A1(n20885), .A2(n20905), .ZN(n20893) );
  NAND2_X1 U23949 ( .A1(n20903), .A2(n20902), .ZN(n20886) );
  NAND2_X1 U23950 ( .A1(n20886), .A2(n20901), .ZN(n20895) );
  NAND2_X1 U23951 ( .A1(n20893), .A2(n20895), .ZN(n20891) );
  AOI222_X1 U23952 ( .A1(n20891), .A2(n20890), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(n20889), .C1(n20888), .C2(n20887), .ZN(n20892) );
  AOI22_X1 U23953 ( .A1(n20917), .A2(n21853), .B1(n20892), .B2(n20918), .ZN(
        P2_U3602) );
  INV_X1 U23954 ( .A(n20893), .ZN(n20898) );
  OAI22_X1 U23955 ( .A1(n20896), .A2(n20895), .B1(n20894), .B2(n20750), .ZN(
        n20897) );
  NOR2_X1 U23956 ( .A1(n20898), .A2(n20897), .ZN(n20899) );
  AOI22_X1 U23957 ( .A1(n20917), .A2(n20900), .B1(n20899), .B2(n20918), .ZN(
        P2_U3603) );
  INV_X1 U23958 ( .A(n20901), .ZN(n20913) );
  NOR2_X1 U23959 ( .A1(n20913), .A2(n20902), .ZN(n20904) );
  MUX2_X1 U23960 ( .A(n20905), .B(n20904), .S(n20903), .Z(n20906) );
  AOI21_X1 U23961 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n20907), .A(n20906), 
        .ZN(n20908) );
  AOI22_X1 U23962 ( .A1(n20917), .A2(n20909), .B1(n20908), .B2(n20918), .ZN(
        P2_U3604) );
  INV_X1 U23963 ( .A(n20910), .ZN(n20912) );
  OAI22_X1 U23964 ( .A1(n20914), .A2(n20913), .B1(n20912), .B2(n20911), .ZN(
        n20915) );
  AOI21_X1 U23965 ( .B1(n20919), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n20915), 
        .ZN(n20916) );
  OAI22_X1 U23966 ( .A1(n20919), .A2(n20918), .B1(n20917), .B2(n20916), .ZN(
        P2_U3605) );
  INV_X1 U23967 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n20920) );
  AOI22_X1 U23968 ( .A1(n20930), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n20920), 
        .B2(n20931), .ZN(P2_U3608) );
  INV_X1 U23969 ( .A(n20921), .ZN(n20926) );
  NAND2_X1 U23970 ( .A1(n20923), .A2(n20922), .ZN(n20924) );
  OAI211_X1 U23971 ( .C1(n20927), .C2(n20926), .A(n20925), .B(n20924), .ZN(
        n20929) );
  MUX2_X1 U23972 ( .A(P2_MORE_REG_SCAN_IN), .B(n20929), .S(n20928), .Z(
        P2_U3609) );
  OAI22_X1 U23973 ( .A1(n20931), .A2(P2_MEMORYFETCH_REG_SCAN_IN), .B1(
        P2_M_IO_N_REG_SCAN_IN), .B2(n20930), .ZN(n20932) );
  INV_X1 U23974 ( .A(n20932), .ZN(P2_U3611) );
  AND2_X1 U23975 ( .A1(n21531), .A2(P1_STATE_REG_0__SCAN_IN), .ZN(n20934) );
  INV_X1 U23976 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n20933) );
  AOI21_X1 U23977 ( .B1(n20934), .B2(n20933), .A(n21625), .ZN(P1_U2802) );
  INV_X1 U23978 ( .A(n20935), .ZN(n20936) );
  OAI21_X1 U23979 ( .B1(n20937), .B2(n20936), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n20938) );
  OAI21_X1 U23980 ( .B1(n20940), .B2(n20939), .A(n20938), .ZN(P1_U2803) );
  NOR2_X1 U23981 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n20942) );
  OAI21_X1 U23982 ( .B1(n20942), .B2(P1_D_C_N_REG_SCAN_IN), .A(n21623), .ZN(
        n20941) );
  OAI21_X1 U23983 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n21623), .A(n20941), 
        .ZN(P1_U2804) );
  AOI21_X1 U23984 ( .B1(P1_STATE_REG_0__SCAN_IN), .B2(n21531), .A(n21625), 
        .ZN(n21591) );
  OAI21_X1 U23985 ( .B1(BS16), .B2(n20942), .A(n21591), .ZN(n21589) );
  OAI21_X1 U23986 ( .B1(n21591), .B2(n21468), .A(n21589), .ZN(P1_U2805) );
  OAI21_X1 U23987 ( .B1(n20945), .B2(n20944), .A(n20943), .ZN(P1_U2806) );
  NOR4_X1 U23988 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_20__SCAN_IN), .A3(P1_DATAWIDTH_REG_21__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_22__SCAN_IN), .ZN(n20949) );
  NOR4_X1 U23989 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_16__SCAN_IN), .A3(P1_DATAWIDTH_REG_17__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_18__SCAN_IN), .ZN(n20948) );
  NOR4_X1 U23990 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_28__SCAN_IN), .A3(P1_DATAWIDTH_REG_29__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n20947) );
  NOR4_X1 U23991 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_24__SCAN_IN), .A3(P1_DATAWIDTH_REG_25__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_26__SCAN_IN), .ZN(n20946) );
  NAND4_X1 U23992 ( .A1(n20949), .A2(n20948), .A3(n20947), .A4(n20946), .ZN(
        n20955) );
  NOR4_X1 U23993 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_3__SCAN_IN), .A3(P1_DATAWIDTH_REG_4__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_5__SCAN_IN), .ZN(n20953) );
  AOI211_X1 U23994 ( .C1(P1_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_12__SCAN_IN), .B(
        P1_DATAWIDTH_REG_30__SCAN_IN), .ZN(n20952) );
  NOR4_X1 U23995 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_11__SCAN_IN), .A3(P1_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_14__SCAN_IN), .ZN(n20951) );
  NOR4_X1 U23996 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_7__SCAN_IN), .A3(P1_DATAWIDTH_REG_8__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_9__SCAN_IN), .ZN(n20950) );
  NAND4_X1 U23997 ( .A1(n20953), .A2(n20952), .A3(n20951), .A4(n20950), .ZN(
        n20954) );
  NOR2_X1 U23998 ( .A1(n20955), .A2(n20954), .ZN(n21610) );
  INV_X1 U23999 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20957) );
  NOR3_X1 U24000 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n20958) );
  OAI21_X1 U24001 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n20958), .A(n21610), .ZN(
        n20956) );
  OAI21_X1 U24002 ( .B1(n21610), .B2(n20957), .A(n20956), .ZN(P1_U2807) );
  INV_X1 U24003 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n21590) );
  AOI21_X1 U24004 ( .B1(n21603), .B2(n21590), .A(n20958), .ZN(n20960) );
  INV_X1 U24005 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20959) );
  INV_X1 U24006 ( .A(n21610), .ZN(n21605) );
  AOI22_X1 U24007 ( .A1(n21610), .A2(n20960), .B1(n20959), .B2(n21605), .ZN(
        P1_U2808) );
  NOR2_X1 U24008 ( .A1(n20999), .A2(n20961), .ZN(n20994) );
  NAND3_X1 U24009 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .A3(n20994), .ZN(n20965) );
  INV_X1 U24010 ( .A(n20962), .ZN(n20963) );
  AOI22_X1 U24011 ( .A1(n21024), .A2(P1_EBX_REG_7__SCAN_IN), .B1(n20992), .B2(
        n20963), .ZN(n20964) );
  OAI21_X1 U24012 ( .B1(P1_REIP_REG_7__SCAN_IN), .B2(n20965), .A(n20964), .ZN(
        n20966) );
  AOI211_X1 U24013 ( .C1(n21019), .C2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n21009), .B(n20966), .ZN(n20973) );
  NAND2_X1 U24014 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .ZN(n20969) );
  NAND2_X1 U24015 ( .A1(n20970), .A2(n20969), .ZN(n20980) );
  NAND2_X1 U24016 ( .A1(n21011), .A2(n20980), .ZN(n20975) );
  AOI22_X1 U24017 ( .A1(n20971), .A2(n20982), .B1(P1_REIP_REG_7__SCAN_IN), 
        .B2(n20975), .ZN(n20972) );
  OAI211_X1 U24018 ( .C1(n20974), .C2(n21015), .A(n20973), .B(n20972), .ZN(
        P1_U2833) );
  NAND2_X1 U24019 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(n21011), .ZN(n20993) );
  AOI22_X1 U24020 ( .A1(n20992), .A2(n20976), .B1(P1_REIP_REG_6__SCAN_IN), 
        .B2(n20975), .ZN(n20977) );
  OAI211_X1 U24021 ( .C1(n21001), .C2(n10142), .A(n20977), .B(n20986), .ZN(
        n20978) );
  AOI21_X1 U24022 ( .B1(n21024), .B2(P1_EBX_REG_6__SCAN_IN), .A(n20978), .ZN(
        n20979) );
  OAI21_X1 U24023 ( .B1(n20980), .B2(n20993), .A(n20979), .ZN(n20981) );
  AOI21_X1 U24024 ( .B1(n20983), .B2(n20982), .A(n20981), .ZN(n20984) );
  OAI21_X1 U24025 ( .B1(n20985), .B2(n21015), .A(n20984), .ZN(P1_U2834) );
  INV_X1 U24026 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n21909) );
  NAND2_X1 U24027 ( .A1(n21024), .A2(P1_EBX_REG_5__SCAN_IN), .ZN(n20987) );
  OAI211_X1 U24028 ( .C1(n21001), .C2(n21909), .A(n20987), .B(n20986), .ZN(
        n20990) );
  NOR2_X1 U24029 ( .A1(n21010), .A2(n20988), .ZN(n20989) );
  AOI211_X1 U24030 ( .C1(n20992), .C2(n20991), .A(n20990), .B(n20989), .ZN(
        n20996) );
  OAI21_X1 U24031 ( .B1(P1_REIP_REG_5__SCAN_IN), .B2(n20994), .A(n20993), .ZN(
        n20995) );
  OAI211_X1 U24032 ( .C1(n21015), .C2(n20997), .A(n20996), .B(n20995), .ZN(
        P1_U2835) );
  NAND3_X1 U24033 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(P1_REIP_REG_1__SCAN_IN), 
        .A3(P1_REIP_REG_2__SCAN_IN), .ZN(n20998) );
  NOR3_X1 U24034 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(n20999), .A3(n20998), .ZN(
        n21008) );
  INV_X1 U24035 ( .A(n21000), .ZN(n21002) );
  OAI22_X1 U24036 ( .A1(n21002), .A2(n21021), .B1(n12057), .B2(n21001), .ZN(
        n21007) );
  OAI22_X1 U24037 ( .A1(n21026), .A2(n21005), .B1(n21004), .B2(n21003), .ZN(
        n21006) );
  NOR4_X1 U24038 ( .A1(n21009), .A2(n21008), .A3(n21007), .A4(n21006), .ZN(
        n21014) );
  INV_X1 U24039 ( .A(n21010), .ZN(n21018) );
  INV_X1 U24040 ( .A(n21011), .ZN(n21012) );
  AOI22_X1 U24041 ( .A1(n21018), .A2(n21093), .B1(n21012), .B2(
        P1_REIP_REG_4__SCAN_IN), .ZN(n21013) );
  OAI211_X1 U24042 ( .C1(n21099), .C2(n21015), .A(n21014), .B(n21013), .ZN(
        P1_U2836) );
  NAND2_X1 U24043 ( .A1(n21016), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n21029) );
  NAND2_X1 U24044 ( .A1(n21019), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n21020) );
  OAI21_X1 U24045 ( .B1(n21022), .B2(n21021), .A(n21020), .ZN(n21023) );
  AOI21_X1 U24046 ( .B1(n21024), .B2(P1_EBX_REG_2__SCAN_IN), .A(n21023), .ZN(
        n21025) );
  AOI22_X1 U24047 ( .A1(P1_EAX_REG_15__SCAN_IN), .A2(n21035), .B1(n21053), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n21031) );
  OAI21_X1 U24048 ( .B1(n21032), .B2(n21615), .A(n21031), .ZN(P1_U2921) );
  INV_X1 U24049 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n21034) );
  AOI22_X1 U24050 ( .A1(P1_LWORD_REG_14__SCAN_IN), .A2(n21054), .B1(n21053), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n21033) );
  OAI21_X1 U24051 ( .B1(n21034), .B2(n21060), .A(n21033), .ZN(P1_U2922) );
  INV_X1 U24052 ( .A(P1_LWORD_REG_13__SCAN_IN), .ZN(n21837) );
  AOI22_X1 U24053 ( .A1(P1_EAX_REG_13__SCAN_IN), .A2(n21035), .B1(n21053), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n21036) );
  OAI21_X1 U24054 ( .B1(n21837), .B2(n21615), .A(n21036), .ZN(P1_U2923) );
  AOI22_X1 U24055 ( .A1(P1_LWORD_REG_12__SCAN_IN), .A2(n21054), .B1(n21053), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n21037) );
  OAI21_X1 U24056 ( .B1(n15284), .B2(n21060), .A(n21037), .ZN(P1_U2924) );
  INV_X1 U24057 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n21039) );
  AOI22_X1 U24058 ( .A1(P1_LWORD_REG_11__SCAN_IN), .A2(n21054), .B1(n21053), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n21038) );
  OAI21_X1 U24059 ( .B1(n21039), .B2(n21060), .A(n21038), .ZN(P1_U2925) );
  AOI22_X1 U24060 ( .A1(P1_LWORD_REG_10__SCAN_IN), .A2(n21054), .B1(n21053), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n21040) );
  OAI21_X1 U24061 ( .B1(n15290), .B2(n21060), .A(n21040), .ZN(P1_U2926) );
  AOI22_X1 U24062 ( .A1(P1_LWORD_REG_9__SCAN_IN), .A2(n21054), .B1(n21053), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n21041) );
  OAI21_X1 U24063 ( .B1(n15291), .B2(n21060), .A(n21041), .ZN(P1_U2927) );
  AOI22_X1 U24064 ( .A1(P1_LWORD_REG_8__SCAN_IN), .A2(n21054), .B1(n21053), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n21042) );
  OAI21_X1 U24065 ( .B1(n21043), .B2(n21060), .A(n21042), .ZN(P1_U2928) );
  INV_X1 U24066 ( .A(P1_LWORD_REG_7__SCAN_IN), .ZN(n21893) );
  OAI222_X1 U24067 ( .A1(n21058), .A2(n21747), .B1(n21060), .B2(n12052), .C1(
        n21615), .C2(n21893), .ZN(P1_U2929) );
  AOI22_X1 U24068 ( .A1(P1_LWORD_REG_6__SCAN_IN), .A2(n21054), .B1(n21053), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n21044) );
  OAI21_X1 U24069 ( .B1(n21045), .B2(n21060), .A(n21044), .ZN(P1_U2930) );
  AOI22_X1 U24070 ( .A1(P1_LWORD_REG_5__SCAN_IN), .A2(n21054), .B1(n21053), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n21046) );
  OAI21_X1 U24071 ( .B1(n12116), .B2(n21060), .A(n21046), .ZN(P1_U2931) );
  AOI22_X1 U24072 ( .A1(P1_LWORD_REG_4__SCAN_IN), .A2(n21054), .B1(n21053), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n21047) );
  OAI21_X1 U24073 ( .B1(n21048), .B2(n21060), .A(n21047), .ZN(P1_U2932) );
  AOI22_X1 U24074 ( .A1(P1_LWORD_REG_3__SCAN_IN), .A2(n21054), .B1(n21053), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n21049) );
  OAI21_X1 U24075 ( .B1(n21050), .B2(n21060), .A(n21049), .ZN(P1_U2933) );
  AOI22_X1 U24076 ( .A1(P1_LWORD_REG_2__SCAN_IN), .A2(n21054), .B1(n21053), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n21051) );
  OAI21_X1 U24077 ( .B1(n21052), .B2(n21060), .A(n21051), .ZN(P1_U2934) );
  AOI22_X1 U24078 ( .A1(P1_LWORD_REG_1__SCAN_IN), .A2(n21054), .B1(n21053), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n21055) );
  OAI21_X1 U24079 ( .B1(n21056), .B2(n21060), .A(n21055), .ZN(P1_U2935) );
  INV_X1 U24080 ( .A(P1_LWORD_REG_0__SCAN_IN), .ZN(n21866) );
  OAI222_X1 U24081 ( .A1(n21615), .A2(n21866), .B1(n21060), .B2(n21059), .C1(
        n21058), .C2(n21057), .ZN(P1_U2936) );
  AOI22_X1 U24082 ( .A1(n21084), .A2(P1_EAX_REG_26__SCAN_IN), .B1(
        P1_UWORD_REG_10__SCAN_IN), .B2(n21077), .ZN(n21063) );
  INV_X1 U24083 ( .A(n21061), .ZN(n21062) );
  NAND2_X1 U24084 ( .A1(n21071), .A2(n21062), .ZN(n21075) );
  NAND2_X1 U24085 ( .A1(n21063), .A2(n21075), .ZN(P1_U2947) );
  AOI22_X1 U24086 ( .A1(n21084), .A2(P1_EAX_REG_27__SCAN_IN), .B1(
        P1_UWORD_REG_11__SCAN_IN), .B2(n21077), .ZN(n21065) );
  NAND2_X1 U24087 ( .A1(n21071), .A2(n21064), .ZN(n21078) );
  NAND2_X1 U24088 ( .A1(n21065), .A2(n21078), .ZN(P1_U2948) );
  AOI22_X1 U24089 ( .A1(n21084), .A2(P1_EAX_REG_29__SCAN_IN), .B1(
        P1_UWORD_REG_13__SCAN_IN), .B2(n21077), .ZN(n21068) );
  INV_X1 U24090 ( .A(n21066), .ZN(n21067) );
  NAND2_X1 U24091 ( .A1(n21071), .A2(n21067), .ZN(n21082) );
  NAND2_X1 U24092 ( .A1(n21068), .A2(n21082), .ZN(P1_U2950) );
  AOI22_X1 U24093 ( .A1(n21084), .A2(P1_EAX_REG_30__SCAN_IN), .B1(
        P1_UWORD_REG_14__SCAN_IN), .B2(n21077), .ZN(n21072) );
  INV_X1 U24094 ( .A(n21069), .ZN(n21070) );
  NAND2_X1 U24095 ( .A1(n21071), .A2(n21070), .ZN(n21085) );
  NAND2_X1 U24096 ( .A1(n21072), .A2(n21085), .ZN(P1_U2951) );
  AOI22_X1 U24097 ( .A1(n21084), .A2(P1_EAX_REG_9__SCAN_IN), .B1(
        P1_LWORD_REG_9__SCAN_IN), .B2(n21077), .ZN(n21074) );
  NAND2_X1 U24098 ( .A1(n21074), .A2(n21073), .ZN(P1_U2961) );
  AOI22_X1 U24099 ( .A1(n21084), .A2(P1_EAX_REG_10__SCAN_IN), .B1(
        P1_LWORD_REG_10__SCAN_IN), .B2(n21077), .ZN(n21076) );
  NAND2_X1 U24100 ( .A1(n21076), .A2(n21075), .ZN(P1_U2962) );
  AOI22_X1 U24101 ( .A1(n21084), .A2(P1_EAX_REG_11__SCAN_IN), .B1(
        P1_LWORD_REG_11__SCAN_IN), .B2(n21077), .ZN(n21079) );
  NAND2_X1 U24102 ( .A1(n21079), .A2(n21078), .ZN(P1_U2963) );
  AOI22_X1 U24103 ( .A1(n21084), .A2(P1_EAX_REG_12__SCAN_IN), .B1(
        P1_LWORD_REG_12__SCAN_IN), .B2(n21077), .ZN(n21081) );
  NAND2_X1 U24104 ( .A1(n21081), .A2(n21080), .ZN(P1_U2964) );
  AOI22_X1 U24105 ( .A1(n21084), .A2(P1_EAX_REG_13__SCAN_IN), .B1(
        P1_LWORD_REG_13__SCAN_IN), .B2(n21077), .ZN(n21083) );
  NAND2_X1 U24106 ( .A1(n21083), .A2(n21082), .ZN(P1_U2965) );
  AOI22_X1 U24107 ( .A1(n21084), .A2(P1_EAX_REG_14__SCAN_IN), .B1(
        P1_LWORD_REG_14__SCAN_IN), .B2(n21077), .ZN(n21086) );
  NAND2_X1 U24108 ( .A1(n21086), .A2(n21085), .ZN(P1_U2966) );
  INV_X1 U24109 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n21087) );
  NOR2_X1 U24110 ( .A1(n21123), .A2(n21087), .ZN(n21102) );
  AOI21_X1 U24111 ( .B1(n21088), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n21102), .ZN(n21097) );
  AOI21_X1 U24112 ( .B1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n15500), .A(
        n21089), .ZN(n21092) );
  XNOR2_X1 U24113 ( .A(n21090), .B(n10109), .ZN(n21091) );
  XNOR2_X1 U24114 ( .A(n21092), .B(n21091), .ZN(n21106) );
  AOI22_X1 U24115 ( .A1(n21106), .A2(n21095), .B1(n21094), .B2(n21093), .ZN(
        n21096) );
  OAI211_X1 U24116 ( .C1(n21099), .C2(n21098), .A(n21097), .B(n21096), .ZN(
        P1_U2995) );
  NOR2_X1 U24117 ( .A1(n21117), .A2(n21100), .ZN(n21127) );
  AOI211_X1 U24118 ( .C1(n21121), .C2(n21101), .A(n21127), .B(n21119), .ZN(
        n21113) );
  AOI21_X1 U24119 ( .B1(n21135), .B2(n21103), .A(n21102), .ZN(n21108) );
  AOI211_X1 U24120 ( .C1(n10109), .C2(n21114), .A(n21104), .B(n21115), .ZN(
        n21105) );
  AOI21_X1 U24121 ( .B1(n21106), .B2(n21110), .A(n21105), .ZN(n21107) );
  OAI211_X1 U24122 ( .C1(n21113), .C2(n10109), .A(n21108), .B(n21107), .ZN(
        P1_U3027) );
  AOI222_X1 U24123 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(n15496), .B1(n21135), 
        .B2(n21111), .C1(n21110), .C2(n21109), .ZN(n21112) );
  OAI221_X1 U24124 ( .B1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n21115), .C1(
        n21114), .C2(n21113), .A(n21112), .ZN(P1_U3028) );
  OR2_X1 U24125 ( .A1(n21144), .A2(n21116), .ZN(n21132) );
  NOR3_X1 U24126 ( .A1(n21118), .A2(n21144), .A3(n21117), .ZN(n21120) );
  AOI211_X1 U24127 ( .C1(n21144), .C2(n21121), .A(n21120), .B(n21119), .ZN(
        n21130) );
  NOR2_X1 U24128 ( .A1(n21122), .A2(n21139), .ZN(n21128) );
  OAI22_X1 U24129 ( .A1(n21125), .A2(n21124), .B1(n14277), .B2(n21123), .ZN(
        n21126) );
  AOI211_X1 U24130 ( .C1(n21128), .C2(n14275), .A(n21127), .B(n21126), .ZN(
        n21129) );
  OAI221_X1 U24131 ( .B1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n21132), .C1(
        n21131), .C2(n21130), .A(n21129), .ZN(P1_U3029) );
  AOI21_X1 U24132 ( .B1(n21135), .B2(n21134), .A(n21133), .ZN(n21143) );
  NAND3_X1 U24133 ( .A1(n21137), .A2(n21144), .A3(n21136), .ZN(n21138) );
  OAI21_X1 U24134 ( .B1(n21140), .B2(n21139), .A(n21138), .ZN(n21141) );
  INV_X1 U24135 ( .A(n21141), .ZN(n21142) );
  OAI211_X1 U24136 ( .C1(n21145), .C2(n21144), .A(n21143), .B(n21142), .ZN(
        P1_U3030) );
  NOR2_X1 U24137 ( .A1(n21147), .A2(n21146), .ZN(P1_U3032) );
  OAI22_X1 U24138 ( .A1(n21167), .A2(n21486), .B1(n21166), .B2(n21313), .ZN(
        n21148) );
  INV_X1 U24139 ( .A(n21148), .ZN(n21150) );
  AOI22_X1 U24140 ( .A1(n21482), .A2(n21170), .B1(n21169), .B2(n21483), .ZN(
        n21149) );
  OAI211_X1 U24141 ( .C1(n21173), .C2(n11812), .A(n21150), .B(n21149), .ZN(
        P1_U3034) );
  OAI22_X1 U24142 ( .A1(n21167), .A2(n21490), .B1(n21166), .B2(n21317), .ZN(
        n21151) );
  INV_X1 U24143 ( .A(n21151), .ZN(n21153) );
  INV_X1 U24144 ( .A(n21936), .ZN(n21487) );
  AOI22_X1 U24145 ( .A1(n21487), .A2(n21170), .B1(n21169), .B2(n21931), .ZN(
        n21152) );
  OAI211_X1 U24146 ( .C1(n21173), .C2(n21154), .A(n21153), .B(n21152), .ZN(
        P1_U3035) );
  INV_X1 U24147 ( .A(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n21158) );
  OAI22_X1 U24148 ( .A1(n21167), .A2(n21496), .B1(n21166), .B2(n21321), .ZN(
        n21155) );
  INV_X1 U24149 ( .A(n21155), .ZN(n21157) );
  AOI22_X1 U24150 ( .A1(n21492), .A2(n21170), .B1(n21169), .B2(n21493), .ZN(
        n21156) );
  OAI211_X1 U24151 ( .C1(n21173), .C2(n21158), .A(n21157), .B(n21156), .ZN(
        P1_U3036) );
  OAI22_X1 U24152 ( .A1(n21167), .A2(n21502), .B1(n21166), .B2(n21325), .ZN(
        n21159) );
  INV_X1 U24153 ( .A(n21159), .ZN(n21161) );
  INV_X1 U24154 ( .A(n21403), .ZN(n21498) );
  AOI22_X1 U24155 ( .A1(n21498), .A2(n21170), .B1(n21169), .B2(n21499), .ZN(
        n21160) );
  OAI211_X1 U24156 ( .C1(n21173), .C2(n21162), .A(n21161), .B(n21160), .ZN(
        P1_U3037) );
  OAI22_X1 U24157 ( .A1(n21167), .A2(n21508), .B1(n21166), .B2(n21329), .ZN(
        n21163) );
  INV_X1 U24158 ( .A(n21163), .ZN(n21165) );
  INV_X1 U24159 ( .A(n21406), .ZN(n21504) );
  AOI22_X1 U24160 ( .A1(n21504), .A2(n21170), .B1(n21169), .B2(n21505), .ZN(
        n21164) );
  OAI211_X1 U24161 ( .C1(n21173), .C2(n12018), .A(n21165), .B(n21164), .ZN(
        P1_U3038) );
  OAI22_X1 U24162 ( .A1(n21167), .A2(n21525), .B1(n21166), .B2(n21337), .ZN(
        n21168) );
  INV_X1 U24163 ( .A(n21168), .ZN(n21172) );
  INV_X1 U24164 ( .A(n21412), .ZN(n21517) );
  AOI22_X1 U24165 ( .A1(n21517), .A2(n21170), .B1(n21169), .B2(n21519), .ZN(
        n21171) );
  OAI211_X1 U24166 ( .C1(n21173), .C2(n12046), .A(n21172), .B(n21171), .ZN(
        P1_U3040) );
  INV_X1 U24167 ( .A(n21174), .ZN(n21347) );
  NOR2_X1 U24168 ( .A1(n21240), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n21180) );
  INV_X1 U24169 ( .A(n21180), .ZN(n21176) );
  NOR2_X1 U24170 ( .A1(n21414), .A2(n21176), .ZN(n21196) );
  AOI21_X1 U24171 ( .B1(n21175), .B2(n21347), .A(n21196), .ZN(n21177) );
  OAI22_X1 U24172 ( .A1(n21177), .A2(n21417), .B1(n21176), .B2(n21349), .ZN(
        n21197) );
  AOI22_X1 U24173 ( .A1(n21197), .A2(n21466), .B1(n21465), .B2(n21196), .ZN(
        n21183) );
  INV_X1 U24174 ( .A(n21233), .ZN(n21178) );
  OAI21_X1 U24175 ( .B1(n21178), .B2(n21468), .A(n21177), .ZN(n21179) );
  OAI221_X1 U24176 ( .B1(n21376), .B2(n21180), .C1(n21417), .C2(n21179), .A(
        n21422), .ZN(n21198) );
  AOI22_X1 U24177 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n21198), .B1(
        n21226), .B2(n21477), .ZN(n21182) );
  OAI211_X1 U24178 ( .C1(n21480), .C2(n21201), .A(n21183), .B(n21182), .ZN(
        P1_U3041) );
  AOI22_X1 U24179 ( .A1(n21197), .A2(n21482), .B1(n21481), .B2(n21196), .ZN(
        n21185) );
  AOI22_X1 U24180 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n21198), .B1(
        n21226), .B2(n21483), .ZN(n21184) );
  OAI211_X1 U24181 ( .C1(n21486), .C2(n21201), .A(n21185), .B(n21184), .ZN(
        P1_U3042) );
  AOI22_X1 U24182 ( .A1(n21197), .A2(n21487), .B1(n21928), .B2(n21196), .ZN(
        n21187) );
  AOI22_X1 U24183 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n21198), .B1(
        n21226), .B2(n21931), .ZN(n21186) );
  OAI211_X1 U24184 ( .C1(n21490), .C2(n21201), .A(n21187), .B(n21186), .ZN(
        P1_U3043) );
  AOI22_X1 U24185 ( .A1(n21197), .A2(n21492), .B1(n21491), .B2(n21196), .ZN(
        n21189) );
  AOI22_X1 U24186 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n21198), .B1(
        n21226), .B2(n21493), .ZN(n21188) );
  OAI211_X1 U24187 ( .C1(n21496), .C2(n21201), .A(n21189), .B(n21188), .ZN(
        P1_U3044) );
  AOI22_X1 U24188 ( .A1(n21197), .A2(n21498), .B1(n21497), .B2(n21196), .ZN(
        n21191) );
  AOI22_X1 U24189 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n21198), .B1(
        n21226), .B2(n21499), .ZN(n21190) );
  OAI211_X1 U24190 ( .C1(n21502), .C2(n21201), .A(n21191), .B(n21190), .ZN(
        P1_U3045) );
  AOI22_X1 U24191 ( .A1(n21197), .A2(n21504), .B1(n21503), .B2(n21196), .ZN(
        n21193) );
  AOI22_X1 U24192 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n21198), .B1(
        n21226), .B2(n21505), .ZN(n21192) );
  OAI211_X1 U24193 ( .C1(n21508), .C2(n21201), .A(n21193), .B(n21192), .ZN(
        P1_U3046) );
  AOI22_X1 U24194 ( .A1(n21197), .A2(n21510), .B1(n21509), .B2(n21196), .ZN(
        n21195) );
  AOI22_X1 U24195 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n21198), .B1(
        n21226), .B2(n21511), .ZN(n21194) );
  OAI211_X1 U24196 ( .C1(n21514), .C2(n21201), .A(n21195), .B(n21194), .ZN(
        P1_U3047) );
  AOI22_X1 U24197 ( .A1(n21197), .A2(n21517), .B1(n21516), .B2(n21196), .ZN(
        n21200) );
  AOI22_X1 U24198 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n21198), .B1(
        n21226), .B2(n21519), .ZN(n21199) );
  OAI211_X1 U24199 ( .C1(n21525), .C2(n21201), .A(n21200), .B(n21199), .ZN(
        P1_U3048) );
  NOR3_X1 U24200 ( .A1(n21226), .A2(n21262), .A3(n21417), .ZN(n21203) );
  INV_X1 U24201 ( .A(n21377), .ZN(n21296) );
  NOR2_X1 U24202 ( .A1(n21203), .A2(n21296), .ZN(n21210) );
  INV_X1 U24203 ( .A(n21210), .ZN(n21204) );
  NOR2_X1 U24204 ( .A1(n21237), .A2(n13944), .ZN(n21209) );
  NAND2_X1 U24205 ( .A1(n21380), .A2(n15793), .ZN(n21207) );
  INV_X1 U24206 ( .A(n21207), .ZN(n21299) );
  NOR3_X2 U24207 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21681), .A3(
        n21240), .ZN(n21225) );
  AOI22_X1 U24208 ( .A1(n21226), .A2(n21425), .B1(n21465), .B2(n21225), .ZN(
        n21212) );
  INV_X1 U24209 ( .A(n21225), .ZN(n21206) );
  INV_X1 U24210 ( .A(n21386), .ZN(n21205) );
  AOI21_X1 U24211 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n21206), .A(n21205), 
        .ZN(n21208) );
  NAND2_X1 U24212 ( .A1(n21207), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n21305) );
  AOI22_X1 U24213 ( .A1(n21227), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n21262), .B2(n21477), .ZN(n21211) );
  OAI211_X1 U24214 ( .C1(n21230), .C2(n21394), .A(n21212), .B(n21211), .ZN(
        P1_U3049) );
  AOI22_X1 U24215 ( .A1(n21226), .A2(n21429), .B1(n21481), .B2(n21225), .ZN(
        n21214) );
  AOI22_X1 U24216 ( .A1(n21227), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n21262), .B2(n21483), .ZN(n21213) );
  OAI211_X1 U24217 ( .C1(n21230), .C2(n21397), .A(n21214), .B(n21213), .ZN(
        P1_U3050) );
  AOI22_X1 U24218 ( .A1(n21226), .A2(n21929), .B1(n21928), .B2(n21225), .ZN(
        n21216) );
  AOI22_X1 U24219 ( .A1(n21227), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n21262), .B2(n21931), .ZN(n21215) );
  OAI211_X1 U24220 ( .C1(n21230), .C2(n21936), .A(n21216), .B(n21215), .ZN(
        P1_U3051) );
  AOI22_X1 U24221 ( .A1(n21226), .A2(n21436), .B1(n21491), .B2(n21225), .ZN(
        n21218) );
  AOI22_X1 U24222 ( .A1(n21227), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n21262), .B2(n21493), .ZN(n21217) );
  OAI211_X1 U24223 ( .C1(n21230), .C2(n21400), .A(n21218), .B(n21217), .ZN(
        P1_U3052) );
  AOI22_X1 U24224 ( .A1(n21226), .A2(n21440), .B1(n21497), .B2(n21225), .ZN(
        n21220) );
  AOI22_X1 U24225 ( .A1(n21227), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n21262), .B2(n21499), .ZN(n21219) );
  OAI211_X1 U24226 ( .C1(n21230), .C2(n21403), .A(n21220), .B(n21219), .ZN(
        P1_U3053) );
  AOI22_X1 U24227 ( .A1(n21226), .A2(n21444), .B1(n21503), .B2(n21225), .ZN(
        n21222) );
  AOI22_X1 U24228 ( .A1(n21227), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n21262), .B2(n21505), .ZN(n21221) );
  OAI211_X1 U24229 ( .C1(n21230), .C2(n21406), .A(n21222), .B(n21221), .ZN(
        P1_U3054) );
  AOI22_X1 U24230 ( .A1(n21226), .A2(n21448), .B1(n21509), .B2(n21225), .ZN(
        n21224) );
  AOI22_X1 U24231 ( .A1(n21227), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n21262), .B2(n21511), .ZN(n21223) );
  OAI211_X1 U24232 ( .C1(n21230), .C2(n21409), .A(n21224), .B(n21223), .ZN(
        P1_U3055) );
  AOI22_X1 U24233 ( .A1(n21226), .A2(n21454), .B1(n21516), .B2(n21225), .ZN(
        n21229) );
  AOI22_X1 U24234 ( .A1(n21227), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n21262), .B2(n21519), .ZN(n21228) );
  OAI211_X1 U24235 ( .C1(n21230), .C2(n21412), .A(n21229), .B(n21228), .ZN(
        P1_U3056) );
  NOR2_X1 U24236 ( .A1(n21681), .A2(n21240), .ZN(n21238) );
  INV_X1 U24237 ( .A(n21231), .ZN(n21232) );
  AOI21_X1 U24238 ( .B1(n21233), .B2(n21232), .A(n21417), .ZN(n21239) );
  INV_X1 U24239 ( .A(n21240), .ZN(n21234) );
  NAND2_X1 U24240 ( .A1(n21235), .A2(n21234), .ZN(n21246) );
  OAI21_X1 U24241 ( .B1(n21237), .B2(n21236), .A(n21246), .ZN(n21242) );
  INV_X1 U24242 ( .A(n21246), .ZN(n21260) );
  AOI22_X1 U24243 ( .A1(n21261), .A2(n21477), .B1(n21260), .B2(n21465), .ZN(
        n21245) );
  INV_X1 U24244 ( .A(n21239), .ZN(n21243) );
  OAI21_X1 U24245 ( .B1(n21681), .B2(n21240), .A(n21417), .ZN(n21241) );
  OAI211_X1 U24246 ( .C1(n21243), .C2(n21242), .A(n21422), .B(n21241), .ZN(
        n21263) );
  AOI22_X1 U24247 ( .A1(n21263), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n21262), .B2(n21425), .ZN(n21244) );
  OAI211_X1 U24248 ( .C1(n21266), .C2(n21394), .A(n21245), .B(n21244), .ZN(
        P1_U3057) );
  NOR2_X1 U24249 ( .A1(n21313), .A2(n21246), .ZN(n21247) );
  AOI21_X1 U24250 ( .B1(n21262), .B2(n21429), .A(n21247), .ZN(n21249) );
  AOI22_X1 U24251 ( .A1(n21263), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n21261), .B2(n21483), .ZN(n21248) );
  OAI211_X1 U24252 ( .C1(n21266), .C2(n21397), .A(n21249), .B(n21248), .ZN(
        P1_U3058) );
  AOI22_X1 U24253 ( .A1(n21261), .A2(n21931), .B1(n21260), .B2(n21928), .ZN(
        n21251) );
  AOI22_X1 U24254 ( .A1(n21263), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n21262), .B2(n21929), .ZN(n21250) );
  OAI211_X1 U24255 ( .C1(n21266), .C2(n21936), .A(n21251), .B(n21250), .ZN(
        P1_U3059) );
  AOI22_X1 U24256 ( .A1(n21261), .A2(n21493), .B1(n21260), .B2(n21491), .ZN(
        n21253) );
  AOI22_X1 U24257 ( .A1(n21263), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n21262), .B2(n21436), .ZN(n21252) );
  OAI211_X1 U24258 ( .C1(n21266), .C2(n21400), .A(n21253), .B(n21252), .ZN(
        P1_U3060) );
  AOI22_X1 U24259 ( .A1(n21262), .A2(n21440), .B1(n21497), .B2(n21260), .ZN(
        n21255) );
  AOI22_X1 U24260 ( .A1(n21263), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n21261), .B2(n21499), .ZN(n21254) );
  OAI211_X1 U24261 ( .C1(n21266), .C2(n21403), .A(n21255), .B(n21254), .ZN(
        P1_U3061) );
  AOI22_X1 U24262 ( .A1(n21261), .A2(n21505), .B1(n21260), .B2(n21503), .ZN(
        n21257) );
  AOI22_X1 U24263 ( .A1(n21263), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n21262), .B2(n21444), .ZN(n21256) );
  OAI211_X1 U24264 ( .C1(n21266), .C2(n21406), .A(n21257), .B(n21256), .ZN(
        P1_U3062) );
  AOI22_X1 U24265 ( .A1(n21262), .A2(n21448), .B1(n21509), .B2(n21260), .ZN(
        n21259) );
  AOI22_X1 U24266 ( .A1(n21263), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n21261), .B2(n21511), .ZN(n21258) );
  OAI211_X1 U24267 ( .C1(n21266), .C2(n21409), .A(n21259), .B(n21258), .ZN(
        P1_U3063) );
  AOI22_X1 U24268 ( .A1(n21261), .A2(n21519), .B1(n21260), .B2(n21516), .ZN(
        n21265) );
  AOI22_X1 U24269 ( .A1(n21263), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n21262), .B2(n21454), .ZN(n21264) );
  OAI211_X1 U24270 ( .C1(n21266), .C2(n21412), .A(n21265), .B(n21264), .ZN(
        P1_U3064) );
  NOR2_X1 U24271 ( .A1(n21269), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n21275) );
  INV_X1 U24272 ( .A(n21275), .ZN(n21271) );
  NOR2_X1 U24273 ( .A1(n21414), .A2(n21271), .ZN(n21290) );
  AOI21_X1 U24274 ( .B1(n21270), .B2(n21347), .A(n21290), .ZN(n21272) );
  OAI22_X1 U24275 ( .A1(n21272), .A2(n21417), .B1(n21271), .B2(n21349), .ZN(
        n21291) );
  AOI22_X1 U24276 ( .A1(n21291), .A2(n21466), .B1(n21465), .B2(n21290), .ZN(
        n21277) );
  OAI21_X1 U24277 ( .B1(n21273), .B2(n21468), .A(n21272), .ZN(n21274) );
  OAI221_X1 U24278 ( .B1(n21376), .B2(n21275), .C1(n21417), .C2(n21274), .A(
        n21422), .ZN(n21293) );
  AOI22_X1 U24279 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n21293), .B1(
        n21292), .B2(n21425), .ZN(n21276) );
  OAI211_X1 U24280 ( .C1(n21428), .C2(n21339), .A(n21277), .B(n21276), .ZN(
        P1_U3073) );
  AOI22_X1 U24281 ( .A1(n21291), .A2(n21482), .B1(n21481), .B2(n21290), .ZN(
        n21279) );
  AOI22_X1 U24282 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n21293), .B1(
        n21292), .B2(n21429), .ZN(n21278) );
  OAI211_X1 U24283 ( .C1(n21432), .C2(n21339), .A(n21279), .B(n21278), .ZN(
        P1_U3074) );
  AOI22_X1 U24284 ( .A1(n21291), .A2(n21487), .B1(n21928), .B2(n21290), .ZN(
        n21281) );
  AOI22_X1 U24285 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n21293), .B1(
        n21292), .B2(n21929), .ZN(n21280) );
  OAI211_X1 U24286 ( .C1(n21435), .C2(n21339), .A(n21281), .B(n21280), .ZN(
        P1_U3075) );
  AOI22_X1 U24287 ( .A1(n21291), .A2(n21492), .B1(n21491), .B2(n21290), .ZN(
        n21283) );
  AOI22_X1 U24288 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n21293), .B1(
        n21292), .B2(n21436), .ZN(n21282) );
  OAI211_X1 U24289 ( .C1(n21439), .C2(n21339), .A(n21283), .B(n21282), .ZN(
        P1_U3076) );
  AOI22_X1 U24290 ( .A1(n21291), .A2(n21498), .B1(n21497), .B2(n21290), .ZN(
        n21285) );
  AOI22_X1 U24291 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n21293), .B1(
        n21292), .B2(n21440), .ZN(n21284) );
  OAI211_X1 U24292 ( .C1(n21443), .C2(n21339), .A(n21285), .B(n21284), .ZN(
        P1_U3077) );
  AOI22_X1 U24293 ( .A1(n21291), .A2(n21504), .B1(n21503), .B2(n21290), .ZN(
        n21287) );
  AOI22_X1 U24294 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n21293), .B1(
        n21292), .B2(n21444), .ZN(n21286) );
  OAI211_X1 U24295 ( .C1(n21447), .C2(n21339), .A(n21287), .B(n21286), .ZN(
        P1_U3078) );
  AOI22_X1 U24296 ( .A1(n21291), .A2(n21510), .B1(n21509), .B2(n21290), .ZN(
        n21289) );
  AOI22_X1 U24297 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n21293), .B1(
        n21292), .B2(n21448), .ZN(n21288) );
  OAI211_X1 U24298 ( .C1(n21451), .C2(n21339), .A(n21289), .B(n21288), .ZN(
        P1_U3079) );
  AOI22_X1 U24299 ( .A1(n21291), .A2(n21517), .B1(n21516), .B2(n21290), .ZN(
        n21295) );
  AOI22_X1 U24300 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n21293), .B1(
        n21292), .B2(n21454), .ZN(n21294) );
  OAI211_X1 U24301 ( .C1(n21459), .C2(n21339), .A(n21295), .B(n21294), .ZN(
        P1_U3080) );
  NOR2_X1 U24302 ( .A1(n21341), .A2(n21417), .ZN(n21297) );
  AOI21_X1 U24303 ( .B1(n21297), .B2(n21339), .A(n21296), .ZN(n21310) );
  INV_X1 U24304 ( .A(n21310), .ZN(n21300) );
  NOR2_X1 U24305 ( .A1(n21298), .A2(n13944), .ZN(n21309) );
  INV_X1 U24306 ( .A(n21301), .ZN(n21302) );
  NOR2_X1 U24307 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21302), .ZN(
        n21306) );
  INV_X1 U24308 ( .A(n21306), .ZN(n21338) );
  OAI22_X1 U24309 ( .A1(n21339), .A2(n21480), .B1(n21303), .B2(n21338), .ZN(
        n21304) );
  INV_X1 U24310 ( .A(n21304), .ZN(n21312) );
  OAI211_X1 U24311 ( .C1(n21306), .C2(n21719), .A(n21473), .B(n21305), .ZN(
        n21307) );
  INV_X1 U24312 ( .A(n21307), .ZN(n21308) );
  AOI22_X1 U24313 ( .A1(n21342), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n21341), .B2(n21477), .ZN(n21311) );
  OAI211_X1 U24314 ( .C1(n21345), .C2(n21394), .A(n21312), .B(n21311), .ZN(
        P1_U3081) );
  OAI22_X1 U24315 ( .A1(n21339), .A2(n21486), .B1(n21338), .B2(n21313), .ZN(
        n21314) );
  INV_X1 U24316 ( .A(n21314), .ZN(n21316) );
  AOI22_X1 U24317 ( .A1(n21342), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n21341), .B2(n21483), .ZN(n21315) );
  OAI211_X1 U24318 ( .C1(n21345), .C2(n21397), .A(n21316), .B(n21315), .ZN(
        P1_U3082) );
  OAI22_X1 U24319 ( .A1(n21339), .A2(n21490), .B1(n21338), .B2(n21317), .ZN(
        n21318) );
  INV_X1 U24320 ( .A(n21318), .ZN(n21320) );
  AOI22_X1 U24321 ( .A1(n21342), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n21341), .B2(n21931), .ZN(n21319) );
  OAI211_X1 U24322 ( .C1(n21345), .C2(n21936), .A(n21320), .B(n21319), .ZN(
        P1_U3083) );
  OAI22_X1 U24323 ( .A1(n21339), .A2(n21496), .B1(n21338), .B2(n21321), .ZN(
        n21322) );
  INV_X1 U24324 ( .A(n21322), .ZN(n21324) );
  AOI22_X1 U24325 ( .A1(n21342), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n21341), .B2(n21493), .ZN(n21323) );
  OAI211_X1 U24326 ( .C1(n21345), .C2(n21400), .A(n21324), .B(n21323), .ZN(
        P1_U3084) );
  OAI22_X1 U24327 ( .A1(n21339), .A2(n21502), .B1(n21338), .B2(n21325), .ZN(
        n21326) );
  INV_X1 U24328 ( .A(n21326), .ZN(n21328) );
  AOI22_X1 U24329 ( .A1(n21342), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n21341), .B2(n21499), .ZN(n21327) );
  OAI211_X1 U24330 ( .C1(n21345), .C2(n21403), .A(n21328), .B(n21327), .ZN(
        P1_U3085) );
  OAI22_X1 U24331 ( .A1(n21339), .A2(n21508), .B1(n21338), .B2(n21329), .ZN(
        n21330) );
  INV_X1 U24332 ( .A(n21330), .ZN(n21332) );
  AOI22_X1 U24333 ( .A1(n21342), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n21341), .B2(n21505), .ZN(n21331) );
  OAI211_X1 U24334 ( .C1(n21345), .C2(n21406), .A(n21332), .B(n21331), .ZN(
        P1_U3086) );
  OAI22_X1 U24335 ( .A1(n21339), .A2(n21514), .B1(n21333), .B2(n21338), .ZN(
        n21334) );
  INV_X1 U24336 ( .A(n21334), .ZN(n21336) );
  AOI22_X1 U24337 ( .A1(n21342), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n21341), .B2(n21511), .ZN(n21335) );
  OAI211_X1 U24338 ( .C1(n21345), .C2(n21409), .A(n21336), .B(n21335), .ZN(
        P1_U3087) );
  OAI22_X1 U24339 ( .A1(n21339), .A2(n21525), .B1(n21338), .B2(n21337), .ZN(
        n21340) );
  INV_X1 U24340 ( .A(n21340), .ZN(n21344) );
  AOI22_X1 U24341 ( .A1(n21342), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n21341), .B2(n21519), .ZN(n21343) );
  OAI211_X1 U24342 ( .C1(n21345), .C2(n21412), .A(n21344), .B(n21343), .ZN(
        P1_U3088) );
  NOR2_X1 U24343 ( .A1(n21346), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n21353) );
  INV_X1 U24344 ( .A(n21353), .ZN(n21350) );
  NOR2_X1 U24345 ( .A1(n21414), .A2(n21350), .ZN(n21370) );
  AOI21_X1 U24346 ( .B1(n21348), .B2(n21347), .A(n21370), .ZN(n21351) );
  OAI22_X1 U24347 ( .A1(n21351), .A2(n21417), .B1(n21350), .B2(n21349), .ZN(
        n21371) );
  AOI22_X1 U24348 ( .A1(n21371), .A2(n21466), .B1(n21465), .B2(n21370), .ZN(
        n21357) );
  OAI21_X1 U24349 ( .B1(n21355), .B2(n21468), .A(n21351), .ZN(n21352) );
  OAI221_X1 U24350 ( .B1(n21376), .B2(n21353), .C1(n21417), .C2(n21352), .A(
        n21422), .ZN(n21372) );
  AOI22_X1 U24351 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n21372), .B1(
        n21930), .B2(n21477), .ZN(n21356) );
  OAI211_X1 U24352 ( .C1(n21480), .C2(n21375), .A(n21357), .B(n21356), .ZN(
        P1_U3105) );
  AOI22_X1 U24353 ( .A1(n21371), .A2(n21482), .B1(n21481), .B2(n21370), .ZN(
        n21359) );
  AOI22_X1 U24354 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n21372), .B1(
        n21930), .B2(n21483), .ZN(n21358) );
  OAI211_X1 U24355 ( .C1(n21486), .C2(n21375), .A(n21359), .B(n21358), .ZN(
        P1_U3106) );
  AOI22_X1 U24356 ( .A1(n21371), .A2(n21487), .B1(n21928), .B2(n21370), .ZN(
        n21361) );
  AOI22_X1 U24357 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n21372), .B1(
        n21930), .B2(n21931), .ZN(n21360) );
  OAI211_X1 U24358 ( .C1(n21490), .C2(n21375), .A(n21361), .B(n21360), .ZN(
        P1_U3107) );
  AOI22_X1 U24359 ( .A1(n21371), .A2(n21492), .B1(n21491), .B2(n21370), .ZN(
        n21363) );
  AOI22_X1 U24360 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n21372), .B1(
        n21930), .B2(n21493), .ZN(n21362) );
  OAI211_X1 U24361 ( .C1(n21496), .C2(n21375), .A(n21363), .B(n21362), .ZN(
        P1_U3108) );
  AOI22_X1 U24362 ( .A1(n21371), .A2(n21498), .B1(n21497), .B2(n21370), .ZN(
        n21365) );
  AOI22_X1 U24363 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n21372), .B1(
        n21930), .B2(n21499), .ZN(n21364) );
  OAI211_X1 U24364 ( .C1(n21502), .C2(n21375), .A(n21365), .B(n21364), .ZN(
        P1_U3109) );
  AOI22_X1 U24365 ( .A1(n21371), .A2(n21504), .B1(n21503), .B2(n21370), .ZN(
        n21367) );
  AOI22_X1 U24366 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n21372), .B1(
        n21930), .B2(n21505), .ZN(n21366) );
  OAI211_X1 U24367 ( .C1(n21508), .C2(n21375), .A(n21367), .B(n21366), .ZN(
        P1_U3110) );
  AOI22_X1 U24368 ( .A1(n21371), .A2(n21510), .B1(n21509), .B2(n21370), .ZN(
        n21369) );
  AOI22_X1 U24369 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n21372), .B1(
        n21930), .B2(n21511), .ZN(n21368) );
  OAI211_X1 U24370 ( .C1(n21514), .C2(n21375), .A(n21369), .B(n21368), .ZN(
        P1_U3111) );
  AOI22_X1 U24371 ( .A1(n21371), .A2(n21517), .B1(n21516), .B2(n21370), .ZN(
        n21374) );
  AOI22_X1 U24372 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n21372), .B1(
        n21930), .B2(n21519), .ZN(n21373) );
  OAI211_X1 U24373 ( .C1(n21525), .C2(n21375), .A(n21374), .B(n21373), .ZN(
        P1_U3112) );
  NAND2_X1 U24374 ( .A1(n21391), .A2(n21376), .ZN(n21378) );
  OAI21_X1 U24375 ( .B1(n21930), .B2(n21378), .A(n21377), .ZN(n21389) );
  OR2_X1 U24376 ( .A1(n21379), .A2(n13944), .ZN(n21388) );
  INV_X1 U24377 ( .A(n21388), .ZN(n21383) );
  NAND2_X1 U24378 ( .A1(n21380), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n21461) );
  INV_X1 U24379 ( .A(n21461), .ZN(n21381) );
  INV_X1 U24380 ( .A(n21384), .ZN(n21385) );
  NOR2_X1 U24381 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21385), .ZN(
        n21927) );
  AOI22_X1 U24382 ( .A1(n21930), .A2(n21425), .B1(n21465), .B2(n21927), .ZN(
        n21393) );
  NAND2_X1 U24383 ( .A1(n21461), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n21474) );
  OAI211_X1 U24384 ( .C1(n21719), .C2(n21927), .A(n21386), .B(n21474), .ZN(
        n21387) );
  AOI21_X1 U24385 ( .B1(n21389), .B2(n21388), .A(n21387), .ZN(n21390) );
  AOI22_X1 U24386 ( .A1(n21933), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n21932), .B2(n21477), .ZN(n21392) );
  OAI211_X1 U24387 ( .C1(n21937), .C2(n21394), .A(n21393), .B(n21392), .ZN(
        P1_U3113) );
  AOI22_X1 U24388 ( .A1(n21930), .A2(n21429), .B1(n21481), .B2(n21927), .ZN(
        n21396) );
  AOI22_X1 U24389 ( .A1(n21933), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n21932), .B2(n21483), .ZN(n21395) );
  OAI211_X1 U24390 ( .C1(n21937), .C2(n21397), .A(n21396), .B(n21395), .ZN(
        P1_U3114) );
  AOI22_X1 U24391 ( .A1(n21930), .A2(n21436), .B1(n21491), .B2(n21927), .ZN(
        n21399) );
  AOI22_X1 U24392 ( .A1(n21933), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n21932), .B2(n21493), .ZN(n21398) );
  OAI211_X1 U24393 ( .C1(n21937), .C2(n21400), .A(n21399), .B(n21398), .ZN(
        P1_U3116) );
  AOI22_X1 U24394 ( .A1(n21930), .A2(n21440), .B1(n21497), .B2(n21927), .ZN(
        n21402) );
  AOI22_X1 U24395 ( .A1(n21933), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n21932), .B2(n21499), .ZN(n21401) );
  OAI211_X1 U24396 ( .C1(n21937), .C2(n21403), .A(n21402), .B(n21401), .ZN(
        P1_U3117) );
  AOI22_X1 U24397 ( .A1(n21930), .A2(n21444), .B1(n21503), .B2(n21927), .ZN(
        n21405) );
  AOI22_X1 U24398 ( .A1(n21933), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n21932), .B2(n21505), .ZN(n21404) );
  OAI211_X1 U24399 ( .C1(n21937), .C2(n21406), .A(n21405), .B(n21404), .ZN(
        P1_U3118) );
  AOI22_X1 U24400 ( .A1(n21930), .A2(n21448), .B1(n21509), .B2(n21927), .ZN(
        n21408) );
  AOI22_X1 U24401 ( .A1(n21933), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n21932), .B2(n21511), .ZN(n21407) );
  OAI211_X1 U24402 ( .C1(n21937), .C2(n21409), .A(n21408), .B(n21407), .ZN(
        P1_U3119) );
  AOI22_X1 U24403 ( .A1(n21930), .A2(n21454), .B1(n21516), .B2(n21927), .ZN(
        n21411) );
  AOI22_X1 U24404 ( .A1(n21933), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n21932), .B2(n21519), .ZN(n21410) );
  OAI211_X1 U24405 ( .C1(n21937), .C2(n21412), .A(n21411), .B(n21410), .ZN(
        P1_U3120) );
  NOR2_X1 U24406 ( .A1(n21464), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n21423) );
  INV_X1 U24407 ( .A(n21423), .ZN(n21416) );
  NOR2_X1 U24408 ( .A1(n21414), .A2(n21416), .ZN(n21452) );
  INV_X1 U24409 ( .A(n21452), .ZN(n21418) );
  INV_X1 U24410 ( .A(n21415), .ZN(n21463) );
  OAI222_X1 U24411 ( .A1(n21418), .A2(n21417), .B1(n21349), .B2(n21416), .C1(
        n21174), .C2(n21463), .ZN(n21453) );
  AOI22_X1 U24412 ( .A1(n21453), .A2(n21466), .B1(n21465), .B2(n21452), .ZN(
        n21427) );
  INV_X1 U24413 ( .A(n21419), .ZN(n21421) );
  NOR2_X1 U24414 ( .A1(n21421), .A2(n21420), .ZN(n21424) );
  AOI22_X1 U24415 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n21456), .B1(
        n21455), .B2(n21425), .ZN(n21426) );
  OAI211_X1 U24416 ( .C1(n21428), .C2(n21524), .A(n21427), .B(n21426), .ZN(
        P1_U3137) );
  AOI22_X1 U24417 ( .A1(n21453), .A2(n21482), .B1(n21481), .B2(n21452), .ZN(
        n21431) );
  AOI22_X1 U24418 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n21456), .B1(
        n21455), .B2(n21429), .ZN(n21430) );
  OAI211_X1 U24419 ( .C1(n21432), .C2(n21524), .A(n21431), .B(n21430), .ZN(
        P1_U3138) );
  AOI22_X1 U24420 ( .A1(n21453), .A2(n21487), .B1(n21928), .B2(n21452), .ZN(
        n21434) );
  AOI22_X1 U24421 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n21456), .B1(
        n21455), .B2(n21929), .ZN(n21433) );
  OAI211_X1 U24422 ( .C1(n21435), .C2(n21524), .A(n21434), .B(n21433), .ZN(
        P1_U3139) );
  AOI22_X1 U24423 ( .A1(n21453), .A2(n21492), .B1(n21491), .B2(n21452), .ZN(
        n21438) );
  AOI22_X1 U24424 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n21456), .B1(
        n21455), .B2(n21436), .ZN(n21437) );
  OAI211_X1 U24425 ( .C1(n21439), .C2(n21524), .A(n21438), .B(n21437), .ZN(
        P1_U3140) );
  AOI22_X1 U24426 ( .A1(n21453), .A2(n21498), .B1(n21497), .B2(n21452), .ZN(
        n21442) );
  AOI22_X1 U24427 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n21456), .B1(
        n21455), .B2(n21440), .ZN(n21441) );
  OAI211_X1 U24428 ( .C1(n21443), .C2(n21524), .A(n21442), .B(n21441), .ZN(
        P1_U3141) );
  AOI22_X1 U24429 ( .A1(n21453), .A2(n21504), .B1(n21503), .B2(n21452), .ZN(
        n21446) );
  AOI22_X1 U24430 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n21456), .B1(
        n21455), .B2(n21444), .ZN(n21445) );
  OAI211_X1 U24431 ( .C1(n21447), .C2(n21524), .A(n21446), .B(n21445), .ZN(
        P1_U3142) );
  AOI22_X1 U24432 ( .A1(n21453), .A2(n21510), .B1(n21509), .B2(n21452), .ZN(
        n21450) );
  AOI22_X1 U24433 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n21456), .B1(
        n21455), .B2(n21448), .ZN(n21449) );
  OAI211_X1 U24434 ( .C1(n21451), .C2(n21524), .A(n21450), .B(n21449), .ZN(
        P1_U3143) );
  AOI22_X1 U24435 ( .A1(n21453), .A2(n21517), .B1(n21516), .B2(n21452), .ZN(
        n21458) );
  AOI22_X1 U24436 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n21456), .B1(
        n21455), .B2(n21454), .ZN(n21457) );
  OAI211_X1 U24437 ( .C1(n21459), .C2(n21524), .A(n21458), .B(n21457), .ZN(
        P1_U3144) );
  INV_X1 U24438 ( .A(n21460), .ZN(n21462) );
  OAI22_X1 U24439 ( .A1(n21463), .A2(n13944), .B1(n21462), .B2(n21461), .ZN(
        n21518) );
  NOR3_X2 U24440 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21681), .A3(
        n21464), .ZN(n21515) );
  AOI22_X1 U24441 ( .A1(n21518), .A2(n21466), .B1(n21465), .B2(n21515), .ZN(
        n21479) );
  INV_X1 U24442 ( .A(n21467), .ZN(n21470) );
  AOI21_X1 U24443 ( .B1(n21524), .B2(n21476), .A(n21468), .ZN(n21469) );
  AOI21_X1 U24444 ( .B1(n21471), .B2(n21470), .A(n21469), .ZN(n21472) );
  NOR2_X1 U24445 ( .A1(n21472), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n21475) );
  AOI22_X1 U24446 ( .A1(n21521), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n21520), .B2(n21477), .ZN(n21478) );
  OAI211_X1 U24447 ( .C1(n21480), .C2(n21524), .A(n21479), .B(n21478), .ZN(
        P1_U3145) );
  AOI22_X1 U24448 ( .A1(n21518), .A2(n21482), .B1(n21481), .B2(n21515), .ZN(
        n21485) );
  AOI22_X1 U24449 ( .A1(n21521), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n21520), .B2(n21483), .ZN(n21484) );
  OAI211_X1 U24450 ( .C1(n21486), .C2(n21524), .A(n21485), .B(n21484), .ZN(
        P1_U3146) );
  AOI22_X1 U24451 ( .A1(n21518), .A2(n21487), .B1(n21928), .B2(n21515), .ZN(
        n21489) );
  AOI22_X1 U24452 ( .A1(n21521), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n21520), .B2(n21931), .ZN(n21488) );
  OAI211_X1 U24453 ( .C1(n21490), .C2(n21524), .A(n21489), .B(n21488), .ZN(
        P1_U3147) );
  AOI22_X1 U24454 ( .A1(n21518), .A2(n21492), .B1(n21491), .B2(n21515), .ZN(
        n21495) );
  AOI22_X1 U24455 ( .A1(n21521), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n21520), .B2(n21493), .ZN(n21494) );
  OAI211_X1 U24456 ( .C1(n21496), .C2(n21524), .A(n21495), .B(n21494), .ZN(
        P1_U3148) );
  AOI22_X1 U24457 ( .A1(n21518), .A2(n21498), .B1(n21497), .B2(n21515), .ZN(
        n21501) );
  AOI22_X1 U24458 ( .A1(n21521), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n21520), .B2(n21499), .ZN(n21500) );
  OAI211_X1 U24459 ( .C1(n21502), .C2(n21524), .A(n21501), .B(n21500), .ZN(
        P1_U3149) );
  AOI22_X1 U24460 ( .A1(n21518), .A2(n21504), .B1(n21503), .B2(n21515), .ZN(
        n21507) );
  AOI22_X1 U24461 ( .A1(n21521), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n21520), .B2(n21505), .ZN(n21506) );
  OAI211_X1 U24462 ( .C1(n21508), .C2(n21524), .A(n21507), .B(n21506), .ZN(
        P1_U3150) );
  AOI22_X1 U24463 ( .A1(n21518), .A2(n21510), .B1(n21509), .B2(n21515), .ZN(
        n21513) );
  AOI22_X1 U24464 ( .A1(n21521), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n21520), .B2(n21511), .ZN(n21512) );
  OAI211_X1 U24465 ( .C1(n21514), .C2(n21524), .A(n21513), .B(n21512), .ZN(
        P1_U3151) );
  AOI22_X1 U24466 ( .A1(n21518), .A2(n21517), .B1(n21516), .B2(n21515), .ZN(
        n21523) );
  AOI22_X1 U24467 ( .A1(n21521), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n21520), .B2(n21519), .ZN(n21522) );
  OAI211_X1 U24468 ( .C1(n21525), .C2(n21524), .A(n21523), .B(n21522), .ZN(
        P1_U3152) );
  AND2_X1 U24469 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n21526), .ZN(
        P1_U3164) );
  INV_X1 U24470 ( .A(P1_DATAWIDTH_REG_30__SCAN_IN), .ZN(n21838) );
  NOR2_X1 U24471 ( .A1(n21591), .A2(n21838), .ZN(P1_U3165) );
  AND2_X1 U24472 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n21526), .ZN(
        P1_U3166) );
  AND2_X1 U24473 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n21526), .ZN(
        P1_U3167) );
  AND2_X1 U24474 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n21526), .ZN(
        P1_U3168) );
  AND2_X1 U24475 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n21526), .ZN(
        P1_U3169) );
  AND2_X1 U24476 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n21526), .ZN(
        P1_U3170) );
  AND2_X1 U24477 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n21526), .ZN(
        P1_U3171) );
  AND2_X1 U24478 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n21526), .ZN(
        P1_U3172) );
  AND2_X1 U24479 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n21526), .ZN(
        P1_U3173) );
  AND2_X1 U24480 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n21526), .ZN(
        P1_U3174) );
  AND2_X1 U24481 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n21526), .ZN(
        P1_U3175) );
  AND2_X1 U24482 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n21526), .ZN(
        P1_U3176) );
  AND2_X1 U24483 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n21526), .ZN(
        P1_U3177) );
  AND2_X1 U24484 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n21526), .ZN(
        P1_U3178) );
  AND2_X1 U24485 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n21526), .ZN(
        P1_U3179) );
  AND2_X1 U24486 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n21526), .ZN(
        P1_U3180) );
  AND2_X1 U24487 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n21526), .ZN(
        P1_U3181) );
  AND2_X1 U24488 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n21526), .ZN(
        P1_U3182) );
  INV_X1 U24489 ( .A(P1_DATAWIDTH_REG_12__SCAN_IN), .ZN(n21834) );
  NOR2_X1 U24490 ( .A1(n21591), .A2(n21834), .ZN(P1_U3183) );
  AND2_X1 U24491 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n21526), .ZN(
        P1_U3184) );
  AND2_X1 U24492 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n21526), .ZN(
        P1_U3185) );
  AND2_X1 U24493 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n21526), .ZN(P1_U3186) );
  AND2_X1 U24494 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n21526), .ZN(P1_U3187) );
  AND2_X1 U24495 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n21526), .ZN(P1_U3188) );
  AND2_X1 U24496 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n21526), .ZN(P1_U3189) );
  AND2_X1 U24497 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n21526), .ZN(P1_U3190) );
  AND2_X1 U24498 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n21526), .ZN(P1_U3191) );
  AND2_X1 U24499 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n21526), .ZN(P1_U3192) );
  AND2_X1 U24500 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n21526), .ZN(P1_U3193) );
  AOI21_X1 U24501 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n21533), .A(n21527), 
        .ZN(n21534) );
  OAI21_X1 U24502 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(P1_STATE_REG_2__SCAN_IN), 
        .A(HOLD), .ZN(n21528) );
  OAI211_X1 U24503 ( .C1(P1_STATE_REG_0__SCAN_IN), .C2(n21536), .A(n21528), 
        .B(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n21529) );
  INV_X1 U24504 ( .A(n21529), .ZN(n21530) );
  OAI22_X1 U24505 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n21534), .B1(n21625), 
        .B2(n21530), .ZN(P1_U3194) );
  AOI21_X1 U24506 ( .B1(n21533), .B2(n21536), .A(n21531), .ZN(n21540) );
  INV_X1 U24507 ( .A(n21532), .ZN(n21533) );
  NAND4_X1 U24508 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .A3(P1_REQUESTPENDING_REG_SCAN_IN), .A4(n21533), .ZN(n21539) );
  INV_X1 U24509 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n21621) );
  OAI211_X1 U24510 ( .C1(P1_STATE_REG_2__SCAN_IN), .C2(n21621), .A(
        P1_STATE_REG_0__SCAN_IN), .B(HOLD), .ZN(n21538) );
  INV_X1 U24511 ( .A(n21534), .ZN(n21535) );
  OAI211_X1 U24512 ( .C1(P1_STATE_REG_1__SCAN_IN), .C2(n21536), .A(
        P1_STATE_REG_2__SCAN_IN), .B(n21535), .ZN(n21537) );
  OAI221_X1 U24513 ( .B1(n21540), .B2(n21539), .C1(n21540), .C2(n21538), .A(
        n21537), .ZN(P1_U3196) );
  INV_X1 U24514 ( .A(n21581), .ZN(n21566) );
  NOR2_X2 U24515 ( .A1(n21541), .A2(n21623), .ZN(n21577) );
  OAI222_X1 U24516 ( .A1(n21566), .A2(n14277), .B1(n21542), .B2(n21625), .C1(
        n21603), .C2(n21583), .ZN(P1_U3197) );
  AOI222_X1 U24517 ( .A1(n21577), .A2(P1_REIP_REG_2__SCAN_IN), .B1(
        P1_ADDRESS_REG_1__SCAN_IN), .B2(n21576), .C1(P1_REIP_REG_3__SCAN_IN), 
        .C2(n21581), .ZN(n21543) );
  INV_X1 U24518 ( .A(n21543), .ZN(P1_U3198) );
  AOI22_X1 U24519 ( .A1(P1_ADDRESS_REG_2__SCAN_IN), .A2(n21623), .B1(
        P1_REIP_REG_4__SCAN_IN), .B2(n21581), .ZN(n21544) );
  OAI21_X1 U24520 ( .B1(n21545), .B2(n21583), .A(n21544), .ZN(P1_U3199) );
  AOI22_X1 U24521 ( .A1(P1_ADDRESS_REG_3__SCAN_IN), .A2(n21576), .B1(
        P1_REIP_REG_5__SCAN_IN), .B2(n21581), .ZN(n21546) );
  OAI21_X1 U24522 ( .B1(n21087), .B2(n21583), .A(n21546), .ZN(P1_U3200) );
  AOI22_X1 U24523 ( .A1(P1_ADDRESS_REG_4__SCAN_IN), .A2(n21576), .B1(
        P1_REIP_REG_6__SCAN_IN), .B2(n21581), .ZN(n21547) );
  OAI21_X1 U24524 ( .B1(n18022), .B2(n21583), .A(n21547), .ZN(P1_U3201) );
  INV_X1 U24525 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n21550) );
  AOI22_X1 U24526 ( .A1(P1_ADDRESS_REG_5__SCAN_IN), .A2(n21576), .B1(
        P1_REIP_REG_6__SCAN_IN), .B2(n21577), .ZN(n21548) );
  OAI21_X1 U24527 ( .B1(n21550), .B2(n21566), .A(n21548), .ZN(P1_U3202) );
  AOI22_X1 U24528 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(n21576), .B1(
        P1_REIP_REG_8__SCAN_IN), .B2(n21581), .ZN(n21549) );
  OAI21_X1 U24529 ( .B1(n21550), .B2(n21583), .A(n21549), .ZN(P1_U3203) );
  AOI22_X1 U24530 ( .A1(P1_ADDRESS_REG_7__SCAN_IN), .A2(n21576), .B1(
        P1_REIP_REG_8__SCAN_IN), .B2(n21577), .ZN(n21551) );
  OAI21_X1 U24531 ( .B1(n15104), .B2(n21566), .A(n21551), .ZN(P1_U3204) );
  AOI22_X1 U24532 ( .A1(P1_ADDRESS_REG_8__SCAN_IN), .A2(n21576), .B1(
        P1_REIP_REG_10__SCAN_IN), .B2(n21581), .ZN(n21552) );
  OAI21_X1 U24533 ( .B1(n15104), .B2(n21583), .A(n21552), .ZN(P1_U3205) );
  AOI22_X1 U24534 ( .A1(P1_ADDRESS_REG_9__SCAN_IN), .A2(n21623), .B1(
        P1_REIP_REG_10__SCAN_IN), .B2(n21577), .ZN(n21553) );
  OAI21_X1 U24535 ( .B1(n21554), .B2(n21566), .A(n21553), .ZN(P1_U3206) );
  AOI222_X1 U24536 ( .A1(n21577), .A2(P1_REIP_REG_11__SCAN_IN), .B1(
        P1_ADDRESS_REG_10__SCAN_IN), .B2(n21576), .C1(P1_REIP_REG_12__SCAN_IN), 
        .C2(n21581), .ZN(n21555) );
  INV_X1 U24537 ( .A(n21555), .ZN(P1_U3207) );
  AOI222_X1 U24538 ( .A1(n21577), .A2(P1_REIP_REG_12__SCAN_IN), .B1(
        P1_ADDRESS_REG_11__SCAN_IN), .B2(n21576), .C1(P1_REIP_REG_13__SCAN_IN), 
        .C2(n21581), .ZN(n21556) );
  INV_X1 U24539 ( .A(n21556), .ZN(P1_U3208) );
  INV_X1 U24540 ( .A(P1_ADDRESS_REG_12__SCAN_IN), .ZN(n21873) );
  OAI222_X1 U24541 ( .A1(n21583), .A2(n21558), .B1(n21873), .B2(n21625), .C1(
        n21557), .C2(n21566), .ZN(P1_U3209) );
  AOI222_X1 U24542 ( .A1(n21581), .A2(P1_REIP_REG_15__SCAN_IN), .B1(
        P1_ADDRESS_REG_13__SCAN_IN), .B2(n21576), .C1(P1_REIP_REG_14__SCAN_IN), 
        .C2(n21577), .ZN(n21559) );
  INV_X1 U24543 ( .A(n21559), .ZN(P1_U3210) );
  AOI22_X1 U24544 ( .A1(P1_ADDRESS_REG_14__SCAN_IN), .A2(n21576), .B1(
        P1_REIP_REG_16__SCAN_IN), .B2(n21581), .ZN(n21560) );
  OAI21_X1 U24545 ( .B1(n21561), .B2(n21583), .A(n21560), .ZN(P1_U3211) );
  AOI22_X1 U24546 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(n21623), .B1(
        P1_REIP_REG_16__SCAN_IN), .B2(n21577), .ZN(n21562) );
  OAI21_X1 U24547 ( .B1(n21564), .B2(n21566), .A(n21562), .ZN(P1_U3212) );
  AOI22_X1 U24548 ( .A1(P1_ADDRESS_REG_16__SCAN_IN), .A2(n21576), .B1(
        P1_REIP_REG_18__SCAN_IN), .B2(n21581), .ZN(n21563) );
  OAI21_X1 U24549 ( .B1(n21564), .B2(n21583), .A(n21563), .ZN(P1_U3213) );
  AOI22_X1 U24550 ( .A1(P1_ADDRESS_REG_17__SCAN_IN), .A2(n21623), .B1(
        P1_REIP_REG_18__SCAN_IN), .B2(n21577), .ZN(n21565) );
  OAI21_X1 U24551 ( .B1(n21567), .B2(n21566), .A(n21565), .ZN(P1_U3214) );
  INV_X1 U24552 ( .A(P1_ADDRESS_REG_18__SCAN_IN), .ZN(n21821) );
  INV_X1 U24553 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n21850) );
  OAI222_X1 U24554 ( .A1(n21583), .A2(n21567), .B1(n21821), .B2(n21625), .C1(
        n21850), .C2(n21566), .ZN(P1_U3215) );
  AOI222_X1 U24555 ( .A1(n21577), .A2(P1_REIP_REG_20__SCAN_IN), .B1(
        P1_ADDRESS_REG_19__SCAN_IN), .B2(n21576), .C1(P1_REIP_REG_21__SCAN_IN), 
        .C2(n21581), .ZN(n21568) );
  INV_X1 U24556 ( .A(n21568), .ZN(P1_U3216) );
  AOI222_X1 U24557 ( .A1(n21581), .A2(P1_REIP_REG_22__SCAN_IN), .B1(
        P1_ADDRESS_REG_20__SCAN_IN), .B2(n21576), .C1(P1_REIP_REG_21__SCAN_IN), 
        .C2(n21577), .ZN(n21569) );
  INV_X1 U24558 ( .A(n21569), .ZN(P1_U3217) );
  AOI222_X1 U24559 ( .A1(n21577), .A2(P1_REIP_REG_22__SCAN_IN), .B1(
        P1_ADDRESS_REG_21__SCAN_IN), .B2(n21576), .C1(P1_REIP_REG_23__SCAN_IN), 
        .C2(n21581), .ZN(n21570) );
  INV_X1 U24560 ( .A(n21570), .ZN(P1_U3218) );
  AOI222_X1 U24561 ( .A1(n21577), .A2(P1_REIP_REG_23__SCAN_IN), .B1(
        P1_ADDRESS_REG_22__SCAN_IN), .B2(n21576), .C1(P1_REIP_REG_24__SCAN_IN), 
        .C2(n21581), .ZN(n21571) );
  INV_X1 U24562 ( .A(n21571), .ZN(P1_U3219) );
  AOI222_X1 U24563 ( .A1(n21577), .A2(P1_REIP_REG_24__SCAN_IN), .B1(
        P1_ADDRESS_REG_23__SCAN_IN), .B2(n21576), .C1(P1_REIP_REG_25__SCAN_IN), 
        .C2(n21581), .ZN(n21572) );
  INV_X1 U24564 ( .A(n21572), .ZN(P1_U3220) );
  AOI22_X1 U24565 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(n21581), .B1(
        P1_ADDRESS_REG_24__SCAN_IN), .B2(n21623), .ZN(n21573) );
  OAI21_X1 U24566 ( .B1(n21835), .B2(n21583), .A(n21573), .ZN(P1_U3221) );
  AOI222_X1 U24567 ( .A1(n21577), .A2(P1_REIP_REG_26__SCAN_IN), .B1(
        P1_ADDRESS_REG_25__SCAN_IN), .B2(n21576), .C1(P1_REIP_REG_27__SCAN_IN), 
        .C2(n21581), .ZN(n21574) );
  INV_X1 U24568 ( .A(n21574), .ZN(P1_U3222) );
  AOI222_X1 U24569 ( .A1(n21577), .A2(P1_REIP_REG_27__SCAN_IN), .B1(
        P1_ADDRESS_REG_26__SCAN_IN), .B2(n21576), .C1(P1_REIP_REG_28__SCAN_IN), 
        .C2(n21581), .ZN(n21575) );
  INV_X1 U24570 ( .A(n21575), .ZN(P1_U3223) );
  AOI222_X1 U24571 ( .A1(n21577), .A2(P1_REIP_REG_28__SCAN_IN), .B1(
        P1_ADDRESS_REG_27__SCAN_IN), .B2(n21576), .C1(P1_REIP_REG_29__SCAN_IN), 
        .C2(n21581), .ZN(n21578) );
  INV_X1 U24572 ( .A(n21578), .ZN(P1_U3224) );
  AOI22_X1 U24573 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(n21581), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n21623), .ZN(n21579) );
  OAI21_X1 U24574 ( .B1(n21580), .B2(n21583), .A(n21579), .ZN(P1_U3225) );
  AOI22_X1 U24575 ( .A1(P1_REIP_REG_31__SCAN_IN), .A2(n21581), .B1(
        P1_ADDRESS_REG_29__SCAN_IN), .B2(n21623), .ZN(n21582) );
  OAI21_X1 U24576 ( .B1(n12858), .B2(n21583), .A(n21582), .ZN(P1_U3226) );
  OAI22_X1 U24577 ( .A1(n21623), .A2(P1_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P1_BE_N_REG_3__SCAN_IN), .B2(n21625), .ZN(n21584) );
  INV_X1 U24578 ( .A(n21584), .ZN(P1_U3458) );
  OAI22_X1 U24579 ( .A1(n21623), .A2(P1_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P1_BE_N_REG_2__SCAN_IN), .B2(n21625), .ZN(n21585) );
  INV_X1 U24580 ( .A(n21585), .ZN(P1_U3459) );
  OAI22_X1 U24581 ( .A1(n21623), .A2(P1_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P1_BE_N_REG_1__SCAN_IN), .B2(n21625), .ZN(n21586) );
  INV_X1 U24582 ( .A(n21586), .ZN(P1_U3460) );
  OAI22_X1 U24583 ( .A1(n21623), .A2(P1_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P1_BE_N_REG_0__SCAN_IN), .B2(n21625), .ZN(n21587) );
  INV_X1 U24584 ( .A(n21587), .ZN(P1_U3461) );
  OAI21_X1 U24585 ( .B1(P1_DATAWIDTH_REG_0__SCAN_IN), .B2(n21591), .A(n21589), 
        .ZN(n21588) );
  INV_X1 U24586 ( .A(n21588), .ZN(P1_U3464) );
  OAI21_X1 U24587 ( .B1(n21591), .B2(n21590), .A(n21589), .ZN(P1_U3465) );
  INV_X1 U24588 ( .A(n21592), .ZN(n21593) );
  AOI21_X1 U24589 ( .B1(n21593), .B2(n21719), .A(P1_STATE2_REG_1__SCAN_IN), 
        .ZN(n21595) );
  OAI22_X1 U24590 ( .A1(n21596), .A2(n21595), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n21594), .ZN(n21598) );
  AOI22_X1 U24591 ( .A1(n21599), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n21598), .B2(n21597), .ZN(n21600) );
  OAI21_X1 U24592 ( .B1(n21602), .B2(n21601), .A(n21600), .ZN(P1_U3474) );
  AOI21_X1 U24593 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n21604) );
  AOI22_X1 U24594 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .B1(n21604), .B2(n21603), .ZN(n21607) );
  INV_X1 U24595 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n21606) );
  AOI22_X1 U24596 ( .A1(n21610), .A2(n21607), .B1(n21606), .B2(n21605), .ZN(
        P1_U3481) );
  INV_X1 U24597 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n21609) );
  OAI21_X1 U24598 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(P1_REIP_REG_0__SCAN_IN), 
        .A(n21610), .ZN(n21608) );
  OAI21_X1 U24599 ( .B1(n21610), .B2(n21609), .A(n21608), .ZN(P1_U3482) );
  AOI22_X1 U24600 ( .A1(n21625), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n21884), 
        .B2(n21623), .ZN(P1_U3483) );
  INV_X1 U24601 ( .A(n21611), .ZN(n21614) );
  INV_X1 U24602 ( .A(n21612), .ZN(n21613) );
  OAI211_X1 U24603 ( .C1(n21615), .C2(n21533), .A(n21614), .B(n21613), .ZN(
        n21622) );
  OAI211_X1 U24604 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n21617), .A(n21616), 
        .B(P1_STATE2_REG_2__SCAN_IN), .ZN(n21618) );
  NAND3_X1 U24605 ( .A1(n21622), .A2(n21619), .A3(n21618), .ZN(n21620) );
  OAI21_X1 U24606 ( .B1(n21622), .B2(n21621), .A(n21620), .ZN(P1_U3485) );
  AOI22_X1 U24607 ( .A1(n21625), .A2(n21624), .B1(n21689), .B2(n21623), .ZN(
        P1_U3486) );
  NOR4_X1 U24608 ( .A1(P2_REIP_REG_20__SCAN_IN), .A2(P2_DATAO_REG_2__SCAN_IN), 
        .A3(P3_ADDRESS_REG_9__SCAN_IN), .A4(n15212), .ZN(n21629) );
  NOR4_X1 U24609 ( .A1(P2_ADDRESS_REG_13__SCAN_IN), .A2(n21819), .A3(n21818), 
        .A4(n21826), .ZN(n21628) );
  INV_X1 U24610 ( .A(DATAI_25_), .ZN(n21808) );
  NOR4_X1 U24611 ( .A1(P1_REIP_REG_20__SCAN_IN), .A2(BUF1_REG_7__SCAN_IN), 
        .A3(n21808), .A4(n21849), .ZN(n21627) );
  NOR4_X1 U24612 ( .A1(P1_EAX_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A3(P3_ADDRESS_REG_24__SCAN_IN), 
        .A4(n21805), .ZN(n21626) );
  NAND4_X1 U24613 ( .A1(n21629), .A2(n21628), .A3(n21627), .A4(n21626), .ZN(
        n21645) );
  NOR4_X1 U24614 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A3(BUF2_REG_1__SCAN_IN), .A4(
        n11004), .ZN(n21633) );
  NOR4_X1 U24615 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(
        P3_INSTQUEUE_REG_12__0__SCAN_IN), .A3(P3_ADDRESS_REG_3__SCAN_IN), .A4(
        n21866), .ZN(n21632) );
  NOR4_X1 U24616 ( .A1(P2_REIP_REG_22__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A3(P1_LWORD_REG_7__SCAN_IN), 
        .A4(P3_LWORD_REG_2__SCAN_IN), .ZN(n21631) );
  NOR4_X1 U24617 ( .A1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n10812), .A3(
        n21896), .A4(n21894), .ZN(n21630) );
  NAND4_X1 U24618 ( .A1(n21633), .A2(n21632), .A3(n21631), .A4(n21630), .ZN(
        n21644) );
  NOR4_X1 U24619 ( .A1(P2_EAX_REG_29__SCAN_IN), .A2(P1_EBX_REG_25__SCAN_IN), 
        .A3(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A4(n21696), .ZN(n21637) );
  NOR4_X1 U24620 ( .A1(P2_LWORD_REG_11__SCAN_IN), .A2(n21690), .A3(n21683), 
        .A4(n21689), .ZN(n21636) );
  NOR4_X1 U24621 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n16823), .A3(n21714), .A4(
        n21716), .ZN(n21635) );
  NOR4_X1 U24622 ( .A1(BUF2_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(P3_REIP_REG_6__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n21634) );
  NAND4_X1 U24623 ( .A1(n21637), .A2(n21636), .A3(n21635), .A4(n21634), .ZN(
        n21643) );
  NOR4_X1 U24624 ( .A1(P3_REIP_REG_21__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_12__SCAN_IN), .A3(n21852), .A4(n21835), .ZN(n21641)
         );
  NOR4_X1 U24625 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P2_EBX_REG_9__SCAN_IN), .A3(P2_DATAO_REG_18__SCAN_IN), .A4(n13728), 
        .ZN(n21640) );
  NOR4_X1 U24626 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(
        P1_LWORD_REG_13__SCAN_IN), .A3(P3_EAX_REG_25__SCAN_IN), .A4(n21684), 
        .ZN(n21639) );
  NOR4_X1 U24627 ( .A1(n21840), .A2(n15234), .A3(n15104), .A4(n21838), .ZN(
        n21638) );
  NAND4_X1 U24628 ( .A1(n21641), .A2(n21640), .A3(n21639), .A4(n21638), .ZN(
        n21642) );
  NOR4_X1 U24629 ( .A1(n21645), .A2(n21644), .A3(n21643), .A4(n21642), .ZN(
        n21678) );
  NAND4_X1 U24630 ( .A1(P2_LWORD_REG_1__SCAN_IN), .A2(P1_DATAO_REG_7__SCAN_IN), 
        .A3(n16835), .A4(n21745), .ZN(n21646) );
  NOR3_X1 U24631 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(
        P2_UWORD_REG_11__SCAN_IN), .A3(n21646), .ZN(n21652) );
  NAND4_X1 U24632 ( .A1(P3_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_UWORD_REG_3__SCAN_IN), .A3(n21776), .A4(n21772), .ZN(n21650) );
  NAND4_X1 U24633 ( .A1(P2_DATAO_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUE_REG_14__4__SCAN_IN), .A3(P3_LWORD_REG_12__SCAN_IN), .A4(
        n21765), .ZN(n21649) );
  NAND4_X1 U24634 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_1__2__SCAN_IN), .A3(P3_UWORD_REG_14__SCAN_IN), .A4(
        n13316), .ZN(n21648) );
  NAND4_X1 U24635 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(BS16), .A3(
        n21778), .A4(n21792), .ZN(n21647) );
  NOR4_X1 U24636 ( .A1(n21650), .A2(n21649), .A3(n21648), .A4(n21647), .ZN(
        n21651) );
  AND4_X1 U24637 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_INSTQUEUE_REG_1__0__SCAN_IN), .A3(n21652), .A4(n21651), .ZN(n21676)
         );
  INV_X1 U24638 ( .A(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n21704) );
  NOR4_X1 U24639 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(
        P1_INSTQUEUE_REG_10__6__SCAN_IN), .A3(n21704), .A4(n21653), .ZN(n21675) );
  AND4_X1 U24640 ( .A1(n21654), .A2(P1_ADDRESS_REG_12__SCAN_IN), .A3(
        P3_EAX_REG_1__SCAN_IN), .A4(n21821), .ZN(n21669) );
  NAND4_X1 U24641 ( .A1(n21656), .A2(n21655), .A3(
        P2_INSTQUEUE_REG_8__2__SCAN_IN), .A4(BUF1_REG_27__SCAN_IN), .ZN(n21657) );
  NOR2_X1 U24642 ( .A1(n21658), .A2(n21657), .ZN(n21668) );
  INV_X1 U24643 ( .A(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n21788) );
  NOR4_X1 U24644 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(
        P1_MORE_REG_SCAN_IN), .A3(n21681), .A4(n12613), .ZN(n21659) );
  NAND3_X1 U24645 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n21659), .A3(
        n11096), .ZN(n21660) );
  NOR2_X1 U24646 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n21660), .ZN(n21663) );
  INV_X1 U24647 ( .A(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n21662) );
  INV_X1 U24648 ( .A(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n21661) );
  NAND3_X1 U24649 ( .A1(n21663), .A2(n21662), .A3(n21661), .ZN(n21666) );
  INV_X1 U24650 ( .A(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n21664) );
  NAND4_X1 U24651 ( .A1(n21664), .A2(n21728), .A3(
        P1_INSTQUEUE_REG_0__0__SCAN_IN), .A4(P1_INSTQUEUE_REG_15__7__SCAN_IN), 
        .ZN(n21665) );
  NOR2_X1 U24652 ( .A1(n21666), .A2(n21665), .ZN(n21667) );
  AND3_X1 U24653 ( .A1(n21669), .A2(n21668), .A3(n21667), .ZN(n21674) );
  NAND4_X1 U24654 ( .A1(DATAI_19_), .A2(P3_DATAO_REG_31__SCAN_IN), .A3(n21670), 
        .A4(n21869), .ZN(n21672) );
  NAND4_X1 U24655 ( .A1(P2_EAX_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_12__1__SCAN_IN), .A3(P3_DATAWIDTH_REG_10__SCAN_IN), 
        .A4(n21732), .ZN(n21671) );
  INV_X1 U24656 ( .A(P1_ADDRESS_REG_25__SCAN_IN), .ZN(n21910) );
  NOR3_X1 U24657 ( .A1(n21672), .A2(n21671), .A3(n21910), .ZN(n21673) );
  AND4_X1 U24658 ( .A1(n21676), .A2(n21675), .A3(n21674), .A4(n21673), .ZN(
        n21677) );
  AOI21_X1 U24659 ( .B1(n21678), .B2(n21677), .A(P1_W_R_N_REG_SCAN_IN), .ZN(
        n21926) );
  AOI22_X1 U24660 ( .A1(n21681), .A2(keyinput93), .B1(keyinput92), .B2(n21680), 
        .ZN(n21679) );
  OAI221_X1 U24661 ( .B1(n21681), .B2(keyinput93), .C1(n21680), .C2(keyinput92), .A(n21679), .ZN(n21687) );
  AOI22_X1 U24662 ( .A1(n21684), .A2(keyinput34), .B1(n21683), .B2(keyinput28), 
        .ZN(n21682) );
  OAI221_X1 U24663 ( .B1(n21684), .B2(keyinput34), .C1(n21683), .C2(keyinput28), .A(n21682), .ZN(n21686) );
  XOR2_X1 U24664 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B(keyinput40), .Z(
        n21685) );
  OR3_X1 U24665 ( .A1(n21687), .A2(n21686), .A3(n21685), .ZN(n21694) );
  AOI22_X1 U24666 ( .A1(n21690), .A2(keyinput85), .B1(keyinput71), .B2(n21689), 
        .ZN(n21688) );
  OAI221_X1 U24667 ( .B1(n21690), .B2(keyinput85), .C1(n21689), .C2(keyinput71), .A(n21688), .ZN(n21693) );
  XNOR2_X1 U24668 ( .A(n21691), .B(keyinput79), .ZN(n21692) );
  NOR3_X1 U24669 ( .A1(n21694), .A2(n21693), .A3(n21692), .ZN(n21740) );
  AOI22_X1 U24670 ( .A1(n21697), .A2(keyinput91), .B1(keyinput10), .B2(n21696), 
        .ZN(n21695) );
  OAI221_X1 U24671 ( .B1(n21697), .B2(keyinput91), .C1(n21696), .C2(keyinput10), .A(n21695), .ZN(n21709) );
  AOI22_X1 U24672 ( .A1(n21700), .A2(keyinput19), .B1(keyinput104), .B2(n21699), .ZN(n21698) );
  OAI221_X1 U24673 ( .B1(n21700), .B2(keyinput19), .C1(n21699), .C2(
        keyinput104), .A(n21698), .ZN(n21708) );
  AOI22_X1 U24674 ( .A1(n21702), .A2(keyinput90), .B1(keyinput36), .B2(n13646), 
        .ZN(n21701) );
  OAI221_X1 U24675 ( .B1(n21702), .B2(keyinput90), .C1(n13646), .C2(keyinput36), .A(n21701), .ZN(n21707) );
  AOI22_X1 U24676 ( .A1(n21705), .A2(keyinput31), .B1(n21704), .B2(keyinput4), 
        .ZN(n21703) );
  OAI221_X1 U24677 ( .B1(n21705), .B2(keyinput31), .C1(n21704), .C2(keyinput4), 
        .A(n21703), .ZN(n21706) );
  NOR4_X1 U24678 ( .A1(n21709), .A2(n21708), .A3(n21707), .A4(n21706), .ZN(
        n21739) );
  AOI22_X1 U24679 ( .A1(n21712), .A2(keyinput124), .B1(keyinput75), .B2(n21711), .ZN(n21710) );
  OAI221_X1 U24680 ( .B1(n21712), .B2(keyinput124), .C1(n21711), .C2(
        keyinput75), .A(n21710), .ZN(n21723) );
  AOI22_X1 U24681 ( .A1(n21714), .A2(keyinput70), .B1(n16787), .B2(keyinput74), 
        .ZN(n21713) );
  OAI221_X1 U24682 ( .B1(n21714), .B2(keyinput70), .C1(n16787), .C2(keyinput74), .A(n21713), .ZN(n21722) );
  AOI22_X1 U24683 ( .A1(n16823), .A2(keyinput58), .B1(keyinput16), .B2(n21716), 
        .ZN(n21715) );
  OAI221_X1 U24684 ( .B1(n16823), .B2(keyinput58), .C1(n21716), .C2(keyinput16), .A(n21715), .ZN(n21721) );
  AOI22_X1 U24685 ( .A1(n21719), .A2(keyinput123), .B1(n21718), .B2(keyinput11), .ZN(n21717) );
  OAI221_X1 U24686 ( .B1(n21719), .B2(keyinput123), .C1(n21718), .C2(
        keyinput11), .A(n21717), .ZN(n21720) );
  NOR4_X1 U24687 ( .A1(n21723), .A2(n21722), .A3(n21721), .A4(n21720), .ZN(
        n21738) );
  AOI22_X1 U24688 ( .A1(n21726), .A2(keyinput110), .B1(keyinput32), .B2(n21725), .ZN(n21724) );
  OAI221_X1 U24689 ( .B1(n21726), .B2(keyinput110), .C1(n21725), .C2(
        keyinput32), .A(n21724), .ZN(n21736) );
  AOI22_X1 U24690 ( .A1(n21728), .A2(keyinput118), .B1(n11096), .B2(keyinput81), .ZN(n21727) );
  OAI221_X1 U24691 ( .B1(n21728), .B2(keyinput118), .C1(n11096), .C2(
        keyinput81), .A(n21727), .ZN(n21735) );
  XNOR2_X1 U24692 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(keyinput96), 
        .ZN(n21731) );
  XNOR2_X1 U24693 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B(keyinput5), .ZN(
        n21730) );
  XNOR2_X1 U24694 ( .A(keyinput94), .B(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n21729) );
  NAND3_X1 U24695 ( .A1(n21731), .A2(n21730), .A3(n21729), .ZN(n21734) );
  XNOR2_X1 U24696 ( .A(n21732), .B(keyinput114), .ZN(n21733) );
  NOR4_X1 U24697 ( .A1(n21736), .A2(n21735), .A3(n21734), .A4(n21733), .ZN(
        n21737) );
  NAND4_X1 U24698 ( .A1(n21740), .A2(n21739), .A3(n21738), .A4(n21737), .ZN(
        n21924) );
  AOI22_X1 U24699 ( .A1(n21743), .A2(keyinput127), .B1(keyinput48), .B2(n21742), .ZN(n21741) );
  OAI221_X1 U24700 ( .B1(n21743), .B2(keyinput127), .C1(n21742), .C2(
        keyinput48), .A(n21741), .ZN(n21755) );
  AOI22_X1 U24701 ( .A1(n16835), .A2(keyinput24), .B1(keyinput125), .B2(n21745), .ZN(n21744) );
  OAI221_X1 U24702 ( .B1(n16835), .B2(keyinput24), .C1(n21745), .C2(
        keyinput125), .A(n21744), .ZN(n21754) );
  AOI22_X1 U24703 ( .A1(n21748), .A2(keyinput3), .B1(keyinput46), .B2(n21747), 
        .ZN(n21746) );
  OAI221_X1 U24704 ( .B1(n21748), .B2(keyinput3), .C1(n21747), .C2(keyinput46), 
        .A(n21746), .ZN(n21753) );
  XOR2_X1 U24705 ( .A(n21749), .B(keyinput116), .Z(n21751) );
  XNOR2_X1 U24706 ( .A(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B(keyinput8), .ZN(
        n21750) );
  NAND2_X1 U24707 ( .A1(n21751), .A2(n21750), .ZN(n21752) );
  NOR4_X1 U24708 ( .A1(n21755), .A2(n21754), .A3(n21753), .A4(n21752), .ZN(
        n21802) );
  AOI22_X1 U24709 ( .A1(n11587), .A2(keyinput60), .B1(keyinput83), .B2(n21757), 
        .ZN(n21756) );
  OAI221_X1 U24710 ( .B1(n11587), .B2(keyinput60), .C1(n21757), .C2(keyinput83), .A(n21756), .ZN(n21770) );
  AOI22_X1 U24711 ( .A1(n21760), .A2(keyinput106), .B1(n21759), .B2(keyinput0), 
        .ZN(n21758) );
  OAI221_X1 U24712 ( .B1(n21760), .B2(keyinput106), .C1(n21759), .C2(keyinput0), .A(n21758), .ZN(n21769) );
  AOI22_X1 U24713 ( .A1(n21763), .A2(keyinput35), .B1(keyinput27), .B2(n21762), 
        .ZN(n21761) );
  OAI221_X1 U24714 ( .B1(n21763), .B2(keyinput35), .C1(n21762), .C2(keyinput27), .A(n21761), .ZN(n21768) );
  AOI22_X1 U24715 ( .A1(n21766), .A2(keyinput18), .B1(keyinput43), .B2(n21765), 
        .ZN(n21764) );
  OAI221_X1 U24716 ( .B1(n21766), .B2(keyinput18), .C1(n21765), .C2(keyinput43), .A(n21764), .ZN(n21767) );
  NOR4_X1 U24717 ( .A1(n21770), .A2(n21769), .A3(n21768), .A4(n21767), .ZN(
        n21801) );
  AOI22_X1 U24718 ( .A1(n21773), .A2(keyinput20), .B1(n21772), .B2(keyinput44), 
        .ZN(n21771) );
  OAI221_X1 U24719 ( .B1(n21773), .B2(keyinput20), .C1(n21772), .C2(keyinput44), .A(n21771), .ZN(n21785) );
  AOI22_X1 U24720 ( .A1(n21776), .A2(keyinput66), .B1(keyinput126), .B2(n21775), .ZN(n21774) );
  OAI221_X1 U24721 ( .B1(n21776), .B2(keyinput66), .C1(n21775), .C2(
        keyinput126), .A(n21774), .ZN(n21784) );
  AOI22_X1 U24722 ( .A1(n21779), .A2(keyinput50), .B1(n21778), .B2(keyinput103), .ZN(n21777) );
  OAI221_X1 U24723 ( .B1(n21779), .B2(keyinput50), .C1(n21778), .C2(
        keyinput103), .A(n21777), .ZN(n21783) );
  XOR2_X1 U24724 ( .A(n21662), .B(keyinput95), .Z(n21781) );
  XNOR2_X1 U24725 ( .A(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B(keyinput84), .ZN(
        n21780) );
  NAND2_X1 U24726 ( .A1(n21781), .A2(n21780), .ZN(n21782) );
  NOR4_X1 U24727 ( .A1(n21785), .A2(n21784), .A3(n21783), .A4(n21782), .ZN(
        n21800) );
  AOI22_X1 U24728 ( .A1(n13316), .A2(keyinput65), .B1(keyinput15), .B2(n14165), 
        .ZN(n21786) );
  OAI221_X1 U24729 ( .B1(n13316), .B2(keyinput65), .C1(n14165), .C2(keyinput15), .A(n21786), .ZN(n21798) );
  AOI22_X1 U24730 ( .A1(n21789), .A2(keyinput42), .B1(n21788), .B2(keyinput55), 
        .ZN(n21787) );
  OAI221_X1 U24731 ( .B1(n21789), .B2(keyinput42), .C1(n21788), .C2(keyinput55), .A(n21787), .ZN(n21797) );
  AOI22_X1 U24732 ( .A1(n21792), .A2(keyinput76), .B1(n21791), .B2(keyinput73), 
        .ZN(n21790) );
  OAI221_X1 U24733 ( .B1(n21792), .B2(keyinput76), .C1(n21791), .C2(keyinput73), .A(n21790), .ZN(n21796) );
  XNOR2_X1 U24734 ( .A(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B(keyinput122), .ZN(
        n21794) );
  XNOR2_X1 U24735 ( .A(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B(keyinput30), .ZN(
        n21793) );
  NAND2_X1 U24736 ( .A1(n21794), .A2(n21793), .ZN(n21795) );
  NOR4_X1 U24737 ( .A1(n21798), .A2(n21797), .A3(n21796), .A4(n21795), .ZN(
        n21799) );
  NAND4_X1 U24738 ( .A1(n21802), .A2(n21801), .A3(n21800), .A4(n21799), .ZN(
        n21923) );
  AOI22_X1 U24739 ( .A1(n21805), .A2(keyinput108), .B1(n21804), .B2(keyinput47), .ZN(n21803) );
  OAI221_X1 U24740 ( .B1(n21805), .B2(keyinput108), .C1(n21804), .C2(
        keyinput47), .A(n21803), .ZN(n21816) );
  AOI22_X1 U24741 ( .A1(n11462), .A2(keyinput98), .B1(keyinput68), .B2(n15212), 
        .ZN(n21806) );
  OAI221_X1 U24742 ( .B1(n11462), .B2(keyinput98), .C1(n15212), .C2(keyinput68), .A(n21806), .ZN(n21815) );
  AOI22_X1 U24743 ( .A1(n21809), .A2(keyinput97), .B1(n21808), .B2(keyinput12), 
        .ZN(n21807) );
  OAI221_X1 U24744 ( .B1(n21809), .B2(keyinput97), .C1(n21808), .C2(keyinput12), .A(n21807), .ZN(n21814) );
  AOI22_X1 U24745 ( .A1(n21812), .A2(keyinput121), .B1(n21811), .B2(keyinput62), .ZN(n21810) );
  OAI221_X1 U24746 ( .B1(n21812), .B2(keyinput121), .C1(n21811), .C2(
        keyinput62), .A(n21810), .ZN(n21813) );
  NOR4_X1 U24747 ( .A1(n21816), .A2(n21815), .A3(n21814), .A4(n21813), .ZN(
        n21863) );
  AOI22_X1 U24748 ( .A1(n21819), .A2(keyinput17), .B1(keyinput26), .B2(n21818), 
        .ZN(n21817) );
  OAI221_X1 U24749 ( .B1(n21819), .B2(keyinput17), .C1(n21818), .C2(keyinput26), .A(n21817), .ZN(n21830) );
  AOI22_X1 U24750 ( .A1(n21821), .A2(keyinput120), .B1(n12613), .B2(keyinput61), .ZN(n21820) );
  OAI221_X1 U24751 ( .B1(n21821), .B2(keyinput120), .C1(n12613), .C2(
        keyinput61), .A(n21820), .ZN(n21829) );
  AOI22_X1 U24752 ( .A1(n21661), .A2(keyinput53), .B1(keyinput38), .B2(n21823), 
        .ZN(n21822) );
  OAI221_X1 U24753 ( .B1(n21661), .B2(keyinput53), .C1(n21823), .C2(keyinput38), .A(n21822), .ZN(n21828) );
  AOI22_X1 U24754 ( .A1(n21826), .A2(keyinput39), .B1(keyinput13), .B2(n21825), 
        .ZN(n21824) );
  OAI221_X1 U24755 ( .B1(n21826), .B2(keyinput39), .C1(n21825), .C2(keyinput13), .A(n21824), .ZN(n21827) );
  NOR4_X1 U24756 ( .A1(n21830), .A2(n21829), .A3(n21828), .A4(n21827), .ZN(
        n21862) );
  AOI22_X1 U24757 ( .A1(n21832), .A2(keyinput109), .B1(n15104), .B2(keyinput88), .ZN(n21831) );
  OAI221_X1 U24758 ( .B1(n21832), .B2(keyinput109), .C1(n15104), .C2(
        keyinput88), .A(n21831), .ZN(n21844) );
  AOI22_X1 U24759 ( .A1(n21835), .A2(keyinput115), .B1(keyinput72), .B2(n21834), .ZN(n21833) );
  OAI221_X1 U24760 ( .B1(n21835), .B2(keyinput115), .C1(n21834), .C2(
        keyinput72), .A(n21833), .ZN(n21843) );
  AOI22_X1 U24761 ( .A1(n21838), .A2(keyinput69), .B1(keyinput117), .B2(n21837), .ZN(n21836) );
  OAI221_X1 U24762 ( .B1(n21838), .B2(keyinput69), .C1(n21837), .C2(
        keyinput117), .A(n21836), .ZN(n21842) );
  AOI22_X1 U24763 ( .A1(n21840), .A2(keyinput2), .B1(keyinput9), .B2(n15234), 
        .ZN(n21839) );
  OAI221_X1 U24764 ( .B1(n21840), .B2(keyinput2), .C1(n15234), .C2(keyinput9), 
        .A(n21839), .ZN(n21841) );
  NOR4_X1 U24765 ( .A1(n21844), .A2(n21843), .A3(n21842), .A4(n21841), .ZN(
        n21861) );
  INV_X1 U24766 ( .A(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n21846) );
  AOI22_X1 U24767 ( .A1(n21847), .A2(keyinput23), .B1(keyinput57), .B2(n21846), 
        .ZN(n21845) );
  OAI221_X1 U24768 ( .B1(n21847), .B2(keyinput23), .C1(n21846), .C2(keyinput57), .A(n21845), .ZN(n21859) );
  AOI22_X1 U24769 ( .A1(n21850), .A2(keyinput1), .B1(keyinput67), .B2(n21849), 
        .ZN(n21848) );
  OAI221_X1 U24770 ( .B1(n21850), .B2(keyinput1), .C1(n21849), .C2(keyinput67), 
        .A(n21848), .ZN(n21858) );
  AOI22_X1 U24771 ( .A1(n21853), .A2(keyinput99), .B1(keyinput119), .B2(n21852), .ZN(n21851) );
  OAI221_X1 U24772 ( .B1(n21853), .B2(keyinput99), .C1(n21852), .C2(
        keyinput119), .A(n21851), .ZN(n21857) );
  AOI22_X1 U24773 ( .A1(n13728), .A2(keyinput25), .B1(keyinput7), .B2(n21855), 
        .ZN(n21854) );
  OAI221_X1 U24774 ( .B1(n13728), .B2(keyinput25), .C1(n21855), .C2(keyinput7), 
        .A(n21854), .ZN(n21856) );
  NOR4_X1 U24775 ( .A1(n21859), .A2(n21858), .A3(n21857), .A4(n21856), .ZN(
        n21860) );
  NAND4_X1 U24776 ( .A1(n21863), .A2(n21862), .A3(n21861), .A4(n21860), .ZN(
        n21922) );
  AOI22_X1 U24777 ( .A1(n21866), .A2(keyinput112), .B1(keyinput59), .B2(n21865), .ZN(n21864) );
  OAI221_X1 U24778 ( .B1(n21866), .B2(keyinput112), .C1(n21865), .C2(
        keyinput59), .A(n21864), .ZN(n21877) );
  AOI22_X1 U24779 ( .A1(n21869), .A2(keyinput80), .B1(n21868), .B2(keyinput89), 
        .ZN(n21867) );
  OAI221_X1 U24780 ( .B1(n21869), .B2(keyinput80), .C1(n21868), .C2(keyinput89), .A(n21867), .ZN(n21876) );
  XNOR2_X1 U24781 ( .A(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B(keyinput86), .ZN(
        n21872) );
  XNOR2_X1 U24782 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B(keyinput101), .ZN(
        n21871) );
  XNOR2_X1 U24783 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B(keyinput37), .ZN(
        n21870) );
  NAND3_X1 U24784 ( .A1(n21872), .A2(n21871), .A3(n21870), .ZN(n21875) );
  XNOR2_X1 U24785 ( .A(n21873), .B(keyinput64), .ZN(n21874) );
  NOR4_X1 U24786 ( .A1(n21877), .A2(n21876), .A3(n21875), .A4(n21874), .ZN(
        n21920) );
  INV_X1 U24787 ( .A(DATAI_19_), .ZN(n21880) );
  AOI22_X1 U24788 ( .A1(n21880), .A2(keyinput21), .B1(keyinput6), .B2(n21879), 
        .ZN(n21878) );
  OAI221_X1 U24789 ( .B1(n21880), .B2(keyinput21), .C1(n21879), .C2(keyinput6), 
        .A(n21878), .ZN(n21891) );
  AOI22_X1 U24790 ( .A1(n21883), .A2(keyinput111), .B1(keyinput63), .B2(n21882), .ZN(n21881) );
  OAI221_X1 U24791 ( .B1(n21883), .B2(keyinput111), .C1(n21882), .C2(
        keyinput63), .A(n21881), .ZN(n21890) );
  AOI22_X1 U24792 ( .A1(keyinput14), .A2(n21656), .B1(keyinput49), .B2(n21884), 
        .ZN(n21885) );
  OAI21_X1 U24793 ( .B1(n21656), .B2(keyinput14), .A(n21885), .ZN(n21889) );
  XNOR2_X1 U24794 ( .A(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B(keyinput52), .ZN(
        n21887) );
  XNOR2_X1 U24795 ( .A(keyinput105), .B(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n21886) );
  NAND2_X1 U24796 ( .A1(n21887), .A2(n21886), .ZN(n21888) );
  NOR4_X1 U24797 ( .A1(n21891), .A2(n21890), .A3(n21889), .A4(n21888), .ZN(
        n21919) );
  AOI22_X1 U24798 ( .A1(n21894), .A2(keyinput22), .B1(keyinput29), .B2(n21893), 
        .ZN(n21892) );
  OAI221_X1 U24799 ( .B1(n21894), .B2(keyinput22), .C1(n21893), .C2(keyinput29), .A(n21892), .ZN(n21904) );
  AOI22_X1 U24800 ( .A1(n10812), .A2(keyinput100), .B1(keyinput41), .B2(n21896), .ZN(n21895) );
  OAI221_X1 U24801 ( .B1(n10812), .B2(keyinput100), .C1(n21896), .C2(
        keyinput41), .A(n21895), .ZN(n21903) );
  AOI22_X1 U24802 ( .A1(n13142), .A2(keyinput51), .B1(n21898), .B2(keyinput45), 
        .ZN(n21897) );
  OAI221_X1 U24803 ( .B1(n13142), .B2(keyinput51), .C1(n21898), .C2(keyinput45), .A(n21897), .ZN(n21902) );
  AOI22_X1 U24804 ( .A1(n16949), .A2(keyinput82), .B1(keyinput87), .B2(n21900), 
        .ZN(n21899) );
  OAI221_X1 U24805 ( .B1(n16949), .B2(keyinput82), .C1(n21900), .C2(keyinput87), .A(n21899), .ZN(n21901) );
  NOR4_X1 U24806 ( .A1(n21904), .A2(n21903), .A3(n21902), .A4(n21901), .ZN(
        n21918) );
  AOI22_X1 U24807 ( .A1(n21906), .A2(keyinput33), .B1(n10968), .B2(keyinput107), .ZN(n21905) );
  OAI221_X1 U24808 ( .B1(n21906), .B2(keyinput33), .C1(n10968), .C2(
        keyinput107), .A(n21905), .ZN(n21916) );
  AOI22_X1 U24809 ( .A1(n13632), .A2(keyinput56), .B1(n11004), .B2(keyinput102), .ZN(n21907) );
  OAI221_X1 U24810 ( .B1(n13632), .B2(keyinput56), .C1(n11004), .C2(
        keyinput102), .A(n21907), .ZN(n21915) );
  AOI22_X1 U24811 ( .A1(n21910), .A2(keyinput78), .B1(n21909), .B2(keyinput77), 
        .ZN(n21908) );
  OAI221_X1 U24812 ( .B1(n21910), .B2(keyinput78), .C1(n21909), .C2(keyinput77), .A(n21908), .ZN(n21914) );
  XOR2_X1 U24813 ( .A(n21664), .B(keyinput113), .Z(n21912) );
  XNOR2_X1 U24814 ( .A(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B(keyinput54), .ZN(
        n21911) );
  NAND2_X1 U24815 ( .A1(n21912), .A2(n21911), .ZN(n21913) );
  NOR4_X1 U24816 ( .A1(n21916), .A2(n21915), .A3(n21914), .A4(n21913), .ZN(
        n21917) );
  NAND4_X1 U24817 ( .A1(n21920), .A2(n21919), .A3(n21918), .A4(n21917), .ZN(
        n21921) );
  NOR4_X1 U24818 ( .A1(n21924), .A2(n21923), .A3(n21922), .A4(n21921), .ZN(
        n21925) );
  OAI21_X1 U24819 ( .B1(keyinput49), .B2(n21926), .A(n21925), .ZN(n21939) );
  AOI22_X1 U24820 ( .A1(n21930), .A2(n21929), .B1(n21928), .B2(n21927), .ZN(
        n21935) );
  AOI22_X1 U24821 ( .A1(n21933), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n21932), .B2(n21931), .ZN(n21934) );
  OAI211_X1 U24822 ( .C1(n21937), .C2(n21936), .A(n21935), .B(n21934), .ZN(
        n21938) );
  XNOR2_X1 U24823 ( .A(n21939), .B(n21938), .ZN(P1_U3115) );
  INV_X2 U11597 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11000) );
  AND2_X1 U11295 ( .A1(n14443), .A2(n13950), .ZN(n11797) );
  NAND2_X1 U13100 ( .A1(n10727), .A2(n9861), .ZN(n11202) );
  NAND4_X1 U15172 ( .A1(n11863), .A2(n11854), .A3(n11891), .A4(n13440), .ZN(
        n14459) );
  CLKBUF_X1 U11151 ( .A(n9691), .Z(n9706) );
  OR2_X1 U13386 ( .A1(n11600), .A2(n11599), .ZN(n10372) );
  NOR2_X1 U11252 ( .A1(n16905), .A2(n10406), .ZN(n17208) );
  AND2_X1 U11186 ( .A1(n10732), .A2(n10734), .ZN(n10721) );
  AND2_X1 U11193 ( .A1(n11741), .A2(n14443), .ZN(n11823) );
  CLKBUF_X1 U11200 ( .A(n10726), .Z(n12821) );
  CLKBUF_X1 U11287 ( .A(n11223), .Z(n12779) );
  CLKBUF_X1 U11519 ( .A(n14864), .Z(n14875) );
  CLKBUF_X1 U11621 ( .A(n10784), .Z(n10797) );
  CLKBUF_X1 U12289 ( .A(n11229), .Z(n9702) );
  CLKBUF_X1 U12779 ( .A(n11009), .Z(n12958) );
  CLKBUF_X1 U13948 ( .A(n11869), .Z(n12634) );
  CLKBUF_X1 U15094 ( .A(n14901), .Z(n14902) );
  INV_X1 U18576 ( .A(n10734), .ZN(n11170) );
endmodule

