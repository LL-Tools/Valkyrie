

module b21_C_2inp_gates_syn ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, 
        ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, 
        ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, 
        ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, 
        ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, P1_U3352, P1_U3351, 
        P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, 
        P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, 
        P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, 
        P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, 
        P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, 
        P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, 
        P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, 
        P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, 
        P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, 
        P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, 
        P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, 
        P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, 
        P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, 
        P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, 
        P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, 
        P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, 
        P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, 
        P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, 
        P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, 
        P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, 
        P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, 
        P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, 
        P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, 
        P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, 
        P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, 
        P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, 
        P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, 
        P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, 
        P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, 
        P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, 
        P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, 
        P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, 
        P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, 
        P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, 
        P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, 
        P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, 
        P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, 
        P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, 
        P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, 
        P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, 
        P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, 
        P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, 
        P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, 
        P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, 
        P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, 
        P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, 
        P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, 
        P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3152, P2_U3151, P2_U3966, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9382, n9383,
         n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393,
         n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403,
         n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413,
         n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423,
         n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433,
         n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443,
         n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453,
         n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463,
         n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473,
         n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483,
         n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493,
         n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503,
         n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513,
         n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523,
         n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533,
         n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543,
         n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553,
         n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563,
         n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573,
         n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583,
         n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593,
         n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603,
         n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613,
         n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623,
         n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633,
         n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643,
         n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653,
         n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663,
         n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673,
         n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683,
         n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693,
         n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703,
         n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713,
         n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723,
         n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733,
         n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743,
         n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753,
         n9754, n9755, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764,
         n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774,
         n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784,
         n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794,
         n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804,
         n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814,
         n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824,
         n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834,
         n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844,
         n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854,
         n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864,
         n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874,
         n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884,
         n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894,
         n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904,
         n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914,
         n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924,
         n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934,
         n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944,
         n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954,
         n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964,
         n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974,
         n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984,
         n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994,
         n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003,
         n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011,
         n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019,
         n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027,
         n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035,
         n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043,
         n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051,
         n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059,
         n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067,
         n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075,
         n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083,
         n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091,
         n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099,
         n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107,
         n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115,
         n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123,
         n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131,
         n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139,
         n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147,
         n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155,
         n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163,
         n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171,
         n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179,
         n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187,
         n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195,
         n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203,
         n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211,
         n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219,
         n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227,
         n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235,
         n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243,
         n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251,
         n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259,
         n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267,
         n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275,
         n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283,
         n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291,
         n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299,
         n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307,
         n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315,
         n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323,
         n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331,
         n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339,
         n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347,
         n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355,
         n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363,
         n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371,
         n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379,
         n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387,
         n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395,
         n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403,
         n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411,
         n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419,
         n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427,
         n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435,
         n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443,
         n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451,
         n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459,
         n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467,
         n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475,
         n10476, n10477, n10478;

  NAND2_X1 U4878 ( .A1(n9152), .A2(n9222), .ZN(n9212) );
  INV_X1 U4879 ( .A(n9702), .ZN(n4379) );
  NAND2_X1 U4880 ( .A1(n8986), .A2(n8765), .ZN(n8900) );
  XNOR2_X1 U4881 ( .A(n5634), .B(n5633), .ZN(n8132) );
  INV_X1 U4882 ( .A(n10158), .ZN(n10011) );
  INV_X1 U4883 ( .A(n6800), .ZN(n6871) );
  AND2_X1 U4884 ( .A1(n7373), .A2(n5002), .ZN(n4422) );
  INV_X1 U4885 ( .A(n6382), .ZN(n6246) );
  INV_X1 U4886 ( .A(n7422), .ZN(n7372) );
  INV_X2 U4887 ( .A(n5877), .ZN(n5911) );
  BUF_X2 U4888 ( .A(n7007), .Z(n4376) );
  INV_X2 U4889 ( .A(n5581), .ZN(n5635) );
  CLKBUF_X3 U4890 ( .A(n5538), .Z(n4375) );
  INV_X1 U4891 ( .A(n7543), .ZN(n5926) );
  INV_X1 U4892 ( .A(n9361), .ZN(n7537) );
  AND2_X1 U4893 ( .A1(n5537), .A2(n5764), .ZN(n9361) );
  NAND2_X1 U4894 ( .A1(n5768), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5770) );
  NAND4_X1 U4895 ( .A1(n5970), .A2(n5969), .A3(n6018), .A4(n5968), .ZN(n5971)
         );
  AOI21_X1 U4896 ( .B1(n9850), .B2(n10087), .A(n10334), .ZN(n4570) );
  AND4_X1 U4897 ( .A1(n6203), .A2(n6188), .A3(n6186), .A4(n6168), .ZN(n5970)
         );
  NOR2_X1 U4898 ( .A1(n8804), .A2(n4889), .ZN(n8949) );
  OAI21_X1 U4899 ( .B1(n4379), .B2(n4669), .A(n4671), .ZN(n6870) );
  INV_X1 U4900 ( .A(n6139), .ZN(n4798) );
  NOR2_X1 U4901 ( .A1(n5063), .A2(n9398), .ZN(n5062) );
  AND2_X1 U4902 ( .A1(n8613), .A2(n5836), .ZN(n4748) );
  NAND2_X1 U4903 ( .A1(n5282), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5321) );
  OR2_X1 U4904 ( .A1(n10394), .A2(n9035), .ZN(n5779) );
  BUF_X1 U4905 ( .A(n5298), .Z(n5454) );
  INV_X2 U4906 ( .A(n6977), .ZN(n6245) );
  NAND2_X1 U4907 ( .A1(n9933), .A2(n9910), .ZN(n9906) );
  NAND2_X1 U4908 ( .A1(n4400), .A2(n7372), .ZN(n7470) );
  OR2_X1 U4909 ( .A1(n5495), .A2(n8989), .ZN(n5542) );
  INV_X1 U4911 ( .A(n6913), .ZN(n6734) );
  NOR2_X1 U4912 ( .A1(n9906), .A2(n5053), .ZN(n9864) );
  NAND3_X1 U4913 ( .A1(n6585), .A2(n6584), .A3(n7447), .ZN(n7442) );
  AND2_X1 U4914 ( .A1(n9851), .A2(n9850), .ZN(n10101) );
  INV_X1 U4915 ( .A(n7711), .ZN(n10333) );
  AND2_X1 U4916 ( .A1(n7138), .A2(n7554), .ZN(n7564) );
  AND4_X1 U4917 ( .A1(n5271), .A2(n5270), .A3(n5269), .A4(n5268), .ZN(n7671)
         );
  NAND2_X1 U4918 ( .A1(n8862), .A2(n7757), .ZN(n7554) );
  AND4_X1 U4919 ( .A1(n6112), .A2(n6111), .A3(n6110), .A4(n6109), .ZN(n8207)
         );
  NAND2_X1 U4920 ( .A1(n10086), .A2(n9841), .ZN(n10082) );
  AOI21_X1 U4921 ( .B1(n8842), .B2(n10099), .A(n8841), .ZN(n10109) );
  AND2_X1 U4922 ( .A1(n6908), .A2(n7323), .ZN(n10057) );
  XNOR2_X1 U4923 ( .A(n5620), .B(n5647), .ZN(n8518) );
  INV_X1 U4924 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n6188) );
  INV_X1 U4925 ( .A(n4399), .ZN(n6964) );
  NAND2_X1 U4926 ( .A1(n4580), .A2(n10268), .ZN(n10269) );
  AND4_X1 U4927 ( .A1(n5247), .A2(n5248), .A3(n5249), .A4(n5246), .ZN(n7782)
         );
  XNOR2_X1 U4928 ( .A(n5132), .B(n9585), .ZN(n8857) );
  NAND4_X1 U4929 ( .A1(n6069), .A2(n6068), .A3(n6067), .A4(n6066), .ZN(n9777)
         );
  INV_X1 U4931 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5133) );
  INV_X1 U4932 ( .A(n5207), .ZN(n5538) );
  AND2_X1 U4933 ( .A1(n4432), .A2(n4926), .ZN(n4373) );
  OAI21_X2 U4934 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10437), .ZN(n10435) );
  NAND2_X1 U4935 ( .A1(n5138), .A2(n8693), .ZN(n4374) );
  NAND2_X2 U4936 ( .A1(n5138), .A2(n8693), .ZN(n5260) );
  NAND2_X1 U4937 ( .A1(n9358), .A2(n4994), .ZN(n4991) );
  NAND2_X1 U4938 ( .A1(n5430), .A2(n5429), .ZN(n5448) );
  NAND2_X2 U4939 ( .A1(n8500), .A2(n8511), .ZN(n8499) );
  NAND2_X2 U4940 ( .A1(n7355), .A2(n5780), .ZN(n8500) );
  OAI21_X2 U4941 ( .B1(n10054), .B2(n6657), .A(n6656), .ZN(n10034) );
  AOI21_X2 U4942 ( .B1(n8617), .B2(n9054), .A(n9053), .ZN(n9077) );
  NOR2_X2 U4943 ( .A1(n8679), .A2(n8678), .ZN(n9053) );
  XNOR2_X2 U4944 ( .A(n9067), .B(n9068), .ZN(n9060) );
  OAI21_X2 U4945 ( .B1(P2_REG1_REG_14__SCAN_IN), .B2(n9059), .A(n9058), .ZN(
        n9067) );
  AND2_X2 U4946 ( .A1(n6102), .A2(n4434), .ZN(n7046) );
  NAND2_X2 U4947 ( .A1(n4635), .A2(n4633), .ZN(n9474) );
  OAI21_X1 U4948 ( .B1(n5815), .B2(n4591), .A(n4590), .ZN(n4589) );
  NAND2_X2 U4949 ( .A1(n8076), .A2(n8075), .ZN(n8550) );
  NOR2_X1 U4950 ( .A1(n9055), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n9079) );
  XNOR2_X2 U4951 ( .A(n5985), .B(n5981), .ZN(n10245) );
  NAND2_X2 U4952 ( .A1(n7967), .A2(n4583), .ZN(n8076) );
  OAI21_X2 U4953 ( .B1(n5015), .B2(n5014), .A(n5012), .ZN(n5309) );
  NAND2_X2 U4954 ( .A1(n4987), .A2(n7789), .ZN(n7932) );
  NAND2_X2 U4955 ( .A1(n7784), .A2(n7783), .ZN(n7789) );
  NAND2_X2 U4956 ( .A1(n4991), .A2(n4992), .ZN(n9304) );
  INV_X1 U4957 ( .A(n9777), .ZN(n7484) );
  AND2_X4 U4958 ( .A1(n5002), .A2(n6974), .ZN(n6918) );
  OAI21_X1 U4959 ( .B1(n9205), .B2(n4983), .A(n4466), .ZN(n9446) );
  AOI21_X2 U4960 ( .B1(n7229), .B2(P2_REG1_REG_4__SCAN_IN), .A(n7270), .ZN(
        n7284) );
  NOR4_X2 U4961 ( .A1(n6453), .A2(n6688), .A3(n6452), .A4(n6451), .ZN(n6570)
         );
  XNOR2_X2 U4962 ( .A(n5770), .B(n5769), .ZN(n8862) );
  NAND2_X2 U4963 ( .A1(n7932), .A2(n7790), .ZN(n7985) );
  XNOR2_X2 U4964 ( .A(n4838), .B(n6035), .ZN(n7006) );
  AND2_X1 U4965 ( .A1(n4381), .A2(n9859), .ZN(n10104) );
  NAND2_X1 U4966 ( .A1(n4383), .A2(n4378), .ZN(n10105) );
  INV_X1 U4967 ( .A(n10098), .ZN(n4378) );
  NAND2_X1 U4968 ( .A1(n4572), .A2(n9151), .ZN(n9205) );
  NAND2_X1 U4969 ( .A1(n9854), .A2(n4941), .ZN(n4940) );
  NAND2_X1 U4970 ( .A1(n5892), .A2(n5890), .ZN(n9208) );
  NOR2_X1 U4971 ( .A1(n9079), .A2(n9080), .ZN(n9083) );
  NAND2_X1 U4972 ( .A1(n9495), .A2(n9349), .ZN(n9309) );
  AND2_X1 U4973 ( .A1(n6273), .A2(n6272), .ZN(n10131) );
  NAND2_X1 U4974 ( .A1(n7536), .A2(n5635), .ZN(n4618) );
  NAND2_X1 U4975 ( .A1(n6643), .A2(n6543), .ZN(n7514) );
  INV_X4 U4976 ( .A(n4422), .ZN(n6806) );
  NAND4_X1 U4977 ( .A1(n6579), .A2(n6578), .A3(n6577), .A4(n6576), .ZN(n6580)
         );
  BUF_X2 U4978 ( .A(n6266), .Z(n4380) );
  NAND4_X2 U4980 ( .A1(n5174), .A2(n5176), .A3(n5175), .A4(n5177), .ZN(n7141)
         );
  CLKBUF_X1 U4981 ( .A(n7322), .Z(n4594) );
  INV_X1 U4982 ( .A(n5260), .ZN(n5482) );
  INV_X1 U4983 ( .A(n7595), .ZN(n5070) );
  BUF_X1 U4984 ( .A(n5244), .Z(n4394) );
  INV_X2 U4985 ( .A(n5581), .ZN(n5183) );
  CLKBUF_X2 U4986 ( .A(n5227), .Z(n5285) );
  NAND2_X1 U4988 ( .A1(n5138), .A2(n5136), .ZN(n5244) );
  NAND2_X2 U4989 ( .A1(n7169), .A2(n7168), .ZN(n7249) );
  NAND4_X1 U4990 ( .A1(n5948), .A2(n5129), .A3(n5127), .A4(n5128), .ZN(n5143)
         );
  NOR2_X1 U4991 ( .A1(P2_IR_REG_26__SCAN_IN), .A2(P2_IR_REG_25__SCAN_IN), .ZN(
        n5127) );
  INV_X1 U4992 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n6050) );
  OAI211_X1 U4993 ( .C1(n10105), .C2(n10188), .A(n10104), .B(n10103), .ZN(
        n10216) );
  AOI21_X1 U4994 ( .B1(n9877), .B2(n10099), .A(n9876), .ZN(n10114) );
  NAND2_X1 U4995 ( .A1(n4382), .A2(n10099), .ZN(n4381) );
  NOR2_X1 U4996 ( .A1(n4568), .A2(n4567), .ZN(n4566) );
  OR2_X1 U4997 ( .A1(n10110), .A2(n10188), .ZN(n4573) );
  NOR2_X1 U4998 ( .A1(n9157), .A2(n9439), .ZN(n9158) );
  NAND2_X1 U4999 ( .A1(n9182), .A2(n9181), .ZN(n9450) );
  NAND2_X1 U5000 ( .A1(n6896), .A2(n6895), .ZN(n9740) );
  XNOR2_X1 U5001 ( .A(n9160), .B(n9159), .ZN(n9164) );
  OAI21_X1 U5002 ( .B1(n9863), .B2(n4942), .A(n4384), .ZN(n4383) );
  AND2_X1 U5003 ( .A1(n8808), .A2(n8807), .ZN(n4513) );
  AOI21_X1 U5004 ( .B1(n4548), .B2(n10099), .A(n4546), .ZN(n10119) );
  AOI21_X1 U5005 ( .B1(n4944), .B2(n4403), .A(n6623), .ZN(n8832) );
  INV_X1 U5006 ( .A(n9739), .ZN(n6896) );
  NAND2_X1 U5007 ( .A1(n9205), .A2(n9208), .ZN(n4986) );
  BUF_X1 U5008 ( .A(n9862), .Z(n9863) );
  AND2_X1 U5009 ( .A1(n5941), .A2(n7091), .ZN(n4508) );
  AND2_X1 U5010 ( .A1(n6517), .A2(n6400), .ZN(n6562) );
  NAND2_X1 U5011 ( .A1(n4890), .A2(n8801), .ZN(n8804) );
  OAI21_X2 U5012 ( .B1(n9892), .B2(n6620), .A(n6619), .ZN(n9881) );
  OR2_X1 U5013 ( .A1(n6441), .A2(n6516), .ZN(n6442) );
  AND2_X1 U5014 ( .A1(n9155), .A2(n4981), .ZN(n4980) );
  NAND2_X1 U5015 ( .A1(n6870), .A2(n5023), .ZN(n5022) );
  NAND2_X1 U5016 ( .A1(n9250), .A2(n9254), .ZN(n9249) );
  AND2_X1 U5017 ( .A1(n5066), .A2(n9189), .ZN(n9183) );
  NOR3_X1 U5018 ( .A1(n9212), .A2(n9432), .A3(n5064), .ZN(n9133) );
  NAND2_X1 U5019 ( .A1(n4417), .A2(n9854), .ZN(n4939) );
  NAND2_X1 U5020 ( .A1(n4571), .A2(n5918), .ZN(n9250) );
  AOI21_X1 U5021 ( .B1(n4673), .B2(n4672), .A(n4430), .ZN(n4671) );
  NOR2_X1 U5022 ( .A1(n4417), .A2(n9854), .ZN(n4384) );
  AND2_X1 U5023 ( .A1(n4388), .A2(n4386), .ZN(n4385) );
  OAI21_X1 U5024 ( .B1(n4428), .B2(n4697), .A(n4695), .ZN(n4694) );
  NOR2_X1 U5025 ( .A1(n4531), .A2(n5052), .ZN(n9882) );
  INV_X1 U5026 ( .A(n4669), .ZN(n4673) );
  NAND2_X1 U5027 ( .A1(n4388), .A2(n4387), .ZN(n4389) );
  AND2_X1 U5028 ( .A1(n9858), .A2(n9857), .ZN(n9859) );
  NAND2_X1 U5029 ( .A1(n9968), .A2(n6615), .ZN(n4388) );
  AOI21_X1 U5030 ( .B1(n6343), .B2(n6342), .A(n6341), .ZN(n6356) );
  OAI21_X1 U5031 ( .B1(n5003), .B2(n4408), .A(n6849), .ZN(n4669) );
  NAND2_X1 U5032 ( .A1(n8763), .A2(n8982), .ZN(n8986) );
  NAND2_X1 U5033 ( .A1(n5737), .A2(n5736), .ZN(n9432) );
  OAI21_X1 U5034 ( .B1(n6660), .B2(n6484), .A(n4406), .ZN(n4960) );
  NAND2_X1 U5035 ( .A1(n5004), .A2(n6839), .ZN(n5003) );
  AND2_X1 U5036 ( .A1(n5058), .A2(n5057), .ZN(n5056) );
  NOR2_X1 U5037 ( .A1(n9242), .A2(n5034), .ZN(n5033) );
  NAND2_X1 U5038 ( .A1(n6680), .A2(n6682), .ZN(n9871) );
  OR2_X1 U5039 ( .A1(n10116), .A2(n9744), .ZN(n9869) );
  NAND2_X1 U5040 ( .A1(n10116), .A2(n9744), .ZN(n6679) );
  AND2_X1 U5041 ( .A1(n9291), .A2(n5874), .ZN(n9274) );
  AND2_X1 U5042 ( .A1(n5883), .A2(n5879), .ZN(n9254) );
  OR2_X1 U5043 ( .A1(n10121), .A2(n9652), .ZN(n6677) );
  NOR2_X2 U5044 ( .A1(n9320), .A2(n9489), .ZN(n9305) );
  NAND2_X2 U5045 ( .A1(n6316), .A2(n6315), .ZN(n10116) );
  OR2_X1 U5046 ( .A1(n6838), .A2(n9676), .ZN(n6839) );
  AND2_X1 U5047 ( .A1(n6675), .A2(n6414), .ZN(n9916) );
  CLKBUF_X1 U5048 ( .A(n10027), .Z(n4532) );
  INV_X1 U5049 ( .A(n6340), .ZN(n6680) );
  NAND2_X1 U5050 ( .A1(n5637), .A2(n5636), .ZN(n9468) );
  NAND2_X1 U5051 ( .A1(n8518), .A2(n6381), .ZN(n6316) );
  NAND2_X2 U5052 ( .A1(n6293), .A2(n6292), .ZN(n10121) );
  OR2_X1 U5053 ( .A1(n5569), .A2(n5570), .ZN(n9275) );
  OR2_X1 U5054 ( .A1(n10126), .A2(n9720), .ZN(n6675) );
  CLKBUF_X1 U5055 ( .A(n8549), .Z(n4510) );
  NAND2_X1 U5056 ( .A1(n8132), .A2(n6381), .ZN(n6293) );
  AOI21_X1 U5057 ( .B1(n5847), .B2(n5846), .A(n9388), .ZN(n5848) );
  NAND2_X1 U5058 ( .A1(n6303), .A2(n6302), .ZN(n10126) );
  NOR2_X1 U5059 ( .A1(n10144), .A2(n9979), .ZN(n6616) );
  AND2_X1 U5060 ( .A1(n4390), .A2(n10035), .ZN(n6612) );
  NAND2_X2 U5061 ( .A1(n5563), .A2(n9309), .ZN(n9328) );
  NAND2_X1 U5062 ( .A1(n5615), .A2(n5648), .ZN(n5620) );
  AND2_X1 U5063 ( .A1(n5062), .A2(n9345), .ZN(n5061) );
  OR2_X1 U5064 ( .A1(n9489), .A2(n8918), .ZN(n9292) );
  NAND2_X1 U5065 ( .A1(n5632), .A2(n5600), .ZN(n8018) );
  NAND2_X1 U5066 ( .A1(n5516), .A2(n5515), .ZN(n9489) );
  NAND2_X1 U5067 ( .A1(n6254), .A2(n6253), .ZN(n10144) );
  NAND2_X1 U5068 ( .A1(n8607), .A2(n6606), .ZN(n4390) );
  AOI21_X1 U5069 ( .B1(n4748), .B2(n5932), .A(n4746), .ZN(n4745) );
  NAND2_X1 U5070 ( .A1(n6248), .A2(n6247), .ZN(n10148) );
  NAND2_X1 U5071 ( .A1(n4618), .A2(n5540), .ZN(n9495) );
  NOR2_X1 U5072 ( .A1(n6662), .A2(n4959), .ZN(n4958) );
  AND2_X1 U5073 ( .A1(n9345), .A2(n9333), .ZN(n9329) );
  OR2_X1 U5074 ( .A1(n6610), .A2(n6609), .ZN(n10035) );
  OR2_X1 U5075 ( .A1(n9508), .A2(n9522), .ZN(n5063) );
  AND2_X1 U5076 ( .A1(n8184), .A2(n5827), .ZN(n5074) );
  OR2_X1 U5077 ( .A1(n9508), .A2(n9387), .ZN(n5849) );
  OR2_X1 U5078 ( .A1(n8554), .A2(n8553), .ZN(n5100) );
  INV_X1 U5079 ( .A(n8613), .ZN(n8622) );
  INV_X1 U5080 ( .A(n8179), .ZN(n8184) );
  NAND2_X1 U5081 ( .A1(n8095), .A2(n8096), .ZN(n8607) );
  NAND2_X1 U5082 ( .A1(n5492), .A2(n5491), .ZN(n9508) );
  NAND2_X1 U5083 ( .A1(n6263), .A2(n6262), .ZN(n10140) );
  NAND2_X1 U5084 ( .A1(n5036), .A2(n5552), .ZN(n9484) );
  AND2_X1 U5085 ( .A1(n8179), .A2(n8176), .ZN(n8554) );
  AND2_X1 U5086 ( .A1(n6822), .A2(n6821), .ZN(n9700) );
  NAND2_X1 U5087 ( .A1(n6218), .A2(n6217), .ZN(n10158) );
  OR2_X1 U5088 ( .A1(n10164), .A2(n9759), .ZN(n6464) );
  NAND2_X1 U5089 ( .A1(n5834), .A2(n5828), .ZN(n8179) );
  NAND2_X1 U5090 ( .A1(n6234), .A2(n6233), .ZN(n10154) );
  NAND2_X1 U5091 ( .A1(n8683), .A2(n8682), .ZN(n8684) );
  INV_X1 U5092 ( .A(n9280), .ZN(n9313) );
  XNOR2_X1 U5093 ( .A(n5532), .B(n5531), .ZN(n7536) );
  OR2_X1 U5094 ( .A1(n9398), .A2(n9027), .ZN(n5850) );
  AND2_X1 U5095 ( .A1(n5845), .A2(n5844), .ZN(n9408) );
  OR2_X1 U5096 ( .A1(n9526), .A2(n9012), .ZN(n5839) );
  OR2_X1 U5097 ( .A1(n5576), .A2(n5575), .ZN(n4732) );
  NAND2_X1 U5098 ( .A1(n7798), .A2(n5923), .ZN(n5079) );
  XNOR2_X1 U5099 ( .A(n5486), .B(n5487), .ZN(n7296) );
  NAND2_X1 U5100 ( .A1(n6205), .A2(n6204), .ZN(n10164) );
  NAND2_X1 U5101 ( .A1(n6157), .A2(n6156), .ZN(n10174) );
  NAND2_X1 U5102 ( .A1(n5067), .A2(n8973), .ZN(n5834) );
  INV_X1 U5103 ( .A(n10048), .ZN(n10168) );
  NAND2_X1 U5104 ( .A1(n10184), .A2(n9706), .ZN(n8597) );
  OAI21_X1 U5105 ( .B1(n7945), .B2(n6604), .A(n6603), .ZN(n8095) );
  AOI21_X1 U5106 ( .B1(n4684), .B2(n4683), .A(n4457), .ZN(n4682) );
  INV_X1 U5107 ( .A(n8590), .ZN(n10184) );
  NAND2_X1 U5108 ( .A1(n5438), .A2(n5437), .ZN(n9522) );
  AND2_X1 U5109 ( .A1(n6192), .A2(n6191), .ZN(n10048) );
  INV_X1 U5110 ( .A(n8723), .ZN(n9531) );
  NAND2_X1 U5111 ( .A1(n5603), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5638) );
  NAND2_X1 U5112 ( .A1(n4516), .A2(n4735), .ZN(n7798) );
  AND2_X1 U5113 ( .A1(n5390), .A2(n5389), .ZN(n8723) );
  INV_X1 U5114 ( .A(n5605), .ZN(n5603) );
  NAND2_X2 U5115 ( .A1(n6170), .A2(n6169), .ZN(n10178) );
  AND2_X1 U5116 ( .A1(n6125), .A2(n6124), .ZN(n8590) );
  XNOR2_X1 U5117 ( .A(n5402), .B(n5423), .ZN(n7113) );
  AND2_X1 U5118 ( .A1(n4912), .A2(n4911), .ZN(n8141) );
  OAI21_X2 U5119 ( .B1(n7893), .B2(n6599), .A(n6598), .ZN(n8034) );
  NAND2_X1 U5120 ( .A1(n5448), .A2(n5446), .ZN(n4703) );
  OAI21_X1 U5121 ( .B1(n5448), .B2(n5447), .A(n5446), .ZN(n5467) );
  NOR2_X1 U5122 ( .A1(n6763), .A2(n4690), .ZN(n4689) );
  OR2_X1 U5123 ( .A1(n10196), .A2(n7950), .ZN(n6649) );
  OR2_X1 U5124 ( .A1(n6763), .A2(n6764), .ZN(n4688) );
  NOR2_X2 U5125 ( .A1(n7837), .A2(n10201), .ZN(n8039) );
  XNOR2_X1 U5126 ( .A(n5400), .B(n5399), .ZN(n7109) );
  NAND2_X1 U5127 ( .A1(n5351), .A2(n5350), .ZN(n9541) );
  AND2_X1 U5128 ( .A1(n9547), .A2(n8159), .ZN(n5818) );
  NAND2_X1 U5129 ( .A1(n6142), .A2(n6141), .ZN(n7958) );
  AOI21_X1 U5130 ( .B1(n4874), .B2(n4876), .A(n4446), .ZN(n4873) );
  NAND2_X1 U5131 ( .A1(n5979), .A2(n5978), .ZN(n10196) );
  OR2_X1 U5132 ( .A1(n6762), .A2(n6761), .ZN(n6763) );
  OAI21_X1 U5133 ( .B1(n5426), .B2(n5425), .A(n5095), .ZN(n5430) );
  NAND2_X1 U5134 ( .A1(n5426), .A2(n5418), .ZN(n5400) );
  AND2_X2 U5135 ( .A1(n6698), .A2(n7848), .ZN(n5045) );
  NAND2_X1 U5136 ( .A1(n8060), .A2(n4444), .ZN(n7997) );
  NAND2_X1 U5137 ( .A1(n5811), .A2(n5812), .ZN(n7988) );
  XNOR2_X1 U5138 ( .A(n5345), .B(n5089), .ZN(n6995) );
  OR2_X1 U5139 ( .A1(n9775), .A2(n7748), .ZN(n6643) );
  OR2_X1 U5140 ( .A1(n10206), .A2(n8530), .ZN(n6646) );
  NAND2_X1 U5141 ( .A1(n6000), .A2(n5999), .ZN(n10201) );
  NAND2_X1 U5142 ( .A1(n5302), .A2(n5301), .ZN(n9552) );
  NAND2_X1 U5143 ( .A1(n5281), .A2(n5280), .ZN(n10407) );
  NAND2_X1 U5144 ( .A1(n6012), .A2(n6011), .ZN(n10206) );
  AND2_X1 U5145 ( .A1(n6115), .A2(n6114), .ZN(n7748) );
  NAND2_X1 U5146 ( .A1(n6585), .A2(n6584), .ZN(n7443) );
  NAND2_X1 U5147 ( .A1(n8506), .A2(n7671), .ZN(n5805) );
  OR2_X1 U5148 ( .A1(n9776), .A2(n10345), .ZN(n6497) );
  XNOR2_X1 U5149 ( .A(n5291), .B(n5014), .ZN(n6962) );
  NAND2_X1 U5150 ( .A1(n5259), .A2(n5258), .ZN(n8506) );
  AND2_X2 U5151 ( .A1(n7420), .A2(n6918), .ZN(n6913) );
  AND2_X1 U5152 ( .A1(n4976), .A2(n4478), .ZN(n7848) );
  AND2_X2 U5153 ( .A1(n5779), .A2(n7350), .ZN(n8065) );
  NOR2_X1 U5154 ( .A1(n7874), .A2(n7533), .ZN(n8058) );
  INV_X1 U5155 ( .A(n8207), .ZN(n9775) );
  NAND2_X1 U5156 ( .A1(n5243), .A2(n4754), .ZN(n4809) );
  NAND2_X1 U5157 ( .A1(n4841), .A2(n4445), .ZN(n7077) );
  NAND2_X1 U5158 ( .A1(n5164), .A2(n5163), .ZN(n5790) );
  OR2_X1 U5159 ( .A1(n9779), .A2(n7458), .ZN(n7702) );
  INV_X1 U5160 ( .A(n6696), .ZN(n4400) );
  NAND4_X2 U5162 ( .A1(n6098), .A2(n6097), .A3(n6096), .A4(n6095), .ZN(n9776)
         );
  NAND2_X1 U5163 ( .A1(n5071), .A2(n5070), .ZN(n7594) );
  NAND2_X1 U5164 ( .A1(n5256), .A2(n5255), .ZN(n5275) );
  NAND2_X1 U5165 ( .A1(n4612), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5412) );
  OR2_X1 U5166 ( .A1(n7027), .A2(n4842), .ZN(n4841) );
  NAND2_X1 U5167 ( .A1(n9035), .A2(n10394), .ZN(n7350) );
  AND4_X1 U5168 ( .A1(n6579), .A2(n6578), .A3(n6577), .A4(n6576), .ZN(n7483)
         );
  OR2_X1 U5169 ( .A1(n7872), .A2(n10389), .ZN(n7874) );
  XNOR2_X1 U5170 ( .A(n6024), .B(P1_IR_REG_22__SCAN_IN), .ZN(n6688) );
  NAND4_X2 U5171 ( .A1(n5231), .A2(n5230), .A3(n5229), .A4(n5228), .ZN(n9035)
         );
  INV_X1 U5172 ( .A(n9036), .ZN(n5164) );
  NAND2_X2 U5173 ( .A1(n7315), .A2(n4895), .ZN(n8788) );
  AND3_X1 U5174 ( .A1(n6064), .A2(n6063), .A3(n6062), .ZN(n7458) );
  INV_X1 U5175 ( .A(n5393), .ZN(n4612) );
  NAND4_X1 U5176 ( .A1(n6058), .A2(n6057), .A3(n6056), .A4(n6055), .ZN(n9779)
         );
  NAND2_X1 U5177 ( .A1(n6520), .A2(n7625), .ZN(n5002) );
  INV_X1 U5178 ( .A(n7318), .ZN(n5071) );
  OAI211_X1 U5179 ( .C1(n6977), .C2(n4376), .A(n6053), .B(n6052), .ZN(n7469)
         );
  CLKBUF_X1 U5180 ( .A(n6126), .Z(n6385) );
  XNOR2_X1 U5181 ( .A(n10267), .B(n4530), .ZN(n10460) );
  NAND2_X1 U5182 ( .A1(n5379), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5393) );
  AND2_X1 U5183 ( .A1(n6411), .A2(n6410), .ZN(n6520) );
  NAND4_X2 U5184 ( .A1(n5142), .A2(n5141), .A3(n5140), .A4(n5139), .ZN(n9036)
         );
  NAND4_X2 U5185 ( .A1(n5168), .A2(n5169), .A3(n5167), .A4(n5170), .ZN(n7318)
         );
  NAND2_X1 U5186 ( .A1(n5482), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5230) );
  NAND2_X1 U5187 ( .A1(n5239), .A2(n5238), .ZN(n5253) );
  NAND2_X2 U5188 ( .A1(n6530), .A2(n6951), .ZN(n6974) );
  AND2_X1 U5189 ( .A1(n8861), .A2(n6030), .ZN(n6126) );
  NAND2_X2 U5190 ( .A1(n4397), .A2(n6964), .ZN(n6382) );
  NOR2_X1 U5191 ( .A1(n10462), .A2(n10266), .ZN(n10267) );
  OR2_X1 U5192 ( .A1(n4395), .A2(n8248), .ZN(n5141) );
  INV_X1 U5193 ( .A(n5380), .ZN(n5379) );
  XNOR2_X1 U5194 ( .A(n6529), .B(P1_IR_REG_26__SCAN_IN), .ZN(n6951) );
  NAND2_X1 U5195 ( .A1(n4608), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5380) );
  OR2_X1 U5196 ( .A1(n7543), .A2(n7757), .ZN(n7884) );
  CLKBUF_X2 U5197 ( .A(n5244), .Z(n4395) );
  OR2_X1 U5198 ( .A1(n4374), .A2(n7164), .ZN(n5177) );
  XNOR2_X1 U5199 ( .A(n6444), .B(n6443), .ZN(n7625) );
  OR2_X1 U5200 ( .A1(n5514), .A2(n6986), .ZN(n5186) );
  INV_X1 U5201 ( .A(n5353), .ZN(n4608) );
  NAND2_X1 U5202 ( .A1(n6528), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6529) );
  NAND2_X1 U5203 ( .A1(n10237), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5983) );
  NAND2_X1 U5204 ( .A1(n4609), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5353) );
  MUX2_X1 U5205 ( .A(n10359), .B(n9592), .S(n5207), .Z(n7595) );
  NAND2_X1 U5206 ( .A1(n4574), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5985) );
  AND2_X2 U5207 ( .A1(n8857), .A2(n5136), .ZN(n5225) );
  NAND2_X1 U5208 ( .A1(n6028), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6444) );
  INV_X1 U5209 ( .A(n8857), .ZN(n5138) );
  NAND2_X2 U5210 ( .A1(n5956), .A2(n8847), .ZN(n5207) );
  XNOR2_X1 U5211 ( .A(n5751), .B(n5750), .ZN(n7757) );
  NAND2_X1 U5212 ( .A1(n5980), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5975) );
  INV_X1 U5213 ( .A(n5136), .ZN(n8693) );
  INV_X1 U5214 ( .A(n5339), .ZN(n4609) );
  NAND2_X2 U5215 ( .A1(n6964), .A2(P1_U3084), .ZN(n10251) );
  AND2_X1 U5216 ( .A1(n5042), .A2(n4798), .ZN(n4797) );
  OAI21_X1 U5217 ( .B1(n5143), .B2(P2_IR_REG_27__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n4734) );
  XNOR2_X1 U5218 ( .A(n5254), .B(SI_5_), .ZN(n5251) );
  OR2_X1 U5219 ( .A1(n5134), .A2(n5133), .ZN(n5135) );
  CLKBUF_X1 U5220 ( .A(n5949), .Z(n4537) );
  NAND2_X1 U5221 ( .A1(n5090), .A2(n5159), .ZN(n7223) );
  AND2_X1 U5222 ( .A1(n5043), .A2(n5972), .ZN(n5042) );
  XNOR2_X1 U5223 ( .A(n5203), .B(n5209), .ZN(n7253) );
  XNOR2_X1 U5224 ( .A(n6051), .B(n6050), .ZN(n7007) );
  NAND2_X2 U5225 ( .A1(n4653), .A2(n5184), .ZN(n7204) );
  CLKBUF_X3 U5226 ( .A(n5470), .Z(n4398) );
  INV_X1 U5227 ( .A(n5283), .ZN(n5282) );
  CLKBUF_X3 U5228 ( .A(n5470), .Z(n4399) );
  AND2_X1 U5229 ( .A1(n4656), .A2(n4654), .ZN(n4653) );
  NAND2_X1 U5230 ( .A1(n5265), .A2(n5264), .ZN(n5283) );
  AND2_X1 U5231 ( .A1(n4900), .A2(n5533), .ZN(n4899) );
  INV_X1 U5232 ( .A(n4392), .ZN(n4391) );
  INV_X1 U5233 ( .A(n5965), .ZN(n5976) );
  NOR2_X1 U5234 ( .A1(n5973), .A2(P1_IR_REG_27__SCAN_IN), .ZN(n5043) );
  NAND3_X1 U5235 ( .A1(n4641), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n4640) );
  NAND3_X1 U5236 ( .A1(n4645), .A2(n4644), .A3(n4643), .ZN(n4642) );
  INV_X1 U5237 ( .A(n5263), .ZN(n5265) );
  AND2_X1 U5238 ( .A1(n5458), .A2(n5477), .ZN(n4900) );
  NAND4_X1 U5239 ( .A1(n4808), .A2(n5120), .A3(n5121), .A4(n5122), .ZN(n5298)
         );
  OR2_X1 U5240 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), .ZN(
        n5973) );
  INV_X1 U5241 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n6186) );
  AND2_X1 U5242 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_REG3_REG_6__SCAN_IN), 
        .ZN(n5264) );
  INV_X1 U5243 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n6168) );
  INV_X1 U5244 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n6164) );
  BUF_X2 U5245 ( .A(P2_IR_REG_0__SCAN_IN), .Z(n10367) );
  INV_X4 U5246 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  NOR2_X1 U5247 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n5968) );
  INV_X1 U5248 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n5995) );
  INV_X1 U5249 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5458) );
  NOR2_X1 U5250 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n5122) );
  NOR2_X2 U5251 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n4808) );
  NOR2_X1 U5252 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n5123) );
  INV_X1 U5253 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n5982) );
  NOR2_X1 U5254 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n5121) );
  NOR2_X1 U5255 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n5124) );
  INV_X4 U5256 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  NOR2_X1 U5257 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n5120) );
  INV_X1 U5258 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5477) );
  NOR2_X1 U5259 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n5125) );
  INV_X1 U5260 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4643) );
  INV_X1 U5261 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4645) );
  INV_X1 U5262 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4641) );
  INV_X1 U5263 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4644) );
  OAI21_X2 U5264 ( .B1(n9862), .B2(n4940), .A(n4939), .ZN(n10098) );
  XNOR2_X1 U5265 ( .A(n9855), .B(n9854), .ZN(n4382) );
  OAI21_X2 U5266 ( .B1(n9870), .B2(n4964), .A(n4961), .ZN(n9855) );
  INV_X1 U5267 ( .A(n6614), .ZN(n4386) );
  NOR2_X1 U5268 ( .A1(n6614), .A2(n6616), .ZN(n4387) );
  NAND2_X1 U5269 ( .A1(n9941), .A2(n4931), .ZN(n4927) );
  NAND2_X1 U5270 ( .A1(n4389), .A2(n6617), .ZN(n9941) );
  OAI22_X2 U5271 ( .A1(n6612), .A2(n6611), .B1(n10168), .B2(n10056), .ZN(
        n10028) );
  NOR2_X1 U5272 ( .A1(n7442), .A2(n6589), .ZN(n7767) );
  NAND2_X2 U5273 ( .A1(n4391), .A2(n5976), .ZN(n6139) );
  NAND4_X1 U5274 ( .A1(n6049), .A2(n5962), .A3(n5995), .A4(n6050), .ZN(n4392)
         );
  NOR2_X2 U5275 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n5963) );
  AND2_X2 U5276 ( .A1(n7349), .A2(n7348), .ZN(n7784) );
  OAI21_X2 U5277 ( .B1(n7860), .B2(n7861), .A(n4865), .ZN(n4867) );
  OR2_X1 U5278 ( .A1(n5744), .A2(n7217), .ZN(n5231) );
  OAI21_X1 U5279 ( .B1(n5848), .B2(n4817), .A(n4815), .ZN(n4819) );
  INV_X1 U5280 ( .A(n10245), .ZN(n6030) );
  INV_X2 U5281 ( .A(n7583), .ZN(n8787) );
  NAND2_X2 U5282 ( .A1(n9383), .A2(n9146), .ZN(n9358) );
  AOI21_X2 U5283 ( .B1(P2_REG1_REG_8__SCAN_IN), .B2(n7494), .A(n7490), .ZN(
        n7492) );
  AND3_X2 U5284 ( .A1(n6700), .A2(n10061), .A3(n5048), .ZN(n9998) );
  NAND2_X4 U5285 ( .A1(n4642), .A2(n4640), .ZN(n5470) );
  NAND2_X1 U5286 ( .A1(n5143), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4733) );
  OAI21_X2 U5287 ( .B1(n10027), .B2(n4921), .A(n4920), .ZN(n9968) );
  OAI21_X2 U5288 ( .B1(n8621), .B2(n4990), .A(n4988), .ZN(n9144) );
  NAND2_X2 U5289 ( .A1(n8556), .A2(n5932), .ZN(n8621) );
  AND2_X1 U5290 ( .A1(n8058), .A2(n10394), .ZN(n8060) );
  NOR2_X2 U5291 ( .A1(n9212), .A2(n9454), .ZN(n5066) );
  AND2_X2 U5292 ( .A1(n8039), .A2(n8043), .ZN(n7956) );
  OAI21_X2 U5293 ( .B1(n9241), .B2(n5679), .A(n5678), .ZN(n5680) );
  NAND2_X1 U5294 ( .A1(n9474), .A2(n9220), .ZN(n9236) );
  NOR2_X2 U5295 ( .A1(n4846), .A2(n4844), .ZN(n4843) );
  AND2_X1 U5296 ( .A1(n5776), .A2(n8862), .ZN(n5877) );
  NAND2_X1 U5297 ( .A1(n5188), .A2(n5189), .ZN(n5786) );
  INV_X2 U5298 ( .A(n5189), .ZN(n7316) );
  NAND3_X2 U5299 ( .A1(n5187), .A2(n5186), .A3(n5185), .ZN(n5189) );
  NAND2_X1 U5300 ( .A1(n6531), .A2(n7322), .ZN(n4396) );
  NAND2_X1 U5301 ( .A1(n6531), .A2(n7322), .ZN(n4397) );
  NAND2_X2 U5302 ( .A1(n6531), .A2(n7322), .ZN(n6977) );
  NAND2_X2 U5303 ( .A1(n5045), .A2(n4418), .ZN(n7837) );
  XNOR2_X2 U5304 ( .A(n5135), .B(P2_IR_REG_29__SCAN_IN), .ZN(n5136) );
  NOR2_X4 U5305 ( .A1(n5103), .A2(n10140), .ZN(n9931) );
  AND2_X4 U5306 ( .A1(n6713), .A2(n6974), .ZN(n6800) );
  NOR2_X4 U5307 ( .A1(n9850), .A2(n10087), .ZN(n9841) );
  OR2_X2 U5308 ( .A1(n9969), .A2(n10144), .ZN(n5103) );
  CLKBUF_X2 U5309 ( .A(n6696), .Z(n4401) );
  NOR2_X2 U5310 ( .A1(n7470), .A2(n7469), .ZN(n7454) );
  OAI211_X1 U5311 ( .C1(n7006), .C2(n6977), .A(n6038), .B(n6037), .ZN(n6696)
         );
  AND2_X1 U5312 ( .A1(n7139), .A2(n7138), .ZN(n9406) );
  INV_X1 U5313 ( .A(n9406), .ZN(n4402) );
  NAND2_X1 U5314 ( .A1(n4708), .A2(n4707), .ZN(n4706) );
  INV_X1 U5315 ( .A(n5446), .ZN(n4707) );
  AND2_X1 U5316 ( .A1(n4785), .A2(n4788), .ZN(n4784) );
  INV_X1 U5317 ( .A(n4789), .ZN(n4788) );
  NAND2_X1 U5318 ( .A1(n4786), .A2(n6243), .ZN(n4785) );
  OAI21_X1 U5319 ( .B1(n6467), .B2(n4791), .A(n4790), .ZN(n4789) );
  NAND2_X1 U5320 ( .A1(n10107), .A2(n9745), .ZN(n6412) );
  AND2_X1 U5321 ( .A1(n6869), .A2(n4469), .ZN(n5023) );
  NAND2_X1 U5322 ( .A1(n6370), .A2(n6369), .ZN(n10087) );
  NOR2_X1 U5323 ( .A1(n6618), .A2(n4936), .ZN(n4935) );
  INV_X1 U5324 ( .A(n5092), .ZN(n4936) );
  OR2_X1 U5325 ( .A1(n10102), .A2(n9596), .ZN(n6684) );
  NAND2_X1 U5326 ( .A1(n10102), .A2(n9596), .ZN(n6685) );
  INV_X1 U5327 ( .A(n4702), .ZN(n4701) );
  OAI21_X1 U5328 ( .B1(n4705), .B2(n4708), .A(n5016), .ZN(n4702) );
  AND2_X1 U5329 ( .A1(n5646), .A2(n5645), .ZN(n8954) );
  NAND2_X1 U5330 ( .A1(n5764), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5765) );
  INV_X1 U5331 ( .A(n9888), .ZN(n9655) );
  NAND2_X1 U5332 ( .A1(n5857), .A2(n5856), .ZN(n5858) );
  INV_X1 U5333 ( .A(n5855), .ZN(n5857) );
  AND2_X1 U5334 ( .A1(n4824), .A2(n4441), .ZN(n4509) );
  NOR2_X1 U5335 ( .A1(n4826), .A2(n4825), .ZN(n4824) );
  NAND2_X1 U5336 ( .A1(n5887), .A2(n5892), .ZN(n4825) );
  NOR2_X1 U5337 ( .A1(n9452), .A2(n9198), .ZN(n5897) );
  AND2_X1 U5338 ( .A1(n7965), .A2(n7986), .ZN(n5816) );
  OAI21_X1 U5339 ( .B1(n4784), .B2(n4969), .A(n9912), .ZN(n4783) );
  OAI21_X1 U5340 ( .B1(n4399), .B2(n4554), .A(n4553), .ZN(n5292) );
  NAND2_X1 U5341 ( .A1(n4399), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n4553) );
  NAND2_X1 U5342 ( .A1(n8815), .A2(n8816), .ZN(n4888) );
  NOR2_X1 U5343 ( .A1(n5638), .A2(n8958), .ZN(n4617) );
  AND2_X1 U5344 ( .A1(n7387), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n4915) );
  OR2_X1 U5345 ( .A1(n9475), .A2(n9281), .ZN(n5883) );
  OR2_X1 U5346 ( .A1(n5593), .A2(n8916), .ZN(n5919) );
  NAND2_X1 U5347 ( .A1(n4997), .A2(n9328), .ZN(n4996) );
  INV_X1 U5348 ( .A(n4998), .ZN(n4997) );
  OR2_X1 U5349 ( .A1(n9522), .A2(n9385), .ZN(n5845) );
  NOR2_X1 U5350 ( .A1(n5928), .A2(n4743), .ZN(n4742) );
  INV_X1 U5351 ( .A(n5805), .ZN(n4743) );
  NOR2_X2 U5352 ( .A1(n5454), .A2(n5453), .ZN(n5949) );
  OR2_X1 U5353 ( .A1(n5241), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n5278) );
  NAND2_X1 U5354 ( .A1(n6448), .A2(n5042), .ZN(n5980) );
  OAI21_X1 U5355 ( .B1(n6746), .B2(n4685), .A(n4682), .ZN(n6772) );
  INV_X1 U5356 ( .A(n4689), .ZN(n4683) );
  OR2_X1 U5357 ( .A1(n6862), .A2(n9641), .ZN(n6868) );
  OR2_X1 U5358 ( .A1(n6290), .A2(n4791), .ZN(n4764) );
  INV_X1 U5359 ( .A(n4767), .ZN(n4766) );
  NAND2_X1 U5360 ( .A1(n4544), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n6317) );
  AND2_X1 U5361 ( .A1(n10121), .A2(n9919), .ZN(n6620) );
  OR2_X1 U5362 ( .A1(n10140), .A2(n6857), .ZN(n6468) );
  NAND2_X1 U5363 ( .A1(n4924), .A2(n9990), .ZN(n4923) );
  NAND2_X1 U5364 ( .A1(n4373), .A2(n4925), .ZN(n4924) );
  INV_X1 U5365 ( .A(n4424), .ZN(n4925) );
  OR2_X1 U5366 ( .A1(n4569), .A2(n9841), .ZN(n10090) );
  INV_X1 U5367 ( .A(n4570), .ZN(n4569) );
  OR2_X1 U5368 ( .A1(n5658), .A2(n4485), .ZN(n4728) );
  INV_X1 U5369 ( .A(n5972), .ZN(n5041) );
  AND2_X1 U5370 ( .A1(n5018), .A2(n5504), .ZN(n5017) );
  OR2_X1 U5371 ( .A1(n5020), .A2(n4404), .ZN(n5018) );
  NAND2_X1 U5372 ( .A1(n4617), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n5669) );
  INV_X1 U5373 ( .A(n4617), .ZN(n5640) );
  NAND2_X1 U5374 ( .A1(n7142), .A2(n9361), .ZN(n7138) );
  INV_X1 U5375 ( .A(n4395), .ZN(n5698) );
  INV_X1 U5376 ( .A(n5285), .ZN(n5707) );
  XNOR2_X1 U5377 ( .A(n7204), .B(P2_REG1_REG_1__SCAN_IN), .ZN(n7197) );
  OR2_X1 U5378 ( .A1(n7220), .A2(n7219), .ZN(n4919) );
  NAND2_X1 U5379 ( .A1(n7260), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n4918) );
  INV_X1 U5380 ( .A(n7256), .ZN(n4916) );
  OR2_X1 U5381 ( .A1(n4916), .A2(n4915), .ZN(n4663) );
  NAND2_X1 U5382 ( .A1(n4919), .A2(n4664), .ZN(n4662) );
  NOR2_X1 U5383 ( .A1(n4915), .A2(n4665), .ZN(n4664) );
  INV_X1 U5384 ( .A(n4918), .ZN(n4665) );
  NAND2_X1 U5385 ( .A1(n8684), .A2(n8685), .ZN(n9058) );
  AND2_X1 U5386 ( .A1(n7142), .A2(n5955), .ZN(n7589) );
  AND2_X1 U5387 ( .A1(n5714), .A2(n4441), .ZN(n9179) );
  NAND2_X1 U5388 ( .A1(n9249), .A2(n5879), .ZN(n9241) );
  NAND2_X1 U5389 ( .A1(n8499), .A2(n4742), .ZN(n4741) );
  NAND2_X1 U5390 ( .A1(n5538), .A2(n7287), .ZN(n4756) );
  AND2_X1 U5391 ( .A1(n7589), .A2(n7140), .ZN(n9411) );
  OR2_X1 U5392 ( .A1(n7554), .A2(n7543), .ZN(n9518) );
  INV_X1 U5393 ( .A(n10403), .ZN(n10408) );
  OR2_X1 U5394 ( .A1(n7554), .A2(n7315), .ZN(n10403) );
  NAND2_X1 U5395 ( .A1(n7601), .A2(n7602), .ZN(n6746) );
  OAI22_X1 U5396 ( .A1(n4681), .A2(n4410), .B1(n4423), .B2(n4680), .ZN(n4679)
         );
  NOR2_X1 U5397 ( .A1(n6895), .A2(n4410), .ZN(n4680) );
  OR2_X1 U5398 ( .A1(n6317), .A2(n9651), .ZN(n6330) );
  AND2_X1 U5399 ( .A1(n6367), .A2(n6366), .ZN(n9596) );
  OR2_X1 U5400 ( .A1(n9847), .A2(n6371), .ZN(n6367) );
  INV_X1 U5401 ( .A(n6307), .ZN(n6371) );
  OAI21_X1 U5402 ( .B1(n7071), .B2(n4854), .A(n4461), .ZN(n4853) );
  INV_X1 U5403 ( .A(n4855), .ZN(n4854) );
  NAND2_X1 U5404 ( .A1(n7329), .A2(n4848), .ZN(n4852) );
  INV_X1 U5405 ( .A(n7071), .ZN(n4848) );
  AOI21_X1 U5406 ( .B1(n4843), .B2(n4840), .A(n5114), .ZN(n4839) );
  INV_X1 U5407 ( .A(n7026), .ZN(n4840) );
  OR2_X1 U5408 ( .A1(n9833), .A2(n9832), .ZN(n4836) );
  NAND2_X1 U5409 ( .A1(n4836), .A2(n4835), .ZN(n4834) );
  NAND2_X1 U5410 ( .A1(n9829), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n4835) );
  OR2_X1 U5411 ( .A1(n10293), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n4559) );
  AOI21_X1 U5412 ( .B1(n4722), .B2(n4724), .A(n4489), .ZN(n4721) );
  INV_X1 U5413 ( .A(n4725), .ZN(n4722) );
  INV_X1 U5414 ( .A(n4724), .ZN(n4723) );
  NAND2_X1 U5415 ( .A1(n5731), .A2(n5108), .ZN(n5734) );
  AOI21_X1 U5416 ( .B1(n4935), .B2(n4933), .A(n4463), .ZN(n4932) );
  CLKBUF_X1 U5417 ( .A(n6382), .Z(n4525) );
  OR2_X1 U5418 ( .A1(n10201), .A2(n9773), .ZN(n6598) );
  INV_X1 U5419 ( .A(n9952), .ZN(n10055) );
  INV_X1 U5420 ( .A(n9002), .ZN(n9014) );
  NAND2_X1 U5421 ( .A1(n5912), .A2(n5911), .ZN(n4827) );
  INV_X1 U5422 ( .A(n9596), .ZN(n9769) );
  NAND2_X1 U5423 ( .A1(n6337), .A2(n6336), .ZN(n9888) );
  NAND2_X1 U5424 ( .A1(n4527), .A2(n5911), .ZN(n4526) );
  NAND2_X1 U5425 ( .A1(n5799), .A2(n7350), .ZN(n4527) );
  OAI21_X1 U5426 ( .B1(n4777), .B2(n4791), .A(n4774), .ZN(n4772) );
  INV_X1 U5427 ( .A(n4779), .ZN(n4776) );
  AOI21_X1 U5428 ( .B1(n5858), .B2(n5921), .A(n4816), .ZN(n4815) );
  NAND2_X1 U5429 ( .A1(n5859), .A2(n5921), .ZN(n4817) );
  AOI21_X1 U5430 ( .B1(n5868), .B2(n5867), .A(n5866), .ZN(n5878) );
  INV_X1 U5431 ( .A(n6469), .ZN(n4792) );
  NAND2_X1 U5432 ( .A1(n4803), .A2(n4442), .ZN(n4802) );
  NAND2_X1 U5433 ( .A1(n6482), .A2(n4803), .ZN(n4799) );
  INV_X1 U5434 ( .A(n5033), .ZN(n5030) );
  INV_X1 U5435 ( .A(n6826), .ZN(n5008) );
  NAND2_X1 U5436 ( .A1(n4782), .A2(n4784), .ZN(n6286) );
  AND2_X1 U5437 ( .A1(n5650), .A2(n5653), .ZN(n5651) );
  INV_X1 U5438 ( .A(n5098), .ZN(n4709) );
  NAND2_X1 U5439 ( .A1(n5312), .A2(n5311), .ZN(n5329) );
  NAND2_X1 U5440 ( .A1(n5295), .A2(n5294), .ZN(n5307) );
  NOR2_X1 U5441 ( .A1(n7774), .A2(n4877), .ZN(n4876) );
  INV_X1 U5442 ( .A(n7669), .ZN(n4877) );
  INV_X1 U5443 ( .A(n8805), .ZN(n4889) );
  INV_X1 U5444 ( .A(n5088), .ZN(n5087) );
  AND2_X1 U5445 ( .A1(n5915), .A2(n5714), .ZN(n5088) );
  NOR2_X1 U5446 ( .A1(n5085), .A2(n9432), .ZN(n5084) );
  NOR4_X1 U5447 ( .A1(n9311), .A2(n9328), .A3(n9347), .A4(n5934), .ZN(n5935)
         );
  NOR2_X1 U5448 ( .A1(n9440), .A2(n5938), .ZN(n4523) );
  NAND2_X1 U5449 ( .A1(n5065), .A2(n4985), .ZN(n5064) );
  NOR2_X1 U5450 ( .A1(n9438), .A2(n9452), .ZN(n5065) );
  NAND2_X1 U5451 ( .A1(n4615), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5605) );
  AOI21_X1 U5452 ( .B1(n9328), .B2(n4652), .A(n4464), .ZN(n4651) );
  INV_X1 U5453 ( .A(n4999), .ZN(n4652) );
  INV_X1 U5454 ( .A(n4996), .ZN(n4994) );
  INV_X1 U5455 ( .A(n4744), .ZN(n4740) );
  NOR2_X1 U5456 ( .A1(n8506), .A2(n4809), .ZN(n5060) );
  NAND2_X1 U5457 ( .A1(n8825), .A2(n4985), .ZN(n4984) );
  NAND2_X1 U5458 ( .A1(n4982), .A2(n9154), .ZN(n4981) );
  INV_X1 U5459 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5130) );
  NAND2_X1 U5460 ( .A1(n5771), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5945) );
  NAND2_X1 U5461 ( .A1(n9716), .A2(n5025), .ZN(n5024) );
  NAND2_X1 U5462 ( .A1(n6877), .A2(n4696), .ZN(n4695) );
  INV_X1 U5463 ( .A(n5024), .ZN(n4696) );
  INV_X1 U5464 ( .A(n9619), .ZN(n4697) );
  OR2_X1 U5465 ( .A1(n6782), .A2(n8575), .ZN(n6786) );
  OR2_X1 U5466 ( .A1(n6747), .A2(n6748), .ZN(n4691) );
  INV_X1 U5467 ( .A(n6339), .ZN(n4760) );
  NAND2_X1 U5468 ( .A1(n6390), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n6040) );
  AND2_X1 U5469 ( .A1(n4866), .A2(n4493), .ZN(n4865) );
  OR2_X1 U5470 ( .A1(n7861), .A2(n7859), .ZN(n4866) );
  NAND2_X1 U5471 ( .A1(n6347), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n6360) );
  INV_X1 U5472 ( .A(n4942), .ZN(n4941) );
  NAND2_X1 U5473 ( .A1(n5054), .A2(n9868), .ZN(n5053) );
  NOR2_X1 U5474 ( .A1(n10116), .A2(n10121), .ZN(n5054) );
  INV_X1 U5475 ( .A(n4544), .ZN(n6306) );
  AND2_X1 U5476 ( .A1(n10131), .A2(n9918), .ZN(n6671) );
  NOR2_X1 U5477 ( .A1(n6454), .A2(n6668), .ZN(n4971) );
  NOR2_X1 U5478 ( .A1(n9947), .A2(n4969), .ZN(n4968) );
  NAND2_X1 U5479 ( .A1(n7446), .A2(n7702), .ZN(n6076) );
  OAI21_X1 U5480 ( .B1(n7463), .B2(n7369), .A(n7483), .ZN(n6572) );
  AOI21_X1 U5481 ( .B1(n7461), .B2(n7464), .A(n6054), .ZN(n7448) );
  XNOR2_X1 U5482 ( .A(n4401), .B(n9780), .ZN(n6422) );
  NAND2_X1 U5483 ( .A1(n5720), .A2(n5719), .ZN(n5729) );
  NOR2_X2 U5484 ( .A1(n5971), .A2(n6139), .ZN(n6448) );
  INV_X1 U5485 ( .A(n5475), .ZN(n5019) );
  AOI21_X1 U5486 ( .B1(n5290), .B2(n5013), .A(n4429), .ZN(n5012) );
  NAND2_X1 U5487 ( .A1(n4470), .A2(n4888), .ZN(n4883) );
  AND2_X1 U5488 ( .A1(n4407), .A2(n4440), .ZN(n4882) );
  INV_X1 U5489 ( .A(n4876), .ZN(n4875) );
  INV_X1 U5490 ( .A(n7662), .ZN(n4550) );
  NOR2_X1 U5491 ( .A1(n8814), .A2(n4887), .ZN(n4886) );
  INV_X1 U5492 ( .A(n8807), .ZN(n4887) );
  OR2_X1 U5493 ( .A1(n8844), .A2(n8849), .ZN(n5775) );
  AND4_X1 U5494 ( .A1(n5306), .A2(n5305), .A3(n5304), .A4(n5303), .ZN(n7936)
         );
  NAND2_X1 U5495 ( .A1(n7198), .A2(n7153), .ZN(n7157) );
  OAI21_X1 U5496 ( .B1(n7223), .B2(P2_REG1_REG_2__SCAN_IN), .A(n4904), .ZN(
        n7158) );
  NAND2_X1 U5497 ( .A1(n7223), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n4904) );
  AND2_X1 U5498 ( .A1(n4903), .A2(n4902), .ZN(n7244) );
  NAND2_X1 U5499 ( .A1(n7214), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n4902) );
  AND2_X1 U5500 ( .A1(n4662), .A2(n4483), .ZN(n7490) );
  INV_X1 U5501 ( .A(n7385), .ZN(n4661) );
  NAND2_X1 U5502 ( .A1(n4667), .A2(n4666), .ZN(n4914) );
  INV_X1 U5503 ( .A(n7728), .ZN(n4666) );
  AND2_X1 U5504 ( .A1(n4914), .A2(n4913), .ZN(n9040) );
  NAND2_X1 U5505 ( .A1(n8142), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n4913) );
  OR2_X1 U5506 ( .A1(n9040), .A2(n9039), .ZN(n4912) );
  NAND2_X1 U5507 ( .A1(n8648), .A2(n4901), .ZN(n8650) );
  OR2_X1 U5508 ( .A1(n8649), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n4901) );
  NOR2_X1 U5509 ( .A1(n9069), .A2(n9070), .ZN(n9072) );
  NAND2_X1 U5510 ( .A1(n9093), .A2(n8442), .ZN(n4905) );
  NAND2_X1 U5511 ( .A1(n9072), .A2(n9071), .ZN(n9086) );
  AND2_X1 U5512 ( .A1(n9086), .A2(n4658), .ZN(n9106) );
  AND2_X1 U5513 ( .A1(n4659), .A2(n4905), .ZN(n4658) );
  INV_X1 U5514 ( .A(n9088), .ZN(n4659) );
  NOR2_X1 U5515 ( .A1(n9106), .A2(n4660), .ZN(n9118) );
  OAI211_X1 U5516 ( .C1(n9118), .C2(n4909), .A(n4907), .B(n4906), .ZN(n9123)
         );
  AOI21_X1 U5517 ( .B1(n4908), .B2(n4910), .A(n4497), .ZN(n4907) );
  INV_X1 U5518 ( .A(n4910), .ZN(n4909) );
  OR2_X1 U5519 ( .A1(n9106), .A2(n4498), .ZN(n4906) );
  AND2_X1 U5520 ( .A1(n5713), .A2(n5712), .ZN(n9198) );
  OR2_X1 U5521 ( .A1(n9185), .A2(n4394), .ZN(n5713) );
  INV_X1 U5522 ( .A(n9025), .ZN(n9197) );
  NAND2_X1 U5523 ( .A1(n9461), .A2(n9197), .ZN(n5890) );
  AND2_X1 U5524 ( .A1(n5668), .A2(n5667), .ZN(n9152) );
  NOR2_X1 U5525 ( .A1(n9468), .A2(n9475), .ZN(n5058) );
  AND2_X1 U5526 ( .A1(n5630), .A2(n5629), .ZN(n9243) );
  OR2_X1 U5527 ( .A1(n9224), .A2(n4394), .ZN(n5630) );
  OR2_X1 U5528 ( .A1(n5593), .A2(n9299), .ZN(n4637) );
  AND2_X1 U5529 ( .A1(n4636), .A2(n4631), .ZN(n4630) );
  NAND2_X1 U5530 ( .A1(n4632), .A2(n4639), .ZN(n4631) );
  INV_X1 U5531 ( .A(n9149), .ZN(n4632) );
  NAND2_X1 U5532 ( .A1(n5568), .A2(n4427), .ZN(n4571) );
  NAND2_X1 U5533 ( .A1(n9148), .A2(n5001), .ZN(n4998) );
  NAND2_X1 U5534 ( .A1(n9499), .A2(n9333), .ZN(n4999) );
  NOR2_X1 U5535 ( .A1(n9358), .A2(n9357), .ZN(n9356) );
  AND4_X1 U5536 ( .A1(n5445), .A2(n5444), .A3(n5443), .A4(n5442), .ZN(n9385)
         );
  INV_X1 U5537 ( .A(n5839), .ZN(n4746) );
  NAND2_X1 U5538 ( .A1(n4611), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5440) );
  INV_X1 U5539 ( .A(n5412), .ZN(n4611) );
  NAND2_X1 U5540 ( .A1(n4510), .A2(n8557), .ZN(n8548) );
  NAND2_X1 U5541 ( .A1(n5076), .A2(n5077), .ZN(n5075) );
  INV_X1 U5542 ( .A(n8077), .ZN(n5076) );
  AND2_X1 U5543 ( .A1(n5075), .A2(n5827), .ZN(n8183) );
  AND2_X1 U5544 ( .A1(n7970), .A2(n5922), .ZN(n5078) );
  NAND2_X1 U5545 ( .A1(n4741), .A2(n4744), .ZN(n7989) );
  INV_X1 U5546 ( .A(n7782), .ZN(n4810) );
  INV_X1 U5547 ( .A(n9411), .ZN(n9384) );
  OR2_X1 U5548 ( .A1(n7568), .A2(n5188), .ZN(n7342) );
  INV_X1 U5549 ( .A(n9466), .ZN(n4628) );
  INV_X1 U5550 ( .A(n9465), .ZN(n4627) );
  AND3_X1 U5551 ( .A1(n7134), .A2(n7541), .A3(n7133), .ZN(n7362) );
  AND2_X1 U5552 ( .A1(n7121), .A2(n8193), .ZN(n10371) );
  AND2_X1 U5553 ( .A1(n4899), .A2(n5749), .ZN(n4898) );
  XNOR2_X1 U5554 ( .A(n5257), .B(P2_IR_REG_6__SCAN_IN), .ZN(n7260) );
  AND2_X1 U5555 ( .A1(n5242), .A2(n5278), .ZN(n7287) );
  INV_X1 U5556 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5157) );
  NAND2_X1 U5557 ( .A1(n4808), .A2(n5157), .ZN(n5208) );
  INV_X1 U5558 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n4655) );
  AND2_X1 U5559 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n4657) );
  OAI21_X1 U5560 ( .B1(n6521), .B2(n5973), .A(n4467), .ZN(n4950) );
  NOR2_X1 U5561 ( .A1(n4949), .A2(n4948), .ZN(n4947) );
  XNOR2_X1 U5562 ( .A(n6856), .B(n6806), .ZN(n6861) );
  NAND2_X1 U5563 ( .A1(n5987), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n6108) );
  INV_X1 U5564 ( .A(n6106), .ZN(n5987) );
  NAND2_X1 U5565 ( .A1(n6158), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n6173) );
  INV_X1 U5566 ( .A(n6171), .ZN(n6158) );
  NAND2_X1 U5567 ( .A1(n6868), .A2(n4426), .ZN(n6869) );
  OR2_X1 U5568 ( .A1(n6330), .A2(n9742), .ZN(n6349) );
  AND2_X1 U5569 ( .A1(n6377), .A2(n6376), .ZN(n9768) );
  AND2_X1 U5570 ( .A1(n6271), .A2(n6270), .ZN(n6857) );
  NAND2_X1 U5571 ( .A1(n7065), .A2(n7066), .ZN(n7064) );
  NAND2_X1 U5572 ( .A1(n4852), .A2(n4850), .ZN(n9790) );
  NOR2_X1 U5573 ( .A1(n4853), .A2(n4851), .ZN(n4850) );
  NOR2_X1 U5574 ( .A1(n7430), .A2(n4863), .ZN(n4862) );
  INV_X1 U5575 ( .A(n7410), .ZN(n4863) );
  NAND2_X1 U5576 ( .A1(n7412), .A2(n4864), .ZN(n4861) );
  OAI21_X1 U5577 ( .B1(n7411), .B2(n4860), .A(n4857), .ZN(n7718) );
  INV_X1 U5578 ( .A(n4861), .ZN(n4860) );
  AOI21_X1 U5579 ( .B1(n4859), .B2(n4861), .A(n4858), .ZN(n4857) );
  INV_X1 U5580 ( .A(n4862), .ZN(n4859) );
  OR2_X1 U5581 ( .A1(n7179), .A2(n7180), .ZN(n7411) );
  OR2_X1 U5582 ( .A1(n7721), .A2(n7722), .ZN(n7860) );
  XNOR2_X1 U5583 ( .A(n4867), .B(n8709), .ZN(n8635) );
  NOR2_X1 U5584 ( .A1(n8634), .A2(n8635), .ZN(n8697) );
  INV_X1 U5585 ( .A(n10290), .ZN(n4833) );
  NAND2_X1 U5586 ( .A1(n6384), .A2(n6383), .ZN(n6437) );
  AND2_X1 U5587 ( .A1(n6512), .A2(n6555), .ZN(n10097) );
  INV_X1 U5588 ( .A(n4965), .ZN(n4964) );
  AOI21_X1 U5589 ( .B1(n4965), .B2(n4963), .A(n4962), .ZN(n4961) );
  NOR2_X1 U5590 ( .A1(n8838), .A2(n6509), .ZN(n4965) );
  NAND2_X1 U5591 ( .A1(n6684), .A2(n6685), .ZN(n9854) );
  NAND2_X1 U5592 ( .A1(n9873), .A2(n10057), .ZN(n9857) );
  NAND2_X1 U5593 ( .A1(n9873), .A2(n10055), .ZN(n9875) );
  OR2_X1 U5594 ( .A1(n6413), .A2(n6620), .ZN(n9899) );
  AOI21_X1 U5595 ( .B1(n4930), .B2(n4932), .A(n4929), .ZN(n4928) );
  NOR2_X1 U5596 ( .A1(n9910), .A2(n9720), .ZN(n4929) );
  INV_X1 U5597 ( .A(n4935), .ZN(n4934) );
  AND2_X1 U5598 ( .A1(n6282), .A2(n6281), .ZN(n9951) );
  AND2_X1 U5599 ( .A1(n6415), .A2(n6666), .ZN(n9977) );
  NAND2_X1 U5600 ( .A1(n4424), .A2(n6613), .ZN(n4926) );
  OAI21_X1 U5601 ( .B1(n7515), .B2(n6597), .A(n6596), .ZN(n7893) );
  OAI21_X1 U5602 ( .B1(n7832), .B2(n4975), .A(n6646), .ZN(n4974) );
  NAND2_X1 U5603 ( .A1(n6076), .A2(n7698), .ZN(n7704) );
  OR2_X1 U5604 ( .A1(n7185), .A2(n7367), .ZN(n10334) );
  OAI211_X1 U5605 ( .C1(n5734), .C2(n4723), .A(n4721), .B(n4717), .ZN(n9583)
         );
  NAND2_X1 U5606 ( .A1(n5665), .A2(n5664), .ZN(n5682) );
  NAND2_X1 U5607 ( .A1(n5632), .A2(n5631), .ZN(n5634) );
  XNOR2_X1 U5608 ( .A(n5576), .B(n5571), .ZN(n6261) );
  AND4_X1 U5609 ( .A1(n5327), .A2(n5326), .A3(n5325), .A4(n5324), .ZN(n7986)
         );
  AND4_X1 U5610 ( .A1(n5358), .A2(n5357), .A3(n5356), .A4(n5355), .ZN(n8657)
         );
  OAI21_X1 U5611 ( .B1(n4512), .B2(n4431), .A(n4511), .ZN(n8811) );
  NAND2_X1 U5612 ( .A1(n4512), .A2(n8810), .ZN(n4511) );
  NAND2_X1 U5613 ( .A1(n8809), .A2(n4513), .ZN(n4512) );
  AND2_X1 U5614 ( .A1(n5640), .A2(n5639), .ZN(n9238) );
  NAND2_X1 U5615 ( .A1(n9468), .A2(n9019), .ZN(n4534) );
  INV_X1 U5616 ( .A(n7554), .ZN(n4895) );
  AND2_X1 U5617 ( .A1(n5612), .A2(n5611), .ZN(n9281) );
  OR2_X1 U5618 ( .A1(n8999), .A2(n9386), .ZN(n9017) );
  NAND2_X1 U5619 ( .A1(n7552), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9002) );
  NAND2_X1 U5620 ( .A1(n5942), .A2(n4508), .ZN(n4507) );
  INV_X1 U5621 ( .A(n9147), .ZN(n9333) );
  AND3_X1 U5622 ( .A1(n5498), .A2(n5497), .A3(n5496), .ZN(n9387) );
  OAI211_X1 U5623 ( .C1(n7204), .C2(n7164), .A(n7165), .B(n4610), .ZN(n7207)
         );
  NAND2_X1 U5624 ( .A1(n7204), .A2(n7164), .ZN(n4610) );
  NAND2_X1 U5625 ( .A1(n7226), .A2(n7225), .ZN(n7277) );
  NAND2_X1 U5626 ( .A1(n8141), .A2(n8140), .ZN(n8648) );
  OR2_X1 U5627 ( .A1(n9126), .A2(n4604), .ZN(n4603) );
  NAND2_X1 U5628 ( .A1(n4606), .A2(n4605), .ZN(n4604) );
  NOR2_X1 U5629 ( .A1(n10362), .A2(n7537), .ZN(n4605) );
  INV_X1 U5630 ( .A(n9152), .ZN(n9461) );
  NAND2_X1 U5631 ( .A1(n5039), .A2(n9211), .ZN(n9459) );
  OAI21_X1 U5632 ( .B1(n5916), .B2(n4454), .A(n4624), .ZN(n4623) );
  NAND2_X1 U5633 ( .A1(n5916), .A2(n4625), .ZN(n4624) );
  INV_X1 U5634 ( .A(n9221), .ZN(n4625) );
  NOR2_X1 U5635 ( .A1(n5916), .A2(n9221), .ZN(n4622) );
  NAND2_X1 U5636 ( .A1(n4619), .A2(n4449), .ZN(n4621) );
  INV_X1 U5637 ( .A(n9236), .ZN(n4619) );
  NAND2_X1 U5638 ( .A1(n10373), .A2(n7556), .ZN(n9373) );
  INV_X1 U5639 ( .A(n9404), .ZN(n9427) );
  INV_X1 U5640 ( .A(n9450), .ZN(n4753) );
  AND2_X1 U5641 ( .A1(n9452), .A2(n10408), .ZN(n4752) );
  NOR2_X1 U5642 ( .A1(n4411), .A2(n9765), .ZN(n4676) );
  NAND2_X1 U5643 ( .A1(n4679), .A2(n4455), .ZN(n4678) );
  NAND2_X1 U5644 ( .A1(n6346), .A2(n6345), .ZN(n10107) );
  OAI22_X1 U5645 ( .A1(n7482), .A2(n7481), .B1(n6745), .B2(n6744), .ZN(n7601)
         );
  INV_X1 U5646 ( .A(n9926), .ZN(n9720) );
  AND2_X1 U5647 ( .A1(n6324), .A2(n6323), .ZN(n9744) );
  INV_X1 U5648 ( .A(n9744), .ZN(n9900) );
  NAND2_X1 U5649 ( .A1(n6301), .A2(n6300), .ZN(n9919) );
  OR2_X1 U5650 ( .A1(n9686), .A2(n6371), .ZN(n6301) );
  INV_X1 U5651 ( .A(n6857), .ZN(n9959) );
  NOR2_X1 U5652 ( .A1(n7331), .A2(n7330), .ZN(n7329) );
  OR2_X1 U5653 ( .A1(n7080), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n7076) );
  NOR2_X1 U5654 ( .A1(n7429), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n4519) );
  NAND2_X1 U5655 ( .A1(n8717), .A2(n10302), .ZN(n4562) );
  INV_X1 U5656 ( .A(n4561), .ZN(n4560) );
  OAI21_X1 U5657 ( .B1(n8719), .B2(n8720), .A(n9632), .ZN(n4868) );
  INV_X1 U5658 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n8720) );
  NAND2_X1 U5659 ( .A1(n6380), .A2(n6379), .ZN(n10079) );
  NAND2_X1 U5660 ( .A1(n4721), .A2(n4723), .ZN(n4718) );
  INV_X1 U5661 ( .A(n10097), .ZN(n10088) );
  NAND2_X1 U5662 ( .A1(n6708), .A2(n6707), .ZN(n6709) );
  NAND2_X1 U5663 ( .A1(n6358), .A2(n6357), .ZN(n10102) );
  NAND2_X1 U5664 ( .A1(n10247), .A2(n6381), .ZN(n6358) );
  XNOR2_X1 U5665 ( .A(n8832), .B(n6436), .ZN(n10110) );
  INV_X1 U5666 ( .A(n8840), .ZN(n8841) );
  AOI21_X1 U5667 ( .B1(n9769), .B2(n10055), .A(n8839), .ZN(n8840) );
  INV_X1 U5668 ( .A(n5824), .ZN(n4590) );
  AND2_X1 U5669 ( .A1(n5816), .A2(n5877), .ZN(n4591) );
  INV_X1 U5670 ( .A(n4773), .ZN(n6119) );
  INV_X1 U5671 ( .A(n4772), .ZN(n4771) );
  NOR2_X1 U5672 ( .A1(n5885), .A2(n4585), .ZN(n4584) );
  NAND2_X1 U5673 ( .A1(n5880), .A2(n5917), .ZN(n4585) );
  NAND2_X1 U5674 ( .A1(n4793), .A2(n4791), .ZN(n4790) );
  NAND2_X1 U5675 ( .A1(n6666), .A2(n6416), .ZN(n4793) );
  NAND2_X1 U5676 ( .A1(n4415), .A2(n4787), .ZN(n4786) );
  NAND2_X1 U5677 ( .A1(n4792), .A2(n7368), .ZN(n4787) );
  OR2_X1 U5678 ( .A1(n5901), .A2(n5902), .ZN(n4592) );
  NAND2_X1 U5679 ( .A1(n7316), .A2(n7141), .ZN(n5925) );
  NAND2_X1 U5680 ( .A1(n5069), .A2(n5925), .ZN(n5784) );
  NAND2_X1 U5681 ( .A1(n7594), .A2(n5786), .ZN(n5069) );
  INV_X1 U5682 ( .A(n7747), .ZN(n4686) );
  NAND2_X1 U5683 ( .A1(n4800), .A2(n4443), .ZN(n6228) );
  AND2_X1 U5684 ( .A1(n9868), .A2(n9888), .ZN(n6340) );
  INV_X1 U5685 ( .A(n6671), .ZN(n6669) );
  NOR2_X1 U5686 ( .A1(n6304), .A2(n8331), .ZN(n4544) );
  NAND2_X1 U5687 ( .A1(n6491), .A2(n6497), .ZN(n4953) );
  AOI21_X1 U5688 ( .B1(n4713), .B2(n5688), .A(n4712), .ZN(n4711) );
  INV_X1 U5689 ( .A(n5715), .ZN(n4712) );
  INV_X1 U5690 ( .A(n5594), .ZN(n4729) );
  AND2_X1 U5691 ( .A1(n6526), .A2(n6447), .ZN(n5972) );
  AOI21_X1 U5692 ( .B1(n5017), .B2(n4404), .A(n5511), .ZN(n5016) );
  NOR2_X1 U5693 ( .A1(n5476), .A2(n5021), .ZN(n5020) );
  INV_X1 U5694 ( .A(n5468), .ZN(n5021) );
  AOI21_X1 U5695 ( .B1(n5422), .B2(n5421), .A(n5420), .ZN(n5424) );
  INV_X1 U5696 ( .A(n5421), .ZN(n5425) );
  NAND2_X1 U5697 ( .A1(n5386), .A2(SI_13_), .ZN(n5421) );
  INV_X1 U5698 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n5310) );
  INV_X1 U5699 ( .A(SI_7_), .ZN(n4699) );
  OAI21_X1 U5700 ( .B1(n4398), .B2(n4539), .A(n4538), .ZN(n5276) );
  NAND2_X1 U5701 ( .A1(n4398), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n4538) );
  OAI21_X1 U5702 ( .B1(n5470), .B2(P1_DATAO_REG_3__SCAN_IN), .A(n4576), .ZN(
        n5218) );
  NAND2_X1 U5703 ( .A1(n5470), .A2(n6944), .ZN(n4576) );
  OAI211_X1 U5704 ( .C1(n5470), .C2(n6987), .A(n5196), .B(n5195), .ZN(n5198)
         );
  NAND2_X1 U5705 ( .A1(n5517), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5544) );
  INV_X1 U5706 ( .A(n5542), .ZN(n5517) );
  AND2_X1 U5707 ( .A1(n9121), .A2(n9122), .ZN(n4910) );
  INV_X1 U5708 ( .A(n9119), .ZN(n4908) );
  NAND2_X1 U5709 ( .A1(n5030), .A2(n9206), .ZN(n5029) );
  AND2_X1 U5710 ( .A1(n9206), .A2(n9254), .ZN(n5032) );
  OR2_X1 U5711 ( .A1(n9464), .A2(n9243), .ZN(n9207) );
  INV_X1 U5712 ( .A(n9139), .ZN(n4990) );
  NOR2_X1 U5713 ( .A1(n5462), .A2(n8304), .ZN(n4616) );
  NAND2_X1 U5714 ( .A1(n5073), .A2(n5834), .ZN(n5072) );
  INV_X1 U5715 ( .A(n5074), .ZN(n5073) );
  INV_X1 U5716 ( .A(n7988), .ZN(n7791) );
  OR2_X1 U5717 ( .A1(n10407), .A2(n7987), .ZN(n4744) );
  OR2_X1 U5718 ( .A1(n5375), .A2(P2_IR_REG_11__SCAN_IN), .ZN(n5388) );
  OR2_X1 U5719 ( .A1(n5454), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n5335) );
  INV_X1 U5720 ( .A(n5980), .ZN(n4949) );
  NOR2_X1 U5721 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .ZN(
        n4948) );
  AND2_X1 U5722 ( .A1(n8219), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n6077) );
  INV_X1 U5723 ( .A(n6974), .ZN(n6725) );
  NOR2_X1 U5724 ( .A1(n9626), .A2(n9727), .ZN(n5010) );
  NAND2_X1 U5725 ( .A1(n5011), .A2(n5007), .ZN(n5004) );
  NOR2_X1 U5726 ( .A1(n9674), .A2(n6838), .ZN(n5011) );
  NAND2_X1 U5727 ( .A1(n5008), .A2(n5009), .ZN(n5007) );
  NOR2_X1 U5728 ( .A1(n6220), .A2(n6219), .ZN(n4599) );
  INV_X1 U5729 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n6408) );
  INV_X1 U5730 ( .A(n7432), .ZN(n4858) );
  NOR2_X1 U5731 ( .A1(n5755), .A2(n4726), .ZN(n4725) );
  INV_X1 U5732 ( .A(n5733), .ZN(n4726) );
  NOR2_X1 U5733 ( .A1(n5758), .A2(n4488), .ZN(n4724) );
  OR2_X1 U5734 ( .A1(n10087), .A2(n9768), .ZN(n6512) );
  INV_X1 U5735 ( .A(n6681), .ZN(n4963) );
  OR2_X1 U5736 ( .A1(n10121), .A2(n9919), .ZN(n6619) );
  AND2_X1 U5737 ( .A1(n4932), .A2(n4439), .ZN(n4931) );
  AND2_X1 U5738 ( .A1(n4439), .A2(n4934), .ZN(n4930) );
  NAND2_X1 U5739 ( .A1(n4600), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n6304) );
  NOR2_X1 U5740 ( .A1(n6264), .A2(n9642), .ZN(n4600) );
  NAND2_X1 U5741 ( .A1(n4956), .A2(n4955), .ZN(n4954) );
  INV_X1 U5742 ( .A(n4958), .ZN(n4955) );
  NAND2_X1 U5743 ( .A1(n6418), .A2(n6654), .ZN(n6653) );
  NAND2_X1 U5744 ( .A1(n4778), .A2(n6587), .ZN(n4777) );
  INV_X1 U5745 ( .A(n4780), .ZN(n4778) );
  AOI21_X1 U5746 ( .B1(n4781), .B2(n6496), .A(n6491), .ZN(n4780) );
  NAND2_X1 U5747 ( .A1(n6496), .A2(n6587), .ZN(n4779) );
  AND2_X1 U5748 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n8219) );
  INV_X1 U5749 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n6447) );
  NOR2_X1 U5750 ( .A1(n5595), .A2(n4731), .ZN(n4730) );
  INV_X1 U5751 ( .A(n5574), .ZN(n4731) );
  AOI21_X1 U5752 ( .B1(n4648), .B2(n4650), .A(n5525), .ZN(n4647) );
  INV_X1 U5753 ( .A(n4649), .ZN(n4648) );
  OAI21_X1 U5754 ( .B1(n4708), .B2(n4650), .A(n5475), .ZN(n4649) );
  INV_X1 U5755 ( .A(n5020), .ZN(n4650) );
  NAND2_X1 U5756 ( .A1(n5432), .A2(n5431), .ZN(n5446) );
  XNOR2_X1 U5757 ( .A(n5427), .B(SI_14_), .ZN(n5423) );
  AND2_X1 U5758 ( .A1(n5368), .A2(n5370), .ZN(n5369) );
  XNOR2_X1 U5759 ( .A(n5366), .B(SI_11_), .ZN(n5361) );
  NAND2_X1 U5760 ( .A1(n5307), .A2(n5297), .ZN(n5308) );
  XNOR2_X1 U5761 ( .A(n5276), .B(SI_6_), .ZN(n5273) );
  INV_X1 U5762 ( .A(n5251), .ZN(n5252) );
  INV_X4 U5763 ( .A(n8787), .ZN(n8820) );
  INV_X1 U5764 ( .A(n4615), .ZN(n5585) );
  OR2_X1 U5765 ( .A1(n7782), .A2(n8819), .ZN(n7613) );
  NAND2_X1 U5766 ( .A1(n4515), .A2(n4514), .ZN(n4892) );
  INV_X1 U5767 ( .A(n7653), .ZN(n4514) );
  INV_X1 U5768 ( .A(n7912), .ZN(n4871) );
  CLKBUF_X1 U5769 ( .A(n7643), .Z(n4552) );
  NAND2_X1 U5770 ( .A1(n4552), .A2(n7644), .ZN(n7670) );
  NAND2_X1 U5771 ( .A1(n5938), .A2(n5911), .ZN(n4829) );
  INV_X1 U5772 ( .A(n5081), .ZN(n5080) );
  OAI22_X1 U5773 ( .A1(n4414), .A2(n4494), .B1(n5088), .B2(n5082), .ZN(n5081)
         );
  INV_X1 U5774 ( .A(n5084), .ZN(n5082) );
  NOR2_X1 U5775 ( .A1(n4412), .A2(n5084), .ZN(n5083) );
  AND2_X1 U5776 ( .A1(n5937), .A2(n4413), .ZN(n5939) );
  AND3_X1 U5777 ( .A1(n5485), .A2(n5484), .A3(n5483), .ZN(n9147) );
  AND3_X1 U5778 ( .A1(n5466), .A2(n5465), .A3(n5464), .ZN(n9027) );
  AND4_X1 U5779 ( .A1(n5344), .A2(n5343), .A3(n5342), .A4(n5341), .ZN(n8159)
         );
  NOR2_X1 U5780 ( .A1(n7244), .A2(n7243), .ZN(n7242) );
  OR2_X1 U5781 ( .A1(n7727), .A2(n4668), .ZN(n4667) );
  AND2_X1 U5782 ( .A1(n7731), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n4668) );
  NAND2_X1 U5783 ( .A1(n7496), .A2(n7495), .ZN(n7737) );
  NAND2_X1 U5784 ( .A1(n8650), .A2(n8651), .ZN(n8683) );
  NAND2_X1 U5785 ( .A1(n9127), .A2(n10366), .ZN(n4606) );
  NAND2_X1 U5786 ( .A1(n4549), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5536) );
  NAND2_X1 U5787 ( .A1(n5949), .A2(n4899), .ZN(n4549) );
  AND2_X1 U5788 ( .A1(n5703), .A2(n5670), .ZN(n9000) );
  NAND2_X1 U5789 ( .A1(n9266), .A2(n9261), .ZN(n9256) );
  INV_X1 U5790 ( .A(n4993), .ZN(n4992) );
  OAI21_X1 U5791 ( .B1(n4996), .B2(n9364), .A(n4651), .ZN(n4993) );
  NAND2_X1 U5792 ( .A1(n4616), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n5495) );
  AND2_X1 U5793 ( .A1(n9391), .A2(n9326), .ZN(n9362) );
  INV_X1 U5794 ( .A(n4616), .ZN(n5493) );
  NOR2_X1 U5795 ( .A1(n9416), .A2(n9522), .ZN(n9417) );
  AND4_X1 U5796 ( .A1(n5385), .A2(n5384), .A3(n5383), .A4(n5382), .ZN(n8661)
         );
  AND4_X1 U5797 ( .A1(n5417), .A2(n5416), .A3(n5415), .A4(n5414), .ZN(n9012)
         );
  AND2_X1 U5798 ( .A1(n4409), .A2(n7980), .ZN(n8564) );
  AND2_X1 U5799 ( .A1(n7968), .A2(n7966), .ZN(n4583) );
  NAND2_X1 U5800 ( .A1(n5079), .A2(n5922), .ZN(n7974) );
  NAND2_X1 U5801 ( .A1(n7980), .A2(n8131), .ZN(n8188) );
  INV_X1 U5802 ( .A(n4736), .ZN(n4735) );
  AND2_X1 U5803 ( .A1(n5923), .A2(n5922), .ZN(n7797) );
  NOR2_X2 U5804 ( .A1(n7997), .A2(n9552), .ZN(n7996) );
  AND2_X1 U5805 ( .A1(n8509), .A2(n8507), .ZN(n7783) );
  AND2_X1 U5806 ( .A1(n8060), .A2(n7781), .ZN(n8504) );
  OR3_X1 U5807 ( .A1(n7870), .A2(n7869), .A3(n7868), .ZN(n7871) );
  CLKBUF_X1 U5808 ( .A(n7314), .Z(n7317) );
  NAND2_X1 U5809 ( .A1(n4982), .A2(n4979), .ZN(n4978) );
  NAND2_X1 U5810 ( .A1(n6261), .A2(n5635), .ZN(n5036) );
  INV_X1 U5811 ( .A(n9518), .ZN(n10409) );
  AOI22_X1 U5812 ( .A1(n4810), .A2(n9412), .B1(n7346), .B2(n9411), .ZN(n8068)
         );
  XNOR2_X1 U5813 ( .A(n5947), .B(P2_IR_REG_24__SCAN_IN), .ZN(n7135) );
  AND2_X1 U5814 ( .A1(n4537), .A2(n5458), .ZN(n5488) );
  AND2_X1 U5815 ( .A1(n5435), .A2(n5408), .ZN(n9059) );
  AND2_X1 U5816 ( .A1(n5210), .A2(n5209), .ZN(n5214) );
  INV_X1 U5817 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5209) );
  INV_X1 U5818 ( .A(n4691), .ZN(n4690) );
  NAND2_X1 U5819 ( .A1(n6077), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n6106) );
  INV_X1 U5820 ( .A(n4423), .ZN(n4681) );
  NOR2_X1 U5821 ( .A1(n6772), .A2(n6771), .ZN(n8107) );
  NAND2_X1 U5822 ( .A1(n6206), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n6220) );
  INV_X1 U5823 ( .A(n6208), .ZN(n6206) );
  NAND2_X1 U5824 ( .A1(n5022), .A2(n4428), .ZN(n9617) );
  NAND2_X1 U5825 ( .A1(n4692), .A2(n6877), .ZN(n9616) );
  NAND2_X1 U5826 ( .A1(n5022), .A2(n5024), .ZN(n4692) );
  NOR2_X1 U5827 ( .A1(n9685), .A2(n4694), .ZN(n4693) );
  NAND2_X1 U5828 ( .A1(n4543), .A2(n4453), .ZN(n6003) );
  INV_X1 U5829 ( .A(n6108), .ZN(n4543) );
  AND2_X1 U5830 ( .A1(n6816), .A2(n6815), .ZN(n9699) );
  NAND2_X1 U5831 ( .A1(n6128), .A2(n6127), .ZN(n6171) );
  INV_X1 U5832 ( .A(n6143), .ZN(n6128) );
  INV_X1 U5833 ( .A(n6918), .ZN(n6874) );
  OR2_X1 U5834 ( .A1(n6791), .A2(n6790), .ZN(n8537) );
  NAND2_X1 U5835 ( .A1(n4542), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n6143) );
  INV_X1 U5836 ( .A(n6003), .ZN(n4542) );
  NAND2_X1 U5837 ( .A1(n4599), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n6249) );
  INV_X1 U5838 ( .A(n4599), .ZN(n6238) );
  NAND2_X1 U5839 ( .A1(n6746), .A2(n4691), .ZN(n8200) );
  INV_X1 U5840 ( .A(n9743), .ZN(n9755) );
  NAND2_X1 U5841 ( .A1(n4598), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n6194) );
  INV_X1 U5842 ( .A(n6173), .ZN(n4598) );
  NAND2_X1 U5843 ( .A1(n4597), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n6208) );
  INV_X1 U5844 ( .A(n6194), .ZN(n4597) );
  NOR2_X1 U5845 ( .A1(n6398), .A2(n4962), .ZN(n6368) );
  OAI21_X1 U5846 ( .B1(n4766), .B2(n4769), .A(n4761), .ZN(n5101) );
  NOR2_X1 U5847 ( .A1(n6356), .A2(n4763), .ZN(n4762) );
  NAND2_X1 U5848 ( .A1(n4768), .A2(n6339), .ZN(n4763) );
  AND2_X1 U5849 ( .A1(n6355), .A2(n6354), .ZN(n9745) );
  OR2_X1 U5850 ( .A1(n8835), .A2(n6371), .ZN(n6355) );
  NAND4_X1 U5851 ( .A1(n6042), .A2(n6041), .A3(n6040), .A4(n6039), .ZN(n6729)
         );
  NAND2_X1 U5852 ( .A1(n6266), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6041) );
  AND2_X1 U5853 ( .A1(n7332), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n4855) );
  NAND2_X1 U5854 ( .A1(n7064), .A2(n4451), .ZN(n9784) );
  NOR2_X1 U5855 ( .A1(n8697), .A2(n8698), .ZN(n8699) );
  AOI21_X1 U5856 ( .B1(n8713), .B2(P1_REG1_REG_16__SCAN_IN), .A(n9812), .ZN(
        n9826) );
  OAI21_X1 U5857 ( .B1(n8716), .B2(n8715), .A(n9818), .ZN(n4561) );
  INV_X1 U5858 ( .A(n10090), .ZN(n10089) );
  NAND2_X1 U5859 ( .A1(n4945), .A2(n4403), .ZN(n4942) );
  AND2_X1 U5860 ( .A1(n8838), .A2(n4946), .ZN(n4943) );
  NOR2_X1 U5861 ( .A1(n9954), .A2(n9655), .ZN(n8839) );
  AND2_X1 U5862 ( .A1(n5051), .A2(n8837), .ZN(n5050) );
  INV_X1 U5863 ( .A(n5053), .ZN(n5051) );
  INV_X1 U5864 ( .A(n5054), .ZN(n5052) );
  INV_X1 U5865 ( .A(n4600), .ZN(n6275) );
  NAND2_X1 U5866 ( .A1(n4541), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n6256) );
  INV_X1 U5867 ( .A(n6249), .ZN(n4541) );
  NAND2_X1 U5868 ( .A1(n4540), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n6264) );
  INV_X1 U5869 ( .A(n6256), .ZN(n4540) );
  NOR2_X1 U5870 ( .A1(n10154), .A2(n10174), .ZN(n5048) );
  NAND2_X1 U5871 ( .A1(n9998), .A2(n9975), .ZN(n9969) );
  NAND2_X1 U5872 ( .A1(n4373), .A2(n4405), .ZN(n4921) );
  NAND2_X1 U5873 ( .A1(n4923), .A2(n4405), .ZN(n4920) );
  NAND2_X1 U5874 ( .A1(n10062), .A2(n6700), .ZN(n10007) );
  NAND2_X1 U5875 ( .A1(n4957), .A2(n6661), .ZN(n10003) );
  NAND2_X1 U5876 ( .A1(n6660), .A2(n4958), .ZN(n4957) );
  AND2_X1 U5877 ( .A1(n6464), .A2(n6661), .ZN(n10029) );
  AND2_X1 U5878 ( .A1(n10061), .A2(n10060), .ZN(n10062) );
  INV_X1 U5879 ( .A(n6653), .ZN(n8608) );
  AND4_X1 U5880 ( .A1(n5993), .A2(n5992), .A3(n5991), .A4(n5990), .ZN(n7950)
         );
  AOI21_X1 U5881 ( .B1(n6590), .B2(n7766), .A(n4465), .ZN(n4938) );
  NAND2_X1 U5882 ( .A1(n5045), .A2(n5046), .ZN(n7839) );
  NOR2_X1 U5883 ( .A1(n7820), .A2(n7819), .ZN(n7822) );
  OAI21_X1 U5884 ( .B1(n6076), .B2(n4779), .A(n4777), .ZN(n7813) );
  INV_X1 U5885 ( .A(n8219), .ZN(n6079) );
  CLKBUF_X1 U5886 ( .A(n7448), .Z(n4517) );
  NAND2_X1 U5887 ( .A1(n6422), .A2(n7376), .ZN(n6047) );
  CLKBUF_X1 U5888 ( .A(n6422), .Z(n7377) );
  NAND2_X1 U5889 ( .A1(n6329), .A2(n6328), .ZN(n10111) );
  INV_X1 U5890 ( .A(n7958), .ZN(n10190) );
  INV_X1 U5891 ( .A(n10134), .ZN(n10188) );
  INV_X1 U5892 ( .A(n10334), .ZN(n10341) );
  XNOR2_X1 U5893 ( .A(n5756), .B(n5735), .ZN(n8856) );
  INV_X1 U5894 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5981) );
  XNOR2_X1 U5895 ( .A(n5729), .B(n5721), .ZN(n8692) );
  AOI21_X1 U5896 ( .B1(n5689), .B2(n4715), .A(n4714), .ZN(n4713) );
  INV_X1 U5897 ( .A(n5681), .ZN(n4715) );
  INV_X1 U5898 ( .A(n5699), .ZN(n4714) );
  CLKBUF_X1 U5899 ( .A(n6531), .Z(n7016) );
  NAND2_X1 U5900 ( .A1(n5690), .A2(n5689), .ZN(n5700) );
  INV_X1 U5901 ( .A(n5690), .ZN(n5687) );
  NAND2_X1 U5902 ( .A1(n6521), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6523) );
  INV_X1 U5903 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n6526) );
  NAND2_X1 U5904 ( .A1(n4727), .A2(n5594), .ZN(n5652) );
  NAND2_X1 U5905 ( .A1(n4732), .A2(n4730), .ZN(n4727) );
  AND2_X1 U5906 ( .A1(n5631), .A2(n5599), .ZN(n5650) );
  NAND2_X1 U5907 ( .A1(n4732), .A2(n5574), .ZN(n5596) );
  OAI21_X1 U5908 ( .B1(n5469), .B2(n4404), .A(n5017), .ZN(n5512) );
  INV_X1 U5909 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5962) );
  NOR2_X1 U5910 ( .A1(n6070), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n6085) );
  NAND2_X1 U5911 ( .A1(n4504), .A2(n4503), .ZN(n6070) );
  OAI21_X1 U5912 ( .B1(n5470), .B2(n5097), .A(n5153), .ZN(n5197) );
  NOR2_X1 U5913 ( .A1(n10264), .A2(n10263), .ZN(n10265) );
  NAND2_X1 U5914 ( .A1(n10460), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n4580) );
  NAND2_X1 U5915 ( .A1(n7670), .A2(n7669), .ZN(n7775) );
  AND2_X1 U5916 ( .A1(n4879), .A2(n4883), .ZN(n8868) );
  AND2_X1 U5917 ( .A1(n5592), .A2(n5591), .ZN(n8916) );
  NAND2_X1 U5918 ( .A1(n4881), .A2(n4407), .ZN(n4880) );
  NAND2_X1 U5919 ( .A1(n4883), .A2(n8867), .ZN(n4881) );
  NAND2_X1 U5920 ( .A1(n10247), .A2(n5635), .ZN(n5702) );
  NAND2_X1 U5921 ( .A1(n4897), .A2(n8788), .ZN(n7569) );
  INV_X1 U5922 ( .A(n7568), .ZN(n4897) );
  NAND2_X1 U5923 ( .A1(n7618), .A2(n7617), .ZN(n7619) );
  AND2_X1 U5924 ( .A1(n4892), .A2(n7582), .ZN(n7588) );
  NOR2_X1 U5925 ( .A1(n8962), .A2(n4894), .ZN(n4893) );
  INV_X1 U5926 ( .A(n8769), .ZN(n4894) );
  NAND2_X1 U5927 ( .A1(n8900), .A2(n8769), .ZN(n8963) );
  INV_X1 U5929 ( .A(n8992), .ZN(n9013) );
  NAND2_X1 U5930 ( .A1(n7660), .A2(n7571), .ZN(n7687) );
  NAND2_X1 U5931 ( .A1(n4885), .A2(n8813), .ZN(n8998) );
  INV_X1 U5932 ( .A(n7677), .ZN(n9011) );
  OAI21_X1 U5933 ( .B1(n8819), .B2(n7137), .A(n7091), .ZN(n5772) );
  INV_X1 U5934 ( .A(n8862), .ZN(n7142) );
  INV_X1 U5935 ( .A(n8954), .ZN(n9251) );
  OR2_X1 U5936 ( .A1(n4374), .A2(n7163), .ZN(n5139) );
  OR2_X1 U5937 ( .A1(n5260), .A2(n5166), .ZN(n5167) );
  INV_X1 U5938 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10258) );
  NAND2_X1 U5939 ( .A1(n7231), .A2(n7230), .ZN(n7292) );
  INV_X1 U5940 ( .A(n4919), .ZN(n7254) );
  NAND2_X1 U5941 ( .A1(n7262), .A2(n7261), .ZN(n7392) );
  INV_X1 U5942 ( .A(n4917), .ZN(n7257) );
  AND2_X1 U5943 ( .A1(n4917), .A2(n4916), .ZN(n7384) );
  NAND2_X1 U5944 ( .A1(n4919), .A2(n4918), .ZN(n4917) );
  NAND2_X1 U5945 ( .A1(n4662), .A2(n4663), .ZN(n7386) );
  NOR2_X1 U5946 ( .A1(n7492), .A2(n7491), .ZN(n7727) );
  INV_X1 U5947 ( .A(n4914), .ZN(n8138) );
  INV_X1 U5948 ( .A(n4667), .ZN(n7729) );
  INV_X1 U5949 ( .A(n4912), .ZN(n9038) );
  NAND2_X1 U5950 ( .A1(n9048), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n4911) );
  NOR2_X1 U5951 ( .A1(n8646), .A2(n8645), .ZN(n8676) );
  NAND2_X1 U5952 ( .A1(n9086), .A2(n4905), .ZN(n9089) );
  INV_X1 U5953 ( .A(n10366), .ZN(n9112) );
  AND2_X1 U5954 ( .A1(n7167), .A2(n8854), .ZN(n10362) );
  NAND2_X1 U5955 ( .A1(n5760), .A2(n5759), .ZN(n8844) );
  NAND2_X1 U5956 ( .A1(n5915), .A2(n5914), .ZN(n9440) );
  NAND2_X1 U5957 ( .A1(n5680), .A2(n5890), .ZN(n9196) );
  NAND2_X1 U5958 ( .A1(n9266), .A2(n5058), .ZN(n9223) );
  NOR2_X1 U5959 ( .A1(n9254), .A2(n4634), .ZN(n4633) );
  INV_X1 U5960 ( .A(n4637), .ZN(n4634) );
  INV_X1 U5961 ( .A(n9484), .ZN(n9290) );
  INV_X1 U5962 ( .A(n9328), .ZN(n9318) );
  INV_X1 U5963 ( .A(n4995), .ZN(n9319) );
  OAI21_X1 U5964 ( .B1(n9356), .B2(n4998), .A(n4999), .ZN(n4995) );
  NOR2_X1 U5965 ( .A1(n9356), .A2(n5000), .ZN(n9339) );
  NAND2_X1 U5966 ( .A1(n9140), .A2(n9139), .ZN(n9405) );
  NAND2_X1 U5967 ( .A1(n8548), .A2(n4748), .ZN(n8612) );
  NAND2_X1 U5968 ( .A1(n5075), .A2(n5074), .ZN(n8182) );
  NAND2_X1 U5969 ( .A1(n4739), .A2(n4741), .ZN(n7991) );
  NAND2_X1 U5970 ( .A1(n8499), .A2(n5805), .ZN(n7935) );
  AOI22_X1 U5971 ( .A1(n4810), .A2(n9411), .B1(n9033), .B2(n9412), .ZN(n8502)
         );
  INV_X1 U5972 ( .A(n4755), .ZN(n4754) );
  OAI21_X1 U5973 ( .B1(n5514), .B2(n4757), .A(n4756), .ZN(n4755) );
  INV_X1 U5974 ( .A(n9425), .ZN(n9354) );
  NAND2_X1 U5975 ( .A1(n9427), .A2(n7886), .ZN(n9429) );
  OAI211_X1 U5976 ( .C1(n10414), .C2(n9462), .A(n5038), .B(n4458), .ZN(n9565)
         );
  INV_X1 U5977 ( .A(n9459), .ZN(n5038) );
  AND2_X1 U5978 ( .A1(n9461), .A2(n10408), .ZN(n5037) );
  NOR2_X1 U5979 ( .A1(n4628), .A2(n4627), .ZN(n4626) );
  INV_X1 U5980 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n9585) );
  AND3_X1 U5981 ( .A1(n4448), .A2(n5127), .A3(n5131), .ZN(n4831) );
  AND2_X1 U5982 ( .A1(n5951), .A2(n5143), .ZN(n8193) );
  NAND2_X1 U5983 ( .A1(n5766), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5751) );
  INV_X1 U5984 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n7115) );
  INV_X1 U5985 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n7095) );
  INV_X1 U5986 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n7025) );
  INV_X1 U5987 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6996) );
  INV_X1 U5988 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6993) );
  INV_X1 U5989 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6971) );
  AND2_X1 U5990 ( .A1(n5208), .A2(n5158), .ZN(n5090) );
  NAND2_X1 U5991 ( .A1(n5133), .A2(n5157), .ZN(n5158) );
  NAND2_X1 U5992 ( .A1(n4657), .A2(n10367), .ZN(n4656) );
  NAND2_X1 U5993 ( .A1(n4655), .A2(n5133), .ZN(n4654) );
  NAND2_X1 U5994 ( .A1(n4687), .A2(n4688), .ZN(n7746) );
  NAND2_X1 U5995 ( .A1(n6746), .A2(n4689), .ZN(n4687) );
  AND4_X1 U5996 ( .A1(n6199), .A2(n6198), .A3(n6197), .A4(n6196), .ZN(n9612)
         );
  AOI22_X1 U5997 ( .A1(n7401), .A2(n7400), .B1(n6739), .B2(n6738), .ZN(n7482)
         );
  NAND2_X1 U5998 ( .A1(n9740), .A2(n5028), .ZN(n6935) );
  NOR2_X1 U5999 ( .A1(n9594), .A2(n4410), .ZN(n5028) );
  XNOR2_X1 U6000 ( .A(n6861), .B(n6860), .ZN(n9641) );
  INV_X1 U6001 ( .A(n6759), .ZN(n7844) );
  NAND2_X1 U6002 ( .A1(n5027), .A2(n9616), .ZN(n9684) );
  NAND2_X1 U6003 ( .A1(n9617), .A2(n9619), .ZN(n5027) );
  AND4_X1 U6004 ( .A1(n6016), .A2(n6015), .A3(n6014), .A4(n6013), .ZN(n8530)
         );
  NAND2_X1 U6005 ( .A1(n5026), .A2(n6873), .ZN(n9713) );
  OR2_X1 U6006 ( .A1(n5026), .A2(n6873), .ZN(n9714) );
  NAND2_X1 U6007 ( .A1(n6870), .A2(n6869), .ZN(n5026) );
  INV_X1 U6008 ( .A(n10131), .ZN(n9934) );
  AND2_X1 U6009 ( .A1(n6349), .A2(n6331), .ZN(n9866) );
  AND4_X1 U6010 ( .A1(n6213), .A2(n6212), .A3(n6211), .A4(n6210), .ZN(n9759)
         );
  NAND2_X1 U6011 ( .A1(n6312), .A2(n6311), .ZN(n9926) );
  INV_X1 U6012 ( .A(n9951), .ZN(n9918) );
  OR2_X1 U6013 ( .A1(n6974), .A2(n6949), .ZN(n9778) );
  NAND2_X1 U6014 ( .A1(n6307), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n6033) );
  XNOR2_X1 U6015 ( .A(n7006), .B(n4837), .ZN(n7059) );
  NOR2_X1 U6016 ( .A1(n7059), .A2(n7060), .ZN(n7058) );
  AOI21_X1 U6017 ( .B1(P1_REG2_REG_1__SCAN_IN), .B2(n7052), .A(n7058), .ZN(
        n7331) );
  NOR2_X1 U6018 ( .A1(n7329), .A2(n4855), .ZN(n7072) );
  NOR2_X1 U6019 ( .A1(n7072), .A2(n7071), .ZN(n7070) );
  INV_X1 U6020 ( .A(n4853), .ZN(n4849) );
  NAND2_X1 U6021 ( .A1(n7027), .A2(n7026), .ZN(n4845) );
  AND2_X1 U6022 ( .A1(n4845), .A2(n4847), .ZN(n7038) );
  AND2_X1 U6023 ( .A1(n4841), .A2(n4839), .ZN(n7012) );
  AOI21_X1 U6024 ( .B1(n7005), .B2(n7004), .A(n7040), .ZN(n7082) );
  NAND2_X1 U6025 ( .A1(n7078), .A2(n7079), .ZN(n7176) );
  NAND2_X1 U6026 ( .A1(n4522), .A2(n4521), .ZN(n4520) );
  INV_X1 U6027 ( .A(n7409), .ZN(n4522) );
  AND2_X1 U6028 ( .A1(n7411), .A2(n7410), .ZN(n7413) );
  NAND2_X1 U6029 ( .A1(n4856), .A2(n4861), .ZN(n7431) );
  NAND2_X1 U6030 ( .A1(n7411), .A2(n4862), .ZN(n4856) );
  AOI22_X1 U6031 ( .A1(n7856), .A2(n7855), .B1(n7854), .B2(n7853), .ZN(n8626)
         );
  NOR2_X1 U6032 ( .A1(n7862), .A2(n7861), .ZN(n8633) );
  AND2_X1 U6033 ( .A1(n7860), .A2(n7859), .ZN(n7862) );
  NOR2_X1 U6034 ( .A1(n9804), .A2(n9805), .ZN(n9803) );
  NOR2_X1 U6035 ( .A1(n9797), .A2(n8712), .ZN(n9814) );
  NOR2_X1 U6036 ( .A1(n9814), .A2(n9813), .ZN(n9812) );
  INV_X1 U6037 ( .A(n4836), .ZN(n9831) );
  INV_X1 U6038 ( .A(n4834), .ZN(n10289) );
  NAND2_X1 U6039 ( .A1(n9856), .A2(n10055), .ZN(n9858) );
  NAND2_X1 U6040 ( .A1(n9875), .A2(n9874), .ZN(n9876) );
  INV_X1 U6041 ( .A(n10111), .ZN(n9868) );
  INV_X1 U6042 ( .A(n4547), .ZN(n4546) );
  AOI22_X1 U6043 ( .A1(n9888), .A2(n10055), .B1(n10057), .B2(n9919), .ZN(n4547) );
  INV_X1 U6044 ( .A(n10116), .ZN(n9885) );
  CLKBUF_X1 U6045 ( .A(n9892), .Z(n9893) );
  OAI21_X1 U6046 ( .B1(n9941), .B2(n4934), .A(n4932), .ZN(n9905) );
  NAND2_X1 U6047 ( .A1(n4937), .A2(n5092), .ZN(n9930) );
  NAND2_X1 U6048 ( .A1(n9941), .A2(n9947), .ZN(n4937) );
  NAND2_X1 U6049 ( .A1(n4967), .A2(n6667), .ZN(n9948) );
  NAND2_X1 U6050 ( .A1(n9976), .A2(n6666), .ZN(n9957) );
  NAND2_X1 U6051 ( .A1(n4922), .A2(n4373), .ZN(n9991) );
  NAND2_X1 U6052 ( .A1(n4532), .A2(n4424), .ZN(n4922) );
  NOR2_X1 U6053 ( .A1(n4532), .A2(n6613), .ZN(n10012) );
  INV_X1 U6054 ( .A(n4977), .ZN(n4976) );
  OAI22_X1 U6055 ( .A1(n6382), .A2(n6959), .B1(n6977), .B2(n7037), .ZN(n4977)
         );
  NAND2_X1 U6056 ( .A1(n7704), .A2(n6496), .ZN(n7759) );
  NAND2_X1 U6057 ( .A1(n4797), .A2(n4795), .ZN(n10237) );
  NOR2_X1 U6058 ( .A1(n5971), .A2(n4796), .ZN(n4795) );
  NAND2_X1 U6059 ( .A1(n5974), .A2(n5981), .ZN(n4796) );
  XNOR2_X1 U6060 ( .A(n5716), .B(n5715), .ZN(n10247) );
  OAI21_X1 U6061 ( .B1(n5682), .B2(n5688), .A(n4713), .ZN(n5716) );
  INV_X1 U6062 ( .A(n6688), .ZN(n7892) );
  INV_X1 U6063 ( .A(n7419), .ZN(n7744) );
  INV_X1 U6064 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n8428) );
  INV_X1 U6065 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6998) );
  XNOR2_X1 U6066 ( .A(n6113), .B(P1_IR_REG_7__SCAN_IN), .ZN(n7080) );
  INV_X1 U6067 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6943) );
  INV_X1 U6068 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6944) );
  INV_X1 U6069 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6958) );
  NAND2_X1 U6070 ( .A1(n4518), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6051) );
  INV_X1 U6071 ( .A(n6049), .ZN(n4518) );
  AND2_X1 U6072 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n10265), .ZN(n10461) );
  XNOR2_X1 U6073 ( .A(n10270), .B(n10269), .ZN(n10472) );
  XNOR2_X1 U6074 ( .A(n10273), .B(n4563), .ZN(n10471) );
  NAND2_X1 U6075 ( .A1(n10435), .A2(n4581), .ZN(n10434) );
  NOR2_X1 U6076 ( .A1(n10433), .A2(n4582), .ZN(n4581) );
  NOR2_X1 U6077 ( .A1(n10284), .A2(n10283), .ZN(n4582) );
  NAND2_X1 U6078 ( .A1(n10434), .A2(n10285), .ZN(n10465) );
  AOI21_X1 U6079 ( .B1(n9019), .B2(n9464), .A(n8812), .ZN(n4564) );
  INV_X1 U6080 ( .A(n8811), .ZN(n4565) );
  AND2_X1 U6081 ( .A1(n8961), .A2(n4534), .ZN(n4533) );
  NAND2_X1 U6082 ( .A1(n8955), .A2(n4536), .ZN(n4535) );
  OAI21_X1 U6083 ( .B1(n7782), .B2(n9037), .A(n4811), .ZN(P2_U3557) );
  NAND2_X1 U6084 ( .A1(n9037), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n4811) );
  INV_X1 U6085 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n9132) );
  NAND2_X1 U6086 ( .A1(n4603), .A2(n4607), .ZN(n9130) );
  NAND2_X1 U6087 ( .A1(n10424), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n4749) );
  NAND2_X1 U6088 ( .A1(n9563), .A2(n10426), .ZN(n4750) );
  NAND2_X1 U6089 ( .A1(n10416), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n4555) );
  NAND2_X1 U6090 ( .A1(n4678), .A2(n8526), .ZN(n4677) );
  INV_X1 U6091 ( .A(n4868), .ZN(n4577) );
  NAND2_X1 U6092 ( .A1(n4869), .A2(n10310), .ZN(n4579) );
  OR2_X1 U6093 ( .A1(n8718), .A2(n10310), .ZN(n4578) );
  AND2_X1 U6094 ( .A1(n10079), .A2(n10064), .ZN(n9839) );
  NOR2_X1 U6095 ( .A1(n6710), .A2(n6709), .ZN(n6711) );
  OAI211_X1 U6096 ( .C1(n10110), .C2(n10074), .A(n4602), .B(n4433), .ZN(
        P1_U3264) );
  XNOR2_X1 U6097 ( .A(n5765), .B(P2_IR_REG_20__SCAN_IN), .ZN(n7543) );
  AND2_X1 U6098 ( .A1(n10111), .A2(n9888), .ZN(n6623) );
  OR2_X1 U6099 ( .A1(n10111), .A2(n9888), .ZN(n4403) );
  INV_X1 U6100 ( .A(n5916), .ZN(n9228) );
  AND2_X1 U6101 ( .A1(n9207), .A2(n5889), .ZN(n5916) );
  NAND2_X1 U6102 ( .A1(n7892), .A2(n10310), .ZN(n7368) );
  INV_X1 U6103 ( .A(n6873), .ZN(n5025) );
  OR2_X1 U6104 ( .A1(n5505), .A2(n5019), .ZN(n4404) );
  NAND2_X1 U6105 ( .A1(n8846), .A2(n5062), .ZN(n9340) );
  NAND2_X1 U6106 ( .A1(n10154), .A2(n10004), .ZN(n4405) );
  AND2_X1 U6107 ( .A1(n4954), .A2(n4452), .ZN(n4406) );
  INV_X1 U6108 ( .A(n5914), .ZN(n5085) );
  INV_X1 U6109 ( .A(n9947), .ZN(n4933) );
  NAND2_X1 U6110 ( .A1(n8817), .A2(n8818), .ZN(n4407) );
  OR2_X1 U6111 ( .A1(n4437), .A2(n5010), .ZN(n4408) );
  AND3_X1 U6112 ( .A1(n8131), .A2(n5068), .A3(n5067), .ZN(n4409) );
  AND2_X1 U6113 ( .A1(n6899), .A2(n6898), .ZN(n4410) );
  NAND2_X1 U6114 ( .A1(n8621), .A2(n4435), .ZN(n9140) );
  NAND2_X1 U6115 ( .A1(n5378), .A2(n5377), .ZN(n9536) );
  INV_X1 U6116 ( .A(n9536), .ZN(n5067) );
  NAND2_X1 U6117 ( .A1(n8209), .A2(n7848), .ZN(n6586) );
  AND2_X1 U6118 ( .A1(n4679), .A2(n4459), .ZN(n4411) );
  INV_X1 U6119 ( .A(n6623), .ZN(n4946) );
  OR2_X1 U6120 ( .A1(n10144), .A2(n9953), .ZN(n6667) );
  INV_X1 U6121 ( .A(n6667), .ZN(n4969) );
  NOR2_X1 U6122 ( .A1(n10079), .A2(n4698), .ZN(n6452) );
  AOI21_X1 U6123 ( .B1(n9193), .B2(n5698), .A(n5697), .ZN(n8825) );
  NOR2_X1 U6124 ( .A1(n5085), .A2(n4494), .ZN(n4412) );
  AOI21_X1 U6125 ( .B1(n5447), .B2(n5446), .A(n4709), .ZN(n4708) );
  AND4_X1 U6126 ( .A1(n5913), .A2(n9179), .A3(n4523), .A4(n9154), .ZN(n4413)
         );
  AND2_X1 U6127 ( .A1(n5909), .A2(n5086), .ZN(n4414) );
  INV_X1 U6128 ( .A(n4983), .ZN(n4982) );
  OAI21_X1 U6129 ( .B1(n9154), .B2(n4436), .A(n4984), .ZN(n4983) );
  NAND2_X1 U6130 ( .A1(n4476), .A2(n4791), .ZN(n4415) );
  AND2_X1 U6131 ( .A1(n4623), .A2(n10399), .ZN(n4416) );
  NOR2_X1 U6132 ( .A1(n4943), .A2(n6624), .ZN(n4417) );
  AND2_X1 U6133 ( .A1(n5046), .A2(n5044), .ZN(n4418) );
  AND2_X1 U6134 ( .A1(n5651), .A2(n4730), .ZN(n4419) );
  OR2_X1 U6135 ( .A1(n4826), .A2(n5890), .ZN(n4420) );
  NAND2_X1 U6136 ( .A1(n5895), .A2(n5898), .ZN(n9195) );
  NAND2_X1 U6137 ( .A1(n7557), .A2(n9373), .ZN(n9019) );
  NAND2_X1 U6138 ( .A1(n7788), .A2(n7789), .ZN(n7931) );
  NAND2_X1 U6139 ( .A1(n5820), .A2(n5817), .ZN(n7968) );
  NAND2_X1 U6140 ( .A1(n9119), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n4421) );
  NAND2_X1 U6141 ( .A1(n5461), .A2(n5460), .ZN(n9398) );
  OR2_X1 U6142 ( .A1(n9595), .A2(n9594), .ZN(n4423) );
  OR2_X1 U6143 ( .A1(n10158), .A2(n10019), .ZN(n4424) );
  NOR2_X1 U6144 ( .A1(n6671), .A2(n9914), .ZN(n4425) );
  OAI21_X1 U6145 ( .B1(n9702), .B2(n5005), .A(n5003), .ZN(n9625) );
  NAND2_X1 U6146 ( .A1(n4973), .A2(n6652), .ZN(n8093) );
  AND2_X1 U6147 ( .A1(n4967), .A2(n4968), .ZN(n9911) );
  INV_X1 U6148 ( .A(n10345), .ZN(n7819) );
  NAND2_X1 U6149 ( .A1(n6030), .A2(n8861), .ZN(n6048) );
  NAND2_X1 U6150 ( .A1(n9638), .A2(n6867), .ZN(n4426) );
  AND3_X1 U6151 ( .A1(n5567), .A2(n9275), .A3(n5919), .ZN(n4427) );
  AND2_X1 U6152 ( .A1(n6876), .A2(n5024), .ZN(n4428) );
  NAND2_X1 U6153 ( .A1(n5446), .A2(n5434), .ZN(n5447) );
  AND2_X1 U6154 ( .A1(n5292), .A2(SI_7_), .ZN(n4429) );
  NAND2_X1 U6155 ( .A1(n9693), .A2(n6868), .ZN(n4430) );
  OR3_X1 U6156 ( .A1(n8814), .A2(n4884), .A3(n7677), .ZN(n4431) );
  INV_X1 U6157 ( .A(n6837), .ZN(n4505) );
  OR2_X1 U6158 ( .A1(n10011), .A2(n9669), .ZN(n4432) );
  OR2_X1 U6159 ( .A1(n10109), .A2(n10317), .ZN(n4433) );
  OR2_X1 U6160 ( .A1(n6100), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n4434) );
  AND2_X1 U6161 ( .A1(n8622), .A2(n8620), .ZN(n4435) );
  OR2_X1 U6162 ( .A1(n9468), .A2(n8954), .ZN(n9206) );
  NAND2_X1 U6163 ( .A1(n9152), .A2(n9197), .ZN(n4436) );
  XNOR2_X1 U6164 ( .A(n5292), .B(n4699), .ZN(n5290) );
  INV_X1 U6165 ( .A(n5290), .ZN(n5014) );
  NOR2_X1 U6166 ( .A1(n8845), .A2(n9526), .ZN(n8846) );
  AND2_X1 U6167 ( .A1(n9629), .A2(n9628), .ZN(n4437) );
  INV_X1 U6168 ( .A(n8813), .ZN(n4884) );
  AOI21_X1 U6169 ( .B1(n5003), .B2(n5005), .A(n4408), .ZN(n4674) );
  NOR2_X1 U6170 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n5749) );
  INV_X1 U6171 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5533) );
  INV_X1 U6172 ( .A(n10407), .ZN(n5059) );
  OR3_X1 U6173 ( .A1(n10088), .A2(n10188), .A3(n10095), .ZN(n4438) );
  AND2_X1 U6174 ( .A1(n9541), .A2(n8657), .ZN(n5819) );
  OR2_X1 U6175 ( .A1(n10126), .A2(n9926), .ZN(n4439) );
  AND2_X1 U6176 ( .A1(n4886), .A2(n4888), .ZN(n4440) );
  NAND2_X1 U6177 ( .A1(n9475), .A2(n9281), .ZN(n5879) );
  INV_X1 U6178 ( .A(n5879), .ZN(n5034) );
  NAND2_X1 U6179 ( .A1(n9452), .A2(n9198), .ZN(n4441) );
  AND2_X1 U6180 ( .A1(n6418), .A2(n6184), .ZN(n4442) );
  AND3_X1 U6181 ( .A1(n10036), .A2(n4804), .A3(n4799), .ZN(n4443) );
  AND2_X1 U6182 ( .A1(n5060), .A2(n5059), .ZN(n4444) );
  NAND2_X1 U6183 ( .A1(n9206), .A2(n5917), .ZN(n9242) );
  NAND2_X1 U6184 ( .A1(n4635), .A2(n4637), .ZN(n9253) );
  AND2_X1 U6185 ( .A1(n4839), .A2(n7013), .ZN(n4445) );
  AND2_X1 U6186 ( .A1(n7773), .A2(n7772), .ZN(n4446) );
  AND2_X1 U6187 ( .A1(n4834), .A2(n4833), .ZN(n4447) );
  AND2_X1 U6188 ( .A1(n5130), .A2(n5144), .ZN(n4448) );
  NAND2_X1 U6189 ( .A1(n5602), .A2(n5601), .ZN(n9475) );
  OR2_X1 U6190 ( .A1(n10107), .A2(n9745), .ZN(n6683) );
  INV_X1 U6191 ( .A(n6683), .ZN(n4962) );
  INV_X1 U6192 ( .A(n5932), .ZN(n8557) );
  AND2_X1 U6193 ( .A1(n5916), .A2(n9242), .ZN(n4449) );
  AND2_X1 U6194 ( .A1(n9249), .A2(n5033), .ZN(n4450) );
  INV_X1 U6195 ( .A(n7968), .ZN(n7970) );
  INV_X1 U6196 ( .A(n5002), .ZN(n6713) );
  NAND2_X1 U6197 ( .A1(n5723), .A2(n5722), .ZN(n9438) );
  INV_X1 U6198 ( .A(n9364), .ZN(n9357) );
  OR2_X1 U6199 ( .A1(n7069), .A2(n7001), .ZN(n4451) );
  NAND2_X1 U6200 ( .A1(n6665), .A2(n6664), .ZN(n4452) );
  AND2_X1 U6201 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_REG3_REG_9__SCAN_IN), 
        .ZN(n4453) );
  INV_X1 U6202 ( .A(n6060), .ZN(n4504) );
  AND2_X1 U6204 ( .A1(n9237), .A2(n4625), .ZN(n4454) );
  NAND2_X1 U6205 ( .A1(n5480), .A2(n5479), .ZN(n9499) );
  INV_X1 U6206 ( .A(n9499), .ZN(n9345) );
  INV_X1 U6207 ( .A(n4809), .ZN(n7781) );
  OR2_X1 U6208 ( .A1(n4423), .A2(n4410), .ZN(n4455) );
  INV_X1 U6209 ( .A(n5001), .ZN(n5000) );
  AND2_X1 U6210 ( .A1(n4953), .A2(n6492), .ZN(n4456) );
  INV_X1 U6211 ( .A(n4639), .ZN(n4638) );
  NAND2_X1 U6212 ( .A1(n9290), .A2(n9280), .ZN(n4639) );
  OR2_X1 U6213 ( .A1(n8209), .A2(n7848), .ZN(n6587) );
  NOR2_X1 U6214 ( .A1(n6769), .A2(n6768), .ZN(n4457) );
  NOR2_X1 U6215 ( .A1(n9460), .A2(n5037), .ZN(n4458) );
  INV_X1 U6216 ( .A(n5055), .ZN(n9894) );
  NOR2_X1 U6217 ( .A1(n4531), .A2(n10121), .ZN(n5055) );
  OR2_X1 U6218 ( .A1(n4681), .A2(n9738), .ZN(n4459) );
  INV_X1 U6219 ( .A(n7430), .ZN(n4864) );
  AND2_X1 U6220 ( .A1(n7429), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n7430) );
  INV_X1 U6221 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n8247) );
  INV_X1 U6222 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n8418) );
  AND2_X1 U6223 ( .A1(n6905), .A2(n6904), .ZN(n9594) );
  NOR2_X1 U6224 ( .A1(n6663), .A2(n6455), .ZN(n4956) );
  NAND2_X1 U6225 ( .A1(n8551), .A2(n8552), .ZN(n4460) );
  NAND2_X1 U6226 ( .A1(n7008), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n4461) );
  AND3_X1 U6227 ( .A1(n5833), .A2(n5911), .A3(n5834), .ZN(n4462) );
  AND2_X1 U6228 ( .A1(n10131), .A2(n9951), .ZN(n4463) );
  AND2_X1 U6229 ( .A1(n9495), .A2(n9312), .ZN(n4464) );
  NAND2_X1 U6230 ( .A1(n10140), .A2(n6857), .ZN(n9912) );
  NAND2_X1 U6231 ( .A1(n6684), .A2(n6683), .ZN(n4769) );
  AND2_X1 U6232 ( .A1(n10345), .A2(n6591), .ZN(n4465) );
  AND2_X1 U6233 ( .A1(n4980), .A2(n4978), .ZN(n4466) );
  AND2_X1 U6234 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .ZN(
        n4467) );
  INV_X1 U6235 ( .A(n4685), .ZN(n4684) );
  NAND2_X1 U6236 ( .A1(n4688), .A2(n4686), .ZN(n4685) );
  INV_X1 U6237 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6968) );
  NAND2_X1 U6238 ( .A1(n5077), .A2(n5834), .ZN(n4468) );
  INV_X1 U6239 ( .A(n6482), .ZN(n4807) );
  NAND2_X1 U6240 ( .A1(n5622), .A2(n5621), .ZN(n9464) );
  INV_X1 U6241 ( .A(n9464), .ZN(n5057) );
  NAND2_X1 U6242 ( .A1(n6683), .A2(n6412), .ZN(n8838) );
  INV_X1 U6243 ( .A(n4705), .ZN(n4704) );
  NAND2_X1 U6244 ( .A1(n5017), .A2(n4706), .ZN(n4705) );
  NOR2_X1 U6245 ( .A1(n9364), .A2(n5852), .ZN(n5859) );
  OR2_X1 U6246 ( .A1(n9716), .A2(n5025), .ZN(n4469) );
  OR2_X1 U6247 ( .A1(n8997), .A2(n4884), .ZN(n4470) );
  OR2_X1 U6248 ( .A1(n10168), .A2(n9612), .ZN(n6659) );
  INV_X1 U6249 ( .A(n9208), .ZN(n4979) );
  AND3_X1 U6250 ( .A1(n9228), .A2(n9242), .A3(n9220), .ZN(n4471) );
  OR2_X1 U6251 ( .A1(n5913), .A2(n5911), .ZN(n4472) );
  OR2_X1 U6252 ( .A1(n9495), .A2(n9349), .ZN(n5563) );
  INV_X1 U6253 ( .A(n5563), .ZN(n4816) );
  AND2_X1 U6254 ( .A1(n10109), .A2(n10108), .ZN(n4473) );
  NAND2_X1 U6255 ( .A1(n5702), .A2(n5701), .ZN(n9452) );
  NOR2_X1 U6256 ( .A1(n6936), .A2(n9737), .ZN(n4474) );
  AND2_X1 U6257 ( .A1(n5361), .A2(n5346), .ZN(n4475) );
  AND2_X1 U6258 ( .A1(n6415), .A2(n6417), .ZN(n4476) );
  AND2_X1 U6259 ( .A1(n4968), .A2(n6669), .ZN(n4477) );
  AND2_X1 U6260 ( .A1(n5919), .A2(n5918), .ZN(n9278) );
  INV_X1 U6261 ( .A(n9278), .ZN(n4636) );
  OR2_X1 U6262 ( .A1(n6991), .A2(n6090), .ZN(n4478) );
  AND2_X1 U6263 ( .A1(n8548), .A2(n5836), .ZN(n4479) );
  NOR2_X1 U6264 ( .A1(n6877), .A2(n9619), .ZN(n4480) );
  AND2_X1 U6265 ( .A1(n4786), .A2(n6667), .ZN(n4481) );
  AND2_X1 U6266 ( .A1(n9154), .A2(n5890), .ZN(n4482) );
  AND2_X1 U6267 ( .A1(n4663), .A2(n4661), .ZN(n4483) );
  AND2_X1 U6268 ( .A1(n9154), .A2(n5894), .ZN(n4484) );
  AND2_X1 U6269 ( .A1(n5651), .A2(n4729), .ZN(n4485) );
  AND2_X1 U6270 ( .A1(n5884), .A2(n5916), .ZN(n4486) );
  NAND2_X1 U6271 ( .A1(n7782), .A2(n4809), .ZN(n5780) );
  INV_X1 U6272 ( .A(n6825), .ZN(n5009) );
  OR2_X1 U6273 ( .A1(n4728), .A2(n5575), .ZN(n4487) );
  AND2_X1 U6274 ( .A1(n5775), .A2(n5907), .ZN(n5913) );
  AOI21_X1 U6275 ( .B1(n9702), .B2(n6826), .A(n6825), .ZN(n5006) );
  NOR2_X1 U6276 ( .A1(n5754), .A2(SI_30_), .ZN(n4488) );
  INV_X1 U6277 ( .A(n4896), .ZN(n7315) );
  NAND2_X1 U6278 ( .A1(n5926), .A2(n7537), .ZN(n4896) );
  AND2_X1 U6279 ( .A1(n7996), .A2(n8008), .ZN(n7980) );
  INV_X1 U6280 ( .A(n6645), .ZN(n4975) );
  AND2_X1 U6281 ( .A1(n6659), .A2(n6658), .ZN(n10036) );
  INV_X1 U6282 ( .A(n10036), .ZN(n4806) );
  INV_X1 U6283 ( .A(n6492), .ZN(n4952) );
  NAND2_X1 U6284 ( .A1(n5693), .A2(n5692), .ZN(n9454) );
  INV_X1 U6285 ( .A(n9454), .ZN(n4985) );
  AND2_X1 U6286 ( .A1(n5758), .A2(n4488), .ZN(n4489) );
  AND2_X1 U6287 ( .A1(n8621), .A2(n8620), .ZN(n4490) );
  NAND2_X1 U6288 ( .A1(n7967), .A2(n7966), .ZN(n7969) );
  INV_X1 U6289 ( .A(n5045), .ZN(n7820) );
  NAND2_X1 U6290 ( .A1(n4537), .A2(n4900), .ZN(n4491) );
  INV_X1 U6291 ( .A(n4720), .ZN(n4719) );
  NAND2_X1 U6292 ( .A1(n4725), .A2(n5758), .ZN(n4720) );
  AND2_X1 U6293 ( .A1(n4720), .A2(n4721), .ZN(n4492) );
  NAND2_X1 U6294 ( .A1(n8632), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4493) );
  INV_X1 U6295 ( .A(n9737), .ZN(n8526) );
  AND2_X1 U6296 ( .A1(n7189), .A2(n6907), .ZN(n10207) );
  NAND2_X1 U6297 ( .A1(n8060), .A2(n5060), .ZN(n7939) );
  INV_X1 U6298 ( .A(n9837), .ZN(n4698) );
  INV_X1 U6299 ( .A(n10399), .ZN(n10414) );
  NOR2_X1 U6300 ( .A1(n7099), .A2(n7757), .ZN(n4494) );
  NAND2_X1 U6301 ( .A1(n6497), .A2(n6492), .ZN(n7812) );
  INV_X1 U6302 ( .A(n7812), .ZN(n4774) );
  INV_X1 U6303 ( .A(n10206), .ZN(n5044) );
  AND2_X1 U6304 ( .A1(n8713), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n4495) );
  INV_X1 U6305 ( .A(n7748), .ZN(n5047) );
  NOR2_X1 U6306 ( .A1(n7413), .A2(n7412), .ZN(n4496) );
  INV_X1 U6307 ( .A(n9541), .ZN(n5068) );
  NOR2_X1 U6308 ( .A1(n9121), .A2(n9122), .ZN(n4497) );
  OR2_X1 U6309 ( .A1(n4421), .A2(n4660), .ZN(n4498) );
  AND2_X1 U6310 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n4499) );
  AND2_X1 U6311 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n4500) );
  INV_X1 U6312 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n4521) );
  NAND2_X1 U6313 ( .A1(n7157), .A2(n7158), .ZN(n4903) );
  NAND2_X1 U6314 ( .A1(n4845), .A2(n4843), .ZN(n4501) );
  INV_X1 U6315 ( .A(n4847), .ZN(n4846) );
  NAND2_X1 U6316 ( .A1(n7037), .A2(n7010), .ZN(n4847) );
  AND2_X1 U6317 ( .A1(n4852), .A2(n4849), .ZN(n4502) );
  INV_X1 U6318 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n4503) );
  INV_X1 U6319 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n4757) );
  INV_X1 U6320 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n4837) );
  INV_X1 U6321 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n4554) );
  INV_X1 U6322 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n4539) );
  INV_X1 U6323 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n4563) );
  INV_X1 U6324 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n4530) );
  AOI21_X1 U6325 ( .B1(n10106), .B2(n10077), .A(n8843), .ZN(n4602) );
  NAND2_X1 U6326 ( .A1(n10089), .A2(n10077), .ZN(n6708) );
  NAND2_X1 U6327 ( .A1(n9210), .A2(n4402), .ZN(n5039) );
  OR2_X1 U6328 ( .A1(n6291), .A2(n7368), .ZN(n4765) );
  OR2_X1 U6329 ( .A1(n6182), .A2(n7368), .ZN(n4804) );
  INV_X1 U6330 ( .A(n7368), .ZN(n4791) );
  OR2_X1 U6331 ( .A1(n6179), .A2(n7368), .ZN(n4805) );
  AND2_X1 U6332 ( .A1(n6656), .A2(n7368), .ZN(n4803) );
  NAND2_X1 U6333 ( .A1(n4776), .A2(n7368), .ZN(n4775) );
  NAND2_X2 U6334 ( .A1(n6690), .A2(n6689), .ZN(n10099) );
  INV_X1 U6335 ( .A(n4843), .ZN(n4842) );
  INV_X1 U6336 ( .A(n7039), .ZN(n4844) );
  NAND2_X1 U6337 ( .A1(n4562), .A2(n4560), .ZN(n4869) );
  AOI21_X1 U6338 ( .B1(n10293), .B2(P1_REG2_REG_18__SCAN_IN), .A(n4447), .ZN(
        n8705) );
  NOR2_X1 U6339 ( .A1(n9809), .A2(n4495), .ZN(n9833) );
  XNOR2_X1 U6340 ( .A(n6836), .B(n4505), .ZN(n9676) );
  NAND2_X1 U6341 ( .A1(n4545), .A2(n4474), .ZN(n6937) );
  NAND2_X1 U6342 ( .A1(n4506), .A2(n4486), .ZN(n5888) );
  NAND3_X1 U6343 ( .A1(n5882), .A2(n5881), .A3(n4584), .ZN(n4506) );
  AOI21_X2 U6344 ( .B1(n4828), .B2(n4827), .A(n7543), .ZN(n5943) );
  NOR2_X1 U6345 ( .A1(n5796), .A2(n4812), .ZN(n5804) );
  OAI22_X1 U6346 ( .A1(n5906), .A2(n5905), .B1(n5914), .B2(n5911), .ZN(n5908)
         );
  NAND2_X1 U6347 ( .A1(n9584), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5132) );
  NAND4_X1 U6348 ( .A1(n4507), .A2(n5960), .A3(n5961), .A4(n5959), .ZN(
        P2_U3244) );
  NAND2_X1 U6349 ( .A1(n5888), .A2(n4509), .ZN(n4821) );
  NAND2_X1 U6350 ( .A1(n5782), .A2(n5877), .ZN(n4528) );
  OAI21_X1 U6351 ( .B1(n5832), .B2(n5831), .A(n4586), .ZN(n5843) );
  AOI21_X2 U6352 ( .B1(n7428), .B2(n7427), .A(n4519), .ZN(n7717) );
  NOR2_X1 U6353 ( .A1(n7041), .A2(n7042), .ZN(n7040) );
  OAI22_X1 U6354 ( .A1(n8626), .A2(n8625), .B1(n8632), .B2(
        P1_REG1_REG_13__SCAN_IN), .ZN(n8629) );
  NOR2_X1 U6355 ( .A1(n9826), .A2(n9825), .ZN(n9824) );
  OAI22_X1 U6356 ( .A1(n7082), .A2(n7081), .B1(n7080), .B2(
        P1_REG1_REG_7__SCAN_IN), .ZN(n7083) );
  NOR2_X1 U6357 ( .A1(n9784), .A2(n9785), .ZN(n9783) );
  AOI21_X1 U6358 ( .B1(P1_REG1_REG_8__SCAN_IN), .B2(n7177), .A(n7172), .ZN(
        n7173) );
  XNOR2_X1 U6359 ( .A(n9802), .B(n8710), .ZN(n9796) );
  AOI21_X1 U6360 ( .B1(n9829), .B2(P1_REG1_REG_17__SCAN_IN), .A(n9824), .ZN(
        n10299) );
  XNOR2_X1 U6361 ( .A(n4558), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n8714) );
  NAND2_X1 U6362 ( .A1(n7407), .A2(n4520), .ZN(n7428) );
  AND2_X2 U6363 ( .A1(n9178), .A2(n5714), .ZN(n9160) );
  NAND2_X1 U6364 ( .A1(n9200), .A2(n5895), .ZN(n9180) );
  NAND2_X1 U6365 ( .A1(n4737), .A2(n4739), .ZN(n4516) );
  AOI21_X1 U6366 ( .B1(n4873), .B2(n4875), .A(n4871), .ZN(n4870) );
  NAND2_X1 U6367 ( .A1(n7918), .A2(n7917), .ZN(n8168) );
  INV_X1 U6368 ( .A(n7654), .ZN(n4515) );
  INV_X1 U6369 ( .A(n7644), .ZN(n4874) );
  NAND2_X1 U6370 ( .A1(n5091), .A2(n7571), .ZN(n7663) );
  NAND2_X1 U6371 ( .A1(n4565), .A2(n4564), .ZN(P2_U3227) );
  OAI21_X1 U6372 ( .B1(n8742), .B2(n8741), .A(n8740), .ZN(n8923) );
  NAND2_X2 U6373 ( .A1(n8893), .A2(n8892), .ZN(n8951) );
  OAI22_X2 U6374 ( .A1(n7985), .A2(n7791), .B1(n7999), .B2(n7936), .ZN(n7794)
         );
  NAND2_X2 U6375 ( .A1(n7793), .A2(n7792), .ZN(n7967) );
  NAND2_X1 U6376 ( .A1(n7642), .A2(n7641), .ZN(n7643) );
  OAI21_X1 U6377 ( .B1(n4986), .B2(n9154), .A(n4982), .ZN(n9177) );
  NAND2_X1 U6378 ( .A1(n4535), .A2(n4533), .ZN(P2_U3231) );
  NAND2_X2 U6379 ( .A1(n7565), .A2(n7884), .ZN(n7583) );
  OR2_X1 U6380 ( .A1(n6090), .A2(n6985), .ZN(n6037) );
  NAND2_X1 U6381 ( .A1(n7947), .A2(n6651), .ZN(n4973) );
  NAND2_X1 U6382 ( .A1(n6542), .A2(n6541), .ZN(n7512) );
  INV_X1 U6383 ( .A(n4974), .ZN(n7894) );
  AOI211_X2 U6384 ( .C1(n10052), .C2(n10112), .A(n9879), .B(n9878), .ZN(n9880)
         );
  NAND2_X1 U6385 ( .A1(n7894), .A2(n6647), .ZN(n8032) );
  NAND2_X1 U6386 ( .A1(n9915), .A2(n6675), .ZN(n9898) );
  NAND2_X1 U6387 ( .A1(n6678), .A2(n6677), .ZN(n9887) );
  NOR2_X1 U6388 ( .A1(n10028), .A2(n10029), .ZN(n10027) );
  NAND2_X2 U6389 ( .A1(n7976), .A2(n5817), .ZN(n8077) );
  NAND2_X1 U6390 ( .A1(n5680), .A2(n4482), .ZN(n9200) );
  INV_X1 U6391 ( .A(n5784), .ZN(n7877) );
  AOI21_X1 U6392 ( .B1(n8145), .B2(n8146), .A(n9047), .ZN(n8148) );
  NOR3_X1 U6393 ( .A1(n10098), .A2(n10097), .A3(n10096), .ZN(n4568) );
  NAND2_X1 U6394 ( .A1(n4797), .A2(n4794), .ZN(n4574) );
  NAND2_X1 U6395 ( .A1(n10094), .A2(n10092), .ZN(n4567) );
  OAI21_X2 U6396 ( .B1(n7887), .B2(n7876), .A(n7344), .ZN(n7523) );
  AOI21_X2 U6397 ( .B1(n9304), .B2(n9311), .A(n5104), .ZN(n9288) );
  OAI21_X2 U6398 ( .B1(n9288), .B2(n4638), .A(n4630), .ZN(n4635) );
  NAND2_X1 U6399 ( .A1(n10298), .A2(n4559), .ZN(n4558) );
  AOI21_X1 U6400 ( .B1(n7002), .B2(n7009), .A(n9783), .ZN(n7030) );
  NAND2_X1 U6401 ( .A1(n5035), .A2(n4475), .ZN(n5371) );
  NAND2_X1 U6402 ( .A1(n4947), .A2(n4950), .ZN(n7322) );
  AND2_X1 U6403 ( .A1(n6537), .A2(n6494), .ZN(n5115) );
  NAND3_X1 U6404 ( .A1(n4524), .A2(n10093), .A3(n4566), .ZN(n10215) );
  NAND2_X1 U6405 ( .A1(n10100), .A2(n10099), .ZN(n4524) );
  NAND2_X1 U6406 ( .A1(n4528), .A2(n4526), .ZN(n5797) );
  NAND2_X1 U6407 ( .A1(n5830), .A2(n4462), .ZN(n4586) );
  XNOR2_X1 U6408 ( .A(n4529), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n9125) );
  OR2_X1 U6409 ( .A1(n9117), .A2(n9116), .ZN(n4529) );
  NAND2_X1 U6410 ( .A1(n4588), .A2(n4472), .ZN(n4587) );
  NAND2_X1 U6411 ( .A1(n4614), .A2(n4613), .ZN(n9105) );
  NAND2_X1 U6412 ( .A1(n4821), .A2(n4822), .ZN(n4593) );
  NAND2_X1 U6413 ( .A1(n9128), .A2(n7537), .ZN(n4607) );
  NAND2_X1 U6414 ( .A1(n10475), .A2(n10476), .ZN(n10261) );
  NAND2_X1 U6415 ( .A1(n10259), .A2(n10260), .ZN(n10475) );
  NOR2_X1 U6416 ( .A1(n10454), .A2(n4499), .ZN(n10453) );
  NOR2_X1 U6417 ( .A1(n10277), .A2(n10468), .ZN(n10459) );
  AOI21_X1 U6418 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10448), .ZN(n10447) );
  AOI21_X1 U6419 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10445), .ZN(n10442) );
  NAND2_X1 U6420 ( .A1(n6592), .A2(n4938), .ZN(n7515) );
  NAND2_X1 U6421 ( .A1(n7619), .A2(n7620), .ZN(n7642) );
  OR2_X2 U6422 ( .A1(n8957), .A2(n8956), .ZN(n4536) );
  NAND2_X1 U6423 ( .A1(n4892), .A2(n4891), .ZN(n7618) );
  OR2_X1 U6424 ( .A1(n7584), .A2(n7585), .ZN(n7586) );
  INV_X1 U6425 ( .A(n5277), .ZN(n5013) );
  NOR2_X1 U6426 ( .A1(n6407), .A2(n6406), .ZN(n6453) );
  NAND2_X1 U6427 ( .A1(n4951), .A2(n4953), .ZN(n6539) );
  NOR2_X1 U6428 ( .A1(n10114), .A2(n10317), .ZN(n9878) );
  NOR2_X1 U6429 ( .A1(n6571), .A2(n6569), .ZN(n4595) );
  NOR2_X2 U6430 ( .A1(n6139), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n6165) );
  INV_X1 U6431 ( .A(n6935), .ZN(n4545) );
  OAI21_X1 U6432 ( .B1(n5309), .B2(n5308), .A(n5307), .ZN(n5328) );
  OAI21_X1 U6433 ( .B1(n5022), .B2(n4480), .A(n4693), .ZN(n9682) );
  INV_X1 U6434 ( .A(n5273), .ZN(n5274) );
  INV_X1 U6435 ( .A(n9508), .ZN(n9372) );
  NAND2_X1 U6436 ( .A1(n5275), .A2(n5274), .ZN(n5015) );
  NAND2_X1 U6437 ( .A1(n8846), .A2(n5061), .ZN(n9341) );
  NOR2_X4 U6438 ( .A1(n9267), .A2(n5593), .ZN(n9266) );
  NAND2_X1 U6439 ( .A1(n4750), .A2(n4749), .ZN(P2_U3548) );
  INV_X1 U6440 ( .A(n5066), .ZN(n9192) );
  NOR2_X1 U6441 ( .A1(n9451), .A2(n4752), .ZN(n4751) );
  AND2_X1 U6442 ( .A1(n5094), .A2(n6652), .ZN(n4972) );
  NAND2_X1 U6443 ( .A1(n5345), .A2(n5089), .ZN(n5035) );
  NAND2_X1 U6444 ( .A1(n10471), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n10274) );
  NAND2_X1 U6445 ( .A1(n10453), .A2(n10452), .ZN(n10451) );
  NAND2_X1 U6446 ( .A1(n4573), .A2(n4473), .ZN(n10217) );
  XNOR2_X1 U6447 ( .A(n9887), .B(n9886), .ZN(n4548) );
  NOR2_X1 U6448 ( .A1(n10456), .A2(n10455), .ZN(n10454) );
  XNOR2_X1 U6449 ( .A(n4601), .B(n6436), .ZN(n8842) );
  INV_X1 U6450 ( .A(n7663), .ZN(n4551) );
  NAND2_X1 U6451 ( .A1(n4551), .A2(n4550), .ZN(n7660) );
  NAND2_X1 U6452 ( .A1(n4556), .A2(n4555), .ZN(P2_U3516) );
  NAND2_X1 U6453 ( .A1(n9563), .A2(n10418), .ZN(n4556) );
  OAI21_X2 U6454 ( .B1(n8555), .B2(n4460), .A(n5100), .ZN(n8556) );
  INV_X1 U6455 ( .A(n5794), .ZN(n7527) );
  NAND2_X1 U6456 ( .A1(n9474), .A2(n4471), .ZN(n4572) );
  XNOR2_X2 U6457 ( .A(n4557), .B(n9154), .ZN(n9458) );
  NAND2_X1 U6458 ( .A1(n4986), .A2(n4436), .ZN(n4557) );
  NAND3_X1 U6459 ( .A1(n4578), .A2(n4579), .A3(n4577), .ZN(P1_U3260) );
  NAND2_X1 U6460 ( .A1(n7334), .A2(n7335), .ZN(n7333) );
  XNOR2_X1 U6461 ( .A(n4376), .B(P1_REG1_REG_2__SCAN_IN), .ZN(n7335) );
  OAI21_X1 U6462 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10451), .ZN(n10449) );
  OAI21_X1 U6463 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10440), .ZN(n10438) );
  OAI21_X1 U6464 ( .B1(n10427), .B2(n10258), .A(n10429), .ZN(n10473) );
  NOR2_X1 U6465 ( .A1(n10457), .A2(n4500), .ZN(n10456) );
  OAI21_X1 U6466 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n10286), .A(n10464), .ZN(
        n10288) );
  NAND2_X1 U6467 ( .A1(n8893), .A2(n8803), .ZN(n8809) );
  NAND2_X1 U6468 ( .A1(n8900), .A2(n4893), .ZN(n8964) );
  OAI21_X1 U6469 ( .B1(n8168), .B2(n8167), .A(n5113), .ZN(n8742) );
  XNOR2_X1 U6470 ( .A(n4734), .B(n5130), .ZN(n5956) );
  AND2_X1 U6471 ( .A1(n7617), .A2(n7586), .ZN(n7587) );
  NAND2_X1 U6472 ( .A1(n8798), .A2(n8797), .ZN(n4890) );
  NAND2_X2 U6473 ( .A1(n5371), .A2(n5369), .ZN(n5426) );
  NAND2_X1 U6474 ( .A1(n5216), .A2(n5217), .ZN(n5221) );
  NAND2_X1 U6475 ( .A1(n5201), .A2(n5200), .ZN(n5216) );
  INV_X1 U6476 ( .A(n4748), .ZN(n4747) );
  OAI21_X1 U6477 ( .B1(n4435), .B2(n4990), .A(n9141), .ZN(n4989) );
  INV_X1 U6478 ( .A(n4989), .ZN(n4988) );
  NAND4_X2 U6479 ( .A1(n6033), .A2(n6031), .A3(n6034), .A4(n6032), .ZN(n9780)
         );
  OAI211_X1 U6480 ( .C1(n9453), .C2(n10414), .A(n4753), .B(n4751), .ZN(n9563)
         );
  XNOR2_X1 U6481 ( .A(n10407), .B(n9033), .ZN(n7934) );
  NOR2_X1 U6482 ( .A1(n10450), .A2(n10449), .ZN(n10448) );
  NOR2_X1 U6483 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10461), .ZN(n10266) );
  AOI211_X1 U6484 ( .C1(P2_ADDR_REG_14__SCAN_IN), .C2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10281), .B(n10447), .ZN(n10445) );
  NAND2_X1 U6485 ( .A1(n7343), .A2(n7342), .ZN(n7887) );
  INV_X1 U6486 ( .A(n5536), .ZN(n5534) );
  NAND2_X1 U6487 ( .A1(n4587), .A2(n5910), .ZN(n4830) );
  AOI21_X1 U6488 ( .B1(n4593), .B2(n5903), .A(n4592), .ZN(n5906) );
  NOR2_X1 U6489 ( .A1(n4818), .A2(n5858), .ZN(n5869) );
  NAND2_X1 U6490 ( .A1(n4589), .A2(n5823), .ZN(n5829) );
  NAND3_X1 U6491 ( .A1(n5908), .A2(n5909), .A3(n5907), .ZN(n4588) );
  NAND3_X1 U6492 ( .A1(n6581), .A2(n6580), .A3(n4401), .ZN(n6582) );
  NAND2_X1 U6493 ( .A1(n4596), .A2(n4595), .ZN(P1_U3240) );
  INV_X1 U6494 ( .A(n6570), .ZN(n4596) );
  OAI21_X1 U6495 ( .B1(n4770), .B2(n6356), .A(n6412), .ZN(n4767) );
  NAND2_X1 U6496 ( .A1(n4758), .A2(n4766), .ZN(n6398) );
  NAND2_X2 U6497 ( .A1(n9978), .A2(n9977), .ZN(n9976) );
  NAND2_X1 U6498 ( .A1(n4966), .A2(n6682), .ZN(n4601) );
  NAND2_X1 U6499 ( .A1(n6644), .A2(n6643), .ZN(n7832) );
  INV_X1 U6500 ( .A(n6539), .ZN(n6537) );
  NOR2_X1 U6501 ( .A1(n6493), .A2(n4952), .ZN(n4951) );
  AOI21_X2 U6502 ( .B1(n9164), .B2(n4402), .A(n9163), .ZN(n9447) );
  NOR2_X1 U6503 ( .A1(n9105), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n9117) );
  NAND2_X1 U6504 ( .A1(n9104), .A2(n9120), .ZN(n4613) );
  INV_X1 U6505 ( .A(n9116), .ZN(n4614) );
  NAND2_X2 U6506 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5263) );
  AND2_X1 U6507 ( .A1(n5891), .A2(n5911), .ZN(n4826) );
  NAND2_X1 U6508 ( .A1(n4830), .A2(n4829), .ZN(n4828) );
  NAND2_X1 U6509 ( .A1(n4484), .A2(n4420), .ZN(n4823) );
  NAND2_X1 U6510 ( .A1(n4823), .A2(n4441), .ZN(n4822) );
  NOR2_X2 U6511 ( .A1(n5554), .A2(n5553), .ZN(n4615) );
  NAND2_X1 U6512 ( .A1(n9236), .A2(n4622), .ZN(n4620) );
  NOR2_X1 U6513 ( .A1(n9236), .A2(n9237), .ZN(n9235) );
  NAND3_X1 U6514 ( .A1(n4621), .A2(n4623), .A3(n4620), .ZN(n9467) );
  NAND3_X1 U6515 ( .A1(n4621), .A2(n4416), .A3(n4620), .ZN(n4629) );
  NAND2_X1 U6516 ( .A1(n4629), .A2(n4626), .ZN(n9566) );
  AOI21_X1 U6517 ( .B1(n9288), .B2(n9149), .A(n4638), .ZN(n9265) );
  NAND2_X1 U6518 ( .A1(n4703), .A2(n4648), .ZN(n4646) );
  OAI21_X1 U6519 ( .B1(n4703), .B2(n4650), .A(n4648), .ZN(n5526) );
  NAND2_X1 U6520 ( .A1(n4646), .A2(n4647), .ZN(n5528) );
  NAND2_X1 U6521 ( .A1(n4703), .A2(n4708), .ZN(n5469) );
  AND2_X1 U6522 ( .A1(n9107), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n4660) );
  NAND2_X1 U6523 ( .A1(n4670), .A2(n4673), .ZN(n9692) );
  NAND2_X1 U6524 ( .A1(n4379), .A2(n4674), .ZN(n4670) );
  INV_X1 U6525 ( .A(n4674), .ZN(n4672) );
  NAND2_X1 U6526 ( .A1(n6896), .A2(n4676), .ZN(n4675) );
  OAI211_X1 U6527 ( .C1(n6896), .C2(n4677), .A(n9601), .B(n4675), .ZN(P1_U3212) );
  NAND2_X1 U6528 ( .A1(n5448), .A2(n4704), .ZN(n4700) );
  NAND2_X1 U6529 ( .A1(n4700), .A2(n4701), .ZN(n5551) );
  NAND2_X1 U6530 ( .A1(n5682), .A2(n4713), .ZN(n4710) );
  NAND2_X1 U6531 ( .A1(n4710), .A2(n4711), .ZN(n5720) );
  NAND2_X1 U6532 ( .A1(n5682), .A2(n5681), .ZN(n5690) );
  NAND2_X1 U6533 ( .A1(n5734), .A2(n4492), .ZN(n4716) );
  NAND2_X1 U6534 ( .A1(n5734), .A2(n4719), .ZN(n4717) );
  OAI211_X1 U6535 ( .C1(n5734), .C2(n4718), .A(n6381), .B(n4716), .ZN(n6380)
         );
  NAND2_X1 U6536 ( .A1(n5734), .A2(n5733), .ZN(n5756) );
  OAI22_X1 U6537 ( .A1(n5576), .A2(n4487), .B1(n4419), .B2(n4728), .ZN(n5662)
         );
  XNOR2_X2 U6538 ( .A(n4733), .B(n5144), .ZN(n8847) );
  OAI21_X1 U6539 ( .B1(n4738), .B2(n7988), .A(n5812), .ZN(n4736) );
  INV_X1 U6540 ( .A(n8499), .ZN(n4737) );
  NOR2_X1 U6541 ( .A1(n7988), .A2(n4740), .ZN(n4739) );
  OR2_X1 U6542 ( .A1(n4742), .A2(n4740), .ZN(n4738) );
  OAI21_X2 U6543 ( .B1(n8549), .B2(n4747), .A(n4745), .ZN(n9409) );
  INV_X2 U6544 ( .A(n5514), .ZN(n5539) );
  NAND3_X1 U6545 ( .A1(n4765), .A2(n4764), .A3(n4759), .ZN(n4758) );
  NOR2_X1 U6546 ( .A1(n6356), .A2(n4760), .ZN(n4759) );
  NAND3_X1 U6547 ( .A1(n4765), .A2(n4764), .A3(n4762), .ZN(n4761) );
  INV_X1 U6548 ( .A(n4769), .ZN(n4768) );
  NOR2_X1 U6549 ( .A1(n6338), .A2(n9871), .ZN(n4770) );
  OAI21_X1 U6550 ( .B1(n6076), .B2(n4775), .A(n4771), .ZN(n4773) );
  INV_X1 U6551 ( .A(n7698), .ZN(n4781) );
  INV_X2 U6552 ( .A(n9780), .ZN(n7463) );
  NAND2_X1 U6553 ( .A1(n6244), .A2(n4786), .ZN(n4782) );
  AOI21_X1 U6554 ( .B1(n6244), .B2(n4481), .A(n4783), .ZN(n6284) );
  NOR2_X1 U6555 ( .A1(n5971), .A2(P1_IR_REG_28__SCAN_IN), .ZN(n4794) );
  OR2_X1 U6556 ( .A1(n6185), .A2(n4801), .ZN(n4800) );
  AND2_X1 U6557 ( .A1(n4805), .A2(n4802), .ZN(n4801) );
  INV_X1 U6558 ( .A(n4808), .ZN(n5184) );
  AND2_X1 U6559 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n5184), .ZN(n5156) );
  OR2_X1 U6560 ( .A1(n7782), .A2(n4809), .ZN(n5799) );
  AOI21_X1 U6561 ( .B1(n4813), .B2(n5805), .A(n5877), .ZN(n4812) );
  NAND2_X1 U6562 ( .A1(n4814), .A2(n5783), .ZN(n4813) );
  NAND2_X1 U6563 ( .A1(n5797), .A2(n5780), .ZN(n4814) );
  NOR2_X1 U6564 ( .A1(n5848), .A2(n4820), .ZN(n4818) );
  INV_X1 U6565 ( .A(n4819), .ZN(n5873) );
  INV_X1 U6566 ( .A(n5859), .ZN(n4820) );
  AND2_X1 U6567 ( .A1(n4448), .A2(n5127), .ZN(n4832) );
  NAND4_X1 U6568 ( .A1(n5948), .A2(n5129), .A3(n5128), .A4(n4831), .ZN(n9584)
         );
  AND4_X1 U6569 ( .A1(n5129), .A2(n5128), .A3(n5948), .A4(n4832), .ZN(n5134)
         );
  NAND2_X1 U6570 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n4838) );
  INV_X1 U6571 ( .A(n9791), .ZN(n4851) );
  INV_X1 U6572 ( .A(n4867), .ZN(n8696) );
  OAI21_X1 U6573 ( .B1(P1_REG2_REG_4__SCAN_IN), .B2(n9789), .A(n9790), .ZN(
        n7027) );
  NOR2_X1 U6574 ( .A1(n9811), .A2(n9810), .ZN(n9809) );
  NOR2_X1 U6575 ( .A1(n8700), .A2(n9803), .ZN(n9811) );
  OAI21_X1 U6576 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n7719), .A(n7718), .ZN(
        n7721) );
  OAI21_X1 U6577 ( .B1(n7177), .B2(P1_REG2_REG_8__SCAN_IN), .A(n7176), .ZN(
        n7179) );
  XNOR2_X1 U6578 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n8705), .ZN(n8716) );
  NAND2_X1 U6579 ( .A1(n7077), .A2(n7076), .ZN(n7078) );
  OAI21_X1 U6580 ( .B1(n4552), .B2(n4875), .A(n4873), .ZN(n7913) );
  NAND2_X1 U6581 ( .A1(n4872), .A2(n4870), .ZN(n7918) );
  NAND2_X1 U6582 ( .A1(n7643), .A2(n4873), .ZN(n4872) );
  NAND3_X1 U6583 ( .A1(n8809), .A2(n4882), .A3(n8808), .ZN(n4878) );
  NAND2_X1 U6584 ( .A1(n4878), .A2(n4880), .ZN(n8824) );
  NAND3_X1 U6585 ( .A1(n8809), .A2(n8808), .A3(n4440), .ZN(n4879) );
  NAND3_X1 U6586 ( .A1(n8809), .A2(n8808), .A3(n4886), .ZN(n4885) );
  AND2_X1 U6587 ( .A1(n7587), .A2(n7582), .ZN(n4891) );
  NAND2_X1 U6588 ( .A1(n8964), .A2(n8774), .ZN(n8775) );
  INV_X2 U6589 ( .A(n8788), .ZN(n8819) );
  NAND2_X1 U6590 ( .A1(n5949), .A2(n4898), .ZN(n5766) );
  INV_X1 U6591 ( .A(n9123), .ZN(n9127) );
  NAND2_X1 U6592 ( .A1(n4927), .A2(n4928), .ZN(n9892) );
  AND2_X1 U6593 ( .A1(n7812), .A2(n7809), .ZN(n6590) );
  INV_X1 U6594 ( .A(n9862), .ZN(n4944) );
  INV_X1 U6595 ( .A(n6624), .ZN(n4945) );
  NAND2_X1 U6596 ( .A1(n6660), .A2(n6659), .ZN(n10018) );
  INV_X1 U6597 ( .A(n6659), .ZN(n4959) );
  INV_X1 U6598 ( .A(n4960), .ZN(n9978) );
  NAND2_X1 U6599 ( .A1(n9870), .A2(n6681), .ZN(n4966) );
  NAND2_X1 U6600 ( .A1(n9976), .A2(n4971), .ZN(n4970) );
  NAND2_X1 U6601 ( .A1(n4970), .A2(n4477), .ZN(n6674) );
  CLKBUF_X1 U6602 ( .A(n4970), .Z(n4967) );
  NAND2_X1 U6603 ( .A1(n4973), .A2(n4972), .ZN(n8600) );
  INV_X1 U6604 ( .A(n7848), .ZN(n7903) );
  AND2_X1 U6605 ( .A1(n7788), .A2(n5928), .ZN(n4987) );
  NAND2_X1 U6606 ( .A1(n9372), .A2(n9387), .ZN(n5001) );
  NAND2_X1 U6607 ( .A1(n6839), .A2(n5009), .ZN(n5005) );
  NAND2_X1 U6608 ( .A1(n5015), .A2(n5277), .ZN(n5291) );
  NAND2_X1 U6609 ( .A1(n5469), .A2(n5468), .ZN(n5486) );
  NAND2_X1 U6610 ( .A1(n9250), .A2(n5032), .ZN(n5031) );
  NAND2_X1 U6611 ( .A1(n5031), .A2(n5029), .ZN(n9229) );
  NAND2_X1 U6612 ( .A1(n5035), .A2(n5346), .ZN(n5360) );
  NOR2_X1 U6613 ( .A1(n5971), .A2(n5041), .ZN(n5040) );
  NAND2_X1 U6614 ( .A1(n4798), .A2(n5040), .ZN(n6521) );
  NOR2_X1 U6615 ( .A1(n7819), .A2(n5047), .ZN(n5046) );
  INV_X1 U6616 ( .A(n9906), .ZN(n5049) );
  NAND2_X1 U6617 ( .A1(n5050), .A2(n5049), .ZN(n9849) );
  AND2_X2 U6618 ( .A1(n9266), .A2(n5056), .ZN(n9222) );
  NOR3_X1 U6619 ( .A1(n9398), .A2(n9416), .A3(n9522), .ZN(n9396) );
  OR2_X2 U6620 ( .A1(n9212), .A2(n5064), .ZN(n9167) );
  NAND3_X1 U6621 ( .A1(n4409), .A2(n7980), .A3(n8723), .ZN(n8845) );
  NAND3_X1 U6622 ( .A1(n8131), .A2(n7980), .A3(n5068), .ZN(n5112) );
  OAI21_X2 U6623 ( .B1(n8077), .B2(n4468), .A(n5072), .ZN(n8549) );
  INV_X1 U6624 ( .A(n8551), .ZN(n5077) );
  NAND2_X1 U6625 ( .A1(n5079), .A2(n5078), .ZN(n7976) );
  OAI21_X1 U6626 ( .B1(n9178), .B2(n5083), .A(n5080), .ZN(n5762) );
  NAND2_X1 U6627 ( .A1(n5087), .A2(n5914), .ZN(n5086) );
  CLKBUF_X1 U6628 ( .A(n6520), .Z(n7419) );
  INV_X1 U6629 ( .A(n6727), .ZN(n6728) );
  NAND2_X1 U6630 ( .A1(n5652), .A2(n5650), .ZN(n5632) );
  INV_X1 U6631 ( .A(n7707), .ZN(n6698) );
  XNOR2_X1 U6632 ( .A(n6731), .B(n6732), .ZN(n7305) );
  NAND2_X1 U6633 ( .A1(n6697), .A2(n10333), .ZN(n7707) );
  INV_X1 U6634 ( .A(n5989), .ZN(n5986) );
  CLKBUF_X1 U6635 ( .A(n5989), .Z(n8861) );
  OR2_X1 U6636 ( .A1(n5244), .A2(n7668), .ZN(n5174) );
  OAI211_X1 U6637 ( .C1(n10344), .C2(n6705), .A(n4438), .B(n10090), .ZN(n10091) );
  INV_X1 U6638 ( .A(n7708), .ZN(n6697) );
  NAND2_X1 U6639 ( .A1(n7318), .A2(n5070), .ZN(n7568) );
  NAND2_X1 U6640 ( .A1(n6701), .A2(n9992), .ZN(n10315) );
  AND2_X1 U6641 ( .A1(n5346), .A2(n5334), .ZN(n5089) );
  OR2_X1 U6642 ( .A1(n7567), .A2(n7566), .ZN(n5091) );
  OR2_X1 U6643 ( .A1(n9942), .A2(n6857), .ZN(n5092) );
  NOR2_X1 U6644 ( .A1(n6792), .A2(n8537), .ZN(n5093) );
  NOR2_X1 U6645 ( .A1(n8596), .A2(n6653), .ZN(n5094) );
  NAND2_X1 U6646 ( .A1(n6536), .A2(n7444), .ZN(n7446) );
  AND2_X1 U6647 ( .A1(n5424), .A2(n5423), .ZN(n5095) );
  OR3_X1 U6648 ( .A1(n7590), .A2(n7589), .A3(n10408), .ZN(n7677) );
  AND2_X1 U6649 ( .A1(n5585), .A2(n5555), .ZN(n5096) );
  AND2_X1 U6650 ( .A1(n5152), .A2(n5151), .ZN(n5097) );
  AND2_X1 U6651 ( .A1(n5468), .A2(n5452), .ZN(n5098) );
  OR2_X1 U6652 ( .A1(n6226), .A2(n10013), .ZN(n5099) );
  AND2_X1 U6653 ( .A1(n5329), .A2(n5314), .ZN(n5102) );
  AND2_X1 U6654 ( .A1(n5503), .A2(n5529), .ZN(n5504) );
  AND2_X1 U6655 ( .A1(n9489), .A2(n9332), .ZN(n5104) );
  OR3_X1 U6656 ( .A1(n6402), .A2(n7368), .A3(n6512), .ZN(n5105) );
  NAND2_X1 U6657 ( .A1(n9440), .A2(n10399), .ZN(n5106) );
  OR2_X1 U6658 ( .A1(n5805), .A2(n5911), .ZN(n5107) );
  OR2_X1 U6659 ( .A1(n5732), .A2(SI_29_), .ZN(n5108) );
  AND3_X1 U6660 ( .A1(n6515), .A2(n6555), .A3(n6514), .ZN(n5109) );
  AND4_X1 U6661 ( .A1(n10097), .A2(n6436), .A3(n6435), .A4(n6434), .ZN(n5110)
         );
  AND2_X1 U6662 ( .A1(n7934), .A2(n5107), .ZN(n5111) );
  AND2_X1 U6663 ( .A1(n8166), .A2(n8165), .ZN(n5113) );
  INV_X1 U6664 ( .A(n5819), .ZN(n5827) );
  AND2_X1 U6665 ( .A1(n7046), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5114) );
  INV_X1 U6666 ( .A(n7447), .ZN(n7444) );
  NAND2_X1 U6667 ( .A1(n7305), .A2(n7306), .ZN(n7304) );
  NOR4_X1 U6668 ( .A1(n6138), .A2(n6137), .A3(n8596), .A4(n6136), .ZN(n6148)
         );
  INV_X1 U6669 ( .A(n9329), .ZN(n5856) );
  NAND2_X1 U6670 ( .A1(n5919), .A2(n5864), .ZN(n5865) );
  OAI21_X1 U6671 ( .B1(n5919), .B2(n5877), .A(n5865), .ZN(n5866) );
  AOI21_X1 U6672 ( .B1(n6228), .B2(n6227), .A(n5099), .ZN(n6244) );
  NAND2_X1 U6673 ( .A1(n5886), .A2(n5877), .ZN(n5887) );
  NAND2_X1 U6674 ( .A1(n5893), .A2(n5911), .ZN(n5894) );
  INV_X1 U6675 ( .A(n5419), .ZN(n5420) );
  NOR2_X1 U6676 ( .A1(n7527), .A2(n8065), .ZN(n7345) );
  AND2_X1 U6677 ( .A1(n5649), .A2(n5648), .ZN(n5653) );
  OAI21_X1 U6678 ( .B1(n8952), .B2(n9251), .A(n8892), .ZN(n8802) );
  AND2_X1 U6679 ( .A1(n6725), .A2(P1_IR_REG_0__SCAN_IN), .ZN(n6726) );
  INV_X1 U6680 ( .A(n9776), .ZN(n6591) );
  OR2_X1 U6681 ( .A1(n5655), .A2(n5654), .ZN(n5657) );
  NOR2_X1 U6682 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n6018) );
  INV_X1 U6683 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n5293) );
  INV_X1 U6684 ( .A(n7888), .ZN(n5163) );
  AOI21_X1 U6685 ( .B1(n6800), .B2(n7422), .A(n6726), .ZN(n6727) );
  OAI211_X1 U6686 ( .C1(n7368), .C2(n6558), .A(n5105), .B(n6400), .ZN(n6401)
         );
  AND2_X1 U6687 ( .A1(n5633), .A2(n5631), .ZN(n5654) );
  NAND2_X1 U6688 ( .A1(n6023), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6409) );
  AND2_X1 U6689 ( .A1(n8889), .A2(n8739), .ZN(n8740) );
  AND2_X1 U6690 ( .A1(n8902), .A2(n8764), .ZN(n8765) );
  NAND2_X1 U6691 ( .A1(n8952), .A2(n8806), .ZN(n8807) );
  OR2_X1 U6692 ( .A1(n8681), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n8682) );
  AND2_X1 U6694 ( .A1(n7542), .A2(n7541), .ZN(n7867) );
  INV_X1 U6695 ( .A(n8556), .ZN(n8558) );
  INV_X1 U6696 ( .A(n5488), .ZN(n5489) );
  INV_X1 U6697 ( .A(n6877), .ZN(n6876) );
  AOI21_X1 U6698 ( .B1(n8105), .B2(n8108), .A(n8107), .ZN(n8524) );
  NAND2_X1 U6699 ( .A1(n9900), .A2(n10057), .ZN(n9874) );
  AND2_X1 U6700 ( .A1(n10164), .A2(n10038), .ZN(n6613) );
  OR2_X1 U6701 ( .A1(n6928), .A2(n6949), .ZN(n6926) );
  NAND2_X1 U6702 ( .A1(n5387), .A2(n8399), .ZN(n5419) );
  NAND2_X1 U6703 ( .A1(n5332), .A2(n5331), .ZN(n5346) );
  INV_X1 U6704 ( .A(n9332), .ZN(n8918) );
  OR2_X1 U6705 ( .A1(n8999), .A2(n9384), .ZN(n8992) );
  OR2_X1 U6706 ( .A1(n7590), .A2(n4896), .ZN(n8999) );
  INV_X1 U6707 ( .A(n7757), .ZN(n5955) );
  INV_X1 U6708 ( .A(n9195), .ZN(n9154) );
  NOR2_X1 U6709 ( .A1(n9606), .A2(n9605), .ZN(n9662) );
  INV_X1 U6710 ( .A(n6859), .ZN(n6860) );
  OR2_X1 U6711 ( .A1(n6909), .A2(n7194), .ZN(n6927) );
  INV_X1 U6712 ( .A(n9770), .ZN(n9706) );
  OR2_X1 U6713 ( .A1(n6924), .A2(n7323), .ZN(n9758) );
  OR2_X1 U6714 ( .A1(n9650), .A2(n6371), .ZN(n6324) );
  INV_X1 U6715 ( .A(n10107), .ZN(n8837) );
  INV_X1 U6716 ( .A(n10126), .ZN(n9910) );
  NOR2_X1 U6717 ( .A1(n10148), .A2(n9988), .ZN(n6614) );
  NAND2_X1 U6718 ( .A1(n10095), .A2(n10134), .ZN(n10096) );
  AND2_X1 U6719 ( .A1(n7375), .A2(n7374), .ZN(n10040) );
  INV_X1 U6720 ( .A(n9017), .ZN(n8990) );
  AND2_X1 U6721 ( .A1(n5728), .A2(n5727), .ZN(n8826) );
  AND2_X1 U6722 ( .A1(n5549), .A2(n5548), .ZN(n9349) );
  AND2_X1 U6723 ( .A1(n7156), .A2(n7155), .ZN(n10366) );
  INV_X1 U6724 ( .A(n9124), .ZN(n10361) );
  INV_X1 U6725 ( .A(n9386), .ZN(n9412) );
  AND2_X1 U6726 ( .A1(n9383), .A2(n9382), .ZN(n9511) );
  INV_X1 U6727 ( .A(n9427), .ZN(n9421) );
  NAND2_X1 U6728 ( .A1(n9427), .A2(n7883), .ZN(n9371) );
  INV_X1 U6729 ( .A(n9371), .ZN(n9422) );
  AOI21_X1 U6730 ( .B1(n10371), .B2(n10381), .A(n10382), .ZN(n7870) );
  OR2_X1 U6731 ( .A1(n9446), .A2(n5106), .ZN(n9449) );
  AND2_X1 U6732 ( .A1(n8186), .A2(n8185), .ZN(n9539) );
  NAND2_X1 U6733 ( .A1(n8560), .A2(n9556), .ZN(n10399) );
  AND2_X1 U6734 ( .A1(n7548), .A2(n10385), .ZN(n10373) );
  INV_X1 U6735 ( .A(n6390), .ZN(n6388) );
  AND3_X1 U6736 ( .A1(n6242), .A2(n6241), .A3(n6240), .ZN(n6714) );
  AND2_X1 U6737 ( .A1(n7014), .A2(n6981), .ZN(n10302) );
  NAND2_X1 U6738 ( .A1(n9869), .A2(n6679), .ZN(n9886) );
  NAND2_X1 U6739 ( .A1(n6468), .A2(n9912), .ZN(n9947) );
  AND2_X1 U6740 ( .A1(n10315), .A2(n7421), .ZN(n10052) );
  OR3_X1 U6741 ( .A1(n10334), .A2(n9962), .A3(n6946), .ZN(n9992) );
  OR2_X1 U6742 ( .A1(n7368), .A2(n7367), .ZN(n10211) );
  AND2_X1 U6743 ( .A1(n7193), .A2(n7192), .ZN(n7211) );
  AND2_X1 U6744 ( .A1(n5998), .A2(n5997), .ZN(n7409) );
  XNOR2_X1 U6745 ( .A(n6010), .B(P1_IR_REG_8__SCAN_IN), .ZN(n7177) );
  INV_X1 U6746 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n10256) );
  INV_X1 U6747 ( .A(n9131), .ZN(n10358) );
  INV_X1 U6748 ( .A(n9019), .ZN(n8996) );
  INV_X1 U6749 ( .A(n9243), .ZN(n9026) );
  INV_X1 U6750 ( .A(n8916), .ZN(n9299) );
  INV_X1 U6751 ( .A(n10362), .ZN(n9101) );
  AND2_X1 U6752 ( .A1(n8615), .A2(n8614), .ZN(n9529) );
  AND2_X1 U6753 ( .A1(n7871), .A2(n9373), .ZN(n9404) );
  INV_X1 U6754 ( .A(n10426), .ZN(n10424) );
  INV_X1 U6755 ( .A(n10418), .ZN(n10416) );
  NAND2_X1 U6756 ( .A1(n10373), .A2(n10372), .ZN(n10383) );
  INV_X1 U6757 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n7117) );
  INV_X1 U6758 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n8236) );
  INV_X1 U6759 ( .A(n9734), .ZN(n9760) );
  INV_X1 U6760 ( .A(n8526), .ZN(n9765) );
  INV_X1 U6761 ( .A(n9745), .ZN(n9873) );
  INV_X1 U6762 ( .A(n6714), .ZN(n10004) );
  INV_X1 U6763 ( .A(n6437), .ZN(n10086) );
  INV_X1 U6764 ( .A(n10357), .ZN(n10355) );
  OR3_X1 U6765 ( .A1(n10194), .A2(n10193), .A3(n10192), .ZN(n10233) );
  XNOR2_X1 U6766 ( .A(n6527), .B(n6526), .ZN(n8133) );
  INV_X1 U6767 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n7119) );
  INV_X1 U6768 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n8414) );
  XNOR2_X1 U6769 ( .A(n6088), .B(n6087), .ZN(n7037) );
  NOR2_X1 U6770 ( .A1(n10470), .A2(n10469), .ZN(n10468) );
  NOR2_X1 U6771 ( .A1(n10459), .A2(n10458), .ZN(n10457) );
  INV_X1 U6772 ( .A(n9037), .ZN(P2_U3966) );
  INV_X1 U6773 ( .A(n9778), .ZN(P1_U4006) );
  OAI21_X1 U6774 ( .B1(n6712), .B2(n10074), .A(n6711), .ZN(P1_U3355) );
  NOR2_X1 U6775 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .ZN(
        n5117) );
  INV_X1 U6776 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5116) );
  NAND3_X1 U6777 ( .A1(n5749), .A2(n5117), .A3(n5116), .ZN(n5119) );
  INV_X2 U6778 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5769) );
  NAND4_X1 U6779 ( .A1(n5458), .A2(n5477), .A3(n5533), .A4(n5769), .ZN(n5118)
         );
  NOR2_X2 U6780 ( .A1(n5119), .A2(n5118), .ZN(n5948) );
  INV_X1 U6781 ( .A(n5298), .ZN(n5129) );
  NOR2_X1 U6782 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n5126) );
  NAND4_X1 U6783 ( .A1(n5126), .A2(n5125), .A3(n5124), .A4(n5123), .ZN(n5453)
         );
  INV_X1 U6784 ( .A(n5453), .ZN(n5128) );
  INV_X1 U6785 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5131) );
  NAND2_X1 U6786 ( .A1(n5225), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5142) );
  INV_X1 U6787 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n8248) );
  NAND2_X1 U6788 ( .A1(n8857), .A2(n8693), .ZN(n5227) );
  INV_X1 U6789 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n5137) );
  OR2_X1 U6790 ( .A1(n5227), .A2(n5137), .ZN(n5140) );
  INV_X1 U6791 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n7163) );
  INV_X1 U6792 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5144) );
  NAND2_X2 U6793 ( .A1(n5207), .A2(n6964), .ZN(n5581) );
  NAND2_X1 U6794 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5146) );
  INV_X1 U6795 ( .A(SI_1_), .ZN(n5178) );
  NAND2_X1 U6796 ( .A1(n5146), .A2(n5178), .ZN(n5145) );
  NAND2_X1 U6797 ( .A1(n5145), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n5149) );
  INV_X1 U6798 ( .A(n5146), .ZN(n5147) );
  NAND2_X1 U6799 ( .A1(n5147), .A2(SI_1_), .ZN(n5148) );
  NAND2_X1 U6800 ( .A1(n5149), .A2(n5148), .ZN(n5150) );
  NAND2_X1 U6801 ( .A1(n5470), .A2(n5150), .ZN(n5153) );
  OAI211_X1 U6802 ( .C1(SI_1_), .C2(P1_DATAO_REG_1__SCAN_IN), .A(SI_0_), .B(
        P1_DATAO_REG_0__SCAN_IN), .ZN(n5152) );
  NAND2_X1 U6803 ( .A1(SI_1_), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5151) );
  INV_X1 U6804 ( .A(SI_2_), .ZN(n5195) );
  XNOR2_X1 U6805 ( .A(n5197), .B(n5195), .ZN(n5155) );
  MUX2_X1 U6806 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .S(n4398), .Z(n5154) );
  XNOR2_X1 U6807 ( .A(n5155), .B(n5154), .ZN(n6988) );
  OR2_X1 U6808 ( .A1(n5581), .A2(n6988), .ZN(n5162) );
  NAND2_X4 U6809 ( .A1(n5207), .A2(n4399), .ZN(n5514) );
  INV_X1 U6810 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6987) );
  OR2_X1 U6811 ( .A1(n5514), .A2(n6987), .ZN(n5161) );
  NAND2_X1 U6812 ( .A1(n5156), .A2(P2_IR_REG_2__SCAN_IN), .ZN(n5159) );
  OR2_X1 U6813 ( .A1(n7154), .A2(n7223), .ZN(n5160) );
  AND3_X2 U6814 ( .A1(n5162), .A2(n5161), .A3(n5160), .ZN(n7888) );
  NAND2_X1 U6815 ( .A1(n9036), .A2(n7888), .ZN(n5788) );
  NAND2_X1 U6816 ( .A1(n5788), .A2(n5790), .ZN(n5924) );
  INV_X1 U6817 ( .A(n5924), .ZN(n7876) );
  NAND2_X1 U6818 ( .A1(n5225), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5170) );
  INV_X1 U6819 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n8025) );
  OR2_X1 U6820 ( .A1(n4395), .A2(n8025), .ZN(n5169) );
  INV_X1 U6821 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n5165) );
  OR2_X1 U6822 ( .A1(n5227), .A2(n5165), .ZN(n5168) );
  INV_X1 U6823 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n5166) );
  INV_X1 U6824 ( .A(n10367), .ZN(n10359) );
  NAND2_X1 U6825 ( .A1(n6964), .A2(SI_0_), .ZN(n5172) );
  INV_X1 U6826 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5171) );
  XNOR2_X1 U6827 ( .A(n5172), .B(n5171), .ZN(n9592) );
  INV_X1 U6828 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n7164) );
  INV_X1 U6829 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n5173) );
  OR2_X1 U6830 ( .A1(n5227), .A2(n5173), .ZN(n5176) );
  NAND2_X1 U6831 ( .A1(n5225), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5175) );
  INV_X1 U6832 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n7668) );
  INV_X1 U6833 ( .A(n7141), .ZN(n5188) );
  MUX2_X1 U6834 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n5470), .Z(n5179) );
  XNOR2_X1 U6835 ( .A(n5179), .B(n5178), .ZN(n5182) );
  MUX2_X1 U6836 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(P2_DATAO_REG_0__SCAN_IN), 
        .S(n4398), .Z(n5180) );
  NAND2_X1 U6837 ( .A1(n5180), .A2(SI_0_), .ZN(n5181) );
  XNOR2_X1 U6838 ( .A(n5182), .B(n5181), .ZN(n6036) );
  NAND2_X1 U6839 ( .A1(n5183), .A2(n6036), .ZN(n5187) );
  INV_X1 U6840 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6986) );
  OR2_X1 U6841 ( .A1(n5207), .A2(n7204), .ZN(n5185) );
  NAND2_X1 U6842 ( .A1(n7876), .A2(n7877), .ZN(n7875) );
  NAND2_X1 U6843 ( .A1(n7875), .A2(n5790), .ZN(n7526) );
  NAND2_X1 U6844 ( .A1(n5225), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5194) );
  INV_X1 U6845 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n5190) );
  OR2_X1 U6846 ( .A1(n5285), .A2(n5190), .ZN(n5193) );
  INV_X1 U6847 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n7224) );
  OR2_X1 U6848 ( .A1(n5260), .A2(n7224), .ZN(n5192) );
  OR2_X1 U6849 ( .A1(n4394), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5191) );
  NAND4_X2 U6850 ( .A1(n5194), .A2(n5193), .A3(n5192), .A4(n5191), .ZN(n7346)
         );
  NAND2_X1 U6851 ( .A1(n5470), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5196) );
  NAND2_X1 U6852 ( .A1(n5198), .A2(n5197), .ZN(n5201) );
  NAND2_X1 U6853 ( .A1(n5470), .A2(n6958), .ZN(n5199) );
  OAI211_X1 U6854 ( .C1(n5470), .C2(P1_DATAO_REG_2__SCAN_IN), .A(n5199), .B(
        SI_2_), .ZN(n5200) );
  XNOR2_X1 U6855 ( .A(n5218), .B(SI_3_), .ZN(n5217) );
  INV_X1 U6856 ( .A(n5217), .ZN(n5202) );
  XNOR2_X1 U6857 ( .A(n5216), .B(n5202), .ZN(n6059) );
  NAND2_X1 U6858 ( .A1(n5635), .A2(n6059), .ZN(n5206) );
  NAND2_X1 U6859 ( .A1(n5208), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5203) );
  OR2_X1 U6860 ( .A1(n7154), .A2(n7253), .ZN(n5205) );
  OR2_X1 U6861 ( .A1(n5514), .A2(n6968), .ZN(n5204) );
  AND3_X2 U6862 ( .A1(n5206), .A2(n5205), .A3(n5204), .ZN(n8491) );
  OR2_X1 U6863 ( .A1(n7346), .A2(n8491), .ZN(n8064) );
  NAND2_X1 U6864 ( .A1(n7346), .A2(n8491), .ZN(n5798) );
  NAND2_X1 U6865 ( .A1(n8064), .A2(n5798), .ZN(n5794) );
  NAND2_X1 U6866 ( .A1(n7526), .A2(n7527), .ZN(n7525) );
  INV_X1 U6867 ( .A(n5208), .ZN(n5210) );
  INV_X1 U6868 ( .A(n5214), .ZN(n5211) );
  NAND2_X1 U6869 ( .A1(n5211), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5212) );
  MUX2_X1 U6870 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5212), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n5215) );
  INV_X1 U6871 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5213) );
  NAND2_X1 U6872 ( .A1(n5214), .A2(n5213), .ZN(n5241) );
  NAND2_X1 U6873 ( .A1(n5215), .A2(n5241), .ZN(n7281) );
  INV_X1 U6874 ( .A(n7281), .ZN(n7229) );
  AOI22_X1 U6875 ( .A1(n5539), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n4375), .B2(
        n7229), .ZN(n5224) );
  INV_X1 U6876 ( .A(n5218), .ZN(n5219) );
  NAND2_X1 U6877 ( .A1(n5219), .A2(SI_3_), .ZN(n5220) );
  NAND2_X1 U6878 ( .A1(n5221), .A2(n5220), .ZN(n5235) );
  MUX2_X1 U6879 ( .A(n6971), .B(n6943), .S(n5470), .Z(n5236) );
  XNOR2_X1 U6880 ( .A(n5236), .B(SI_4_), .ZN(n5234) );
  INV_X1 U6881 ( .A(n5234), .ZN(n5222) );
  XNOR2_X1 U6882 ( .A(n5235), .B(n5222), .ZN(n6073) );
  NAND2_X1 U6883 ( .A1(n6073), .A2(n5635), .ZN(n5223) );
  AND2_X2 U6884 ( .A1(n5224), .A2(n5223), .ZN(n10394) );
  INV_X1 U6885 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n7217) );
  OAI21_X1 U6886 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(P2_REG3_REG_4__SCAN_IN), 
        .A(n5263), .ZN(n8061) );
  OR2_X1 U6887 ( .A1(n4394), .A2(n8061), .ZN(n5229) );
  INV_X1 U6888 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n5226) );
  OR2_X1 U6889 ( .A1(n5227), .A2(n5226), .ZN(n5228) );
  INV_X1 U6890 ( .A(n8065), .ZN(n5232) );
  INV_X1 U6891 ( .A(n8064), .ZN(n5781) );
  NOR2_X1 U6892 ( .A1(n5232), .A2(n5781), .ZN(n5233) );
  NAND2_X1 U6893 ( .A1(n7525), .A2(n5233), .ZN(n7351) );
  NAND2_X1 U6894 ( .A1(n5235), .A2(n5234), .ZN(n5239) );
  INV_X1 U6895 ( .A(n5236), .ZN(n5237) );
  NAND2_X1 U6896 ( .A1(n5237), .A2(SI_4_), .ZN(n5238) );
  MUX2_X1 U6897 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n5470), .Z(n5254) );
  XNOR2_X1 U6898 ( .A(n5253), .B(n5251), .ZN(n6089) );
  NAND2_X1 U6899 ( .A1(n6089), .A2(n5635), .ZN(n5243) );
  NAND2_X1 U6900 ( .A1(n5241), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5240) );
  MUX2_X1 U6901 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5240), .S(
        P2_IR_REG_5__SCAN_IN), .Z(n5242) );
  NAND2_X1 U6902 ( .A1(n5225), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5249) );
  INV_X1 U6903 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n8088) );
  OR2_X1 U6904 ( .A1(n5260), .A2(n8088), .ZN(n5248) );
  INV_X1 U6905 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5262) );
  XNOR2_X1 U6906 ( .A(n5263), .B(n5262), .ZN(n8086) );
  OR2_X1 U6907 ( .A1(n4394), .A2(n8086), .ZN(n5247) );
  INV_X1 U6908 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n5245) );
  OR2_X1 U6909 ( .A1(n5285), .A2(n5245), .ZN(n5246) );
  AND2_X2 U6910 ( .A1(n5780), .A2(n5799), .ZN(n7785) );
  AND2_X1 U6911 ( .A1(n7350), .A2(n7785), .ZN(n5250) );
  NAND2_X1 U6912 ( .A1(n7351), .A2(n5250), .ZN(n7355) );
  NAND2_X1 U6913 ( .A1(n5253), .A2(n5252), .ZN(n5256) );
  NAND2_X1 U6914 ( .A1(n5254), .A2(SI_5_), .ZN(n5255) );
  XNOR2_X1 U6915 ( .A(n5275), .B(n5273), .ZN(n6099) );
  NAND2_X1 U6916 ( .A1(n6099), .A2(n5635), .ZN(n5259) );
  NAND2_X1 U6917 ( .A1(n5278), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5257) );
  AOI22_X1 U6918 ( .A1(n5539), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n4375), .B2(
        n7260), .ZN(n5258) );
  NAND2_X1 U6919 ( .A1(n5225), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5271) );
  INV_X1 U6920 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7232) );
  OR2_X1 U6921 ( .A1(n5260), .A2(n7232), .ZN(n5270) );
  INV_X1 U6922 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n5261) );
  OAI21_X1 U6923 ( .B1(n5263), .B2(n5262), .A(n5261), .ZN(n5266) );
  NAND2_X1 U6924 ( .A1(n5266), .A2(n5283), .ZN(n7646) );
  OR2_X1 U6925 ( .A1(n4395), .A2(n7646), .ZN(n5269) );
  INV_X1 U6926 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n5267) );
  OR2_X1 U6927 ( .A1(n5285), .A2(n5267), .ZN(n5268) );
  NOR2_X2 U6928 ( .A1(n8506), .A2(n7671), .ZN(n5803) );
  INV_X1 U6929 ( .A(n5803), .ZN(n5272) );
  NAND2_X2 U6930 ( .A1(n5272), .A2(n5805), .ZN(n8509) );
  INV_X1 U6931 ( .A(n8509), .ZN(n8511) );
  NAND2_X1 U6932 ( .A1(n5276), .A2(SI_6_), .ZN(n5277) );
  NAND2_X1 U6933 ( .A1(n6962), .A2(n5635), .ZN(n5281) );
  OAI21_X1 U6934 ( .B1(n5278), .B2(P2_IR_REG_6__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5279) );
  XNOR2_X1 U6935 ( .A(n5279), .B(P2_IR_REG_7__SCAN_IN), .ZN(n7387) );
  AOI22_X1 U6936 ( .A1(n5539), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n4375), .B2(
        n7387), .ZN(n5280) );
  NAND2_X1 U6937 ( .A1(n5225), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5289) );
  INV_X1 U6938 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n7938) );
  OR2_X1 U6939 ( .A1(n5260), .A2(n7938), .ZN(n5288) );
  INV_X1 U6940 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n8444) );
  NAND2_X1 U6941 ( .A1(n5283), .A2(n8444), .ZN(n5284) );
  NAND2_X1 U6942 ( .A1(n5321), .A2(n5284), .ZN(n7941) );
  OR2_X1 U6943 ( .A1(n4395), .A2(n7941), .ZN(n5287) );
  OR2_X1 U6944 ( .A1(n5285), .A2(n10417), .ZN(n5286) );
  NAND4_X1 U6945 ( .A1(n5289), .A2(n5288), .A3(n5287), .A4(n5286), .ZN(n9033)
         );
  INV_X1 U6946 ( .A(n7934), .ZN(n5928) );
  INV_X1 U6947 ( .A(n9033), .ZN(n7987) );
  MUX2_X1 U6948 ( .A(n8236), .B(n5293), .S(n4399), .Z(n5295) );
  INV_X1 U6949 ( .A(SI_8_), .ZN(n5294) );
  INV_X1 U6950 ( .A(n5295), .ZN(n5296) );
  NAND2_X1 U6951 ( .A1(n5296), .A2(SI_8_), .ZN(n5297) );
  XNOR2_X1 U6952 ( .A(n5309), .B(n5308), .ZN(n6960) );
  NAND2_X1 U6953 ( .A1(n6960), .A2(n5635), .ZN(n5302) );
  NAND2_X1 U6954 ( .A1(n5454), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5299) );
  MUX2_X1 U6955 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5299), .S(
        P2_IR_REG_8__SCAN_IN), .Z(n5300) );
  AND2_X1 U6956 ( .A1(n5300), .A2(n5335), .ZN(n7494) );
  AOI22_X1 U6957 ( .A1(n5539), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n4375), .B2(
        n7494), .ZN(n5301) );
  NAND2_X1 U6958 ( .A1(n5225), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5306) );
  INV_X1 U6959 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7995) );
  OR2_X1 U6960 ( .A1(n5260), .A2(n7995), .ZN(n5305) );
  INV_X1 U6961 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n5319) );
  XNOR2_X1 U6962 ( .A(n5321), .B(n5319), .ZN(n7998) );
  OR2_X1 U6963 ( .A1(n4394), .A2(n7998), .ZN(n5304) );
  INV_X1 U6964 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n8405) );
  OR2_X1 U6965 ( .A1(n5285), .A2(n8405), .ZN(n5303) );
  OR2_X1 U6966 ( .A1(n9552), .A2(n7936), .ZN(n5811) );
  NAND2_X1 U6967 ( .A1(n9552), .A2(n7936), .ZN(n5812) );
  MUX2_X1 U6968 ( .A(n6993), .B(n5310), .S(n4399), .Z(n5312) );
  INV_X1 U6969 ( .A(SI_9_), .ZN(n5311) );
  INV_X1 U6970 ( .A(n5312), .ZN(n5313) );
  NAND2_X1 U6971 ( .A1(n5313), .A2(SI_9_), .ZN(n5314) );
  XNOR2_X1 U6972 ( .A(n5328), .B(n5102), .ZN(n6989) );
  NAND2_X1 U6973 ( .A1(n6989), .A2(n5635), .ZN(n5317) );
  NAND2_X1 U6974 ( .A1(n5335), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5315) );
  XNOR2_X1 U6975 ( .A(n5315), .B(P2_IR_REG_9__SCAN_IN), .ZN(n7731) );
  AOI22_X1 U6976 ( .A1(n5539), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n4375), .B2(
        n7731), .ZN(n5316) );
  NAND2_X1 U6977 ( .A1(n5317), .A2(n5316), .ZN(n7965) );
  NAND2_X1 U6978 ( .A1(n5225), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5327) );
  INV_X1 U6979 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n8005) );
  OR2_X1 U6980 ( .A1(n5260), .A2(n8005), .ZN(n5326) );
  INV_X1 U6981 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5318) );
  OAI21_X1 U6982 ( .B1(n5321), .B2(n5319), .A(n5318), .ZN(n5322) );
  NAND2_X1 U6983 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_REG3_REG_9__SCAN_IN), 
        .ZN(n5320) );
  OR2_X2 U6984 ( .A1(n5321), .A2(n5320), .ZN(n5339) );
  NAND2_X1 U6985 ( .A1(n5322), .A2(n5339), .ZN(n8007) );
  OR2_X1 U6986 ( .A1(n4395), .A2(n8007), .ZN(n5325) );
  INV_X1 U6987 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n5323) );
  OR2_X1 U6988 ( .A1(n5285), .A2(n5323), .ZN(n5324) );
  OR2_X1 U6989 ( .A1(n7965), .A2(n7986), .ZN(n5923) );
  INV_X1 U6990 ( .A(n5816), .ZN(n5922) );
  NAND2_X1 U6991 ( .A1(n5328), .A2(n5102), .ZN(n5330) );
  NAND2_X1 U6992 ( .A1(n5330), .A2(n5329), .ZN(n5345) );
  MUX2_X1 U6993 ( .A(n6996), .B(n6998), .S(n4398), .Z(n5332) );
  INV_X1 U6994 ( .A(SI_10_), .ZN(n5331) );
  INV_X1 U6995 ( .A(n5332), .ZN(n5333) );
  NAND2_X1 U6996 ( .A1(n5333), .A2(SI_10_), .ZN(n5334) );
  NAND2_X1 U6997 ( .A1(n6995), .A2(n5635), .ZN(n5338) );
  NOR2_X1 U6998 ( .A1(n5335), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n5348) );
  OR2_X1 U6999 ( .A1(n5348), .A2(n5133), .ZN(n5336) );
  XNOR2_X1 U7000 ( .A(n5336), .B(P2_IR_REG_10__SCAN_IN), .ZN(n8142) );
  AOI22_X1 U7001 ( .A1(n5539), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n4375), .B2(
        n8142), .ZN(n5337) );
  NAND2_X1 U7002 ( .A1(n5338), .A2(n5337), .ZN(n9547) );
  NAND2_X1 U7003 ( .A1(n5707), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5344) );
  INV_X1 U7004 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7732) );
  OR2_X1 U7005 ( .A1(n5260), .A2(n7732), .ZN(n5343) );
  INV_X1 U7006 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n8398) );
  OR2_X1 U7007 ( .A1(n5744), .A2(n8398), .ZN(n5342) );
  NAND2_X1 U7008 ( .A1(n5339), .A2(n8247), .ZN(n5340) );
  NAND2_X1 U7009 ( .A1(n5353), .A2(n5340), .ZN(n8126) );
  OR2_X1 U7010 ( .A1(n4394), .A2(n8126), .ZN(n5341) );
  OR2_X1 U7011 ( .A1(n9547), .A2(n8159), .ZN(n5817) );
  INV_X1 U7012 ( .A(n5818), .ZN(n5820) );
  MUX2_X1 U7013 ( .A(n7025), .B(n8414), .S(n4399), .Z(n5366) );
  XNOR2_X1 U7014 ( .A(n5360), .B(n5361), .ZN(n7022) );
  NAND2_X1 U7015 ( .A1(n7022), .A2(n5635), .ZN(n5351) );
  INV_X1 U7016 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5347) );
  NAND2_X1 U7017 ( .A1(n5348), .A2(n5347), .ZN(n5375) );
  NAND2_X1 U7018 ( .A1(n5375), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5349) );
  XNOR2_X1 U7019 ( .A(n5349), .B(P2_IR_REG_11__SCAN_IN), .ZN(n9048) );
  AOI22_X1 U7020 ( .A1(n5539), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n4375), .B2(
        n9048), .ZN(n5350) );
  NAND2_X1 U7021 ( .A1(n5225), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5358) );
  INV_X1 U7022 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n5352) );
  OR2_X1 U7023 ( .A1(n5285), .A2(n5352), .ZN(n5357) );
  INV_X1 U7024 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n9042) );
  NAND2_X1 U7025 ( .A1(n5353), .A2(n9042), .ZN(n5354) );
  NAND2_X1 U7026 ( .A1(n5380), .A2(n5354), .ZN(n8171) );
  OR2_X1 U7027 ( .A1(n4394), .A2(n8171), .ZN(n5356) );
  INV_X1 U7028 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n8145) );
  OR2_X1 U7029 ( .A1(n5260), .A2(n8145), .ZN(n5355) );
  NOR2_X1 U7030 ( .A1(n9541), .A2(n8657), .ZN(n5825) );
  INV_X1 U7031 ( .A(n5825), .ZN(n5359) );
  NAND2_X1 U7032 ( .A1(n5359), .A2(n5827), .ZN(n8551) );
  INV_X1 U7033 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n5362) );
  MUX2_X1 U7034 ( .A(n7095), .B(n5362), .S(n4398), .Z(n5363) );
  INV_X1 U7035 ( .A(SI_12_), .ZN(n8456) );
  NAND2_X1 U7036 ( .A1(n5363), .A2(n8456), .ZN(n5418) );
  INV_X1 U7037 ( .A(n5363), .ZN(n5364) );
  NAND2_X1 U7038 ( .A1(n5364), .A2(SI_12_), .ZN(n5365) );
  NAND2_X1 U7039 ( .A1(n5418), .A2(n5365), .ZN(n5372) );
  INV_X1 U7040 ( .A(n5372), .ZN(n5368) );
  INV_X1 U7041 ( .A(n5366), .ZN(n5367) );
  NAND2_X1 U7042 ( .A1(n5367), .A2(SI_11_), .ZN(n5370) );
  NAND2_X1 U7043 ( .A1(n5371), .A2(n5370), .ZN(n5373) );
  NAND2_X1 U7044 ( .A1(n5373), .A2(n5372), .ZN(n5374) );
  NAND2_X1 U7045 ( .A1(n5426), .A2(n5374), .ZN(n7094) );
  NAND2_X1 U7046 ( .A1(n7094), .A2(n5635), .ZN(n5378) );
  NAND2_X1 U7047 ( .A1(n5388), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5376) );
  XNOR2_X1 U7048 ( .A(n5376), .B(P2_IR_REG_12__SCAN_IN), .ZN(n8649) );
  AOI22_X1 U7049 ( .A1(n5539), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n8649), .B2(
        n4375), .ZN(n5377) );
  NAND2_X1 U7050 ( .A1(n5707), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5385) );
  INV_X1 U7051 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n8139) );
  OR2_X1 U7052 ( .A1(n5744), .A2(n8139), .ZN(n5384) );
  INV_X1 U7053 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n8187) );
  OR2_X1 U7054 ( .A1(n5260), .A2(n8187), .ZN(n5383) );
  INV_X1 U7055 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n8149) );
  NAND2_X1 U7056 ( .A1(n5380), .A2(n8149), .ZN(n5381) );
  NAND2_X1 U7057 ( .A1(n5393), .A2(n5381), .ZN(n8663) );
  OR2_X1 U7058 ( .A1(n4395), .A2(n8663), .ZN(n5382) );
  INV_X1 U7059 ( .A(n8661), .ZN(n8973) );
  NAND2_X1 U7060 ( .A1(n9536), .A2(n8661), .ZN(n5828) );
  MUX2_X1 U7061 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n4398), .Z(n5386) );
  INV_X1 U7062 ( .A(n5386), .ZN(n5387) );
  INV_X1 U7063 ( .A(SI_13_), .ZN(n8399) );
  AND2_X1 U7064 ( .A1(n5421), .A2(n5419), .ZN(n5399) );
  NAND2_X1 U7065 ( .A1(n7109), .A2(n5635), .ZN(n5390) );
  OAI21_X1 U7066 ( .B1(n5388), .B2(P2_IR_REG_12__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5404) );
  XNOR2_X1 U7067 ( .A(n5404), .B(P2_IR_REG_13__SCAN_IN), .ZN(n8681) );
  AOI22_X1 U7068 ( .A1(n8681), .A2(n4375), .B1(n5539), .B2(
        P1_DATAO_REG_13__SCAN_IN), .ZN(n5389) );
  NAND2_X1 U7069 ( .A1(n5707), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5398) );
  INV_X1 U7070 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n5391) );
  OR2_X1 U7071 ( .A1(n5260), .A2(n5391), .ZN(n5397) );
  INV_X1 U7072 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n8647) );
  OR2_X1 U7073 ( .A1(n5744), .A2(n8647), .ZN(n5396) );
  INV_X1 U7074 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5392) );
  NAND2_X1 U7075 ( .A1(n5393), .A2(n5392), .ZN(n5394) );
  NAND2_X1 U7076 ( .A1(n5412), .A2(n5394), .ZN(n8975) );
  OR2_X1 U7077 ( .A1(n4395), .A2(n8975), .ZN(n5395) );
  NAND4_X1 U7078 ( .A1(n5398), .A2(n5397), .A3(n5396), .A4(n5395), .ZN(n9028)
         );
  NAND2_X1 U7079 ( .A1(n8723), .A2(n9028), .ZN(n5833) );
  INV_X1 U7080 ( .A(n9028), .ZN(n8879) );
  NAND2_X1 U7081 ( .A1(n9531), .A2(n8879), .ZN(n5836) );
  NAND2_X1 U7082 ( .A1(n5833), .A2(n5836), .ZN(n5932) );
  NAND2_X1 U7083 ( .A1(n5400), .A2(n5399), .ZN(n5401) );
  NAND2_X1 U7084 ( .A1(n5401), .A2(n5419), .ZN(n5402) );
  MUX2_X1 U7085 ( .A(n7115), .B(n8428), .S(n4399), .Z(n5427) );
  NAND2_X1 U7086 ( .A1(n7113), .A2(n5635), .ZN(n5410) );
  INV_X1 U7087 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5403) );
  NAND2_X1 U7088 ( .A1(n5404), .A2(n5403), .ZN(n5405) );
  NAND2_X1 U7089 ( .A1(n5405), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5407) );
  INV_X1 U7090 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5406) );
  NAND2_X1 U7091 ( .A1(n5407), .A2(n5406), .ZN(n5435) );
  OR2_X1 U7092 ( .A1(n5407), .A2(n5406), .ZN(n5408) );
  AOI22_X1 U7093 ( .A1(n9059), .A2(n4375), .B1(n5539), .B2(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n5409) );
  NAND2_X2 U7094 ( .A1(n5410), .A2(n5409), .ZN(n9526) );
  NAND2_X1 U7095 ( .A1(n5707), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5417) );
  INV_X1 U7096 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8680) );
  OR2_X1 U7097 ( .A1(n5744), .A2(n8680), .ZN(n5416) );
  INV_X1 U7098 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n8617) );
  OR2_X1 U7099 ( .A1(n5260), .A2(n8617), .ZN(n5415) );
  INV_X1 U7100 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n5411) );
  NAND2_X1 U7101 ( .A1(n5412), .A2(n5411), .ZN(n5413) );
  NAND2_X1 U7102 ( .A1(n5440), .A2(n5413), .ZN(n8885) );
  OR2_X1 U7103 ( .A1(n4394), .A2(n8885), .ZN(n5414) );
  NAND2_X1 U7104 ( .A1(n9526), .A2(n9012), .ZN(n5840) );
  AND2_X2 U7105 ( .A1(n5839), .A2(n5840), .ZN(n8613) );
  INV_X1 U7106 ( .A(n5418), .ZN(n5422) );
  INV_X1 U7107 ( .A(n5427), .ZN(n5428) );
  NAND2_X1 U7108 ( .A1(n5428), .A2(SI_14_), .ZN(n5429) );
  MUX2_X1 U7109 ( .A(n7117), .B(n7119), .S(n4399), .Z(n5432) );
  INV_X1 U7110 ( .A(SI_15_), .ZN(n5431) );
  INV_X1 U7111 ( .A(n5432), .ZN(n5433) );
  NAND2_X1 U7112 ( .A1(n5433), .A2(SI_15_), .ZN(n5434) );
  XNOR2_X1 U7113 ( .A(n5448), .B(n5447), .ZN(n7116) );
  NAND2_X1 U7114 ( .A1(n7116), .A2(n5183), .ZN(n5438) );
  NAND2_X1 U7115 ( .A1(n5435), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5436) );
  XNOR2_X1 U7116 ( .A(n5436), .B(P2_IR_REG_15__SCAN_IN), .ZN(n9078) );
  AOI22_X1 U7117 ( .A1(n9078), .A2(n4375), .B1(n5539), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n5437) );
  INV_X1 U7118 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n5439) );
  OR2_X2 U7119 ( .A1(n5440), .A2(n5439), .ZN(n5462) );
  NAND2_X1 U7120 ( .A1(n5440), .A2(n5439), .ZN(n5441) );
  AND2_X1 U7121 ( .A1(n5462), .A2(n5441), .ZN(n9420) );
  NAND2_X1 U7122 ( .A1(n9420), .A2(n5698), .ZN(n5445) );
  NAND2_X1 U7123 ( .A1(n5707), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5444) );
  INV_X1 U7124 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n9061) );
  OR2_X1 U7125 ( .A1(n5744), .A2(n9061), .ZN(n5443) );
  INV_X1 U7126 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8249) );
  OR2_X1 U7127 ( .A1(n5260), .A2(n8249), .ZN(n5442) );
  NAND2_X1 U7128 ( .A1(n9522), .A2(n9385), .ZN(n5844) );
  NAND2_X1 U7129 ( .A1(n9409), .A2(n9408), .ZN(n9407) );
  NAND2_X1 U7130 ( .A1(n9407), .A2(n5845), .ZN(n9389) );
  INV_X1 U7131 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7301) );
  INV_X1 U7132 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n7303) );
  MUX2_X1 U7133 ( .A(n7301), .B(n7303), .S(n4398), .Z(n5450) );
  INV_X1 U7134 ( .A(SI_16_), .ZN(n5449) );
  NAND2_X1 U7135 ( .A1(n5450), .A2(n5449), .ZN(n5468) );
  INV_X1 U7136 ( .A(n5450), .ZN(n5451) );
  NAND2_X1 U7137 ( .A1(n5451), .A2(SI_16_), .ZN(n5452) );
  XNOR2_X1 U7138 ( .A(n5467), .B(n5098), .ZN(n7300) );
  NAND2_X1 U7139 ( .A1(n7300), .A2(n5635), .ZN(n5461) );
  INV_X1 U7140 ( .A(n4537), .ZN(n5455) );
  NAND2_X1 U7141 ( .A1(n5455), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5456) );
  MUX2_X1 U7142 ( .A(n5456), .B(P2_IR_REG_31__SCAN_IN), .S(n5458), .Z(n5457)
         );
  INV_X1 U7143 ( .A(n5457), .ZN(n5459) );
  NOR2_X1 U7144 ( .A1(n5459), .A2(n5488), .ZN(n9087) );
  AOI22_X1 U7145 ( .A1(n5539), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n4375), .B2(
        n9087), .ZN(n5460) );
  AOI22_X1 U7146 ( .A1(n5225), .A2(P2_REG1_REG_16__SCAN_IN), .B1(n5707), .B2(
        P2_REG0_REG_16__SCAN_IN), .ZN(n5466) );
  INV_X1 U7147 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n8304) );
  NAND2_X1 U7148 ( .A1(n5462), .A2(n8304), .ZN(n5463) );
  AND2_X1 U7149 ( .A1(n5493), .A2(n5463), .ZN(n9397) );
  NAND2_X1 U7150 ( .A1(n9397), .A2(n5698), .ZN(n5465) );
  INV_X1 U7151 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n9081) );
  OR2_X1 U7152 ( .A1(n5260), .A2(n9081), .ZN(n5464) );
  NAND2_X1 U7153 ( .A1(n9398), .A2(n9027), .ZN(n9363) );
  NAND2_X1 U7154 ( .A1(n5850), .A2(n9363), .ZN(n9388) );
  OR2_X2 U7155 ( .A1(n9389), .A2(n9388), .ZN(n9391) );
  INV_X1 U7156 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n5472) );
  INV_X1 U7157 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n5471) );
  MUX2_X1 U7158 ( .A(n5472), .B(n5471), .S(n4399), .Z(n5473) );
  XNOR2_X1 U7159 ( .A(n5473), .B(SI_17_), .ZN(n5487) );
  INV_X1 U7160 ( .A(n5487), .ZN(n5476) );
  INV_X1 U7161 ( .A(n5473), .ZN(n5474) );
  NAND2_X1 U7162 ( .A1(n5474), .A2(SI_17_), .ZN(n5475) );
  MUX2_X1 U7163 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n4399), .Z(n5499) );
  XNOR2_X1 U7164 ( .A(n5499), .B(SI_18_), .ZN(n5525) );
  XNOR2_X1 U7165 ( .A(n5526), .B(n5525), .ZN(n7439) );
  NAND2_X1 U7166 ( .A1(n7439), .A2(n5635), .ZN(n5480) );
  NAND2_X1 U7167 ( .A1(n4491), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5478) );
  XNOR2_X1 U7168 ( .A(n5478), .B(P2_IR_REG_18__SCAN_IN), .ZN(n9120) );
  AOI22_X1 U7169 ( .A1(n5539), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n4375), .B2(
        n9120), .ZN(n5479) );
  INV_X1 U7170 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n8989) );
  NAND2_X1 U7171 ( .A1(n5495), .A2(n8989), .ZN(n5481) );
  AND2_X1 U7172 ( .A1(n5542), .A2(n5481), .ZN(n9343) );
  NAND2_X1 U7173 ( .A1(n9343), .A2(n5698), .ZN(n5485) );
  AOI22_X1 U7174 ( .A1(n5225), .A2(P2_REG1_REG_18__SCAN_IN), .B1(n4393), .B2(
        P2_REG2_REG_18__SCAN_IN), .ZN(n5484) );
  NAND2_X1 U7175 ( .A1(n5707), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n5483) );
  NAND2_X1 U7176 ( .A1(n9499), .A2(n9147), .ZN(n5921) );
  NAND2_X1 U7177 ( .A1(n7296), .A2(n5635), .ZN(n5492) );
  NAND2_X1 U7178 ( .A1(n5489), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5490) );
  XNOR2_X1 U7179 ( .A(n5490), .B(P2_IR_REG_17__SCAN_IN), .ZN(n9107) );
  AOI22_X1 U7180 ( .A1(n5539), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n4375), .B2(
        n9107), .ZN(n5491) );
  INV_X1 U7181 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8944) );
  NAND2_X1 U7182 ( .A1(n5493), .A2(n8944), .ZN(n5494) );
  NAND2_X1 U7183 ( .A1(n5495), .A2(n5494), .ZN(n9374) );
  OR2_X1 U7184 ( .A1(n9374), .A2(n4395), .ZN(n5498) );
  AOI22_X1 U7185 ( .A1(n5225), .A2(P2_REG1_REG_17__SCAN_IN), .B1(n4393), .B2(
        P2_REG2_REG_17__SCAN_IN), .ZN(n5497) );
  NAND2_X1 U7186 ( .A1(n5707), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5496) );
  NAND2_X1 U7187 ( .A1(n9508), .A2(n9387), .ZN(n5853) );
  AND3_X1 U7188 ( .A1(n5921), .A2(n5853), .A3(n9363), .ZN(n9271) );
  NAND2_X1 U7189 ( .A1(n5499), .A2(SI_18_), .ZN(n5527) );
  MUX2_X1 U7190 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(P2_DATAO_REG_19__SCAN_IN), 
        .S(n4399), .Z(n5501) );
  NAND2_X1 U7191 ( .A1(n5501), .A2(SI_19_), .ZN(n5530) );
  NAND2_X1 U7192 ( .A1(n5527), .A2(n5530), .ZN(n5505) );
  NOR2_X1 U7193 ( .A1(n5499), .A2(SI_18_), .ZN(n5500) );
  NAND2_X1 U7194 ( .A1(n5500), .A2(n5530), .ZN(n5503) );
  INV_X1 U7195 ( .A(n5501), .ZN(n5502) );
  INV_X1 U7196 ( .A(SI_19_), .ZN(n8344) );
  NAND2_X1 U7197 ( .A1(n5502), .A2(n8344), .ZN(n5529) );
  INV_X1 U7198 ( .A(n5512), .ZN(n5510) );
  INV_X1 U7199 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n8454) );
  INV_X1 U7200 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7627) );
  MUX2_X1 U7201 ( .A(n8454), .B(n7627), .S(n4398), .Z(n5507) );
  INV_X1 U7202 ( .A(SI_20_), .ZN(n5506) );
  NAND2_X1 U7203 ( .A1(n5507), .A2(n5506), .ZN(n5550) );
  INV_X1 U7204 ( .A(n5507), .ZN(n5508) );
  NAND2_X1 U7205 ( .A1(n5508), .A2(SI_20_), .ZN(n5509) );
  NAND2_X1 U7206 ( .A1(n5550), .A2(n5509), .ZN(n5511) );
  NAND2_X1 U7207 ( .A1(n5510), .A2(n5511), .ZN(n5513) );
  NAND2_X1 U7208 ( .A1(n5513), .A2(n5551), .ZN(n7624) );
  NAND2_X1 U7209 ( .A1(n7624), .A2(n5183), .ZN(n5516) );
  OR2_X1 U7210 ( .A1(n5514), .A2(n8454), .ZN(n5515) );
  INV_X1 U7211 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n8305) );
  OR2_X2 U7212 ( .A1(n5544), .A2(n8305), .ZN(n5554) );
  NAND2_X1 U7213 ( .A1(n5544), .A2(n8305), .ZN(n5518) );
  NAND2_X1 U7214 ( .A1(n5554), .A2(n5518), .ZN(n8966) );
  OR2_X1 U7215 ( .A1(n8966), .A2(n4394), .ZN(n5524) );
  INV_X1 U7216 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n5521) );
  NAND2_X1 U7217 ( .A1(n5707), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n5520) );
  NAND2_X1 U7218 ( .A1(n4393), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n5519) );
  OAI211_X1 U7219 ( .C1(n5744), .C2(n5521), .A(n5520), .B(n5519), .ZN(n5522)
         );
  INV_X1 U7220 ( .A(n5522), .ZN(n5523) );
  NAND2_X1 U7221 ( .A1(n5524), .A2(n5523), .ZN(n9332) );
  NAND2_X1 U7222 ( .A1(n9489), .A2(n8918), .ZN(n5920) );
  NAND2_X1 U7223 ( .A1(n5528), .A2(n5527), .ZN(n5532) );
  NAND2_X1 U7224 ( .A1(n5530), .A2(n5529), .ZN(n5531) );
  NAND2_X1 U7225 ( .A1(n5534), .A2(P2_IR_REG_19__SCAN_IN), .ZN(n5537) );
  INV_X1 U7226 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5535) );
  NAND2_X1 U7227 ( .A1(n5536), .A2(n5535), .ZN(n5764) );
  AOI22_X1 U7228 ( .A1(n5539), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n9361), .B2(
        n4375), .ZN(n5540) );
  INV_X1 U7229 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n5541) );
  NAND2_X1 U7230 ( .A1(n5542), .A2(n5541), .ZN(n5543) );
  NAND2_X1 U7231 ( .A1(n5544), .A2(n5543), .ZN(n8904) );
  OR2_X1 U7232 ( .A1(n8904), .A2(n4394), .ZN(n5549) );
  INV_X1 U7233 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n9122) );
  NAND2_X1 U7234 ( .A1(n5707), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n5546) );
  NAND2_X1 U7235 ( .A1(n4393), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n5545) );
  OAI211_X1 U7236 ( .C1(n5744), .C2(n9122), .A(n5546), .B(n5545), .ZN(n5547)
         );
  INV_X1 U7237 ( .A(n5547), .ZN(n5548) );
  NAND2_X1 U7238 ( .A1(n5920), .A2(n9309), .ZN(n5872) );
  INV_X1 U7239 ( .A(n5872), .ZN(n9291) );
  NAND2_X1 U7240 ( .A1(n5551), .A2(n5550), .ZN(n5576) );
  INV_X1 U7241 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7758) );
  INV_X1 U7242 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7745) );
  MUX2_X1 U7243 ( .A(n7758), .B(n7745), .S(n4398), .Z(n5572) );
  XNOR2_X1 U7244 ( .A(n5572), .B(SI_21_), .ZN(n5571) );
  OR2_X1 U7245 ( .A1(n5514), .A2(n7758), .ZN(n5552) );
  INV_X1 U7246 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n5553) );
  NAND2_X1 U7247 ( .A1(n5554), .A2(n5553), .ZN(n5555) );
  NAND2_X1 U7248 ( .A1(n5096), .A2(n5698), .ZN(n5561) );
  INV_X1 U7249 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n5558) );
  NAND2_X1 U7250 ( .A1(n4393), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n5557) );
  NAND2_X1 U7251 ( .A1(n5707), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n5556) );
  OAI211_X1 U7252 ( .C1(n5744), .C2(n5558), .A(n5557), .B(n5556), .ZN(n5559)
         );
  INV_X1 U7253 ( .A(n5559), .ZN(n5560) );
  AND2_X2 U7254 ( .A1(n5561), .A2(n5560), .ZN(n9280) );
  NAND2_X1 U7255 ( .A1(n9484), .A2(n9280), .ZN(n5874) );
  AND2_X1 U7256 ( .A1(n9271), .A2(n9274), .ZN(n5562) );
  NAND2_X1 U7257 ( .A1(n9391), .A2(n5562), .ZN(n5568) );
  INV_X1 U7258 ( .A(n9274), .ZN(n5566) );
  INV_X1 U7259 ( .A(n5849), .ZN(n9327) );
  NAND2_X1 U7260 ( .A1(n5921), .A2(n9327), .ZN(n5564) );
  NAND2_X1 U7261 ( .A1(n5564), .A2(n5856), .ZN(n5565) );
  NOR2_X1 U7262 ( .A1(n9328), .A2(n5565), .ZN(n9272) );
  OR2_X1 U7263 ( .A1(n5566), .A2(n9272), .ZN(n5567) );
  INV_X1 U7264 ( .A(n5874), .ZN(n5570) );
  XNOR2_X1 U7265 ( .A(n9484), .B(n9313), .ZN(n9297) );
  AND2_X1 U7266 ( .A1(n9292), .A2(n9297), .ZN(n5569) );
  INV_X1 U7267 ( .A(n5571), .ZN(n5575) );
  INV_X1 U7268 ( .A(n5572), .ZN(n5573) );
  NAND2_X1 U7269 ( .A1(n5573), .A2(SI_21_), .ZN(n5574) );
  INV_X1 U7270 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n8865) );
  INV_X1 U7271 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8379) );
  MUX2_X1 U7272 ( .A(n8865), .B(n8379), .S(n4398), .Z(n5578) );
  INV_X1 U7273 ( .A(SI_22_), .ZN(n5577) );
  NAND2_X1 U7274 ( .A1(n5578), .A2(n5577), .ZN(n5594) );
  INV_X1 U7275 ( .A(n5578), .ZN(n5579) );
  NAND2_X1 U7276 ( .A1(n5579), .A2(SI_22_), .ZN(n5580) );
  NAND2_X1 U7277 ( .A1(n5594), .A2(n5580), .ZN(n5595) );
  XNOR2_X1 U7278 ( .A(n5596), .B(n5595), .ZN(n7891) );
  NAND2_X1 U7279 ( .A1(n7891), .A2(n5183), .ZN(n5583) );
  OR2_X1 U7280 ( .A1(n5514), .A2(n8865), .ZN(n5582) );
  NAND2_X1 U7281 ( .A1(n5583), .A2(n5582), .ZN(n5593) );
  INV_X1 U7282 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n5584) );
  NAND2_X1 U7283 ( .A1(n5585), .A2(n5584), .ZN(n5586) );
  AND2_X1 U7284 ( .A1(n5605), .A2(n5586), .ZN(n9268) );
  NAND2_X1 U7285 ( .A1(n9268), .A2(n5698), .ZN(n5592) );
  INV_X1 U7286 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n5589) );
  NAND2_X1 U7287 ( .A1(n5707), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n5588) );
  NAND2_X1 U7288 ( .A1(n4393), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n5587) );
  OAI211_X1 U7289 ( .C1(n5744), .C2(n5589), .A(n5588), .B(n5587), .ZN(n5590)
         );
  INV_X1 U7290 ( .A(n5590), .ZN(n5591) );
  NAND2_X1 U7291 ( .A1(n5593), .A2(n8916), .ZN(n5918) );
  INV_X1 U7292 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n8017) );
  INV_X1 U7293 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n8022) );
  MUX2_X1 U7294 ( .A(n8017), .B(n8022), .S(n4399), .Z(n5597) );
  INV_X1 U7295 ( .A(SI_23_), .ZN(n8430) );
  NAND2_X1 U7296 ( .A1(n5597), .A2(n8430), .ZN(n5631) );
  INV_X1 U7297 ( .A(n5597), .ZN(n5598) );
  NAND2_X1 U7298 ( .A1(n5598), .A2(SI_23_), .ZN(n5599) );
  OR2_X1 U7299 ( .A1(n5652), .A2(n5650), .ZN(n5600) );
  NAND2_X1 U7300 ( .A1(n8018), .A2(n5183), .ZN(n5602) );
  OR2_X1 U7301 ( .A1(n5514), .A2(n8017), .ZN(n5601) );
  INV_X1 U7302 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n5604) );
  NAND2_X1 U7303 ( .A1(n5605), .A2(n5604), .ZN(n5606) );
  NAND2_X1 U7304 ( .A1(n5638), .A2(n5606), .ZN(n8895) );
  OR2_X1 U7305 ( .A1(n8895), .A2(n4395), .ZN(n5612) );
  INV_X1 U7306 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n5609) );
  NAND2_X1 U7307 ( .A1(n4393), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n5608) );
  NAND2_X1 U7308 ( .A1(n5707), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n5607) );
  OAI211_X1 U7309 ( .C1(n5744), .C2(n5609), .A(n5608), .B(n5607), .ZN(n5610)
         );
  INV_X1 U7310 ( .A(n5610), .ZN(n5611) );
  INV_X1 U7311 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n8135) );
  INV_X1 U7312 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n8134) );
  MUX2_X1 U7313 ( .A(n8135), .B(n8134), .S(n4398), .Z(n5613) );
  XNOR2_X1 U7314 ( .A(n5613), .B(SI_24_), .ZN(n5633) );
  NAND2_X1 U7315 ( .A1(n5632), .A2(n5654), .ZN(n5615) );
  INV_X1 U7316 ( .A(n5613), .ZN(n5614) );
  NAND2_X1 U7317 ( .A1(n5614), .A2(SI_24_), .ZN(n5648) );
  INV_X1 U7318 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n8523) );
  INV_X1 U7319 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n8520) );
  MUX2_X1 U7320 ( .A(n8523), .B(n8520), .S(n4399), .Z(n5617) );
  INV_X1 U7321 ( .A(SI_25_), .ZN(n5616) );
  NAND2_X1 U7322 ( .A1(n5617), .A2(n5616), .ZN(n5656) );
  INV_X1 U7323 ( .A(n5617), .ZN(n5618) );
  NAND2_X1 U7324 ( .A1(n5618), .A2(SI_25_), .ZN(n5619) );
  NAND2_X1 U7325 ( .A1(n5656), .A2(n5619), .ZN(n5647) );
  NAND2_X1 U7326 ( .A1(n8518), .A2(n5635), .ZN(n5622) );
  OR2_X1 U7327 ( .A1(n5514), .A2(n8523), .ZN(n5621) );
  INV_X1 U7328 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n8958) );
  INV_X1 U7329 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n5623) );
  NAND2_X1 U7330 ( .A1(n5640), .A2(n5623), .ZN(n5624) );
  NAND2_X1 U7331 ( .A1(n5669), .A2(n5624), .ZN(n9224) );
  INV_X1 U7332 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n5627) );
  NAND2_X1 U7333 ( .A1(n5225), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n5626) );
  NAND2_X1 U7334 ( .A1(n5707), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n5625) );
  OAI211_X1 U7335 ( .C1(n5260), .C2(n5627), .A(n5626), .B(n5625), .ZN(n5628)
         );
  INV_X1 U7336 ( .A(n5628), .ZN(n5629) );
  NAND2_X1 U7337 ( .A1(n9464), .A2(n9243), .ZN(n5889) );
  NAND2_X1 U7338 ( .A1(n8132), .A2(n5635), .ZN(n5637) );
  OR2_X1 U7339 ( .A1(n5514), .A2(n8135), .ZN(n5636) );
  NAND2_X1 U7340 ( .A1(n5638), .A2(n8958), .ZN(n5639) );
  NAND2_X1 U7341 ( .A1(n9238), .A2(n5698), .ZN(n5646) );
  INV_X1 U7342 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n5643) );
  NAND2_X1 U7343 ( .A1(n4393), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n5642) );
  NAND2_X1 U7344 ( .A1(n5707), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n5641) );
  OAI211_X1 U7345 ( .C1(n5744), .C2(n5643), .A(n5642), .B(n5641), .ZN(n5644)
         );
  INV_X1 U7346 ( .A(n5644), .ZN(n5645) );
  NAND2_X1 U7347 ( .A1(n9468), .A2(n8954), .ZN(n5917) );
  NAND2_X1 U7348 ( .A1(n5889), .A2(n5917), .ZN(n5679) );
  INV_X1 U7349 ( .A(n5889), .ZN(n5676) );
  INV_X1 U7350 ( .A(n5647), .ZN(n5649) );
  INV_X1 U7351 ( .A(n5653), .ZN(n5655) );
  NAND2_X1 U7352 ( .A1(n5657), .A2(n5656), .ZN(n5658) );
  INV_X1 U7353 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n8195) );
  INV_X1 U7354 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n8198) );
  MUX2_X1 U7355 ( .A(n8195), .B(n8198), .S(n4398), .Z(n5659) );
  INV_X1 U7356 ( .A(SI_26_), .ZN(n8315) );
  NAND2_X1 U7357 ( .A1(n5659), .A2(n8315), .ZN(n5681) );
  INV_X1 U7358 ( .A(n5659), .ZN(n5660) );
  NAND2_X1 U7359 ( .A1(n5660), .A2(SI_26_), .ZN(n5661) );
  NAND2_X1 U7360 ( .A1(n5681), .A2(n5661), .ZN(n5663) );
  NAND2_X1 U7361 ( .A1(n5662), .A2(n5663), .ZN(n5666) );
  INV_X1 U7362 ( .A(n5662), .ZN(n5665) );
  INV_X1 U7363 ( .A(n5663), .ZN(n5664) );
  NAND2_X1 U7364 ( .A1(n5666), .A2(n5682), .ZN(n8192) );
  NAND2_X1 U7365 ( .A1(n8192), .A2(n5635), .ZN(n5668) );
  OR2_X1 U7366 ( .A1(n5514), .A2(n8195), .ZN(n5667) );
  INV_X1 U7367 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n9001) );
  OR2_X2 U7368 ( .A1(n5669), .A2(n9001), .ZN(n5703) );
  NAND2_X1 U7369 ( .A1(n5669), .A2(n9001), .ZN(n5670) );
  NAND2_X1 U7370 ( .A1(n9000), .A2(n5698), .ZN(n5675) );
  INV_X1 U7371 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8401) );
  NAND2_X1 U7372 ( .A1(n4393), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n5672) );
  NAND2_X1 U7373 ( .A1(n5707), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n5671) );
  OAI211_X1 U7374 ( .C1(n5744), .C2(n8401), .A(n5672), .B(n5671), .ZN(n5673)
         );
  INV_X1 U7375 ( .A(n5673), .ZN(n5674) );
  NAND2_X1 U7376 ( .A1(n5675), .A2(n5674), .ZN(n9025) );
  NAND2_X1 U7377 ( .A1(n9152), .A2(n9025), .ZN(n5892) );
  OAI211_X1 U7378 ( .C1(n5676), .C2(n9206), .A(n4979), .B(n9207), .ZN(n5677)
         );
  INV_X1 U7379 ( .A(n5677), .ZN(n5678) );
  INV_X1 U7380 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n8675) );
  INV_X1 U7381 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n6344) );
  MUX2_X1 U7382 ( .A(n8675), .B(n6344), .S(n4399), .Z(n5684) );
  INV_X1 U7383 ( .A(SI_27_), .ZN(n5683) );
  NAND2_X1 U7384 ( .A1(n5684), .A2(n5683), .ZN(n5699) );
  INV_X1 U7385 ( .A(n5684), .ZN(n5685) );
  NAND2_X1 U7386 ( .A1(n5685), .A2(SI_27_), .ZN(n5686) );
  NAND2_X1 U7387 ( .A1(n5699), .A2(n5686), .ZN(n5688) );
  NAND2_X1 U7388 ( .A1(n5687), .A2(n5688), .ZN(n5691) );
  INV_X1 U7389 ( .A(n5688), .ZN(n5689) );
  NAND2_X1 U7390 ( .A1(n5691), .A2(n5700), .ZN(n8640) );
  NAND2_X1 U7391 ( .A1(n8640), .A2(n5183), .ZN(n5693) );
  OR2_X1 U7392 ( .A1(n5514), .A2(n8675), .ZN(n5692) );
  XNOR2_X1 U7393 ( .A(n5703), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n9193) );
  INV_X1 U7394 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n5696) );
  NAND2_X1 U7395 ( .A1(n4393), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n5695) );
  NAND2_X1 U7396 ( .A1(n5707), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n5694) );
  OAI211_X1 U7397 ( .C1(n5744), .C2(n5696), .A(n5695), .B(n5694), .ZN(n5697)
         );
  OR2_X2 U7398 ( .A1(n9454), .A2(n8825), .ZN(n5895) );
  NAND2_X1 U7399 ( .A1(n9454), .A2(n8825), .ZN(n5898) );
  INV_X1 U7400 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8855) );
  INV_X1 U7401 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n10250) );
  MUX2_X1 U7402 ( .A(n8855), .B(n10250), .S(n4398), .Z(n5718) );
  XNOR2_X1 U7403 ( .A(n5718), .B(SI_28_), .ZN(n5715) );
  OR2_X1 U7404 ( .A1(n5514), .A2(n8855), .ZN(n5701) );
  INV_X1 U7405 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n8869) );
  INV_X1 U7406 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n8827) );
  OAI21_X1 U7407 ( .B1(n5703), .B2(n8869), .A(n8827), .ZN(n5706) );
  INV_X1 U7408 ( .A(n5703), .ZN(n5705) );
  AND2_X1 U7409 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(P2_REG3_REG_28__SCAN_IN), 
        .ZN(n5704) );
  NAND2_X1 U7410 ( .A1(n5705), .A2(n5704), .ZN(n9168) );
  NAND2_X1 U7411 ( .A1(n5706), .A2(n9168), .ZN(n9185) );
  INV_X1 U7412 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n5710) );
  NAND2_X1 U7413 ( .A1(n4393), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n5709) );
  NAND2_X1 U7414 ( .A1(n5707), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n5708) );
  OAI211_X1 U7415 ( .C1(n5744), .C2(n5710), .A(n5709), .B(n5708), .ZN(n5711)
         );
  INV_X1 U7416 ( .A(n5711), .ZN(n5712) );
  INV_X1 U7417 ( .A(n5897), .ZN(n5714) );
  NAND2_X1 U7418 ( .A1(n9180), .A2(n9179), .ZN(n9178) );
  INV_X1 U7419 ( .A(SI_28_), .ZN(n5717) );
  NAND2_X1 U7420 ( .A1(n5718), .A2(n5717), .ZN(n5719) );
  INV_X1 U7421 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8694) );
  INV_X1 U7422 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n10242) );
  MUX2_X1 U7423 ( .A(n8694), .B(n10242), .S(n4398), .Z(n5730) );
  XNOR2_X1 U7424 ( .A(n5730), .B(SI_29_), .ZN(n5721) );
  NAND2_X1 U7425 ( .A1(n8692), .A2(n5635), .ZN(n5723) );
  OR2_X1 U7426 ( .A1(n5514), .A2(n8694), .ZN(n5722) );
  OR2_X1 U7427 ( .A1(n9168), .A2(n4395), .ZN(n5728) );
  INV_X1 U7428 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n8403) );
  NAND2_X1 U7429 ( .A1(n4393), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n5725) );
  INV_X1 U7430 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n8283) );
  OR2_X1 U7431 ( .A1(n5285), .A2(n8283), .ZN(n5724) );
  OAI211_X1 U7432 ( .C1(n5744), .C2(n8403), .A(n5725), .B(n5724), .ZN(n5726)
         );
  INV_X1 U7433 ( .A(n5726), .ZN(n5727) );
  NOR2_X1 U7434 ( .A1(n9438), .A2(n8826), .ZN(n5902) );
  INV_X1 U7435 ( .A(n5902), .ZN(n5915) );
  NAND2_X1 U7436 ( .A1(n9438), .A2(n8826), .ZN(n5914) );
  INV_X1 U7437 ( .A(n5729), .ZN(n5731) );
  INV_X1 U7438 ( .A(n5730), .ZN(n5732) );
  NAND2_X1 U7439 ( .A1(n5732), .A2(SI_29_), .ZN(n5733) );
  MUX2_X1 U7440 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .S(n4399), .Z(n5754) );
  XNOR2_X1 U7441 ( .A(n5754), .B(SI_30_), .ZN(n5735) );
  NAND2_X1 U7442 ( .A1(n8856), .A2(n5183), .ZN(n5737) );
  INV_X1 U7443 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8858) );
  OR2_X1 U7444 ( .A1(n5514), .A2(n8858), .ZN(n5736) );
  INV_X1 U7445 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n5738) );
  OR2_X1 U7446 ( .A1(n5744), .A2(n5738), .ZN(n5742) );
  INV_X1 U7447 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n9135) );
  OR2_X1 U7448 ( .A1(n5260), .A2(n9135), .ZN(n5741) );
  INV_X1 U7449 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n5739) );
  OR2_X1 U7450 ( .A1(n5285), .A2(n5739), .ZN(n5740) );
  AND3_X1 U7451 ( .A1(n5742), .A2(n5741), .A3(n5740), .ZN(n9162) );
  OR2_X1 U7452 ( .A1(n9432), .A2(n9162), .ZN(n5909) );
  INV_X1 U7453 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n5743) );
  OR2_X1 U7454 ( .A1(n5744), .A2(n5743), .ZN(n5748) );
  INV_X1 U7455 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n8850) );
  OR2_X1 U7456 ( .A1(n5260), .A2(n8850), .ZN(n5747) );
  INV_X1 U7457 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n5745) );
  OR2_X1 U7458 ( .A1(n5285), .A2(n5745), .ZN(n5746) );
  AND3_X1 U7459 ( .A1(n5748), .A2(n5747), .A3(n5746), .ZN(n8849) );
  INV_X1 U7460 ( .A(n8849), .ZN(n7099) );
  INV_X1 U7461 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5750) );
  INV_X1 U7462 ( .A(n5754), .ZN(n5753) );
  INV_X1 U7463 ( .A(SI_30_), .ZN(n5752) );
  NOR2_X1 U7464 ( .A1(n5753), .A2(n5752), .ZN(n5755) );
  INV_X1 U7465 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n9587) );
  INV_X1 U7466 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n6378) );
  MUX2_X1 U7467 ( .A(n9587), .B(n6378), .S(n4399), .Z(n5757) );
  XNOR2_X1 U7468 ( .A(n5757), .B(SI_31_), .ZN(n5758) );
  NAND2_X1 U7469 ( .A1(n9583), .A2(n5635), .ZN(n5760) );
  OR2_X1 U7470 ( .A1(n5514), .A2(n9587), .ZN(n5759) );
  NAND2_X1 U7471 ( .A1(n9432), .A2(n9162), .ZN(n5907) );
  NAND2_X1 U7472 ( .A1(n8844), .A2(n8849), .ZN(n5910) );
  INV_X1 U7473 ( .A(n5910), .ZN(n5761) );
  AOI21_X1 U7474 ( .B1(n5762), .B2(n5913), .A(n5761), .ZN(n5763) );
  XNOR2_X1 U7475 ( .A(n5763), .B(n7537), .ZN(n5774) );
  INV_X1 U7476 ( .A(n5766), .ZN(n5767) );
  NAND2_X1 U7477 ( .A1(n5767), .A2(n5750), .ZN(n5768) );
  AND2_X1 U7478 ( .A1(n7543), .A2(n5955), .ZN(n7137) );
  NAND2_X1 U7479 ( .A1(n5770), .A2(n5769), .ZN(n5771) );
  XNOR2_X1 U7480 ( .A(n5945), .B(P2_IR_REG_23__SCAN_IN), .ZN(n7545) );
  AND2_X1 U7481 ( .A1(n7545), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7091) );
  INV_X1 U7482 ( .A(n5772), .ZN(n5773) );
  NAND2_X1 U7483 ( .A1(n5774), .A2(n5773), .ZN(n5961) );
  INV_X1 U7484 ( .A(n5775), .ZN(n5912) );
  AND2_X1 U7485 ( .A1(n5955), .A2(n9361), .ZN(n5776) );
  INV_X1 U7486 ( .A(n5919), .ZN(n5778) );
  NOR2_X1 U7487 ( .A1(n9484), .A2(n9280), .ZN(n5870) );
  NAND2_X1 U7488 ( .A1(n9292), .A2(n5877), .ZN(n5777) );
  NOR4_X1 U7489 ( .A1(n5778), .A2(n5870), .A3(n4816), .A4(n5777), .ZN(n5868)
         );
  NAND2_X1 U7490 ( .A1(n5780), .A2(n5779), .ZN(n5782) );
  OR2_X1 U7491 ( .A1(n5782), .A2(n5781), .ZN(n5783) );
  NAND2_X1 U7492 ( .A1(n7318), .A2(n7595), .ZN(n7597) );
  NAND2_X1 U7493 ( .A1(n7597), .A2(n5925), .ZN(n5787) );
  OAI211_X1 U7494 ( .C1(n5787), .C2(n7757), .A(n5784), .B(n5790), .ZN(n5785)
         );
  NAND2_X1 U7495 ( .A1(n5785), .A2(n5788), .ZN(n5793) );
  NAND2_X1 U7496 ( .A1(n5787), .A2(n5786), .ZN(n5789) );
  NAND2_X1 U7497 ( .A1(n5789), .A2(n5788), .ZN(n5791) );
  NAND2_X1 U7498 ( .A1(n5791), .A2(n5790), .ZN(n5792) );
  MUX2_X1 U7499 ( .A(n5793), .B(n5792), .S(n5877), .Z(n5795) );
  NOR3_X1 U7500 ( .A1(n5795), .A2(n5797), .A3(n5794), .ZN(n5796) );
  AOI21_X1 U7501 ( .B1(n7350), .B2(n5798), .A(n5797), .ZN(n5801) );
  INV_X1 U7502 ( .A(n5799), .ZN(n5800) );
  NOR3_X1 U7503 ( .A1(n5801), .A2(n5803), .A3(n5800), .ZN(n5802) );
  OAI22_X1 U7504 ( .A1(n5804), .A2(n5803), .B1(n5911), .B2(n5802), .ZN(n5806)
         );
  NAND2_X1 U7505 ( .A1(n5806), .A2(n5111), .ZN(n5810) );
  NAND2_X1 U7506 ( .A1(n10407), .A2(n5911), .ZN(n5808) );
  NAND2_X1 U7507 ( .A1(n5059), .A2(n5877), .ZN(n5807) );
  MUX2_X1 U7508 ( .A(n5808), .B(n5807), .S(n9033), .Z(n5809) );
  NAND3_X1 U7509 ( .A1(n5810), .A2(n7791), .A3(n5809), .ZN(n5814) );
  MUX2_X1 U7510 ( .A(n5812), .B(n5811), .S(n5911), .Z(n5813) );
  AOI211_X1 U7511 ( .C1(n5814), .C2(n5813), .A(n5818), .B(n5816), .ZN(n5815)
         );
  NAND2_X1 U7512 ( .A1(n5817), .A2(n5923), .ZN(n5824) );
  NOR2_X1 U7513 ( .A1(n5819), .A2(n5818), .ZN(n5822) );
  AOI21_X1 U7514 ( .B1(n5820), .B2(n5824), .A(n5825), .ZN(n5821) );
  MUX2_X1 U7515 ( .A(n5822), .B(n5821), .S(n5911), .Z(n5823) );
  INV_X1 U7516 ( .A(n5829), .ZN(n5826) );
  NOR2_X1 U7517 ( .A1(n5826), .A2(n5825), .ZN(n5832) );
  NAND3_X1 U7518 ( .A1(n5836), .A2(n5877), .A3(n5828), .ZN(n5831) );
  NAND3_X1 U7519 ( .A1(n5829), .A2(n5828), .A3(n5827), .ZN(n5830) );
  MUX2_X1 U7520 ( .A(n5833), .B(n5836), .S(n5911), .Z(n5838) );
  INV_X1 U7521 ( .A(n5834), .ZN(n5835) );
  NAND3_X1 U7522 ( .A1(n5836), .A2(n5835), .A3(n5877), .ZN(n5837) );
  NAND3_X1 U7523 ( .A1(n8613), .A2(n5838), .A3(n5837), .ZN(n5842) );
  MUX2_X1 U7524 ( .A(n5840), .B(n5839), .S(n5911), .Z(n5841) );
  OAI211_X1 U7525 ( .C1(n5843), .C2(n5842), .A(n9408), .B(n5841), .ZN(n5847)
         );
  MUX2_X1 U7526 ( .A(n5845), .B(n5844), .S(n5911), .Z(n5846) );
  NAND2_X1 U7527 ( .A1(n5849), .A2(n5853), .ZN(n9364) );
  INV_X1 U7528 ( .A(n5850), .ZN(n5851) );
  INV_X1 U7529 ( .A(n9363), .ZN(n9325) );
  MUX2_X1 U7530 ( .A(n5851), .B(n9325), .S(n5911), .Z(n5852) );
  NAND2_X1 U7531 ( .A1(n5921), .A2(n5853), .ZN(n5854) );
  MUX2_X1 U7532 ( .A(n5854), .B(n9327), .S(n5911), .Z(n5855) );
  OAI21_X1 U7533 ( .B1(n5869), .B2(n9329), .A(n9309), .ZN(n5867) );
  NOR2_X1 U7534 ( .A1(n9332), .A2(n5911), .ZN(n5860) );
  AND2_X1 U7535 ( .A1(n9489), .A2(n5860), .ZN(n5861) );
  AOI21_X1 U7536 ( .B1(n5877), .B2(n9280), .A(n5861), .ZN(n5863) );
  INV_X1 U7537 ( .A(n5861), .ZN(n5862) );
  OAI22_X1 U7538 ( .A1(n5863), .A2(n9290), .B1(n5862), .B2(n9313), .ZN(n5864)
         );
  INV_X1 U7539 ( .A(n5870), .ZN(n5871) );
  OAI211_X1 U7540 ( .C1(n5873), .C2(n5872), .A(n9292), .B(n5871), .ZN(n5875)
         );
  NAND3_X1 U7541 ( .A1(n5875), .A2(n5918), .A3(n5874), .ZN(n5876) );
  NAND4_X1 U7542 ( .A1(n5878), .A2(n5883), .A3(n5911), .A4(n5876), .ZN(n5882)
         );
  NAND4_X1 U7543 ( .A1(n5878), .A2(n5877), .A3(n5918), .A4(n5879), .ZN(n5881)
         );
  NAND2_X1 U7544 ( .A1(n5034), .A2(n5911), .ZN(n5880) );
  AOI21_X1 U7545 ( .B1(n9206), .B2(n5883), .A(n5911), .ZN(n5885) );
  MUX2_X1 U7546 ( .A(n5917), .B(n9206), .S(n5911), .Z(n5884) );
  INV_X1 U7547 ( .A(n9207), .ZN(n5886) );
  NAND2_X1 U7548 ( .A1(n5890), .A2(n5889), .ZN(n5891) );
  INV_X1 U7549 ( .A(n5892), .ZN(n5893) );
  INV_X1 U7550 ( .A(n5895), .ZN(n5896) );
  NOR2_X1 U7551 ( .A1(n5897), .A2(n5896), .ZN(n5899) );
  MUX2_X1 U7552 ( .A(n5899), .B(n5898), .S(n5911), .Z(n5903) );
  INV_X1 U7553 ( .A(n9452), .ZN(n9189) );
  NAND2_X1 U7554 ( .A1(n9189), .A2(n5911), .ZN(n5900) );
  AOI22_X1 U7555 ( .A1(n5900), .A2(n4441), .B1(n9198), .B2(n5911), .ZN(n5901)
         );
  NOR2_X1 U7556 ( .A1(n8826), .A2(n5911), .ZN(n5904) );
  MUX2_X1 U7557 ( .A(n5904), .B(n8826), .S(n9438), .Z(n5905) );
  NAND2_X1 U7558 ( .A1(n5910), .A2(n5909), .ZN(n5938) );
  INV_X1 U7559 ( .A(n5943), .ZN(n5942) );
  NAND2_X1 U7560 ( .A1(n9292), .A2(n5920), .ZN(n9311) );
  NAND2_X1 U7561 ( .A1(n5856), .A2(n5921), .ZN(n9347) );
  INV_X1 U7562 ( .A(n9388), .ZN(n9380) );
  NAND2_X1 U7563 ( .A1(n7594), .A2(n7597), .ZN(n8023) );
  NAND2_X1 U7564 ( .A1(n5786), .A2(n5925), .ZN(n7314) );
  NOR4_X1 U7565 ( .A1(n5924), .A2(n8023), .A3(n7317), .A4(n5926), .ZN(n5927)
         );
  NAND4_X1 U7566 ( .A1(n5927), .A2(n7785), .A3(n8065), .A4(n7527), .ZN(n5929)
         );
  NOR4_X1 U7567 ( .A1(n5929), .A2(n7988), .A3(n5928), .A4(n8509), .ZN(n5930)
         );
  NAND4_X1 U7568 ( .A1(n8184), .A2(n7970), .A3(n7797), .A4(n5930), .ZN(n5931)
         );
  NOR4_X1 U7569 ( .A1(n8622), .A2(n5932), .A3(n5931), .A4(n8551), .ZN(n5933)
         );
  NAND4_X1 U7570 ( .A1(n9357), .A2(n9380), .A3(n9408), .A4(n5933), .ZN(n5934)
         );
  NAND4_X1 U7571 ( .A1(n9254), .A2(n9278), .A3(n5935), .A4(n9297), .ZN(n5936)
         );
  NOR4_X1 U7572 ( .A1(n9208), .A2(n9228), .A3(n9242), .A4(n5936), .ZN(n5937)
         );
  XOR2_X1 U7573 ( .A(n7537), .B(n5939), .Z(n5940) );
  OAI22_X1 U7574 ( .A1(n5940), .A2(n5955), .B1(n7543), .B2(n7138), .ZN(n5941)
         );
  NAND3_X1 U7575 ( .A1(n5943), .A2(n7091), .A3(n7564), .ZN(n5960) );
  INV_X1 U7576 ( .A(n7091), .ZN(n8015) );
  INV_X1 U7577 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5944) );
  NAND2_X1 U7578 ( .A1(n5945), .A2(n5944), .ZN(n5946) );
  NAND2_X1 U7579 ( .A1(n5946), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5947) );
  NAND2_X1 U7580 ( .A1(n4537), .A2(n5948), .ZN(n5952) );
  OAI21_X1 U7581 ( .B1(n5952), .B2(P2_IR_REG_25__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5950) );
  MUX2_X1 U7582 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5950), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n5951) );
  NAND2_X1 U7583 ( .A1(n5952), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5953) );
  XNOR2_X1 U7584 ( .A(n5953), .B(P2_IR_REG_25__SCAN_IN), .ZN(n7122) );
  AND2_X1 U7585 ( .A1(n8193), .A2(n7122), .ZN(n5954) );
  NAND2_X1 U7586 ( .A1(n7135), .A2(n5954), .ZN(n7548) );
  NOR2_X1 U7587 ( .A1(n7545), .A2(P2_U3152), .ZN(n10385) );
  INV_X1 U7588 ( .A(n8847), .ZN(n5957) );
  INV_X1 U7589 ( .A(n5956), .ZN(n7140) );
  NAND4_X1 U7590 ( .A1(n10373), .A2(n5957), .A3(n9411), .A4(n7315), .ZN(n5958)
         );
  OAI211_X1 U7591 ( .C1(n7142), .C2(n8015), .A(n5958), .B(P2_B_REG_SCAN_IN), 
        .ZN(n5959) );
  NOR2_X4 U7592 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n6049) );
  NOR2_X2 U7593 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n5964) );
  INV_X2 U7594 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n6088) );
  NAND4_X1 U7595 ( .A1(n5964), .A2(n5963), .A3(n6088), .A4(n8279), .ZN(n5965)
         );
  INV_X2 U7596 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n6203) );
  NOR2_X1 U7597 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n5967) );
  NOR2_X1 U7598 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n5966) );
  AND2_X1 U7599 ( .A1(n5967), .A2(n5966), .ZN(n5969) );
  INV_X1 U7600 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5974) );
  XNOR2_X2 U7601 ( .A(n5975), .B(n5974), .ZN(n6531) );
  NAND2_X2 U7602 ( .A1(n4396), .A2(n4399), .ZN(n6090) );
  INV_X4 U7603 ( .A(n6090), .ZN(n6381) );
  NAND2_X1 U7604 ( .A1(n6995), .A2(n6381), .ZN(n5979) );
  NAND2_X1 U7605 ( .A1(n6049), .A2(n6050), .ZN(n6060) );
  NAND2_X1 U7606 ( .A1(n5976), .A2(n4504), .ZN(n5994) );
  OR2_X1 U7607 ( .A1(n5994), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n5997) );
  NAND2_X1 U7608 ( .A1(n5997), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5977) );
  XNOR2_X1 U7609 ( .A(n5977), .B(P1_IR_REG_10__SCAN_IN), .ZN(n7429) );
  AOI22_X1 U7610 ( .A1(n6246), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6245), .B2(
        n7429), .ZN(n5978) );
  XNOR2_X2 U7611 ( .A(n5983), .B(n5982), .ZN(n5989) );
  INV_X1 U7612 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5984) );
  INV_X2 U7613 ( .A(n6048), .ZN(n6389) );
  NAND2_X1 U7614 ( .A1(n6389), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5993) );
  AND2_X2 U7615 ( .A1(n5986), .A2(n10245), .ZN(n6266) );
  NAND2_X1 U7616 ( .A1(n6266), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5992) );
  AND2_X4 U7617 ( .A1(n6030), .A2(n5986), .ZN(n6307) );
  NAND2_X1 U7618 ( .A1(n6003), .A2(n8418), .ZN(n5988) );
  NAND2_X1 U7619 ( .A1(n6143), .A2(n5988), .ZN(n8579) );
  INV_X1 U7620 ( .A(n8579), .ZN(n8041) );
  NAND2_X1 U7621 ( .A1(n6307), .A2(n8041), .ZN(n5991) );
  AND2_X4 U7622 ( .A1(n10245), .A2(n5989), .ZN(n6390) );
  NAND2_X1 U7623 ( .A1(n6390), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5990) );
  NAND2_X1 U7624 ( .A1(n10196), .A2(n7950), .ZN(n6421) );
  NAND2_X1 U7625 ( .A1(n6989), .A2(n6381), .ZN(n6000) );
  NAND2_X1 U7626 ( .A1(n5994), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5996) );
  MUX2_X1 U7627 ( .A(n5996), .B(P1_IR_REG_31__SCAN_IN), .S(n5995), .Z(n5998)
         );
  AOI22_X1 U7628 ( .A1(n6246), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n6245), .B2(
        n7409), .ZN(n5999) );
  NAND2_X1 U7629 ( .A1(n6266), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6008) );
  NAND2_X1 U7630 ( .A1(n6389), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6007) );
  INV_X1 U7631 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n6002) );
  INV_X1 U7632 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n6001) );
  OAI21_X1 U7633 ( .B1(n6108), .B2(n6002), .A(n6001), .ZN(n6004) );
  AND2_X1 U7634 ( .A1(n6004), .A2(n6003), .ZN(n8532) );
  NAND2_X1 U7635 ( .A1(n6307), .A2(n8532), .ZN(n6006) );
  NAND2_X1 U7636 ( .A1(n6390), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n6005) );
  NAND4_X1 U7637 ( .A1(n6008), .A2(n6007), .A3(n6006), .A4(n6005), .ZN(n9773)
         );
  INV_X1 U7638 ( .A(n9773), .ZN(n8114) );
  NAND2_X1 U7639 ( .A1(n10201), .A2(n8114), .ZN(n8031) );
  AND2_X1 U7640 ( .A1(n6421), .A2(n8031), .ZN(n6648) );
  INV_X1 U7641 ( .A(n6649), .ZN(n6009) );
  NOR2_X1 U7642 ( .A1(n6648), .A2(n6009), .ZN(n6457) );
  NAND2_X1 U7643 ( .A1(n6960), .A2(n6381), .ZN(n6012) );
  NAND2_X1 U7644 ( .A1(n6085), .A2(n6088), .ZN(n6100) );
  OAI21_X1 U7645 ( .B1(n4434), .B2(P1_IR_REG_7__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6010) );
  AOI22_X1 U7646 ( .A1(n6246), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n6245), .B2(
        n7177), .ZN(n6011) );
  INV_X1 U7647 ( .A(n6048), .ZN(n6091) );
  NAND2_X1 U7648 ( .A1(n6091), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6016) );
  NAND2_X1 U7649 ( .A1(n6266), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6015) );
  XNOR2_X1 U7650 ( .A(n6108), .B(P1_REG3_REG_8__SCAN_IN), .ZN(n8111) );
  NAND2_X1 U7651 ( .A1(n6307), .A2(n8111), .ZN(n6014) );
  NAND2_X1 U7652 ( .A1(n6390), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n6013) );
  NAND2_X1 U7653 ( .A1(n10206), .A2(n8530), .ZN(n6645) );
  NAND2_X1 U7654 ( .A1(n6188), .A2(n6186), .ZN(n6200) );
  INV_X1 U7655 ( .A(n6200), .ZN(n6017) );
  NAND3_X1 U7656 ( .A1(n6018), .A2(n6017), .A3(n6203), .ZN(n6020) );
  AND2_X1 U7657 ( .A1(n6164), .A2(n6168), .ZN(n6154) );
  INV_X1 U7658 ( .A(n6154), .ZN(n6019) );
  NOR2_X1 U7659 ( .A1(n6020), .A2(n6019), .ZN(n6025) );
  INV_X1 U7660 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n6021) );
  AND2_X1 U7661 ( .A1(n6025), .A2(n6021), .ZN(n6022) );
  NAND2_X1 U7662 ( .A1(n6022), .A2(n6165), .ZN(n6028) );
  INV_X1 U7663 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n6443) );
  NAND2_X1 U7664 ( .A1(n6444), .A2(n6443), .ZN(n6023) );
  NAND2_X1 U7665 ( .A1(n6409), .A2(n6408), .ZN(n6410) );
  NAND2_X1 U7666 ( .A1(n6410), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6024) );
  NAND2_X1 U7667 ( .A1(n6025), .A2(n6165), .ZN(n6026) );
  NAND2_X1 U7668 ( .A1(n6026), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6027) );
  MUX2_X1 U7669 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6027), .S(
        P1_IR_REG_19__SCAN_IN), .Z(n6029) );
  NAND2_X1 U7670 ( .A1(n6029), .A2(n6028), .ZN(n9962) );
  INV_X1 U7671 ( .A(n9962), .ZN(n10310) );
  NOR3_X1 U7672 ( .A1(n6457), .A2(n4975), .A3(n7368), .ZN(n6153) );
  NAND2_X1 U7673 ( .A1(n6266), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6034) );
  NAND2_X1 U7674 ( .A1(n6390), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n6032) );
  NAND2_X1 U7675 ( .A1(n6126), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6031) );
  INV_X1 U7676 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n6035) );
  INV_X1 U7677 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6954) );
  OR2_X1 U7678 ( .A1(n6382), .A2(n6954), .ZN(n6038) );
  INV_X1 U7679 ( .A(n6036), .ZN(n6985) );
  NAND2_X1 U7680 ( .A1(n6307), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n6042) );
  NAND2_X1 U7681 ( .A1(n6126), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6039) );
  INV_X1 U7682 ( .A(SI_0_), .ZN(n6043) );
  NOR2_X1 U7683 ( .A1(n6964), .A2(n6043), .ZN(n6045) );
  INV_X1 U7684 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n6044) );
  XNOR2_X1 U7685 ( .A(n6045), .B(n6044), .ZN(n10252) );
  MUX2_X1 U7686 ( .A(P1_IR_REG_0__SCAN_IN), .B(n10252), .S(n6977), .Z(n7422)
         );
  NOR2_X1 U7687 ( .A1(n4575), .A2(n7372), .ZN(n7376) );
  NAND2_X1 U7688 ( .A1(n7463), .A2(n4401), .ZN(n6046) );
  NAND2_X1 U7689 ( .A1(n6047), .A2(n6046), .ZN(n7461) );
  NAND2_X1 U7690 ( .A1(n6266), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6579) );
  NAND2_X1 U7691 ( .A1(n6307), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n6578) );
  NAND2_X1 U7692 ( .A1(n6390), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n6577) );
  NAND2_X1 U7693 ( .A1(n6091), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6576) );
  OR2_X1 U7694 ( .A1(n6090), .A2(n6988), .ZN(n6053) );
  OR2_X1 U7695 ( .A1(n6382), .A2(n6958), .ZN(n6052) );
  XNOR2_X1 U7696 ( .A(n6580), .B(n7469), .ZN(n7464) );
  INV_X1 U7697 ( .A(n7469), .ZN(n7506) );
  NOR2_X1 U7698 ( .A1(n6580), .A2(n7506), .ZN(n6054) );
  INV_X1 U7699 ( .A(n7448), .ZN(n6536) );
  NAND2_X1 U7700 ( .A1(n6266), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6058) );
  NAND2_X1 U7701 ( .A1(n6390), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n6057) );
  NAND2_X1 U7702 ( .A1(n6307), .A2(n8466), .ZN(n6056) );
  NAND2_X1 U7703 ( .A1(n6126), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6055) );
  INV_X1 U7704 ( .A(n6059), .ZN(n6967) );
  OR2_X1 U7705 ( .A1(n6090), .A2(n6967), .ZN(n6064) );
  OR2_X1 U7706 ( .A1(n6382), .A2(n6944), .ZN(n6063) );
  NAND2_X1 U7707 ( .A1(n6060), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6061) );
  XNOR2_X1 U7708 ( .A(n6061), .B(P1_IR_REG_3__SCAN_IN), .ZN(n7008) );
  NAND2_X1 U7709 ( .A1(n6245), .A2(n7008), .ZN(n6062) );
  NAND2_X1 U7710 ( .A1(n9779), .A2(n7458), .ZN(n6494) );
  NAND2_X1 U7711 ( .A1(n7702), .A2(n6494), .ZN(n7447) );
  NAND2_X1 U7712 ( .A1(n6266), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6069) );
  NAND2_X1 U7713 ( .A1(n6091), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6068) );
  OAI21_X1 U7714 ( .B1(P1_REG3_REG_3__SCAN_IN), .B2(P1_REG3_REG_4__SCAN_IN), 
        .A(n6079), .ZN(n6065) );
  INV_X1 U7715 ( .A(n6065), .ZN(n7710) );
  NAND2_X1 U7716 ( .A1(n6307), .A2(n7710), .ZN(n6067) );
  NAND2_X1 U7717 ( .A1(n6390), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n6066) );
  NAND2_X1 U7718 ( .A1(n6070), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6072) );
  INV_X1 U7719 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n6071) );
  XNOR2_X1 U7720 ( .A(n6072), .B(n6071), .ZN(n7009) );
  INV_X1 U7721 ( .A(n6073), .ZN(n6970) );
  OR2_X1 U7722 ( .A1(n6090), .A2(n6970), .ZN(n6075) );
  OR2_X1 U7723 ( .A1(n6382), .A2(n6943), .ZN(n6074) );
  OAI211_X1 U7724 ( .C1(n6977), .C2(n7009), .A(n6075), .B(n6074), .ZN(n7711)
         );
  XNOR2_X1 U7725 ( .A(n7711), .B(n9777), .ZN(n7698) );
  NAND2_X1 U7726 ( .A1(n7484), .A2(n7711), .ZN(n6496) );
  NAND2_X1 U7727 ( .A1(n6266), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6084) );
  NAND2_X1 U7728 ( .A1(n6091), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6083) );
  INV_X1 U7729 ( .A(n6077), .ZN(n6093) );
  INV_X1 U7730 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n6078) );
  NAND2_X1 U7731 ( .A1(n6079), .A2(n6078), .ZN(n6080) );
  AND2_X1 U7732 ( .A1(n6093), .A2(n6080), .ZN(n7850) );
  NAND2_X1 U7733 ( .A1(n6307), .A2(n7850), .ZN(n6082) );
  NAND2_X1 U7734 ( .A1(n6390), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n6081) );
  NAND4_X2 U7735 ( .A1(n6084), .A2(n6083), .A3(n6082), .A4(n6081), .ZN(n8209)
         );
  INV_X1 U7736 ( .A(n6085), .ZN(n6086) );
  NAND2_X1 U7737 ( .A1(n6086), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6087) );
  INV_X1 U7738 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6959) );
  INV_X1 U7739 ( .A(n6089), .ZN(n6991) );
  NAND2_X1 U7740 ( .A1(n6091), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6098) );
  NAND2_X1 U7741 ( .A1(n6266), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6097) );
  INV_X1 U7742 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6092) );
  NAND2_X1 U7743 ( .A1(n6093), .A2(n6092), .ZN(n6094) );
  AND2_X1 U7744 ( .A1(n6106), .A2(n6094), .ZN(n8212) );
  NAND2_X1 U7745 ( .A1(n6307), .A2(n8212), .ZN(n6096) );
  NAND2_X1 U7746 ( .A1(n6390), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n6095) );
  NAND2_X1 U7747 ( .A1(n6099), .A2(n6381), .ZN(n6105) );
  NAND2_X1 U7748 ( .A1(n6100), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6101) );
  MUX2_X1 U7749 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6101), .S(
        P1_IR_REG_6__SCAN_IN), .Z(n6102) );
  NAND2_X1 U7750 ( .A1(n6245), .A2(n7046), .ZN(n6104) );
  INV_X1 U7751 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6945) );
  OR2_X1 U7752 ( .A1(n6382), .A2(n6945), .ZN(n6103) );
  AND3_X2 U7753 ( .A1(n6105), .A2(n6104), .A3(n6103), .ZN(n10345) );
  NAND2_X1 U7754 ( .A1(n9776), .A2(n10345), .ZN(n6492) );
  AOI21_X1 U7755 ( .B1(n6119), .B2(n7813), .A(n4952), .ZN(n6116) );
  NAND2_X1 U7756 ( .A1(n4380), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6112) );
  NAND2_X1 U7757 ( .A1(n6389), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6111) );
  INV_X1 U7758 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n8264) );
  NAND2_X1 U7759 ( .A1(n6106), .A2(n8264), .ZN(n6107) );
  AND2_X1 U7760 ( .A1(n6108), .A2(n6107), .ZN(n7753) );
  NAND2_X1 U7761 ( .A1(n6307), .A2(n7753), .ZN(n6110) );
  NAND2_X1 U7762 ( .A1(n6390), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n6109) );
  NAND2_X1 U7763 ( .A1(n6962), .A2(n6381), .ZN(n6115) );
  NAND2_X1 U7764 ( .A1(n4434), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6113) );
  AOI22_X1 U7765 ( .A1(n6246), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n6245), .B2(
        n7080), .ZN(n6114) );
  INV_X1 U7766 ( .A(n6643), .ZN(n6118) );
  NAND2_X1 U7767 ( .A1(n7748), .A2(n9775), .ZN(n6543) );
  OAI21_X1 U7768 ( .B1(n6116), .B2(n6118), .A(n6543), .ZN(n6152) );
  INV_X1 U7769 ( .A(n6497), .ZN(n6117) );
  NOR3_X1 U7770 ( .A1(n6119), .A2(n6118), .A3(n6117), .ZN(n6150) );
  OR2_X1 U7771 ( .A1(n10201), .A2(n8114), .ZN(n6647) );
  NAND2_X1 U7772 ( .A1(n6649), .A2(n6647), .ZN(n6122) );
  INV_X1 U7773 ( .A(n6122), .ZN(n6120) );
  NAND4_X1 U7774 ( .A1(n6120), .A2(n6646), .A3(n6543), .A4(n7368), .ZN(n6149)
         );
  INV_X1 U7775 ( .A(n6646), .ZN(n6121) );
  NOR2_X1 U7776 ( .A1(n6122), .A2(n6121), .ZN(n6458) );
  NOR3_X1 U7777 ( .A1(n6457), .A2(n6458), .A3(n7368), .ZN(n6138) );
  AOI211_X1 U7778 ( .C1(n6645), .C2(n8031), .A(n4791), .B(n6122), .ZN(n6137)
         );
  NAND2_X1 U7779 ( .A1(n7094), .A2(n6381), .ZN(n6125) );
  NOR2_X1 U7780 ( .A1(n6165), .A2(n5984), .ZN(n6123) );
  XNOR2_X1 U7781 ( .A(n6123), .B(n6164), .ZN(n7858) );
  AOI22_X1 U7782 ( .A1(n6246), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n6245), .B2(
        n7858), .ZN(n6124) );
  NAND2_X1 U7783 ( .A1(n4380), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n6135) );
  NAND2_X1 U7784 ( .A1(n6385), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n6134) );
  AND2_X1 U7785 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_REG3_REG_12__SCAN_IN), 
        .ZN(n6127) );
  INV_X1 U7786 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n6130) );
  INV_X1 U7787 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n6129) );
  OAI21_X1 U7788 ( .B1(n6143), .B2(n6130), .A(n6129), .ZN(n6131) );
  AND2_X1 U7789 ( .A1(n6171), .A2(n6131), .ZN(n8593) );
  NAND2_X1 U7790 ( .A1(n6307), .A2(n8593), .ZN(n6133) );
  NAND2_X1 U7791 ( .A1(n6390), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n6132) );
  NAND4_X1 U7792 ( .A1(n6135), .A2(n6134), .A3(n6133), .A4(n6132), .ZN(n9770)
         );
  NAND2_X1 U7793 ( .A1(n8590), .A2(n9770), .ZN(n6419) );
  INV_X1 U7794 ( .A(n6419), .ZN(n8596) );
  OAI21_X1 U7795 ( .B1(n4791), .B2(n6421), .A(n8597), .ZN(n6136) );
  NAND2_X1 U7796 ( .A1(n7022), .A2(n6381), .ZN(n6142) );
  NAND2_X1 U7797 ( .A1(n6139), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6140) );
  XNOR2_X1 U7798 ( .A(n6140), .B(P1_IR_REG_11__SCAN_IN), .ZN(n7719) );
  AOI22_X1 U7799 ( .A1(n6246), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n6245), .B2(
        n7719), .ZN(n6141) );
  NAND2_X1 U7800 ( .A1(n6385), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n6147) );
  NAND2_X1 U7801 ( .A1(n4380), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6146) );
  XNOR2_X1 U7802 ( .A(n6143), .B(P1_REG3_REG_11__SCAN_IN), .ZN(n8545) );
  NAND2_X1 U7803 ( .A1(n6307), .A2(n8545), .ZN(n6145) );
  NAND2_X1 U7804 ( .A1(n6390), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n6144) );
  NAND4_X1 U7805 ( .A1(n6147), .A2(n6146), .A3(n6145), .A4(n6144), .ZN(n9771)
         );
  XNOR2_X1 U7806 ( .A(n7958), .B(n9771), .ZN(n6420) );
  OAI211_X1 U7807 ( .C1(n6150), .C2(n6149), .A(n6148), .B(n6420), .ZN(n6151)
         );
  AOI21_X1 U7808 ( .B1(n6153), .B2(n6152), .A(n6151), .ZN(n6185) );
  NAND2_X1 U7809 ( .A1(n7113), .A2(n6381), .ZN(n6157) );
  NAND2_X1 U7810 ( .A1(n6165), .A2(n6154), .ZN(n6155) );
  NAND2_X1 U7811 ( .A1(n6155), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6202) );
  XNOR2_X1 U7812 ( .A(n6202), .B(P1_IR_REG_14__SCAN_IN), .ZN(n8709) );
  AOI22_X1 U7813 ( .A1(n6246), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n6245), .B2(
        n8709), .ZN(n6156) );
  NAND2_X1 U7814 ( .A1(n6266), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n6163) );
  NAND2_X1 U7815 ( .A1(n6390), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n6162) );
  INV_X1 U7816 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n8630) );
  NAND2_X1 U7817 ( .A1(n6173), .A2(n8630), .ZN(n6159) );
  AND2_X1 U7818 ( .A1(n6194), .A2(n6159), .ZN(n10065) );
  NAND2_X1 U7819 ( .A1(n6307), .A2(n10065), .ZN(n6161) );
  NAND2_X1 U7820 ( .A1(n6385), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n6160) );
  NAND4_X1 U7821 ( .A1(n6163), .A2(n6162), .A3(n6161), .A4(n6160), .ZN(n10037)
         );
  INV_X1 U7822 ( .A(n10037), .ZN(n6428) );
  NAND2_X1 U7823 ( .A1(n10174), .A2(n6428), .ZN(n6180) );
  NAND2_X1 U7824 ( .A1(n7109), .A2(n6381), .ZN(n6170) );
  AND2_X1 U7825 ( .A1(n6165), .A2(n6164), .ZN(n6166) );
  NOR2_X1 U7826 ( .A1(n6166), .A2(n5984), .ZN(n6167) );
  XNOR2_X1 U7827 ( .A(n6168), .B(n6167), .ZN(n8632) );
  AOI22_X1 U7828 ( .A1(n6246), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n6245), .B2(
        n8632), .ZN(n6169) );
  NAND2_X1 U7829 ( .A1(n4380), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n6177) );
  NAND2_X1 U7830 ( .A1(n6385), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n6176) );
  INV_X1 U7831 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n8263) );
  NAND2_X1 U7832 ( .A1(n6171), .A2(n8263), .ZN(n6172) );
  AND2_X1 U7833 ( .A1(n6173), .A2(n6172), .ZN(n9710) );
  NAND2_X1 U7834 ( .A1(n6307), .A2(n9710), .ZN(n6175) );
  NAND2_X1 U7835 ( .A1(n6390), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n6174) );
  NAND4_X1 U7836 ( .A1(n6177), .A2(n6176), .A3(n6175), .A4(n6174), .ZN(n10058)
         );
  INV_X1 U7837 ( .A(n10058), .ZN(n6607) );
  NAND2_X1 U7838 ( .A1(n10178), .A2(n6607), .ZN(n6654) );
  NAND2_X1 U7839 ( .A1(n6180), .A2(n6654), .ZN(n6482) );
  INV_X1 U7840 ( .A(n9771), .ZN(n8589) );
  NAND2_X1 U7841 ( .A1(n7958), .A2(n8589), .ZN(n6651) );
  NAND2_X1 U7842 ( .A1(n8597), .A2(n6651), .ZN(n6456) );
  AND2_X1 U7843 ( .A1(n6456), .A2(n6419), .ZN(n6178) );
  OR2_X1 U7844 ( .A1(n6482), .A2(n6178), .ZN(n6179) );
  OR2_X1 U7845 ( .A1(n10174), .A2(n6428), .ZN(n6656) );
  INV_X1 U7846 ( .A(n10178), .ZN(n9707) );
  NAND2_X1 U7847 ( .A1(n9707), .A2(n10058), .ZN(n6418) );
  NAND2_X1 U7848 ( .A1(n6656), .A2(n6418), .ZN(n6181) );
  NAND2_X1 U7849 ( .A1(n6181), .A2(n6180), .ZN(n6182) );
  OR2_X1 U7850 ( .A1(n7958), .A2(n8589), .ZN(n6652) );
  NAND2_X1 U7851 ( .A1(n6419), .A2(n6652), .ZN(n6183) );
  NAND2_X1 U7852 ( .A1(n6183), .A2(n8597), .ZN(n6184) );
  NAND2_X1 U7853 ( .A1(n7116), .A2(n6381), .ZN(n6192) );
  NAND2_X1 U7854 ( .A1(n6202), .A2(n6186), .ZN(n6187) );
  NAND2_X1 U7855 ( .A1(n6187), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6189) );
  XNOR2_X1 U7856 ( .A(n6189), .B(n6188), .ZN(n9802) );
  INV_X1 U7857 ( .A(n9802), .ZN(n6190) );
  AOI22_X1 U7858 ( .A1(n6246), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n6245), .B2(
        n6190), .ZN(n6191) );
  NAND2_X1 U7859 ( .A1(n4380), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n6199) );
  NAND2_X1 U7860 ( .A1(n6390), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n6198) );
  INV_X1 U7861 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n6193) );
  NAND2_X1 U7862 ( .A1(n6194), .A2(n6193), .ZN(n6195) );
  AND2_X1 U7863 ( .A1(n6208), .A2(n6195), .ZN(n10045) );
  NAND2_X1 U7864 ( .A1(n6307), .A2(n10045), .ZN(n6197) );
  NAND2_X1 U7865 ( .A1(n6389), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n6196) );
  NAND2_X1 U7866 ( .A1(n10168), .A2(n9612), .ZN(n6658) );
  NAND2_X1 U7867 ( .A1(n7300), .A2(n6381), .ZN(n6205) );
  NAND2_X1 U7868 ( .A1(n6200), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6201) );
  NAND2_X1 U7869 ( .A1(n6202), .A2(n6201), .ZN(n6215) );
  XNOR2_X1 U7870 ( .A(n6215), .B(n6203), .ZN(n8713) );
  AOI22_X1 U7871 ( .A1(n6246), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n6245), .B2(
        n8713), .ZN(n6204) );
  NAND2_X1 U7872 ( .A1(n4380), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n6213) );
  NAND2_X1 U7873 ( .A1(n6385), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n6212) );
  INV_X1 U7874 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n6207) );
  NAND2_X1 U7875 ( .A1(n6208), .A2(n6207), .ZN(n6209) );
  AND2_X1 U7876 ( .A1(n6220), .A2(n6209), .ZN(n10023) );
  NAND2_X1 U7877 ( .A1(n6307), .A2(n10023), .ZN(n6211) );
  NAND2_X1 U7878 ( .A1(n6390), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n6210) );
  NAND2_X1 U7879 ( .A1(n10164), .A2(n9759), .ZN(n6661) );
  INV_X1 U7880 ( .A(n10029), .ZN(n10017) );
  INV_X1 U7881 ( .A(n6658), .ZN(n6481) );
  MUX2_X1 U7882 ( .A(n6481), .B(n4959), .S(n7368), .Z(n6214) );
  NOR2_X1 U7883 ( .A1(n10017), .A2(n6214), .ZN(n6227) );
  INV_X1 U7884 ( .A(n6464), .ZN(n6662) );
  INV_X1 U7885 ( .A(n6661), .ZN(n6455) );
  MUX2_X1 U7886 ( .A(n6662), .B(n6455), .S(n7368), .Z(n6226) );
  NAND2_X1 U7887 ( .A1(n7296), .A2(n6381), .ZN(n6218) );
  OR2_X1 U7888 ( .A1(n6215), .A2(P1_IR_REG_16__SCAN_IN), .ZN(n6216) );
  NAND2_X1 U7889 ( .A1(n6216), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6230) );
  XNOR2_X1 U7890 ( .A(n6230), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9829) );
  AOI22_X1 U7891 ( .A1(n6246), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n6245), .B2(
        n9829), .ZN(n6217) );
  NAND2_X1 U7892 ( .A1(n4380), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n6225) );
  NAND2_X1 U7893 ( .A1(n6390), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n6224) );
  INV_X1 U7894 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n6219) );
  NAND2_X1 U7895 ( .A1(n6220), .A2(n6219), .ZN(n6221) );
  AND2_X1 U7896 ( .A1(n6238), .A2(n6221), .ZN(n10009) );
  NAND2_X1 U7897 ( .A1(n6307), .A2(n10009), .ZN(n6223) );
  NAND2_X1 U7898 ( .A1(n6389), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n6222) );
  NAND4_X1 U7899 ( .A1(n6225), .A2(n6224), .A3(n6223), .A4(n6222), .ZN(n10019)
         );
  INV_X1 U7900 ( .A(n10019), .ZN(n9669) );
  OR2_X1 U7901 ( .A1(n10158), .A2(n9669), .ZN(n9985) );
  NAND2_X1 U7902 ( .A1(n10158), .A2(n9669), .ZN(n9984) );
  NAND2_X1 U7903 ( .A1(n9985), .A2(n9984), .ZN(n10013) );
  NAND2_X1 U7904 ( .A1(n7439), .A2(n6381), .ZN(n6234) );
  INV_X1 U7905 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n6229) );
  NAND2_X1 U7906 ( .A1(n6230), .A2(n6229), .ZN(n6231) );
  NAND2_X1 U7907 ( .A1(n6231), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6232) );
  XNOR2_X1 U7908 ( .A(n6232), .B(P1_IR_REG_18__SCAN_IN), .ZN(n10293) );
  AOI22_X1 U7909 ( .A1(n6246), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n10293), 
        .B2(n6245), .ZN(n6233) );
  NAND2_X1 U7910 ( .A1(n4380), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n6236) );
  NAND2_X1 U7911 ( .A1(n6385), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n6235) );
  AND2_X1 U7912 ( .A1(n6236), .A2(n6235), .ZN(n6242) );
  INV_X1 U7913 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n6237) );
  NAND2_X1 U7914 ( .A1(n6238), .A2(n6237), .ZN(n6239) );
  NAND2_X1 U7915 ( .A1(n6249), .A2(n6239), .ZN(n9993) );
  OR2_X1 U7916 ( .A1(n9993), .A2(n6371), .ZN(n6241) );
  NAND2_X1 U7917 ( .A1(n6390), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n6240) );
  NAND2_X1 U7918 ( .A1(n10154), .A2(n6714), .ZN(n6664) );
  NAND2_X1 U7919 ( .A1(n6664), .A2(n9984), .ZN(n6663) );
  OR2_X1 U7920 ( .A1(n10154), .A2(n6714), .ZN(n6417) );
  NAND2_X1 U7921 ( .A1(n6417), .A2(n9985), .ZN(n6665) );
  MUX2_X1 U7922 ( .A(n6663), .B(n6665), .S(n7368), .Z(n6243) );
  NAND2_X1 U7923 ( .A1(n7536), .A2(n6381), .ZN(n6248) );
  AOI22_X1 U7924 ( .A1(n6246), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n10310), 
        .B2(n6245), .ZN(n6247) );
  INV_X1 U7925 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n8343) );
  NAND2_X1 U7926 ( .A1(n6249), .A2(n8343), .ZN(n6250) );
  NAND2_X1 U7927 ( .A1(n6256), .A2(n6250), .ZN(n9972) );
  AOI22_X1 U7928 ( .A1(n6389), .A2(P1_REG1_REG_19__SCAN_IN), .B1(n4380), .B2(
        P1_REG2_REG_19__SCAN_IN), .ZN(n6252) );
  NAND2_X1 U7929 ( .A1(n6390), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n6251) );
  OAI211_X1 U7930 ( .C1(n9972), .C2(n6371), .A(n6252), .B(n6251), .ZN(n9988)
         );
  INV_X1 U7931 ( .A(n9988), .ZN(n9729) );
  OR2_X1 U7932 ( .A1(n10148), .A2(n9729), .ZN(n6415) );
  NAND2_X1 U7933 ( .A1(n7624), .A2(n6381), .ZN(n6254) );
  OR2_X1 U7934 ( .A1(n4525), .A2(n7627), .ZN(n6253) );
  INV_X1 U7935 ( .A(n6385), .ZN(n6260) );
  INV_X1 U7936 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n8413) );
  INV_X1 U7937 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n6255) );
  NAND2_X1 U7938 ( .A1(n6256), .A2(n6255), .ZN(n6257) );
  NAND2_X1 U7939 ( .A1(n6264), .A2(n6257), .ZN(n9964) );
  OR2_X1 U7940 ( .A1(n9964), .A2(n6371), .ZN(n6259) );
  AOI22_X1 U7941 ( .A1(n6390), .A2(P1_REG0_REG_20__SCAN_IN), .B1(n4380), .B2(
        P1_REG2_REG_20__SCAN_IN), .ZN(n6258) );
  OAI211_X1 U7942 ( .C1(n6260), .C2(n8413), .A(n6259), .B(n6258), .ZN(n9979)
         );
  INV_X1 U7943 ( .A(n9979), .ZN(n9953) );
  AND2_X1 U7944 ( .A1(n10144), .A2(n9953), .ZN(n6668) );
  INV_X1 U7945 ( .A(n6668), .ZN(n6416) );
  NAND2_X1 U7946 ( .A1(n10148), .A2(n9729), .ZN(n6666) );
  NAND2_X1 U7947 ( .A1(n6666), .A2(n6664), .ZN(n6469) );
  AND2_X1 U7948 ( .A1(n6667), .A2(n6415), .ZN(n6467) );
  NAND2_X1 U7949 ( .A1(n6261), .A2(n6381), .ZN(n6263) );
  OR2_X1 U7950 ( .A1(n4525), .A2(n7745), .ZN(n6262) );
  INV_X1 U7951 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n9642) );
  NAND2_X1 U7952 ( .A1(n6264), .A2(n9642), .ZN(n6265) );
  NAND2_X1 U7953 ( .A1(n6275), .A2(n6265), .ZN(n9943) );
  OR2_X1 U7954 ( .A1(n9943), .A2(n6371), .ZN(n6271) );
  INV_X1 U7955 ( .A(n6266), .ZN(n6364) );
  INV_X1 U7956 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n9944) );
  NAND2_X1 U7957 ( .A1(n6390), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n6268) );
  NAND2_X1 U7958 ( .A1(n6389), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n6267) );
  OAI211_X1 U7959 ( .C1(n6364), .C2(n9944), .A(n6268), .B(n6267), .ZN(n6269)
         );
  INV_X1 U7960 ( .A(n6269), .ZN(n6270) );
  NAND2_X1 U7961 ( .A1(n7891), .A2(n6381), .ZN(n6273) );
  OR2_X1 U7962 ( .A1(n4525), .A2(n8379), .ZN(n6272) );
  INV_X1 U7963 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n6274) );
  NAND2_X1 U7964 ( .A1(n6275), .A2(n6274), .ZN(n6276) );
  NAND2_X1 U7965 ( .A1(n6304), .A2(n6276), .ZN(n9717) );
  OR2_X1 U7966 ( .A1(n9717), .A2(n6371), .ZN(n6282) );
  INV_X1 U7967 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n6279) );
  NAND2_X1 U7968 ( .A1(n6389), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n6278) );
  NAND2_X1 U7969 ( .A1(n4380), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n6277) );
  OAI211_X1 U7970 ( .C1(n6279), .C2(n6388), .A(n6278), .B(n6277), .ZN(n6280)
         );
  INV_X1 U7971 ( .A(n6280), .ZN(n6281) );
  NAND2_X1 U7972 ( .A1(n6669), .A2(n6468), .ZN(n6283) );
  NAND2_X1 U7973 ( .A1(n9934), .A2(n9951), .ZN(n6670) );
  OAI21_X1 U7974 ( .B1(n6284), .B2(n6283), .A(n6670), .ZN(n6291) );
  INV_X1 U7975 ( .A(n6468), .ZN(n6285) );
  NOR2_X1 U7976 ( .A1(n6286), .A2(n6285), .ZN(n6289) );
  NAND2_X1 U7977 ( .A1(n6468), .A2(n6668), .ZN(n6287) );
  AND2_X1 U7978 ( .A1(n6287), .A2(n9912), .ZN(n6288) );
  NAND2_X1 U7979 ( .A1(n6288), .A2(n6670), .ZN(n6473) );
  OAI21_X1 U7980 ( .B1(n6289), .B2(n6473), .A(n6669), .ZN(n6290) );
  OR2_X1 U7981 ( .A1(n4525), .A2(n8134), .ZN(n6292) );
  INV_X1 U7982 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n8331) );
  INV_X1 U7983 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n6294) );
  NAND2_X1 U7984 ( .A1(n6306), .A2(n6294), .ZN(n6295) );
  NAND2_X1 U7985 ( .A1(n6317), .A2(n6295), .ZN(n9686) );
  INV_X1 U7986 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n6298) );
  NAND2_X1 U7987 ( .A1(n4380), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n6297) );
  NAND2_X1 U7988 ( .A1(n6389), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n6296) );
  OAI211_X1 U7989 ( .C1(n6388), .C2(n6298), .A(n6297), .B(n6296), .ZN(n6299)
         );
  INV_X1 U7990 ( .A(n6299), .ZN(n6300) );
  INV_X1 U7991 ( .A(n9919), .ZN(n9652) );
  INV_X1 U7992 ( .A(n6677), .ZN(n6314) );
  NAND2_X1 U7993 ( .A1(n10121), .A2(n9652), .ZN(n6676) );
  NAND2_X1 U7994 ( .A1(n8018), .A2(n6381), .ZN(n6303) );
  OR2_X1 U7995 ( .A1(n4525), .A2(n8022), .ZN(n6302) );
  NAND2_X1 U7996 ( .A1(n6304), .A2(n8331), .ZN(n6305) );
  AND2_X1 U7997 ( .A1(n6306), .A2(n6305), .ZN(n9908) );
  NAND2_X1 U7998 ( .A1(n9908), .A2(n6307), .ZN(n6312) );
  INV_X1 U7999 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n8262) );
  NAND2_X1 U8000 ( .A1(n6390), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n6309) );
  NAND2_X1 U8001 ( .A1(n6385), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n6308) );
  OAI211_X1 U8002 ( .C1(n6364), .C2(n8262), .A(n6309), .B(n6308), .ZN(n6310)
         );
  INV_X1 U8003 ( .A(n6310), .ZN(n6311) );
  NAND2_X1 U8004 ( .A1(n10126), .A2(n9720), .ZN(n6414) );
  NAND2_X1 U8005 ( .A1(n6676), .A2(n6414), .ZN(n6502) );
  INV_X1 U8006 ( .A(n6675), .ZN(n6313) );
  NOR3_X1 U8007 ( .A1(n6314), .A2(n6502), .A3(n6313), .ZN(n6339) );
  OR2_X1 U8008 ( .A1(n4525), .A2(n8520), .ZN(n6315) );
  INV_X1 U8009 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n9651) );
  NAND2_X1 U8010 ( .A1(n6317), .A2(n9651), .ZN(n6318) );
  NAND2_X1 U8011 ( .A1(n6330), .A2(n6318), .ZN(n9650) );
  INV_X1 U8012 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n6321) );
  NAND2_X1 U8013 ( .A1(n4380), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n6320) );
  NAND2_X1 U8014 ( .A1(n6385), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n6319) );
  OAI211_X1 U8015 ( .C1(n6321), .C2(n6388), .A(n6320), .B(n6319), .ZN(n6322)
         );
  INV_X1 U8016 ( .A(n6322), .ZN(n6323) );
  NAND2_X1 U8017 ( .A1(n6502), .A2(n6677), .ZN(n6325) );
  NAND2_X1 U8018 ( .A1(n6679), .A2(n6325), .ZN(n6535) );
  INV_X1 U8019 ( .A(n6676), .ZN(n6326) );
  AND2_X1 U8020 ( .A1(n9869), .A2(n6677), .ZN(n6504) );
  OAI21_X1 U8021 ( .B1(n6326), .B2(n6675), .A(n6504), .ZN(n6327) );
  MUX2_X1 U8022 ( .A(n6535), .B(n6327), .S(n7368), .Z(n6338) );
  NAND2_X1 U8023 ( .A1(n8192), .A2(n6381), .ZN(n6329) );
  OR2_X1 U8024 ( .A1(n4525), .A2(n8198), .ZN(n6328) );
  INV_X1 U8025 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n9742) );
  NAND2_X1 U8026 ( .A1(n6330), .A2(n9742), .ZN(n6331) );
  NAND2_X1 U8027 ( .A1(n9866), .A2(n6307), .ZN(n6337) );
  INV_X1 U8028 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n6334) );
  NAND2_X1 U8029 ( .A1(n6390), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n6333) );
  NAND2_X1 U8030 ( .A1(n6389), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n6332) );
  OAI211_X1 U8031 ( .C1(n6364), .C2(n6334), .A(n6333), .B(n6332), .ZN(n6335)
         );
  INV_X1 U8032 ( .A(n6335), .ZN(n6336) );
  NAND2_X1 U8033 ( .A1(n10111), .A2(n9655), .ZN(n6682) );
  INV_X1 U8034 ( .A(n9871), .ZN(n6343) );
  MUX2_X1 U8035 ( .A(n9869), .B(n6679), .S(n7368), .Z(n6342) );
  INV_X1 U8036 ( .A(n6682), .ZN(n6509) );
  MUX2_X1 U8037 ( .A(n6509), .B(n6340), .S(n7368), .Z(n6341) );
  NAND2_X1 U8038 ( .A1(n8640), .A2(n6381), .ZN(n6346) );
  OR2_X1 U8039 ( .A1(n4525), .A2(n6344), .ZN(n6345) );
  INV_X1 U8040 ( .A(n6349), .ZN(n6347) );
  INV_X1 U8041 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n6348) );
  NAND2_X1 U8042 ( .A1(n6349), .A2(n6348), .ZN(n6350) );
  NAND2_X1 U8043 ( .A1(n6360), .A2(n6350), .ZN(n8835) );
  INV_X1 U8044 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n8340) );
  NAND2_X1 U8045 ( .A1(n4380), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n6352) );
  NAND2_X1 U8046 ( .A1(n6389), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n6351) );
  OAI211_X1 U8047 ( .C1(n8340), .C2(n6388), .A(n6352), .B(n6351), .ZN(n6353)
         );
  INV_X1 U8048 ( .A(n6353), .ZN(n6354) );
  OR2_X1 U8049 ( .A1(n4525), .A2(n10250), .ZN(n6357) );
  INV_X1 U8050 ( .A(n6360), .ZN(n6359) );
  NAND2_X1 U8051 ( .A1(n6359), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n6702) );
  INV_X1 U8052 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n8362) );
  NAND2_X1 U8053 ( .A1(n6360), .A2(n8362), .ZN(n6361) );
  NAND2_X1 U8054 ( .A1(n6702), .A2(n6361), .ZN(n9847) );
  INV_X1 U8055 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n9846) );
  NAND2_X1 U8056 ( .A1(n6385), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n6363) );
  NAND2_X1 U8057 ( .A1(n6390), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n6362) );
  OAI211_X1 U8058 ( .C1(n6364), .C2(n9846), .A(n6363), .B(n6362), .ZN(n6365)
         );
  INV_X1 U8059 ( .A(n6365), .ZN(n6366) );
  NAND2_X1 U8060 ( .A1(n6685), .A2(n6412), .ZN(n6511) );
  OAI211_X1 U8061 ( .C1(n6368), .C2(n6511), .A(n6684), .B(n7368), .ZN(n6397)
         );
  NAND2_X1 U8062 ( .A1(n8692), .A2(n6381), .ZN(n6370) );
  OR2_X1 U8063 ( .A1(n4525), .A2(n10242), .ZN(n6369) );
  OR2_X1 U8064 ( .A1(n6702), .A2(n6371), .ZN(n6377) );
  INV_X1 U8065 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n6374) );
  NAND2_X1 U8066 ( .A1(n6389), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n6373) );
  NAND2_X1 U8067 ( .A1(n4380), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n6372) );
  OAI211_X1 U8068 ( .C1(n6374), .C2(n6388), .A(n6373), .B(n6372), .ZN(n6375)
         );
  INV_X1 U8069 ( .A(n6375), .ZN(n6376) );
  NAND2_X1 U8070 ( .A1(n10087), .A2(n9768), .ZN(n6555) );
  NAND2_X1 U8071 ( .A1(n10088), .A2(n7368), .ZN(n6396) );
  OR2_X1 U8072 ( .A1(n4525), .A2(n6378), .ZN(n6379) );
  NAND2_X1 U8073 ( .A1(n8856), .A2(n6381), .ZN(n6384) );
  INV_X1 U8074 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8859) );
  OR2_X1 U8075 ( .A1(n4525), .A2(n8859), .ZN(n6383) );
  INV_X1 U8076 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n8282) );
  NAND2_X1 U8077 ( .A1(n4380), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n6387) );
  NAND2_X1 U8078 ( .A1(n6385), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n6386) );
  OAI211_X1 U8079 ( .C1(n6388), .C2(n8282), .A(n6387), .B(n6386), .ZN(n9767)
         );
  INV_X1 U8080 ( .A(n9767), .ZN(n6438) );
  OR2_X1 U8081 ( .A1(n6437), .A2(n6438), .ZN(n6439) );
  NAND2_X1 U8082 ( .A1(n6389), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n6393) );
  NAND2_X1 U8083 ( .A1(n4380), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6392) );
  NAND2_X1 U8084 ( .A1(n6390), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6391) );
  NAND3_X1 U8085 ( .A1(n6393), .A2(n6392), .A3(n6391), .ZN(n9837) );
  NAND2_X1 U8086 ( .A1(n6439), .A2(n9837), .ZN(n6394) );
  NAND2_X1 U8087 ( .A1(n10079), .A2(n6394), .ZN(n6558) );
  NAND2_X1 U8088 ( .A1(n6558), .A2(n6512), .ZN(n6395) );
  AOI21_X1 U8089 ( .B1(n6397), .B2(n6396), .A(n6395), .ZN(n6407) );
  NAND2_X1 U8090 ( .A1(n9837), .A2(n9767), .ZN(n6399) );
  AND2_X1 U8091 ( .A1(n6437), .A2(n6399), .ZN(n6402) );
  INV_X1 U8092 ( .A(n6402), .ZN(n6554) );
  NAND4_X1 U8093 ( .A1(n6554), .A2(n4791), .A3(n6555), .A4(n6685), .ZN(n6405)
         );
  INV_X1 U8094 ( .A(n6452), .ZN(n6400) );
  INV_X1 U8095 ( .A(n6401), .ZN(n6404) );
  NAND2_X1 U8096 ( .A1(n10079), .A2(n4698), .ZN(n6440) );
  NAND3_X1 U8097 ( .A1(n6440), .A2(n6402), .A3(n7368), .ZN(n6403) );
  OAI211_X1 U8098 ( .C1(n5101), .C2(n6405), .A(n6404), .B(n6403), .ZN(n6406)
         );
  OR2_X1 U8099 ( .A1(n6409), .A2(n6408), .ZN(n6411) );
  NAND2_X1 U8100 ( .A1(n6688), .A2(n7419), .ZN(n6940) );
  INV_X1 U8101 ( .A(n6940), .ZN(n6908) );
  NAND2_X1 U8102 ( .A1(n6453), .A2(n6908), .ZN(n6450) );
  INV_X1 U8103 ( .A(n8838), .ZN(n6436) );
  INV_X1 U8104 ( .A(n9854), .ZN(n6435) );
  INV_X1 U8105 ( .A(n6619), .ZN(n6413) );
  INV_X1 U8106 ( .A(n6670), .ZN(n9914) );
  NAND2_X1 U8107 ( .A1(n6416), .A2(n6667), .ZN(n9958) );
  NAND2_X1 U8108 ( .A1(n6417), .A2(n6664), .ZN(n9990) );
  NAND2_X1 U8109 ( .A1(n6419), .A2(n8597), .ZN(n8096) );
  INV_X1 U8110 ( .A(n6420), .ZN(n7948) );
  NAND2_X1 U8111 ( .A1(n6649), .A2(n6421), .ZN(n6600) );
  INV_X1 U8112 ( .A(n6600), .ZN(n8035) );
  NAND2_X1 U8113 ( .A1(n6646), .A2(n6645), .ZN(n6594) );
  INV_X1 U8114 ( .A(n6594), .ZN(n7831) );
  AND2_X1 U8115 ( .A1(n4575), .A2(n7372), .ZN(n6487) );
  NOR2_X1 U8116 ( .A1(n7376), .A2(n6487), .ZN(n7188) );
  NAND4_X1 U8117 ( .A1(n7188), .A2(n7444), .A3(n7377), .A4(n7698), .ZN(n6424)
         );
  AND2_X1 U8118 ( .A1(n6587), .A2(n6586), .ZN(n7764) );
  NAND2_X1 U8119 ( .A1(n7764), .A2(n7464), .ZN(n6423) );
  NOR4_X1 U8120 ( .A1(n6424), .A2(n6423), .A3(n7812), .A4(n7514), .ZN(n6425)
         );
  AND2_X1 U8121 ( .A1(n6647), .A2(n8031), .ZN(n7895) );
  NAND4_X1 U8122 ( .A1(n8035), .A2(n7831), .A3(n6425), .A4(n7895), .ZN(n6426)
         );
  NOR3_X1 U8123 ( .A1(n8096), .A2(n7948), .A3(n6426), .ZN(n6427) );
  AND2_X1 U8124 ( .A1(n8608), .A2(n6427), .ZN(n6429) );
  XNOR2_X1 U8125 ( .A(n10174), .B(n6428), .ZN(n6657) );
  INV_X1 U8126 ( .A(n6657), .ZN(n10072) );
  NAND4_X1 U8127 ( .A1(n10029), .A2(n10036), .A3(n6429), .A4(n10072), .ZN(
        n6430) );
  NOR4_X1 U8128 ( .A1(n9958), .A2(n9990), .A3(n10013), .A4(n6430), .ZN(n6431)
         );
  AND4_X1 U8129 ( .A1(n9916), .A2(n9977), .A3(n4933), .A4(n6431), .ZN(n6432)
         );
  NAND3_X1 U8130 ( .A1(n9899), .A2(n4425), .A3(n6432), .ZN(n6433) );
  NOR3_X1 U8131 ( .A1(n9871), .A2(n9886), .A3(n6433), .ZN(n6434) );
  NAND2_X1 U8132 ( .A1(n6437), .A2(n6438), .ZN(n6514) );
  NAND3_X1 U8133 ( .A1(n6400), .A2(n5110), .A3(n6514), .ZN(n6441) );
  NAND2_X1 U8134 ( .A1(n6440), .A2(n6439), .ZN(n6516) );
  NAND2_X1 U8135 ( .A1(n6442), .A2(n7744), .ZN(n6561) );
  INV_X1 U8136 ( .A(n6448), .ZN(n6445) );
  NAND2_X1 U8137 ( .A1(n6445), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6446) );
  MUX2_X1 U8138 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6446), .S(
        P1_IR_REG_23__SCAN_IN), .Z(n6449) );
  NAND2_X1 U8139 ( .A1(n6448), .A2(n6447), .ZN(n6525) );
  NAND2_X1 U8140 ( .A1(n6449), .A2(n6525), .ZN(n6972) );
  NOR2_X1 U8141 ( .A1(n6972), .A2(P1_U3084), .ZN(n8019) );
  NAND2_X1 U8142 ( .A1(n10310), .A2(n8019), .ZN(n6518) );
  AOI211_X1 U8143 ( .C1(n6450), .C2(n6561), .A(n4377), .B(n6518), .ZN(n6571)
         );
  INV_X1 U8144 ( .A(n4377), .ZN(n7367) );
  NAND3_X1 U8145 ( .A1(n7419), .A2(n7367), .A3(n8019), .ZN(n6451) );
  INV_X1 U8146 ( .A(n6666), .ZN(n6454) );
  NOR2_X1 U8147 ( .A1(n6473), .A2(n6454), .ZN(n6486) );
  NOR2_X1 U8148 ( .A1(n6663), .A2(n6455), .ZN(n6477) );
  INV_X1 U8149 ( .A(n6456), .ZN(n6479) );
  INV_X1 U8150 ( .A(n6457), .ZN(n6478) );
  INV_X1 U8151 ( .A(n6458), .ZN(n6459) );
  NAND3_X1 U8152 ( .A1(n6479), .A2(n6478), .A3(n6459), .ZN(n6460) );
  NAND2_X1 U8153 ( .A1(n4442), .A2(n6460), .ZN(n6461) );
  NAND2_X1 U8154 ( .A1(n4807), .A2(n6461), .ZN(n6462) );
  NAND2_X1 U8155 ( .A1(n6462), .A2(n6656), .ZN(n6463) );
  NAND2_X1 U8156 ( .A1(n6463), .A2(n6658), .ZN(n6465) );
  NAND3_X1 U8157 ( .A1(n6465), .A2(n6464), .A3(n6659), .ZN(n6466) );
  NAND3_X1 U8158 ( .A1(n6486), .A2(n6477), .A3(n6466), .ZN(n6476) );
  INV_X1 U8159 ( .A(n6665), .ZN(n6470) );
  OAI211_X1 U8160 ( .C1(n6470), .C2(n6469), .A(n6468), .B(n6467), .ZN(n6471)
         );
  INV_X1 U8161 ( .A(n6471), .ZN(n6472) );
  OAI211_X1 U8162 ( .C1(n6473), .C2(n6472), .A(n6669), .B(n6675), .ZN(n6474)
         );
  INV_X1 U8163 ( .A(n6474), .ZN(n6475) );
  AND2_X1 U8164 ( .A1(n6476), .A2(n6475), .ZN(n6544) );
  INV_X1 U8165 ( .A(n6477), .ZN(n6484) );
  NAND4_X1 U8166 ( .A1(n6479), .A2(n6645), .A3(n6643), .A4(n6478), .ZN(n6480)
         );
  OR3_X1 U8167 ( .A1(n6482), .A2(n6481), .A3(n6480), .ZN(n6483) );
  NOR2_X1 U8168 ( .A1(n6484), .A2(n6483), .ZN(n6485) );
  NAND2_X1 U8169 ( .A1(n6486), .A2(n6485), .ZN(n6545) );
  OAI21_X1 U8170 ( .B1(n7463), .B2(n4401), .A(n7419), .ZN(n6490) );
  INV_X1 U8171 ( .A(n6487), .ZN(n6488) );
  OAI21_X1 U8172 ( .B1(n7483), .B2(n7469), .A(n6488), .ZN(n6489) );
  OAI211_X1 U8173 ( .C1(n6490), .C2(n6489), .A(n4517), .B(n7702), .ZN(n6495)
         );
  INV_X1 U8174 ( .A(n6586), .ZN(n6491) );
  AND2_X1 U8175 ( .A1(n9777), .A2(n10333), .ZN(n6493) );
  NAND2_X1 U8176 ( .A1(n6495), .A2(n5115), .ZN(n6500) );
  NAND3_X1 U8177 ( .A1(n6497), .A2(n6587), .A3(n6496), .ZN(n6498) );
  NAND2_X1 U8178 ( .A1(n4456), .A2(n6498), .ZN(n6538) );
  INV_X1 U8179 ( .A(n6543), .ZN(n6499) );
  AOI21_X1 U8180 ( .B1(n6500), .B2(n6538), .A(n6499), .ZN(n6501) );
  OR2_X1 U8181 ( .A1(n6545), .A2(n6501), .ZN(n6503) );
  AOI21_X1 U8182 ( .B1(n6544), .B2(n6503), .A(n6502), .ZN(n6506) );
  INV_X1 U8183 ( .A(n6504), .ZN(n6505) );
  OAI21_X1 U8184 ( .B1(n6506), .B2(n6505), .A(n6679), .ZN(n6507) );
  NAND2_X1 U8185 ( .A1(n6680), .A2(n6507), .ZN(n6508) );
  NOR2_X1 U8186 ( .A1(n8838), .A2(n6508), .ZN(n6513) );
  AND2_X1 U8187 ( .A1(n6683), .A2(n6509), .ZN(n6510) );
  OR2_X1 U8188 ( .A1(n6511), .A2(n6510), .ZN(n6534) );
  AND2_X1 U8189 ( .A1(n6512), .A2(n6684), .ZN(n6552) );
  OAI21_X1 U8190 ( .B1(n6513), .B2(n6534), .A(n6552), .ZN(n6515) );
  OR2_X1 U8191 ( .A1(n6516), .A2(n5109), .ZN(n6517) );
  INV_X1 U8192 ( .A(n6518), .ZN(n6519) );
  NAND3_X1 U8193 ( .A1(n6562), .A2(n6519), .A3(n4377), .ZN(n6568) );
  NAND2_X1 U8194 ( .A1(n6688), .A2(n9962), .ZN(n7373) );
  OR2_X1 U8195 ( .A1(n7373), .A2(n5002), .ZN(n7186) );
  INV_X1 U8196 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n6522) );
  NAND2_X1 U8197 ( .A1(n6523), .A2(n6522), .ZN(n6528) );
  OR2_X1 U8198 ( .A1(n6523), .A2(n6522), .ZN(n6524) );
  NAND2_X1 U8199 ( .A1(n6528), .A2(n6524), .ZN(n8519) );
  NAND2_X1 U8200 ( .A1(n6525), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6527) );
  NOR2_X1 U8201 ( .A1(n8519), .A2(n8133), .ZN(n6530) );
  NAND2_X1 U8202 ( .A1(n6972), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6949) );
  INV_X1 U8203 ( .A(n6949), .ZN(n6956) );
  NAND2_X1 U8204 ( .A1(n6974), .A2(n6956), .ZN(n6946) );
  OR3_X1 U8205 ( .A1(n4594), .A2(n6946), .A3(n7016), .ZN(n6533) );
  INV_X1 U8206 ( .A(P1_B_REG_SCAN_IN), .ZN(n6692) );
  AOI21_X1 U8207 ( .B1(n7892), .B2(n8019), .A(n6692), .ZN(n6532) );
  OAI21_X1 U8208 ( .B1(n7186), .B2(n6533), .A(n6532), .ZN(n6567) );
  AND2_X1 U8209 ( .A1(n9962), .A2(n8019), .ZN(n6563) );
  INV_X1 U8210 ( .A(n6534), .ZN(n6551) );
  INV_X1 U8211 ( .A(n6535), .ZN(n6548) );
  NAND2_X1 U8212 ( .A1(n6536), .A2(n5115), .ZN(n6542) );
  OAI21_X1 U8213 ( .B1(n6539), .B2(n7702), .A(n6538), .ZN(n6540) );
  INV_X1 U8214 ( .A(n6540), .ZN(n6541) );
  NAND2_X1 U8215 ( .A1(n7512), .A2(n6543), .ZN(n6644) );
  INV_X1 U8216 ( .A(n6644), .ZN(n6546) );
  OAI211_X1 U8217 ( .C1(n6546), .C2(n6545), .A(n6544), .B(n6677), .ZN(n6547)
         );
  NAND2_X1 U8218 ( .A1(n6548), .A2(n6547), .ZN(n6549) );
  NAND4_X1 U8219 ( .A1(n6683), .A2(n6680), .A3(n9869), .A4(n6549), .ZN(n6550)
         );
  NAND2_X1 U8220 ( .A1(n6551), .A2(n6550), .ZN(n6553) );
  NAND2_X1 U8221 ( .A1(n6553), .A2(n6552), .ZN(n6556) );
  NAND3_X1 U8222 ( .A1(n6556), .A2(n6555), .A3(n6554), .ZN(n6557) );
  NAND2_X1 U8223 ( .A1(n6558), .A2(n6557), .ZN(n6559) );
  NAND3_X1 U8224 ( .A1(n6559), .A2(n7419), .A3(n6400), .ZN(n6560) );
  NAND4_X1 U8225 ( .A1(n6561), .A2(n7367), .A3(n6563), .A4(n6560), .ZN(n6566)
         );
  INV_X1 U8226 ( .A(n6562), .ZN(n6564) );
  NAND3_X1 U8227 ( .A1(n6564), .A2(n6563), .A3(n4377), .ZN(n6565) );
  NAND4_X1 U8228 ( .A1(n6568), .A2(n6567), .A3(n6566), .A4(n6565), .ZN(n6569)
         );
  NAND2_X1 U8229 ( .A1(n6729), .A2(n7422), .ZN(n7369) );
  NAND2_X1 U8230 ( .A1(n7369), .A2(n7463), .ZN(n6581) );
  NAND2_X1 U8231 ( .A1(n6581), .A2(n4401), .ZN(n6574) );
  INV_X1 U8232 ( .A(n6572), .ZN(n6573) );
  NAND2_X1 U8233 ( .A1(n6574), .A2(n6573), .ZN(n6575) );
  NAND2_X1 U8234 ( .A1(n6575), .A2(n7469), .ZN(n6585) );
  INV_X1 U8235 ( .A(n7369), .ZN(n7370) );
  NAND3_X1 U8236 ( .A1(n7370), .A2(n9780), .A3(n6580), .ZN(n6583) );
  AND2_X1 U8237 ( .A1(n6582), .A2(n6583), .ZN(n6584) );
  AND2_X1 U8238 ( .A1(n9777), .A2(n7711), .ZN(n6589) );
  NAND2_X1 U8239 ( .A1(n8209), .A2(n7903), .ZN(n7809) );
  NAND2_X1 U8240 ( .A1(n7767), .A2(n6590), .ZN(n6592) );
  INV_X1 U8241 ( .A(n7458), .ZN(n7629) );
  OR2_X1 U8242 ( .A1(n9779), .A2(n7629), .ZN(n7697) );
  NAND2_X1 U8243 ( .A1(n6587), .A2(n6586), .ZN(n6588) );
  NAND2_X1 U8244 ( .A1(n7484), .A2(n10333), .ZN(n7762) );
  OAI211_X1 U8245 ( .C1(n6589), .C2(n7697), .A(n6588), .B(n7762), .ZN(n7766)
         );
  NAND2_X1 U8246 ( .A1(n8207), .A2(n7748), .ZN(n7828) );
  NAND2_X1 U8247 ( .A1(n6594), .A2(n7828), .ZN(n6597) );
  INV_X1 U8248 ( .A(n7828), .ZN(n6593) );
  NOR2_X1 U8249 ( .A1(n7514), .A2(n6593), .ZN(n6595) );
  INV_X1 U8250 ( .A(n8530), .ZN(n9774) );
  AOI22_X1 U8251 ( .A1(n6595), .A2(n6594), .B1(n10206), .B2(n9774), .ZN(n6596)
         );
  AND2_X1 U8252 ( .A1(n10201), .A2(n9773), .ZN(n6599) );
  NAND2_X1 U8253 ( .A1(n8034), .A2(n6600), .ZN(n6602) );
  INV_X1 U8254 ( .A(n7950), .ZN(n9772) );
  OR2_X1 U8255 ( .A1(n10196), .A2(n9772), .ZN(n6601) );
  NAND2_X1 U8256 ( .A1(n6602), .A2(n6601), .ZN(n7945) );
  NOR2_X1 U8257 ( .A1(n7958), .A2(n9771), .ZN(n6604) );
  NAND2_X1 U8258 ( .A1(n7958), .A2(n9771), .ZN(n6603) );
  AND2_X1 U8259 ( .A1(n10178), .A2(n10058), .ZN(n10068) );
  AND2_X1 U8260 ( .A1(n10174), .A2(n10037), .ZN(n6610) );
  NOR2_X1 U8261 ( .A1(n10068), .A2(n6610), .ZN(n6605) );
  NAND2_X1 U8262 ( .A1(n10184), .A2(n9770), .ZN(n8606) );
  AND2_X1 U8263 ( .A1(n6605), .A2(n8606), .ZN(n6606) );
  NAND2_X1 U8264 ( .A1(n9707), .A2(n6607), .ZN(n10070) );
  OR2_X1 U8265 ( .A1(n10174), .A2(n10037), .ZN(n6608) );
  AND2_X1 U8266 ( .A1(n10070), .A2(n6608), .ZN(n6609) );
  NOR2_X1 U8267 ( .A1(n10048), .A2(n9612), .ZN(n6611) );
  INV_X1 U8268 ( .A(n9612), .ZN(n10056) );
  INV_X1 U8269 ( .A(n9759), .ZN(n10038) );
  NAND2_X1 U8270 ( .A1(n10148), .A2(n9988), .ZN(n6615) );
  INV_X1 U8271 ( .A(n10148), .ZN(n9975) );
  INV_X1 U8272 ( .A(n10144), .ZN(n6853) );
  NAND2_X1 U8273 ( .A1(n10144), .A2(n9979), .ZN(n6617) );
  INV_X1 U8274 ( .A(n10140), .ZN(n9942) );
  NOR2_X1 U8275 ( .A1(n10131), .A2(n9951), .ZN(n6618) );
  NAND2_X1 U8276 ( .A1(n9881), .A2(n9886), .ZN(n6622) );
  NAND2_X1 U8277 ( .A1(n9885), .A2(n9744), .ZN(n6621) );
  NAND2_X1 U8278 ( .A1(n6622), .A2(n6621), .ZN(n9862) );
  NOR2_X1 U8279 ( .A1(n10107), .A2(n9873), .ZN(n6624) );
  NAND2_X1 U8280 ( .A1(n10102), .A2(n9769), .ZN(n10095) );
  NAND2_X1 U8281 ( .A1(n4378), .A2(n10095), .ZN(n6625) );
  XNOR2_X1 U8282 ( .A(n6625), .B(n10088), .ZN(n6712) );
  AND2_X1 U8283 ( .A1(n9962), .A2(n4377), .ZN(n6906) );
  OR2_X1 U8284 ( .A1(n6940), .A2(n6906), .ZN(n6626) );
  NAND2_X1 U8285 ( .A1(n6626), .A2(n6974), .ZN(n6928) );
  INV_X1 U8286 ( .A(n6926), .ZN(n7101) );
  NAND2_X1 U8287 ( .A1(n8519), .A2(P1_B_REG_SCAN_IN), .ZN(n6628) );
  INV_X1 U8288 ( .A(n8133), .ZN(n6627) );
  MUX2_X1 U8289 ( .A(n6628), .B(P1_B_REG_SCAN_IN), .S(n6627), .Z(n6629) );
  NAND2_X1 U8290 ( .A1(n6629), .A2(n6951), .ZN(n6947) );
  INV_X1 U8291 ( .A(n8519), .ZN(n6950) );
  OAI22_X1 U8292 ( .A1(n6947), .A2(P1_D_REG_1__SCAN_IN), .B1(n6951), .B2(n6950), .ZN(n7191) );
  INV_X1 U8293 ( .A(n7191), .ZN(n6639) );
  INV_X1 U8294 ( .A(n6947), .ZN(n6640) );
  NOR4_X1 U8295 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_2__SCAN_IN), .A4(P1_D_REG_4__SCAN_IN), .ZN(n6637) );
  NOR4_X1 U8296 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_20__SCAN_IN), .A3(
        P1_D_REG_30__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n6636) );
  INV_X1 U8297 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n10323) );
  INV_X1 U8298 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n10321) );
  INV_X1 U8299 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n10325) );
  INV_X1 U8300 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n10326) );
  NAND4_X1 U8301 ( .A1(n10323), .A2(n10321), .A3(n10325), .A4(n10326), .ZN(
        n8225) );
  NOR4_X1 U8302 ( .A1(P1_D_REG_8__SCAN_IN), .A2(P1_D_REG_9__SCAN_IN), .A3(
        P1_D_REG_11__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n6633) );
  NOR4_X1 U8303 ( .A1(P1_D_REG_5__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_7__SCAN_IN), .A4(P1_D_REG_10__SCAN_IN), .ZN(n6632) );
  NOR4_X1 U8304 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_25__SCAN_IN), .A4(P1_D_REG_26__SCAN_IN), .ZN(n6631) );
  NOR4_X1 U8305 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_16__SCAN_IN), .A3(
        P1_D_REG_23__SCAN_IN), .A4(P1_D_REG_19__SCAN_IN), .ZN(n6630) );
  NAND4_X1 U8306 ( .A1(n6633), .A2(n6632), .A3(n6631), .A4(n6630), .ZN(n6634)
         );
  NOR4_X1 U8307 ( .A1(P1_D_REG_31__SCAN_IN), .A2(P1_D_REG_28__SCAN_IN), .A3(
        n8225), .A4(n6634), .ZN(n6635) );
  NAND3_X1 U8308 ( .A1(n6637), .A2(n6636), .A3(n6635), .ZN(n6638) );
  NAND2_X1 U8309 ( .A1(n6640), .A2(n6638), .ZN(n7190) );
  NAND2_X1 U8310 ( .A1(n6639), .A2(n7190), .ZN(n6909) );
  INV_X1 U8311 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n6957) );
  INV_X1 U8312 ( .A(n6951), .ZN(n8196) );
  AND2_X1 U8313 ( .A1(n8196), .A2(n8133), .ZN(n6955) );
  AOI21_X1 U8314 ( .B1(n6640), .B2(n6957), .A(n6955), .ZN(n7210) );
  NOR2_X1 U8315 ( .A1(n6909), .A2(n7210), .ZN(n6641) );
  NAND2_X1 U8316 ( .A1(n7101), .A2(n6641), .ZN(n6701) );
  NAND2_X1 U8317 ( .A1(n7892), .A2(n7744), .ZN(n7185) );
  AND2_X1 U8318 ( .A1(n7186), .A2(n6806), .ZN(n6642) );
  NAND2_X1 U8319 ( .A1(n10315), .A2(n6642), .ZN(n10074) );
  NAND2_X1 U8320 ( .A1(n8032), .A2(n6648), .ZN(n6650) );
  NAND2_X1 U8321 ( .A1(n6650), .A2(n6649), .ZN(n7947) );
  OR2_X1 U8322 ( .A1(n6653), .A2(n8597), .ZN(n8599) );
  AND2_X1 U8323 ( .A1(n8599), .A2(n6654), .ZN(n6655) );
  NAND2_X1 U8324 ( .A1(n8600), .A2(n6655), .ZN(n10054) );
  NAND2_X1 U8325 ( .A1(n10034), .A2(n6658), .ZN(n6660) );
  OAI211_X1 U8326 ( .C1(n6671), .C2(n9912), .A(n9916), .B(n6670), .ZN(n6672)
         );
  INV_X1 U8327 ( .A(n6672), .ZN(n6673) );
  NAND2_X1 U8328 ( .A1(n6674), .A2(n6673), .ZN(n9915) );
  NAND2_X1 U8329 ( .A1(n9898), .A2(n6676), .ZN(n6678) );
  NAND2_X1 U8330 ( .A1(n9887), .A2(n6679), .ZN(n9870) );
  AND2_X1 U8331 ( .A1(n9869), .A2(n6680), .ZN(n6681) );
  INV_X1 U8332 ( .A(n6684), .ZN(n6686) );
  OAI21_X1 U8333 ( .B1(n9855), .B2(n6686), .A(n6685), .ZN(n6687) );
  XNOR2_X1 U8334 ( .A(n6687), .B(n10097), .ZN(n10100) );
  NAND2_X1 U8335 ( .A1(n6688), .A2(n10310), .ZN(n6690) );
  OR2_X1 U8336 ( .A1(n7744), .A2(n4377), .ZN(n6689) );
  INV_X2 U8337 ( .A(n10315), .ZN(n10317) );
  AND2_X1 U8338 ( .A1(n10099), .A2(n10315), .ZN(n6691) );
  NAND2_X1 U8339 ( .A1(n10100), .A2(n6691), .ZN(n6695) );
  INV_X1 U8340 ( .A(n7016), .ZN(n7323) );
  OR2_X1 U8341 ( .A1(n6940), .A2(n7323), .ZN(n9952) );
  NOR2_X1 U8342 ( .A1(n4594), .A2(n6692), .ZN(n6693) );
  NOR2_X1 U8343 ( .A1(n9952), .A2(n6693), .ZN(n9838) );
  AOI22_X1 U8344 ( .A1(n9769), .A2(n10057), .B1(n9838), .B2(n9767), .ZN(n10092) );
  OR2_X1 U8345 ( .A1(n10317), .A2(n10092), .ZN(n6694) );
  NAND2_X1 U8346 ( .A1(n6695), .A2(n6694), .ZN(n6710) );
  NAND2_X1 U8347 ( .A1(n7454), .A2(n7458), .ZN(n7708) );
  INV_X1 U8348 ( .A(n10196), .ZN(n8043) );
  NAND2_X1 U8349 ( .A1(n7956), .A2(n10190), .ZN(n7955) );
  OR2_X2 U8350 ( .A1(n7955), .A2(n10184), .ZN(n8604) );
  NOR2_X4 U8351 ( .A1(n8604), .A2(n10178), .ZN(n10061) );
  INV_X1 U8352 ( .A(n10174), .ZN(n10060) );
  INV_X1 U8353 ( .A(n10164), .ZN(n6699) );
  AND2_X1 U8354 ( .A1(n6699), .A2(n10048), .ZN(n10006) );
  AND2_X1 U8355 ( .A1(n10006), .A2(n10011), .ZN(n6700) );
  AND2_X2 U8356 ( .A1(n9931), .A2(n10131), .ZN(n9933) );
  OR2_X2 U8357 ( .A1(n9849), .A2(n10102), .ZN(n9850) );
  NOR2_X1 U8358 ( .A1(n6701), .A2(n10310), .ZN(n10077) );
  INV_X1 U8359 ( .A(n10087), .ZN(n6705) );
  NOR2_X1 U8360 ( .A1(n7185), .A2(n4377), .ZN(n10306) );
  NAND2_X1 U8361 ( .A1(n10315), .A2(n10306), .ZN(n10047) );
  INV_X1 U8362 ( .A(n6702), .ZN(n6703) );
  INV_X1 U8363 ( .A(n9992), .ZN(n10307) );
  AOI22_X1 U8364 ( .A1(n6703), .A2(n10307), .B1(P1_REG2_REG_29__SCAN_IN), .B2(
        n10317), .ZN(n6704) );
  OAI21_X1 U8365 ( .B1(n6705), .B2(n10047), .A(n6704), .ZN(n6706) );
  INV_X1 U8366 ( .A(n6706), .ZN(n6707) );
  NAND2_X1 U8367 ( .A1(n7892), .A2(n6906), .ZN(n7420) );
  NOR2_X1 U8368 ( .A1(n6714), .A2(n6734), .ZN(n6715) );
  AOI21_X1 U8369 ( .B1(n10154), .B2(n6800), .A(n6715), .ZN(n9727) );
  NAND2_X1 U8370 ( .A1(n10154), .A2(n6918), .ZN(n6717) );
  NAND2_X1 U8371 ( .A1(n10004), .A2(n6800), .ZN(n6716) );
  NAND2_X1 U8372 ( .A1(n6717), .A2(n6716), .ZN(n6718) );
  XNOR2_X1 U8373 ( .A(n6718), .B(n4422), .ZN(n9626) );
  NAND2_X1 U8374 ( .A1(n9777), .A2(n6800), .ZN(n6720) );
  NAND2_X1 U8375 ( .A1(n6918), .A2(n7711), .ZN(n6719) );
  NAND2_X1 U8376 ( .A1(n6720), .A2(n6719), .ZN(n6721) );
  XNOR2_X1 U8377 ( .A(n6721), .B(n6806), .ZN(n6748) );
  OAI22_X1 U8378 ( .A1(n7484), .A2(n6734), .B1(n10333), .B2(n6871), .ZN(n6747)
         );
  INV_X1 U8379 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n6982) );
  NOR2_X1 U8380 ( .A1(n6974), .A2(n6982), .ZN(n6722) );
  AOI21_X1 U8381 ( .B1(n6918), .B2(n7422), .A(n6722), .ZN(n6724) );
  NAND2_X1 U8382 ( .A1(n4575), .A2(n6800), .ZN(n6723) );
  NAND2_X1 U8383 ( .A1(n6724), .A2(n6723), .ZN(n7104) );
  AOI21_X1 U8384 ( .B1(n6913), .B2(n4575), .A(n6728), .ZN(n7105) );
  NAND2_X1 U8385 ( .A1(n7105), .A2(n7104), .ZN(n7103) );
  OAI21_X1 U8386 ( .B1(n4422), .B2(n7104), .A(n7103), .ZN(n6731) );
  INV_X1 U8387 ( .A(n6731), .ZN(n6733) );
  INV_X1 U8388 ( .A(n6800), .ZN(n6777) );
  OAI22_X1 U8389 ( .A1(n7463), .A2(n6777), .B1(n4400), .B2(n6874), .ZN(n6730)
         );
  XNOR2_X1 U8390 ( .A(n6730), .B(n6806), .ZN(n6732) );
  AOI22_X1 U8391 ( .A1(n9780), .A2(n6913), .B1(n6800), .B2(n4401), .ZN(n7306)
         );
  OAI21_X1 U8392 ( .B1(n6733), .B2(n6732), .A(n7304), .ZN(n7401) );
  OAI22_X1 U8393 ( .A1(n7483), .A2(n6734), .B1(n7506), .B2(n6871), .ZN(n6737)
         );
  OAI22_X1 U8394 ( .A1(n7483), .A2(n6777), .B1(n7506), .B2(n6874), .ZN(n6735)
         );
  XNOR2_X1 U8395 ( .A(n6735), .B(n6806), .ZN(n6736) );
  XOR2_X1 U8396 ( .A(n6737), .B(n6736), .Z(n7400) );
  INV_X1 U8397 ( .A(n6736), .ZN(n6739) );
  INV_X1 U8398 ( .A(n6737), .ZN(n6738) );
  AOI22_X1 U8399 ( .A1(n6913), .A2(n9779), .B1(n6800), .B2(n7629), .ZN(n6743)
         );
  NAND2_X1 U8400 ( .A1(n9779), .A2(n6800), .ZN(n6741) );
  NAND2_X1 U8401 ( .A1(n7629), .A2(n6918), .ZN(n6740) );
  NAND2_X1 U8402 ( .A1(n6741), .A2(n6740), .ZN(n6742) );
  XNOR2_X1 U8403 ( .A(n6742), .B(n6806), .ZN(n6745) );
  XOR2_X1 U8404 ( .A(n6743), .B(n6745), .Z(n7481) );
  INV_X1 U8405 ( .A(n6743), .ZN(n6744) );
  XOR2_X1 U8406 ( .A(n6748), .B(n6747), .Z(n7602) );
  AOI22_X1 U8407 ( .A1(n6913), .A2(n9776), .B1(n7819), .B2(n6800), .ZN(n8202)
         );
  INV_X1 U8408 ( .A(n8202), .ZN(n6757) );
  NAND2_X1 U8409 ( .A1(n7819), .A2(n6918), .ZN(n6750) );
  NAND2_X1 U8410 ( .A1(n9776), .A2(n6800), .ZN(n6749) );
  NAND2_X1 U8411 ( .A1(n6750), .A2(n6749), .ZN(n6751) );
  XNOR2_X1 U8412 ( .A(n6751), .B(n6806), .ZN(n8203) );
  NAND2_X1 U8413 ( .A1(n8209), .A2(n6800), .ZN(n6753) );
  NAND2_X1 U8414 ( .A1(n6918), .A2(n7903), .ZN(n6752) );
  NAND2_X1 U8415 ( .A1(n6753), .A2(n6752), .ZN(n6754) );
  XNOR2_X1 U8416 ( .A(n6754), .B(n4422), .ZN(n8201) );
  INV_X1 U8417 ( .A(n8201), .ZN(n6758) );
  NAND2_X1 U8418 ( .A1(n6913), .A2(n8209), .ZN(n6756) );
  NAND2_X1 U8419 ( .A1(n6800), .A2(n7903), .ZN(n6755) );
  AND2_X1 U8420 ( .A1(n6756), .A2(n6755), .ZN(n6759) );
  AOI22_X1 U8421 ( .A1(n6757), .A2(n8203), .B1(n6758), .B2(n7844), .ZN(n6764)
         );
  NOR3_X1 U8422 ( .A1(n6758), .A2(n6757), .A3(n7844), .ZN(n6762) );
  AOI21_X1 U8423 ( .B1(n8201), .B2(n6759), .A(n8202), .ZN(n6760) );
  NOR2_X1 U8424 ( .A1(n6760), .A2(n8203), .ZN(n6761) );
  OR2_X1 U8425 ( .A1(n8207), .A2(n6734), .ZN(n6766) );
  OR2_X1 U8426 ( .A1(n7748), .A2(n6871), .ZN(n6765) );
  NAND2_X1 U8427 ( .A1(n6766), .A2(n6765), .ZN(n6769) );
  OAI22_X1 U8428 ( .A1(n8207), .A2(n6871), .B1(n7748), .B2(n6874), .ZN(n6767)
         );
  XNOR2_X1 U8429 ( .A(n6767), .B(n6806), .ZN(n6768) );
  XNOR2_X1 U8430 ( .A(n6769), .B(n6768), .ZN(n7747) );
  AOI22_X1 U8431 ( .A1(n9774), .A2(n6913), .B1(n6800), .B2(n10206), .ZN(n6771)
         );
  NAND2_X1 U8432 ( .A1(n6772), .A2(n6771), .ZN(n8105) );
  AOI22_X1 U8433 ( .A1(n9774), .A2(n6800), .B1(n10206), .B2(n6918), .ZN(n6770)
         );
  XOR2_X1 U8434 ( .A(n6806), .B(n6770), .Z(n8108) );
  AOI22_X1 U8435 ( .A1(n10201), .A2(n6800), .B1(n6913), .B2(n9773), .ZN(n6787)
         );
  AOI22_X1 U8436 ( .A1(n10201), .A2(n6918), .B1(n6800), .B2(n9773), .ZN(n6773)
         );
  XNOR2_X1 U8437 ( .A(n6773), .B(n6806), .ZN(n6788) );
  XOR2_X1 U8438 ( .A(n6787), .B(n6788), .Z(n8525) );
  NAND2_X1 U8439 ( .A1(n10196), .A2(n6918), .ZN(n6775) );
  OR2_X1 U8440 ( .A1(n7950), .A2(n6871), .ZN(n6774) );
  NAND2_X1 U8441 ( .A1(n6775), .A2(n6774), .ZN(n6776) );
  XNOR2_X1 U8442 ( .A(n6776), .B(n6806), .ZN(n6780) );
  INV_X1 U8443 ( .A(n6780), .ZN(n6779) );
  OAI22_X1 U8444 ( .A1(n8043), .A2(n6777), .B1(n7950), .B2(n6734), .ZN(n6781)
         );
  INV_X1 U8445 ( .A(n6781), .ZN(n6778) );
  NAND2_X1 U8446 ( .A1(n6779), .A2(n6778), .ZN(n6789) );
  INV_X1 U8447 ( .A(n6789), .ZN(n6782) );
  XOR2_X1 U8448 ( .A(n6781), .B(n6780), .Z(n8575) );
  AND2_X1 U8449 ( .A1(n8525), .A2(n6786), .ZN(n8536) );
  OAI22_X1 U8450 ( .A1(n10190), .A2(n6871), .B1(n8589), .B2(n6734), .ZN(n6795)
         );
  NAND2_X1 U8451 ( .A1(n7958), .A2(n6918), .ZN(n6784) );
  NAND2_X1 U8452 ( .A1(n9771), .A2(n6800), .ZN(n6783) );
  NAND2_X1 U8453 ( .A1(n6784), .A2(n6783), .ZN(n6785) );
  XNOR2_X1 U8454 ( .A(n6785), .B(n6806), .ZN(n6794) );
  XOR2_X1 U8455 ( .A(n6795), .B(n6794), .Z(n8540) );
  AND2_X1 U8456 ( .A1(n8536), .A2(n8540), .ZN(n6793) );
  INV_X1 U8457 ( .A(n8540), .ZN(n6792) );
  INV_X1 U8458 ( .A(n6786), .ZN(n6791) );
  NAND2_X1 U8459 ( .A1(n6788), .A2(n6787), .ZN(n8572) );
  AND2_X1 U8460 ( .A1(n8572), .A2(n6789), .ZN(n6790) );
  AOI21_X1 U8461 ( .B1(n8524), .B2(n6793), .A(n5093), .ZN(n6799) );
  INV_X1 U8462 ( .A(n6794), .ZN(n6797) );
  INV_X1 U8463 ( .A(n6795), .ZN(n6796) );
  NAND2_X1 U8464 ( .A1(n6797), .A2(n6796), .ZN(n6798) );
  NAND2_X1 U8465 ( .A1(n6799), .A2(n6798), .ZN(n8586) );
  OAI22_X1 U8466 ( .A1(n8590), .A2(n6874), .B1(n9706), .B2(n6871), .ZN(n6801)
         );
  XNOR2_X1 U8467 ( .A(n6801), .B(n6806), .ZN(n8584) );
  OAI22_X1 U8468 ( .A1(n8590), .A2(n6871), .B1(n9706), .B2(n6734), .ZN(n8583)
         );
  NOR2_X1 U8469 ( .A1(n8584), .A2(n8583), .ZN(n6803) );
  NAND2_X1 U8470 ( .A1(n8584), .A2(n8583), .ZN(n6802) );
  OAI21_X2 U8471 ( .B1(n8586), .B2(n6803), .A(n6802), .ZN(n9702) );
  NAND2_X1 U8472 ( .A1(n10174), .A2(n6918), .ZN(n6805) );
  NAND2_X1 U8473 ( .A1(n10037), .A2(n6800), .ZN(n6804) );
  NAND2_X1 U8474 ( .A1(n6805), .A2(n6804), .ZN(n6807) );
  XNOR2_X1 U8475 ( .A(n6807), .B(n6806), .ZN(n9603) );
  INV_X1 U8476 ( .A(n9603), .ZN(n9605) );
  NAND2_X1 U8477 ( .A1(n10174), .A2(n6800), .ZN(n6809) );
  NAND2_X1 U8478 ( .A1(n6913), .A2(n10037), .ZN(n6808) );
  NAND2_X1 U8479 ( .A1(n6809), .A2(n6808), .ZN(n9607) );
  INV_X1 U8480 ( .A(n9607), .ZN(n9659) );
  NAND2_X1 U8481 ( .A1(n10178), .A2(n6918), .ZN(n6811) );
  NAND2_X1 U8482 ( .A1(n10058), .A2(n6800), .ZN(n6810) );
  NAND2_X1 U8483 ( .A1(n6811), .A2(n6810), .ZN(n6812) );
  XNOR2_X1 U8484 ( .A(n6812), .B(n6806), .ZN(n6822) );
  INV_X1 U8485 ( .A(n6822), .ZN(n6816) );
  NAND2_X1 U8486 ( .A1(n10178), .A2(n6800), .ZN(n6814) );
  NAND2_X1 U8487 ( .A1(n6913), .A2(n10058), .ZN(n6813) );
  NAND2_X1 U8488 ( .A1(n6814), .A2(n6813), .ZN(n6821) );
  INV_X1 U8489 ( .A(n6821), .ZN(n6815) );
  AOI21_X1 U8490 ( .B1(n9605), .B2(n9659), .A(n9699), .ZN(n6826) );
  NAND2_X1 U8491 ( .A1(n10164), .A2(n6918), .ZN(n6818) );
  OR2_X1 U8492 ( .A1(n9759), .A2(n6871), .ZN(n6817) );
  NAND2_X1 U8493 ( .A1(n6818), .A2(n6817), .ZN(n6819) );
  XNOR2_X1 U8494 ( .A(n6819), .B(n4422), .ZN(n6829) );
  AOI22_X1 U8495 ( .A1(n10164), .A2(n6800), .B1(n6913), .B2(n10038), .ZN(n9664) );
  OAI22_X1 U8496 ( .A1(n10048), .A2(n6874), .B1(n9612), .B2(n6871), .ZN(n6820)
         );
  XNOR2_X1 U8497 ( .A(n6820), .B(n6806), .ZN(n9661) );
  OAI22_X1 U8498 ( .A1(n10048), .A2(n6871), .B1(n9612), .B2(n6734), .ZN(n6827)
         );
  AOI22_X1 U8499 ( .A1(n9661), .A2(n6827), .B1(n9700), .B2(n9607), .ZN(n6824)
         );
  OAI21_X1 U8500 ( .B1(n9700), .B2(n9607), .A(n9603), .ZN(n6823) );
  OAI211_X1 U8501 ( .C1(n6829), .C2(n9664), .A(n6824), .B(n6823), .ZN(n6825)
         );
  INV_X1 U8502 ( .A(n6827), .ZN(n9753) );
  INV_X1 U8503 ( .A(n9661), .ZN(n6828) );
  AOI21_X1 U8504 ( .B1(n9753), .B2(n6828), .A(n9664), .ZN(n6831) );
  INV_X1 U8505 ( .A(n6829), .ZN(n9665) );
  NAND2_X1 U8506 ( .A1(n9664), .A2(n9753), .ZN(n6830) );
  OAI22_X1 U8507 ( .A1(n6831), .A2(n9665), .B1(n9661), .B2(n6830), .ZN(n9674)
         );
  NAND2_X1 U8508 ( .A1(n10158), .A2(n6918), .ZN(n6833) );
  NAND2_X1 U8509 ( .A1(n10019), .A2(n6800), .ZN(n6832) );
  NAND2_X1 U8510 ( .A1(n6833), .A2(n6832), .ZN(n6834) );
  XNOR2_X1 U8511 ( .A(n6834), .B(n6806), .ZN(n6836) );
  INV_X1 U8512 ( .A(n6836), .ZN(n6835) );
  OAI22_X1 U8513 ( .A1(n10011), .A2(n6871), .B1(n9669), .B2(n6734), .ZN(n6837)
         );
  AND2_X1 U8514 ( .A1(n6835), .A2(n4505), .ZN(n6838) );
  NAND2_X1 U8515 ( .A1(n10148), .A2(n6918), .ZN(n6841) );
  NAND2_X1 U8516 ( .A1(n9988), .A2(n6800), .ZN(n6840) );
  NAND2_X1 U8517 ( .A1(n6841), .A2(n6840), .ZN(n6842) );
  XNOR2_X1 U8518 ( .A(n6842), .B(n6806), .ZN(n9629) );
  NAND2_X1 U8519 ( .A1(n10148), .A2(n6800), .ZN(n6844) );
  NAND2_X1 U8520 ( .A1(n9988), .A2(n6913), .ZN(n6843) );
  NAND2_X1 U8521 ( .A1(n6844), .A2(n6843), .ZN(n9628) );
  NAND2_X1 U8522 ( .A1(n9626), .A2(n9727), .ZN(n6845) );
  INV_X1 U8523 ( .A(n6845), .ZN(n6848) );
  INV_X1 U8524 ( .A(n9628), .ZN(n6847) );
  AOI21_X1 U8525 ( .B1(n9628), .B2(n6845), .A(n9629), .ZN(n6846) );
  AOI21_X1 U8526 ( .B1(n6848), .B2(n6847), .A(n6846), .ZN(n6849) );
  NAND2_X1 U8527 ( .A1(n10144), .A2(n6918), .ZN(n6851) );
  NAND2_X1 U8528 ( .A1(n9979), .A2(n6800), .ZN(n6850) );
  NAND2_X1 U8529 ( .A1(n6851), .A2(n6850), .ZN(n6852) );
  XNOR2_X1 U8530 ( .A(n6852), .B(n6806), .ZN(n6863) );
  OAI22_X1 U8531 ( .A1(n6853), .A2(n6871), .B1(n9953), .B2(n6734), .ZN(n6864)
         );
  XOR2_X1 U8532 ( .A(n6863), .B(n6864), .Z(n9693) );
  NAND2_X1 U8533 ( .A1(n10140), .A2(n6918), .ZN(n6855) );
  NAND2_X1 U8534 ( .A1(n9959), .A2(n6800), .ZN(n6854) );
  NAND2_X1 U8535 ( .A1(n6855), .A2(n6854), .ZN(n6856) );
  INV_X1 U8536 ( .A(n6861), .ZN(n6858) );
  OAI22_X1 U8537 ( .A1(n9942), .A2(n6871), .B1(n6857), .B2(n6734), .ZN(n6859)
         );
  NAND2_X1 U8538 ( .A1(n6858), .A2(n6860), .ZN(n6867) );
  INV_X1 U8539 ( .A(n6867), .ZN(n6862) );
  INV_X1 U8540 ( .A(n6863), .ZN(n6866) );
  INV_X1 U8541 ( .A(n6864), .ZN(n6865) );
  NAND2_X1 U8542 ( .A1(n6866), .A2(n6865), .ZN(n9638) );
  AOI22_X1 U8543 ( .A1(n9934), .A2(n6800), .B1(n6913), .B2(n9918), .ZN(n6873)
         );
  OAI22_X1 U8544 ( .A1(n10131), .A2(n6874), .B1(n9951), .B2(n6871), .ZN(n6872)
         );
  XNOR2_X1 U8545 ( .A(n6872), .B(n6806), .ZN(n9716) );
  OAI22_X1 U8546 ( .A1(n9910), .A2(n6874), .B1(n9720), .B2(n6871), .ZN(n6875)
         );
  XNOR2_X1 U8547 ( .A(n6875), .B(n6806), .ZN(n6877) );
  OAI22_X1 U8548 ( .A1(n9910), .A2(n6871), .B1(n9720), .B2(n6734), .ZN(n9619)
         );
  AOI22_X1 U8549 ( .A1(n10121), .A2(n6918), .B1(n6800), .B2(n9919), .ZN(n6878)
         );
  XNOR2_X1 U8550 ( .A(n6878), .B(n6806), .ZN(n6880) );
  AOI22_X1 U8551 ( .A1(n10121), .A2(n6800), .B1(n6913), .B2(n9919), .ZN(n6879)
         );
  XNOR2_X1 U8552 ( .A(n6880), .B(n6879), .ZN(n9685) );
  NAND2_X1 U8553 ( .A1(n6880), .A2(n6879), .ZN(n6881) );
  NAND2_X1 U8554 ( .A1(n9682), .A2(n6881), .ZN(n9648) );
  OAI22_X1 U8555 ( .A1(n9885), .A2(n6871), .B1(n9744), .B2(n6734), .ZN(n6886)
         );
  NAND2_X1 U8556 ( .A1(n10116), .A2(n6918), .ZN(n6883) );
  NAND2_X1 U8557 ( .A1(n9900), .A2(n6800), .ZN(n6882) );
  NAND2_X1 U8558 ( .A1(n6883), .A2(n6882), .ZN(n6884) );
  XNOR2_X1 U8559 ( .A(n6884), .B(n6806), .ZN(n6885) );
  XOR2_X1 U8560 ( .A(n6886), .B(n6885), .Z(n9649) );
  NAND2_X1 U8561 ( .A1(n9648), .A2(n9649), .ZN(n6890) );
  INV_X1 U8562 ( .A(n6885), .ZN(n6888) );
  INV_X1 U8563 ( .A(n6886), .ZN(n6887) );
  NAND2_X1 U8564 ( .A1(n6888), .A2(n6887), .ZN(n6889) );
  NAND2_X1 U8565 ( .A1(n6890), .A2(n6889), .ZN(n9739) );
  NAND2_X1 U8566 ( .A1(n10111), .A2(n6918), .ZN(n6892) );
  NAND2_X1 U8567 ( .A1(n9888), .A2(n6800), .ZN(n6891) );
  NAND2_X1 U8568 ( .A1(n6892), .A2(n6891), .ZN(n6893) );
  XNOR2_X1 U8569 ( .A(n6893), .B(n6806), .ZN(n6899) );
  AND2_X1 U8570 ( .A1(n9888), .A2(n6913), .ZN(n6894) );
  AOI21_X1 U8571 ( .B1(n10111), .B2(n6800), .A(n6894), .ZN(n6897) );
  XOR2_X1 U8572 ( .A(n6899), .B(n6897), .Z(n9738) );
  INV_X1 U8573 ( .A(n9738), .ZN(n6895) );
  INV_X1 U8574 ( .A(n6897), .ZN(n6898) );
  NAND2_X1 U8575 ( .A1(n10107), .A2(n6918), .ZN(n6901) );
  NAND2_X1 U8576 ( .A1(n9873), .A2(n6800), .ZN(n6900) );
  NAND2_X1 U8577 ( .A1(n6901), .A2(n6900), .ZN(n6902) );
  XNOR2_X1 U8578 ( .A(n6902), .B(n4422), .ZN(n6912) );
  INV_X1 U8579 ( .A(n6912), .ZN(n6905) );
  NOR2_X1 U8580 ( .A1(n9745), .A2(n6734), .ZN(n6903) );
  AOI21_X1 U8581 ( .B1(n10107), .B2(n6800), .A(n6903), .ZN(n6911) );
  INV_X1 U8582 ( .A(n6911), .ZN(n6904) );
  INV_X1 U8583 ( .A(n7185), .ZN(n7189) );
  INV_X1 U8584 ( .A(n6906), .ZN(n6907) );
  NOR2_X1 U8585 ( .A1(n10207), .A2(n6908), .ZN(n6910) );
  INV_X1 U8586 ( .A(n7210), .ZN(n7194) );
  NOR2_X1 U8587 ( .A1(n6927), .A2(n6946), .ZN(n6923) );
  NAND2_X1 U8588 ( .A1(n6910), .A2(n6923), .ZN(n9737) );
  AND2_X1 U8589 ( .A1(n6912), .A2(n6911), .ZN(n9595) );
  INV_X1 U8590 ( .A(n9595), .ZN(n6932) );
  NAND2_X1 U8591 ( .A1(n10102), .A2(n6800), .ZN(n6915) );
  NAND2_X1 U8592 ( .A1(n9769), .A2(n6913), .ZN(n6914) );
  NAND2_X1 U8593 ( .A1(n6915), .A2(n6914), .ZN(n6916) );
  XNOR2_X1 U8594 ( .A(n6916), .B(n4422), .ZN(n6920) );
  NOR2_X1 U8595 ( .A1(n9596), .A2(n6777), .ZN(n6917) );
  AOI21_X1 U8596 ( .B1(n10102), .B2(n6918), .A(n6917), .ZN(n6919) );
  XNOR2_X1 U8597 ( .A(n6920), .B(n6919), .ZN(n6936) );
  NAND4_X1 U8598 ( .A1(n6935), .A2(n8526), .A3(n6932), .A4(n6936), .ZN(n6939)
         );
  NAND2_X1 U8599 ( .A1(n6923), .A2(n10306), .ZN(n6921) );
  NAND2_X1 U8600 ( .A1(n6921), .A2(n9992), .ZN(n9734) );
  INV_X1 U8601 ( .A(n7186), .ZN(n6922) );
  NAND2_X1 U8602 ( .A1(n6923), .A2(n6922), .ZN(n6924) );
  OR2_X1 U8603 ( .A1(n6924), .A2(n7016), .ZN(n9743) );
  NOR2_X1 U8604 ( .A1(n10334), .A2(n9962), .ZN(n6925) );
  NOR2_X1 U8605 ( .A1(n6926), .A2(n6925), .ZN(n7193) );
  NAND2_X1 U8606 ( .A1(n7193), .A2(n6927), .ZN(n7102) );
  AOI21_X1 U8607 ( .B1(n6928), .B2(P1_STATE_REG_SCAN_IN), .A(n8019), .ZN(n6929) );
  NAND2_X1 U8608 ( .A1(n7102), .A2(n6929), .ZN(n9763) );
  INV_X1 U8609 ( .A(n9763), .ZN(n9732) );
  OAI22_X1 U8610 ( .A1(n9847), .A2(n9732), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8362), .ZN(n6930) );
  AOI21_X1 U8611 ( .B1(n9873), .B2(n9755), .A(n6930), .ZN(n6931) );
  OAI21_X1 U8612 ( .B1(n9768), .B2(n9758), .A(n6931), .ZN(n6934) );
  NOR3_X1 U8613 ( .A1(n6936), .A2(n6932), .A3(n9765), .ZN(n6933) );
  AOI211_X1 U8614 ( .C1(n9734), .C2(n10102), .A(n6934), .B(n6933), .ZN(n6938)
         );
  NAND3_X1 U8615 ( .A1(n6939), .A2(n6938), .A3(n6937), .ZN(P1_U3218) );
  OR2_X1 U8616 ( .A1(n7548), .A2(P2_U3152), .ZN(n7148) );
  OR2_X2 U8617 ( .A1(n7148), .A2(n7545), .ZN(n9037) );
  NAND2_X1 U8618 ( .A1(n6940), .A2(n6974), .ZN(n6941) );
  NAND2_X1 U8619 ( .A1(n6941), .A2(n6972), .ZN(n7014) );
  NAND2_X1 U8620 ( .A1(n7014), .A2(n6977), .ZN(n6942) );
  NAND2_X1 U8621 ( .A1(n6942), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  AND2_X1 U8622 ( .A1(n4399), .A2(P1_U3084), .ZN(n10246) );
  INV_X2 U8623 ( .A(n10246), .ZN(n10244) );
  OAI222_X1 U8624 ( .A1(n10251), .A2(n6943), .B1(n10244), .B2(n6970), .C1(
        P1_U3084), .C2(n7009), .ZN(P1_U3349) );
  INV_X1 U8625 ( .A(n7008), .ZN(n7069) );
  OAI222_X1 U8626 ( .A1(n10251), .A2(n6944), .B1(n10244), .B2(n6967), .C1(
        P1_U3084), .C2(n7069), .ZN(P1_U3350) );
  INV_X1 U8627 ( .A(n6099), .ZN(n6969) );
  INV_X1 U8628 ( .A(n7046), .ZN(n7004) );
  OAI222_X1 U8629 ( .A1(n10251), .A2(n6945), .B1(n10244), .B2(n6969), .C1(
        P1_U3084), .C2(n7004), .ZN(P1_U3347) );
  INV_X1 U8630 ( .A(n6946), .ZN(n6948) );
  NAND2_X1 U8631 ( .A1(n6948), .A2(n6947), .ZN(n10328) );
  INV_X1 U8632 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n6953) );
  NOR3_X1 U8633 ( .A1(n6951), .A2(n6950), .A3(n6949), .ZN(n6952) );
  AOI21_X1 U8634 ( .B1(n10328), .B2(n6953), .A(n6952), .ZN(P1_U3441) );
  OAI222_X1 U8635 ( .A1(P1_U3084), .A2(n7006), .B1(n10251), .B2(n6954), .C1(
        n10244), .C2(n6985), .ZN(P1_U3352) );
  AOI22_X1 U8636 ( .A1(n10328), .A2(n6957), .B1(n6956), .B2(n6955), .ZN(
        P1_U3440) );
  OAI222_X1 U8637 ( .A1(n4376), .A2(P1_U3084), .B1(n10244), .B2(n6988), .C1(
        n6958), .C2(n10251), .ZN(P1_U3351) );
  OAI222_X1 U8638 ( .A1(n10251), .A2(n6959), .B1(n10244), .B2(n6991), .C1(
        P1_U3084), .C2(n7037), .ZN(P1_U3348) );
  INV_X1 U8639 ( .A(n6960), .ZN(n6966) );
  INV_X1 U8640 ( .A(n10251), .ZN(n10239) );
  AOI22_X1 U8641 ( .A1(n7177), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n10239), .ZN(n6961) );
  OAI21_X1 U8642 ( .B1(n6966), .B2(n10244), .A(n6961), .ZN(P1_U3345) );
  INV_X1 U8643 ( .A(n6962), .ZN(n6965) );
  AOI22_X1 U8644 ( .A1(n7080), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n10239), .ZN(n6963) );
  OAI21_X1 U8645 ( .B1(n6965), .B2(n10244), .A(n6963), .ZN(P1_U3346) );
  NAND2_X1 U8646 ( .A1(n4398), .A2(P2_U3152), .ZN(n8866) );
  INV_X1 U8647 ( .A(n8866), .ZN(n7440) );
  INV_X1 U8648 ( .A(n7440), .ZN(n9586) );
  NAND2_X1 U8649 ( .A1(n6964), .A2(P2_U3152), .ZN(n8864) );
  INV_X1 U8650 ( .A(n7387), .ZN(n7269) );
  OAI222_X1 U8651 ( .A1(n9586), .A2(n4554), .B1(n8864), .B2(n6965), .C1(
        P2_U3152), .C2(n7269), .ZN(P2_U3351) );
  INV_X1 U8652 ( .A(n8864), .ZN(n8014) );
  INV_X1 U8653 ( .A(n8014), .ZN(n9591) );
  INV_X1 U8654 ( .A(n7494), .ZN(n7399) );
  OAI222_X1 U8655 ( .A1(n9586), .A2(n8236), .B1(n9591), .B2(n6966), .C1(
        P2_U3152), .C2(n7399), .ZN(P2_U3350) );
  OAI222_X1 U8656 ( .A1(n9586), .A2(n6968), .B1(n9591), .B2(n6967), .C1(
        P2_U3152), .C2(n7253), .ZN(P2_U3355) );
  INV_X1 U8657 ( .A(n7260), .ZN(n7240) );
  OAI222_X1 U8658 ( .A1(n9586), .A2(n4539), .B1(n9591), .B2(n6969), .C1(
        P2_U3152), .C2(n7240), .ZN(P2_U3352) );
  OAI222_X1 U8659 ( .A1(n9586), .A2(n6971), .B1(n9591), .B2(n6970), .C1(
        P2_U3152), .C2(n7281), .ZN(P2_U3354) );
  INV_X1 U8660 ( .A(n6972), .ZN(n6973) );
  NOR2_X1 U8661 ( .A1(n6974), .A2(n6973), .ZN(n6975) );
  OR2_X1 U8662 ( .A1(P1_U3083), .A2(n6975), .ZN(n8719) );
  INV_X1 U8663 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n10431) );
  INV_X1 U8664 ( .A(n4594), .ZN(n6980) );
  INV_X1 U8665 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n7425) );
  AOI21_X1 U8666 ( .B1(n6980), .B2(n7425), .A(n7016), .ZN(n6976) );
  XNOR2_X1 U8667 ( .A(n6976), .B(P1_IR_REG_0__SCAN_IN), .ZN(n7326) );
  OAI211_X1 U8668 ( .C1(n6980), .C2(P1_REG1_REG_0__SCAN_IN), .A(n6977), .B(
        P1_STATE_REG_SCAN_IN), .ZN(n6978) );
  NOR2_X1 U8669 ( .A1(n7326), .A2(n6978), .ZN(n6979) );
  AOI22_X1 U8670 ( .A1(n7014), .A2(n6979), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        P1_U3084), .ZN(n6984) );
  OR2_X1 U8671 ( .A1(n7016), .A2(P1_U3084), .ZN(n10248) );
  NOR2_X1 U8672 ( .A1(n10248), .A2(n6980), .ZN(n6981) );
  NAND3_X1 U8673 ( .A1(n10302), .A2(P1_IR_REG_0__SCAN_IN), .A3(n6982), .ZN(
        n6983) );
  OAI211_X1 U8674 ( .C1(n8719), .C2(n10431), .A(n6984), .B(n6983), .ZN(
        P1_U3241) );
  OAI222_X1 U8675 ( .A1(P2_U3152), .A2(n7204), .B1(n9586), .B2(n6986), .C1(
        n9591), .C2(n6985), .ZN(P2_U3357) );
  OAI222_X1 U8676 ( .A1(n7223), .A2(P2_U3152), .B1(n9591), .B2(n6988), .C1(
        n6987), .C2(n9586), .ZN(P2_U3356) );
  INV_X1 U8677 ( .A(n6989), .ZN(n6992) );
  AOI22_X1 U8678 ( .A1(n7409), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n10239), .ZN(n6990) );
  OAI21_X1 U8679 ( .B1(n6992), .B2(n10244), .A(n6990), .ZN(P1_U3344) );
  INV_X1 U8680 ( .A(n7287), .ZN(n7295) );
  OAI222_X1 U8681 ( .A1(n9586), .A2(n4757), .B1(n9591), .B2(n6991), .C1(
        P2_U3152), .C2(n7295), .ZN(P2_U3353) );
  INV_X1 U8682 ( .A(n7731), .ZN(n7503) );
  OAI222_X1 U8683 ( .A1(n8866), .A2(n6993), .B1(n9591), .B2(n6992), .C1(n7503), 
        .C2(P2_U3152), .ZN(P2_U3349) );
  NAND2_X1 U8684 ( .A1(n9837), .A2(P1_U4006), .ZN(n6994) );
  OAI21_X1 U8685 ( .B1(P1_U4006), .B2(n9587), .A(n6994), .ZN(P1_U3586) );
  INV_X1 U8686 ( .A(n6995), .ZN(n6997) );
  INV_X1 U8687 ( .A(n8142), .ZN(n7741) );
  OAI222_X1 U8688 ( .A1(n8866), .A2(n6996), .B1(n8864), .B2(n6997), .C1(n7741), 
        .C2(P2_U3152), .ZN(P2_U3348) );
  INV_X1 U8689 ( .A(n7429), .ZN(n7426) );
  OAI222_X1 U8690 ( .A1(n10251), .A2(n6998), .B1(n10244), .B2(n6997), .C1(
        n7426), .C2(P1_U3084), .ZN(P1_U3343) );
  INV_X1 U8691 ( .A(n10302), .ZN(n9823) );
  XNOR2_X1 U8692 ( .A(n7080), .B(P1_REG1_REG_7__SCAN_IN), .ZN(n7081) );
  INV_X1 U8693 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n7005) );
  INV_X1 U8694 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n7003) );
  INV_X1 U8695 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n7002) );
  INV_X1 U8696 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n7001) );
  XNOR2_X1 U8697 ( .A(n7006), .B(P1_REG1_REG_1__SCAN_IN), .ZN(n7055) );
  AND2_X1 U8698 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n7054) );
  NAND2_X1 U8699 ( .A1(n7055), .A2(n7054), .ZN(n7053) );
  INV_X1 U8700 ( .A(n7006), .ZN(n7052) );
  NAND2_X1 U8701 ( .A1(n7052), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6999) );
  NAND2_X1 U8702 ( .A1(n7053), .A2(n6999), .ZN(n7334) );
  INV_X1 U8703 ( .A(n4376), .ZN(n7332) );
  NAND2_X1 U8704 ( .A1(n7332), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n7000) );
  NAND2_X1 U8705 ( .A1(n7333), .A2(n7000), .ZN(n7065) );
  XNOR2_X1 U8706 ( .A(n7008), .B(n7001), .ZN(n7066) );
  INV_X1 U8707 ( .A(n7009), .ZN(n9789) );
  XNOR2_X1 U8708 ( .A(n9789), .B(P1_REG1_REG_4__SCAN_IN), .ZN(n9785) );
  XNOR2_X1 U8709 ( .A(n7037), .B(P1_REG1_REG_5__SCAN_IN), .ZN(n7031) );
  NAND2_X1 U8710 ( .A1(n7030), .A2(n7031), .ZN(n7029) );
  OAI21_X1 U8711 ( .B1(n7037), .B2(n7003), .A(n7029), .ZN(n7041) );
  MUX2_X1 U8712 ( .A(n7005), .B(P1_REG1_REG_6__SCAN_IN), .S(n7046), .Z(n7042)
         );
  XOR2_X1 U8713 ( .A(n7081), .B(n7082), .Z(n7021) );
  XOR2_X1 U8714 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n7080), .Z(n7013) );
  NAND2_X1 U8715 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n7060) );
  XOR2_X1 U8716 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n4376), .Z(n7330) );
  XNOR2_X1 U8717 ( .A(n7008), .B(P1_REG2_REG_3__SCAN_IN), .ZN(n7071) );
  XNOR2_X1 U8718 ( .A(n7009), .B(P1_REG2_REG_4__SCAN_IN), .ZN(n9791) );
  XNOR2_X1 U8719 ( .A(n7037), .B(P1_REG2_REG_5__SCAN_IN), .ZN(n7026) );
  INV_X1 U8720 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n7010) );
  INV_X1 U8721 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n7011) );
  MUX2_X1 U8722 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n7011), .S(n7046), .Z(n7039)
         );
  OAI21_X1 U8723 ( .B1(n7013), .B2(n7012), .A(n7077), .ZN(n7015) );
  NOR2_X1 U8724 ( .A1(n4594), .A2(P1_U3084), .ZN(n8641) );
  NAND2_X1 U8725 ( .A1(n7014), .A2(n8641), .ZN(n8715) );
  INV_X1 U8726 ( .A(n8715), .ZN(n7017) );
  AND2_X1 U8727 ( .A1(n7017), .A2(n7323), .ZN(n10292) );
  INV_X1 U8728 ( .A(n8719), .ZN(n10301) );
  AOI22_X1 U8729 ( .A1(n7015), .A2(n10292), .B1(n10301), .B2(
        P1_ADDR_REG_7__SCAN_IN), .ZN(n7020) );
  AND2_X1 U8730 ( .A1(n7017), .A2(n7016), .ZN(n10294) );
  NAND2_X1 U8731 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3084), .ZN(n7749) );
  INV_X1 U8732 ( .A(n7749), .ZN(n7018) );
  AOI21_X1 U8733 ( .B1(n10294), .B2(n7080), .A(n7018), .ZN(n7019) );
  OAI211_X1 U8734 ( .C1(n9823), .C2(n7021), .A(n7020), .B(n7019), .ZN(P1_U3248) );
  INV_X1 U8735 ( .A(n7022), .ZN(n7024) );
  INV_X1 U8736 ( .A(n7719), .ZN(n7023) );
  OAI222_X1 U8737 ( .A1(n10251), .A2(n8414), .B1(n10244), .B2(n7024), .C1(
        n7023), .C2(P1_U3084), .ZN(P1_U3342) );
  INV_X1 U8738 ( .A(n9048), .ZN(n8146) );
  OAI222_X1 U8739 ( .A1(n9586), .A2(n7025), .B1(n9591), .B2(n7024), .C1(n8146), 
        .C2(P2_U3152), .ZN(P2_U3347) );
  INV_X1 U8740 ( .A(n10294), .ZN(n9818) );
  XNOR2_X1 U8741 ( .A(n7027), .B(n7026), .ZN(n7028) );
  AOI22_X1 U8742 ( .A1(n7028), .A2(n10292), .B1(n10301), .B2(
        P1_ADDR_REG_5__SCAN_IN), .ZN(n7036) );
  OAI211_X1 U8743 ( .C1(n7031), .C2(n7030), .A(n10302), .B(n7029), .ZN(n7032)
         );
  INV_X1 U8744 ( .A(n7032), .ZN(n7034) );
  NAND2_X1 U8745 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3084), .ZN(n7846) );
  INV_X1 U8746 ( .A(n7846), .ZN(n7033) );
  NOR2_X1 U8747 ( .A1(n7034), .A2(n7033), .ZN(n7035) );
  OAI211_X1 U8748 ( .C1(n7037), .C2(n9818), .A(n7036), .B(n7035), .ZN(P1_U3246) );
  OAI211_X1 U8749 ( .C1(n7039), .C2(n7038), .A(n4501), .B(n10292), .ZN(n7048)
         );
  NAND2_X1 U8750 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_U3084), .ZN(n8206) );
  INV_X1 U8751 ( .A(n8206), .ZN(n7045) );
  AOI21_X1 U8752 ( .B1(n7042), .B2(n7041), .A(n7040), .ZN(n7043) );
  NOR2_X1 U8753 ( .A1(n7043), .A2(n9823), .ZN(n7044) );
  AOI211_X1 U8754 ( .C1(n10294), .C2(n7046), .A(n7045), .B(n7044), .ZN(n7047)
         );
  OAI211_X1 U8755 ( .C1(n8719), .C2(n4530), .A(n7048), .B(n7047), .ZN(P1_U3247) );
  NAND2_X1 U8756 ( .A1(n8209), .A2(P1_U4006), .ZN(n7049) );
  OAI21_X1 U8757 ( .B1(P1_U4006), .B2(n4757), .A(n7049), .ZN(P1_U3560) );
  NAND2_X1 U8758 ( .A1(n9037), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n7050) );
  OAI21_X1 U8759 ( .B1(n9037), .B2(n9162), .A(n7050), .ZN(P2_U3582) );
  NAND2_X1 U8760 ( .A1(n9037), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n7051) );
  OAI21_X1 U8761 ( .B1(n9037), .B2(n9387), .A(n7051), .ZN(P2_U3569) );
  INV_X1 U8762 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n7312) );
  NAND2_X1 U8763 ( .A1(n10294), .A2(n7052), .ZN(n7057) );
  OAI211_X1 U8764 ( .C1(n7055), .C2(n7054), .A(n10302), .B(n7053), .ZN(n7056)
         );
  OAI211_X1 U8765 ( .C1(P1_STATE_REG_SCAN_IN), .C2(n7312), .A(n7057), .B(n7056), .ZN(n7062) );
  INV_X1 U8766 ( .A(n10292), .ZN(n9830) );
  AOI211_X1 U8767 ( .C1(n7060), .C2(n7059), .A(n7058), .B(n9830), .ZN(n7061)
         );
  AOI211_X1 U8768 ( .C1(n10301), .C2(P1_ADDR_REG_1__SCAN_IN), .A(n7062), .B(
        n7061), .ZN(n7063) );
  INV_X1 U8769 ( .A(n7063), .ZN(P1_U3242) );
  INV_X1 U8770 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n8466) );
  NOR2_X1 U8771 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8466), .ZN(n7486) );
  INV_X1 U8772 ( .A(n7486), .ZN(n7068) );
  OAI211_X1 U8773 ( .C1(n7066), .C2(n7065), .A(n10302), .B(n7064), .ZN(n7067)
         );
  OAI211_X1 U8774 ( .C1(n9818), .C2(n7069), .A(n7068), .B(n7067), .ZN(n7074)
         );
  AOI211_X1 U8775 ( .C1(n7072), .C2(n7071), .A(n7070), .B(n9830), .ZN(n7073)
         );
  AOI211_X1 U8776 ( .C1(n10301), .C2(P1_ADDR_REG_3__SCAN_IN), .A(n7074), .B(
        n7073), .ZN(n7075) );
  INV_X1 U8777 ( .A(n7075), .ZN(P1_U3244) );
  INV_X1 U8778 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n7836) );
  MUX2_X1 U8779 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n7836), .S(n7177), .Z(n7079)
         );
  OAI21_X1 U8780 ( .B1(n7079), .B2(n7078), .A(n7176), .ZN(n7088) );
  XNOR2_X1 U8781 ( .A(n7177), .B(P1_REG1_REG_8__SCAN_IN), .ZN(n7084) );
  NOR2_X1 U8782 ( .A1(n7083), .A2(n7084), .ZN(n7172) );
  AOI211_X1 U8783 ( .C1(n7084), .C2(n7083), .A(n9823), .B(n7172), .ZN(n7087)
         );
  AND2_X1 U8784 ( .A1(P1_U3084), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n8110) );
  AOI21_X1 U8785 ( .B1(n10294), .B2(n7177), .A(n8110), .ZN(n7085) );
  OAI21_X1 U8786 ( .B1(n8719), .B2(n4563), .A(n7085), .ZN(n7086) );
  AOI211_X1 U8787 ( .C1(n7088), .C2(n10292), .A(n7087), .B(n7086), .ZN(n7089)
         );
  INV_X1 U8788 ( .A(n7089), .ZN(P1_U3249) );
  NAND2_X1 U8789 ( .A1(n10373), .A2(n7589), .ZN(n7090) );
  NAND2_X1 U8790 ( .A1(n7090), .A2(n7154), .ZN(n7093) );
  OR2_X1 U8791 ( .A1(n10373), .A2(n7091), .ZN(n7092) );
  NAND2_X1 U8792 ( .A1(n7093), .A2(n7092), .ZN(n9131) );
  NOR2_X1 U8793 ( .A1(n10358), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U8794 ( .A(n7094), .ZN(n7096) );
  INV_X1 U8795 ( .A(n8649), .ZN(n8644) );
  OAI222_X1 U8796 ( .A1(n9586), .A2(n7095), .B1(n8864), .B2(n7096), .C1(
        P2_U3152), .C2(n8644), .ZN(P2_U3346) );
  INV_X1 U8797 ( .A(n7858), .ZN(n7854) );
  OAI222_X1 U8798 ( .A1(P1_U3084), .A2(n7854), .B1(n10244), .B2(n7096), .C1(
        n10251), .C2(n5362), .ZN(P1_U3341) );
  NAND2_X1 U8799 ( .A1(P2_U3966), .A2(n7318), .ZN(n7097) );
  OAI21_X1 U8800 ( .B1(P2_U3966), .B2(n6044), .A(n7097), .ZN(P2_U3552) );
  NAND2_X1 U8801 ( .A1(P2_U3966), .A2(n8973), .ZN(n7098) );
  OAI21_X1 U8802 ( .B1(P2_U3966), .B2(n5362), .A(n7098), .ZN(P2_U3564) );
  NAND2_X1 U8803 ( .A1(P2_U3966), .A2(n7099), .ZN(n7100) );
  OAI21_X1 U8804 ( .B1(P2_U3966), .B2(n6378), .A(n7100), .ZN(P2_U3583) );
  NAND2_X1 U8805 ( .A1(n7102), .A2(n7101), .ZN(n7404) );
  INV_X1 U8806 ( .A(n7404), .ZN(n7313) );
  INV_X1 U8807 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n7108) );
  OAI21_X1 U8808 ( .B1(n7105), .B2(n7104), .A(n7103), .ZN(n7324) );
  OAI22_X1 U8809 ( .A1(n9760), .A2(n7372), .B1(n9758), .B2(n7463), .ZN(n7106)
         );
  AOI21_X1 U8810 ( .B1(n7324), .B2(n8526), .A(n7106), .ZN(n7107) );
  OAI21_X1 U8811 ( .B1(n7313), .B2(n7108), .A(n7107), .ZN(P1_U3230) );
  INV_X1 U8812 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n7110) );
  INV_X1 U8813 ( .A(n7109), .ZN(n7111) );
  INV_X1 U8814 ( .A(n8632), .ZN(n7857) );
  OAI222_X1 U8815 ( .A1(n10251), .A2(n7110), .B1(n10244), .B2(n7111), .C1(
        n7857), .C2(P1_U3084), .ZN(P1_U3340) );
  INV_X1 U8816 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n7112) );
  INV_X1 U8817 ( .A(n8681), .ZN(n8677) );
  OAI222_X1 U8818 ( .A1(n9586), .A2(n7112), .B1(n8864), .B2(n7111), .C1(n8677), 
        .C2(P2_U3152), .ZN(P2_U3345) );
  INV_X1 U8819 ( .A(n8709), .ZN(n8695) );
  INV_X1 U8820 ( .A(n7113), .ZN(n7114) );
  OAI222_X1 U8821 ( .A1(P1_U3084), .A2(n8695), .B1(n10244), .B2(n7114), .C1(
        n8428), .C2(n10251), .ZN(P1_U3339) );
  INV_X1 U8822 ( .A(n9059), .ZN(n9054) );
  OAI222_X1 U8823 ( .A1(n9586), .A2(n7115), .B1(n8864), .B2(n7114), .C1(n9054), 
        .C2(P2_U3152), .ZN(P2_U3344) );
  INV_X1 U8824 ( .A(n7116), .ZN(n7118) );
  INV_X1 U8825 ( .A(n9078), .ZN(n9068) );
  OAI222_X1 U8826 ( .A1(n9586), .A2(n7117), .B1(n8864), .B2(n7118), .C1(
        P2_U3152), .C2(n9068), .ZN(P2_U3343) );
  OAI222_X1 U8827 ( .A1(n10251), .A2(n7119), .B1(n10244), .B2(n7118), .C1(
        P1_U3084), .C2(n9802), .ZN(P1_U3338) );
  INV_X1 U8828 ( .A(n7135), .ZN(n8137) );
  INV_X1 U8829 ( .A(P2_B_REG_SCAN_IN), .ZN(n7120) );
  INV_X1 U8830 ( .A(n7122), .ZN(n8521) );
  OAI221_X1 U8831 ( .B1(n7135), .B2(P2_B_REG_SCAN_IN), .C1(n8137), .C2(n7120), 
        .A(n8521), .ZN(n7121) );
  INV_X1 U8832 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n10384) );
  NOR2_X1 U8833 ( .A1(n8193), .A2(n7122), .ZN(n10386) );
  AOI21_X1 U8834 ( .B1(n10371), .B2(n10384), .A(n10386), .ZN(n7542) );
  INV_X1 U8835 ( .A(n7542), .ZN(n7134) );
  NOR4_X1 U8836 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_16__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_18__SCAN_IN), .ZN(n7126) );
  NOR4_X1 U8837 ( .A1(P2_D_REG_13__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_11__SCAN_IN), .A4(P2_D_REG_14__SCAN_IN), .ZN(n7125) );
  NOR4_X1 U8838 ( .A1(P2_D_REG_25__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n7124) );
  NOR4_X1 U8839 ( .A1(P2_D_REG_19__SCAN_IN), .A2(P2_D_REG_20__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_23__SCAN_IN), .ZN(n7123) );
  NAND4_X1 U8840 ( .A1(n7126), .A2(n7125), .A3(n7124), .A4(n7123), .ZN(n7132)
         );
  NOR2_X1 U8841 ( .A1(P2_D_REG_12__SCAN_IN), .A2(P2_D_REG_8__SCAN_IN), .ZN(
        n7130) );
  NOR4_X1 U8842 ( .A1(P2_D_REG_28__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_3__SCAN_IN), .A4(P2_D_REG_29__SCAN_IN), .ZN(n7129) );
  NOR4_X1 U8843 ( .A1(P2_D_REG_5__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_7__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n7128) );
  NOR4_X1 U8844 ( .A1(P2_D_REG_24__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_2__SCAN_IN), .A4(P2_D_REG_4__SCAN_IN), .ZN(n7127) );
  NAND4_X1 U8845 ( .A1(n7130), .A2(n7129), .A3(n7128), .A4(n7127), .ZN(n7131)
         );
  OAI21_X1 U8846 ( .B1(n7132), .B2(n7131), .A(n10371), .ZN(n7541) );
  NAND2_X1 U8847 ( .A1(n7589), .A2(n4896), .ZN(n7546) );
  NAND2_X1 U8848 ( .A1(n10373), .A2(n7546), .ZN(n7869) );
  NOR2_X1 U8849 ( .A1(n9518), .A2(n7537), .ZN(n7556) );
  NOR2_X1 U8850 ( .A1(n7869), .A2(n7556), .ZN(n7133) );
  INV_X1 U8851 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n10381) );
  NOR2_X1 U8852 ( .A1(n7135), .A2(n8193), .ZN(n10382) );
  INV_X1 U8853 ( .A(n7870), .ZN(n7136) );
  AND2_X2 U8854 ( .A1(n7362), .A2(n7136), .ZN(n10418) );
  INV_X1 U8855 ( .A(n7137), .ZN(n7139) );
  INV_X1 U8856 ( .A(n7140), .ZN(n8854) );
  NAND2_X1 U8857 ( .A1(n7589), .A2(n8854), .ZN(n9386) );
  AOI22_X1 U8858 ( .A1(n8023), .A2(n4402), .B1(n9412), .B2(n7141), .ZN(n8024)
         );
  XNOR2_X1 U8859 ( .A(n7142), .B(n7884), .ZN(n7143) );
  NAND2_X1 U8860 ( .A1(n7143), .A2(n7537), .ZN(n8560) );
  NOR2_X1 U8861 ( .A1(n7543), .A2(n7537), .ZN(n7144) );
  NAND2_X1 U8862 ( .A1(n7144), .A2(n8862), .ZN(n9556) );
  NAND2_X1 U8863 ( .A1(n10399), .A2(n8023), .ZN(n7145) );
  OAI211_X1 U8864 ( .C1(n7554), .C2(n7595), .A(n8024), .B(n7145), .ZN(n9559)
         );
  NAND2_X1 U8865 ( .A1(n10418), .A2(n9559), .ZN(n7146) );
  OAI21_X1 U8866 ( .B1(n10418), .B2(n5165), .A(n7146), .ZN(P2_U3451) );
  INV_X1 U8867 ( .A(n7223), .ZN(n7214) );
  INV_X1 U8868 ( .A(n7589), .ZN(n7147) );
  NAND2_X1 U8869 ( .A1(n10373), .A2(n7147), .ZN(n7150) );
  AND2_X1 U8870 ( .A1(n7148), .A2(n8015), .ZN(n7149) );
  NAND2_X1 U8871 ( .A1(n7150), .A2(n7149), .ZN(n7156) );
  NAND2_X1 U8872 ( .A1(n7156), .A2(n7154), .ZN(n7151) );
  NAND2_X1 U8873 ( .A1(n7151), .A2(n9037), .ZN(n7167) );
  INV_X1 U8874 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n7161) );
  INV_X1 U8875 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10419) );
  NAND2_X1 U8876 ( .A1(n10367), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n10365) );
  INV_X1 U8877 ( .A(n10365), .ZN(n7152) );
  NAND2_X1 U8878 ( .A1(n7197), .A2(n7152), .ZN(n7198) );
  INV_X1 U8879 ( .A(n7204), .ZN(n7203) );
  NAND2_X1 U8880 ( .A1(n7203), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n7153) );
  AND2_X1 U8881 ( .A1(n7154), .A2(n8847), .ZN(n7155) );
  OAI211_X1 U8882 ( .C1(n7158), .C2(n7157), .A(n10366), .B(n4903), .ZN(n7160)
         );
  NAND2_X1 U8883 ( .A1(P2_U3152), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n7159) );
  OAI211_X1 U8884 ( .C1(n9131), .C2(n7161), .A(n7160), .B(n7159), .ZN(n7162)
         );
  AOI21_X1 U8885 ( .B1(n7214), .B2(n10362), .A(n7162), .ZN(n7171) );
  MUX2_X1 U8886 ( .A(n7163), .B(P2_REG2_REG_2__SCAN_IN), .S(n7223), .Z(n7169)
         );
  AND2_X1 U8887 ( .A1(P2_REG2_REG_0__SCAN_IN), .A2(n10367), .ZN(n7165) );
  OAI21_X1 U8888 ( .B1(n7164), .B2(n7204), .A(n7207), .ZN(n7168) );
  NOR2_X1 U8889 ( .A1(n8854), .A2(n8847), .ZN(n7166) );
  NAND2_X1 U8890 ( .A1(n7167), .A2(n7166), .ZN(n9124) );
  OAI211_X1 U8891 ( .C1(n7169), .C2(n7168), .A(n10361), .B(n7249), .ZN(n7170)
         );
  NAND2_X1 U8892 ( .A1(n7171), .A2(n7170), .ZN(P2_U3247) );
  XOR2_X1 U8893 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n7409), .Z(n7174) );
  NAND2_X1 U8894 ( .A1(n7173), .A2(n7174), .ZN(n7407) );
  OAI21_X1 U8895 ( .B1(n7174), .B2(n7173), .A(n7407), .ZN(n7183) );
  INV_X1 U8896 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10470) );
  NAND2_X1 U8897 ( .A1(n10294), .A2(n7409), .ZN(n7175) );
  NAND2_X1 U8898 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n8528) );
  OAI211_X1 U8899 ( .C1(n8719), .C2(n10470), .A(n7175), .B(n8528), .ZN(n7182)
         );
  XNOR2_X1 U8900 ( .A(n7409), .B(P1_REG2_REG_9__SCAN_IN), .ZN(n7180) );
  INV_X1 U8901 ( .A(n7411), .ZN(n7178) );
  AOI211_X1 U8902 ( .C1(n7180), .C2(n7179), .A(n9830), .B(n7178), .ZN(n7181)
         );
  AOI211_X1 U8903 ( .C1(n10302), .C2(n7183), .A(n7182), .B(n7181), .ZN(n7184)
         );
  INV_X1 U8904 ( .A(n7184), .ZN(P1_U3250) );
  NAND2_X1 U8905 ( .A1(n7186), .A2(n7185), .ZN(n7187) );
  OAI22_X1 U8906 ( .A1(n7188), .A2(n7187), .B1(n7463), .B2(n9952), .ZN(n7418)
         );
  AOI21_X1 U8907 ( .B1(n7422), .B2(n7189), .A(n7418), .ZN(n7213) );
  AND2_X1 U8908 ( .A1(n7191), .A2(n7190), .ZN(n7192) );
  AND2_X2 U8909 ( .A1(n7211), .A2(n7194), .ZN(n10353) );
  INV_X1 U8910 ( .A(n10353), .ZN(n10351) );
  INV_X1 U8911 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n7195) );
  OR2_X1 U8912 ( .A1(n10353), .A2(n7195), .ZN(n7196) );
  OAI21_X1 U8913 ( .B1(n7213), .B2(n10351), .A(n7196), .ZN(P1_U3454) );
  OAI22_X1 U8914 ( .A1(n9131), .A2(n10258), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7668), .ZN(n7202) );
  INV_X1 U8915 ( .A(n7197), .ZN(n7200) );
  INV_X1 U8916 ( .A(n7198), .ZN(n7199) );
  AOI211_X1 U8917 ( .C1(n10365), .C2(n7200), .A(n7199), .B(n9112), .ZN(n7201)
         );
  AOI211_X1 U8918 ( .C1(n10362), .C2(n7203), .A(n7202), .B(n7201), .ZN(n7209)
         );
  MUX2_X1 U8919 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n7164), .S(n7204), .Z(n7205)
         );
  OAI21_X1 U8920 ( .B1(n5166), .B2(n10359), .A(n7205), .ZN(n7206) );
  NAND3_X1 U8921 ( .A1(n10361), .A2(n7207), .A3(n7206), .ZN(n7208) );
  NAND2_X1 U8922 ( .A1(n7209), .A2(n7208), .ZN(P2_U3246) );
  AND2_X2 U8923 ( .A1(n7211), .A2(n7210), .ZN(n10357) );
  NAND2_X1 U8924 ( .A1(n10355), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n7212) );
  OAI21_X1 U8925 ( .B1(n7213), .B2(n10355), .A(n7212), .ZN(P1_U3523) );
  NAND2_X1 U8926 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3152), .ZN(n7647) );
  INV_X1 U8927 ( .A(n7647), .ZN(n7222) );
  INV_X1 U8928 ( .A(n7253), .ZN(n7216) );
  INV_X1 U8929 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n7215) );
  MUX2_X1 U8930 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n7215), .S(n7253), .Z(n7243)
         );
  AOI21_X1 U8931 ( .B1(n7216), .B2(P2_REG1_REG_3__SCAN_IN), .A(n7242), .ZN(
        n7272) );
  MUX2_X1 U8932 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n7217), .S(n7281), .Z(n7271)
         );
  NOR2_X1 U8933 ( .A1(n7272), .A2(n7271), .ZN(n7270) );
  INV_X1 U8934 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n7218) );
  MUX2_X1 U8935 ( .A(n7218), .B(P2_REG1_REG_5__SCAN_IN), .S(n7287), .Z(n7283)
         );
  NOR2_X1 U8936 ( .A1(n7284), .A2(n7283), .ZN(n7282) );
  AOI21_X1 U8937 ( .B1(n7287), .B2(P2_REG1_REG_5__SCAN_IN), .A(n7282), .ZN(
        n7220) );
  XNOR2_X1 U8938 ( .A(n7260), .B(P2_REG1_REG_6__SCAN_IN), .ZN(n7219) );
  AOI211_X1 U8939 ( .C1(n7220), .C2(n7219), .A(n9112), .B(n7254), .ZN(n7221)
         );
  AOI211_X1 U8940 ( .C1(n10358), .C2(P2_ADDR_REG_6__SCAN_IN), .A(n7222), .B(
        n7221), .ZN(n7239) );
  OR2_X1 U8941 ( .A1(n7223), .A2(n7163), .ZN(n7248) );
  NAND2_X1 U8942 ( .A1(n7249), .A2(n7248), .ZN(n7226) );
  MUX2_X1 U8943 ( .A(n7224), .B(P2_REG2_REG_3__SCAN_IN), .S(n7253), .Z(n7225)
         );
  OR2_X1 U8944 ( .A1(n7253), .A2(n7224), .ZN(n7276) );
  NAND2_X1 U8945 ( .A1(n7277), .A2(n7276), .ZN(n7228) );
  INV_X1 U8946 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n8070) );
  MUX2_X1 U8947 ( .A(n8070), .B(P2_REG2_REG_4__SCAN_IN), .S(n7281), .Z(n7227)
         );
  NAND2_X1 U8948 ( .A1(n7228), .A2(n7227), .ZN(n7290) );
  NAND2_X1 U8949 ( .A1(n7229), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n7289) );
  NAND2_X1 U8950 ( .A1(n7290), .A2(n7289), .ZN(n7231) );
  MUX2_X1 U8951 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n8088), .S(n7287), .Z(n7230)
         );
  NAND2_X1 U8952 ( .A1(n7287), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n7236) );
  NAND2_X1 U8953 ( .A1(n7292), .A2(n7236), .ZN(n7234) );
  MUX2_X1 U8954 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n7232), .S(n7260), .Z(n7233)
         );
  NAND2_X1 U8955 ( .A1(n7234), .A2(n7233), .ZN(n7265) );
  MUX2_X1 U8956 ( .A(n7232), .B(P2_REG2_REG_6__SCAN_IN), .S(n7260), .Z(n7235)
         );
  NAND3_X1 U8957 ( .A1(n7292), .A2(n7236), .A3(n7235), .ZN(n7237) );
  NAND3_X1 U8958 ( .A1(n10361), .A2(n7265), .A3(n7237), .ZN(n7238) );
  OAI211_X1 U8959 ( .C1(n9101), .C2(n7240), .A(n7239), .B(n7238), .ZN(P2_U3251) );
  INV_X1 U8960 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n7241) );
  NOR2_X1 U8961 ( .A1(n9131), .A2(n7241), .ZN(n7246) );
  AOI211_X1 U8962 ( .C1(n7244), .C2(n7243), .A(n7242), .B(n9112), .ZN(n7245)
         );
  AOI211_X1 U8963 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(P2_U3152), .A(n7246), .B(
        n7245), .ZN(n7252) );
  MUX2_X1 U8964 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n7224), .S(n7253), .Z(n7247)
         );
  NAND3_X1 U8965 ( .A1(n7249), .A2(n7248), .A3(n7247), .ZN(n7250) );
  NAND3_X1 U8966 ( .A1(n10361), .A2(n7277), .A3(n7250), .ZN(n7251) );
  OAI211_X1 U8967 ( .C1(n9101), .C2(n7253), .A(n7252), .B(n7251), .ZN(P2_U3248) );
  NOR2_X1 U8968 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8444), .ZN(n7259) );
  INV_X1 U8969 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n7255) );
  MUX2_X1 U8970 ( .A(n7255), .B(P2_REG1_REG_7__SCAN_IN), .S(n7387), .Z(n7256)
         );
  AOI211_X1 U8971 ( .C1(n7257), .C2(n7256), .A(n9112), .B(n7384), .ZN(n7258)
         );
  AOI211_X1 U8972 ( .C1(n10358), .C2(P2_ADDR_REG_7__SCAN_IN), .A(n7259), .B(
        n7258), .ZN(n7268) );
  NAND2_X1 U8973 ( .A1(n7260), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n7264) );
  NAND2_X1 U8974 ( .A1(n7265), .A2(n7264), .ZN(n7262) );
  MUX2_X1 U8975 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n7938), .S(n7387), .Z(n7261)
         );
  MUX2_X1 U8976 ( .A(n7938), .B(P2_REG2_REG_7__SCAN_IN), .S(n7387), .Z(n7263)
         );
  NAND3_X1 U8977 ( .A1(n7265), .A2(n7264), .A3(n7263), .ZN(n7266) );
  NAND3_X1 U8978 ( .A1(n10361), .A2(n7392), .A3(n7266), .ZN(n7267) );
  OAI211_X1 U8979 ( .C1(n9101), .C2(n7269), .A(n7268), .B(n7267), .ZN(P2_U3252) );
  NAND2_X1 U8980 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3152), .ZN(n7558) );
  INV_X1 U8981 ( .A(n7558), .ZN(n7274) );
  AOI211_X1 U8982 ( .C1(n7272), .C2(n7271), .A(n7270), .B(n9112), .ZN(n7273)
         );
  AOI211_X1 U8983 ( .C1(n10358), .C2(P2_ADDR_REG_4__SCAN_IN), .A(n7274), .B(
        n7273), .ZN(n7280) );
  MUX2_X1 U8984 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n8070), .S(n7281), .Z(n7275)
         );
  NAND3_X1 U8985 ( .A1(n7277), .A2(n7276), .A3(n7275), .ZN(n7278) );
  NAND3_X1 U8986 ( .A1(n10361), .A2(n7290), .A3(n7278), .ZN(n7279) );
  OAI211_X1 U8987 ( .C1(n9101), .C2(n7281), .A(n7280), .B(n7279), .ZN(P2_U3249) );
  NAND2_X1 U8988 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3152), .ZN(n7607) );
  INV_X1 U8989 ( .A(n7607), .ZN(n7286) );
  AOI211_X1 U8990 ( .C1(n7284), .C2(n7283), .A(n9112), .B(n7282), .ZN(n7285)
         );
  AOI211_X1 U8991 ( .C1(n10358), .C2(P2_ADDR_REG_5__SCAN_IN), .A(n7286), .B(
        n7285), .ZN(n7294) );
  MUX2_X1 U8992 ( .A(n8088), .B(P2_REG2_REG_5__SCAN_IN), .S(n7287), .Z(n7288)
         );
  NAND3_X1 U8993 ( .A1(n7290), .A2(n7289), .A3(n7288), .ZN(n7291) );
  NAND3_X1 U8994 ( .A1(n10361), .A2(n7292), .A3(n7291), .ZN(n7293) );
  OAI211_X1 U8995 ( .C1(n9101), .C2(n7295), .A(n7294), .B(n7293), .ZN(P2_U3250) );
  INV_X1 U8996 ( .A(n7296), .ZN(n7299) );
  AOI22_X1 U8997 ( .A1(n9107), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n7440), .ZN(n7297) );
  OAI21_X1 U8998 ( .B1(n7299), .B2(n9591), .A(n7297), .ZN(P2_U3341) );
  AOI22_X1 U8999 ( .A1(n9829), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n10239), .ZN(n7298) );
  OAI21_X1 U9000 ( .B1(n7299), .B2(n10244), .A(n7298), .ZN(P1_U3336) );
  INV_X1 U9001 ( .A(n7300), .ZN(n7302) );
  INV_X1 U9002 ( .A(n9087), .ZN(n9093) );
  OAI222_X1 U9003 ( .A1(n9586), .A2(n7301), .B1(n9591), .B2(n7302), .C1(n9093), 
        .C2(P2_U3152), .ZN(P2_U3342) );
  INV_X1 U9004 ( .A(n8713), .ZN(n9817) );
  OAI222_X1 U9005 ( .A1(n10251), .A2(n7303), .B1(P1_U3084), .B2(n9817), .C1(
        n7302), .C2(n10244), .ZN(P1_U3337) );
  OAI21_X1 U9006 ( .B1(n7306), .B2(n7305), .A(n7304), .ZN(n7307) );
  NAND2_X1 U9007 ( .A1(n7307), .A2(n8526), .ZN(n7311) );
  INV_X1 U9008 ( .A(n9758), .ZN(n9703) );
  INV_X1 U9009 ( .A(n4575), .ZN(n7308) );
  OAI22_X1 U9010 ( .A1(n9760), .A2(n4400), .B1(n9743), .B2(n7308), .ZN(n7309)
         );
  AOI21_X1 U9011 ( .B1(n9703), .B2(n6580), .A(n7309), .ZN(n7310) );
  OAI211_X1 U9012 ( .C1(n7313), .C2(n7312), .A(n7311), .B(n7310), .ZN(P1_U3220) );
  NAND2_X1 U9013 ( .A1(n7314), .A2(n7568), .ZN(n7341) );
  OAI21_X1 U9014 ( .B1(n7317), .B2(n7568), .A(n7341), .ZN(n8051) );
  NAND2_X1 U9015 ( .A1(n7316), .A2(n7595), .ZN(n7872) );
  OAI211_X1 U9016 ( .C1(n7316), .C2(n7595), .A(n10409), .B(n7872), .ZN(n8047)
         );
  OAI21_X1 U9017 ( .B1(n7316), .B2(n10403), .A(n8047), .ZN(n7320) );
  XOR2_X1 U9018 ( .A(n7317), .B(n7594), .Z(n7319) );
  AOI22_X1 U9019 ( .A1(n9412), .A2(n9036), .B1(n9411), .B2(n7318), .ZN(n7664)
         );
  OAI21_X1 U9020 ( .B1(n7319), .B2(n9406), .A(n7664), .ZN(n8050) );
  AOI211_X1 U9021 ( .C1(n10399), .C2(n8051), .A(n7320), .B(n8050), .ZN(n7366)
         );
  NAND2_X1 U9022 ( .A1(n10416), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n7321) );
  OAI21_X1 U9023 ( .B1(n10416), .B2(n7366), .A(n7321), .ZN(P2_U3454) );
  NAND2_X1 U9024 ( .A1(n7323), .A2(n4594), .ZN(n7327) );
  NOR2_X1 U9025 ( .A1(n7324), .A2(n7327), .ZN(n7325) );
  AOI211_X1 U9026 ( .C1(n7327), .C2(n7326), .A(n9778), .B(n7325), .ZN(n9781)
         );
  INV_X1 U9027 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n7328) );
  NOR2_X1 U9028 ( .A1(n8719), .A2(n7328), .ZN(n7340) );
  AOI211_X1 U9029 ( .C1(n7331), .C2(n7330), .A(n7329), .B(n9830), .ZN(n7339)
         );
  INV_X1 U9030 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n7472) );
  NAND2_X1 U9031 ( .A1(n10294), .A2(n7332), .ZN(n7337) );
  OAI211_X1 U9032 ( .C1(n7335), .C2(n7334), .A(n10302), .B(n7333), .ZN(n7336)
         );
  OAI211_X1 U9033 ( .C1(P1_STATE_REG_SCAN_IN), .C2(n7472), .A(n7337), .B(n7336), .ZN(n7338) );
  OR4_X1 U9034 ( .A1(n9781), .A2(n7340), .A3(n7339), .A4(n7338), .ZN(P1_U3243)
         );
  NAND2_X1 U9035 ( .A1(n7341), .A2(n5189), .ZN(n7343) );
  INV_X1 U9036 ( .A(n7888), .ZN(n10389) );
  OR2_X1 U9037 ( .A1(n9036), .A2(n10389), .ZN(n7344) );
  NAND2_X1 U9038 ( .A1(n7345), .A2(n7523), .ZN(n7349) );
  INV_X1 U9039 ( .A(n8491), .ZN(n7533) );
  OR2_X1 U9040 ( .A1(n7346), .A2(n7533), .ZN(n8054) );
  INV_X1 U9041 ( .A(n10394), .ZN(n8063) );
  OAI22_X1 U9042 ( .A1(n8065), .A2(n8054), .B1(n9035), .B2(n8063), .ZN(n7347)
         );
  INV_X1 U9043 ( .A(n7347), .ZN(n7348) );
  XNOR2_X1 U9044 ( .A(n7784), .B(n7785), .ZN(n8082) );
  NAND2_X1 U9045 ( .A1(n7351), .A2(n7350), .ZN(n7353) );
  INV_X1 U9046 ( .A(n7785), .ZN(n7352) );
  NAND2_X1 U9047 ( .A1(n7353), .A2(n7352), .ZN(n7354) );
  NAND2_X1 U9048 ( .A1(n7355), .A2(n7354), .ZN(n7358) );
  NAND2_X1 U9049 ( .A1(n9411), .A2(n9035), .ZN(n7356) );
  OAI21_X1 U9050 ( .B1(n7671), .B2(n9386), .A(n7356), .ZN(n7357) );
  AOI21_X1 U9051 ( .B1(n7358), .B2(n4402), .A(n7357), .ZN(n8089) );
  OAI21_X1 U9052 ( .B1(n8060), .B2(n7781), .A(n10409), .ZN(n7359) );
  OR2_X1 U9053 ( .A1(n8504), .A2(n7359), .ZN(n8083) );
  OAI211_X1 U9054 ( .C1(n7781), .C2(n10403), .A(n8089), .B(n8083), .ZN(n7360)
         );
  AOI21_X1 U9055 ( .B1(n10399), .B2(n8082), .A(n7360), .ZN(n7364) );
  OR2_X1 U9056 ( .A1(n10418), .A2(n5245), .ZN(n7361) );
  OAI21_X1 U9057 ( .B1(n7364), .B2(n10416), .A(n7361), .ZN(P2_U3466) );
  AND2_X2 U9058 ( .A1(n7362), .A2(n7870), .ZN(n10426) );
  NAND2_X1 U9059 ( .A1(n10424), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n7363) );
  OAI21_X1 U9060 ( .B1(n7364), .B2(n10424), .A(n7363), .ZN(P2_U3525) );
  NAND2_X1 U9061 ( .A1(n10424), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n7365) );
  OAI21_X1 U9062 ( .B1(n10424), .B2(n7366), .A(n7365), .ZN(P2_U3521) );
  INV_X1 U9063 ( .A(n10211), .ZN(n10347) );
  INV_X1 U9064 ( .A(n7377), .ZN(n7371) );
  OR2_X1 U9065 ( .A1(n7377), .A2(n7369), .ZN(n7462) );
  OAI21_X1 U9066 ( .B1(n7371), .B2(n7370), .A(n7462), .ZN(n7381) );
  INV_X1 U9067 ( .A(n7381), .ZN(n10313) );
  INV_X1 U9068 ( .A(n10207), .ZN(n10344) );
  OAI211_X1 U9069 ( .C1(n4400), .C2(n7372), .A(n10341), .B(n7470), .ZN(n10309)
         );
  OAI21_X1 U9070 ( .B1(n10344), .B2(n4400), .A(n10309), .ZN(n7382) );
  OR2_X1 U9071 ( .A1(n7373), .A2(n6713), .ZN(n7375) );
  OR2_X1 U9072 ( .A1(n7420), .A2(n7744), .ZN(n7374) );
  AOI22_X1 U9073 ( .A1(n6580), .A2(n10055), .B1(n10057), .B2(n4575), .ZN(n7380) );
  XNOR2_X1 U9074 ( .A(n7377), .B(n7376), .ZN(n7378) );
  NAND2_X1 U9075 ( .A1(n7378), .A2(n10099), .ZN(n7379) );
  OAI211_X1 U9076 ( .C1(n7381), .C2(n10040), .A(n7380), .B(n7379), .ZN(n10311)
         );
  AOI211_X1 U9077 ( .C1(n10347), .C2(n10313), .A(n7382), .B(n10311), .ZN(
        n10330) );
  NAND2_X1 U9078 ( .A1(n10355), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n7383) );
  OAI21_X1 U9079 ( .B1(n10330), .B2(n10355), .A(n7383), .ZN(P1_U3524) );
  XNOR2_X1 U9080 ( .A(n7494), .B(P2_REG1_REG_8__SCAN_IN), .ZN(n7385) );
  AOI211_X1 U9081 ( .C1(n7386), .C2(n7385), .A(n9112), .B(n7490), .ZN(n7395)
         );
  NAND2_X1 U9082 ( .A1(n7387), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n7391) );
  NAND2_X1 U9083 ( .A1(n7392), .A2(n7391), .ZN(n7389) );
  MUX2_X1 U9084 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n7995), .S(n7494), .Z(n7388)
         );
  NAND2_X1 U9085 ( .A1(n7389), .A2(n7388), .ZN(n7499) );
  MUX2_X1 U9086 ( .A(n7995), .B(P2_REG2_REG_8__SCAN_IN), .S(n7494), .Z(n7390)
         );
  NAND3_X1 U9087 ( .A1(n7392), .A2(n7391), .A3(n7390), .ZN(n7393) );
  AND3_X1 U9088 ( .A1(n10361), .A2(n7499), .A3(n7393), .ZN(n7394) );
  NOR2_X1 U9089 ( .A1(n7395), .A2(n7394), .ZN(n7398) );
  NAND2_X1 U9090 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3152), .ZN(n7776) );
  INV_X1 U9091 ( .A(n7776), .ZN(n7396) );
  AOI21_X1 U9092 ( .B1(n10358), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n7396), .ZN(
        n7397) );
  OAI211_X1 U9093 ( .C1(n7399), .C2(n9101), .A(n7398), .B(n7397), .ZN(P2_U3253) );
  XOR2_X1 U9094 ( .A(n7401), .B(n7400), .Z(n7406) );
  INV_X1 U9095 ( .A(n9779), .ZN(n7701) );
  AOI22_X1 U9096 ( .A1(n9755), .A2(n9780), .B1(n7469), .B2(n9734), .ZN(n7402)
         );
  OAI21_X1 U9097 ( .B1(n7701), .B2(n9758), .A(n7402), .ZN(n7403) );
  AOI21_X1 U9098 ( .B1(P1_REG3_REG_2__SCAN_IN), .B2(n7404), .A(n7403), .ZN(
        n7405) );
  OAI21_X1 U9099 ( .B1(n7406), .B2(n9765), .A(n7405), .ZN(P1_U3235) );
  XOR2_X1 U9100 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n7429), .Z(n7427) );
  XOR2_X1 U9101 ( .A(n7428), .B(n7427), .Z(n7417) );
  NAND2_X1 U9102 ( .A1(n10294), .A2(n7429), .ZN(n7408) );
  NAND2_X1 U9103 ( .A1(P1_U3084), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n8576) );
  NAND2_X1 U9104 ( .A1(n7408), .A2(n8576), .ZN(n7415) );
  NAND2_X1 U9105 ( .A1(n7409), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n7410) );
  XNOR2_X1 U9106 ( .A(n7429), .B(P1_REG2_REG_10__SCAN_IN), .ZN(n7412) );
  AOI211_X1 U9107 ( .C1(n7413), .C2(n7412), .A(n9830), .B(n4496), .ZN(n7414)
         );
  AOI211_X1 U9108 ( .C1(n10301), .C2(P1_ADDR_REG_10__SCAN_IN), .A(n7415), .B(
        n7414), .ZN(n7416) );
  OAI21_X1 U9109 ( .B1(n9823), .B2(n7417), .A(n7416), .ZN(P1_U3251) );
  AOI22_X1 U9110 ( .A1(n7418), .A2(n10315), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        n10307), .ZN(n7424) );
  INV_X1 U9111 ( .A(n10047), .ZN(n10064) );
  NOR2_X1 U9112 ( .A1(n7420), .A2(n7419), .ZN(n7421) );
  OAI21_X1 U9113 ( .B1(n10064), .B2(n10052), .A(n7422), .ZN(n7423) );
  OAI211_X1 U9114 ( .C1(n10315), .C2(n7425), .A(n7424), .B(n7423), .ZN(
        P1_U3291) );
  XNOR2_X1 U9115 ( .A(n7719), .B(P1_REG1_REG_11__SCAN_IN), .ZN(n7716) );
  INV_X1 U9116 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n8380) );
  XOR2_X1 U9117 ( .A(n7717), .B(n7716), .Z(n7438) );
  XOR2_X1 U9118 ( .A(P1_REG2_REG_11__SCAN_IN), .B(n7719), .Z(n7432) );
  OAI21_X1 U9119 ( .B1(n7432), .B2(n7431), .A(n7718), .ZN(n7436) );
  INV_X1 U9120 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n7434) );
  NAND2_X1 U9121 ( .A1(n10294), .A2(n7719), .ZN(n7433) );
  NAND2_X1 U9122 ( .A1(P1_U3084), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n8541) );
  OAI211_X1 U9123 ( .C1(n8719), .C2(n7434), .A(n7433), .B(n8541), .ZN(n7435)
         );
  AOI21_X1 U9124 ( .B1(n7436), .B2(n10292), .A(n7435), .ZN(n7437) );
  OAI21_X1 U9125 ( .B1(n9823), .B2(n7438), .A(n7437), .ZN(P1_U3252) );
  INV_X1 U9126 ( .A(n7439), .ZN(n7480) );
  AOI22_X1 U9127 ( .A1(n9120), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n7440), .ZN(n7441) );
  OAI21_X1 U9128 ( .B1(n7480), .B2(n9591), .A(n7441), .ZN(P2_U3340) );
  INV_X1 U9129 ( .A(n10040), .ZN(n7946) );
  NAND2_X1 U9130 ( .A1(n7443), .A2(n7444), .ZN(n7445) );
  NAND2_X1 U9131 ( .A1(n7442), .A2(n7445), .ZN(n7628) );
  INV_X1 U9132 ( .A(n10057), .ZN(n9954) );
  OAI22_X1 U9133 ( .A1(n7483), .A2(n9954), .B1(n7484), .B2(n9952), .ZN(n7451)
         );
  NAND2_X1 U9134 ( .A1(n4517), .A2(n7447), .ZN(n7449) );
  INV_X1 U9135 ( .A(n10099), .ZN(n9950) );
  AOI21_X1 U9136 ( .B1(n7446), .B2(n7449), .A(n9950), .ZN(n7450) );
  AOI211_X1 U9137 ( .C1(n7946), .C2(n7628), .A(n7451), .B(n7450), .ZN(n7632)
         );
  AND2_X1 U9138 ( .A1(n6713), .A2(n10310), .ZN(n10314) );
  NAND2_X1 U9139 ( .A1(n10315), .A2(n10314), .ZN(n10049) );
  INV_X1 U9140 ( .A(n10049), .ZN(n7962) );
  INV_X1 U9141 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n7452) );
  OAI22_X1 U9142 ( .A1(n10315), .A2(n7452), .B1(n9992), .B2(
        P1_REG3_REG_3__SCAN_IN), .ZN(n7453) );
  INV_X1 U9143 ( .A(n7453), .ZN(n7457) );
  OR2_X1 U9144 ( .A1(n7454), .A2(n7458), .ZN(n7455) );
  AND2_X1 U9145 ( .A1(n7708), .A2(n7455), .ZN(n7630) );
  NAND2_X1 U9146 ( .A1(n10052), .A2(n7630), .ZN(n7456) );
  OAI211_X1 U9147 ( .C1(n7458), .C2(n10047), .A(n7457), .B(n7456), .ZN(n7459)
         );
  AOI21_X1 U9148 ( .B1(n7962), .B2(n7628), .A(n7459), .ZN(n7460) );
  OAI21_X1 U9149 ( .B1(n7632), .B2(n10317), .A(n7460), .ZN(P1_U3288) );
  XOR2_X1 U9150 ( .A(n7461), .B(n7464), .Z(n7468) );
  AOI22_X1 U9151 ( .A1(n9780), .A2(n10057), .B1(n10055), .B2(n9779), .ZN(n7467) );
  OAI21_X1 U9152 ( .B1(n4400), .B2(n7463), .A(n7462), .ZN(n7465) );
  XNOR2_X1 U9153 ( .A(n7465), .B(n7464), .ZN(n7510) );
  NAND2_X1 U9154 ( .A1(n7510), .A2(n7946), .ZN(n7466) );
  OAI211_X1 U9155 ( .C1(n7468), .C2(n9950), .A(n7467), .B(n7466), .ZN(n7508)
         );
  AND2_X1 U9156 ( .A1(n7470), .A2(n7469), .ZN(n7471) );
  OR2_X1 U9157 ( .A1(n7471), .A2(n7454), .ZN(n7507) );
  INV_X1 U9158 ( .A(n7507), .ZN(n7475) );
  INV_X1 U9159 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n7473) );
  OAI22_X1 U9160 ( .A1(n10315), .A2(n7473), .B1(n7472), .B2(n9992), .ZN(n7474)
         );
  AOI21_X1 U9161 ( .B1(n10052), .B2(n7475), .A(n7474), .ZN(n7477) );
  NAND2_X1 U9162 ( .A1(n7510), .A2(n7962), .ZN(n7476) );
  OAI211_X1 U9163 ( .C1(n7506), .C2(n10047), .A(n7477), .B(n7476), .ZN(n7478)
         );
  AOI21_X1 U9164 ( .B1(n10315), .B2(n7508), .A(n7478), .ZN(n7479) );
  INV_X1 U9165 ( .A(n7479), .ZN(P1_U3289) );
  INV_X1 U9166 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n8329) );
  INV_X1 U9167 ( .A(n10293), .ZN(n8707) );
  OAI222_X1 U9168 ( .A1(n10251), .A2(n8329), .B1(n10244), .B2(n7480), .C1(
        P1_U3084), .C2(n8707), .ZN(P1_U3335) );
  XOR2_X1 U9169 ( .A(n7482), .B(n7481), .Z(n7489) );
  OAI22_X1 U9170 ( .A1(n7484), .A2(n9758), .B1(n9743), .B2(n7483), .ZN(n7485)
         );
  AOI211_X1 U9171 ( .C1(n7629), .C2(n9734), .A(n7486), .B(n7485), .ZN(n7488)
         );
  NAND2_X1 U9172 ( .A1(n9763), .A2(n8466), .ZN(n7487) );
  OAI211_X1 U9173 ( .C1(n7489), .C2(n9737), .A(n7488), .B(n7487), .ZN(P1_U3216) );
  XNOR2_X1 U9174 ( .A(n7731), .B(P2_REG1_REG_9__SCAN_IN), .ZN(n7491) );
  AOI211_X1 U9175 ( .C1(n7492), .C2(n7491), .A(n9112), .B(n7727), .ZN(n7505)
         );
  NAND2_X1 U9176 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3152), .ZN(n7925) );
  INV_X1 U9177 ( .A(n7925), .ZN(n7493) );
  AOI21_X1 U9178 ( .B1(n10358), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n7493), .ZN(
        n7502) );
  NAND2_X1 U9179 ( .A1(n7494), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n7498) );
  NAND2_X1 U9180 ( .A1(n7499), .A2(n7498), .ZN(n7496) );
  MUX2_X1 U9181 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n8005), .S(n7731), .Z(n7495)
         );
  MUX2_X1 U9182 ( .A(n8005), .B(P2_REG2_REG_9__SCAN_IN), .S(n7731), .Z(n7497)
         );
  NAND3_X1 U9183 ( .A1(n7499), .A2(n7498), .A3(n7497), .ZN(n7500) );
  NAND3_X1 U9184 ( .A1(n10361), .A2(n7737), .A3(n7500), .ZN(n7501) );
  OAI211_X1 U9185 ( .C1(n9101), .C2(n7503), .A(n7502), .B(n7501), .ZN(n7504)
         );
  OR2_X1 U9186 ( .A1(n7505), .A2(n7504), .ZN(P2_U3254) );
  OAI22_X1 U9187 ( .A1(n7507), .A2(n10334), .B1(n7506), .B2(n10344), .ZN(n7509) );
  AOI211_X1 U9188 ( .C1(n10347), .C2(n7510), .A(n7509), .B(n7508), .ZN(n10332)
         );
  NAND2_X1 U9189 ( .A1(n10355), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n7511) );
  OAI21_X1 U9190 ( .B1(n10332), .B2(n10355), .A(n7511), .ZN(P1_U3525) );
  XOR2_X1 U9191 ( .A(n7512), .B(n7514), .Z(n7513) );
  AOI222_X1 U9192 ( .A1(n10099), .A2(n7513), .B1(n9776), .B2(n10057), .C1(
        n9774), .C2(n10055), .ZN(n7683) );
  NAND2_X1 U9193 ( .A1(n7515), .A2(n7514), .ZN(n7829) );
  OAI21_X1 U9194 ( .B1(n7515), .B2(n7514), .A(n7829), .ZN(n7681) );
  INV_X1 U9195 ( .A(n10074), .ZN(n9938) );
  OAI211_X1 U9196 ( .C1(n7822), .C2(n7748), .A(n10341), .B(n7839), .ZN(n7679)
         );
  INV_X1 U9197 ( .A(n10077), .ZN(n7520) );
  INV_X1 U9198 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n7517) );
  INV_X1 U9199 ( .A(n7753), .ZN(n7516) );
  OAI22_X1 U9200 ( .A1(n10315), .A2(n7517), .B1(n7516), .B2(n9992), .ZN(n7518)
         );
  AOI21_X1 U9201 ( .B1(n10064), .B2(n5047), .A(n7518), .ZN(n7519) );
  OAI21_X1 U9202 ( .B1(n7679), .B2(n7520), .A(n7519), .ZN(n7521) );
  AOI21_X1 U9203 ( .B1(n7681), .B2(n9938), .A(n7521), .ZN(n7522) );
  OAI21_X1 U9204 ( .B1(n7683), .B2(n10317), .A(n7522), .ZN(P1_U3284) );
  INV_X1 U9205 ( .A(n7523), .ZN(n7524) );
  NOR2_X1 U9206 ( .A1(n7524), .A2(n7527), .ZN(n8056) );
  AOI21_X1 U9207 ( .B1(n7524), .B2(n7527), .A(n8056), .ZN(n8492) );
  OAI21_X1 U9208 ( .B1(n7527), .B2(n7526), .A(n7525), .ZN(n7530) );
  INV_X1 U9209 ( .A(n9035), .ZN(n7655) );
  OAI22_X1 U9210 ( .A1(n9384), .A2(n5164), .B1(n7655), .B2(n9386), .ZN(n7529)
         );
  NOR2_X1 U9211 ( .A1(n8492), .A2(n8560), .ZN(n7528) );
  AOI211_X1 U9212 ( .C1(n4402), .C2(n7530), .A(n7529), .B(n7528), .ZN(n8498)
         );
  NAND2_X1 U9213 ( .A1(n7874), .A2(n7533), .ZN(n7531) );
  NAND2_X1 U9214 ( .A1(n7531), .A2(n10409), .ZN(n7532) );
  NOR2_X1 U9215 ( .A1(n8058), .A2(n7532), .ZN(n8496) );
  AOI21_X1 U9216 ( .B1(n10408), .B2(n7533), .A(n8496), .ZN(n7534) );
  OAI211_X1 U9217 ( .C1(n8492), .C2(n9556), .A(n8498), .B(n7534), .ZN(n9558)
         );
  NAND2_X1 U9218 ( .A1(n9558), .A2(n10418), .ZN(n7535) );
  OAI21_X1 U9219 ( .B1(n10418), .B2(n5190), .A(n7535), .ZN(P2_U3460) );
  INV_X1 U9220 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7538) );
  INV_X1 U9221 ( .A(n7536), .ZN(n7539) );
  OAI222_X1 U9222 ( .A1(n8866), .A2(n7538), .B1(n9591), .B2(n7539), .C1(n7537), 
        .C2(P2_U3152), .ZN(P2_U3339) );
  INV_X1 U9223 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7540) );
  OAI222_X1 U9224 ( .A1(n10251), .A2(n7540), .B1(n10244), .B2(n7539), .C1(
        P1_U3084), .C2(n9962), .ZN(P1_U3334) );
  INV_X1 U9225 ( .A(n8061), .ZN(n7563) );
  NAND2_X1 U9226 ( .A1(n7870), .A2(n7867), .ZN(n7544) );
  NAND2_X1 U9227 ( .A1(n7544), .A2(n10403), .ZN(n7551) );
  NAND2_X1 U9228 ( .A1(n7544), .A2(n7543), .ZN(n7550) );
  INV_X1 U9229 ( .A(n7545), .ZN(n7547) );
  AND3_X1 U9230 ( .A1(n7548), .A2(n7547), .A3(n7546), .ZN(n7549) );
  NAND3_X1 U9231 ( .A1(n7551), .A2(n7550), .A3(n7549), .ZN(n7552) );
  AND2_X1 U9232 ( .A1(n10373), .A2(n7867), .ZN(n7553) );
  NAND2_X1 U9233 ( .A1(n7870), .A2(n7553), .ZN(n7590) );
  NOR2_X1 U9234 ( .A1(n7554), .A2(n5926), .ZN(n7883) );
  INV_X1 U9235 ( .A(n7883), .ZN(n7555) );
  OR2_X1 U9236 ( .A1(n7590), .A2(n7555), .ZN(n7557) );
  NAND2_X1 U9237 ( .A1(n9019), .A2(n8063), .ZN(n7559) );
  NAND2_X1 U9238 ( .A1(n7559), .A2(n7558), .ZN(n7562) );
  INV_X1 U9239 ( .A(n7346), .ZN(n7560) );
  OAI22_X1 U9240 ( .A1(n7560), .A2(n8992), .B1(n9017), .B2(n7782), .ZN(n7561)
         );
  AOI211_X1 U9241 ( .C1(n7563), .C2(n9014), .A(n7562), .B(n7561), .ZN(n7593)
         );
  NAND2_X1 U9242 ( .A1(n7564), .A2(n7757), .ZN(n7565) );
  XNOR2_X1 U9243 ( .A(n7583), .B(n7316), .ZN(n7567) );
  NAND2_X1 U9244 ( .A1(n8788), .A2(n7141), .ZN(n7566) );
  NAND2_X1 U9245 ( .A1(n7567), .A2(n7566), .ZN(n7571) );
  OR2_X1 U9246 ( .A1(n7583), .A2(n5070), .ZN(n7570) );
  NAND2_X1 U9247 ( .A1(n7570), .A2(n7569), .ZN(n7662) );
  XNOR2_X1 U9248 ( .A(n7888), .B(n7583), .ZN(n7572) );
  NAND2_X1 U9249 ( .A1(n8788), .A2(n9036), .ZN(n7573) );
  NAND2_X1 U9250 ( .A1(n7572), .A2(n7573), .ZN(n7577) );
  INV_X1 U9251 ( .A(n7572), .ZN(n7575) );
  INV_X1 U9252 ( .A(n7573), .ZN(n7574) );
  NAND2_X1 U9253 ( .A1(n7575), .A2(n7574), .ZN(n7576) );
  AND2_X1 U9254 ( .A1(n7577), .A2(n7576), .ZN(n7688) );
  NAND2_X1 U9255 ( .A1(n7687), .A2(n7688), .ZN(n7686) );
  NAND2_X1 U9256 ( .A1(n7686), .A2(n7577), .ZN(n7654) );
  XNOR2_X1 U9257 ( .A(n7583), .B(n8491), .ZN(n7578) );
  NAND2_X1 U9258 ( .A1(n8788), .A2(n7346), .ZN(n7579) );
  XNOR2_X1 U9259 ( .A(n7578), .B(n7579), .ZN(n7653) );
  INV_X1 U9260 ( .A(n7578), .ZN(n7581) );
  INV_X1 U9261 ( .A(n7579), .ZN(n7580) );
  NAND2_X1 U9262 ( .A1(n7581), .A2(n7580), .ZN(n7582) );
  XNOR2_X1 U9263 ( .A(n8820), .B(n10394), .ZN(n7584) );
  NAND2_X1 U9264 ( .A1(n8788), .A2(n9035), .ZN(n7585) );
  NAND2_X1 U9265 ( .A1(n7584), .A2(n7585), .ZN(n7617) );
  OAI21_X1 U9266 ( .B1(n7588), .B2(n7587), .A(n7618), .ZN(n7591) );
  NAND2_X1 U9267 ( .A1(n7591), .A2(n9011), .ZN(n7592) );
  NAND2_X1 U9268 ( .A1(n7593), .A2(n7592), .ZN(P2_U3232) );
  NOR2_X1 U9269 ( .A1(n9014), .A2(P2_U3152), .ZN(n7693) );
  OAI21_X1 U9270 ( .B1(n8788), .B2(n7595), .A(n7594), .ZN(n7596) );
  AOI22_X1 U9271 ( .A1(n9011), .A2(n7596), .B1(n9019), .B2(n5070), .ZN(n7600)
         );
  NAND2_X1 U9272 ( .A1(n9011), .A2(n8788), .ZN(n8984) );
  INV_X1 U9273 ( .A(n8984), .ZN(n8790) );
  INV_X1 U9274 ( .A(n7597), .ZN(n7598) );
  AOI22_X1 U9275 ( .A1(n8790), .A2(n7598), .B1(n8990), .B2(n7141), .ZN(n7599)
         );
  OAI211_X1 U9276 ( .C1(n7693), .C2(n8025), .A(n7600), .B(n7599), .ZN(P2_U3234) );
  XOR2_X1 U9277 ( .A(n7602), .B(n7601), .Z(n7606) );
  AOI22_X1 U9278 ( .A1(n9703), .A2(n8209), .B1(n9755), .B2(n9779), .ZN(n7603)
         );
  NAND2_X1 U9279 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3084), .ZN(n9782) );
  OAI211_X1 U9280 ( .C1(n10333), .C2(n9760), .A(n7603), .B(n9782), .ZN(n7604)
         );
  AOI21_X1 U9281 ( .B1(n7710), .B2(n9763), .A(n7604), .ZN(n7605) );
  OAI21_X1 U9282 ( .B1(n7606), .B2(n9737), .A(n7605), .ZN(P1_U3228) );
  INV_X1 U9283 ( .A(n8086), .ZN(n7611) );
  NAND2_X1 U9284 ( .A1(n9019), .A2(n4809), .ZN(n7608) );
  NAND2_X1 U9285 ( .A1(n7608), .A2(n7607), .ZN(n7610) );
  OAI22_X1 U9286 ( .A1(n7655), .A2(n8992), .B1(n9017), .B2(n7671), .ZN(n7609)
         );
  AOI211_X1 U9287 ( .C1(n7611), .C2(n9014), .A(n7610), .B(n7609), .ZN(n7623)
         );
  XNOR2_X1 U9288 ( .A(n8820), .B(n7781), .ZN(n7612) );
  NAND2_X1 U9289 ( .A1(n7612), .A2(n7613), .ZN(n7641) );
  INV_X1 U9290 ( .A(n7612), .ZN(n7615) );
  INV_X1 U9291 ( .A(n7613), .ZN(n7614) );
  NAND2_X1 U9292 ( .A1(n7615), .A2(n7614), .ZN(n7616) );
  AND2_X1 U9293 ( .A1(n7641), .A2(n7616), .ZN(n7620) );
  OAI21_X1 U9294 ( .B1(n7620), .B2(n7619), .A(n7642), .ZN(n7621) );
  NAND2_X1 U9295 ( .A1(n7621), .A2(n9011), .ZN(n7622) );
  NAND2_X1 U9296 ( .A1(n7623), .A2(n7622), .ZN(P2_U3229) );
  INV_X1 U9297 ( .A(n7624), .ZN(n7626) );
  OAI222_X1 U9298 ( .A1(n8866), .A2(n8454), .B1(n9591), .B2(n7626), .C1(
        P2_U3152), .C2(n5926), .ZN(P2_U3338) );
  OAI222_X1 U9299 ( .A1(n10251), .A2(n7627), .B1(n10244), .B2(n7626), .C1(
        P1_U3084), .C2(n4377), .ZN(P1_U3333) );
  INV_X1 U9300 ( .A(n7628), .ZN(n7633) );
  AOI22_X1 U9301 ( .A1(n7630), .A2(n10341), .B1(n10207), .B2(n7629), .ZN(n7631) );
  OAI211_X1 U9302 ( .C1(n7633), .C2(n10211), .A(n7632), .B(n7631), .ZN(n7635)
         );
  NAND2_X1 U9303 ( .A1(n7635), .A2(n10357), .ZN(n7634) );
  OAI21_X1 U9304 ( .B1(n10357), .B2(n7001), .A(n7634), .ZN(P1_U3526) );
  INV_X1 U9305 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n7637) );
  NAND2_X1 U9306 ( .A1(n7635), .A2(n10353), .ZN(n7636) );
  OAI21_X1 U9307 ( .B1(n10353), .B2(n7637), .A(n7636), .ZN(P1_U3463) );
  XNOR2_X1 U9308 ( .A(n8820), .B(n8506), .ZN(n7639) );
  NOR2_X1 U9309 ( .A1(n7671), .A2(n8819), .ZN(n7638) );
  OR2_X1 U9310 ( .A1(n7639), .A2(n7638), .ZN(n7669) );
  NAND2_X1 U9311 ( .A1(n7639), .A2(n7638), .ZN(n7640) );
  AND2_X1 U9312 ( .A1(n7669), .A2(n7640), .ZN(n7644) );
  OAI21_X1 U9313 ( .B1(n7644), .B2(n4552), .A(n7670), .ZN(n7645) );
  NAND2_X1 U9314 ( .A1(n7645), .A2(n9011), .ZN(n7652) );
  INV_X1 U9315 ( .A(n7646), .ZN(n8505) );
  NAND2_X1 U9316 ( .A1(n9019), .A2(n8506), .ZN(n7648) );
  NAND2_X1 U9317 ( .A1(n7648), .A2(n7647), .ZN(n7650) );
  OAI22_X1 U9318 ( .A1(n7782), .A2(n8992), .B1(n9017), .B2(n7987), .ZN(n7649)
         );
  AOI211_X1 U9319 ( .C1(n8505), .C2(n9014), .A(n7650), .B(n7649), .ZN(n7651)
         );
  NAND2_X1 U9320 ( .A1(n7652), .A2(n7651), .ZN(P2_U3241) );
  XNOR2_X1 U9321 ( .A(n7654), .B(n7653), .ZN(n7659) );
  OAI22_X1 U9322 ( .A1(n8996), .A2(n8491), .B1(n9017), .B2(n7655), .ZN(n7657)
         );
  MUX2_X1 U9323 ( .A(n9014), .B(P2_U3152), .S(P2_REG3_REG_3__SCAN_IN), .Z(
        n7656) );
  AOI211_X1 U9324 ( .C1(n9013), .C2(n9036), .A(n7657), .B(n7656), .ZN(n7658)
         );
  OAI21_X1 U9325 ( .B1(n7659), .B2(n7677), .A(n7658), .ZN(P2_U3220) );
  INV_X1 U9326 ( .A(n7660), .ZN(n7661) );
  AOI21_X1 U9327 ( .B1(n7663), .B2(n7662), .A(n7661), .ZN(n7665) );
  OAI22_X1 U9328 ( .A1(n7665), .A2(n7677), .B1(n8999), .B2(n7664), .ZN(n7666)
         );
  AOI21_X1 U9329 ( .B1(n5189), .B2(n9019), .A(n7666), .ZN(n7667) );
  OAI21_X1 U9330 ( .B1(n7693), .B2(n7668), .A(n7667), .ZN(P2_U3224) );
  XNOR2_X1 U9331 ( .A(n10407), .B(n8820), .ZN(n7773) );
  NOR2_X1 U9332 ( .A1(n7987), .A2(n8819), .ZN(n7772) );
  XNOR2_X1 U9333 ( .A(n7773), .B(n7772), .ZN(n7774) );
  XNOR2_X1 U9334 ( .A(n7775), .B(n7774), .ZN(n7678) );
  INV_X1 U9335 ( .A(n7941), .ZN(n7675) );
  INV_X1 U9336 ( .A(n7671), .ZN(n9034) );
  NAND2_X1 U9337 ( .A1(n9013), .A2(n9034), .ZN(n7673) );
  AOI22_X1 U9338 ( .A1(n9019), .A2(n10407), .B1(P2_REG3_REG_7__SCAN_IN), .B2(
        P2_U3152), .ZN(n7672) );
  OAI211_X1 U9339 ( .C1(n7936), .C2(n9017), .A(n7673), .B(n7672), .ZN(n7674)
         );
  AOI21_X1 U9340 ( .B1(n7675), .B2(n9014), .A(n7674), .ZN(n7676) );
  OAI21_X1 U9341 ( .B1(n7678), .B2(n7677), .A(n7676), .ZN(P2_U3215) );
  INV_X1 U9342 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n7685) );
  NAND2_X1 U9343 ( .A1(n10040), .A2(n10211), .ZN(n10134) );
  OAI21_X1 U9344 ( .B1(n7748), .B2(n10344), .A(n7679), .ZN(n7680) );
  AOI21_X1 U9345 ( .B1(n7681), .B2(n10134), .A(n7680), .ZN(n7682) );
  NAND2_X1 U9346 ( .A1(n7683), .A2(n7682), .ZN(n7694) );
  NAND2_X1 U9347 ( .A1(n7694), .A2(n10357), .ZN(n7684) );
  OAI21_X1 U9348 ( .B1(n10357), .B2(n7685), .A(n7684), .ZN(P1_U3530) );
  OAI21_X1 U9349 ( .B1(n7688), .B2(n7687), .A(n7686), .ZN(n7691) );
  AOI22_X1 U9350 ( .A1(n8990), .A2(n7346), .B1(n10389), .B2(n9019), .ZN(n7689)
         );
  OAI21_X1 U9351 ( .B1(n5188), .B2(n8992), .A(n7689), .ZN(n7690) );
  AOI21_X1 U9352 ( .B1(n9011), .B2(n7691), .A(n7690), .ZN(n7692) );
  OAI21_X1 U9353 ( .B1(n7693), .B2(n8248), .A(n7692), .ZN(P2_U3239) );
  INV_X1 U9354 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n7696) );
  NAND2_X1 U9355 ( .A1(n7694), .A2(n10353), .ZN(n7695) );
  OAI21_X1 U9356 ( .B1(n10353), .B2(n7696), .A(n7695), .ZN(P1_U3475) );
  NAND2_X1 U9357 ( .A1(n7442), .A2(n7697), .ZN(n7699) );
  NAND2_X1 U9358 ( .A1(n7699), .A2(n4781), .ZN(n7763) );
  OAI21_X1 U9359 ( .B1(n7699), .B2(n4781), .A(n7763), .ZN(n10339) );
  INV_X1 U9360 ( .A(n8209), .ZN(n7700) );
  OAI22_X1 U9361 ( .A1(n7701), .A2(n9954), .B1(n7700), .B2(n9952), .ZN(n7706)
         );
  NAND3_X1 U9362 ( .A1(n7446), .A2(n4781), .A3(n7702), .ZN(n7703) );
  AOI21_X1 U9363 ( .B1(n7704), .B2(n7703), .A(n9950), .ZN(n7705) );
  AOI211_X1 U9364 ( .C1(n7946), .C2(n10339), .A(n7706), .B(n7705), .ZN(n10336)
         );
  INV_X1 U9365 ( .A(n10052), .ZN(n9936) );
  NAND2_X1 U9366 ( .A1(n7708), .A2(n7711), .ZN(n7709) );
  NAND2_X1 U9367 ( .A1(n7707), .A2(n7709), .ZN(n10335) );
  AOI22_X1 U9368 ( .A1(n10317), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n7710), .B2(
        n10307), .ZN(n7713) );
  NAND2_X1 U9369 ( .A1(n10064), .A2(n7711), .ZN(n7712) );
  OAI211_X1 U9370 ( .C1(n9936), .C2(n10335), .A(n7713), .B(n7712), .ZN(n7714)
         );
  AOI21_X1 U9371 ( .B1(n10339), .B2(n7962), .A(n7714), .ZN(n7715) );
  OAI21_X1 U9372 ( .B1(n10336), .B2(n10317), .A(n7715), .ZN(P1_U3287) );
  XOR2_X1 U9373 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n7858), .Z(n7855) );
  OAI22_X1 U9374 ( .A1(n7717), .A2(n7716), .B1(P1_REG1_REG_11__SCAN_IN), .B2(
        n7719), .ZN(n7856) );
  XOR2_X1 U9375 ( .A(n7855), .B(n7856), .Z(n7726) );
  NAND2_X1 U9376 ( .A1(P1_U3084), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n8587) );
  OAI21_X1 U9377 ( .B1(n9818), .B2(n7854), .A(n8587), .ZN(n7724) );
  XNOR2_X1 U9378 ( .A(n7858), .B(P1_REG2_REG_12__SCAN_IN), .ZN(n7722) );
  INV_X1 U9379 ( .A(n7860), .ZN(n7720) );
  AOI211_X1 U9380 ( .C1(n7722), .C2(n7721), .A(n9830), .B(n7720), .ZN(n7723)
         );
  AOI211_X1 U9381 ( .C1(n10301), .C2(P1_ADDR_REG_12__SCAN_IN), .A(n7724), .B(
        n7723), .ZN(n7725) );
  OAI21_X1 U9382 ( .B1(n9823), .B2(n7726), .A(n7725), .ZN(P1_U3253) );
  XNOR2_X1 U9383 ( .A(n8142), .B(P2_REG1_REG_10__SCAN_IN), .ZN(n7728) );
  AOI211_X1 U9384 ( .C1(n7729), .C2(n7728), .A(n9112), .B(n8138), .ZN(n7743)
         );
  NOR2_X1 U9385 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8247), .ZN(n7730) );
  AOI21_X1 U9386 ( .B1(n10358), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n7730), .ZN(
        n7740) );
  NAND2_X1 U9387 ( .A1(n7731), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n7736) );
  NAND2_X1 U9388 ( .A1(n7737), .A2(n7736), .ZN(n7734) );
  MUX2_X1 U9389 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n7732), .S(n8142), .Z(n7733)
         );
  NAND2_X1 U9390 ( .A1(n7734), .A2(n7733), .ZN(n8144) );
  MUX2_X1 U9391 ( .A(n7732), .B(P2_REG2_REG_10__SCAN_IN), .S(n8142), .Z(n7735)
         );
  NAND3_X1 U9392 ( .A1(n7737), .A2(n7736), .A3(n7735), .ZN(n7738) );
  NAND3_X1 U9393 ( .A1(n10361), .A2(n8144), .A3(n7738), .ZN(n7739) );
  OAI211_X1 U9394 ( .C1(n9101), .C2(n7741), .A(n7740), .B(n7739), .ZN(n7742)
         );
  OR2_X1 U9395 ( .A1(n7743), .A2(n7742), .ZN(P2_U3255) );
  INV_X1 U9396 ( .A(n6261), .ZN(n7756) );
  OAI222_X1 U9397 ( .A1(n10251), .A2(n7745), .B1(n10244), .B2(n7756), .C1(
        n7744), .C2(P1_U3084), .ZN(P1_U3332) );
  XOR2_X1 U9398 ( .A(n7747), .B(n7746), .Z(n7755) );
  NOR2_X1 U9399 ( .A1(n9760), .A2(n7748), .ZN(n7752) );
  NAND2_X1 U9400 ( .A1(n9755), .A2(n9776), .ZN(n7750) );
  OAI211_X1 U9401 ( .C1(n8530), .C2(n9758), .A(n7750), .B(n7749), .ZN(n7751)
         );
  AOI211_X1 U9402 ( .C1(n7753), .C2(n9763), .A(n7752), .B(n7751), .ZN(n7754)
         );
  OAI21_X1 U9403 ( .B1(n7755), .B2(n9765), .A(n7754), .ZN(P1_U3211) );
  OAI222_X1 U9404 ( .A1(n8866), .A2(n7758), .B1(P2_U3152), .B2(n7757), .C1(
        n9591), .C2(n7756), .ZN(P2_U3337) );
  XNOR2_X1 U9405 ( .A(n7759), .B(n7764), .ZN(n7760) );
  AOI222_X1 U9406 ( .A1(n10099), .A2(n7760), .B1(n9777), .B2(n10057), .C1(
        n9776), .C2(n10055), .ZN(n7906) );
  AOI21_X1 U9407 ( .B1(n7903), .B2(n7707), .A(n5045), .ZN(n7904) );
  AOI22_X1 U9408 ( .A1(n10317), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n7850), .B2(
        n10307), .ZN(n7761) );
  OAI21_X1 U9409 ( .B1(n7848), .B2(n10047), .A(n7761), .ZN(n7770) );
  NAND2_X1 U9410 ( .A1(n7763), .A2(n7762), .ZN(n7765) );
  NAND2_X1 U9411 ( .A1(n7765), .A2(n7764), .ZN(n7768) );
  OR2_X1 U9412 ( .A1(n7767), .A2(n7766), .ZN(n7810) );
  NAND2_X1 U9413 ( .A1(n7768), .A2(n7810), .ZN(n7907) );
  NOR2_X1 U9414 ( .A1(n7907), .A2(n10074), .ZN(n7769) );
  AOI211_X1 U9415 ( .C1(n7904), .C2(n10052), .A(n7770), .B(n7769), .ZN(n7771)
         );
  OAI21_X1 U9416 ( .B1(n7906), .B2(n10317), .A(n7771), .ZN(P1_U3286) );
  XNOR2_X1 U9417 ( .A(n9552), .B(n8787), .ZN(n7914) );
  NOR2_X1 U9418 ( .A1(n7936), .A2(n8819), .ZN(n7915) );
  XNOR2_X1 U9419 ( .A(n7914), .B(n7915), .ZN(n7912) );
  XNOR2_X1 U9420 ( .A(n7913), .B(n7912), .ZN(n7780) );
  OAI21_X1 U9421 ( .B1(n9017), .B2(n7986), .A(n7776), .ZN(n7778) );
  INV_X1 U9422 ( .A(n9552), .ZN(n7999) );
  OAI22_X1 U9423 ( .A1(n7999), .A2(n8996), .B1(n9002), .B2(n7998), .ZN(n7777)
         );
  AOI211_X1 U9424 ( .C1(n9013), .C2(n9033), .A(n7778), .B(n7777), .ZN(n7779)
         );
  OAI21_X1 U9425 ( .B1(n7780), .B2(n7677), .A(n7779), .ZN(P2_U3223) );
  INV_X1 U9426 ( .A(n9556), .ZN(n7805) );
  NAND2_X1 U9427 ( .A1(n7782), .A2(n7781), .ZN(n8507) );
  NAND3_X1 U9428 ( .A1(n8509), .A2(n7785), .A3(n4809), .ZN(n7787) );
  NAND2_X1 U9429 ( .A1(n9034), .A2(n8506), .ZN(n7786) );
  AND2_X1 U9430 ( .A1(n7787), .A2(n7786), .ZN(n7788) );
  OR2_X1 U9431 ( .A1(n10407), .A2(n9033), .ZN(n7790) );
  INV_X1 U9432 ( .A(n7794), .ZN(n7793) );
  INV_X1 U9433 ( .A(n7797), .ZN(n7792) );
  NAND2_X1 U9434 ( .A1(n7794), .A2(n7797), .ZN(n7795) );
  NAND2_X1 U9435 ( .A1(n7967), .A2(n7795), .ZN(n8003) );
  INV_X1 U9436 ( .A(n8506), .ZN(n10404) );
  INV_X1 U9437 ( .A(n7965), .ZN(n8008) );
  NOR2_X1 U9438 ( .A1(n7996), .A2(n8008), .ZN(n7796) );
  OR2_X1 U9439 ( .A1(n7980), .A2(n7796), .ZN(n8006) );
  OAI22_X1 U9440 ( .A1(n8006), .A2(n9518), .B1(n8008), .B2(n10403), .ZN(n7804)
         );
  XNOR2_X1 U9441 ( .A(n7798), .B(n7797), .ZN(n7799) );
  NAND2_X1 U9442 ( .A1(n7799), .A2(n4402), .ZN(n7802) );
  INV_X1 U9443 ( .A(n8560), .ZN(n9394) );
  OAI22_X1 U9444 ( .A1(n9384), .A2(n7936), .B1(n8159), .B2(n9386), .ZN(n7800)
         );
  AOI21_X1 U9445 ( .B1(n8003), .B2(n9394), .A(n7800), .ZN(n7801) );
  AND2_X1 U9446 ( .A1(n7802), .A2(n7801), .ZN(n8004) );
  INV_X1 U9447 ( .A(n8004), .ZN(n7803) );
  AOI211_X1 U9448 ( .C1(n7805), .C2(n8003), .A(n7804), .B(n7803), .ZN(n7808)
         );
  NAND2_X1 U9449 ( .A1(n10416), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n7806) );
  OAI21_X1 U9450 ( .B1(n7808), .B2(n10416), .A(n7806), .ZN(P2_U3478) );
  NAND2_X1 U9451 ( .A1(n10424), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n7807) );
  OAI21_X1 U9452 ( .B1(n7808), .B2(n10424), .A(n7807), .ZN(P2_U3529) );
  NAND2_X1 U9453 ( .A1(n7810), .A2(n7809), .ZN(n7811) );
  XNOR2_X1 U9454 ( .A(n7811), .B(n4774), .ZN(n10348) );
  INV_X1 U9455 ( .A(n10348), .ZN(n7827) );
  XNOR2_X1 U9456 ( .A(n7813), .B(n7812), .ZN(n7814) );
  NAND2_X1 U9457 ( .A1(n7814), .A2(n10099), .ZN(n7818) );
  NAND2_X1 U9458 ( .A1(n10057), .A2(n8209), .ZN(n7815) );
  OAI21_X1 U9459 ( .B1(n8207), .B2(n9952), .A(n7815), .ZN(n7816) );
  AOI21_X1 U9460 ( .B1(n10348), .B2(n7946), .A(n7816), .ZN(n7817) );
  AND2_X1 U9461 ( .A1(n7818), .A2(n7817), .ZN(n10350) );
  MUX2_X1 U9462 ( .A(n10350), .B(n7011), .S(n10317), .Z(n7826) );
  AND2_X1 U9463 ( .A1(n7820), .A2(n7819), .ZN(n7821) );
  NOR2_X1 U9464 ( .A1(n7822), .A2(n7821), .ZN(n10342) );
  INV_X1 U9465 ( .A(n8212), .ZN(n7823) );
  OAI22_X1 U9466 ( .A1(n10047), .A2(n10345), .B1(n7823), .B2(n9992), .ZN(n7824) );
  AOI21_X1 U9467 ( .B1(n10342), .B2(n10052), .A(n7824), .ZN(n7825) );
  OAI211_X1 U9468 ( .C1(n7827), .C2(n10049), .A(n7826), .B(n7825), .ZN(
        P1_U3285) );
  NAND2_X1 U9469 ( .A1(n7829), .A2(n7828), .ZN(n7830) );
  XNOR2_X1 U9470 ( .A(n7830), .B(n7831), .ZN(n10212) );
  XNOR2_X1 U9471 ( .A(n7832), .B(n7831), .ZN(n7835) );
  AOI22_X1 U9472 ( .A1(n9775), .A2(n10057), .B1(n10055), .B2(n9773), .ZN(n7833) );
  OAI21_X1 U9473 ( .B1(n10212), .B2(n10040), .A(n7833), .ZN(n7834) );
  AOI21_X1 U9474 ( .B1(n7835), .B2(n10099), .A(n7834), .ZN(n10210) );
  MUX2_X1 U9475 ( .A(n7836), .B(n10210), .S(n10315), .Z(n7843) );
  INV_X1 U9476 ( .A(n7837), .ZN(n7838) );
  AOI21_X1 U9477 ( .B1(n10206), .B2(n7839), .A(n7838), .ZN(n10208) );
  INV_X1 U9478 ( .A(n8111), .ZN(n7840) );
  OAI22_X1 U9479 ( .A1(n10047), .A2(n5044), .B1(n9992), .B2(n7840), .ZN(n7841)
         );
  AOI21_X1 U9480 ( .B1(n10208), .B2(n10052), .A(n7841), .ZN(n7842) );
  OAI211_X1 U9481 ( .C1(n10212), .C2(n10049), .A(n7843), .B(n7842), .ZN(
        P1_U3283) );
  XNOR2_X1 U9482 ( .A(n8200), .B(n8201), .ZN(n7845) );
  NOR2_X1 U9483 ( .A1(n7845), .A2(n7844), .ZN(n8199) );
  AOI21_X1 U9484 ( .B1(n7845), .B2(n7844), .A(n8199), .ZN(n7852) );
  AOI22_X1 U9485 ( .A1(n9703), .A2(n9776), .B1(n9755), .B2(n9777), .ZN(n7847)
         );
  OAI211_X1 U9486 ( .C1(n7848), .C2(n9760), .A(n7847), .B(n7846), .ZN(n7849)
         );
  AOI21_X1 U9487 ( .B1(n7850), .B2(n9763), .A(n7849), .ZN(n7851) );
  OAI21_X1 U9488 ( .B1(n7852), .B2(n9737), .A(n7851), .ZN(P1_U3225) );
  XNOR2_X1 U9489 ( .A(n8632), .B(P1_REG1_REG_13__SCAN_IN), .ZN(n8625) );
  INV_X1 U9490 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n7853) );
  XOR2_X1 U9491 ( .A(n8625), .B(n8626), .Z(n7866) );
  NAND2_X1 U9492 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9704) );
  OAI21_X1 U9493 ( .B1(n9818), .B2(n7857), .A(n9704), .ZN(n7864) );
  NAND2_X1 U9494 ( .A1(n7858), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n7859) );
  XNOR2_X1 U9495 ( .A(n8632), .B(P1_REG2_REG_13__SCAN_IN), .ZN(n7861) );
  AOI211_X1 U9496 ( .C1(n7862), .C2(n7861), .A(n9830), .B(n8633), .ZN(n7863)
         );
  AOI211_X1 U9497 ( .C1(n10301), .C2(P1_ADDR_REG_13__SCAN_IN), .A(n7864), .B(
        n7863), .ZN(n7865) );
  OAI21_X1 U9498 ( .B1(n9823), .B2(n7866), .A(n7865), .ZN(P1_U3254) );
  INV_X1 U9499 ( .A(n7867), .ZN(n7868) );
  NOR2_X1 U9500 ( .A1(n7871), .A2(n9361), .ZN(n9184) );
  NAND2_X1 U9501 ( .A1(n7872), .A2(n10389), .ZN(n7873) );
  AND3_X1 U9502 ( .A1(n10409), .A2(n7874), .A3(n7873), .ZN(n10388) );
  INV_X1 U9503 ( .A(n9373), .ZN(n9419) );
  AOI22_X1 U9504 ( .A1(n9184), .A2(n10388), .B1(P2_REG3_REG_2__SCAN_IN), .B2(
        n9419), .ZN(n7882) );
  OAI21_X1 U9505 ( .B1(n7877), .B2(n7876), .A(n7875), .ZN(n7878) );
  NAND2_X1 U9506 ( .A1(n7878), .A2(n4402), .ZN(n7880) );
  AOI22_X1 U9507 ( .A1(n9412), .A2(n7346), .B1(n9411), .B2(n7141), .ZN(n7879)
         );
  NAND2_X1 U9508 ( .A1(n7880), .A2(n7879), .ZN(n10387) );
  NAND2_X1 U9509 ( .A1(n9427), .A2(n10387), .ZN(n7881) );
  OAI211_X1 U9510 ( .C1(n7163), .C2(n9427), .A(n7882), .B(n7881), .ZN(n7890)
         );
  INV_X1 U9511 ( .A(n7884), .ZN(n7885) );
  NAND2_X1 U9512 ( .A1(n7885), .A2(n9361), .ZN(n7972) );
  NAND2_X1 U9513 ( .A1(n8560), .A2(n7972), .ZN(n7886) );
  XNOR2_X1 U9514 ( .A(n7887), .B(n5924), .ZN(n10391) );
  OAI22_X1 U9515 ( .A1(n7888), .A2(n9371), .B1(n9429), .B2(n10391), .ZN(n7889)
         );
  OR2_X1 U9516 ( .A1(n7890), .A2(n7889), .ZN(P2_U3294) );
  INV_X1 U9517 ( .A(n7891), .ZN(n8863) );
  OAI222_X1 U9518 ( .A1(n10251), .A2(n8379), .B1(n10244), .B2(n8863), .C1(
        P1_U3084), .C2(n7892), .ZN(P1_U3331) );
  XNOR2_X1 U9519 ( .A(n7893), .B(n7895), .ZN(n10200) );
  OAI22_X1 U9520 ( .A1(n8530), .A2(n9954), .B1(n7950), .B2(n9952), .ZN(n7898)
         );
  XOR2_X1 U9521 ( .A(n7894), .B(n7895), .Z(n7896) );
  NOR2_X1 U9522 ( .A1(n7896), .A2(n9950), .ZN(n7897) );
  AOI211_X1 U9523 ( .C1(n10200), .C2(n7946), .A(n7898), .B(n7897), .ZN(n10204)
         );
  INV_X1 U9524 ( .A(n10201), .ZN(n8535) );
  AOI21_X1 U9525 ( .B1(n10201), .B2(n7837), .A(n8039), .ZN(n10202) );
  NAND2_X1 U9526 ( .A1(n10202), .A2(n10052), .ZN(n7900) );
  AOI22_X1 U9527 ( .A1(n10317), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n8532), .B2(
        n10307), .ZN(n7899) );
  OAI211_X1 U9528 ( .C1(n8535), .C2(n10047), .A(n7900), .B(n7899), .ZN(n7901)
         );
  AOI21_X1 U9529 ( .B1(n7962), .B2(n10200), .A(n7901), .ZN(n7902) );
  OAI21_X1 U9530 ( .B1(n10204), .B2(n10317), .A(n7902), .ZN(P1_U3282) );
  AOI22_X1 U9531 ( .A1(n7904), .A2(n10341), .B1(n10207), .B2(n7903), .ZN(n7905) );
  OAI211_X1 U9532 ( .C1(n10188), .C2(n7907), .A(n7906), .B(n7905), .ZN(n7909)
         );
  NAND2_X1 U9533 ( .A1(n7909), .A2(n10357), .ZN(n7908) );
  OAI21_X1 U9534 ( .B1(n10357), .B2(n7003), .A(n7908), .ZN(P1_U3528) );
  INV_X1 U9535 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n7911) );
  NAND2_X1 U9536 ( .A1(n7909), .A2(n10353), .ZN(n7910) );
  OAI21_X1 U9537 ( .B1(n10353), .B2(n7911), .A(n7910), .ZN(P1_U3469) );
  INV_X1 U9538 ( .A(n7914), .ZN(n7916) );
  NAND2_X1 U9539 ( .A1(n7916), .A2(n7915), .ZN(n7917) );
  XNOR2_X1 U9540 ( .A(n7965), .B(n8820), .ZN(n7922) );
  INV_X1 U9541 ( .A(n7922), .ZN(n7920) );
  NOR2_X1 U9542 ( .A1(n7986), .A2(n8819), .ZN(n7921) );
  INV_X1 U9543 ( .A(n7921), .ZN(n7919) );
  NAND2_X1 U9544 ( .A1(n7920), .A2(n7919), .ZN(n8122) );
  INV_X1 U9545 ( .A(n8122), .ZN(n7923) );
  AND2_X1 U9546 ( .A1(n7922), .A2(n7921), .ZN(n8162) );
  NOR2_X1 U9547 ( .A1(n7923), .A2(n8162), .ZN(n7924) );
  XNOR2_X1 U9548 ( .A(n8168), .B(n7924), .ZN(n7930) );
  NOR2_X1 U9549 ( .A1(n9002), .A2(n8007), .ZN(n7928) );
  INV_X1 U9550 ( .A(n8159), .ZN(n9030) );
  NAND2_X1 U9551 ( .A1(n8990), .A2(n9030), .ZN(n7926) );
  OAI211_X1 U9552 ( .C1(n7936), .C2(n8992), .A(n7926), .B(n7925), .ZN(n7927)
         );
  AOI211_X1 U9553 ( .C1(n7965), .C2(n9019), .A(n7928), .B(n7927), .ZN(n7929)
         );
  OAI21_X1 U9554 ( .B1(n7930), .B2(n7677), .A(n7929), .ZN(P2_U3233) );
  INV_X1 U9555 ( .A(n7932), .ZN(n7933) );
  AOI21_X1 U9556 ( .B1(n7934), .B2(n7931), .A(n7933), .ZN(n10413) );
  XNOR2_X1 U9557 ( .A(n7935), .B(n7934), .ZN(n7937) );
  INV_X1 U9558 ( .A(n7936), .ZN(n9032) );
  AOI222_X1 U9559 ( .A1(n4402), .A2(n7937), .B1(n9032), .B2(n9412), .C1(n9034), 
        .C2(n9411), .ZN(n10412) );
  MUX2_X1 U9560 ( .A(n7938), .B(n10412), .S(n9427), .Z(n7944) );
  NAND2_X1 U9561 ( .A1(n9184), .A2(n10409), .ZN(n9425) );
  INV_X1 U9562 ( .A(n7997), .ZN(n7940) );
  AOI21_X1 U9563 ( .B1(n10407), .B2(n7939), .A(n7940), .ZN(n10410) );
  OAI22_X1 U9564 ( .A1(n9371), .A2(n5059), .B1(n9373), .B2(n7941), .ZN(n7942)
         );
  AOI21_X1 U9565 ( .B1(n9354), .B2(n10410), .A(n7942), .ZN(n7943) );
  OAI211_X1 U9566 ( .C1(n10413), .C2(n9429), .A(n7944), .B(n7943), .ZN(
        P2_U3289) );
  XNOR2_X1 U9567 ( .A(n7945), .B(n7948), .ZN(n10189) );
  NAND2_X1 U9568 ( .A1(n10189), .A2(n7946), .ZN(n7954) );
  XNOR2_X1 U9569 ( .A(n7947), .B(n7948), .ZN(n7952) );
  NAND2_X1 U9570 ( .A1(n10055), .A2(n9770), .ZN(n7949) );
  OAI21_X1 U9571 ( .B1(n9954), .B2(n7950), .A(n7949), .ZN(n7951) );
  AOI21_X1 U9572 ( .B1(n7952), .B2(n10099), .A(n7951), .ZN(n7953) );
  NAND2_X1 U9573 ( .A1(n7954), .A2(n7953), .ZN(n10194) );
  INV_X1 U9574 ( .A(n10194), .ZN(n7964) );
  OR2_X1 U9575 ( .A1(n7956), .A2(n10190), .ZN(n7957) );
  NAND2_X1 U9576 ( .A1(n7955), .A2(n7957), .ZN(n10191) );
  AOI22_X1 U9577 ( .A1(n10317), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n8545), .B2(
        n10307), .ZN(n7960) );
  NAND2_X1 U9578 ( .A1(n7958), .A2(n10064), .ZN(n7959) );
  OAI211_X1 U9579 ( .C1(n10191), .C2(n9936), .A(n7960), .B(n7959), .ZN(n7961)
         );
  AOI21_X1 U9580 ( .B1(n10189), .B2(n7962), .A(n7961), .ZN(n7963) );
  OAI21_X1 U9581 ( .B1(n7964), .B2(n10317), .A(n7963), .ZN(P1_U3280) );
  INV_X1 U9582 ( .A(n7986), .ZN(n9031) );
  OR2_X1 U9583 ( .A1(n7965), .A2(n9031), .ZN(n7966) );
  NAND2_X1 U9584 ( .A1(n7969), .A2(n7970), .ZN(n7971) );
  NAND2_X1 U9585 ( .A1(n8076), .A2(n7971), .ZN(n9551) );
  NOR2_X1 U9586 ( .A1(n9421), .A2(n7972), .ZN(n9402) );
  INV_X1 U9587 ( .A(n9402), .ZN(n8493) );
  OAI22_X1 U9588 ( .A1(n9384), .A2(n7986), .B1(n8657), .B2(n9386), .ZN(n7973)
         );
  INV_X1 U9589 ( .A(n7973), .ZN(n7978) );
  NAND2_X1 U9590 ( .A1(n7974), .A2(n7968), .ZN(n7975) );
  NAND3_X1 U9591 ( .A1(n7976), .A2(n4402), .A3(n7975), .ZN(n7977) );
  OAI211_X1 U9592 ( .C1(n9551), .C2(n8560), .A(n7978), .B(n7977), .ZN(n9546)
         );
  MUX2_X1 U9593 ( .A(n9546), .B(P2_REG2_REG_10__SCAN_IN), .S(n9404), .Z(n7979)
         );
  INV_X1 U9594 ( .A(n7979), .ZN(n7984) );
  INV_X1 U9595 ( .A(n9547), .ZN(n8131) );
  OR2_X1 U9596 ( .A1(n7980), .A2(n8131), .ZN(n7981) );
  AND2_X1 U9597 ( .A1(n8188), .A2(n7981), .ZN(n9548) );
  OAI22_X1 U9598 ( .A1(n9371), .A2(n8131), .B1(n9373), .B2(n8126), .ZN(n7982)
         );
  AOI21_X1 U9599 ( .B1(n9548), .B2(n9354), .A(n7982), .ZN(n7983) );
  OAI211_X1 U9600 ( .C1(n9551), .C2(n8493), .A(n7984), .B(n7983), .ZN(P2_U3286) );
  XNOR2_X1 U9601 ( .A(n7985), .B(n7988), .ZN(n7994) );
  INV_X1 U9602 ( .A(n7994), .ZN(n9557) );
  OAI22_X1 U9603 ( .A1(n9384), .A2(n7987), .B1(n7986), .B2(n9386), .ZN(n7993)
         );
  NAND2_X1 U9604 ( .A1(n7989), .A2(n7988), .ZN(n7990) );
  AOI21_X1 U9605 ( .B1(n7991), .B2(n7990), .A(n9406), .ZN(n7992) );
  AOI211_X1 U9606 ( .C1(n9394), .C2(n7994), .A(n7993), .B(n7992), .ZN(n9555)
         );
  MUX2_X1 U9607 ( .A(n7995), .B(n9555), .S(n9427), .Z(n8002) );
  AOI21_X1 U9608 ( .B1(n9552), .B2(n7997), .A(n7996), .ZN(n9553) );
  OAI22_X1 U9609 ( .A1(n9371), .A2(n7999), .B1(n9373), .B2(n7998), .ZN(n8000)
         );
  AOI21_X1 U9610 ( .B1(n9354), .B2(n9553), .A(n8000), .ZN(n8001) );
  OAI211_X1 U9611 ( .C1(n9557), .C2(n8493), .A(n8002), .B(n8001), .ZN(P2_U3288) );
  INV_X1 U9612 ( .A(n8003), .ZN(n8013) );
  MUX2_X1 U9613 ( .A(n8005), .B(n8004), .S(n9427), .Z(n8012) );
  INV_X1 U9614 ( .A(n8006), .ZN(n8010) );
  OAI22_X1 U9615 ( .A1(n9371), .A2(n8008), .B1(n8007), .B2(n9373), .ZN(n8009)
         );
  AOI21_X1 U9616 ( .B1(n8010), .B2(n9354), .A(n8009), .ZN(n8011) );
  OAI211_X1 U9617 ( .C1(n8013), .C2(n8493), .A(n8012), .B(n8011), .ZN(P2_U3287) );
  NAND2_X1 U9618 ( .A1(n8018), .A2(n8014), .ZN(n8016) );
  OAI211_X1 U9619 ( .C1(n8017), .C2(n9586), .A(n8016), .B(n8015), .ZN(P2_U3335) );
  NAND2_X1 U9620 ( .A1(n8018), .A2(n10246), .ZN(n8021) );
  INV_X1 U9621 ( .A(n8019), .ZN(n8020) );
  OAI211_X1 U9622 ( .C1(n8022), .C2(n10251), .A(n8021), .B(n8020), .ZN(
        P1_U3330) );
  INV_X1 U9623 ( .A(n8023), .ZN(n8030) );
  OAI21_X1 U9624 ( .B1(n9373), .B2(n8025), .A(n8024), .ZN(n8027) );
  NOR2_X1 U9625 ( .A1(n9427), .A2(n5166), .ZN(n8026) );
  AOI21_X1 U9626 ( .B1(n9427), .B2(n8027), .A(n8026), .ZN(n8029) );
  OAI21_X1 U9627 ( .B1(n9354), .B2(n9422), .A(n5070), .ZN(n8028) );
  OAI211_X1 U9628 ( .C1(n8030), .C2(n9429), .A(n8029), .B(n8028), .ZN(P2_U3296) );
  NAND2_X1 U9629 ( .A1(n8032), .A2(n8031), .ZN(n8033) );
  XNOR2_X1 U9630 ( .A(n8033), .B(n8035), .ZN(n8038) );
  XNOR2_X1 U9631 ( .A(n8034), .B(n8035), .ZN(n10199) );
  AOI22_X1 U9632 ( .A1(n10055), .A2(n9771), .B1(n10057), .B2(n9773), .ZN(n8036) );
  OAI21_X1 U9633 ( .B1(n10199), .B2(n10040), .A(n8036), .ZN(n8037) );
  AOI21_X1 U9634 ( .B1(n8038), .B2(n10099), .A(n8037), .ZN(n10198) );
  INV_X1 U9635 ( .A(n8039), .ZN(n8040) );
  AOI211_X1 U9636 ( .C1(n10196), .C2(n8040), .A(n10334), .B(n7956), .ZN(n10195) );
  AOI22_X1 U9637 ( .A1(n10317), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n8041), .B2(
        n10307), .ZN(n8042) );
  OAI21_X1 U9638 ( .B1(n8043), .B2(n10047), .A(n8042), .ZN(n8045) );
  NOR2_X1 U9639 ( .A1(n10199), .A2(n10049), .ZN(n8044) );
  AOI211_X1 U9640 ( .C1(n10195), .C2(n10077), .A(n8045), .B(n8044), .ZN(n8046)
         );
  OAI21_X1 U9641 ( .B1(n10317), .B2(n10198), .A(n8046), .ZN(P1_U3281) );
  NOR2_X1 U9642 ( .A1(n9427), .A2(n7164), .ZN(n8049) );
  INV_X1 U9643 ( .A(n9184), .ZN(n8515) );
  OAI22_X1 U9644 ( .A1(n8515), .A2(n8047), .B1(n7668), .B2(n9373), .ZN(n8048)
         );
  AOI211_X1 U9645 ( .C1(n9427), .C2(n8050), .A(n8049), .B(n8048), .ZN(n8053)
         );
  INV_X1 U9646 ( .A(n9429), .ZN(n9255) );
  AOI22_X1 U9647 ( .A1(n9255), .A2(n8051), .B1(n9422), .B2(n5189), .ZN(n8052)
         );
  NAND2_X1 U9648 ( .A1(n8053), .A2(n8052), .ZN(P2_U3295) );
  INV_X1 U9649 ( .A(n8054), .ZN(n8055) );
  NOR2_X1 U9650 ( .A1(n8056), .A2(n8055), .ZN(n8057) );
  XNOR2_X1 U9651 ( .A(n8057), .B(n8065), .ZN(n10397) );
  INV_X1 U9652 ( .A(n10397), .ZN(n8074) );
  OAI21_X1 U9653 ( .B1(n8058), .B2(n10394), .A(n10409), .ZN(n8059) );
  OR2_X1 U9654 ( .A1(n8060), .A2(n8059), .ZN(n10393) );
  OAI22_X1 U9655 ( .A1(n8515), .A2(n10393), .B1(n8061), .B2(n9373), .ZN(n8062)
         );
  AOI21_X1 U9656 ( .B1(n9422), .B2(n8063), .A(n8062), .ZN(n8073) );
  NAND2_X1 U9657 ( .A1(n7525), .A2(n8064), .ZN(n8066) );
  XNOR2_X1 U9658 ( .A(n8066), .B(n8065), .ZN(n8067) );
  NAND2_X1 U9659 ( .A1(n8067), .A2(n4402), .ZN(n8069) );
  NAND2_X1 U9660 ( .A1(n8069), .A2(n8068), .ZN(n10396) );
  INV_X1 U9661 ( .A(n10396), .ZN(n8071) );
  MUX2_X1 U9662 ( .A(n8071), .B(n8070), .S(n9421), .Z(n8072) );
  OAI211_X1 U9663 ( .C1(n8074), .C2(n9429), .A(n8073), .B(n8072), .ZN(P2_U3292) );
  NAND2_X1 U9664 ( .A1(n9547), .A2(n9030), .ZN(n8075) );
  NAND2_X1 U9665 ( .A1(n8550), .A2(n8551), .ZN(n8177) );
  OAI21_X1 U9666 ( .B1(n8550), .B2(n8551), .A(n8177), .ZN(n9545) );
  XNOR2_X1 U9667 ( .A(n8077), .B(n8551), .ZN(n8078) );
  AOI222_X1 U9668 ( .A1(n4402), .A2(n8078), .B1(n8973), .B2(n9412), .C1(n9030), 
        .C2(n9411), .ZN(n9544) );
  MUX2_X1 U9669 ( .A(n8145), .B(n9544), .S(n9427), .Z(n8081) );
  XNOR2_X1 U9670 ( .A(n8188), .B(n5068), .ZN(n9542) );
  OAI22_X1 U9671 ( .A1(n5068), .A2(n9371), .B1(n8171), .B2(n9373), .ZN(n8079)
         );
  AOI21_X1 U9672 ( .B1(n9542), .B2(n9354), .A(n8079), .ZN(n8080) );
  OAI211_X1 U9673 ( .C1(n9429), .C2(n9545), .A(n8081), .B(n8080), .ZN(P2_U3285) );
  INV_X1 U9674 ( .A(n8082), .ZN(n8092) );
  NOR2_X1 U9675 ( .A1(n9421), .A2(n9361), .ZN(n9337) );
  INV_X1 U9676 ( .A(n8083), .ZN(n8084) );
  NAND2_X1 U9677 ( .A1(n9337), .A2(n8084), .ZN(n8085) );
  OAI21_X1 U9678 ( .B1(n9373), .B2(n8086), .A(n8085), .ZN(n8087) );
  AOI21_X1 U9679 ( .B1(n9422), .B2(n4809), .A(n8087), .ZN(n8091) );
  MUX2_X1 U9680 ( .A(n8089), .B(n8088), .S(n9421), .Z(n8090) );
  OAI211_X1 U9681 ( .C1(n8092), .C2(n9429), .A(n8091), .B(n8090), .ZN(P2_U3291) );
  XNOR2_X1 U9682 ( .A(n8093), .B(n8096), .ZN(n8094) );
  AOI222_X1 U9683 ( .A1(n10099), .A2(n8094), .B1(n9771), .B2(n10057), .C1(
        n10058), .C2(n10055), .ZN(n10186) );
  XNOR2_X1 U9684 ( .A(n8095), .B(n8096), .ZN(n10187) );
  INV_X1 U9685 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n8098) );
  INV_X1 U9686 ( .A(n8593), .ZN(n8097) );
  OAI22_X1 U9687 ( .A1(n10315), .A2(n8098), .B1(n8097), .B2(n9992), .ZN(n8099)
         );
  AOI21_X1 U9688 ( .B1(n10184), .B2(n10064), .A(n8099), .ZN(n8102) );
  AOI21_X1 U9689 ( .B1(n7955), .B2(n10184), .A(n10334), .ZN(n8100) );
  AND2_X1 U9690 ( .A1(n8100), .A2(n8604), .ZN(n10183) );
  NAND2_X1 U9691 ( .A1(n10183), .A2(n10077), .ZN(n8101) );
  OAI211_X1 U9692 ( .C1(n10187), .C2(n10074), .A(n8102), .B(n8101), .ZN(n8103)
         );
  INV_X1 U9693 ( .A(n8103), .ZN(n8104) );
  OAI21_X1 U9694 ( .B1(n10186), .B2(n10317), .A(n8104), .ZN(P1_U3279) );
  INV_X1 U9695 ( .A(n8105), .ZN(n8106) );
  NOR2_X1 U9696 ( .A1(n8107), .A2(n8106), .ZN(n8109) );
  XNOR2_X1 U9697 ( .A(n8109), .B(n8108), .ZN(n8117) );
  AOI21_X1 U9698 ( .B1(n9755), .B2(n9775), .A(n8110), .ZN(n8113) );
  NAND2_X1 U9699 ( .A1(n9763), .A2(n8111), .ZN(n8112) );
  OAI211_X1 U9700 ( .C1(n8114), .C2(n9758), .A(n8113), .B(n8112), .ZN(n8115)
         );
  AOI21_X1 U9701 ( .B1(n10206), .B2(n9734), .A(n8115), .ZN(n8116) );
  OAI21_X1 U9702 ( .B1(n8117), .B2(n9737), .A(n8116), .ZN(P1_U3219) );
  XNOR2_X1 U9703 ( .A(n9547), .B(n8820), .ZN(n8118) );
  NOR2_X1 U9704 ( .A1(n8159), .A2(n8819), .ZN(n8119) );
  NAND2_X1 U9705 ( .A1(n8118), .A2(n8119), .ZN(n8161) );
  INV_X1 U9706 ( .A(n8118), .ZN(n8160) );
  INV_X1 U9707 ( .A(n8119), .ZN(n8120) );
  NAND2_X1 U9708 ( .A1(n8160), .A2(n8120), .ZN(n8121) );
  AND2_X1 U9709 ( .A1(n8161), .A2(n8121), .ZN(n8125) );
  OR2_X1 U9710 ( .A1(n8168), .A2(n8162), .ZN(n8123) );
  AND2_X1 U9711 ( .A1(n8123), .A2(n8122), .ZN(n8124) );
  AND2_X1 U9712 ( .A1(n8125), .A2(n8122), .ZN(n8163) );
  NAND2_X1 U9713 ( .A1(n8123), .A2(n8163), .ZN(n8158) );
  OAI211_X1 U9714 ( .C1(n8125), .C2(n8124), .A(n8158), .B(n9011), .ZN(n8130)
         );
  OAI22_X1 U9715 ( .A1(n9017), .A2(n8657), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8247), .ZN(n8128) );
  NOR2_X1 U9716 ( .A1(n9002), .A2(n8126), .ZN(n8127) );
  AOI211_X1 U9717 ( .C1(n9013), .C2(n9031), .A(n8128), .B(n8127), .ZN(n8129)
         );
  OAI211_X1 U9718 ( .C1(n8131), .C2(n8996), .A(n8130), .B(n8129), .ZN(P2_U3219) );
  INV_X1 U9719 ( .A(n8132), .ZN(n8136) );
  OAI222_X1 U9720 ( .A1(n10251), .A2(n8134), .B1(n10244), .B2(n8136), .C1(
        n8133), .C2(P1_U3084), .ZN(P1_U3329) );
  OAI222_X1 U9721 ( .A1(n8137), .A2(P2_U3152), .B1(n9591), .B2(n8136), .C1(
        n8135), .C2(n9586), .ZN(P2_U3334) );
  XNOR2_X1 U9722 ( .A(n9048), .B(P2_REG1_REG_11__SCAN_IN), .ZN(n9039) );
  XNOR2_X1 U9723 ( .A(n8649), .B(n8139), .ZN(n8140) );
  OAI21_X1 U9724 ( .B1(n8141), .B2(n8140), .A(n8648), .ZN(n8153) );
  NAND2_X1 U9725 ( .A1(n8142), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n8143) );
  NAND2_X1 U9726 ( .A1(n8144), .A2(n8143), .ZN(n9045) );
  MUX2_X1 U9727 ( .A(n8145), .B(P2_REG2_REG_11__SCAN_IN), .S(n9048), .Z(n9044)
         );
  NOR2_X1 U9728 ( .A1(n9045), .A2(n9044), .ZN(n9047) );
  MUX2_X1 U9729 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n8187), .S(n8649), .Z(n8147)
         );
  NAND2_X1 U9730 ( .A1(n8147), .A2(n8148), .ZN(n8643) );
  OAI211_X1 U9731 ( .C1(n8148), .C2(n8147), .A(n10361), .B(n8643), .ZN(n8151)
         );
  NOR2_X1 U9732 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8149), .ZN(n8664) );
  AOI21_X1 U9733 ( .B1(n10358), .B2(P2_ADDR_REG_12__SCAN_IN), .A(n8664), .ZN(
        n8150) );
  OAI211_X1 U9734 ( .C1(n9101), .C2(n8644), .A(n8151), .B(n8150), .ZN(n8152)
         );
  AOI21_X1 U9735 ( .B1(n8153), .B2(n10366), .A(n8152), .ZN(n8154) );
  INV_X1 U9736 ( .A(n8154), .ZN(P2_U3257) );
  XNOR2_X1 U9737 ( .A(n9541), .B(n8820), .ZN(n8731) );
  NOR2_X1 U9738 ( .A1(n8657), .A2(n8819), .ZN(n8730) );
  NAND2_X1 U9739 ( .A1(n8731), .A2(n8730), .ZN(n8725) );
  INV_X1 U9740 ( .A(n8731), .ZN(n8658) );
  INV_X1 U9741 ( .A(n8730), .ZN(n8155) );
  NAND2_X1 U9742 ( .A1(n8658), .A2(n8155), .ZN(n8156) );
  AND2_X1 U9743 ( .A1(n8725), .A2(n8156), .ZN(n8165) );
  INV_X1 U9744 ( .A(n8165), .ZN(n8157) );
  AOI21_X1 U9745 ( .B1(n8158), .B2(n8157), .A(n7677), .ZN(n8170) );
  NOR3_X1 U9746 ( .A1(n8984), .A2(n8160), .A3(n8159), .ZN(n8169) );
  INV_X1 U9747 ( .A(n8161), .ZN(n8164) );
  OR2_X1 U9748 ( .A1(n8162), .A2(n8164), .ZN(n8167) );
  OR2_X1 U9749 ( .A1(n8164), .A2(n8163), .ZN(n8166) );
  OAI21_X1 U9750 ( .B1(n8170), .B2(n8169), .A(n8662), .ZN(n8175) );
  OAI22_X1 U9751 ( .A1(n9017), .A2(n8661), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9042), .ZN(n8173) );
  NOR2_X1 U9752 ( .A1(n9002), .A2(n8171), .ZN(n8172) );
  AOI211_X1 U9753 ( .C1(n9013), .C2(n9030), .A(n8173), .B(n8172), .ZN(n8174)
         );
  OAI211_X1 U9754 ( .C1(n5068), .C2(n8996), .A(n8175), .B(n8174), .ZN(P2_U3238) );
  INV_X1 U9755 ( .A(n8657), .ZN(n9029) );
  NAND2_X1 U9756 ( .A1(n9541), .A2(n9029), .ZN(n8176) );
  AND2_X1 U9757 ( .A1(n8177), .A2(n8176), .ZN(n8180) );
  NAND2_X1 U9758 ( .A1(n8177), .A2(n8554), .ZN(n8178) );
  OAI21_X1 U9759 ( .B1(n8180), .B2(n8179), .A(n8178), .ZN(n8181) );
  INV_X1 U9760 ( .A(n8181), .ZN(n9540) );
  OAI211_X1 U9761 ( .C1(n8184), .C2(n8183), .A(n8182), .B(n4402), .ZN(n8186)
         );
  AOI22_X1 U9762 ( .A1(n9029), .A2(n9411), .B1(n9412), .B2(n9028), .ZN(n8185)
         );
  MUX2_X1 U9763 ( .A(n9539), .B(n8187), .S(n9421), .Z(n8191) );
  AOI21_X1 U9764 ( .B1(n9536), .B2(n5112), .A(n8564), .ZN(n9537) );
  OAI22_X1 U9765 ( .A1(n5067), .A2(n9371), .B1(n9373), .B2(n8663), .ZN(n8189)
         );
  AOI21_X1 U9766 ( .B1(n9537), .B2(n9354), .A(n8189), .ZN(n8190) );
  OAI211_X1 U9767 ( .C1(n9540), .C2(n9429), .A(n8191), .B(n8190), .ZN(P2_U3284) );
  INV_X1 U9768 ( .A(n8192), .ZN(n8197) );
  INV_X1 U9769 ( .A(n8193), .ZN(n8194) );
  OAI222_X1 U9770 ( .A1(n8866), .A2(n8195), .B1(n8864), .B2(n8197), .C1(n8194), 
        .C2(P2_U3152), .ZN(P2_U3332) );
  OAI222_X1 U9771 ( .A1(n10251), .A2(n8198), .B1(n10244), .B2(n8197), .C1(
        P1_U3084), .C2(n8196), .ZN(P1_U3327) );
  AOI21_X1 U9772 ( .B1(n8201), .B2(n8200), .A(n8199), .ZN(n8205) );
  XNOR2_X1 U9773 ( .A(n8203), .B(n8202), .ZN(n8204) );
  XNOR2_X1 U9774 ( .A(n8205), .B(n8204), .ZN(n8214) );
  OAI21_X1 U9775 ( .B1(n9758), .B2(n8207), .A(n8206), .ZN(n8208) );
  AOI21_X1 U9776 ( .B1(n9755), .B2(n8209), .A(n8208), .ZN(n8210) );
  OAI21_X1 U9777 ( .B1(n10345), .B2(n9760), .A(n8210), .ZN(n8211) );
  AOI21_X1 U9778 ( .B1(n8212), .B2(n9763), .A(n8211), .ZN(n8213) );
  OAI21_X1 U9779 ( .B1(n8214), .B2(n9765), .A(n8213), .ZN(n8490) );
  INV_X1 U9780 ( .A(keyinput15), .ZN(n8488) );
  INV_X1 U9781 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n10270) );
  OR4_X1 U9782 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .A3(n10256), .A4(n10270), .ZN(n8226) );
  NOR2_X1 U9783 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n10433) );
  INV_X1 U9784 ( .A(n10433), .ZN(n10285) );
  INV_X1 U9785 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n8445) );
  INV_X1 U9786 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8442) );
  AND4_X1 U9787 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P2_REG3_REG_7__SCAN_IN), .A3(
        n8445), .A4(n8442), .ZN(n8215) );
  INV_X1 U9788 ( .A(P1_WR_REG_SCAN_IN), .ZN(n8434) );
  NAND2_X1 U9789 ( .A1(n8215), .A2(n8434), .ZN(n8217) );
  INV_X1 U9790 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10340) );
  NAND4_X1 U9791 ( .A1(SI_23_), .A2(P2_D_REG_12__SCAN_IN), .A3(n10340), .A4(
        n8428), .ZN(n8216) );
  NOR2_X1 U9792 ( .A1(n8217), .A2(n8216), .ZN(n8223) );
  NOR2_X1 U9793 ( .A1(P1_ADDR_REG_14__SCAN_IN), .A2(P2_ADDR_REG_14__SCAN_IN), 
        .ZN(n10281) );
  INV_X1 U9794 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n8440) );
  NAND4_X1 U9795 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), 
        .A3(P2_ADDR_REG_10__SCAN_IN), .A4(n8440), .ZN(n8221) );
  NOR2_X1 U9796 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(P2_DATAO_REG_6__SCAN_IN), 
        .ZN(n8218) );
  NAND4_X1 U9797 ( .A1(n8219), .A2(P2_REG2_REG_3__SCAN_IN), .A3(n8218), .A4(
        n10359), .ZN(n8220) );
  NOR2_X1 U9798 ( .A1(n8221), .A2(n8220), .ZN(n8222) );
  NAND3_X1 U9799 ( .A1(n8223), .A2(n10281), .A3(n8222), .ZN(n8224) );
  NOR4_X1 U9800 ( .A1(n8226), .A2(n10285), .A3(n8225), .A4(n8224), .ZN(n8277)
         );
  INV_X1 U9801 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n8291) );
  NAND4_X1 U9802 ( .A1(P1_REG2_REG_14__SCAN_IN), .A2(P1_REG2_REG_10__SCAN_IN), 
        .A3(P2_REG1_REG_13__SCAN_IN), .A4(n8291), .ZN(n8234) );
  INV_X1 U9803 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n8228) );
  INV_X1 U9804 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n8227) );
  NAND4_X1 U9805 ( .A1(n8228), .A2(n8227), .A3(P2_REG1_REG_21__SCAN_IN), .A4(
        P2_D_REG_24__SCAN_IN), .ZN(n8233) );
  INV_X1 U9806 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n8229) );
  INV_X1 U9807 ( .A(P2_RD_REG_SCAN_IN), .ZN(n8302) );
  NAND4_X1 U9808 ( .A1(n8229), .A2(n7255), .A3(P1_D_REG_17__SCAN_IN), .A4(
        n8302), .ZN(n8232) );
  INV_X1 U9809 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n8230) );
  NAND4_X1 U9810 ( .A1(n8230), .A2(n8305), .A3(SI_26_), .A4(
        P2_REG3_REG_16__SCAN_IN), .ZN(n8231) );
  NOR4_X1 U9811 ( .A1(n8234), .A2(n8233), .A3(n8232), .A4(n8231), .ZN(n8276)
         );
  INV_X1 U9812 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n10374) );
  NAND4_X1 U9813 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), 
        .A3(P2_REG3_REG_1__SCAN_IN), .A4(n10374), .ZN(n8240) );
  NOR2_X1 U9814 ( .A1(P2_REG0_REG_29__SCAN_IN), .A2(P1_REG0_REG_30__SCAN_IN), 
        .ZN(n8237) );
  AND4_X1 U9815 ( .A1(SI_13_), .A2(P2_REG1_REG_29__SCAN_IN), .A3(
        P2_REG0_REG_8__SCAN_IN), .A4(P2_REG1_REG_10__SCAN_IN), .ZN(n8235) );
  NAND4_X1 U9816 ( .A1(n8237), .A2(n6334), .A3(n8236), .A4(n8235), .ZN(n8239)
         );
  INV_X1 U9817 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n8416) );
  NAND4_X1 U9818 ( .A1(P2_REG1_REG_26__SCAN_IN), .A2(P2_REG2_REG_6__SCAN_IN), 
        .A3(P2_D_REG_3__SCAN_IN), .A4(n8416), .ZN(n8238) );
  NOR3_X1 U9819 ( .A1(n8240), .A2(n8239), .A3(n8238), .ZN(n8275) );
  NAND4_X1 U9820 ( .A1(P1_DATAO_REG_7__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), 
        .A3(P2_REG3_REG_19__SCAN_IN), .A4(n9651), .ZN(n8244) );
  NAND4_X1 U9821 ( .A1(P1_D_REG_20__SCAN_IN), .A2(P2_DATAO_REG_22__SCAN_IN), 
        .A3(P1_REG1_REG_10__SCAN_IN), .A4(P2_STATE_REG_SCAN_IN), .ZN(n8243) );
  NAND4_X1 U9822 ( .A1(P1_D_REG_24__SCAN_IN), .A2(P1_REG3_REG_10__SCAN_IN), 
        .A3(P2_REG0_REG_1__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n8242) );
  NAND4_X1 U9823 ( .A1(P1_D_REG_30__SCAN_IN), .A2(P1_REG1_REG_20__SCAN_IN), 
        .A3(P2_IR_REG_12__SCAN_IN), .A4(n8414), .ZN(n8241) );
  NOR4_X1 U9824 ( .A1(n8244), .A2(n8243), .A3(n8242), .A4(n8241), .ZN(n8273)
         );
  NOR4_X1 U9825 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_DATAO_REG_12__SCAN_IN), 
        .A3(n6203), .A4(n9061), .ZN(n8272) );
  NAND4_X1 U9826 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(P1_REG3_REG_23__SCAN_IN), 
        .A3(P1_REG0_REG_6__SCAN_IN), .A4(P1_REG2_REG_5__SCAN_IN), .ZN(n8245)
         );
  NOR3_X1 U9827 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(n10419), .A3(n8245), .ZN(
        n8270) );
  INV_X1 U9828 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n8246) );
  NAND4_X1 U9829 ( .A1(n8247), .A2(n9587), .A3(n8246), .A4(
        P2_IR_REG_31__SCAN_IN), .ZN(n8251) );
  NAND4_X1 U9830 ( .A1(n8249), .A2(n8248), .A3(P2_REG0_REG_16__SCAN_IN), .A4(
        P2_REG1_REG_0__SCAN_IN), .ZN(n8250) );
  NOR2_X1 U9831 ( .A1(n8251), .A2(n8250), .ZN(n8269) );
  NAND4_X1 U9832 ( .A1(n8454), .A2(n8344), .A3(SI_5_), .A4(SI_9_), .ZN(n8260)
         );
  INV_X1 U9833 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n8258) );
  INV_X1 U9834 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n8316) );
  NAND3_X1 U9835 ( .A1(P1_REG1_REG_6__SCAN_IN), .A2(P1_REG2_REG_21__SCAN_IN), 
        .A3(n8316), .ZN(n8256) );
  INV_X1 U9836 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n8471) );
  AND4_X1 U9837 ( .A1(P1_REG0_REG_8__SCAN_IN), .A2(SI_12_), .A3(
        P1_REG0_REG_15__SCAN_IN), .A4(n8471), .ZN(n8254) );
  NOR4_X1 U9838 ( .A1(P1_REG3_REG_28__SCAN_IN), .A2(P1_REG3_REG_6__SCAN_IN), 
        .A3(P1_REG1_REG_9__SCAN_IN), .A4(n7836), .ZN(n8253) );
  NOR4_X1 U9839 ( .A1(P2_REG2_REG_25__SCAN_IN), .A2(n10242), .A3(n8340), .A4(
        n7218), .ZN(n8252) );
  NAND4_X1 U9840 ( .A1(n8254), .A2(n9846), .A3(n8253), .A4(n8252), .ZN(n8255)
         );
  NOR2_X1 U9841 ( .A1(n8256), .A2(n8255), .ZN(n8257) );
  NAND3_X1 U9842 ( .A1(n8258), .A2(P2_D_REG_22__SCAN_IN), .A3(n8257), .ZN(
        n8259) );
  NOR2_X1 U9843 ( .A1(n8260), .A2(n8259), .ZN(n8268) );
  INV_X1 U9844 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n8261) );
  INV_X1 U9845 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n8392) );
  NAND4_X1 U9846 ( .A1(n8262), .A2(n8261), .A3(n8392), .A4(
        P1_REG1_REG_2__SCAN_IN), .ZN(n8266) );
  NAND4_X1 U9847 ( .A1(n8264), .A2(n8263), .A3(n8343), .A4(
        P2_DATAO_REG_3__SCAN_IN), .ZN(n8265) );
  NOR2_X1 U9848 ( .A1(n8266), .A2(n8265), .ZN(n8267) );
  AND4_X1 U9849 ( .A1(n8270), .A2(n8269), .A3(n8268), .A4(n8267), .ZN(n8271)
         );
  AND3_X1 U9850 ( .A1(n8273), .A2(n8272), .A3(n8271), .ZN(n8274) );
  NAND4_X1 U9851 ( .A1(n8277), .A2(n8276), .A3(n8275), .A4(n8274), .ZN(n8487)
         );
  INV_X1 U9852 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n8279) );
  AOI22_X1 U9853 ( .A1(n8279), .A2(keyinput34), .B1(keyinput20), .B2(n10374), 
        .ZN(n8278) );
  OAI221_X1 U9854 ( .B1(n4503), .B2(keyinput34), .C1(n10374), .C2(keyinput20), 
        .A(n8278), .ZN(n8289) );
  AOI22_X1 U9855 ( .A1(n10256), .A2(keyinput37), .B1(n5171), .B2(keyinput118), 
        .ZN(n8280) );
  OAI221_X1 U9856 ( .B1(n10256), .B2(keyinput37), .C1(n5171), .C2(keyinput118), 
        .A(n8280), .ZN(n8288) );
  AOI22_X1 U9857 ( .A1(n8283), .A2(keyinput18), .B1(keyinput72), .B2(n8282), 
        .ZN(n8281) );
  OAI221_X1 U9858 ( .B1(n8283), .B2(keyinput18), .C1(n8282), .C2(keyinput72), 
        .A(n8281), .ZN(n8287) );
  XOR2_X1 U9859 ( .A(n6334), .B(keyinput82), .Z(n8285) );
  XNOR2_X1 U9860 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(keyinput16), .ZN(n8284) );
  NAND2_X1 U9861 ( .A1(n8285), .A2(n8284), .ZN(n8286) );
  NOR4_X1 U9862 ( .A1(n8289), .A2(n8288), .A3(n8287), .A4(n8286), .ZN(n8327)
         );
  AOI22_X1 U9863 ( .A1(n8647), .A2(keyinput104), .B1(n8291), .B2(keyinput94), 
        .ZN(n8290) );
  OAI221_X1 U9864 ( .B1(n8647), .B2(keyinput104), .C1(n8291), .C2(keyinput94), 
        .A(n8290), .ZN(n8294) );
  XOR2_X1 U9865 ( .A(P1_REG1_REG_1__SCAN_IN), .B(keyinput57), .Z(n8293) );
  XNOR2_X1 U9866 ( .A(n10431), .B(keyinput7), .ZN(n8292) );
  OR3_X1 U9867 ( .A1(n8294), .A2(n8293), .A3(n8292), .ZN(n8300) );
  AOI22_X1 U9868 ( .A1(n7255), .A2(keyinput40), .B1(n10321), .B2(keyinput83), 
        .ZN(n8295) );
  OAI221_X1 U9869 ( .B1(n7255), .B2(keyinput40), .C1(n10321), .C2(keyinput83), 
        .A(n8295), .ZN(n8299) );
  INV_X1 U9870 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n8634) );
  INV_X1 U9871 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n8297) );
  AOI22_X1 U9872 ( .A1(n8634), .A2(keyinput53), .B1(keyinput80), .B2(n8297), 
        .ZN(n8296) );
  OAI221_X1 U9873 ( .B1(n8634), .B2(keyinput53), .C1(n8297), .C2(keyinput80), 
        .A(n8296), .ZN(n8298) );
  NOR3_X1 U9874 ( .A1(n8300), .A2(n8299), .A3(n8298), .ZN(n8326) );
  INV_X1 U9875 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n10283) );
  AOI22_X1 U9876 ( .A1(n8302), .A2(keyinput47), .B1(keyinput71), .B2(n10283), 
        .ZN(n8301) );
  OAI221_X1 U9877 ( .B1(n8302), .B2(keyinput47), .C1(n10283), .C2(keyinput71), 
        .A(n8301), .ZN(n8312) );
  AOI22_X1 U9878 ( .A1(n8305), .A2(keyinput103), .B1(keyinput60), .B2(n8304), 
        .ZN(n8303) );
  OAI221_X1 U9879 ( .B1(n8305), .B2(keyinput103), .C1(n8304), .C2(keyinput60), 
        .A(n8303), .ZN(n8311) );
  INV_X1 U9880 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n10324) );
  XOR2_X1 U9881 ( .A(n10324), .B(keyinput32), .Z(n8309) );
  INV_X1 U9882 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n10375) );
  XOR2_X1 U9883 ( .A(n10375), .B(keyinput111), .Z(n8308) );
  XNOR2_X1 U9884 ( .A(P2_REG3_REG_4__SCAN_IN), .B(keyinput50), .ZN(n8307) );
  XNOR2_X1 U9885 ( .A(P1_IR_REG_0__SCAN_IN), .B(keyinput6), .ZN(n8306) );
  NAND4_X1 U9886 ( .A1(n8309), .A2(n8308), .A3(n8307), .A4(n8306), .ZN(n8310)
         );
  NOR3_X1 U9887 ( .A1(n8312), .A2(n8311), .A3(n8310), .ZN(n8325) );
  AOI22_X1 U9888 ( .A1(n5403), .A2(keyinput97), .B1(keyinput63), .B2(n10419), 
        .ZN(n8313) );
  OAI221_X1 U9889 ( .B1(n5403), .B2(keyinput97), .C1(n10419), .C2(keyinput63), 
        .A(n8313), .ZN(n8323) );
  AOI22_X1 U9890 ( .A1(n8315), .A2(keyinput108), .B1(n10325), .B2(keyinput25), 
        .ZN(n8314) );
  OAI221_X1 U9891 ( .B1(n8315), .B2(keyinput108), .C1(n10325), .C2(keyinput25), 
        .A(n8314), .ZN(n8322) );
  XOR2_X1 U9892 ( .A(n8316), .B(keyinput109), .Z(n8320) );
  XNOR2_X1 U9893 ( .A(P2_REG1_REG_1__SCAN_IN), .B(keyinput74), .ZN(n8319) );
  XNOR2_X1 U9894 ( .A(P2_REG1_REG_21__SCAN_IN), .B(keyinput100), .ZN(n8318) );
  XNOR2_X1 U9895 ( .A(P2_REG3_REG_3__SCAN_IN), .B(keyinput13), .ZN(n8317) );
  NAND4_X1 U9896 ( .A1(n8320), .A2(n8319), .A3(n8318), .A4(n8317), .ZN(n8321)
         );
  NOR3_X1 U9897 ( .A1(n8323), .A2(n8322), .A3(n8321), .ZN(n8324) );
  NAND4_X1 U9898 ( .A1(n8327), .A2(n8326), .A3(n8325), .A4(n8324), .ZN(n8485)
         );
  INV_X1 U9899 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10352) );
  AOI22_X1 U9900 ( .A1(n8329), .A2(keyinput95), .B1(keyinput17), .B2(n10352), 
        .ZN(n8328) );
  OAI221_X1 U9901 ( .B1(n8329), .B2(keyinput95), .C1(n10352), .C2(keyinput17), 
        .A(n8328), .ZN(n8338) );
  AOI22_X1 U9902 ( .A1(n8331), .A2(keyinput110), .B1(keyinput88), .B2(n7010), 
        .ZN(n8330) );
  OAI221_X1 U9903 ( .B1(n8331), .B2(keyinput110), .C1(n7010), .C2(keyinput88), 
        .A(n8330), .ZN(n8337) );
  AOI22_X1 U9904 ( .A1(n8261), .A2(keyinput119), .B1(n10326), .B2(keyinput81), 
        .ZN(n8332) );
  OAI221_X1 U9905 ( .B1(n8261), .B2(keyinput119), .C1(n10326), .C2(keyinput81), 
        .A(n8332), .ZN(n8336) );
  XNOR2_X1 U9906 ( .A(SI_5_), .B(keyinput68), .ZN(n8334) );
  XNOR2_X1 U9907 ( .A(keyinput10), .B(P1_REG2_REG_21__SCAN_IN), .ZN(n8333) );
  NAND2_X1 U9908 ( .A1(n8334), .A2(n8333), .ZN(n8335) );
  NOR4_X1 U9909 ( .A1(n8338), .A2(n8337), .A3(n8336), .A4(n8335), .ZN(n8372)
         );
  AOI22_X1 U9910 ( .A1(n8340), .A2(keyinput55), .B1(keyinput122), .B2(n5627), 
        .ZN(n8339) );
  OAI221_X1 U9911 ( .B1(n8340), .B2(keyinput55), .C1(n5627), .C2(keyinput122), 
        .A(n8339), .ZN(n8350) );
  INV_X1 U9912 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n10444) );
  AOI22_X1 U9913 ( .A1(n10444), .A2(keyinput35), .B1(n8249), .B2(keyinput8), 
        .ZN(n8341) );
  OAI221_X1 U9914 ( .B1(n10444), .B2(keyinput35), .C1(n8249), .C2(keyinput8), 
        .A(n8341), .ZN(n8349) );
  AOI22_X1 U9915 ( .A1(n8344), .A2(keyinput79), .B1(keyinput106), .B2(n8343), 
        .ZN(n8342) );
  OAI221_X1 U9916 ( .B1(n8344), .B2(keyinput79), .C1(n8343), .C2(keyinput106), 
        .A(n8342), .ZN(n8348) );
  INV_X1 U9917 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n10376) );
  XOR2_X1 U9918 ( .A(n10376), .B(keyinput91), .Z(n8346) );
  XNOR2_X1 U9919 ( .A(P2_IR_REG_31__SCAN_IN), .B(keyinput117), .ZN(n8345) );
  NAND2_X1 U9920 ( .A1(n8346), .A2(n8345), .ZN(n8347) );
  NOR4_X1 U9921 ( .A1(n8350), .A2(n8349), .A3(n8348), .A4(n8347), .ZN(n8371)
         );
  AOI22_X1 U9922 ( .A1(n10242), .A2(keyinput84), .B1(keyinput52), .B2(n7218), 
        .ZN(n8351) );
  OAI221_X1 U9923 ( .B1(n10242), .B2(keyinput84), .C1(n7218), .C2(keyinput52), 
        .A(n8351), .ZN(n8359) );
  AOI22_X1 U9924 ( .A1(n6203), .A2(keyinput49), .B1(keyinput102), .B2(n5209), 
        .ZN(n8352) );
  OAI221_X1 U9925 ( .B1(n6203), .B2(keyinput49), .C1(n5209), .C2(keyinput102), 
        .A(n8352), .ZN(n8358) );
  XNOR2_X1 U9926 ( .A(P2_REG3_REG_2__SCAN_IN), .B(keyinput93), .ZN(n8356) );
  XNOR2_X1 U9927 ( .A(P2_REG1_REG_0__SCAN_IN), .B(keyinput124), .ZN(n8355) );
  XNOR2_X1 U9928 ( .A(P1_REG3_REG_13__SCAN_IN), .B(keyinput107), .ZN(n8354) );
  XNOR2_X1 U9929 ( .A(SI_9_), .B(keyinput75), .ZN(n8353) );
  NAND4_X1 U9930 ( .A1(n8356), .A2(n8355), .A3(n8354), .A4(n8353), .ZN(n8357)
         );
  NOR3_X1 U9931 ( .A1(n8359), .A2(n8358), .A3(n8357), .ZN(n8370) );
  INV_X1 U9932 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n10255) );
  AOI22_X1 U9933 ( .A1(n9061), .A2(keyinput56), .B1(keyinput96), .B2(n10255), 
        .ZN(n8360) );
  OAI221_X1 U9934 ( .B1(n9061), .B2(keyinput56), .C1(n10255), .C2(keyinput96), 
        .A(n8360), .ZN(n8368) );
  AOI22_X1 U9935 ( .A1(n5362), .A2(keyinput105), .B1(keyinput9), .B2(n8362), 
        .ZN(n8361) );
  OAI221_X1 U9936 ( .B1(n5362), .B2(keyinput105), .C1(n8362), .C2(keyinput9), 
        .A(n8361), .ZN(n8367) );
  AOI22_X1 U9937 ( .A1(n6092), .A2(keyinput76), .B1(keyinput24), .B2(n7836), 
        .ZN(n8363) );
  OAI221_X1 U9938 ( .B1(n6092), .B2(keyinput76), .C1(n7836), .C2(keyinput24), 
        .A(n8363), .ZN(n8366) );
  AOI22_X1 U9939 ( .A1(n4521), .A2(keyinput73), .B1(n8520), .B2(keyinput120), 
        .ZN(n8364) );
  OAI221_X1 U9940 ( .B1(n4521), .B2(keyinput73), .C1(n8520), .C2(keyinput120), 
        .A(n8364), .ZN(n8365) );
  NOR4_X1 U9941 ( .A1(n8368), .A2(n8367), .A3(n8366), .A4(n8365), .ZN(n8369)
         );
  NAND4_X1 U9942 ( .A1(n8372), .A2(n8371), .A3(n8370), .A4(n8369), .ZN(n8484)
         );
  AOI22_X1 U9943 ( .A1(n5541), .A2(keyinput30), .B1(n9651), .B2(keyinput114), 
        .ZN(n8373) );
  OAI221_X1 U9944 ( .B1(n5541), .B2(keyinput30), .C1(n9651), .C2(keyinput114), 
        .A(n8373), .ZN(n8374) );
  INV_X1 U9945 ( .A(n8374), .ZN(n8386) );
  XNOR2_X1 U9946 ( .A(P2_IR_REG_12__SCAN_IN), .B(keyinput46), .ZN(n8377) );
  XNOR2_X1 U9947 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(keyinput121), .ZN(n8376) );
  XNOR2_X1 U9948 ( .A(keyinput90), .B(P1_IR_REG_15__SCAN_IN), .ZN(n8375) );
  AND3_X1 U9949 ( .A1(n8377), .A2(n8376), .A3(n8375), .ZN(n8385) );
  AOI22_X1 U9950 ( .A1(n8380), .A2(keyinput29), .B1(n8379), .B2(keyinput12), 
        .ZN(n8378) );
  OAI221_X1 U9951 ( .B1(n8380), .B2(keyinput29), .C1(n8379), .C2(keyinput12), 
        .A(n8378), .ZN(n8381) );
  INV_X1 U9952 ( .A(n8381), .ZN(n8384) );
  INV_X1 U9953 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n10318) );
  INV_X1 U9954 ( .A(keyinput42), .ZN(n8382) );
  XNOR2_X1 U9955 ( .A(n10318), .B(n8382), .ZN(n8383) );
  AND4_X1 U9956 ( .A1(n8386), .A2(n8385), .A3(n8384), .A4(n8383), .ZN(n8426)
         );
  INV_X1 U9957 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n10443) );
  AOI22_X1 U9958 ( .A1(n10443), .A2(keyinput39), .B1(P2_U3152), .B2(keyinput11), .ZN(n8387) );
  OAI221_X1 U9959 ( .B1(n10443), .B2(keyinput39), .C1(P2_U3152), .C2(
        keyinput11), .A(n8387), .ZN(n8390) );
  INV_X1 U9960 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n10322) );
  XNOR2_X1 U9961 ( .A(n10322), .B(keyinput38), .ZN(n8389) );
  XOR2_X1 U9962 ( .A(P1_REG1_REG_2__SCAN_IN), .B(keyinput87), .Z(n8388) );
  OR3_X1 U9963 ( .A1(n8390), .A2(n8389), .A3(n8388), .ZN(n8396) );
  AOI22_X1 U9964 ( .A1(n8392), .A2(keyinput64), .B1(keyinput67), .B2(n7005), 
        .ZN(n8391) );
  OAI221_X1 U9965 ( .B1(n8392), .B2(keyinput64), .C1(n7005), .C2(keyinput67), 
        .A(n8391), .ZN(n8395) );
  INV_X1 U9966 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n10254) );
  AOI22_X1 U9967 ( .A1(n10270), .A2(keyinput36), .B1(keyinput19), .B2(n10254), 
        .ZN(n8393) );
  OAI221_X1 U9968 ( .B1(n10270), .B2(keyinput36), .C1(n10254), .C2(keyinput19), 
        .A(n8393), .ZN(n8394) );
  NOR3_X1 U9969 ( .A1(n8396), .A2(n8395), .A3(n8394), .ZN(n8425) );
  AOI22_X1 U9970 ( .A1(n8399), .A2(keyinput61), .B1(keyinput92), .B2(n8398), 
        .ZN(n8397) );
  OAI221_X1 U9971 ( .B1(n8399), .B2(keyinput61), .C1(n8398), .C2(keyinput92), 
        .A(n8397), .ZN(n8410) );
  AOI22_X1 U9972 ( .A1(n8401), .A2(keyinput62), .B1(keyinput28), .B2(n7232), 
        .ZN(n8400) );
  OAI221_X1 U9973 ( .B1(n8401), .B2(keyinput62), .C1(n7232), .C2(keyinput28), 
        .A(n8400), .ZN(n8409) );
  AOI22_X1 U9974 ( .A1(n8403), .A2(keyinput125), .B1(keyinput33), .B2(n7668), 
        .ZN(n8402) );
  OAI221_X1 U9975 ( .B1(n8403), .B2(keyinput125), .C1(n7668), .C2(keyinput33), 
        .A(n8402), .ZN(n8408) );
  INV_X1 U9976 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n8406) );
  AOI22_X1 U9977 ( .A1(n8406), .A2(keyinput5), .B1(n8405), .B2(keyinput70), 
        .ZN(n8404) );
  OAI221_X1 U9978 ( .B1(n8406), .B2(keyinput5), .C1(n8405), .C2(keyinput70), 
        .A(n8404), .ZN(n8407) );
  NOR4_X1 U9979 ( .A1(n8410), .A2(n8409), .A3(n8408), .A4(n8407), .ZN(n8424)
         );
  INV_X1 U9980 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n10320) );
  AOI22_X1 U9981 ( .A1(n10320), .A2(keyinput3), .B1(keyinput45), .B2(n5173), 
        .ZN(n8411) );
  OAI221_X1 U9982 ( .B1(n10320), .B2(keyinput3), .C1(n5173), .C2(keyinput45), 
        .A(n8411), .ZN(n8422) );
  AOI22_X1 U9983 ( .A1(n8414), .A2(keyinput59), .B1(keyinput112), .B2(n8413), 
        .ZN(n8412) );
  OAI221_X1 U9984 ( .B1(n8414), .B2(keyinput59), .C1(n8413), .C2(keyinput112), 
        .A(n8412), .ZN(n8421) );
  INV_X1 U9985 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n10379) );
  AOI22_X1 U9986 ( .A1(n8416), .A2(keyinput1), .B1(keyinput85), .B2(n10379), 
        .ZN(n8415) );
  OAI221_X1 U9987 ( .B1(n8416), .B2(keyinput1), .C1(n10379), .C2(keyinput85), 
        .A(n8415), .ZN(n8420) );
  INV_X1 U9988 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n10378) );
  AOI22_X1 U9989 ( .A1(n8418), .A2(keyinput41), .B1(keyinput126), .B2(n10378), 
        .ZN(n8417) );
  OAI221_X1 U9990 ( .B1(n8418), .B2(keyinput41), .C1(n10378), .C2(keyinput126), 
        .A(n8417), .ZN(n8419) );
  NOR4_X1 U9991 ( .A1(n8422), .A2(n8421), .A3(n8420), .A4(n8419), .ZN(n8423)
         );
  NAND4_X1 U9992 ( .A1(n8426), .A2(n8425), .A3(n8424), .A4(n8423), .ZN(n8483)
         );
  INV_X1 U9993 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n10377) );
  AOI22_X1 U9994 ( .A1(n8428), .A2(keyinput23), .B1(keyinput43), .B2(n10377), 
        .ZN(n8427) );
  OAI221_X1 U9995 ( .B1(n8428), .B2(keyinput23), .C1(n10377), .C2(keyinput43), 
        .A(n8427), .ZN(n8438) );
  AOI22_X1 U9996 ( .A1(n10340), .A2(keyinput44), .B1(n8430), .B2(keyinput127), 
        .ZN(n8429) );
  OAI221_X1 U9997 ( .B1(n10340), .B2(keyinput44), .C1(n8430), .C2(keyinput127), 
        .A(n8429), .ZN(n8437) );
  XNOR2_X1 U9998 ( .A(n10367), .B(keyinput69), .ZN(n8433) );
  XNOR2_X1 U9999 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(keyinput78), .ZN(n8432) );
  XNOR2_X1 U10000 ( .A(keyinput54), .B(P2_REG2_REG_3__SCAN_IN), .ZN(n8431) );
  NAND3_X1 U10001 ( .A1(n8433), .A2(n8432), .A3(n8431), .ZN(n8436) );
  XNOR2_X1 U10002 ( .A(n8434), .B(keyinput22), .ZN(n8435) );
  NOR4_X1 U10003 ( .A1(n8438), .A2(n8437), .A3(n8436), .A4(n8435), .ZN(n8481)
         );
  AOI22_X1 U10004 ( .A1(n10323), .A2(keyinput0), .B1(keyinput115), .B2(n8440), 
        .ZN(n8439) );
  OAI221_X1 U10005 ( .B1(n10323), .B2(keyinput0), .C1(n8440), .C2(keyinput115), 
        .A(n8439), .ZN(n8451) );
  INV_X1 U10006 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n10319) );
  AOI22_X1 U10007 ( .A1(n8442), .A2(keyinput98), .B1(n10319), .B2(keyinput116), 
        .ZN(n8441) );
  OAI221_X1 U10008 ( .B1(n8442), .B2(keyinput98), .C1(n10319), .C2(keyinput116), .A(n8441), .ZN(n8450) );
  AOI22_X1 U10009 ( .A1(n8445), .A2(keyinput89), .B1(keyinput113), .B2(n8444), 
        .ZN(n8443) );
  OAI221_X1 U10010 ( .B1(n8445), .B2(keyinput89), .C1(n8444), .C2(keyinput113), 
        .A(n8443), .ZN(n8449) );
  INV_X1 U10011 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n8447) );
  XNOR2_X1 U10012 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput65), .ZN(n8446) );
  OAI21_X1 U10013 ( .B1(n8447), .B2(keyinput15), .A(n8446), .ZN(n8448) );
  NOR4_X1 U10014 ( .A1(n8451), .A2(n8450), .A3(n8449), .A4(n8448), .ZN(n8480)
         );
  INV_X1 U10015 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n8453) );
  AOI22_X1 U10016 ( .A1(n8454), .A2(keyinput99), .B1(keyinput51), .B2(n8453), 
        .ZN(n8452) );
  OAI221_X1 U10017 ( .B1(n8454), .B2(keyinput99), .C1(n8453), .C2(keyinput51), 
        .A(n8452), .ZN(n8464) );
  INV_X1 U10018 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n8457) );
  AOI22_X1 U10019 ( .A1(n8457), .A2(keyinput58), .B1(n8456), .B2(keyinput77), 
        .ZN(n8455) );
  OAI221_X1 U10020 ( .B1(n8457), .B2(keyinput58), .C1(n8456), .C2(keyinput77), 
        .A(n8455), .ZN(n8463) );
  XOR2_X1 U10021 ( .A(n9587), .B(keyinput101), .Z(n8461) );
  XOR2_X1 U10022 ( .A(n8262), .B(keyinput123), .Z(n8460) );
  XNOR2_X1 U10023 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(keyinput26), .ZN(n8459) );
  XNOR2_X1 U10024 ( .A(P1_REG3_REG_7__SCAN_IN), .B(keyinput48), .ZN(n8458) );
  NAND4_X1 U10025 ( .A1(n8461), .A2(n8460), .A3(n8459), .A4(n8458), .ZN(n8462)
         );
  NOR3_X1 U10026 ( .A1(n8464), .A2(n8463), .A3(n8462), .ZN(n8479) );
  AOI22_X1 U10027 ( .A1(n9846), .A2(keyinput66), .B1(keyinput27), .B2(n8466), 
        .ZN(n8465) );
  OAI221_X1 U10028 ( .B1(n9846), .B2(keyinput66), .C1(n8466), .C2(keyinput27), 
        .A(n8465), .ZN(n8477) );
  INV_X1 U10029 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n8468) );
  INV_X1 U10030 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n10284) );
  AOI22_X1 U10031 ( .A1(n8468), .A2(keyinput2), .B1(keyinput21), .B2(n10284), 
        .ZN(n8467) );
  OAI221_X1 U10032 ( .B1(n8468), .B2(keyinput2), .C1(n10284), .C2(keyinput21), 
        .A(n8467), .ZN(n8476) );
  INV_X1 U10033 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n8470) );
  AOI22_X1 U10034 ( .A1(n8471), .A2(keyinput31), .B1(n8470), .B2(keyinput86), 
        .ZN(n8469) );
  OAI221_X1 U10035 ( .B1(n8471), .B2(keyinput31), .C1(n8470), .C2(keyinput86), 
        .A(n8469), .ZN(n8475) );
  XNOR2_X1 U10036 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput4), .ZN(n8473) );
  XNOR2_X1 U10037 ( .A(P2_REG3_REG_10__SCAN_IN), .B(keyinput14), .ZN(n8472) );
  NAND2_X1 U10038 ( .A1(n8473), .A2(n8472), .ZN(n8474) );
  NOR4_X1 U10039 ( .A1(n8477), .A2(n8476), .A3(n8475), .A4(n8474), .ZN(n8478)
         );
  NAND4_X1 U10040 ( .A1(n8481), .A2(n8480), .A3(n8479), .A4(n8478), .ZN(n8482)
         );
  NOR4_X1 U10041 ( .A1(n8485), .A2(n8484), .A3(n8483), .A4(n8482), .ZN(n8486)
         );
  OAI221_X1 U10042 ( .B1(n8488), .B2(P2_IR_REG_25__SCAN_IN), .C1(n8488), .C2(
        n8487), .A(n8486), .ZN(n8489) );
  XNOR2_X1 U10043 ( .A(n8490), .B(n8489), .ZN(P1_U3237) );
  OAI22_X1 U10044 ( .A1(n9427), .A2(n7224), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n9373), .ZN(n8495) );
  OAI22_X1 U10045 ( .A1(n8493), .A2(n8492), .B1(n8491), .B2(n9371), .ZN(n8494)
         );
  AOI211_X1 U10046 ( .C1(n9184), .C2(n8496), .A(n8495), .B(n8494), .ZN(n8497)
         );
  OAI21_X1 U10047 ( .B1(n8498), .B2(n9404), .A(n8497), .ZN(P2_U3293) );
  OAI21_X1 U10048 ( .B1(n8511), .B2(n8500), .A(n8499), .ZN(n8501) );
  NAND2_X1 U10049 ( .A1(n8501), .A2(n4402), .ZN(n8503) );
  NAND2_X1 U10050 ( .A1(n8503), .A2(n8502), .ZN(n10405) );
  MUX2_X1 U10051 ( .A(n10405), .B(P2_REG2_REG_6__SCAN_IN), .S(n9421), .Z(n8517) );
  OAI211_X1 U10052 ( .C1(n8504), .C2(n10404), .A(n10409), .B(n7939), .ZN(
        n10401) );
  AOI22_X1 U10053 ( .A1(n9422), .A2(n8506), .B1(n9419), .B2(n8505), .ZN(n8514)
         );
  OR2_X1 U10054 ( .A1(n7784), .A2(n7785), .ZN(n8508) );
  AND2_X1 U10055 ( .A1(n8508), .A2(n8507), .ZN(n8510) );
  NAND2_X1 U10056 ( .A1(n8510), .A2(n8509), .ZN(n10400) );
  INV_X1 U10057 ( .A(n8510), .ZN(n8512) );
  NAND2_X1 U10058 ( .A1(n8512), .A2(n8511), .ZN(n10398) );
  NAND3_X1 U10059 ( .A1(n10400), .A2(n9255), .A3(n10398), .ZN(n8513) );
  OAI211_X1 U10060 ( .C1(n8515), .C2(n10401), .A(n8514), .B(n8513), .ZN(n8516)
         );
  OR2_X1 U10061 ( .A1(n8517), .A2(n8516), .ZN(P2_U3290) );
  INV_X1 U10062 ( .A(n8518), .ZN(n8522) );
  OAI222_X1 U10063 ( .A1(n10251), .A2(n8520), .B1(n10244), .B2(n8522), .C1(
        P1_U3084), .C2(n8519), .ZN(P1_U3328) );
  OAI222_X1 U10064 ( .A1(n8866), .A2(n8523), .B1(n9591), .B2(n8522), .C1(n8521), .C2(P2_U3152), .ZN(P2_U3333) );
  NAND2_X1 U10065 ( .A1(n8524), .A2(n8525), .ZN(n8573) );
  OAI21_X1 U10066 ( .B1(n8525), .B2(n8524), .A(n8573), .ZN(n8527) );
  NAND2_X1 U10067 ( .A1(n8527), .A2(n8526), .ZN(n8534) );
  NAND2_X1 U10068 ( .A1(n9703), .A2(n9772), .ZN(n8529) );
  OAI211_X1 U10069 ( .C1(n8530), .C2(n9743), .A(n8529), .B(n8528), .ZN(n8531)
         );
  AOI21_X1 U10070 ( .B1(n8532), .B2(n9763), .A(n8531), .ZN(n8533) );
  OAI211_X1 U10071 ( .C1(n8535), .C2(n9760), .A(n8534), .B(n8533), .ZN(
        P1_U3229) );
  NAND2_X1 U10072 ( .A1(n8524), .A2(n8536), .ZN(n8538) );
  NAND2_X1 U10073 ( .A1(n8538), .A2(n8537), .ZN(n8539) );
  XOR2_X1 U10074 ( .A(n8540), .B(n8539), .Z(n8547) );
  NAND2_X1 U10075 ( .A1(n9755), .A2(n9772), .ZN(n8542) );
  OAI211_X1 U10076 ( .C1(n9706), .C2(n9758), .A(n8542), .B(n8541), .ZN(n8544)
         );
  NOR2_X1 U10077 ( .A1(n10190), .A2(n9760), .ZN(n8543) );
  AOI211_X1 U10078 ( .C1(n8545), .C2(n9763), .A(n8544), .B(n8543), .ZN(n8546)
         );
  OAI21_X1 U10079 ( .B1(n8547), .B2(n9765), .A(n8546), .ZN(P1_U3234) );
  OAI21_X1 U10080 ( .B1(n8557), .B2(n4510), .A(n8548), .ZN(n8563) );
  OAI22_X1 U10081 ( .A1(n9384), .A2(n8661), .B1(n9012), .B2(n9386), .ZN(n8562)
         );
  INV_X1 U10082 ( .A(n8550), .ZN(n8555) );
  NAND2_X1 U10083 ( .A1(n5067), .A2(n8661), .ZN(n8552) );
  INV_X1 U10084 ( .A(n8552), .ZN(n8553) );
  NAND2_X1 U10085 ( .A1(n8558), .A2(n8557), .ZN(n8559) );
  NAND2_X1 U10086 ( .A1(n8621), .A2(n8559), .ZN(n9535) );
  NOR2_X1 U10087 ( .A1(n9535), .A2(n8560), .ZN(n8561) );
  AOI211_X1 U10088 ( .C1(n4402), .C2(n8563), .A(n8562), .B(n8561), .ZN(n9534)
         );
  OR2_X1 U10089 ( .A1(n8723), .A2(n8564), .ZN(n8565) );
  AND2_X1 U10090 ( .A1(n8845), .A2(n8565), .ZN(n9532) );
  NOR2_X1 U10091 ( .A1(n9373), .A2(n8975), .ZN(n8566) );
  AOI21_X1 U10092 ( .B1(n9421), .B2(P2_REG2_REG_13__SCAN_IN), .A(n8566), .ZN(
        n8567) );
  OAI21_X1 U10093 ( .B1(n8723), .B2(n9371), .A(n8567), .ZN(n8568) );
  AOI21_X1 U10094 ( .B1(n9532), .B2(n9354), .A(n8568), .ZN(n8571) );
  INV_X1 U10095 ( .A(n9535), .ZN(n8569) );
  NAND2_X1 U10096 ( .A1(n8569), .A2(n9402), .ZN(n8570) );
  OAI211_X1 U10097 ( .C1(n9534), .C2(n9404), .A(n8571), .B(n8570), .ZN(
        P2_U3283) );
  NAND2_X1 U10098 ( .A1(n8573), .A2(n8572), .ZN(n8574) );
  XOR2_X1 U10099 ( .A(n8575), .B(n8574), .Z(n8582) );
  OAI21_X1 U10100 ( .B1(n9758), .B2(n8589), .A(n8576), .ZN(n8577) );
  AOI21_X1 U10101 ( .B1(n9755), .B2(n9773), .A(n8577), .ZN(n8578) );
  OAI21_X1 U10102 ( .B1(n9732), .B2(n8579), .A(n8578), .ZN(n8580) );
  AOI21_X1 U10103 ( .B1(n10196), .B2(n9734), .A(n8580), .ZN(n8581) );
  OAI21_X1 U10104 ( .B1(n8582), .B2(n9737), .A(n8581), .ZN(P1_U3215) );
  XNOR2_X1 U10105 ( .A(n8584), .B(n8583), .ZN(n8585) );
  XNOR2_X1 U10106 ( .A(n8586), .B(n8585), .ZN(n8595) );
  NAND2_X1 U10107 ( .A1(n9703), .A2(n10058), .ZN(n8588) );
  OAI211_X1 U10108 ( .C1(n8589), .C2(n9743), .A(n8588), .B(n8587), .ZN(n8592)
         );
  NOR2_X1 U10109 ( .A1(n8590), .A2(n9760), .ZN(n8591) );
  AOI211_X1 U10110 ( .C1(n8593), .C2(n9763), .A(n8592), .B(n8591), .ZN(n8594)
         );
  OAI21_X1 U10111 ( .B1(n8595), .B2(n9765), .A(n8594), .ZN(P1_U3222) );
  OR2_X1 U10112 ( .A1(n8093), .A2(n8596), .ZN(n8598) );
  NAND2_X1 U10113 ( .A1(n8598), .A2(n8597), .ZN(n8602) );
  AND2_X1 U10114 ( .A1(n8600), .A2(n8599), .ZN(n8601) );
  OAI21_X1 U10115 ( .B1(n8608), .B2(n8602), .A(n8601), .ZN(n8603) );
  AOI222_X1 U10116 ( .A1(n10099), .A2(n8603), .B1(n9770), .B2(n10057), .C1(
        n10037), .C2(n10055), .ZN(n10181) );
  AOI21_X1 U10117 ( .B1(n10178), .B2(n8604), .A(n10061), .ZN(n10179) );
  AOI22_X1 U10118 ( .A1(n10317), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n9710), 
        .B2(n10307), .ZN(n8605) );
  OAI21_X1 U10119 ( .B1(n9707), .B2(n10047), .A(n8605), .ZN(n8610) );
  NAND2_X1 U10120 ( .A1(n8607), .A2(n8606), .ZN(n10069) );
  XOR2_X1 U10121 ( .A(n8608), .B(n10069), .Z(n10182) );
  NOR2_X1 U10122 ( .A1(n10182), .A2(n10074), .ZN(n8609) );
  AOI211_X1 U10123 ( .C1(n10179), .C2(n10052), .A(n8610), .B(n8609), .ZN(n8611) );
  OAI21_X1 U10124 ( .B1(n10317), .B2(n10181), .A(n8611), .ZN(P1_U3278) );
  OAI211_X1 U10125 ( .C1(n4479), .C2(n8613), .A(n8612), .B(n4402), .ZN(n8615)
         );
  INV_X1 U10126 ( .A(n9385), .ZN(n9142) );
  AOI22_X1 U10127 ( .A1(n9142), .A2(n9412), .B1(n9411), .B2(n9028), .ZN(n8614)
         );
  XOR2_X1 U10128 ( .A(n9526), .B(n8845), .Z(n9527) );
  INV_X1 U10129 ( .A(n9526), .ZN(n8616) );
  NOR2_X1 U10130 ( .A1(n8616), .A2(n9371), .ZN(n8619) );
  OAI22_X1 U10131 ( .A1(n9427), .A2(n8617), .B1(n8885), .B2(n9373), .ZN(n8618)
         );
  AOI211_X1 U10132 ( .C1(n9527), .C2(n9354), .A(n8619), .B(n8618), .ZN(n8624)
         );
  NAND2_X1 U10133 ( .A1(n9531), .A2(n9028), .ZN(n8620) );
  OAI21_X1 U10134 ( .B1(n4490), .B2(n8622), .A(n9140), .ZN(n9525) );
  NAND2_X1 U10135 ( .A1(n9525), .A2(n9255), .ZN(n8623) );
  OAI211_X1 U10136 ( .C1(n9529), .C2(n9404), .A(n8624), .B(n8623), .ZN(
        P2_U3282) );
  INV_X1 U10137 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n8627) );
  AOI22_X1 U10138 ( .A1(n8709), .A2(P1_REG1_REG_14__SCAN_IN), .B1(n8627), .B2(
        n8695), .ZN(n8628) );
  NAND2_X1 U10139 ( .A1(n8628), .A2(n8629), .ZN(n8708) );
  OAI21_X1 U10140 ( .B1(n8629), .B2(n8628), .A(n8708), .ZN(n8638) );
  NOR2_X1 U10141 ( .A1(n8630), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9609) );
  AOI21_X1 U10142 ( .B1(n10294), .B2(n8709), .A(n9609), .ZN(n8631) );
  OAI21_X1 U10143 ( .B1(n10443), .B2(n8719), .A(n8631), .ZN(n8637) );
  AOI211_X1 U10144 ( .C1(n8635), .C2(n8634), .A(n8697), .B(n9830), .ZN(n8636)
         );
  AOI211_X1 U10145 ( .C1(n10302), .C2(n8638), .A(n8637), .B(n8636), .ZN(n8639)
         );
  INV_X1 U10146 ( .A(n8639), .ZN(P1_U3255) );
  INV_X1 U10147 ( .A(n8640), .ZN(n8674) );
  AOI21_X1 U10148 ( .B1(n10239), .B2(P2_DATAO_REG_27__SCAN_IN), .A(n8641), 
        .ZN(n8642) );
  OAI21_X1 U10149 ( .B1(n8674), .B2(n10244), .A(n8642), .ZN(P1_U3326) );
  OAI21_X1 U10150 ( .B1(n8644), .B2(n8187), .A(n8643), .ZN(n8646) );
  AOI22_X1 U10151 ( .A1(P2_REG2_REG_13__SCAN_IN), .A2(n8677), .B1(n8681), .B2(
        n5391), .ZN(n8645) );
  AOI21_X1 U10152 ( .B1(n8646), .B2(n8645), .A(n8676), .ZN(n8656) );
  AOI22_X1 U10153 ( .A1(P2_REG1_REG_13__SCAN_IN), .A2(n8681), .B1(n8677), .B2(
        n8647), .ZN(n8651) );
  OAI21_X1 U10154 ( .B1(n8651), .B2(n8650), .A(n8683), .ZN(n8654) );
  NAND2_X1 U10155 ( .A1(P2_U3152), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n8971) );
  NAND2_X1 U10156 ( .A1(n10358), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n8652) );
  OAI211_X1 U10157 ( .C1(n9101), .C2(n8677), .A(n8971), .B(n8652), .ZN(n8653)
         );
  AOI21_X1 U10158 ( .B1(n8654), .B2(n10366), .A(n8653), .ZN(n8655) );
  OAI21_X1 U10159 ( .B1(n8656), .B2(n9124), .A(n8655), .ZN(P2_U3258) );
  INV_X1 U10160 ( .A(n8662), .ZN(n8660) );
  NOR3_X1 U10161 ( .A1(n8658), .A2(n8657), .A3(n8984), .ZN(n8659) );
  AOI21_X1 U10162 ( .B1(n8660), .B2(n9011), .A(n8659), .ZN(n8673) );
  XNOR2_X1 U10163 ( .A(n9536), .B(n8787), .ZN(n8726) );
  OR2_X1 U10164 ( .A1(n8819), .A2(n8661), .ZN(n8724) );
  INV_X1 U10165 ( .A(n8724), .ZN(n8729) );
  XNOR2_X1 U10166 ( .A(n8726), .B(n8729), .ZN(n8672) );
  NAND3_X1 U10167 ( .A1(n8662), .A2(n8725), .A3(n8672), .ZN(n8876) );
  NOR2_X1 U10168 ( .A1(n8876), .A2(n7677), .ZN(n8670) );
  AND2_X1 U10169 ( .A1(n9536), .A2(n9019), .ZN(n8669) );
  NOR2_X1 U10170 ( .A1(n9002), .A2(n8663), .ZN(n8668) );
  NAND2_X1 U10171 ( .A1(n9013), .A2(n9029), .ZN(n8666) );
  INV_X1 U10172 ( .A(n8664), .ZN(n8665) );
  OAI211_X1 U10173 ( .C1(n8879), .C2(n9017), .A(n8666), .B(n8665), .ZN(n8667)
         );
  NOR4_X1 U10174 ( .A1(n8670), .A2(n8669), .A3(n8668), .A4(n8667), .ZN(n8671)
         );
  OAI21_X1 U10175 ( .B1(n8673), .B2(n8672), .A(n8671), .ZN(P2_U3226) );
  OAI222_X1 U10176 ( .A1(n8866), .A2(n8675), .B1(n9591), .B2(n8674), .C1(n8847), .C2(P2_U3152), .ZN(P2_U3331) );
  AOI21_X1 U10177 ( .B1(n5391), .B2(n8677), .A(n8676), .ZN(n8679) );
  AOI22_X1 U10178 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n9054), .B1(n9059), .B2(
        n8617), .ZN(n8678) );
  AOI21_X1 U10179 ( .B1(n8679), .B2(n8678), .A(n9053), .ZN(n8690) );
  AOI22_X1 U10180 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n9059), .B1(n9054), .B2(
        n8680), .ZN(n8685) );
  OAI21_X1 U10181 ( .B1(n8685), .B2(n8684), .A(n9058), .ZN(n8688) );
  NAND2_X1 U10182 ( .A1(P2_U3152), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n8882) );
  NAND2_X1 U10183 ( .A1(n10358), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n8686) );
  OAI211_X1 U10184 ( .C1(n9101), .C2(n9054), .A(n8882), .B(n8686), .ZN(n8687)
         );
  AOI21_X1 U10185 ( .B1(n8688), .B2(n10366), .A(n8687), .ZN(n8689) );
  OAI21_X1 U10186 ( .B1(n8690), .B2(n9124), .A(n8689), .ZN(P2_U3259) );
  NAND2_X1 U10187 ( .A1(n4575), .A2(P1_U4006), .ZN(n8691) );
  OAI21_X1 U10188 ( .B1(P1_U4006), .B2(n5171), .A(n8691), .ZN(P1_U3555) );
  INV_X1 U10189 ( .A(n8692), .ZN(n10243) );
  OAI222_X1 U10190 ( .A1(n8866), .A2(n8694), .B1(P2_U3152), .B2(n8693), .C1(
        n9591), .C2(n10243), .ZN(P2_U3329) );
  NOR2_X1 U10191 ( .A1(n8696), .A2(n8695), .ZN(n8698) );
  NOR2_X1 U10192 ( .A1(n8699), .A2(n9802), .ZN(n8700) );
  INV_X1 U10193 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9804) );
  XNOR2_X1 U10194 ( .A(n8699), .B(n9802), .ZN(n9805) );
  NAND2_X1 U10195 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n8713), .ZN(n8701) );
  OAI21_X1 U10196 ( .B1(n8713), .B2(P1_REG2_REG_16__SCAN_IN), .A(n8701), .ZN(
        n9810) );
  NAND2_X1 U10197 ( .A1(P1_REG2_REG_17__SCAN_IN), .A2(n9829), .ZN(n8702) );
  OAI21_X1 U10198 ( .B1(n9829), .B2(P1_REG2_REG_17__SCAN_IN), .A(n8702), .ZN(
        n9832) );
  OR2_X1 U10199 ( .A1(n10293), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n8704) );
  NAND2_X1 U10200 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n10293), .ZN(n8703) );
  NAND2_X1 U10201 ( .A1(n8704), .A2(n8703), .ZN(n10290) );
  INV_X1 U10202 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n8706) );
  AOI22_X1 U10203 ( .A1(P1_REG1_REG_18__SCAN_IN), .A2(n10293), .B1(n8707), 
        .B2(n8706), .ZN(n10300) );
  OAI21_X1 U10204 ( .B1(n8709), .B2(P1_REG1_REG_14__SCAN_IN), .A(n8708), .ZN(
        n8710) );
  NOR2_X1 U10205 ( .A1(n9802), .A2(n8710), .ZN(n8712) );
  INV_X1 U10206 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n8711) );
  NOR2_X1 U10207 ( .A1(n8711), .A2(n9796), .ZN(n9797) );
  XNOR2_X1 U10208 ( .A(n8713), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n9813) );
  XNOR2_X1 U10209 ( .A(n9829), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n9825) );
  NAND2_X1 U10210 ( .A1(n10300), .A2(n10299), .ZN(n10298) );
  AOI22_X1 U10211 ( .A1(n8716), .A2(n10292), .B1(n10302), .B2(n8714), .ZN(
        n8718) );
  INV_X1 U10212 ( .A(n8714), .ZN(n8717) );
  NAND2_X1 U10213 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9632) );
  AOI22_X1 U10214 ( .A1(n9013), .A2(n9313), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3152), .ZN(n8722) );
  NAND2_X1 U10215 ( .A1(n9014), .A2(n9268), .ZN(n8721) );
  OAI211_X1 U10216 ( .C1(n9281), .C2(n9017), .A(n8722), .B(n8721), .ZN(n8781)
         );
  XNOR2_X1 U10217 ( .A(n8723), .B(n8820), .ZN(n8880) );
  NAND2_X1 U10218 ( .A1(n8788), .A2(n9028), .ZN(n8735) );
  NAND2_X1 U10219 ( .A1(n8880), .A2(n8735), .ZN(n8878) );
  NAND2_X1 U10220 ( .A1(n8726), .A2(n8724), .ZN(n8875) );
  NAND2_X1 U10221 ( .A1(n8878), .A2(n8875), .ZN(n8741) );
  XNOR2_X1 U10222 ( .A(n9526), .B(n8787), .ZN(n8745) );
  NOR2_X1 U10223 ( .A1(n9012), .A2(n8819), .ZN(n8743) );
  XNOR2_X1 U10224 ( .A(n8745), .B(n8743), .ZN(n8889) );
  NAND2_X1 U10225 ( .A1(n8725), .A2(n8724), .ZN(n8728) );
  INV_X1 U10226 ( .A(n8726), .ZN(n8727) );
  NAND2_X1 U10227 ( .A1(n8728), .A2(n8727), .ZN(n8733) );
  NAND3_X1 U10228 ( .A1(n8731), .A2(n8730), .A3(n8729), .ZN(n8732) );
  NAND2_X1 U10229 ( .A1(n8733), .A2(n8732), .ZN(n8734) );
  NAND2_X1 U10230 ( .A1(n8878), .A2(n8734), .ZN(n8738) );
  INV_X1 U10231 ( .A(n8880), .ZN(n8737) );
  INV_X1 U10232 ( .A(n8735), .ZN(n8736) );
  NAND2_X1 U10233 ( .A1(n8737), .A2(n8736), .ZN(n8877) );
  AND2_X1 U10234 ( .A1(n8738), .A2(n8877), .ZN(n8739) );
  XNOR2_X1 U10235 ( .A(n9398), .B(n8787), .ZN(n8930) );
  OR2_X1 U10236 ( .A1(n9027), .A2(n8819), .ZN(n8929) );
  XNOR2_X1 U10237 ( .A(n9522), .B(n8820), .ZN(n8926) );
  NOR2_X1 U10238 ( .A1(n9385), .A2(n8819), .ZN(n8748) );
  INV_X1 U10239 ( .A(n8743), .ZN(n8744) );
  NAND2_X1 U10240 ( .A1(n8745), .A2(n8744), .ZN(n8922) );
  OAI21_X1 U10241 ( .B1(n8926), .B2(n8748), .A(n8922), .ZN(n8746) );
  AOI21_X1 U10242 ( .B1(n8930), .B2(n8929), .A(n8746), .ZN(n8747) );
  NAND2_X1 U10243 ( .A1(n8923), .A2(n8747), .ZN(n8753) );
  INV_X1 U10244 ( .A(n8930), .ZN(n8751) );
  INV_X1 U10245 ( .A(n8926), .ZN(n8924) );
  INV_X1 U10246 ( .A(n8748), .ZN(n9010) );
  OAI21_X1 U10247 ( .B1(n8924), .B2(n9010), .A(n8929), .ZN(n8750) );
  NOR2_X1 U10248 ( .A1(n8929), .A2(n9010), .ZN(n8749) );
  AOI22_X1 U10249 ( .A1(n8751), .A2(n8750), .B1(n8749), .B2(n8926), .ZN(n8752)
         );
  NAND2_X1 U10250 ( .A1(n8753), .A2(n8752), .ZN(n8941) );
  XNOR2_X1 U10251 ( .A(n9508), .B(n8820), .ZN(n8754) );
  NOR2_X1 U10252 ( .A1(n9387), .A2(n8819), .ZN(n8755) );
  NAND2_X1 U10253 ( .A1(n8754), .A2(n8755), .ZN(n8758) );
  INV_X1 U10254 ( .A(n8754), .ZN(n8985) );
  INV_X1 U10255 ( .A(n8755), .ZN(n8756) );
  NAND2_X1 U10256 ( .A1(n8985), .A2(n8756), .ZN(n8757) );
  AND2_X1 U10257 ( .A1(n8758), .A2(n8757), .ZN(n8942) );
  NAND2_X1 U10258 ( .A1(n8941), .A2(n8942), .ZN(n8940) );
  NAND2_X1 U10259 ( .A1(n8940), .A2(n8758), .ZN(n8763) );
  XNOR2_X1 U10260 ( .A(n9499), .B(n8820), .ZN(n8759) );
  NOR2_X1 U10261 ( .A1(n9147), .A2(n8819), .ZN(n8760) );
  NAND2_X1 U10262 ( .A1(n8759), .A2(n8760), .ZN(n8764) );
  INV_X1 U10263 ( .A(n8759), .ZN(n8901) );
  INV_X1 U10264 ( .A(n8760), .ZN(n8761) );
  NAND2_X1 U10265 ( .A1(n8901), .A2(n8761), .ZN(n8762) );
  AND2_X1 U10266 ( .A1(n8764), .A2(n8762), .ZN(n8982) );
  XNOR2_X1 U10267 ( .A(n9495), .B(n8787), .ZN(n8768) );
  NOR2_X1 U10268 ( .A1(n9349), .A2(n8819), .ZN(n8766) );
  XNOR2_X1 U10269 ( .A(n8768), .B(n8766), .ZN(n8902) );
  INV_X1 U10270 ( .A(n8766), .ZN(n8767) );
  NAND2_X1 U10271 ( .A1(n8768), .A2(n8767), .ZN(n8769) );
  XNOR2_X1 U10272 ( .A(n9489), .B(n8820), .ZN(n8770) );
  AND2_X1 U10273 ( .A1(n9332), .A2(n8788), .ZN(n8771) );
  NAND2_X1 U10274 ( .A1(n8770), .A2(n8771), .ZN(n8774) );
  INV_X1 U10275 ( .A(n8770), .ZN(n8913) );
  INV_X1 U10276 ( .A(n8771), .ZN(n8772) );
  NAND2_X1 U10277 ( .A1(n8913), .A2(n8772), .ZN(n8773) );
  NAND2_X1 U10278 ( .A1(n8774), .A2(n8773), .ZN(n8962) );
  XNOR2_X1 U10279 ( .A(n9290), .B(n8820), .ZN(n8776) );
  NOR2_X1 U10280 ( .A1(n9280), .A2(n8819), .ZN(n8777) );
  XNOR2_X1 U10281 ( .A(n8776), .B(n8777), .ZN(n8911) );
  NAND2_X1 U10282 ( .A1(n8775), .A2(n8911), .ZN(n8798) );
  INV_X1 U10283 ( .A(n8776), .ZN(n8778) );
  NAND2_X1 U10284 ( .A1(n8778), .A2(n8777), .ZN(n8795) );
  NAND2_X1 U10285 ( .A1(n8798), .A2(n8795), .ZN(n8779) );
  XNOR2_X1 U10286 ( .A(n5593), .B(n8820), .ZN(n8794) );
  INV_X1 U10287 ( .A(n8794), .ZN(n8800) );
  XNOR2_X1 U10288 ( .A(n8779), .B(n8800), .ZN(n8782) );
  NOR3_X1 U10289 ( .A1(n8782), .A2(n8916), .A3(n8984), .ZN(n8780) );
  AOI211_X1 U10290 ( .C1(n5593), .C2(n9019), .A(n8781), .B(n8780), .ZN(n8784)
         );
  NOR2_X1 U10291 ( .A1(n8916), .A2(n8819), .ZN(n8793) );
  INV_X1 U10292 ( .A(n8793), .ZN(n8799) );
  NAND3_X1 U10293 ( .A1(n8782), .A2(n9011), .A3(n8799), .ZN(n8783) );
  NAND2_X1 U10294 ( .A1(n8784), .A2(n8783), .ZN(P2_U3237) );
  OAI22_X1 U10295 ( .A1(n9197), .A2(n9386), .B1(n8954), .B2(n9384), .ZN(n9230)
         );
  INV_X1 U10296 ( .A(n8999), .ZN(n8785) );
  AOI22_X1 U10297 ( .A1(n9230), .A2(n8785), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3152), .ZN(n8786) );
  OAI21_X1 U10298 ( .B1(n9224), .B2(n9002), .A(n8786), .ZN(n8812) );
  XNOR2_X1 U10299 ( .A(n9464), .B(n8787), .ZN(n8792) );
  NAND2_X1 U10300 ( .A1(n9026), .A2(n8788), .ZN(n8789) );
  NOR2_X1 U10301 ( .A1(n8792), .A2(n8789), .ZN(n8814) );
  NAND2_X1 U10302 ( .A1(n8792), .A2(n8789), .ZN(n8813) );
  NAND2_X1 U10303 ( .A1(n9026), .A2(n8790), .ZN(n8791) );
  OAI22_X1 U10304 ( .A1(n8813), .A2(n7677), .B1(n8792), .B2(n8791), .ZN(n8810)
         );
  NAND2_X1 U10305 ( .A1(n8794), .A2(n8793), .ZN(n8796) );
  AND2_X1 U10306 ( .A1(n8796), .A2(n8795), .ZN(n8797) );
  NAND2_X1 U10307 ( .A1(n8800), .A2(n8799), .ZN(n8801) );
  XNOR2_X1 U10308 ( .A(n9475), .B(n8820), .ZN(n8805) );
  XNOR2_X2 U10309 ( .A(n8804), .B(n8805), .ZN(n8893) );
  XNOR2_X1 U10310 ( .A(n9468), .B(n8820), .ZN(n8952) );
  NOR2_X1 U10311 ( .A1(n9281), .A2(n8819), .ZN(n8892) );
  INV_X1 U10312 ( .A(n8802), .ZN(n8803) );
  NOR2_X1 U10313 ( .A1(n8954), .A2(n8819), .ZN(n8806) );
  OAI21_X1 U10314 ( .B1(n8806), .B2(n8952), .A(n8949), .ZN(n8808) );
  INV_X1 U10315 ( .A(n8806), .ZN(n8956) );
  XNOR2_X1 U10316 ( .A(n9461), .B(n8820), .ZN(n8815) );
  NOR2_X1 U10317 ( .A1(n9197), .A2(n8819), .ZN(n8816) );
  XNOR2_X1 U10318 ( .A(n8815), .B(n8816), .ZN(n8997) );
  NOR2_X1 U10319 ( .A1(n8825), .A2(n8819), .ZN(n8818) );
  XNOR2_X1 U10320 ( .A(n9454), .B(n8820), .ZN(n8817) );
  XOR2_X1 U10321 ( .A(n8818), .B(n8817), .Z(n8867) );
  NOR2_X1 U10322 ( .A1(n9198), .A2(n8819), .ZN(n8821) );
  XNOR2_X1 U10323 ( .A(n8821), .B(n8820), .ZN(n8822) );
  XNOR2_X1 U10324 ( .A(n9452), .B(n8822), .ZN(n8823) );
  XNOR2_X1 U10325 ( .A(n8824), .B(n8823), .ZN(n8831) );
  INV_X1 U10326 ( .A(n8825), .ZN(n9153) );
  INV_X1 U10327 ( .A(n8826), .ZN(n9024) );
  AOI22_X1 U10328 ( .A1(n9153), .A2(n9411), .B1(n9024), .B2(n9412), .ZN(n9181)
         );
  NOR2_X1 U10329 ( .A1(n9181), .A2(n8999), .ZN(n8829) );
  OAI22_X1 U10330 ( .A1(n9185), .A2(n9002), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8827), .ZN(n8828) );
  AOI211_X1 U10331 ( .C1(n9452), .C2(n9019), .A(n8829), .B(n8828), .ZN(n8830)
         );
  OAI21_X1 U10332 ( .B1(n8831), .B2(n7677), .A(n8830), .ZN(P2_U3222) );
  INV_X1 U10333 ( .A(n9864), .ZN(n8834) );
  INV_X1 U10334 ( .A(n9849), .ZN(n8833) );
  AOI211_X1 U10335 ( .C1(n10107), .C2(n8834), .A(n10334), .B(n8833), .ZN(
        n10106) );
  INV_X1 U10336 ( .A(n8835), .ZN(n9597) );
  AOI22_X1 U10337 ( .A1(n9597), .A2(n10307), .B1(P1_REG2_REG_27__SCAN_IN), 
        .B2(n10317), .ZN(n8836) );
  OAI21_X1 U10338 ( .B1(n8837), .B2(n10047), .A(n8836), .ZN(n8843) );
  INV_X1 U10339 ( .A(n9475), .ZN(n9261) );
  INV_X1 U10340 ( .A(n8846), .ZN(n9416) );
  INV_X1 U10341 ( .A(n9398), .ZN(n9512) );
  OR2_X2 U10342 ( .A1(n9341), .A2(n9495), .ZN(n9320) );
  NAND2_X1 U10343 ( .A1(n9305), .A2(n9290), .ZN(n9267) );
  INV_X1 U10344 ( .A(n9438), .ZN(n9171) );
  XOR2_X1 U10345 ( .A(n8844), .B(n9133), .Z(n9431) );
  NOR2_X1 U10346 ( .A1(n8847), .A2(n7120), .ZN(n8848) );
  OR2_X1 U10347 ( .A1(n9386), .A2(n8848), .ZN(n9161) );
  NOR2_X1 U10348 ( .A1(n9161), .A2(n8849), .ZN(n9434) );
  NAND2_X1 U10349 ( .A1(n9427), .A2(n9434), .ZN(n9134) );
  OAI21_X1 U10350 ( .B1(n9427), .B2(n8850), .A(n9134), .ZN(n8851) );
  AOI21_X1 U10351 ( .B1(n8844), .B2(n9422), .A(n8851), .ZN(n8852) );
  OAI21_X1 U10352 ( .B1(n9431), .B2(n9425), .A(n8852), .ZN(P2_U3265) );
  INV_X1 U10353 ( .A(n10247), .ZN(n8853) );
  OAI222_X1 U10354 ( .A1(n8866), .A2(n8855), .B1(P2_U3152), .B2(n8854), .C1(
        n9591), .C2(n8853), .ZN(P2_U3330) );
  INV_X1 U10355 ( .A(n8856), .ZN(n8860) );
  OAI222_X1 U10356 ( .A1(n9586), .A2(n8858), .B1(n9591), .B2(n8860), .C1(n8857), .C2(P2_U3152), .ZN(P2_U3328) );
  OAI222_X1 U10357 ( .A1(P1_U3084), .A2(n8861), .B1(n10244), .B2(n8860), .C1(
        n8859), .C2(n10251), .ZN(P1_U3323) );
  OAI222_X1 U10358 ( .A1(n8866), .A2(n8865), .B1(n8864), .B2(n8863), .C1(
        P2_U3152), .C2(n8862), .ZN(P2_U3336) );
  XNOR2_X1 U10359 ( .A(n8868), .B(n8867), .ZN(n8874) );
  OAI22_X1 U10360 ( .A1(n9197), .A2(n8992), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8869), .ZN(n8871) );
  NOR2_X1 U10361 ( .A1(n9198), .A2(n9017), .ZN(n8870) );
  AOI211_X1 U10362 ( .C1(n9014), .C2(n9193), .A(n8871), .B(n8870), .ZN(n8873)
         );
  NAND2_X1 U10363 ( .A1(n9454), .A2(n9019), .ZN(n8872) );
  OAI211_X1 U10364 ( .C1(n8874), .C2(n7677), .A(n8873), .B(n8872), .ZN(
        P2_U3216) );
  NAND2_X1 U10365 ( .A1(n8876), .A2(n8875), .ZN(n8977) );
  NAND2_X1 U10366 ( .A1(n8878), .A2(n8877), .ZN(n8978) );
  NOR2_X1 U10367 ( .A1(n8977), .A2(n8978), .ZN(n8976) );
  NOR3_X1 U10368 ( .A1(n8880), .A2(n8879), .A3(n8984), .ZN(n8881) );
  AOI21_X1 U10369 ( .B1(n8976), .B2(n9011), .A(n8881), .ZN(n8890) );
  OAI21_X1 U10370 ( .B1(n9017), .B2(n9385), .A(n8882), .ZN(n8883) );
  AOI21_X1 U10371 ( .B1(n9013), .B2(n9028), .A(n8883), .ZN(n8884) );
  OAI21_X1 U10372 ( .B1(n8885), .B2(n9002), .A(n8884), .ZN(n8887) );
  NOR2_X1 U10373 ( .A1(n8923), .A2(n7677), .ZN(n8886) );
  AOI211_X1 U10374 ( .C1(n9526), .C2(n9019), .A(n8887), .B(n8886), .ZN(n8888)
         );
  OAI21_X1 U10375 ( .B1(n8890), .B2(n8889), .A(n8888), .ZN(P2_U3217) );
  INV_X1 U10376 ( .A(n8893), .ZN(n8891) );
  OAI22_X1 U10377 ( .A1(n8891), .A2(n7677), .B1(n9281), .B2(n8984), .ZN(n8894)
         );
  NAND2_X1 U10378 ( .A1(n8894), .A2(n8951), .ZN(n8899) );
  INV_X1 U10379 ( .A(n8895), .ZN(n9259) );
  AOI22_X1 U10380 ( .A1(n9251), .A2(n8990), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3152), .ZN(n8896) );
  OAI21_X1 U10381 ( .B1(n8916), .B2(n8992), .A(n8896), .ZN(n8897) );
  AOI21_X1 U10382 ( .B1(n9259), .B2(n9014), .A(n8897), .ZN(n8898) );
  OAI211_X1 U10383 ( .C1(n9261), .C2(n8996), .A(n8899), .B(n8898), .ZN(
        P2_U3218) );
  OAI21_X1 U10384 ( .B1(n8986), .B2(n8902), .A(n8900), .ZN(n8909) );
  INV_X1 U10385 ( .A(n9495), .ZN(n9324) );
  NOR3_X1 U10386 ( .A1(n8902), .A2(n8901), .A3(n8984), .ZN(n8903) );
  OAI21_X1 U10387 ( .B1(n8903), .B2(n9013), .A(n9333), .ZN(n8907) );
  INV_X1 U10388 ( .A(n8904), .ZN(n9322) );
  NAND2_X1 U10389 ( .A1(P2_U3152), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n9129) );
  OAI21_X1 U10390 ( .B1(n9017), .B2(n8918), .A(n9129), .ZN(n8905) );
  AOI21_X1 U10391 ( .B1(n9322), .B2(n9014), .A(n8905), .ZN(n8906) );
  OAI211_X1 U10392 ( .C1(n9324), .C2(n8996), .A(n8907), .B(n8906), .ZN(n8908)
         );
  AOI21_X1 U10393 ( .B1(n8909), .B2(n9011), .A(n8908), .ZN(n8910) );
  INV_X1 U10394 ( .A(n8910), .ZN(P2_U3221) );
  INV_X1 U10395 ( .A(n8911), .ZN(n8912) );
  AOI21_X1 U10396 ( .B1(n8964), .B2(n8912), .A(n7677), .ZN(n8915) );
  NOR3_X1 U10397 ( .A1(n8913), .A2(n8918), .A3(n8984), .ZN(n8914) );
  OAI21_X1 U10398 ( .B1(n8915), .B2(n8914), .A(n8798), .ZN(n8921) );
  AOI22_X1 U10399 ( .A1(n8990), .A2(n9299), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3152), .ZN(n8917) );
  OAI21_X1 U10400 ( .B1(n8918), .B2(n8992), .A(n8917), .ZN(n8919) );
  AOI21_X1 U10401 ( .B1(n5096), .B2(n9014), .A(n8919), .ZN(n8920) );
  OAI211_X1 U10402 ( .C1(n9290), .C2(n8996), .A(n8921), .B(n8920), .ZN(
        P2_U3225) );
  NAND2_X1 U10403 ( .A1(n8923), .A2(n8922), .ZN(n8925) );
  NOR2_X1 U10404 ( .A1(n8925), .A2(n8924), .ZN(n9007) );
  NOR2_X1 U10405 ( .A1(n8984), .A2(n9385), .ZN(n9009) );
  INV_X1 U10406 ( .A(n8925), .ZN(n8927) );
  NOR2_X1 U10407 ( .A1(n8927), .A2(n8926), .ZN(n9008) );
  INV_X1 U10408 ( .A(n9008), .ZN(n8928) );
  AOI22_X1 U10409 ( .A1(n9007), .A2(n9011), .B1(n9009), .B2(n8928), .ZN(n8939)
         );
  XNOR2_X1 U10410 ( .A(n8930), .B(n8929), .ZN(n8931) );
  INV_X1 U10411 ( .A(n8931), .ZN(n8938) );
  NOR3_X1 U10412 ( .A1(n9007), .A2(n8931), .A3(n7677), .ZN(n8932) );
  OAI21_X1 U10413 ( .B1(n9008), .B2(n9010), .A(n8932), .ZN(n8937) );
  NAND2_X1 U10414 ( .A1(n9013), .A2(n9142), .ZN(n8933) );
  NAND2_X1 U10415 ( .A1(P2_U3152), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n9074) );
  OAI211_X1 U10416 ( .C1(n9387), .C2(n9017), .A(n8933), .B(n9074), .ZN(n8935)
         );
  NOR2_X1 U10417 ( .A1(n9512), .A2(n8996), .ZN(n8934) );
  AOI211_X1 U10418 ( .C1(n9014), .C2(n9397), .A(n8935), .B(n8934), .ZN(n8936)
         );
  OAI211_X1 U10419 ( .C1(n8939), .C2(n8938), .A(n8937), .B(n8936), .ZN(
        P2_U3228) );
  OAI211_X1 U10420 ( .C1(n8942), .C2(n8941), .A(n8940), .B(n9011), .ZN(n8948)
         );
  INV_X1 U10421 ( .A(n9374), .ZN(n8946) );
  NOR2_X1 U10422 ( .A1(n9027), .A2(n9384), .ZN(n8943) );
  AOI21_X1 U10423 ( .B1(n9333), .B2(n9412), .A(n8943), .ZN(n9368) );
  OAI22_X1 U10424 ( .A1(n8999), .A2(n9368), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8944), .ZN(n8945) );
  AOI21_X1 U10425 ( .B1(n9014), .B2(n8946), .A(n8945), .ZN(n8947) );
  OAI211_X1 U10426 ( .C1(n9372), .C2(n8996), .A(n8948), .B(n8947), .ZN(
        P2_U3230) );
  INV_X1 U10427 ( .A(n9468), .ZN(n9240) );
  INV_X1 U10428 ( .A(n8949), .ZN(n8950) );
  NAND2_X1 U10429 ( .A1(n8951), .A2(n8950), .ZN(n8953) );
  XNOR2_X1 U10430 ( .A(n8953), .B(n8952), .ZN(n8957) );
  OAI22_X1 U10431 ( .A1(n8957), .A2(n7677), .B1(n8954), .B2(n8984), .ZN(n8955)
         );
  NOR2_X1 U10432 ( .A1(n8992), .A2(n9281), .ZN(n8960) );
  OAI22_X1 U10433 ( .A1(n9243), .A2(n9017), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8958), .ZN(n8959) );
  AOI211_X1 U10434 ( .C1(n9014), .C2(n9238), .A(n8960), .B(n8959), .ZN(n8961)
         );
  INV_X1 U10435 ( .A(n9489), .ZN(n9308) );
  AOI21_X1 U10436 ( .B1(n8963), .B2(n8962), .A(n7677), .ZN(n8965) );
  NAND2_X1 U10437 ( .A1(n8965), .A2(n8964), .ZN(n8970) );
  INV_X1 U10438 ( .A(n8966), .ZN(n9306) );
  AOI22_X1 U10439 ( .A1(n8990), .A2(n9313), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3152), .ZN(n8967) );
  OAI21_X1 U10440 ( .B1(n9349), .B2(n8992), .A(n8967), .ZN(n8968) );
  AOI21_X1 U10441 ( .B1(n9306), .B2(n9014), .A(n8968), .ZN(n8969) );
  OAI211_X1 U10442 ( .C1(n9308), .C2(n8996), .A(n8970), .B(n8969), .ZN(
        P2_U3235) );
  OAI21_X1 U10443 ( .B1(n9017), .B2(n9012), .A(n8971), .ZN(n8972) );
  AOI21_X1 U10444 ( .B1(n9013), .B2(n8973), .A(n8972), .ZN(n8974) );
  OAI21_X1 U10445 ( .B1(n8975), .B2(n9002), .A(n8974), .ZN(n8980) );
  AOI211_X1 U10446 ( .C1(n8978), .C2(n8977), .A(n7677), .B(n8976), .ZN(n8979)
         );
  AOI211_X1 U10447 ( .C1(n9531), .C2(n9019), .A(n8980), .B(n8979), .ZN(n8981)
         );
  INV_X1 U10448 ( .A(n8981), .ZN(P2_U3236) );
  INV_X1 U10449 ( .A(n8982), .ZN(n8983) );
  AOI21_X1 U10450 ( .B1(n8940), .B2(n8983), .A(n7677), .ZN(n8988) );
  NOR3_X1 U10451 ( .A1(n8985), .A2(n9387), .A3(n8984), .ZN(n8987) );
  OAI21_X1 U10452 ( .B1(n8988), .B2(n8987), .A(n8986), .ZN(n8995) );
  INV_X1 U10453 ( .A(n9349), .ZN(n9312) );
  NOR2_X1 U10454 ( .A1(n8989), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9109) );
  AOI21_X1 U10455 ( .B1(n8990), .B2(n9312), .A(n9109), .ZN(n8991) );
  OAI21_X1 U10456 ( .B1(n9387), .B2(n8992), .A(n8991), .ZN(n8993) );
  AOI21_X1 U10457 ( .B1(n9343), .B2(n9014), .A(n8993), .ZN(n8994) );
  OAI211_X1 U10458 ( .C1(n9345), .C2(n8996), .A(n8995), .B(n8994), .ZN(
        P2_U3240) );
  XNOR2_X1 U10459 ( .A(n8998), .B(n8997), .ZN(n9006) );
  AOI22_X1 U10460 ( .A1(n9153), .A2(n9412), .B1(n9411), .B2(n9026), .ZN(n9211)
         );
  NOR2_X1 U10461 ( .A1(n9211), .A2(n8999), .ZN(n9004) );
  INV_X1 U10462 ( .A(n9000), .ZN(n9215) );
  OAI22_X1 U10463 ( .A1(n9215), .A2(n9002), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9001), .ZN(n9003) );
  AOI211_X1 U10464 ( .C1(n9461), .C2(n9019), .A(n9004), .B(n9003), .ZN(n9005)
         );
  OAI21_X1 U10465 ( .B1(n9006), .B2(n7677), .A(n9005), .ZN(P2_U3242) );
  NOR2_X1 U10466 ( .A1(n9008), .A2(n9007), .ZN(n9023) );
  INV_X1 U10467 ( .A(n9009), .ZN(n9022) );
  NAND3_X1 U10468 ( .A1(n9023), .A2(n9011), .A3(n9010), .ZN(n9021) );
  INV_X1 U10469 ( .A(n9012), .ZN(n9410) );
  AOI22_X1 U10470 ( .A1(n9013), .A2(n9410), .B1(P2_REG3_REG_15__SCAN_IN), .B2(
        P2_U3152), .ZN(n9016) );
  NAND2_X1 U10471 ( .A1(n9014), .A2(n9420), .ZN(n9015) );
  OAI211_X1 U10472 ( .C1(n9027), .C2(n9017), .A(n9016), .B(n9015), .ZN(n9018)
         );
  AOI21_X1 U10473 ( .B1(n9522), .B2(n9019), .A(n9018), .ZN(n9020) );
  OAI211_X1 U10474 ( .C1(n9023), .C2(n9022), .A(n9021), .B(n9020), .ZN(
        P2_U3243) );
  MUX2_X1 U10475 ( .A(n9024), .B(P2_DATAO_REG_29__SCAN_IN), .S(n9037), .Z(
        P2_U3581) );
  INV_X1 U10476 ( .A(n9198), .ZN(n9156) );
  MUX2_X1 U10477 ( .A(n9156), .B(P2_DATAO_REG_28__SCAN_IN), .S(n9037), .Z(
        P2_U3580) );
  MUX2_X1 U10478 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n9153), .S(P2_U3966), .Z(
        P2_U3579) );
  MUX2_X1 U10479 ( .A(n9025), .B(P2_DATAO_REG_26__SCAN_IN), .S(n9037), .Z(
        P2_U3578) );
  MUX2_X1 U10480 ( .A(n9026), .B(P2_DATAO_REG_25__SCAN_IN), .S(n9037), .Z(
        P2_U3577) );
  MUX2_X1 U10481 ( .A(n9251), .B(P2_DATAO_REG_24__SCAN_IN), .S(n9037), .Z(
        P2_U3576) );
  INV_X1 U10482 ( .A(n9281), .ZN(n9150) );
  MUX2_X1 U10483 ( .A(n9150), .B(P2_DATAO_REG_23__SCAN_IN), .S(n9037), .Z(
        P2_U3575) );
  MUX2_X1 U10484 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n9299), .S(P2_U3966), .Z(
        P2_U3574) );
  MUX2_X1 U10485 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n9313), .S(P2_U3966), .Z(
        P2_U3573) );
  MUX2_X1 U10486 ( .A(n9332), .B(P2_DATAO_REG_20__SCAN_IN), .S(n9037), .Z(
        P2_U3572) );
  MUX2_X1 U10487 ( .A(n9312), .B(P2_DATAO_REG_19__SCAN_IN), .S(n9037), .Z(
        P2_U3571) );
  MUX2_X1 U10488 ( .A(n9333), .B(P2_DATAO_REG_18__SCAN_IN), .S(n9037), .Z(
        P2_U3570) );
  INV_X1 U10489 ( .A(n9027), .ZN(n9413) );
  MUX2_X1 U10490 ( .A(n9413), .B(P2_DATAO_REG_16__SCAN_IN), .S(n9037), .Z(
        P2_U3568) );
  MUX2_X1 U10491 ( .A(n9142), .B(P2_DATAO_REG_15__SCAN_IN), .S(n9037), .Z(
        P2_U3567) );
  MUX2_X1 U10492 ( .A(n9410), .B(P2_DATAO_REG_14__SCAN_IN), .S(n9037), .Z(
        P2_U3566) );
  MUX2_X1 U10493 ( .A(n9028), .B(P2_DATAO_REG_13__SCAN_IN), .S(n9037), .Z(
        P2_U3565) );
  MUX2_X1 U10494 ( .A(n9029), .B(P2_DATAO_REG_11__SCAN_IN), .S(n9037), .Z(
        P2_U3563) );
  MUX2_X1 U10495 ( .A(n9030), .B(P2_DATAO_REG_10__SCAN_IN), .S(n9037), .Z(
        P2_U3562) );
  MUX2_X1 U10496 ( .A(n9031), .B(P2_DATAO_REG_9__SCAN_IN), .S(n9037), .Z(
        P2_U3561) );
  MUX2_X1 U10497 ( .A(n9032), .B(P2_DATAO_REG_8__SCAN_IN), .S(n9037), .Z(
        P2_U3560) );
  MUX2_X1 U10498 ( .A(n9033), .B(P2_DATAO_REG_7__SCAN_IN), .S(n9037), .Z(
        P2_U3559) );
  MUX2_X1 U10499 ( .A(n9034), .B(P2_DATAO_REG_6__SCAN_IN), .S(n9037), .Z(
        P2_U3558) );
  MUX2_X1 U10500 ( .A(n9035), .B(P2_DATAO_REG_4__SCAN_IN), .S(n9037), .Z(
        P2_U3556) );
  MUX2_X1 U10501 ( .A(n7346), .B(P2_DATAO_REG_3__SCAN_IN), .S(n9037), .Z(
        P2_U3555) );
  MUX2_X1 U10502 ( .A(n9036), .B(P2_DATAO_REG_2__SCAN_IN), .S(n9037), .Z(
        P2_U3554) );
  MUX2_X1 U10503 ( .A(n7141), .B(P2_DATAO_REG_1__SCAN_IN), .S(n9037), .Z(
        P2_U3553) );
  AOI211_X1 U10504 ( .C1(n9040), .C2(n9039), .A(n9112), .B(n9038), .ZN(n9041)
         );
  INV_X1 U10505 ( .A(n9041), .ZN(n9052) );
  NOR2_X1 U10506 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9042), .ZN(n9043) );
  AOI21_X1 U10507 ( .B1(n10358), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n9043), .ZN(
        n9051) );
  AND2_X1 U10508 ( .A1(n9045), .A2(n9044), .ZN(n9046) );
  OAI21_X1 U10509 ( .B1(n9047), .B2(n9046), .A(n10361), .ZN(n9050) );
  NAND2_X1 U10510 ( .A1(n10362), .A2(n9048), .ZN(n9049) );
  NAND4_X1 U10511 ( .A1(n9052), .A2(n9051), .A3(n9050), .A4(n9049), .ZN(
        P2_U3256) );
  XNOR2_X1 U10512 ( .A(n9077), .B(n9078), .ZN(n9055) );
  AOI21_X1 U10513 ( .B1(n9055), .B2(P2_REG2_REG_15__SCAN_IN), .A(n9079), .ZN(
        n9066) );
  AND2_X1 U10514 ( .A1(P2_U3152), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n9057) );
  NOR2_X1 U10515 ( .A1(n9101), .A2(n9068), .ZN(n9056) );
  AOI211_X1 U10516 ( .C1(n10358), .C2(P2_ADDR_REG_15__SCAN_IN), .A(n9057), .B(
        n9056), .ZN(n9065) );
  INV_X1 U10517 ( .A(n9060), .ZN(n9063) );
  NOR2_X1 U10518 ( .A1(n9061), .A2(n9060), .ZN(n9069) );
  INV_X1 U10519 ( .A(n9069), .ZN(n9062) );
  OAI211_X1 U10520 ( .C1(n9063), .C2(P2_REG1_REG_15__SCAN_IN), .A(n10366), .B(
        n9062), .ZN(n9064) );
  OAI211_X1 U10521 ( .C1(n9066), .C2(n9124), .A(n9065), .B(n9064), .ZN(
        P2_U3260) );
  NOR2_X1 U10522 ( .A1(n9068), .A2(n9067), .ZN(n9070) );
  XOR2_X1 U10523 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n9087), .Z(n9071) );
  OAI21_X1 U10524 ( .B1(n9072), .B2(n9071), .A(n9086), .ZN(n9076) );
  NAND2_X1 U10525 ( .A1(n10358), .A2(P2_ADDR_REG_16__SCAN_IN), .ZN(n9073) );
  OAI211_X1 U10526 ( .C1(n9101), .C2(n9093), .A(n9074), .B(n9073), .ZN(n9075)
         );
  AOI21_X1 U10527 ( .B1(n9076), .B2(n10366), .A(n9075), .ZN(n9085) );
  NOR2_X1 U10528 ( .A1(n9078), .A2(n9077), .ZN(n9080) );
  MUX2_X1 U10529 ( .A(P2_REG2_REG_16__SCAN_IN), .B(n9081), .S(n9087), .Z(n9082) );
  NAND2_X1 U10530 ( .A1(n9082), .A2(n9083), .ZN(n9092) );
  OAI211_X1 U10531 ( .C1(n9083), .C2(n9082), .A(n10361), .B(n9092), .ZN(n9084)
         );
  NAND2_X1 U10532 ( .A1(n9085), .A2(n9084), .ZN(P2_U3261) );
  INV_X1 U10533 ( .A(n9107), .ZN(n9100) );
  AND2_X1 U10534 ( .A1(P2_U3152), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n9091) );
  XNOR2_X1 U10535 ( .A(n9107), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n9088) );
  AOI211_X1 U10536 ( .C1(n9089), .C2(n9088), .A(n9106), .B(n9112), .ZN(n9090)
         );
  AOI211_X1 U10537 ( .C1(n10358), .C2(P2_ADDR_REG_17__SCAN_IN), .A(n9091), .B(
        n9090), .ZN(n9099) );
  OAI21_X1 U10538 ( .B1(n9093), .B2(n9081), .A(n9092), .ZN(n9097) );
  INV_X1 U10539 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n9094) );
  MUX2_X1 U10540 ( .A(n9094), .B(P2_REG2_REG_17__SCAN_IN), .S(n9107), .Z(n9095) );
  INV_X1 U10541 ( .A(n9095), .ZN(n9096) );
  NAND2_X1 U10542 ( .A1(n9096), .A2(n9097), .ZN(n9102) );
  OAI211_X1 U10543 ( .C1(n9097), .C2(n9096), .A(n10361), .B(n9102), .ZN(n9098)
         );
  OAI211_X1 U10544 ( .C1(n9101), .C2(n9100), .A(n9099), .B(n9098), .ZN(
        P2_U3262) );
  NAND2_X1 U10545 ( .A1(P2_REG2_REG_17__SCAN_IN), .A2(n9107), .ZN(n9103) );
  NAND2_X1 U10546 ( .A1(n9103), .A2(n9102), .ZN(n9104) );
  NOR2_X1 U10547 ( .A1(n9104), .A2(n9120), .ZN(n9116) );
  AOI21_X1 U10548 ( .B1(n9105), .B2(P2_REG2_REG_18__SCAN_IN), .A(n9117), .ZN(
        n9115) );
  INV_X1 U10549 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n9108) );
  XNOR2_X1 U10550 ( .A(n9120), .B(n9108), .ZN(n9119) );
  XOR2_X1 U10551 ( .A(n9118), .B(n9119), .Z(n9111) );
  AOI21_X1 U10552 ( .B1(n10358), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n9109), .ZN(
        n9110) );
  OAI21_X1 U10553 ( .B1(n9112), .B2(n9111), .A(n9110), .ZN(n9113) );
  AOI21_X1 U10554 ( .B1(n9120), .B2(n10362), .A(n9113), .ZN(n9114) );
  OAI21_X1 U10555 ( .B1(n9115), .B2(n9124), .A(n9114), .ZN(P2_U3263) );
  OR2_X1 U10556 ( .A1(n9120), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n9121) );
  AOI22_X1 U10557 ( .A1(n9125), .A2(n10361), .B1(n9123), .B2(n10366), .ZN(
        n9128) );
  NOR2_X1 U10558 ( .A1(n9125), .A2(n9124), .ZN(n9126) );
  OAI211_X1 U10559 ( .C1(n9132), .C2(n9131), .A(n9130), .B(n9129), .ZN(
        P2_U3264) );
  AOI21_X1 U10560 ( .B1(n9432), .B2(n9167), .A(n9133), .ZN(n9433) );
  INV_X1 U10561 ( .A(n9433), .ZN(n9138) );
  OAI21_X1 U10562 ( .B1(n9427), .B2(n9135), .A(n9134), .ZN(n9136) );
  AOI21_X1 U10563 ( .B1(n9432), .B2(n9422), .A(n9136), .ZN(n9137) );
  OAI21_X1 U10564 ( .B1(n9138), .B2(n9425), .A(n9137), .ZN(P2_U3266) );
  OR2_X1 U10565 ( .A1(n9526), .A2(n9410), .ZN(n9139) );
  INV_X1 U10566 ( .A(n9408), .ZN(n9141) );
  OR2_X1 U10567 ( .A1(n9522), .A2(n9142), .ZN(n9143) );
  NAND2_X1 U10568 ( .A1(n9144), .A2(n9143), .ZN(n9379) );
  INV_X1 U10569 ( .A(n9379), .ZN(n9145) );
  NAND2_X1 U10570 ( .A1(n9145), .A2(n9388), .ZN(n9383) );
  NAND2_X1 U10571 ( .A1(n9398), .A2(n9413), .ZN(n9146) );
  NAND2_X1 U10572 ( .A1(n9345), .A2(n9147), .ZN(n9148) );
  NAND2_X1 U10573 ( .A1(n9484), .A2(n9313), .ZN(n9149) );
  NAND2_X1 U10574 ( .A1(n9475), .A2(n9150), .ZN(n9220) );
  NOR2_X1 U10575 ( .A1(n9468), .A2(n9251), .ZN(n9221) );
  AOI22_X1 U10576 ( .A1(n9228), .A2(n9221), .B1(n5057), .B2(n9243), .ZN(n9151)
         );
  INV_X1 U10577 ( .A(n9179), .ZN(n9155) );
  INV_X1 U10578 ( .A(n9446), .ZN(n9157) );
  NOR2_X1 U10579 ( .A1(n9452), .A2(n9156), .ZN(n9439) );
  XNOR2_X1 U10580 ( .A(n9158), .B(n9440), .ZN(n9176) );
  INV_X1 U10581 ( .A(n9440), .ZN(n9159) );
  OAI22_X1 U10582 ( .A1(n9198), .A2(n9384), .B1(n9162), .B2(n9161), .ZN(n9163)
         );
  INV_X1 U10583 ( .A(n9447), .ZN(n9174) );
  INV_X1 U10584 ( .A(n9183), .ZN(n9165) );
  NAND2_X1 U10585 ( .A1(n9438), .A2(n9165), .ZN(n9166) );
  NAND2_X1 U10586 ( .A1(n9167), .A2(n9166), .ZN(n9443) );
  NOR2_X1 U10587 ( .A1(n9443), .A2(n9425), .ZN(n9173) );
  INV_X1 U10588 ( .A(n9168), .ZN(n9169) );
  AOI22_X1 U10589 ( .A1(n9169), .A2(n9419), .B1(P2_REG2_REG_29__SCAN_IN), .B2(
        n9404), .ZN(n9170) );
  OAI21_X1 U10590 ( .B1(n9171), .B2(n9371), .A(n9170), .ZN(n9172) );
  AOI211_X1 U10591 ( .C1(n9174), .C2(n9427), .A(n9173), .B(n9172), .ZN(n9175)
         );
  OAI21_X1 U10592 ( .B1(n9176), .B2(n9429), .A(n9175), .ZN(P2_U3267) );
  XNOR2_X1 U10593 ( .A(n9177), .B(n9179), .ZN(n9453) );
  OAI211_X1 U10594 ( .C1(n9180), .C2(n9179), .A(n9178), .B(n4402), .ZN(n9182)
         );
  AOI211_X1 U10595 ( .C1(n9452), .C2(n9192), .A(n9518), .B(n9183), .ZN(n9451)
         );
  NAND2_X1 U10596 ( .A1(n9451), .A2(n9184), .ZN(n9188) );
  INV_X1 U10597 ( .A(n9185), .ZN(n9186) );
  AOI22_X1 U10598 ( .A1(n9186), .A2(n9419), .B1(P2_REG2_REG_28__SCAN_IN), .B2(
        n9404), .ZN(n9187) );
  OAI211_X1 U10599 ( .C1(n9189), .C2(n9371), .A(n9188), .B(n9187), .ZN(n9190)
         );
  AOI21_X1 U10600 ( .B1(n9450), .B2(n9427), .A(n9190), .ZN(n9191) );
  OAI21_X1 U10601 ( .B1(n9453), .B2(n9429), .A(n9191), .ZN(P2_U3268) );
  AOI21_X1 U10602 ( .B1(n9454), .B2(n9212), .A(n5066), .ZN(n9455) );
  AOI22_X1 U10603 ( .A1(n9193), .A2(n9419), .B1(P2_REG2_REG_27__SCAN_IN), .B2(
        n9404), .ZN(n9194) );
  OAI21_X1 U10604 ( .B1(n4985), .B2(n9371), .A(n9194), .ZN(n9203) );
  AOI21_X1 U10605 ( .B1(n9196), .B2(n9195), .A(n9406), .ZN(n9201) );
  OAI22_X1 U10606 ( .A1(n9198), .A2(n9386), .B1(n9197), .B2(n9384), .ZN(n9199)
         );
  AOI21_X1 U10607 ( .B1(n9201), .B2(n9200), .A(n9199), .ZN(n9457) );
  NOR2_X1 U10608 ( .A1(n9457), .A2(n9404), .ZN(n9202) );
  AOI211_X1 U10609 ( .C1(n9354), .C2(n9455), .A(n9203), .B(n9202), .ZN(n9204)
         );
  OAI21_X1 U10610 ( .B1(n9458), .B2(n9429), .A(n9204), .ZN(P2_U3269) );
  XNOR2_X1 U10611 ( .A(n9205), .B(n4979), .ZN(n9462) );
  AOI22_X1 U10612 ( .A1(n9461), .A2(n9422), .B1(P2_REG2_REG_26__SCAN_IN), .B2(
        n9404), .ZN(n9219) );
  NOR2_X1 U10613 ( .A1(n9229), .A2(n9228), .ZN(n9227) );
  NOR2_X1 U10614 ( .A1(n9227), .A2(n5886), .ZN(n9209) );
  XNOR2_X1 U10615 ( .A(n9209), .B(n4979), .ZN(n9210) );
  INV_X1 U10616 ( .A(n9222), .ZN(n9214) );
  INV_X1 U10617 ( .A(n9212), .ZN(n9213) );
  AOI211_X1 U10618 ( .C1(n9461), .C2(n9214), .A(n9518), .B(n9213), .ZN(n9460)
         );
  INV_X1 U10619 ( .A(n9460), .ZN(n9216) );
  OAI22_X1 U10620 ( .A1(n9216), .A2(n9361), .B1(n9373), .B2(n9215), .ZN(n9217)
         );
  OAI21_X1 U10621 ( .B1(n9459), .B2(n9217), .A(n9427), .ZN(n9218) );
  OAI211_X1 U10622 ( .C1(n9462), .C2(n9429), .A(n9219), .B(n9218), .ZN(
        P2_U3270) );
  INV_X1 U10623 ( .A(n9242), .ZN(n9237) );
  AOI211_X1 U10624 ( .C1(n9464), .C2(n9223), .A(n9518), .B(n9222), .ZN(n9463)
         );
  INV_X1 U10625 ( .A(n9224), .ZN(n9225) );
  AOI22_X1 U10626 ( .A1(n9225), .A2(n9419), .B1(P2_REG2_REG_25__SCAN_IN), .B2(
        n9404), .ZN(n9226) );
  OAI21_X1 U10627 ( .B1(n5057), .B2(n9371), .A(n9226), .ZN(n9233) );
  AOI211_X1 U10628 ( .C1(n9229), .C2(n9228), .A(n9406), .B(n9227), .ZN(n9231)
         );
  NOR2_X1 U10629 ( .A1(n9231), .A2(n9230), .ZN(n9466) );
  NOR2_X1 U10630 ( .A1(n9466), .A2(n9404), .ZN(n9232) );
  AOI211_X1 U10631 ( .C1(n9463), .C2(n9337), .A(n9233), .B(n9232), .ZN(n9234)
         );
  OAI21_X1 U10632 ( .B1(n9467), .B2(n9429), .A(n9234), .ZN(P2_U3271) );
  AOI21_X1 U10633 ( .B1(n9237), .B2(n9236), .A(n9235), .ZN(n9472) );
  XOR2_X1 U10634 ( .A(n9256), .B(n9468), .Z(n9469) );
  AOI22_X1 U10635 ( .A1(n9421), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n9238), .B2(
        n9419), .ZN(n9239) );
  OAI21_X1 U10636 ( .B1(n9240), .B2(n9371), .A(n9239), .ZN(n9247) );
  AOI211_X1 U10637 ( .C1(n9242), .C2(n9241), .A(n9406), .B(n4450), .ZN(n9245)
         );
  OAI22_X1 U10638 ( .A1(n9243), .A2(n9386), .B1(n9281), .B2(n9384), .ZN(n9244)
         );
  NOR2_X1 U10639 ( .A1(n9245), .A2(n9244), .ZN(n9471) );
  NOR2_X1 U10640 ( .A1(n9471), .A2(n9404), .ZN(n9246) );
  AOI211_X1 U10641 ( .C1(n9469), .C2(n9354), .A(n9247), .B(n9246), .ZN(n9248)
         );
  OAI21_X1 U10642 ( .B1(n9472), .B2(n9429), .A(n9248), .ZN(P2_U3272) );
  OAI21_X1 U10643 ( .B1(n9254), .B2(n9250), .A(n9249), .ZN(n9252) );
  AOI222_X1 U10644 ( .A1(n4402), .A2(n9252), .B1(n9251), .B2(n9412), .C1(n9299), .C2(n9411), .ZN(n9478) );
  NAND2_X1 U10645 ( .A1(n9253), .A2(n9254), .ZN(n9473) );
  NAND3_X1 U10646 ( .A1(n9474), .A2(n9255), .A3(n9473), .ZN(n9264) );
  INV_X1 U10647 ( .A(n9266), .ZN(n9258) );
  INV_X1 U10648 ( .A(n9256), .ZN(n9257) );
  AOI21_X1 U10649 ( .B1(n9475), .B2(n9258), .A(n9257), .ZN(n9476) );
  AOI22_X1 U10650 ( .A1(n9421), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n9259), .B2(
        n9419), .ZN(n9260) );
  OAI21_X1 U10651 ( .B1(n9261), .B2(n9371), .A(n9260), .ZN(n9262) );
  AOI21_X1 U10652 ( .B1(n9476), .B2(n9354), .A(n9262), .ZN(n9263) );
  OAI211_X1 U10653 ( .C1(n9404), .C2(n9478), .A(n9264), .B(n9263), .ZN(
        P2_U3273) );
  XOR2_X1 U10654 ( .A(n9265), .B(n9278), .Z(n9483) );
  AOI21_X1 U10655 ( .B1(n5593), .B2(n9267), .A(n9266), .ZN(n9480) );
  INV_X1 U10656 ( .A(n5593), .ZN(n9270) );
  AOI22_X1 U10657 ( .A1(n9421), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n9268), .B2(
        n9419), .ZN(n9269) );
  OAI21_X1 U10658 ( .B1(n9270), .B2(n9371), .A(n9269), .ZN(n9286) );
  NAND2_X1 U10659 ( .A1(n9391), .A2(n9271), .ZN(n9273) );
  NAND2_X1 U10660 ( .A1(n9273), .A2(n9272), .ZN(n9330) );
  NAND2_X1 U10661 ( .A1(n9330), .A2(n9274), .ZN(n9276) );
  NAND2_X1 U10662 ( .A1(n9276), .A2(n9275), .ZN(n9279) );
  INV_X1 U10663 ( .A(n9279), .ZN(n9277) );
  AOI21_X1 U10664 ( .B1(n9277), .B2(n4636), .A(n9406), .ZN(n9284) );
  NAND2_X1 U10665 ( .A1(n9279), .A2(n9278), .ZN(n9283) );
  OAI22_X1 U10666 ( .A1(n9281), .A2(n9386), .B1(n9280), .B2(n9384), .ZN(n9282)
         );
  AOI21_X1 U10667 ( .B1(n9284), .B2(n9283), .A(n9282), .ZN(n9482) );
  NOR2_X1 U10668 ( .A1(n9482), .A2(n9404), .ZN(n9285) );
  AOI211_X1 U10669 ( .C1(n9480), .C2(n9354), .A(n9286), .B(n9285), .ZN(n9287)
         );
  OAI21_X1 U10670 ( .B1(n9483), .B2(n9429), .A(n9287), .ZN(P2_U3274) );
  XNOR2_X1 U10671 ( .A(n9288), .B(n9297), .ZN(n9488) );
  XNOR2_X1 U10672 ( .A(n9484), .B(n9305), .ZN(n9485) );
  AOI22_X1 U10673 ( .A1(n9421), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n5096), .B2(
        n9419), .ZN(n9289) );
  OAI21_X1 U10674 ( .B1(n9290), .B2(n9371), .A(n9289), .ZN(n9302) );
  NAND2_X1 U10675 ( .A1(n9330), .A2(n9291), .ZN(n9293) );
  NAND2_X1 U10676 ( .A1(n9293), .A2(n9292), .ZN(n9295) );
  INV_X1 U10677 ( .A(n9295), .ZN(n9298) );
  INV_X1 U10678 ( .A(n9297), .ZN(n9294) );
  OR2_X1 U10679 ( .A1(n9295), .A2(n9294), .ZN(n9296) );
  OAI21_X1 U10680 ( .B1(n9298), .B2(n9297), .A(n9296), .ZN(n9300) );
  AOI222_X1 U10681 ( .A1(n4402), .A2(n9300), .B1(n9299), .B2(n9412), .C1(n9332), .C2(n9411), .ZN(n9487) );
  NOR2_X1 U10682 ( .A1(n9487), .A2(n9404), .ZN(n9301) );
  AOI211_X1 U10683 ( .C1(n9485), .C2(n9354), .A(n9302), .B(n9301), .ZN(n9303)
         );
  OAI21_X1 U10684 ( .B1(n9488), .B2(n9429), .A(n9303), .ZN(P2_U3275) );
  XNOR2_X1 U10685 ( .A(n9304), .B(n9311), .ZN(n9493) );
  AOI21_X1 U10686 ( .B1(n9489), .B2(n9320), .A(n9305), .ZN(n9490) );
  AOI22_X1 U10687 ( .A1(n9421), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n9306), .B2(
        n9419), .ZN(n9307) );
  OAI21_X1 U10688 ( .B1(n9308), .B2(n9371), .A(n9307), .ZN(n9316) );
  NAND2_X1 U10689 ( .A1(n9330), .A2(n9309), .ZN(n9310) );
  XOR2_X1 U10690 ( .A(n9311), .B(n9310), .Z(n9314) );
  AOI222_X1 U10691 ( .A1(n4402), .A2(n9314), .B1(n9313), .B2(n9412), .C1(n9312), .C2(n9411), .ZN(n9492) );
  NOR2_X1 U10692 ( .A1(n9492), .A2(n9404), .ZN(n9315) );
  AOI211_X1 U10693 ( .C1(n9490), .C2(n9354), .A(n9316), .B(n9315), .ZN(n9317)
         );
  OAI21_X1 U10694 ( .B1(n9429), .B2(n9493), .A(n9317), .ZN(P2_U3276) );
  XNOR2_X1 U10695 ( .A(n9319), .B(n9318), .ZN(n9498) );
  INV_X1 U10696 ( .A(n9320), .ZN(n9321) );
  AOI211_X1 U10697 ( .C1(n9495), .C2(n9341), .A(n9518), .B(n9321), .ZN(n9494)
         );
  AOI22_X1 U10698 ( .A1(n9421), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n9322), .B2(
        n9419), .ZN(n9323) );
  OAI21_X1 U10699 ( .B1(n9324), .B2(n9371), .A(n9323), .ZN(n9336) );
  NOR2_X1 U10700 ( .A1(n9364), .A2(n9325), .ZN(n9326) );
  NOR2_X1 U10701 ( .A1(n9362), .A2(n9327), .ZN(n9348) );
  NOR2_X1 U10702 ( .A1(n9348), .A2(n9347), .ZN(n9346) );
  OAI21_X1 U10703 ( .B1(n9346), .B2(n9329), .A(n9328), .ZN(n9331) );
  NAND2_X1 U10704 ( .A1(n9331), .A2(n9330), .ZN(n9334) );
  AOI222_X1 U10705 ( .A1(n4402), .A2(n9334), .B1(n9333), .B2(n9411), .C1(n9332), .C2(n9412), .ZN(n9497) );
  NOR2_X1 U10706 ( .A1(n9497), .A2(n9404), .ZN(n9335) );
  AOI211_X1 U10707 ( .C1(n9494), .C2(n9337), .A(n9336), .B(n9335), .ZN(n9338)
         );
  OAI21_X1 U10708 ( .B1(n9429), .B2(n9498), .A(n9338), .ZN(P2_U3277) );
  XNOR2_X1 U10709 ( .A(n9339), .B(n9347), .ZN(n9503) );
  INV_X1 U10710 ( .A(n9341), .ZN(n9342) );
  AOI21_X1 U10711 ( .B1(n9499), .B2(n9340), .A(n9342), .ZN(n9500) );
  AOI22_X1 U10712 ( .A1(n9421), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n9343), .B2(
        n9419), .ZN(n9344) );
  OAI21_X1 U10713 ( .B1(n9345), .B2(n9371), .A(n9344), .ZN(n9353) );
  AOI211_X1 U10714 ( .C1(n9348), .C2(n9347), .A(n9406), .B(n9346), .ZN(n9351)
         );
  OAI22_X1 U10715 ( .A1(n9349), .A2(n9386), .B1(n9387), .B2(n9384), .ZN(n9350)
         );
  NOR2_X1 U10716 ( .A1(n9351), .A2(n9350), .ZN(n9502) );
  NOR2_X1 U10717 ( .A1(n9502), .A2(n9404), .ZN(n9352) );
  AOI211_X1 U10718 ( .C1(n9500), .C2(n9354), .A(n9353), .B(n9352), .ZN(n9355)
         );
  OAI21_X1 U10719 ( .B1(n9503), .B2(n9429), .A(n9355), .ZN(P2_U3278) );
  INV_X1 U10720 ( .A(n9356), .ZN(n9360) );
  NAND2_X1 U10721 ( .A1(n9358), .A2(n9357), .ZN(n9359) );
  NAND2_X1 U10722 ( .A1(n9360), .A2(n9359), .ZN(n9504) );
  OAI211_X1 U10723 ( .C1(n9396), .C2(n9372), .A(n10409), .B(n9340), .ZN(n9505)
         );
  NOR2_X1 U10724 ( .A1(n9505), .A2(n9361), .ZN(n9370) );
  INV_X1 U10725 ( .A(n9362), .ZN(n9367) );
  NAND2_X1 U10726 ( .A1(n9391), .A2(n9363), .ZN(n9365) );
  NAND2_X1 U10727 ( .A1(n9365), .A2(n9364), .ZN(n9366) );
  NAND3_X1 U10728 ( .A1(n9367), .A2(n4402), .A3(n9366), .ZN(n9369) );
  NAND2_X1 U10729 ( .A1(n9369), .A2(n9368), .ZN(n9506) );
  AOI211_X1 U10730 ( .C1(n9394), .C2(n9504), .A(n9370), .B(n9506), .ZN(n9378)
         );
  NOR2_X1 U10731 ( .A1(n9372), .A2(n9371), .ZN(n9376) );
  OAI22_X1 U10732 ( .A1(n9427), .A2(n9094), .B1(n9374), .B2(n9373), .ZN(n9375)
         );
  AOI211_X1 U10733 ( .C1(n9504), .C2(n9402), .A(n9376), .B(n9375), .ZN(n9377)
         );
  OAI21_X1 U10734 ( .B1(n9378), .B2(n9404), .A(n9377), .ZN(P2_U3279) );
  NAND2_X1 U10735 ( .A1(n9379), .A2(n9380), .ZN(n9382) );
  OAI22_X1 U10736 ( .A1(n9387), .A2(n9386), .B1(n9385), .B2(n9384), .ZN(n9393)
         );
  NAND2_X1 U10737 ( .A1(n9389), .A2(n9388), .ZN(n9390) );
  AOI21_X1 U10738 ( .B1(n9391), .B2(n9390), .A(n9406), .ZN(n9392) );
  AOI211_X1 U10739 ( .C1(n9511), .C2(n9394), .A(n9393), .B(n9392), .ZN(n9516)
         );
  NOR2_X1 U10740 ( .A1(n9417), .A2(n9512), .ZN(n9395) );
  OR2_X1 U10741 ( .A1(n9396), .A2(n9395), .ZN(n9513) );
  AOI22_X1 U10742 ( .A1(n9421), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n9397), .B2(
        n9419), .ZN(n9400) );
  NAND2_X1 U10743 ( .A1(n9398), .A2(n9422), .ZN(n9399) );
  OAI211_X1 U10744 ( .C1(n9513), .C2(n9425), .A(n9400), .B(n9399), .ZN(n9401)
         );
  AOI21_X1 U10745 ( .B1(n9511), .B2(n9402), .A(n9401), .ZN(n9403) );
  OAI21_X1 U10746 ( .B1(n9516), .B2(n9404), .A(n9403), .ZN(P2_U3280) );
  XNOR2_X1 U10747 ( .A(n9405), .B(n9408), .ZN(n9524) );
  OAI211_X1 U10748 ( .C1(n9409), .C2(n9408), .A(n9407), .B(n4402), .ZN(n9415)
         );
  AOI22_X1 U10749 ( .A1(n9413), .A2(n9412), .B1(n9411), .B2(n9410), .ZN(n9414)
         );
  NAND2_X1 U10750 ( .A1(n9415), .A2(n9414), .ZN(n9520) );
  AND2_X1 U10751 ( .A1(n9416), .A2(n9522), .ZN(n9418) );
  OR2_X1 U10752 ( .A1(n9418), .A2(n9417), .ZN(n9519) );
  AOI22_X1 U10753 ( .A1(n9421), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n9420), .B2(
        n9419), .ZN(n9424) );
  NAND2_X1 U10754 ( .A1(n9522), .A2(n9422), .ZN(n9423) );
  OAI211_X1 U10755 ( .C1(n9519), .C2(n9425), .A(n9424), .B(n9423), .ZN(n9426)
         );
  AOI21_X1 U10756 ( .B1(n9520), .B2(n9427), .A(n9426), .ZN(n9428) );
  OAI21_X1 U10757 ( .B1(n9524), .B2(n9429), .A(n9428), .ZN(P2_U3281) );
  AOI21_X1 U10758 ( .B1(n8844), .B2(n10408), .A(n9434), .ZN(n9430) );
  OAI21_X1 U10759 ( .B1(n9431), .B2(n9518), .A(n9430), .ZN(n9560) );
  MUX2_X1 U10760 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n9560), .S(n10426), .Z(
        P2_U3551) );
  INV_X1 U10761 ( .A(n9432), .ZN(n9437) );
  NAND2_X1 U10762 ( .A1(n9433), .A2(n10409), .ZN(n9436) );
  INV_X1 U10763 ( .A(n9434), .ZN(n9435) );
  OAI211_X1 U10764 ( .C1(n9437), .C2(n10403), .A(n9436), .B(n9435), .ZN(n9561)
         );
  MUX2_X1 U10765 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n9561), .S(n10426), .Z(
        P2_U3550) );
  NOR3_X1 U10766 ( .A1(n9440), .A2(n10414), .A3(n9439), .ZN(n9445) );
  NAND2_X1 U10767 ( .A1(n9438), .A2(n10408), .ZN(n9442) );
  NAND3_X1 U10768 ( .A1(n9440), .A2(n9439), .A3(n10399), .ZN(n9441) );
  OAI211_X1 U10769 ( .C1(n9443), .C2(n9518), .A(n9442), .B(n9441), .ZN(n9444)
         );
  AOI21_X1 U10770 ( .B1(n9446), .B2(n9445), .A(n9444), .ZN(n9448) );
  NAND3_X1 U10771 ( .A1(n9449), .A2(n9448), .A3(n9447), .ZN(n9562) );
  MUX2_X1 U10772 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n9562), .S(n10426), .Z(
        P2_U3549) );
  AOI22_X1 U10773 ( .A1(n9455), .A2(n10409), .B1(n10408), .B2(n9454), .ZN(
        n9456) );
  OAI211_X1 U10774 ( .C1(n9458), .C2(n10414), .A(n9457), .B(n9456), .ZN(n9564)
         );
  MUX2_X1 U10775 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n9564), .S(n10426), .Z(
        P2_U3547) );
  MUX2_X1 U10776 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n9565), .S(n10426), .Z(
        P2_U3546) );
  AOI21_X1 U10777 ( .B1(n10408), .B2(n9464), .A(n9463), .ZN(n9465) );
  MUX2_X1 U10778 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n9566), .S(n10426), .Z(
        P2_U3545) );
  AOI22_X1 U10779 ( .A1(n9469), .A2(n10409), .B1(n10408), .B2(n9468), .ZN(
        n9470) );
  OAI211_X1 U10780 ( .C1(n9472), .C2(n10414), .A(n9471), .B(n9470), .ZN(n9567)
         );
  MUX2_X1 U10781 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n9567), .S(n10426), .Z(
        P2_U3544) );
  NAND3_X1 U10782 ( .A1(n9474), .A2(n10399), .A3(n9473), .ZN(n9479) );
  AOI22_X1 U10783 ( .A1(n9476), .A2(n10409), .B1(n10408), .B2(n9475), .ZN(
        n9477) );
  NAND3_X1 U10784 ( .A1(n9479), .A2(n9478), .A3(n9477), .ZN(n9568) );
  MUX2_X1 U10785 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n9568), .S(n10426), .Z(
        P2_U3543) );
  AOI22_X1 U10786 ( .A1(n9480), .A2(n10409), .B1(n10408), .B2(n5593), .ZN(
        n9481) );
  OAI211_X1 U10787 ( .C1(n9483), .C2(n10414), .A(n9482), .B(n9481), .ZN(n9569)
         );
  MUX2_X1 U10788 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n9569), .S(n10426), .Z(
        P2_U3542) );
  AOI22_X1 U10789 ( .A1(n9485), .A2(n10409), .B1(n10408), .B2(n9484), .ZN(
        n9486) );
  OAI211_X1 U10790 ( .C1(n9488), .C2(n10414), .A(n9487), .B(n9486), .ZN(n9570)
         );
  MUX2_X1 U10791 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n9570), .S(n10426), .Z(
        P2_U3541) );
  AOI22_X1 U10792 ( .A1(n9490), .A2(n10409), .B1(n10408), .B2(n9489), .ZN(
        n9491) );
  OAI211_X1 U10793 ( .C1(n9493), .C2(n10414), .A(n9492), .B(n9491), .ZN(n9571)
         );
  MUX2_X1 U10794 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n9571), .S(n10426), .Z(
        P2_U3540) );
  AOI21_X1 U10795 ( .B1(n10408), .B2(n9495), .A(n9494), .ZN(n9496) );
  OAI211_X1 U10796 ( .C1(n10414), .C2(n9498), .A(n9497), .B(n9496), .ZN(n9572)
         );
  MUX2_X1 U10797 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n9572), .S(n10426), .Z(
        P2_U3539) );
  AOI22_X1 U10798 ( .A1(n9500), .A2(n10409), .B1(n10408), .B2(n9499), .ZN(
        n9501) );
  OAI211_X1 U10799 ( .C1(n10414), .C2(n9503), .A(n9502), .B(n9501), .ZN(n9573)
         );
  MUX2_X1 U10800 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n9573), .S(n10426), .Z(
        P2_U3538) );
  INV_X1 U10801 ( .A(n9504), .ZN(n9510) );
  INV_X1 U10802 ( .A(n9505), .ZN(n9507) );
  AOI211_X1 U10803 ( .C1(n10408), .C2(n9508), .A(n9507), .B(n9506), .ZN(n9509)
         );
  OAI21_X1 U10804 ( .B1(n10414), .B2(n9510), .A(n9509), .ZN(n9574) );
  MUX2_X1 U10805 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n9574), .S(n10426), .Z(
        P2_U3537) );
  INV_X1 U10806 ( .A(n9511), .ZN(n9517) );
  OAI22_X1 U10807 ( .A1(n9513), .A2(n9518), .B1(n9512), .B2(n10403), .ZN(n9514) );
  INV_X1 U10808 ( .A(n9514), .ZN(n9515) );
  OAI211_X1 U10809 ( .C1(n9556), .C2(n9517), .A(n9516), .B(n9515), .ZN(n9575)
         );
  MUX2_X1 U10810 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n9575), .S(n10426), .Z(
        P2_U3536) );
  NOR2_X1 U10811 ( .A1(n9519), .A2(n9518), .ZN(n9521) );
  AOI211_X1 U10812 ( .C1(n10408), .C2(n9522), .A(n9521), .B(n9520), .ZN(n9523)
         );
  OAI21_X1 U10813 ( .B1(n10414), .B2(n9524), .A(n9523), .ZN(n9576) );
  MUX2_X1 U10814 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n9576), .S(n10426), .Z(
        P2_U3535) );
  INV_X1 U10815 ( .A(n9525), .ZN(n9530) );
  AOI22_X1 U10816 ( .A1(n9527), .A2(n10409), .B1(n10408), .B2(n9526), .ZN(
        n9528) );
  OAI211_X1 U10817 ( .C1(n10414), .C2(n9530), .A(n9529), .B(n9528), .ZN(n9577)
         );
  MUX2_X1 U10818 ( .A(n9577), .B(P2_REG1_REG_14__SCAN_IN), .S(n10424), .Z(
        P2_U3534) );
  AOI22_X1 U10819 ( .A1(n9532), .A2(n10409), .B1(n10408), .B2(n9531), .ZN(
        n9533) );
  OAI211_X1 U10820 ( .C1(n9556), .C2(n9535), .A(n9534), .B(n9533), .ZN(n9578)
         );
  MUX2_X1 U10821 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n9578), .S(n10426), .Z(
        P2_U3533) );
  AOI22_X1 U10822 ( .A1(n9537), .A2(n10409), .B1(n10408), .B2(n9536), .ZN(
        n9538) );
  OAI211_X1 U10823 ( .C1(n10414), .C2(n9540), .A(n9539), .B(n9538), .ZN(n9579)
         );
  MUX2_X1 U10824 ( .A(n9579), .B(P2_REG1_REG_12__SCAN_IN), .S(n10424), .Z(
        P2_U3532) );
  AOI22_X1 U10825 ( .A1(n9542), .A2(n10409), .B1(n10408), .B2(n9541), .ZN(
        n9543) );
  OAI211_X1 U10826 ( .C1(n10414), .C2(n9545), .A(n9544), .B(n9543), .ZN(n9580)
         );
  MUX2_X1 U10827 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n9580), .S(n10426), .Z(
        P2_U3531) );
  INV_X1 U10828 ( .A(n9546), .ZN(n9550) );
  AOI22_X1 U10829 ( .A1(n9548), .A2(n10409), .B1(n10408), .B2(n9547), .ZN(
        n9549) );
  OAI211_X1 U10830 ( .C1(n9556), .C2(n9551), .A(n9550), .B(n9549), .ZN(n9581)
         );
  MUX2_X1 U10831 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n9581), .S(n10426), .Z(
        P2_U3530) );
  AOI22_X1 U10832 ( .A1(n9553), .A2(n10409), .B1(n10408), .B2(n9552), .ZN(
        n9554) );
  OAI211_X1 U10833 ( .C1(n9557), .C2(n9556), .A(n9555), .B(n9554), .ZN(n9582)
         );
  MUX2_X1 U10834 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n9582), .S(n10426), .Z(
        P2_U3528) );
  MUX2_X1 U10835 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n9558), .S(n10426), .Z(
        P2_U3523) );
  MUX2_X1 U10836 ( .A(P2_REG1_REG_0__SCAN_IN), .B(n9559), .S(n10426), .Z(
        P2_U3520) );
  MUX2_X1 U10837 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n9560), .S(n10418), .Z(
        P2_U3519) );
  MUX2_X1 U10838 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n9561), .S(n10418), .Z(
        P2_U3518) );
  MUX2_X1 U10839 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n9562), .S(n10418), .Z(
        P2_U3517) );
  MUX2_X1 U10840 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n9564), .S(n10418), .Z(
        P2_U3515) );
  MUX2_X1 U10841 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n9565), .S(n10418), .Z(
        P2_U3514) );
  MUX2_X1 U10842 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n9566), .S(n10418), .Z(
        P2_U3513) );
  MUX2_X1 U10843 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n9567), .S(n10418), .Z(
        P2_U3512) );
  MUX2_X1 U10844 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n9568), .S(n10418), .Z(
        P2_U3511) );
  MUX2_X1 U10845 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n9569), .S(n10418), .Z(
        P2_U3510) );
  MUX2_X1 U10846 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n9570), .S(n10418), .Z(
        P2_U3509) );
  MUX2_X1 U10847 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n9571), .S(n10418), .Z(
        P2_U3508) );
  MUX2_X1 U10848 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n9572), .S(n10418), .Z(
        P2_U3507) );
  MUX2_X1 U10849 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n9573), .S(n10418), .Z(
        P2_U3505) );
  MUX2_X1 U10850 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n9574), .S(n10418), .Z(
        P2_U3502) );
  MUX2_X1 U10851 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n9575), .S(n10418), .Z(
        P2_U3499) );
  MUX2_X1 U10852 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n9576), .S(n10418), .Z(
        P2_U3496) );
  MUX2_X1 U10853 ( .A(n9577), .B(P2_REG0_REG_14__SCAN_IN), .S(n10416), .Z(
        P2_U3493) );
  MUX2_X1 U10854 ( .A(P2_REG0_REG_13__SCAN_IN), .B(n9578), .S(n10418), .Z(
        P2_U3490) );
  MUX2_X1 U10855 ( .A(n9579), .B(P2_REG0_REG_12__SCAN_IN), .S(n10416), .Z(
        P2_U3487) );
  MUX2_X1 U10856 ( .A(P2_REG0_REG_11__SCAN_IN), .B(n9580), .S(n10418), .Z(
        P2_U3484) );
  MUX2_X1 U10857 ( .A(P2_REG0_REG_10__SCAN_IN), .B(n9581), .S(n10418), .Z(
        P2_U3481) );
  MUX2_X1 U10858 ( .A(P2_REG0_REG_8__SCAN_IN), .B(n9582), .S(n10418), .Z(
        P2_U3475) );
  INV_X1 U10859 ( .A(n9583), .ZN(n10241) );
  NAND3_X1 U10860 ( .A1(n9585), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .ZN(n9588) );
  OAI22_X1 U10861 ( .A1(n9584), .A2(n9588), .B1(n9587), .B2(n9586), .ZN(n9589)
         );
  INV_X1 U10862 ( .A(n9589), .ZN(n9590) );
  OAI21_X1 U10863 ( .B1(n10241), .B2(n9591), .A(n9590), .ZN(P2_U3327) );
  INV_X1 U10864 ( .A(n9592), .ZN(n9593) );
  MUX2_X1 U10865 ( .A(n9593), .B(n10367), .S(P2_STATE_REG_SCAN_IN), .Z(
        P2_U3358) );
  NOR2_X1 U10866 ( .A1(n9596), .A2(n9758), .ZN(n9600) );
  AOI22_X1 U10867 ( .A1(n9597), .A2(n9763), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3084), .ZN(n9598) );
  OAI21_X1 U10868 ( .B1(n9655), .B2(n9743), .A(n9598), .ZN(n9599) );
  AOI211_X1 U10869 ( .C1(n10107), .C2(n9734), .A(n9600), .B(n9599), .ZN(n9601)
         );
  INV_X1 U10870 ( .A(n9700), .ZN(n9602) );
  AOI21_X1 U10871 ( .B1(n4379), .B2(n9602), .A(n9699), .ZN(n9604) );
  NOR2_X1 U10872 ( .A1(n9604), .A2(n9603), .ZN(n9660) );
  INV_X1 U10873 ( .A(n9604), .ZN(n9606) );
  NOR2_X1 U10874 ( .A1(n9660), .A2(n9662), .ZN(n9608) );
  XNOR2_X1 U10875 ( .A(n9608), .B(n9607), .ZN(n9615) );
  AOI21_X1 U10876 ( .B1(n9755), .B2(n10058), .A(n9609), .ZN(n9611) );
  NAND2_X1 U10877 ( .A1(n9763), .A2(n10065), .ZN(n9610) );
  OAI211_X1 U10878 ( .C1(n9612), .C2(n9758), .A(n9611), .B(n9610), .ZN(n9613)
         );
  AOI21_X1 U10879 ( .B1(n10174), .B2(n9734), .A(n9613), .ZN(n9614) );
  OAI21_X1 U10880 ( .B1(n9615), .B2(n9737), .A(n9614), .ZN(P1_U3213) );
  NAND2_X1 U10881 ( .A1(n9617), .A2(n9616), .ZN(n9618) );
  XOR2_X1 U10882 ( .A(n9619), .B(n9618), .Z(n9624) );
  AOI22_X1 U10883 ( .A1(n9918), .A2(n9755), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3084), .ZN(n9621) );
  NAND2_X1 U10884 ( .A1(n9908), .A2(n9763), .ZN(n9620) );
  OAI211_X1 U10885 ( .C1(n9652), .C2(n9758), .A(n9621), .B(n9620), .ZN(n9622)
         );
  AOI21_X1 U10886 ( .B1(n10126), .B2(n9734), .A(n9622), .ZN(n9623) );
  OAI21_X1 U10887 ( .B1(n9624), .B2(n9737), .A(n9623), .ZN(P1_U3214) );
  INV_X1 U10888 ( .A(n9727), .ZN(n9627) );
  NAND2_X1 U10889 ( .A1(n9625), .A2(n9626), .ZN(n9725) );
  NOR2_X1 U10890 ( .A1(n9625), .A2(n9626), .ZN(n9724) );
  AOI21_X1 U10891 ( .B1(n9627), .B2(n9725), .A(n9724), .ZN(n9631) );
  XNOR2_X1 U10892 ( .A(n9629), .B(n9628), .ZN(n9630) );
  XNOR2_X1 U10893 ( .A(n9631), .B(n9630), .ZN(n9637) );
  OAI21_X1 U10894 ( .B1(n9953), .B2(n9758), .A(n9632), .ZN(n9633) );
  AOI21_X1 U10895 ( .B1(n9755), .B2(n10004), .A(n9633), .ZN(n9634) );
  OAI21_X1 U10896 ( .B1(n9732), .B2(n9972), .A(n9634), .ZN(n9635) );
  AOI21_X1 U10897 ( .B1(n10148), .B2(n9734), .A(n9635), .ZN(n9636) );
  OAI21_X1 U10898 ( .B1(n9637), .B2(n9737), .A(n9636), .ZN(P1_U3217) );
  NAND2_X1 U10899 ( .A1(n9692), .A2(n9693), .ZN(n9639) );
  NAND2_X1 U10900 ( .A1(n9639), .A2(n9638), .ZN(n9640) );
  XOR2_X1 U10901 ( .A(n9641), .B(n9640), .Z(n9647) );
  OAI22_X1 U10902 ( .A1(n9951), .A2(n9758), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9642), .ZN(n9643) );
  AOI21_X1 U10903 ( .B1(n9755), .B2(n9979), .A(n9643), .ZN(n9644) );
  OAI21_X1 U10904 ( .B1(n9732), .B2(n9943), .A(n9644), .ZN(n9645) );
  AOI21_X1 U10905 ( .B1(n10140), .B2(n9734), .A(n9645), .ZN(n9646) );
  OAI21_X1 U10906 ( .B1(n9647), .B2(n9737), .A(n9646), .ZN(P1_U3221) );
  XOR2_X1 U10907 ( .A(n9649), .B(n9648), .Z(n9658) );
  INV_X1 U10908 ( .A(n9650), .ZN(n9883) );
  OAI22_X1 U10909 ( .A1(n9652), .A2(n9743), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9651), .ZN(n9653) );
  AOI21_X1 U10910 ( .B1(n9883), .B2(n9763), .A(n9653), .ZN(n9654) );
  OAI21_X1 U10911 ( .B1(n9655), .B2(n9758), .A(n9654), .ZN(n9656) );
  AOI21_X1 U10912 ( .B1(n10116), .B2(n9734), .A(n9656), .ZN(n9657) );
  OAI21_X1 U10913 ( .B1(n9658), .B2(n9737), .A(n9657), .ZN(P1_U3223) );
  NOR2_X1 U10914 ( .A1(n9660), .A2(n9659), .ZN(n9663) );
  NOR3_X1 U10915 ( .A1(n9663), .A2(n9662), .A3(n9661), .ZN(n9750) );
  OAI21_X1 U10916 ( .B1(n9663), .B2(n9662), .A(n9661), .ZN(n9751) );
  OAI21_X1 U10917 ( .B1(n9750), .B2(n9753), .A(n9751), .ZN(n9667) );
  XNOR2_X1 U10918 ( .A(n9665), .B(n9664), .ZN(n9666) );
  XNOR2_X1 U10919 ( .A(n9667), .B(n9666), .ZN(n9673) );
  NAND2_X1 U10920 ( .A1(n9755), .A2(n10056), .ZN(n9668) );
  NAND2_X1 U10921 ( .A1(P1_U3084), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9815) );
  OAI211_X1 U10922 ( .C1(n9669), .C2(n9758), .A(n9668), .B(n9815), .ZN(n9670)
         );
  AOI21_X1 U10923 ( .B1(n10023), .B2(n9763), .A(n9670), .ZN(n9672) );
  NAND2_X1 U10924 ( .A1(n10164), .A2(n9734), .ZN(n9671) );
  OAI211_X1 U10925 ( .C1(n9673), .C2(n9737), .A(n9672), .B(n9671), .ZN(
        P1_U3224) );
  OR2_X1 U10926 ( .A1(n5006), .A2(n9674), .ZN(n9675) );
  XOR2_X1 U10927 ( .A(n9676), .B(n9675), .Z(n9681) );
  NAND2_X1 U10928 ( .A1(n9703), .A2(n10004), .ZN(n9677) );
  NAND2_X1 U10929 ( .A1(P1_U3084), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9822) );
  OAI211_X1 U10930 ( .C1(n9759), .C2(n9743), .A(n9677), .B(n9822), .ZN(n9679)
         );
  NOR2_X1 U10931 ( .A1(n10011), .A2(n9760), .ZN(n9678) );
  AOI211_X1 U10932 ( .C1(n10009), .C2(n9763), .A(n9679), .B(n9678), .ZN(n9680)
         );
  OAI21_X1 U10933 ( .B1(n9681), .B2(n9737), .A(n9680), .ZN(P1_U3226) );
  INV_X1 U10934 ( .A(n9682), .ZN(n9683) );
  AOI21_X1 U10935 ( .B1(n9685), .B2(n9684), .A(n9683), .ZN(n9691) );
  AOI22_X1 U10936 ( .A1(n9926), .A2(n9755), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3084), .ZN(n9688) );
  INV_X1 U10937 ( .A(n9686), .ZN(n9895) );
  NAND2_X1 U10938 ( .A1(n9895), .A2(n9763), .ZN(n9687) );
  OAI211_X1 U10939 ( .C1(n9744), .C2(n9758), .A(n9688), .B(n9687), .ZN(n9689)
         );
  AOI21_X1 U10940 ( .B1(n10121), .B2(n9734), .A(n9689), .ZN(n9690) );
  OAI21_X1 U10941 ( .B1(n9691), .B2(n9765), .A(n9690), .ZN(P1_U3227) );
  XOR2_X1 U10942 ( .A(n9693), .B(n9692), .Z(n9698) );
  AOI22_X1 U10943 ( .A1(n9959), .A2(n9703), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3084), .ZN(n9695) );
  NAND2_X1 U10944 ( .A1(n9755), .A2(n9988), .ZN(n9694) );
  OAI211_X1 U10945 ( .C1(n9732), .C2(n9964), .A(n9695), .B(n9694), .ZN(n9696)
         );
  AOI21_X1 U10946 ( .B1(n10144), .B2(n9734), .A(n9696), .ZN(n9697) );
  OAI21_X1 U10947 ( .B1(n9698), .B2(n9765), .A(n9697), .ZN(P1_U3231) );
  NOR2_X1 U10948 ( .A1(n9700), .A2(n9699), .ZN(n9701) );
  XNOR2_X1 U10949 ( .A(n9702), .B(n9701), .ZN(n9712) );
  NAND2_X1 U10950 ( .A1(n9703), .A2(n10037), .ZN(n9705) );
  OAI211_X1 U10951 ( .C1(n9706), .C2(n9743), .A(n9705), .B(n9704), .ZN(n9709)
         );
  NOR2_X1 U10952 ( .A1(n9707), .A2(n9760), .ZN(n9708) );
  AOI211_X1 U10953 ( .C1(n9710), .C2(n9763), .A(n9709), .B(n9708), .ZN(n9711)
         );
  OAI21_X1 U10954 ( .B1(n9712), .B2(n9765), .A(n9711), .ZN(P1_U3232) );
  NAND2_X1 U10955 ( .A1(n9714), .A2(n9713), .ZN(n9715) );
  XOR2_X1 U10956 ( .A(n9716), .B(n9715), .Z(n9723) );
  AOI22_X1 U10957 ( .A1(n9959), .A2(n9755), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3084), .ZN(n9719) );
  INV_X1 U10958 ( .A(n9717), .ZN(n9929) );
  NAND2_X1 U10959 ( .A1(n9763), .A2(n9929), .ZN(n9718) );
  OAI211_X1 U10960 ( .C1(n9720), .C2(n9758), .A(n9719), .B(n9718), .ZN(n9721)
         );
  AOI21_X1 U10961 ( .B1(n9934), .B2(n9734), .A(n9721), .ZN(n9722) );
  OAI21_X1 U10962 ( .B1(n9723), .B2(n9765), .A(n9722), .ZN(P1_U3233) );
  INV_X1 U10963 ( .A(n9724), .ZN(n9726) );
  NAND2_X1 U10964 ( .A1(n9726), .A2(n9725), .ZN(n9728) );
  XNOR2_X1 U10965 ( .A(n9728), .B(n9727), .ZN(n9736) );
  NAND2_X1 U10966 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n10295)
         );
  OAI21_X1 U10967 ( .B1(n9758), .B2(n9729), .A(n10295), .ZN(n9730) );
  AOI21_X1 U10968 ( .B1(n9755), .B2(n10019), .A(n9730), .ZN(n9731) );
  OAI21_X1 U10969 ( .B1(n9732), .B2(n9993), .A(n9731), .ZN(n9733) );
  AOI21_X1 U10970 ( .B1(n10154), .B2(n9734), .A(n9733), .ZN(n9735) );
  OAI21_X1 U10971 ( .B1(n9736), .B2(n9765), .A(n9735), .ZN(P1_U3236) );
  AOI21_X1 U10972 ( .B1(n9739), .B2(n9738), .A(n9737), .ZN(n9741) );
  NAND2_X1 U10973 ( .A1(n9741), .A2(n9740), .ZN(n9749) );
  OAI22_X1 U10974 ( .A1(n9744), .A2(n9743), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9742), .ZN(n9747) );
  NOR2_X1 U10975 ( .A1(n9745), .A2(n9758), .ZN(n9746) );
  AOI211_X1 U10976 ( .C1(n9866), .C2(n9763), .A(n9747), .B(n9746), .ZN(n9748)
         );
  OAI211_X1 U10977 ( .C1(n9868), .C2(n9760), .A(n9749), .B(n9748), .ZN(
        P1_U3238) );
  INV_X1 U10978 ( .A(n9750), .ZN(n9752) );
  NAND2_X1 U10979 ( .A1(n9752), .A2(n9751), .ZN(n9754) );
  XNOR2_X1 U10980 ( .A(n9754), .B(n9753), .ZN(n9766) );
  NAND2_X1 U10981 ( .A1(n9755), .A2(n10037), .ZN(n9757) );
  NAND2_X1 U10982 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9801) );
  OAI211_X1 U10983 ( .C1(n9759), .C2(n9758), .A(n9757), .B(n9801), .ZN(n9762)
         );
  NOR2_X1 U10984 ( .A1(n10048), .A2(n9760), .ZN(n9761) );
  AOI211_X1 U10985 ( .C1(n10045), .C2(n9763), .A(n9762), .B(n9761), .ZN(n9764)
         );
  OAI21_X1 U10986 ( .B1(n9766), .B2(n9765), .A(n9764), .ZN(P1_U3239) );
  MUX2_X1 U10987 ( .A(n9767), .B(P1_DATAO_REG_30__SCAN_IN), .S(n9778), .Z(
        P1_U3585) );
  INV_X1 U10988 ( .A(n9768), .ZN(n9856) );
  MUX2_X1 U10989 ( .A(n9856), .B(P1_DATAO_REG_29__SCAN_IN), .S(n9778), .Z(
        P1_U3584) );
  MUX2_X1 U10990 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9769), .S(P1_U4006), .Z(
        P1_U3583) );
  MUX2_X1 U10991 ( .A(n9873), .B(P1_DATAO_REG_27__SCAN_IN), .S(n9778), .Z(
        P1_U3582) );
  MUX2_X1 U10992 ( .A(n9888), .B(P1_DATAO_REG_26__SCAN_IN), .S(n9778), .Z(
        P1_U3581) );
  MUX2_X1 U10993 ( .A(n9900), .B(P1_DATAO_REG_25__SCAN_IN), .S(n9778), .Z(
        P1_U3580) );
  MUX2_X1 U10994 ( .A(n9919), .B(P1_DATAO_REG_24__SCAN_IN), .S(n9778), .Z(
        P1_U3579) );
  MUX2_X1 U10995 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9926), .S(P1_U4006), .Z(
        P1_U3578) );
  MUX2_X1 U10996 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9918), .S(P1_U4006), .Z(
        P1_U3577) );
  MUX2_X1 U10997 ( .A(n9959), .B(P1_DATAO_REG_21__SCAN_IN), .S(n9778), .Z(
        P1_U3576) );
  MUX2_X1 U10998 ( .A(n9979), .B(P1_DATAO_REG_20__SCAN_IN), .S(n9778), .Z(
        P1_U3575) );
  MUX2_X1 U10999 ( .A(n9988), .B(P1_DATAO_REG_19__SCAN_IN), .S(n9778), .Z(
        P1_U3574) );
  MUX2_X1 U11000 ( .A(n10004), .B(P1_DATAO_REG_18__SCAN_IN), .S(n9778), .Z(
        P1_U3573) );
  MUX2_X1 U11001 ( .A(n10019), .B(P1_DATAO_REG_17__SCAN_IN), .S(n9778), .Z(
        P1_U3572) );
  MUX2_X1 U11002 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n10038), .S(P1_U4006), .Z(
        P1_U3571) );
  MUX2_X1 U11003 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n10056), .S(P1_U4006), .Z(
        P1_U3570) );
  MUX2_X1 U11004 ( .A(n10037), .B(P1_DATAO_REG_14__SCAN_IN), .S(n9778), .Z(
        P1_U3569) );
  MUX2_X1 U11005 ( .A(n10058), .B(P1_DATAO_REG_13__SCAN_IN), .S(n9778), .Z(
        P1_U3568) );
  MUX2_X1 U11006 ( .A(n9770), .B(P1_DATAO_REG_12__SCAN_IN), .S(n9778), .Z(
        P1_U3567) );
  MUX2_X1 U11007 ( .A(n9771), .B(P1_DATAO_REG_11__SCAN_IN), .S(n9778), .Z(
        P1_U3566) );
  MUX2_X1 U11008 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9772), .S(P1_U4006), .Z(
        P1_U3565) );
  MUX2_X1 U11009 ( .A(n9773), .B(P1_DATAO_REG_9__SCAN_IN), .S(n9778), .Z(
        P1_U3564) );
  MUX2_X1 U11010 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9774), .S(P1_U4006), .Z(
        P1_U3563) );
  MUX2_X1 U11011 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9775), .S(P1_U4006), .Z(
        P1_U3562) );
  MUX2_X1 U11012 ( .A(n9776), .B(P1_DATAO_REG_6__SCAN_IN), .S(n9778), .Z(
        P1_U3561) );
  MUX2_X1 U11013 ( .A(n9777), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9778), .Z(
        P1_U3559) );
  MUX2_X1 U11014 ( .A(n9779), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9778), .Z(
        P1_U3558) );
  MUX2_X1 U11015 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n6580), .S(P1_U4006), .Z(
        P1_U3557) );
  MUX2_X1 U11016 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n9780), .S(P1_U4006), .Z(
        P1_U3556) );
  INV_X1 U11017 ( .A(n9781), .ZN(n9795) );
  INV_X1 U11018 ( .A(n9782), .ZN(n9788) );
  AOI21_X1 U11019 ( .B1(n9785), .B2(n9784), .A(n9783), .ZN(n9786) );
  NOR2_X1 U11020 ( .A1(n9823), .A2(n9786), .ZN(n9787) );
  AOI211_X1 U11021 ( .C1(n10294), .C2(n9789), .A(n9788), .B(n9787), .ZN(n9794)
         );
  OAI21_X1 U11022 ( .B1(n9791), .B2(n4502), .A(n9790), .ZN(n9792) );
  AOI22_X1 U11023 ( .A1(n10301), .A2(P1_ADDR_REG_4__SCAN_IN), .B1(n9792), .B2(
        n10292), .ZN(n9793) );
  NAND3_X1 U11024 ( .A1(n9795), .A2(n9794), .A3(n9793), .ZN(P1_U3245) );
  INV_X1 U11025 ( .A(n9796), .ZN(n9799) );
  INV_X1 U11026 ( .A(n9797), .ZN(n9798) );
  OAI211_X1 U11027 ( .C1(P1_REG1_REG_15__SCAN_IN), .C2(n9799), .A(n10302), .B(
        n9798), .ZN(n9800) );
  OAI211_X1 U11028 ( .C1(n9818), .C2(n9802), .A(n9801), .B(n9800), .ZN(n9807)
         );
  AOI211_X1 U11029 ( .C1(n9805), .C2(n9804), .A(n9803), .B(n9830), .ZN(n9806)
         );
  AOI211_X1 U11030 ( .C1(n10301), .C2(P1_ADDR_REG_15__SCAN_IN), .A(n9807), .B(
        n9806), .ZN(n9808) );
  INV_X1 U11031 ( .A(n9808), .ZN(P1_U3256) );
  AOI211_X1 U11032 ( .C1(n9811), .C2(n9810), .A(n9809), .B(n9830), .ZN(n9821)
         );
  AOI211_X1 U11033 ( .C1(n9814), .C2(n9813), .A(n9812), .B(n9823), .ZN(n9820)
         );
  NAND2_X1 U11034 ( .A1(n10301), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n9816) );
  OAI211_X1 U11035 ( .C1(n9818), .C2(n9817), .A(n9816), .B(n9815), .ZN(n9819)
         );
  OR3_X1 U11036 ( .A1(n9821), .A2(n9820), .A3(n9819), .ZN(P1_U3257) );
  INV_X1 U11037 ( .A(n9822), .ZN(n9828) );
  AOI211_X1 U11038 ( .C1(n9826), .C2(n9825), .A(n9824), .B(n9823), .ZN(n9827)
         );
  AOI211_X1 U11039 ( .C1(n10294), .C2(n9829), .A(n9828), .B(n9827), .ZN(n9836)
         );
  AOI211_X1 U11040 ( .C1(n9833), .C2(n9832), .A(n9831), .B(n9830), .ZN(n9834)
         );
  AOI21_X1 U11041 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(n10301), .A(n9834), .ZN(
        n9835) );
  NAND2_X1 U11042 ( .A1(n9836), .A2(n9835), .ZN(P1_U3258) );
  XNOR2_X2 U11043 ( .A(n10079), .B(n10082), .ZN(n10081) );
  NAND2_X1 U11044 ( .A1(n9838), .A2(n9837), .ZN(n10084) );
  NOR2_X1 U11045 ( .A1(n10317), .A2(n10084), .ZN(n9843) );
  AOI211_X1 U11046 ( .C1(n10317), .C2(P1_REG2_REG_31__SCAN_IN), .A(n9843), .B(
        n9839), .ZN(n9840) );
  OAI21_X1 U11047 ( .B1(n10081), .B2(n9936), .A(n9840), .ZN(P1_U3261) );
  INV_X1 U11048 ( .A(n9841), .ZN(n9842) );
  NAND2_X1 U11049 ( .A1(n9842), .A2(n6437), .ZN(n10083) );
  NAND3_X1 U11050 ( .A1(n10083), .A2(n10052), .A3(n10082), .ZN(n9845) );
  AOI21_X1 U11051 ( .B1(n10317), .B2(P1_REG2_REG_30__SCAN_IN), .A(n9843), .ZN(
        n9844) );
  OAI211_X1 U11052 ( .C1(n10086), .C2(n10047), .A(n9845), .B(n9844), .ZN(
        P1_U3262) );
  OAI22_X1 U11053 ( .A1(n9847), .A2(n9992), .B1(n9846), .B2(n10315), .ZN(n9848) );
  AOI21_X1 U11054 ( .B1(n10102), .B2(n10064), .A(n9848), .ZN(n9853) );
  AOI21_X1 U11055 ( .B1(n9849), .B2(n10102), .A(n10334), .ZN(n9851) );
  NAND2_X1 U11056 ( .A1(n10101), .A2(n10077), .ZN(n9852) );
  OAI211_X1 U11057 ( .C1(n10105), .C2(n10074), .A(n9853), .B(n9852), .ZN(n9861) );
  NOR2_X1 U11058 ( .A1(n10104), .A2(n10317), .ZN(n9860) );
  OR2_X1 U11059 ( .A1(n9861), .A2(n9860), .ZN(P1_U3263) );
  XOR2_X1 U11060 ( .A(n9871), .B(n9863), .Z(n10115) );
  INV_X1 U11061 ( .A(n9882), .ZN(n9865) );
  AOI21_X1 U11062 ( .B1(n10111), .B2(n9865), .A(n9864), .ZN(n10112) );
  AOI22_X1 U11063 ( .A1(n9866), .A2(n10307), .B1(P1_REG2_REG_26__SCAN_IN), 
        .B2(n10317), .ZN(n9867) );
  OAI21_X1 U11064 ( .B1(n9868), .B2(n10047), .A(n9867), .ZN(n9879) );
  NAND2_X1 U11065 ( .A1(n9870), .A2(n9869), .ZN(n9872) );
  XNOR2_X1 U11066 ( .A(n9872), .B(n9871), .ZN(n9877) );
  OAI21_X1 U11067 ( .B1(n10115), .B2(n10074), .A(n9880), .ZN(P1_U3265) );
  XOR2_X1 U11068 ( .A(n9886), .B(n9881), .Z(n10120) );
  AOI21_X1 U11069 ( .B1(n10116), .B2(n9894), .A(n9882), .ZN(n10117) );
  AOI22_X1 U11070 ( .A1(n9883), .A2(n10307), .B1(P1_REG2_REG_25__SCAN_IN), 
        .B2(n10317), .ZN(n9884) );
  OAI21_X1 U11071 ( .B1(n9885), .B2(n10047), .A(n9884), .ZN(n9890) );
  NOR2_X1 U11072 ( .A1(n10119), .A2(n10317), .ZN(n9889) );
  AOI211_X1 U11073 ( .C1(n10117), .C2(n10052), .A(n9890), .B(n9889), .ZN(n9891) );
  OAI21_X1 U11074 ( .B1(n10120), .B2(n10074), .A(n9891), .ZN(P1_U3266) );
  XOR2_X1 U11075 ( .A(n9899), .B(n9893), .Z(n10125) );
  AOI21_X1 U11076 ( .B1(n10121), .B2(n4531), .A(n5055), .ZN(n10122) );
  INV_X1 U11077 ( .A(n10121), .ZN(n9897) );
  AOI22_X1 U11078 ( .A1(n9895), .A2(n10307), .B1(P1_REG2_REG_24__SCAN_IN), 
        .B2(n10317), .ZN(n9896) );
  OAI21_X1 U11079 ( .B1(n9897), .B2(n10047), .A(n9896), .ZN(n9903) );
  XOR2_X1 U11080 ( .A(n9899), .B(n9898), .Z(n9901) );
  AOI222_X1 U11081 ( .A1(n10099), .A2(n9901), .B1(n9926), .B2(n10057), .C1(
        n9900), .C2(n10055), .ZN(n10124) );
  NOR2_X1 U11082 ( .A1(n10124), .A2(n10317), .ZN(n9902) );
  AOI211_X1 U11083 ( .C1(n10122), .C2(n10052), .A(n9903), .B(n9902), .ZN(n9904) );
  OAI21_X1 U11084 ( .B1(n10125), .B2(n10074), .A(n9904), .ZN(P1_U3267) );
  XNOR2_X1 U11085 ( .A(n9905), .B(n9916), .ZN(n10130) );
  INV_X1 U11086 ( .A(n9933), .ZN(n9907) );
  AOI21_X1 U11087 ( .B1(n10126), .B2(n9907), .A(n5049), .ZN(n10127) );
  AOI22_X1 U11088 ( .A1(n9908), .A2(n10307), .B1(n10317), .B2(
        P1_REG2_REG_23__SCAN_IN), .ZN(n9909) );
  OAI21_X1 U11089 ( .B1(n9910), .B2(n10047), .A(n9909), .ZN(n9923) );
  INV_X1 U11090 ( .A(n9911), .ZN(n9913) );
  NAND2_X1 U11091 ( .A1(n9913), .A2(n9912), .ZN(n9925) );
  AOI21_X1 U11092 ( .B1(n9925), .B2(n4425), .A(n9914), .ZN(n9917) );
  OAI211_X1 U11093 ( .C1(n9917), .C2(n9916), .A(n10099), .B(n9915), .ZN(n9921)
         );
  AOI22_X1 U11094 ( .A1(n9919), .A2(n10055), .B1(n10057), .B2(n9918), .ZN(
        n9920) );
  AND2_X1 U11095 ( .A1(n9921), .A2(n9920), .ZN(n10129) );
  NOR2_X1 U11096 ( .A1(n10129), .A2(n10317), .ZN(n9922) );
  AOI211_X1 U11097 ( .C1(n10127), .C2(n10052), .A(n9923), .B(n9922), .ZN(n9924) );
  OAI21_X1 U11098 ( .B1(n10130), .B2(n10074), .A(n9924), .ZN(P1_U3268) );
  XNOR2_X1 U11099 ( .A(n9925), .B(n4425), .ZN(n9927) );
  AOI222_X1 U11100 ( .A1(n10099), .A2(n9927), .B1(n9926), .B2(n10055), .C1(
        n9959), .C2(n10057), .ZN(n10136) );
  INV_X1 U11101 ( .A(n10136), .ZN(n9928) );
  AOI21_X1 U11102 ( .B1(n9929), .B2(n10307), .A(n9928), .ZN(n9940) );
  XNOR2_X1 U11103 ( .A(n9930), .B(n4425), .ZN(n10135) );
  NOR2_X1 U11104 ( .A1(n9931), .A2(n10131), .ZN(n9932) );
  OR2_X1 U11105 ( .A1(n9933), .A2(n9932), .ZN(n10132) );
  AOI22_X1 U11106 ( .A1(n9934), .A2(n10064), .B1(P1_REG2_REG_22__SCAN_IN), 
        .B2(n10317), .ZN(n9935) );
  OAI21_X1 U11107 ( .B1(n10132), .B2(n9936), .A(n9935), .ZN(n9937) );
  AOI21_X1 U11108 ( .B1(n10135), .B2(n9938), .A(n9937), .ZN(n9939) );
  OAI21_X1 U11109 ( .B1(n10317), .B2(n9940), .A(n9939), .ZN(P1_U3269) );
  XNOR2_X1 U11110 ( .A(n9941), .B(n9947), .ZN(n10142) );
  AOI211_X1 U11111 ( .C1(n10140), .C2(n5103), .A(n10334), .B(n9931), .ZN(
        n10139) );
  NOR2_X1 U11112 ( .A1(n9942), .A2(n10047), .ZN(n9946) );
  OAI22_X1 U11113 ( .A1(n10315), .A2(n9944), .B1(n9943), .B2(n9992), .ZN(n9945) );
  AOI211_X1 U11114 ( .C1(n10139), .C2(n10077), .A(n9946), .B(n9945), .ZN(n9956) );
  AOI21_X1 U11115 ( .B1(n9948), .B2(n9947), .A(n9911), .ZN(n9949) );
  OAI222_X1 U11116 ( .A1(n9954), .A2(n9953), .B1(n9952), .B2(n9951), .C1(n9950), .C2(n9949), .ZN(n10138) );
  NAND2_X1 U11117 ( .A1(n10138), .A2(n10315), .ZN(n9955) );
  OAI211_X1 U11118 ( .C1(n10142), .C2(n10074), .A(n9956), .B(n9955), .ZN(
        P1_U3270) );
  XNOR2_X1 U11119 ( .A(n4385), .B(n9958), .ZN(n10147) );
  AOI22_X1 U11120 ( .A1(n10144), .A2(n10064), .B1(P1_REG2_REG_20__SCAN_IN), 
        .B2(n10317), .ZN(n9967) );
  XOR2_X1 U11121 ( .A(n9958), .B(n9957), .Z(n9960) );
  AOI222_X1 U11122 ( .A1(n10099), .A2(n9960), .B1(n9988), .B2(n10057), .C1(
        n9959), .C2(n10055), .ZN(n10146) );
  AOI21_X1 U11123 ( .B1(n9969), .B2(n10144), .A(n10334), .ZN(n9961) );
  AND2_X1 U11124 ( .A1(n9961), .A2(n5103), .ZN(n10143) );
  NAND2_X1 U11125 ( .A1(n10143), .A2(n9962), .ZN(n9963) );
  OAI211_X1 U11126 ( .C1(n9992), .C2(n9964), .A(n10146), .B(n9963), .ZN(n9965)
         );
  NAND2_X1 U11127 ( .A1(n9965), .A2(n10315), .ZN(n9966) );
  OAI211_X1 U11128 ( .C1(n10147), .C2(n10074), .A(n9967), .B(n9966), .ZN(
        P1_U3271) );
  XNOR2_X1 U11129 ( .A(n9968), .B(n9977), .ZN(n10152) );
  INV_X1 U11130 ( .A(n9998), .ZN(n9971) );
  INV_X1 U11131 ( .A(n9969), .ZN(n9970) );
  AOI21_X1 U11132 ( .B1(n10148), .B2(n9971), .A(n9970), .ZN(n10149) );
  INV_X1 U11133 ( .A(n9972), .ZN(n9973) );
  AOI22_X1 U11134 ( .A1(n10317), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9973), 
        .B2(n10307), .ZN(n9974) );
  OAI21_X1 U11135 ( .B1(n9975), .B2(n10047), .A(n9974), .ZN(n9982) );
  OAI21_X1 U11136 ( .B1(n9978), .B2(n9977), .A(n9976), .ZN(n9980) );
  AOI222_X1 U11137 ( .A1(n10099), .A2(n9980), .B1(n10004), .B2(n10057), .C1(
        n9979), .C2(n10055), .ZN(n10151) );
  NOR2_X1 U11138 ( .A1(n10151), .A2(n10317), .ZN(n9981) );
  AOI211_X1 U11139 ( .C1(n10149), .C2(n10052), .A(n9982), .B(n9981), .ZN(n9983) );
  OAI21_X1 U11140 ( .B1(n10074), .B2(n10152), .A(n9983), .ZN(P1_U3272) );
  INV_X1 U11141 ( .A(n9984), .ZN(n9986) );
  OAI21_X1 U11142 ( .B1(n10003), .B2(n9986), .A(n9985), .ZN(n9987) );
  XNOR2_X1 U11143 ( .A(n9987), .B(n9990), .ZN(n9989) );
  AOI222_X1 U11144 ( .A1(n10099), .A2(n9989), .B1(n10019), .B2(n10057), .C1(
        n9988), .C2(n10055), .ZN(n10156) );
  XNOR2_X1 U11145 ( .A(n9991), .B(n9990), .ZN(n10157) );
  INV_X1 U11146 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9994) );
  OAI22_X1 U11147 ( .A1(n10315), .A2(n9994), .B1(n9993), .B2(n9992), .ZN(n9995) );
  AOI21_X1 U11148 ( .B1(n10154), .B2(n10064), .A(n9995), .ZN(n10000) );
  NAND2_X1 U11149 ( .A1(n10007), .A2(n10154), .ZN(n9996) );
  NAND2_X1 U11150 ( .A1(n9996), .A2(n10341), .ZN(n9997) );
  NOR2_X1 U11151 ( .A1(n9998), .A2(n9997), .ZN(n10153) );
  NAND2_X1 U11152 ( .A1(n10153), .A2(n10077), .ZN(n9999) );
  OAI211_X1 U11153 ( .C1(n10157), .C2(n10074), .A(n10000), .B(n9999), .ZN(
        n10001) );
  INV_X1 U11154 ( .A(n10001), .ZN(n10002) );
  OAI21_X1 U11155 ( .B1(n10317), .B2(n10156), .A(n10002), .ZN(P1_U3273) );
  XOR2_X1 U11156 ( .A(n10003), .B(n10013), .Z(n10005) );
  AOI222_X1 U11157 ( .A1(n10099), .A2(n10005), .B1(n10038), .B2(n10057), .C1(
        n10004), .C2(n10055), .ZN(n10161) );
  NAND2_X1 U11158 ( .A1(n10062), .A2(n10006), .ZN(n10021) );
  INV_X1 U11159 ( .A(n10007), .ZN(n10008) );
  AOI21_X1 U11160 ( .B1(n10158), .B2(n10021), .A(n10008), .ZN(n10159) );
  AOI22_X1 U11161 ( .A1(n10317), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n10009), 
        .B2(n10307), .ZN(n10010) );
  OAI21_X1 U11162 ( .B1(n10011), .B2(n10047), .A(n10010), .ZN(n10015) );
  XOR2_X1 U11163 ( .A(n10013), .B(n10012), .Z(n10162) );
  NOR2_X1 U11164 ( .A1(n10162), .A2(n10074), .ZN(n10014) );
  AOI211_X1 U11165 ( .C1(n10159), .C2(n10052), .A(n10015), .B(n10014), .ZN(
        n10016) );
  OAI21_X1 U11166 ( .B1(n10317), .B2(n10161), .A(n10016), .ZN(P1_U3274) );
  XNOR2_X1 U11167 ( .A(n10018), .B(n10017), .ZN(n10020) );
  AOI222_X1 U11168 ( .A1(n10099), .A2(n10020), .B1(n10056), .B2(n10057), .C1(
        n10019), .C2(n10055), .ZN(n10166) );
  NAND2_X1 U11169 ( .A1(n10062), .A2(n10048), .ZN(n10044) );
  AOI21_X1 U11170 ( .B1(n10044), .B2(n10164), .A(n10334), .ZN(n10022) );
  AND2_X1 U11171 ( .A1(n10022), .A2(n10021), .ZN(n10163) );
  INV_X1 U11172 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n10026) );
  NAND2_X1 U11173 ( .A1(n10164), .A2(n10064), .ZN(n10025) );
  NAND2_X1 U11174 ( .A1(n10307), .A2(n10023), .ZN(n10024) );
  OAI211_X1 U11175 ( .C1(n10315), .C2(n10026), .A(n10025), .B(n10024), .ZN(
        n10032) );
  AOI21_X1 U11176 ( .B1(n10029), .B2(n10028), .A(n4532), .ZN(n10030) );
  INV_X1 U11177 ( .A(n10030), .ZN(n10167) );
  NOR2_X1 U11178 ( .A1(n10167), .A2(n10074), .ZN(n10031) );
  AOI211_X1 U11179 ( .C1(n10163), .C2(n10077), .A(n10032), .B(n10031), .ZN(
        n10033) );
  OAI21_X1 U11180 ( .B1(n10317), .B2(n10166), .A(n10033), .ZN(P1_U3275) );
  XOR2_X1 U11181 ( .A(n10034), .B(n10036), .Z(n10042) );
  XNOR2_X1 U11182 ( .A(n6612), .B(n4806), .ZN(n10172) );
  AOI22_X1 U11183 ( .A1(n10038), .A2(n10055), .B1(n10057), .B2(n10037), .ZN(
        n10039) );
  OAI21_X1 U11184 ( .B1(n10172), .B2(n10040), .A(n10039), .ZN(n10041) );
  AOI21_X1 U11185 ( .B1(n10099), .B2(n10042), .A(n10041), .ZN(n10171) );
  OR2_X1 U11186 ( .A1(n10062), .A2(n10048), .ZN(n10043) );
  AND2_X1 U11187 ( .A1(n10044), .A2(n10043), .ZN(n10169) );
  AOI22_X1 U11188 ( .A1(n10317), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n10045), 
        .B2(n10307), .ZN(n10046) );
  OAI21_X1 U11189 ( .B1(n10048), .B2(n10047), .A(n10046), .ZN(n10051) );
  NOR2_X1 U11190 ( .A1(n10172), .A2(n10049), .ZN(n10050) );
  AOI211_X1 U11191 ( .C1(n10169), .C2(n10052), .A(n10051), .B(n10050), .ZN(
        n10053) );
  OAI21_X1 U11192 ( .B1(n10317), .B2(n10171), .A(n10053), .ZN(P1_U3276) );
  XNOR2_X1 U11193 ( .A(n10054), .B(n10072), .ZN(n10059) );
  AOI222_X1 U11194 ( .A1(n10099), .A2(n10059), .B1(n10058), .B2(n10057), .C1(
        n10056), .C2(n10055), .ZN(n10176) );
  OAI21_X1 U11195 ( .B1(n10061), .B2(n10060), .A(n10341), .ZN(n10063) );
  NOR2_X1 U11196 ( .A1(n10063), .A2(n10062), .ZN(n10173) );
  NAND2_X1 U11197 ( .A1(n10174), .A2(n10064), .ZN(n10067) );
  NAND2_X1 U11198 ( .A1(n10307), .A2(n10065), .ZN(n10066) );
  OAI211_X1 U11199 ( .C1(n10315), .C2(n8634), .A(n10067), .B(n10066), .ZN(
        n10076) );
  OR2_X1 U11200 ( .A1(n10069), .A2(n10068), .ZN(n10071) );
  NAND2_X1 U11201 ( .A1(n10071), .A2(n10070), .ZN(n10073) );
  XNOR2_X1 U11202 ( .A(n10073), .B(n10072), .ZN(n10177) );
  NOR2_X1 U11203 ( .A1(n10177), .A2(n10074), .ZN(n10075) );
  AOI211_X1 U11204 ( .C1(n10173), .C2(n10077), .A(n10076), .B(n10075), .ZN(
        n10078) );
  OAI21_X1 U11205 ( .B1(n10317), .B2(n10176), .A(n10078), .ZN(P1_U3277) );
  NAND2_X1 U11206 ( .A1(n10079), .A2(n10207), .ZN(n10080) );
  OAI211_X1 U11207 ( .C1(n10081), .C2(n10334), .A(n10080), .B(n10084), .ZN(
        n10213) );
  MUX2_X1 U11208 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n10213), .S(n10357), .Z(
        P1_U3554) );
  NAND3_X1 U11209 ( .A1(n10083), .A2(n10341), .A3(n10082), .ZN(n10085) );
  OAI211_X1 U11210 ( .C1(n10086), .C2(n10344), .A(n10085), .B(n10084), .ZN(
        n10214) );
  MUX2_X1 U11211 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n10214), .S(n10357), .Z(
        P1_U3553) );
  NAND3_X1 U11212 ( .A1(n10098), .A2(n10097), .A3(n10134), .ZN(n10094) );
  INV_X1 U11213 ( .A(n10091), .ZN(n10093) );
  MUX2_X1 U11214 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n10215), .S(n10357), .Z(
        P1_U3552) );
  AOI21_X1 U11215 ( .B1(n10207), .B2(n10102), .A(n10101), .ZN(n10103) );
  MUX2_X1 U11216 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n10216), .S(n10357), .Z(
        P1_U3551) );
  AOI21_X1 U11217 ( .B1(n10207), .B2(n10107), .A(n10106), .ZN(n10108) );
  MUX2_X1 U11218 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n10217), .S(n10357), .Z(
        P1_U3550) );
  AOI22_X1 U11219 ( .A1(n10112), .A2(n10341), .B1(n10207), .B2(n10111), .ZN(
        n10113) );
  OAI211_X1 U11220 ( .C1(n10115), .C2(n10188), .A(n10114), .B(n10113), .ZN(
        n10218) );
  MUX2_X1 U11221 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n10218), .S(n10357), .Z(
        P1_U3549) );
  AOI22_X1 U11222 ( .A1(n10117), .A2(n10341), .B1(n10207), .B2(n10116), .ZN(
        n10118) );
  OAI211_X1 U11223 ( .C1(n10120), .C2(n10188), .A(n10119), .B(n10118), .ZN(
        n10219) );
  MUX2_X1 U11224 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n10219), .S(n10357), .Z(
        P1_U3548) );
  AOI22_X1 U11225 ( .A1(n10122), .A2(n10341), .B1(n10207), .B2(n10121), .ZN(
        n10123) );
  OAI211_X1 U11226 ( .C1(n10125), .C2(n10188), .A(n10124), .B(n10123), .ZN(
        n10220) );
  MUX2_X1 U11227 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n10220), .S(n10357), .Z(
        P1_U3547) );
  AOI22_X1 U11228 ( .A1(n10127), .A2(n10341), .B1(n10207), .B2(n10126), .ZN(
        n10128) );
  OAI211_X1 U11229 ( .C1(n10130), .C2(n10188), .A(n10129), .B(n10128), .ZN(
        n10221) );
  MUX2_X1 U11230 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n10221), .S(n10357), .Z(
        P1_U3546) );
  OAI22_X1 U11231 ( .A1(n10132), .A2(n10334), .B1(n10131), .B2(n10344), .ZN(
        n10133) );
  AOI21_X1 U11232 ( .B1(n10135), .B2(n10134), .A(n10133), .ZN(n10137) );
  NAND2_X1 U11233 ( .A1(n10137), .A2(n10136), .ZN(n10222) );
  MUX2_X1 U11234 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n10222), .S(n10357), .Z(
        P1_U3545) );
  AOI211_X1 U11235 ( .C1(n10207), .C2(n10140), .A(n10139), .B(n10138), .ZN(
        n10141) );
  OAI21_X1 U11236 ( .B1(n10188), .B2(n10142), .A(n10141), .ZN(n10223) );
  MUX2_X1 U11237 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n10223), .S(n10357), .Z(
        P1_U3544) );
  AOI21_X1 U11238 ( .B1(n10207), .B2(n10144), .A(n10143), .ZN(n10145) );
  OAI211_X1 U11239 ( .C1(n10147), .C2(n10188), .A(n10146), .B(n10145), .ZN(
        n10224) );
  MUX2_X1 U11240 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n10224), .S(n10357), .Z(
        P1_U3543) );
  AOI22_X1 U11241 ( .A1(n10149), .A2(n10341), .B1(n10207), .B2(n10148), .ZN(
        n10150) );
  OAI211_X1 U11242 ( .C1(n10152), .C2(n10188), .A(n10151), .B(n10150), .ZN(
        n10225) );
  MUX2_X1 U11243 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n10225), .S(n10357), .Z(
        P1_U3542) );
  AOI21_X1 U11244 ( .B1(n10207), .B2(n10154), .A(n10153), .ZN(n10155) );
  OAI211_X1 U11245 ( .C1(n10157), .C2(n10188), .A(n10156), .B(n10155), .ZN(
        n10226) );
  MUX2_X1 U11246 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n10226), .S(n10357), .Z(
        P1_U3541) );
  AOI22_X1 U11247 ( .A1(n10159), .A2(n10341), .B1(n10207), .B2(n10158), .ZN(
        n10160) );
  OAI211_X1 U11248 ( .C1(n10162), .C2(n10188), .A(n10161), .B(n10160), .ZN(
        n10227) );
  MUX2_X1 U11249 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n10227), .S(n10357), .Z(
        P1_U3540) );
  AOI21_X1 U11250 ( .B1(n10207), .B2(n10164), .A(n10163), .ZN(n10165) );
  OAI211_X1 U11251 ( .C1(n10167), .C2(n10188), .A(n10166), .B(n10165), .ZN(
        n10228) );
  MUX2_X1 U11252 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n10228), .S(n10357), .Z(
        P1_U3539) );
  AOI22_X1 U11253 ( .A1(n10169), .A2(n10341), .B1(n10207), .B2(n10168), .ZN(
        n10170) );
  OAI211_X1 U11254 ( .C1(n10211), .C2(n10172), .A(n10171), .B(n10170), .ZN(
        n10229) );
  MUX2_X1 U11255 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n10229), .S(n10357), .Z(
        P1_U3538) );
  AOI21_X1 U11256 ( .B1(n10207), .B2(n10174), .A(n10173), .ZN(n10175) );
  OAI211_X1 U11257 ( .C1(n10188), .C2(n10177), .A(n10176), .B(n10175), .ZN(
        n10230) );
  MUX2_X1 U11258 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n10230), .S(n10357), .Z(
        P1_U3537) );
  AOI22_X1 U11259 ( .A1(n10179), .A2(n10341), .B1(n10207), .B2(n10178), .ZN(
        n10180) );
  OAI211_X1 U11260 ( .C1(n10188), .C2(n10182), .A(n10181), .B(n10180), .ZN(
        n10231) );
  MUX2_X1 U11261 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n10231), .S(n10357), .Z(
        P1_U3536) );
  AOI21_X1 U11262 ( .B1(n10207), .B2(n10184), .A(n10183), .ZN(n10185) );
  OAI211_X1 U11263 ( .C1(n10188), .C2(n10187), .A(n10186), .B(n10185), .ZN(
        n10232) );
  MUX2_X1 U11264 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n10232), .S(n10357), .Z(
        P1_U3535) );
  AND2_X1 U11265 ( .A1(n10189), .A2(n10347), .ZN(n10193) );
  OAI22_X1 U11266 ( .A1(n10191), .A2(n10334), .B1(n10190), .B2(n10344), .ZN(
        n10192) );
  MUX2_X1 U11267 ( .A(n10233), .B(P1_REG1_REG_11__SCAN_IN), .S(n10355), .Z(
        P1_U3534) );
  AOI21_X1 U11268 ( .B1(n10207), .B2(n10196), .A(n10195), .ZN(n10197) );
  OAI211_X1 U11269 ( .C1(n10199), .C2(n10211), .A(n10198), .B(n10197), .ZN(
        n10234) );
  MUX2_X1 U11270 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n10234), .S(n10357), .Z(
        P1_U3533) );
  INV_X1 U11271 ( .A(n10200), .ZN(n10205) );
  AOI22_X1 U11272 ( .A1(n10202), .A2(n10341), .B1(n10207), .B2(n10201), .ZN(
        n10203) );
  OAI211_X1 U11273 ( .C1(n10211), .C2(n10205), .A(n10204), .B(n10203), .ZN(
        n10235) );
  MUX2_X1 U11274 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n10235), .S(n10357), .Z(
        P1_U3532) );
  AOI22_X1 U11275 ( .A1(n10208), .A2(n10341), .B1(n10207), .B2(n10206), .ZN(
        n10209) );
  OAI211_X1 U11276 ( .C1(n10212), .C2(n10211), .A(n10210), .B(n10209), .ZN(
        n10236) );
  MUX2_X1 U11277 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n10236), .S(n10357), .Z(
        P1_U3531) );
  MUX2_X1 U11278 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n10213), .S(n10353), .Z(
        P1_U3522) );
  MUX2_X1 U11279 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n10214), .S(n10353), .Z(
        P1_U3521) );
  MUX2_X1 U11280 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n10215), .S(n10353), .Z(
        P1_U3520) );
  MUX2_X1 U11281 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n10216), .S(n10353), .Z(
        P1_U3519) );
  MUX2_X1 U11282 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n10217), .S(n10353), .Z(
        P1_U3518) );
  MUX2_X1 U11283 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n10218), .S(n10353), .Z(
        P1_U3517) );
  MUX2_X1 U11284 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n10219), .S(n10353), .Z(
        P1_U3516) );
  MUX2_X1 U11285 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n10220), .S(n10353), .Z(
        P1_U3515) );
  MUX2_X1 U11286 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n10221), .S(n10353), .Z(
        P1_U3514) );
  MUX2_X1 U11287 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n10222), .S(n10353), .Z(
        P1_U3513) );
  MUX2_X1 U11288 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n10223), .S(n10353), .Z(
        P1_U3512) );
  MUX2_X1 U11289 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n10224), .S(n10353), .Z(
        P1_U3511) );
  MUX2_X1 U11290 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n10225), .S(n10353), .Z(
        P1_U3510) );
  MUX2_X1 U11291 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n10226), .S(n10353), .Z(
        P1_U3508) );
  MUX2_X1 U11292 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n10227), .S(n10353), .Z(
        P1_U3505) );
  MUX2_X1 U11293 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n10228), .S(n10353), .Z(
        P1_U3502) );
  MUX2_X1 U11294 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n10229), .S(n10353), .Z(
        P1_U3499) );
  MUX2_X1 U11295 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n10230), .S(n10353), .Z(
        P1_U3496) );
  MUX2_X1 U11296 ( .A(P1_REG0_REG_13__SCAN_IN), .B(n10231), .S(n10353), .Z(
        P1_U3493) );
  MUX2_X1 U11297 ( .A(P1_REG0_REG_12__SCAN_IN), .B(n10232), .S(n10353), .Z(
        P1_U3490) );
  MUX2_X1 U11298 ( .A(n10233), .B(P1_REG0_REG_11__SCAN_IN), .S(n10351), .Z(
        P1_U3487) );
  MUX2_X1 U11299 ( .A(P1_REG0_REG_10__SCAN_IN), .B(n10234), .S(n10353), .Z(
        P1_U3484) );
  MUX2_X1 U11300 ( .A(P1_REG0_REG_9__SCAN_IN), .B(n10235), .S(n10353), .Z(
        P1_U3481) );
  MUX2_X1 U11301 ( .A(P1_REG0_REG_8__SCAN_IN), .B(n10236), .S(n10353), .Z(
        P1_U3478) );
  NOR4_X1 U11302 ( .A1(n10237), .A2(P1_IR_REG_30__SCAN_IN), .A3(n5984), .A4(
        P1_U3084), .ZN(n10238) );
  AOI21_X1 U11303 ( .B1(n10239), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n10238), 
        .ZN(n10240) );
  OAI21_X1 U11304 ( .B1(n10241), .B2(n10244), .A(n10240), .ZN(P1_U3322) );
  OAI222_X1 U11305 ( .A1(n10245), .A2(P1_U3084), .B1(n10244), .B2(n10243), 
        .C1(n10242), .C2(n10251), .ZN(P1_U3324) );
  NAND2_X1 U11306 ( .A1(n10247), .A2(n10246), .ZN(n10249) );
  OAI211_X1 U11307 ( .C1(n10251), .C2(n10250), .A(n10249), .B(n10248), .ZN(
        P1_U3325) );
  MUX2_X1 U11308 ( .A(n10252), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  INV_X1 U11309 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10466) );
  NOR2_X1 U11310 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n10253) );
  AOI21_X1 U11311 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n10253), .ZN(n10439) );
  AOI22_X1 U11312 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(n10255), .B1(
        P2_ADDR_REG_13__SCAN_IN), .B2(n10254), .ZN(n10450) );
  NOR2_X1 U11313 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(P1_ADDR_REG_4__SCAN_IN), 
        .ZN(n10264) );
  INV_X1 U11314 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n10257) );
  AOI22_X1 U11315 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(n10257), .B1(
        P1_ADDR_REG_4__SCAN_IN), .B2(n10256), .ZN(n10478) );
  NAND2_X1 U11316 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n10262) );
  XOR2_X1 U11317 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10476) );
  NAND2_X1 U11318 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n10260) );
  XOR2_X1 U11319 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(P1_ADDR_REG_2__SCAN_IN), .Z(
        n10474) );
  AOI21_X1 U11320 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10427) );
  NAND3_X1 U11321 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n10429) );
  NAND2_X1 U11322 ( .A1(n10474), .A2(n10473), .ZN(n10259) );
  NAND2_X1 U11323 ( .A1(n10262), .A2(n10261), .ZN(n10477) );
  NOR2_X1 U11324 ( .A1(n10478), .A2(n10477), .ZN(n10263) );
  NOR2_X1 U11325 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n10265), .ZN(n10462) );
  NAND2_X1 U11326 ( .A1(n10267), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n10268) );
  NAND2_X1 U11327 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n10269), .ZN(n10272) );
  NAND2_X1 U11328 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n10472), .ZN(n10271) );
  NAND2_X1 U11329 ( .A1(n10272), .A2(n10271), .ZN(n10273) );
  NAND2_X1 U11330 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n10273), .ZN(n10275) );
  NAND2_X1 U11331 ( .A1(n10275), .A2(n10274), .ZN(n10276) );
  AND2_X1 U11332 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n10276), .ZN(n10277) );
  XNOR2_X1 U11333 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n10276), .ZN(n10469) );
  NAND2_X1 U11334 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n10278) );
  OAI21_X1 U11335 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10278), .ZN(n10458) );
  NAND2_X1 U11336 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n10279) );
  OAI21_X1 U11337 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n10279), .ZN(n10455) );
  NOR2_X1 U11338 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n10280) );
  AOI21_X1 U11339 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n10280), .ZN(n10452) );
  NOR2_X1 U11340 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n10282) );
  AOI21_X1 U11341 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n10282), .ZN(n10441) );
  NAND2_X1 U11342 ( .A1(n10442), .A2(n10441), .ZN(n10440) );
  NAND2_X1 U11343 ( .A1(n10439), .A2(n10438), .ZN(n10437) );
  NOR2_X1 U11344 ( .A1(n10466), .A2(n10465), .ZN(n10286) );
  NAND2_X1 U11345 ( .A1(n10466), .A2(n10465), .ZN(n10464) );
  XOR2_X1 U11346 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .Z(n10287) );
  XNOR2_X1 U11347 ( .A(n10288), .B(n10287), .ZN(ADD_1071_U4) );
  XNOR2_X1 U11348 ( .A(P1_WR_REG_SCAN_IN), .B(P2_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U11349 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  AOI21_X1 U11350 ( .B1(n10290), .B2(n10289), .A(n4447), .ZN(n10291) );
  NAND2_X1 U11351 ( .A1(n10292), .A2(n10291), .ZN(n10297) );
  NAND2_X1 U11352 ( .A1(n10294), .A2(n10293), .ZN(n10296) );
  AND3_X1 U11353 ( .A1(n10297), .A2(n10296), .A3(n10295), .ZN(n10305) );
  OAI21_X1 U11354 ( .B1(n10300), .B2(n10299), .A(n10298), .ZN(n10303) );
  AOI22_X1 U11355 ( .A1(n10303), .A2(n10302), .B1(n10301), .B2(
        P1_ADDR_REG_18__SCAN_IN), .ZN(n10304) );
  NAND2_X1 U11356 ( .A1(n10305), .A2(n10304), .ZN(P1_U3259) );
  AOI22_X1 U11357 ( .A1(n10307), .A2(P1_REG3_REG_1__SCAN_IN), .B1(n10306), 
        .B2(n4401), .ZN(n10308) );
  OAI21_X1 U11358 ( .B1(n10310), .B2(n10309), .A(n10308), .ZN(n10312) );
  AOI211_X1 U11359 ( .C1(n10314), .C2(n10313), .A(n10312), .B(n10311), .ZN(
        n10316) );
  AOI22_X1 U11360 ( .A1(n10317), .A2(n4837), .B1(n10316), .B2(n10315), .ZN(
        P1_U3290) );
  AND2_X1 U11361 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n10328), .ZN(P1_U3292) );
  INV_X1 U11362 ( .A(n10328), .ZN(n10327) );
  NOR2_X1 U11363 ( .A1(n10327), .A2(n10318), .ZN(P1_U3293) );
  NOR2_X1 U11364 ( .A1(n10327), .A2(n10319), .ZN(P1_U3294) );
  AND2_X1 U11365 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n10328), .ZN(P1_U3295) );
  AND2_X1 U11366 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n10328), .ZN(P1_U3296) );
  AND2_X1 U11367 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n10328), .ZN(P1_U3297) );
  AND2_X1 U11368 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n10328), .ZN(P1_U3298) );
  NOR2_X1 U11369 ( .A1(n10327), .A2(n10320), .ZN(P1_U3299) );
  AND2_X1 U11370 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n10328), .ZN(P1_U3300) );
  AND2_X1 U11371 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n10328), .ZN(P1_U3301) );
  NOR2_X1 U11372 ( .A1(n10327), .A2(n10321), .ZN(P1_U3302) );
  NOR2_X1 U11373 ( .A1(n10327), .A2(n10322), .ZN(P1_U3303) );
  AND2_X1 U11374 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n10328), .ZN(P1_U3304) );
  NOR2_X1 U11375 ( .A1(n10327), .A2(n10323), .ZN(P1_U3305) );
  NOR2_X1 U11376 ( .A1(n10327), .A2(n10324), .ZN(P1_U3306) );
  AND2_X1 U11377 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n10328), .ZN(P1_U3307) );
  AND2_X1 U11378 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n10328), .ZN(P1_U3308) );
  NOR2_X1 U11379 ( .A1(n10327), .A2(n10325), .ZN(P1_U3309) );
  AND2_X1 U11380 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n10328), .ZN(P1_U3310) );
  NOR2_X1 U11381 ( .A1(n10327), .A2(n10326), .ZN(P1_U3311) );
  AND2_X1 U11382 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n10328), .ZN(P1_U3312) );
  AND2_X1 U11383 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n10328), .ZN(P1_U3313) );
  AND2_X1 U11384 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n10328), .ZN(P1_U3314) );
  AND2_X1 U11385 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n10328), .ZN(P1_U3315) );
  AND2_X1 U11386 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n10328), .ZN(P1_U3316) );
  AND2_X1 U11387 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n10328), .ZN(P1_U3317) );
  AND2_X1 U11388 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n10328), .ZN(P1_U3318) );
  AND2_X1 U11389 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n10328), .ZN(P1_U3319) );
  AND2_X1 U11390 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n10328), .ZN(P1_U3320) );
  AND2_X1 U11391 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n10328), .ZN(P1_U3321) );
  INV_X1 U11392 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n10329) );
  AOI22_X1 U11393 ( .A1(n10353), .A2(n10330), .B1(n10329), .B2(n10351), .ZN(
        P1_U3457) );
  INV_X1 U11394 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n10331) );
  AOI22_X1 U11395 ( .A1(n10353), .A2(n10332), .B1(n10331), .B2(n10351), .ZN(
        P1_U3460) );
  OAI22_X1 U11396 ( .A1(n10335), .A2(n10334), .B1(n10333), .B2(n10344), .ZN(
        n10338) );
  INV_X1 U11397 ( .A(n10336), .ZN(n10337) );
  AOI211_X1 U11398 ( .C1(n10347), .C2(n10339), .A(n10338), .B(n10337), .ZN(
        n10354) );
  AOI22_X1 U11399 ( .A1(n10353), .A2(n10354), .B1(n10340), .B2(n10351), .ZN(
        P1_U3466) );
  NAND2_X1 U11400 ( .A1(n10342), .A2(n10341), .ZN(n10343) );
  OAI21_X1 U11401 ( .B1(n10345), .B2(n10344), .A(n10343), .ZN(n10346) );
  AOI21_X1 U11402 ( .B1(n10348), .B2(n10347), .A(n10346), .ZN(n10349) );
  AND2_X1 U11403 ( .A1(n10350), .A2(n10349), .ZN(n10356) );
  AOI22_X1 U11404 ( .A1(n10353), .A2(n10356), .B1(n10352), .B2(n10351), .ZN(
        P1_U3472) );
  AOI22_X1 U11405 ( .A1(n10357), .A2(n10354), .B1(n7002), .B2(n10355), .ZN(
        P1_U3527) );
  AOI22_X1 U11406 ( .A1(n10357), .A2(n10356), .B1(n7005), .B2(n10355), .ZN(
        P1_U3529) );
  AOI22_X1 U11407 ( .A1(n10358), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n10370) );
  NOR2_X1 U11408 ( .A1(n10362), .A2(n5166), .ZN(n10360) );
  MUX2_X1 U11409 ( .A(n10360), .B(n5166), .S(n10359), .Z(n10364) );
  AOI21_X1 U11410 ( .B1(n10367), .B2(n10362), .A(n10361), .ZN(n10363) );
  OR2_X1 U11411 ( .A1(n10364), .A2(n10363), .ZN(n10369) );
  OAI211_X1 U11412 ( .C1(n10367), .C2(P2_REG1_REG_0__SCAN_IN), .A(n10366), .B(
        n10365), .ZN(n10368) );
  NAND3_X1 U11413 ( .A1(n10370), .A2(n10369), .A3(n10368), .ZN(P2_U3245) );
  INV_X1 U11414 ( .A(n10371), .ZN(n10372) );
  AND2_X1 U11415 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n10383), .ZN(P2_U3297) );
  AND2_X1 U11416 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n10383), .ZN(P2_U3298) );
  INV_X1 U11417 ( .A(n10383), .ZN(n10380) );
  NOR2_X1 U11418 ( .A1(n10380), .A2(n10374), .ZN(P2_U3299) );
  AND2_X1 U11419 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n10383), .ZN(P2_U3300) );
  AND2_X1 U11420 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n10383), .ZN(P2_U3301) );
  AND2_X1 U11421 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n10383), .ZN(P2_U3302) );
  AND2_X1 U11422 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n10383), .ZN(P2_U3303) );
  NOR2_X1 U11423 ( .A1(n10380), .A2(n10375), .ZN(P2_U3304) );
  AND2_X1 U11424 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n10383), .ZN(P2_U3305) );
  NOR2_X1 U11425 ( .A1(n10380), .A2(n10376), .ZN(P2_U3306) );
  AND2_X1 U11426 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n10383), .ZN(P2_U3307) );
  AND2_X1 U11427 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n10383), .ZN(P2_U3308) );
  AND2_X1 U11428 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n10383), .ZN(P2_U3309) );
  AND2_X1 U11429 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n10383), .ZN(P2_U3310) );
  AND2_X1 U11430 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n10383), .ZN(P2_U3311) );
  AND2_X1 U11431 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n10383), .ZN(P2_U3312) );
  AND2_X1 U11432 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n10383), .ZN(P2_U3313) );
  AND2_X1 U11433 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n10383), .ZN(P2_U3314) );
  AND2_X1 U11434 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n10383), .ZN(P2_U3315) );
  NOR2_X1 U11435 ( .A1(n10380), .A2(n10377), .ZN(P2_U3316) );
  AND2_X1 U11436 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n10383), .ZN(P2_U3317) );
  AND2_X1 U11437 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n10383), .ZN(P2_U3318) );
  AND2_X1 U11438 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n10383), .ZN(P2_U3319) );
  NOR2_X1 U11439 ( .A1(n10380), .A2(n10378), .ZN(P2_U3320) );
  AND2_X1 U11440 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n10383), .ZN(P2_U3321) );
  AND2_X1 U11441 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n10383), .ZN(P2_U3322) );
  AND2_X1 U11442 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n10383), .ZN(P2_U3323) );
  AND2_X1 U11443 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n10383), .ZN(P2_U3324) );
  NOR2_X1 U11444 ( .A1(n10380), .A2(n10379), .ZN(P2_U3325) );
  AND2_X1 U11445 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n10383), .ZN(P2_U3326) );
  AOI22_X1 U11446 ( .A1(n10382), .A2(n10385), .B1(n10381), .B2(n10383), .ZN(
        P2_U3437) );
  AOI22_X1 U11447 ( .A1(n10386), .A2(n10385), .B1(n10384), .B2(n10383), .ZN(
        P2_U3438) );
  AOI211_X1 U11448 ( .C1(n10408), .C2(n10389), .A(n10388), .B(n10387), .ZN(
        n10390) );
  OAI21_X1 U11449 ( .B1(n10414), .B2(n10391), .A(n10390), .ZN(n10392) );
  INV_X1 U11450 ( .A(n10392), .ZN(n10420) );
  AOI22_X1 U11451 ( .A1(n10418), .A2(n10420), .B1(n5137), .B2(n10416), .ZN(
        P2_U3457) );
  OAI21_X1 U11452 ( .B1(n10394), .B2(n10403), .A(n10393), .ZN(n10395) );
  AOI211_X1 U11453 ( .C1(n10397), .C2(n10399), .A(n10396), .B(n10395), .ZN(
        n10421) );
  AOI22_X1 U11454 ( .A1(n10418), .A2(n10421), .B1(n5226), .B2(n10416), .ZN(
        P2_U3463) );
  NAND3_X1 U11455 ( .A1(n10400), .A2(n10399), .A3(n10398), .ZN(n10402) );
  OAI211_X1 U11456 ( .C1(n10404), .C2(n10403), .A(n10402), .B(n10401), .ZN(
        n10406) );
  NOR2_X1 U11457 ( .A1(n10406), .A2(n10405), .ZN(n10423) );
  AOI22_X1 U11458 ( .A1(n10418), .A2(n10423), .B1(n5267), .B2(n10416), .ZN(
        P2_U3469) );
  AOI22_X1 U11459 ( .A1(n10410), .A2(n10409), .B1(n10408), .B2(n10407), .ZN(
        n10411) );
  OAI211_X1 U11460 ( .C1(n10414), .C2(n10413), .A(n10412), .B(n10411), .ZN(
        n10415) );
  INV_X1 U11461 ( .A(n10415), .ZN(n10425) );
  INV_X1 U11462 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10417) );
  AOI22_X1 U11463 ( .A1(n10418), .A2(n10425), .B1(n10417), .B2(n10416), .ZN(
        P2_U3472) );
  AOI22_X1 U11464 ( .A1(n10426), .A2(n10420), .B1(n10419), .B2(n10424), .ZN(
        P2_U3522) );
  AOI22_X1 U11465 ( .A1(n10426), .A2(n10421), .B1(n7217), .B2(n10424), .ZN(
        P2_U3524) );
  INV_X1 U11466 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10422) );
  AOI22_X1 U11467 ( .A1(n10426), .A2(n10423), .B1(n10422), .B2(n10424), .ZN(
        P2_U3526) );
  AOI22_X1 U11468 ( .A1(n10426), .A2(n10425), .B1(n7255), .B2(n10424), .ZN(
        P2_U3527) );
  INV_X1 U11469 ( .A(n10427), .ZN(n10428) );
  NAND2_X1 U11470 ( .A1(n10429), .A2(n10428), .ZN(n10430) );
  XNOR2_X1 U11471 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n10430), .ZN(ADD_1071_U5)
         );
  INV_X1 U11472 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n10432) );
  AOI22_X1 U11473 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .B1(n10432), .B2(n10431), .ZN(ADD_1071_U46) );
  AOI21_X1 U11474 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n10433), .ZN(n10436) );
  OAI21_X1 U11475 ( .B1(n10436), .B2(n10435), .A(n10434), .ZN(ADD_1071_U56) );
  OAI21_X1 U11476 ( .B1(n10439), .B2(n10438), .A(n10437), .ZN(ADD_1071_U57) );
  OAI21_X1 U11477 ( .B1(n10442), .B2(n10441), .A(n10440), .ZN(ADD_1071_U58) );
  AOI22_X1 U11478 ( .A1(P1_ADDR_REG_14__SCAN_IN), .A2(n10444), .B1(
        P2_ADDR_REG_14__SCAN_IN), .B2(n10443), .ZN(n10446) );
  AOI21_X1 U11479 ( .B1(n10447), .B2(n10446), .A(n10445), .ZN(ADD_1071_U59) );
  AOI21_X1 U11480 ( .B1(n10450), .B2(n10449), .A(n10448), .ZN(ADD_1071_U60) );
  OAI21_X1 U11481 ( .B1(n10453), .B2(n10452), .A(n10451), .ZN(ADD_1071_U61) );
  AOI21_X1 U11482 ( .B1(n10456), .B2(n10455), .A(n10454), .ZN(ADD_1071_U62) );
  AOI21_X1 U11483 ( .B1(n10459), .B2(n10458), .A(n10457), .ZN(ADD_1071_U63) );
  XOR2_X1 U11484 ( .A(n10460), .B(P2_ADDR_REG_6__SCAN_IN), .Z(ADD_1071_U50) );
  NOR2_X1 U11485 ( .A1(n10462), .A2(n10461), .ZN(n10463) );
  XOR2_X1 U11486 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n10463), .Z(ADD_1071_U51) );
  OAI21_X1 U11487 ( .B1(n10466), .B2(n10465), .A(n10464), .ZN(n10467) );
  XNOR2_X1 U11488 ( .A(n10467), .B(P1_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  AOI21_X1 U11489 ( .B1(n10470), .B2(n10469), .A(n10468), .ZN(ADD_1071_U47) );
  XOR2_X1 U11490 ( .A(n10471), .B(P2_ADDR_REG_8__SCAN_IN), .Z(ADD_1071_U48) );
  XOR2_X1 U11491 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(n10472), .Z(ADD_1071_U49) );
  XOR2_X1 U11492 ( .A(n10474), .B(n10473), .Z(ADD_1071_U54) );
  XOR2_X1 U11493 ( .A(n10475), .B(n10476), .Z(ADD_1071_U53) );
  XNOR2_X1 U11494 ( .A(n10478), .B(n10477), .ZN(ADD_1071_U52) );
  CLKBUF_X1 U4910 ( .A(n5482), .Z(n4393) );
  INV_X2 U4930 ( .A(n5225), .ZN(n5744) );
  CLKBUF_X1 U4979 ( .A(n5207), .Z(n7154) );
  CLKBUF_X1 U4987 ( .A(n9906), .Z(n4531) );
  CLKBUF_X1 U5161 ( .A(n8742), .Z(n8662) );
  CLKBUF_X1 U5928 ( .A(n6729), .Z(n4575) );
  CLKBUF_X1 U6203 ( .A(n7625), .Z(n4377) );
endmodule

