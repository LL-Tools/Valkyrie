

module b21_C_gen_AntiSAT_k_128_6 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2, 
        keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7, 
        keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12, 
        keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17, 
        keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22, 
        keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27, 
        keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32, 
        keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37, 
        keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42, 
        keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47, 
        keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52, 
        keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57, 
        keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62, 
        keyinput_f63, keyinput_g0, keyinput_g1, keyinput_g2, keyinput_g3, 
        keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, keyinput_g8, 
        keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, keyinput_g13, 
        keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, keyinput_g18, 
        keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, keyinput_g23, 
        keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, keyinput_g28, 
        keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, keyinput_g33, 
        keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, keyinput_g38, 
        keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, keyinput_g43, 
        keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, keyinput_g48, 
        keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, keyinput_g53, 
        keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, keyinput_g58, 
        keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, keyinput_g63, 
        ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58, 
        ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63, 
        ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51, 
        ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46, 
        U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, 
        P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, 
        P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, 
        P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, 
        P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440, P1_U3441, 
        P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, 
        P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, 
        P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, 
        P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, 
        P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463, P1_U3466, 
        P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484, P1_U3487, 
        P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505, P1_U3508, 
        P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, 
        P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, 
        P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, 
        P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, 
        P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, 
        P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, 
        P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289, P1_U3288, 
        P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, 
        P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, 
        P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, 
        P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262, P1_U3261, 
        P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, 
        P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, 
        P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241, P1_U3555, 
        P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, 
        P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, 
        P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, 
        P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, 
        P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238, P1_U3237, 
        P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, 
        P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, 
        P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, 
        P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084, P1_U3083, 
        P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354, P2_U3353, 
        P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347, P2_U3346, 
        P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340, P2_U3339, 
        P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333, P2_U3332, 
        P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437, P2_U3438, 
        P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, 
        P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, 
        P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, 
        P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, 
        P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, 
        P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, 
        P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502, P2_U3505, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, 
        P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533, P2_U3534, 
        P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, 
        P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, 
        P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294, P2_U3293, 
        P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, 
        P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, 
        P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, 
        P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, 
        P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, 
        P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, 
        P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3552, 
        P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, 
        P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565, P2_U3566, 
        P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572, P2_U3573, 
        P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579, P2_U3580, 
        P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152, P2_U3151, 
        P2_U3966 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2,
         keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7,
         keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12,
         keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17,
         keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22,
         keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27,
         keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32,
         keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37,
         keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42,
         keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47,
         keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52,
         keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57,
         keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62,
         keyinput_f63, keyinput_g0, keyinput_g1, keyinput_g2, keyinput_g3,
         keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, keyinput_g8,
         keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, keyinput_g13,
         keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, keyinput_g18,
         keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, keyinput_g23,
         keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, keyinput_g28,
         keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, keyinput_g33,
         keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, keyinput_g38,
         keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, keyinput_g43,
         keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, keyinput_g48,
         keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, keyinput_g53,
         keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, keyinput_g58,
         keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, keyinput_g63;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319,
         n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329,
         n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339,
         n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349,
         n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359,
         n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369,
         n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379,
         n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389,
         n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399,
         n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409,
         n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419,
         n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429,
         n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439,
         n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449,
         n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459,
         n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469,
         n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479,
         n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489,
         n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499,
         n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509,
         n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519,
         n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529,
         n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539,
         n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549,
         n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559,
         n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569,
         n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579,
         n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589,
         n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599,
         n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609,
         n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619,
         n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
         n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
         n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
         n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
         n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669,
         n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679,
         n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689,
         n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
         n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
         n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719,
         n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729,
         n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739,
         n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749,
         n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759,
         n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769,
         n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779,
         n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789,
         n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799,
         n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809,
         n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819,
         n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829,
         n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839,
         n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849,
         n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859,
         n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869,
         n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879,
         n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889,
         n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899,
         n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909,
         n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919,
         n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929,
         n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939,
         n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949,
         n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959,
         n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969,
         n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979,
         n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989,
         n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999,
         n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009,
         n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019,
         n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029,
         n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039,
         n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049,
         n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059,
         n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069,
         n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079,
         n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089,
         n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099,
         n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109,
         n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119,
         n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129,
         n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139,
         n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149,
         n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159,
         n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169,
         n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179,
         n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189,
         n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199,
         n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209,
         n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219,
         n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229,
         n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239,
         n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249,
         n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259,
         n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269,
         n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279,
         n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289,
         n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299,
         n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309,
         n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319,
         n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329,
         n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339,
         n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349,
         n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359,
         n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369,
         n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379,
         n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389,
         n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399,
         n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409,
         n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419,
         n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429,
         n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439,
         n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449,
         n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459,
         n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469,
         n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479,
         n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489,
         n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499,
         n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509,
         n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519,
         n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529,
         n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539,
         n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549,
         n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559,
         n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5568, n5569, n5570,
         n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580,
         n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590,
         n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600,
         n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610,
         n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620,
         n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630,
         n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640,
         n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650,
         n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660,
         n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670,
         n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680,
         n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690,
         n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700,
         n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710,
         n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720,
         n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730,
         n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740,
         n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750,
         n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760,
         n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770,
         n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780,
         n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790,
         n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800,
         n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810,
         n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820,
         n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830,
         n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840,
         n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850,
         n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860,
         n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870,
         n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880,
         n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890,
         n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900,
         n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910,
         n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920,
         n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930,
         n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940,
         n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950,
         n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960,
         n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970,
         n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980,
         n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990,
         n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000,
         n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010,
         n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020,
         n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030,
         n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040,
         n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050,
         n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060,
         n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070,
         n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080,
         n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090,
         n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100,
         n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110,
         n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120,
         n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130,
         n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140,
         n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150,
         n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160,
         n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170,
         n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180,
         n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190,
         n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200,
         n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210,
         n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220,
         n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230,
         n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240,
         n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250,
         n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260,
         n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270,
         n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280,
         n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290,
         n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300,
         n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310,
         n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320,
         n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330,
         n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340,
         n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350,
         n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360,
         n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370,
         n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380,
         n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390,
         n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400,
         n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410,
         n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420,
         n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430,
         n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440,
         n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450,
         n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460,
         n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470,
         n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480,
         n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490,
         n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500,
         n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510,
         n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520,
         n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530,
         n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540,
         n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550,
         n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560,
         n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570,
         n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580,
         n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590,
         n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600,
         n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610,
         n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620,
         n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630,
         n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640,
         n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650,
         n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660,
         n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670,
         n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680,
         n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690,
         n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700,
         n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710,
         n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720,
         n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730,
         n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740,
         n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750,
         n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760,
         n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770,
         n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780,
         n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790,
         n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800,
         n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810,
         n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820,
         n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830,
         n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840,
         n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850,
         n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860,
         n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870,
         n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880,
         n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890,
         n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900,
         n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910,
         n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920,
         n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930,
         n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940,
         n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950,
         n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960,
         n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970,
         n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980,
         n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990,
         n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000,
         n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010,
         n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020,
         n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030,
         n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040,
         n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050,
         n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060,
         n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070,
         n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080,
         n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090,
         n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100,
         n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110,
         n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120,
         n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130,
         n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140,
         n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150,
         n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160,
         n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170,
         n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180,
         n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190,
         n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200,
         n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210,
         n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220,
         n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230,
         n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240,
         n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250,
         n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260,
         n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270,
         n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280,
         n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290,
         n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300,
         n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310,
         n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320,
         n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330,
         n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340,
         n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350,
         n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360,
         n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370,
         n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380,
         n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390,
         n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400,
         n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410,
         n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420,
         n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430,
         n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440,
         n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450,
         n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460,
         n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470,
         n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480,
         n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490,
         n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500,
         n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510,
         n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520,
         n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530,
         n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540,
         n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550,
         n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560,
         n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570,
         n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580,
         n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590,
         n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600,
         n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610,
         n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620,
         n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630,
         n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640,
         n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650,
         n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660,
         n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670,
         n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680,
         n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690,
         n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700,
         n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710,
         n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720,
         n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730,
         n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740,
         n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750,
         n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760,
         n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770,
         n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780,
         n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790,
         n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800,
         n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810,
         n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820,
         n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830,
         n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840,
         n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850,
         n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860,
         n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870,
         n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880,
         n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890,
         n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900,
         n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910,
         n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920,
         n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930,
         n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940,
         n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950,
         n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960,
         n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970,
         n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980,
         n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990,
         n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000,
         n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010,
         n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020,
         n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030,
         n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040,
         n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050,
         n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060,
         n8061, n8062, n8063, n8064, n8065, n8067, n8068, n8069, n8070, n8071,
         n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081,
         n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091,
         n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101,
         n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111,
         n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121,
         n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131,
         n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141,
         n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151,
         n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161,
         n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171,
         n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181,
         n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191,
         n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201,
         n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211,
         n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221,
         n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231,
         n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241,
         n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251,
         n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261,
         n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271,
         n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281,
         n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291,
         n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301,
         n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311,
         n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321,
         n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331,
         n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341,
         n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351,
         n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361,
         n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371,
         n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381,
         n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391,
         n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401,
         n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411,
         n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421,
         n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431,
         n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441,
         n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451,
         n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461,
         n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471,
         n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481,
         n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491,
         n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501,
         n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511,
         n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521,
         n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531,
         n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541,
         n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551,
         n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561,
         n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571,
         n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581,
         n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591,
         n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601,
         n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611,
         n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621,
         n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631,
         n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641,
         n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651,
         n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661,
         n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671,
         n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681,
         n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691,
         n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701,
         n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711,
         n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721,
         n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731,
         n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741,
         n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751,
         n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761,
         n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771,
         n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781,
         n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791,
         n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801,
         n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811,
         n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821,
         n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831,
         n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841,
         n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851,
         n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861,
         n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871,
         n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881,
         n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891,
         n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901,
         n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911,
         n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921,
         n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931,
         n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941,
         n8942, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081;

  INV_X1 U4815 ( .A(n5818), .ZN(n5242) );
  INV_X1 U4816 ( .A(n5512), .ZN(n5368) );
  XNOR2_X1 U4818 ( .A(n5626), .B(P1_IR_REG_30__SCAN_IN), .ZN(n5631) );
  NAND2_X1 U4819 ( .A1(n5812), .A2(n5811), .ZN(n7926) );
  INV_X1 U4820 ( .A(n7926), .ZN(n7921) );
  INV_X1 U4821 ( .A(n6049), .ZN(n7568) );
  NOR2_X1 U4822 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n4654) );
  AND2_X1 U4823 ( .A1(n5224), .A2(n5223), .ZN(n5471) );
  INV_X1 U4824 ( .A(n5512), .ZN(n5465) );
  INV_X1 U4825 ( .A(n8944), .ZN(n6379) );
  XNOR2_X1 U4826 ( .A(n5557), .B(n5556), .ZN(n5948) );
  AND2_X1 U4827 ( .A1(n4817), .A2(n4747), .ZN(n4310) );
  OR2_X1 U4828 ( .A1(n5013), .A2(n4832), .ZN(n4311) );
  INV_X2 U4829 ( .A(n4667), .ZN(n8616) );
  OAI21_X2 U4830 ( .B1(n8642), .B2(n4664), .A(n4662), .ZN(n4667) );
  NAND3_X2 U4831 ( .A1(n6032), .A2(n6031), .A3(n4815), .ZN(n8891) );
  NAND2_X1 U4832 ( .A1(n6938), .A2(n8790), .ZN(n7094) );
  AND2_X4 U4833 ( .A1(n7937), .A2(n5223), .ZN(n5301) );
  AOI211_X2 U4834 ( .C1(n9278), .C2(n9664), .A(n9277), .B(n9276), .ZN(n9279)
         );
  INV_X2 U4835 ( .A(n5471), .ZN(n4312) );
  INV_X1 U4836 ( .A(n4312), .ZN(n4313) );
  INV_X4 U4837 ( .A(n4312), .ZN(n4314) );
  NAND2_X1 U4838 ( .A1(n9369), .A2(n5630), .ZN(n4315) );
  NAND2_X1 U4839 ( .A1(n9369), .A2(n5630), .ZN(n4316) );
  NAND2_X1 U4840 ( .A1(n9369), .A2(n5630), .ZN(n6044) );
  NOR2_X2 U4841 ( .A1(n5492), .A2(n7699), .ZN(n5491) );
  OAI22_X1 U4842 ( .A1(n8293), .A2(n5395), .B1(n8459), .B2(n8056), .ZN(n8266)
         );
  OAI211_X1 U4843 ( .C1(n7436), .C2(n7435), .A(n7434), .B(n7433), .ZN(n8660)
         );
  NAND2_X1 U4844 ( .A1(n7655), .A2(n7658), .ZN(n7820) );
  INV_X4 U4845 ( .A(n6049), .ZN(n7592) );
  NAND4_X1 U4846 ( .A1(n5248), .A2(n5247), .A3(n5246), .A4(n5245), .ZN(n8068)
         );
  INV_X2 U4847 ( .A(n7564), .ZN(n5923) );
  INV_X1 U4848 ( .A(n7579), .ZN(n6055) );
  INV_X2 U4849 ( .A(n5859), .ZN(n5875) );
  AND2_X1 U4850 ( .A1(n4693), .A2(n4348), .ZN(n6014) );
  NAND4_X1 U4851 ( .A1(n6048), .A2(n6047), .A3(n6046), .A4(n6045), .ZN(n8942)
         );
  CLKBUF_X3 U4852 ( .A(n4333), .Z(n7555) );
  NAND2_X2 U4853 ( .A1(n5948), .A2(n6257), .ZN(n6030) );
  INV_X4 U4854 ( .A(n4829), .ZN(n5918) );
  AND2_X1 U4855 ( .A1(n4447), .A2(n5514), .ZN(n8418) );
  AND2_X1 U4856 ( .A1(n4454), .A2(n4457), .ZN(n4446) );
  NAND2_X1 U4857 ( .A1(n8184), .A2(n7791), .ZN(n8156) );
  AND2_X1 U4858 ( .A1(n4727), .A2(n4726), .ZN(n4725) );
  NAND2_X1 U4859 ( .A1(n8193), .A2(n5506), .ZN(n8197) );
  AND2_X1 U4860 ( .A1(n7784), .A2(n7785), .ZN(n8191) );
  NAND2_X1 U4861 ( .A1(n5164), .A2(n5163), .ZN(n8427) );
  XNOR2_X1 U4862 ( .A(n5166), .B(n5165), .ZN(n7402) );
  NAND2_X1 U4863 ( .A1(n8353), .A2(n8352), .ZN(n8351) );
  AND2_X1 U4864 ( .A1(n8371), .A2(n5356), .ZN(n8353) );
  NAND2_X1 U4865 ( .A1(n4587), .A2(n4928), .ZN(n5154) );
  INV_X1 U4866 ( .A(n5150), .ZN(n4587) );
  NAND2_X1 U4867 ( .A1(n5148), .A2(n5147), .ZN(n8442) );
  OR2_X1 U4868 ( .A1(n7024), .A2(n7834), .ZN(n7026) );
  NAND2_X1 U4869 ( .A1(n5129), .A2(n5128), .ZN(n4907) );
  AOI22_X1 U4870 ( .A1(n9789), .A2(n6932), .B1(n6941), .B2(n8938), .ZN(n6933)
         );
  CLKBUF_X1 U4871 ( .A(n5831), .Z(n8047) );
  NAND2_X1 U4872 ( .A1(n4891), .A2(n4813), .ZN(n5123) );
  NAND2_X1 U4873 ( .A1(n7310), .A2(n7309), .ZN(n9330) );
  INV_X1 U4874 ( .A(n9656), .ZN(n7268) );
  NAND2_X1 U4875 ( .A1(n7077), .A2(n7076), .ZN(n9665) );
  AND2_X1 U4876 ( .A1(n7702), .A2(n7683), .ZN(n7678) );
  AND2_X1 U4877 ( .A1(n7171), .A2(n7170), .ZN(n9656) );
  NAND2_X1 U4878 ( .A1(n5068), .A2(n5067), .ZN(n6955) );
  NAND2_X1 U4879 ( .A1(n4410), .A2(n6429), .ZN(n6510) );
  AND2_X1 U4880 ( .A1(n7695), .A2(n7696), .ZN(n7828) );
  AND2_X1 U4881 ( .A1(n6512), .A2(n8839), .ZN(n8836) );
  AND2_X1 U4882 ( .A1(n6042), .A2(n6043), .ZN(n6102) );
  NAND2_X1 U4883 ( .A1(n6832), .A2(n6831), .ZN(n7066) );
  OAI21_X1 U4884 ( .B1(n6391), .B2(n4638), .A(n4362), .ZN(n8837) );
  AND2_X1 U4885 ( .A1(n6353), .A2(n6352), .ZN(n9892) );
  OR2_X1 U4886 ( .A1(n9827), .A2(n6567), .ZN(n8839) );
  NOR2_X1 U4887 ( .A1(n5853), .A2(n5852), .ZN(n5858) );
  NOR2_X1 U4888 ( .A1(n5927), .A2(n5851), .ZN(n5852) );
  OAI21_X1 U4889 ( .B1(n6055), .B2(n6014), .A(n5920), .ZN(n5921) );
  AND4_X1 U4890 ( .A1(n5232), .A2(n5231), .A3(n5230), .A4(n5229), .ZN(n7623)
         );
  NAND2_X1 U4891 ( .A1(n5850), .A2(n7579), .ZN(n5927) );
  CLKBUF_X1 U4892 ( .A(n5435), .Z(n5508) );
  NAND2_X1 U4893 ( .A1(n4514), .A2(n4837), .ZN(n5034) );
  AND2_X2 U4894 ( .A1(n6256), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U4006) );
  AND3_X1 U4895 ( .A1(n6054), .A2(n6053), .A3(n6052), .ZN(n9863) );
  AND2_X2 U4896 ( .A1(n7937), .A2(n7400), .ZN(n5435) );
  OR3_X2 U4897 ( .A1(n7162), .A2(n7010), .A3(n7064), .ZN(n6090) );
  NAND4_X2 U4898 ( .A1(n5879), .A2(n4756), .A3(n4755), .A4(n4754), .ZN(n6007)
         );
  INV_X1 U4899 ( .A(n5036), .ZN(n5059) );
  XNOR2_X1 U4900 ( .A(n5535), .B(n5553), .ZN(n7162) );
  NAND2_X2 U4901 ( .A1(n5631), .A2(n5630), .ZN(n5933) );
  AOI21_X1 U4902 ( .B1(n4515), .B2(n4518), .A(n4512), .ZN(n4511) );
  AND2_X1 U4903 ( .A1(n4711), .A2(n4516), .ZN(n4515) );
  CLKBUF_X1 U4904 ( .A(n4993), .Z(n7397) );
  XNOR2_X1 U4905 ( .A(n4978), .B(P2_IR_REG_19__SCAN_IN), .ZN(n9946) );
  AOI21_X1 U4906 ( .B1(n4840), .B2(n4714), .A(n4360), .ZN(n4713) );
  NAND2_X1 U4907 ( .A1(n4368), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5537) );
  NAND2_X1 U4908 ( .A1(n5193), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4968) );
  OAI21_X1 U4909 ( .B1(n4483), .B2(n4801), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n4482) );
  NAND2_X1 U4910 ( .A1(n9364), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5626) );
  AOI21_X1 U4911 ( .B1(n6108), .B2(P1_IR_REG_31__SCAN_IN), .A(n4675), .ZN(
        n4674) );
  NAND2_X1 U4912 ( .A1(n4676), .A2(n5544), .ZN(n4675) );
  XNOR2_X1 U4913 ( .A(n4836), .B(n9568), .ZN(n5026) );
  INV_X2 U4914 ( .A(n8530), .ZN(n7939) );
  BUF_X2 U4915 ( .A(n5918), .Z(n4594) );
  AND2_X1 U4916 ( .A1(n4343), .A2(n4959), .ZN(n4752) );
  AND4_X1 U4917 ( .A1(n4653), .A2(n5528), .A3(n4654), .A4(n5568), .ZN(n4652)
         );
  AND4_X1 U4918 ( .A1(n5526), .A2(n5525), .A3(n5604), .A4(n5524), .ZN(n5527)
         );
  INV_X1 U4919 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5661) );
  INV_X2 U4920 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  INV_X1 U4921 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5604) );
  INV_X1 U4922 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5523) );
  INV_X1 U4923 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5528) );
  NOR2_X1 U4924 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n4412) );
  INV_X1 U4925 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5200) );
  AND2_X1 U4926 ( .A1(P1_ADDR_REG_19__SCAN_IN), .A2(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n9592) );
  INV_X1 U4927 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5554) );
  INV_X1 U4928 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5541) );
  INV_X1 U4929 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5553) );
  INV_X1 U4930 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5546) );
  INV_X1 U4931 ( .A(n6298), .ZN(n5851) );
  NAND4_X2 U4932 ( .A1(n5670), .A2(n5669), .A3(n5668), .A4(n5667), .ZN(n6298)
         );
  OAI21_X2 U4933 ( .B1(n7201), .B2(n4670), .A(n4668), .ZN(n7436) );
  OR2_X1 U4934 ( .A1(n8454), .A2(n8247), .ZN(n7768) );
  OR2_X1 U4935 ( .A1(n8497), .A2(n7111), .ZN(n7725) );
  OR2_X1 U4936 ( .A1(n9271), .A2(n9085), .ZN(n9033) );
  NAND2_X1 U4937 ( .A1(n5058), .A2(n5057), .ZN(n4857) );
  INV_X1 U4938 ( .A(n5682), .ZN(n5647) );
  NAND2_X1 U4939 ( .A1(n5682), .A2(n5918), .ZN(n5035) );
  AND2_X1 U4940 ( .A1(n7722), .A2(n7723), .ZN(n4537) );
  INV_X1 U4941 ( .A(n6008), .ZN(n4409) );
  OR2_X1 U4942 ( .A1(n8427), .A2(n8157), .ZN(n7791) );
  XNOR2_X1 U4943 ( .A(n6495), .B(n8068), .ZN(n7821) );
  NOR2_X1 U4944 ( .A1(n4574), .A2(n5019), .ZN(n4573) );
  INV_X1 U4945 ( .A(n4577), .ZN(n4574) );
  OR2_X1 U4946 ( .A1(n8992), .A2(n8772), .ZN(n8877) );
  INV_X1 U4947 ( .A(n9374), .ZN(n5630) );
  OAI21_X1 U4948 ( .B1(n4635), .B2(n4632), .A(n4631), .ZN(n4630) );
  NAND2_X1 U4949 ( .A1(n4635), .A2(n9034), .ZN(n4631) );
  NOR2_X1 U4950 ( .A1(n9051), .A2(n4633), .ZN(n4632) );
  INV_X1 U4951 ( .A(n9034), .ZN(n4633) );
  OR2_X1 U4952 ( .A1(n9061), .A2(n8758), .ZN(n9034) );
  NAND2_X1 U4953 ( .A1(n9100), .A2(n9116), .ZN(n4781) );
  NAND2_X1 U4954 ( .A1(n9281), .A2(n9116), .ZN(n9030) );
  OR2_X1 U4955 ( .A1(n9306), .A2(n9149), .ZN(n7361) );
  OAI21_X1 U4956 ( .B1(n4793), .B2(n4797), .A(n9220), .ZN(n4792) );
  NAND2_X1 U4957 ( .A1(n4409), .A2(n6387), .ZN(n6391) );
  NAND2_X1 U4958 ( .A1(n6030), .A2(n4595), .ZN(n6350) );
  NAND2_X1 U4959 ( .A1(n5553), .A2(n5554), .ZN(n5558) );
  NAND2_X1 U4960 ( .A1(n4940), .A2(n4939), .ZN(n5171) );
  NAND2_X1 U4961 ( .A1(n5166), .A2(n5165), .ZN(n4940) );
  NAND2_X1 U4962 ( .A1(n4588), .A2(n4923), .ZN(n5150) );
  NAND2_X1 U4963 ( .A1(n4921), .A2(n5145), .ZN(n4588) );
  NAND2_X1 U4964 ( .A1(n4902), .A2(n4901), .ZN(n5129) );
  AND2_X1 U4965 ( .A1(n4906), .A2(n4905), .ZN(n5128) );
  NAND2_X1 U4966 ( .A1(n4886), .A2(n4885), .ZN(n5113) );
  NAND2_X1 U4967 ( .A1(n4598), .A2(n4596), .ZN(n4886) );
  AOI21_X1 U4968 ( .B1(n4599), .B2(n4330), .A(n4597), .ZN(n4596) );
  AND2_X1 U4969 ( .A1(n4885), .A2(n4884), .ZN(n5100) );
  INV_X1 U4970 ( .A(n4600), .ZN(n4599) );
  OAI21_X1 U4971 ( .B1(n4603), .B2(n4330), .A(n4880), .ZN(n4600) );
  OAI211_X1 U4972 ( .C1(n4857), .C2(n4606), .A(n4416), .B(n4864), .ZN(n5077)
         );
  NAND2_X1 U4973 ( .A1(n4417), .A2(n4607), .ZN(n4416) );
  INV_X1 U4974 ( .A(n4610), .ZN(n4417) );
  AND2_X1 U4975 ( .A1(n4871), .A2(n4870), .ZN(n5076) );
  NAND2_X1 U4976 ( .A1(n4864), .A2(n4863), .ZN(n5069) );
  XNOR2_X1 U4977 ( .A(n4859), .B(SI_11_), .ZN(n4858) );
  AND2_X1 U4978 ( .A1(n4856), .A2(n4855), .ZN(n5057) );
  NAND2_X1 U4979 ( .A1(n9592), .A2(n4440), .ZN(n4823) );
  INV_X1 U4980 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4821) );
  INV_X1 U4981 ( .A(n8064), .ZN(n6246) );
  NAND2_X1 U4982 ( .A1(n5224), .A2(n7400), .ZN(n5512) );
  NAND2_X1 U4983 ( .A1(n5445), .A2(n4317), .ZN(n4729) );
  NAND2_X1 U4984 ( .A1(n4728), .A2(n4317), .ZN(n4727) );
  INV_X1 U4985 ( .A(n4731), .ZN(n4728) );
  AOI21_X1 U4986 ( .B1(n4732), .B2(n5445), .A(n8172), .ZN(n4731) );
  INV_X1 U4987 ( .A(n5442), .ZN(n4732) );
  AND2_X1 U4988 ( .A1(n5441), .A2(n5440), .ZN(n8181) );
  OR2_X1 U4989 ( .A1(n8202), .A2(n4312), .ZN(n5441) );
  AND2_X1 U4990 ( .A1(n8261), .A2(n7768), .ZN(n4722) );
  XNOR2_X1 U4991 ( .A(n8448), .B(n8229), .ZN(n8261) );
  NAND2_X1 U4992 ( .A1(n4443), .A2(n4441), .ZN(n8277) );
  NOR2_X1 U4993 ( .A1(n8273), .A2(n4442), .ZN(n4441) );
  INV_X1 U4994 ( .A(n7762), .ZN(n4442) );
  AOI21_X1 U4995 ( .B1(n4736), .B2(n4324), .A(n4353), .ZN(n4733) );
  OR2_X1 U4996 ( .A1(n8480), .A2(n8031), .ZN(n7734) );
  NAND2_X1 U4997 ( .A1(n8374), .A2(n7730), .ZN(n4720) );
  NAND2_X1 U4998 ( .A1(n7026), .A2(n4345), .ZN(n5341) );
  NOR2_X1 U4999 ( .A1(n4710), .A2(n4709), .ZN(n4708) );
  NAND2_X1 U5000 ( .A1(n7725), .A2(n5500), .ZN(n4709) );
  OAI21_X1 U5001 ( .B1(n8419), .B2(n8503), .A(n4456), .ZN(n4455) );
  NAND2_X1 U5002 ( .A1(n5044), .A2(n5043), .ZN(n6625) );
  INV_X1 U5003 ( .A(n4581), .ZN(n4580) );
  INV_X1 U5004 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5031) );
  INV_X1 U5005 ( .A(n9313), .ZN(n7348) );
  INV_X1 U5006 ( .A(n4663), .ZN(n4662) );
  OAI21_X1 U5007 ( .B1(n4664), .B2(n4666), .A(n4335), .ZN(n4663) );
  NAND2_X1 U5008 ( .A1(n9019), .A2(n9018), .ZN(n4757) );
  OR2_X1 U5009 ( .A1(n9281), .A2(n9116), .ZN(n9082) );
  AND2_X1 U5010 ( .A1(n9001), .A2(n9000), .ZN(n9004) );
  NAND2_X1 U5011 ( .A1(n7217), .A2(n7216), .ZN(n7302) );
  NAND2_X1 U5012 ( .A1(n7268), .A2(n8934), .ZN(n7216) );
  NAND2_X1 U5013 ( .A1(n4785), .A2(n4783), .ZN(n7214) );
  AND2_X1 U5014 ( .A1(n7095), .A2(n4784), .ZN(n4783) );
  NAND2_X1 U5015 ( .A1(n9672), .A2(n7098), .ZN(n4784) );
  OR2_X1 U5016 ( .A1(n9634), .A2(n9672), .ZN(n4782) );
  INV_X1 U5017 ( .A(n6067), .ZN(n7338) );
  INV_X1 U5018 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5848) );
  NOR2_X1 U5019 ( .A1(n6115), .A2(n6116), .ZN(n6282) );
  AOI21_X1 U5020 ( .B1(n7682), .B2(n7681), .A(n7680), .ZN(n7701) );
  OR2_X1 U5021 ( .A1(n7686), .A2(n7639), .ZN(n7692) );
  INV_X1 U5022 ( .A(n7699), .ZN(n7707) );
  AOI21_X1 U5023 ( .B1(n8690), .B2(n8830), .A(n4497), .ZN(n4496) );
  INV_X1 U5024 ( .A(n8849), .ZN(n4497) );
  AOI21_X1 U5025 ( .B1(n7720), .B2(n7660), .A(n7721), .ZN(n4540) );
  NAND2_X1 U5026 ( .A1(n7719), .A2(n7639), .ZN(n4539) );
  NOR2_X1 U5027 ( .A1(n4431), .A2(n4430), .ZN(n4429) );
  INV_X1 U5028 ( .A(n9240), .ZN(n4430) );
  INV_X1 U5029 ( .A(n8719), .ZN(n4431) );
  NAND2_X1 U5030 ( .A1(n8721), .A2(n4642), .ZN(n4428) );
  AND2_X1 U5031 ( .A1(n4532), .A2(n4375), .ZN(n4531) );
  NAND2_X1 U5032 ( .A1(n4533), .A2(n4534), .ZN(n4532) );
  AND2_X1 U5033 ( .A1(n4535), .A2(n4528), .ZN(n4527) );
  NAND2_X1 U5034 ( .A1(n4531), .A2(n4529), .ZN(n4528) );
  INV_X1 U5035 ( .A(n7787), .ZN(n4535) );
  INV_X1 U5036 ( .A(n4533), .ZN(n4529) );
  NAND2_X1 U5037 ( .A1(n8733), .A2(n8732), .ZN(n4501) );
  NOR2_X1 U5038 ( .A1(n9024), .A2(n8773), .ZN(n4500) );
  NAND2_X1 U5039 ( .A1(n4435), .A2(n8819), .ZN(n4434) );
  NAND2_X1 U5040 ( .A1(n8734), .A2(n8816), .ZN(n4435) );
  NOR2_X1 U5041 ( .A1(n8817), .A2(n8765), .ZN(n4433) );
  AOI21_X1 U5042 ( .B1(n4507), .B2(n4506), .A(n4505), .ZN(n7800) );
  NOR2_X1 U5043 ( .A1(n8422), .A2(n7660), .ZN(n4505) );
  NAND2_X1 U5044 ( .A1(n7797), .A2(n5463), .ZN(n4507) );
  NAND2_X1 U5045 ( .A1(n5255), .A2(n4351), .ZN(n4746) );
  NOR2_X1 U5046 ( .A1(n4746), .A2(n4745), .ZN(n4744) );
  INV_X1 U5047 ( .A(n5249), .ZN(n4745) );
  AND3_X1 U5048 ( .A1(n4974), .A2(n5200), .A3(n4960), .ZN(n4964) );
  AND2_X1 U5049 ( .A1(n4973), .A2(n4972), .ZN(n4586) );
  NAND2_X1 U5050 ( .A1(n9258), .A2(n8777), .ZN(n4488) );
  NAND2_X1 U5051 ( .A1(n8766), .A2(n9053), .ZN(n4491) );
  NOR2_X1 U5052 ( .A1(n9258), .A2(n8765), .ZN(n4490) );
  OR2_X1 U5053 ( .A1(n9626), .A2(n8994), .ZN(n8776) );
  NAND2_X1 U5054 ( .A1(n5530), .A2(n5528), .ZN(n4683) );
  NOR2_X1 U5055 ( .A1(n5041), .A2(n4712), .ZN(n4711) );
  INV_X1 U5056 ( .A(n5033), .ZN(n4712) );
  NAND2_X1 U5057 ( .A1(n4517), .A2(n4837), .ZN(n4516) );
  INV_X1 U5058 ( .A(n5026), .ZN(n4517) );
  INV_X1 U5059 ( .A(n4713), .ZN(n4512) );
  INV_X1 U5060 ( .A(n4839), .ZN(n4714) );
  INV_X1 U5061 ( .A(n4837), .ZN(n4518) );
  NAND2_X1 U5062 ( .A1(n4560), .A2(n4322), .ZN(n7905) );
  AND2_X1 U5063 ( .A1(n5808), .A2(n7635), .ZN(n5816) );
  XNOR2_X1 U5064 ( .A(n7926), .B(n5233), .ZN(n5815) );
  OR2_X1 U5065 ( .A1(n5455), .A2(n7931), .ZN(n5464) );
  NOR2_X1 U5066 ( .A1(n8427), .A2(n8433), .ZN(n4470) );
  OR2_X1 U5067 ( .A1(n8439), .A2(n8042), .ZN(n7780) );
  NOR2_X1 U5068 ( .A1(n8381), .A2(n8480), .ZN(n4463) );
  INV_X1 U5069 ( .A(n7755), .ZN(n7749) );
  INV_X1 U5070 ( .A(n7721), .ZN(n7834) );
  INV_X1 U5071 ( .A(n5309), .ZN(n4750) );
  OAI21_X1 U5072 ( .B1(n4751), .B2(n4750), .A(n7830), .ZN(n4749) );
  AND2_X1 U5073 ( .A1(n6734), .A2(n5300), .ZN(n4751) );
  INV_X1 U5074 ( .A(n5491), .ZN(n6734) );
  AND2_X1 U5075 ( .A1(n4816), .A2(n7683), .ZN(n6816) );
  NOR2_X1 U5076 ( .A1(n6625), .A2(n6814), .ZN(n4461) );
  INV_X1 U5077 ( .A(n6623), .ZN(n4460) );
  NAND2_X1 U5078 ( .A1(n5242), .A2(n5914), .ZN(n7655) );
  INV_X1 U5079 ( .A(n6090), .ZN(n5846) );
  AND2_X1 U5080 ( .A1(n7136), .A2(n7134), .ZN(n4673) );
  OR2_X1 U5081 ( .A1(n7478), .A2(n8568), .ZN(n7501) );
  AND2_X1 U5082 ( .A1(n7489), .A2(n7488), .ZN(n7502) );
  NOR2_X1 U5083 ( .A1(n9061), .A2(n4697), .ZN(n4696) );
  NAND2_X1 U5084 ( .A1(n4699), .A2(n4698), .ZN(n4697) );
  AND2_X1 U5085 ( .A1(n9278), .A2(n8869), .ZN(n9031) );
  AND2_X1 U5086 ( .A1(n8870), .A2(n9082), .ZN(n9032) );
  OR2_X1 U5087 ( .A1(n9278), .A2(n9103), .ZN(n9016) );
  OR2_X1 U5088 ( .A1(n9296), .A2(n9302), .ZN(n4690) );
  AND2_X1 U5089 ( .A1(n9296), .A2(n9006), .ZN(n9024) );
  OR2_X1 U5090 ( .A1(n9302), .A2(n8632), .ZN(n8816) );
  NAND2_X1 U5091 ( .A1(n9330), .A2(n8932), .ZN(n4799) );
  NAND2_X1 U5092 ( .A1(n4642), .A2(n4641), .ZN(n4640) );
  NAND2_X1 U5093 ( .A1(n4370), .A2(n8699), .ZN(n4623) );
  NAND2_X1 U5094 ( .A1(n8698), .A2(n8694), .ZN(n4625) );
  NAND2_X1 U5095 ( .A1(n8699), .A2(n8698), .ZN(n4624) );
  OR2_X1 U5096 ( .A1(n9665), .A2(n9641), .ZN(n8701) );
  NAND2_X1 U5097 ( .A1(n6930), .A2(n4388), .ZN(n9789) );
  AND2_X1 U5098 ( .A1(n5844), .A2(n9154), .ZN(n5883) );
  INV_X1 U5099 ( .A(n4645), .ZN(n4644) );
  NAND2_X1 U5100 ( .A1(n5559), .A2(n4646), .ZN(n4645) );
  NAND2_X1 U5101 ( .A1(n5641), .A2(n5533), .ZN(n5562) );
  NAND2_X1 U5102 ( .A1(n4919), .A2(n4918), .ZN(n5146) );
  NAND2_X1 U5103 ( .A1(n4614), .A2(n4612), .ZN(n4919) );
  AOI21_X1 U5104 ( .B1(n4615), .B2(n4331), .A(n4613), .ZN(n4612) );
  INV_X1 U5105 ( .A(n4875), .ZN(n4601) );
  NOR2_X1 U5106 ( .A1(n4876), .A2(n4604), .ZN(n4603) );
  INV_X1 U5107 ( .A(n4871), .ZN(n4604) );
  NAND2_X1 U5108 ( .A1(n5077), .A2(n5076), .ZN(n4872) );
  NAND2_X1 U5109 ( .A1(n4853), .A2(n4852), .ZN(n4856) );
  INV_X1 U5110 ( .A(SI_6_), .ZN(n9458) );
  OAI211_X1 U5111 ( .C1(n4829), .C2(P1_DATAO_REG_0__SCAN_IN), .A(SI_0_), .B(
        n4508), .ZN(n4824) );
  NAND2_X1 U5112 ( .A1(n4829), .A2(n4509), .ZN(n4508) );
  NAND2_X1 U5113 ( .A1(n5265), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5274) );
  AOI21_X1 U5114 ( .B1(n8028), .B2(n8027), .A(n7887), .ZN(n7954) );
  AND2_X1 U5115 ( .A1(n7986), .A2(n7874), .ZN(n7979) );
  OR2_X1 U5116 ( .A1(n5350), .A2(n9444), .ZN(n5359) );
  NAND2_X1 U5117 ( .A1(n4542), .A2(n4541), .ZN(n6245) );
  AND2_X1 U5118 ( .A1(n6198), .A2(n6192), .ZN(n4541) );
  AOI21_X1 U5119 ( .B1(n6639), .B2(n6638), .A(n6637), .ZN(n6646) );
  OR2_X1 U5120 ( .A1(n5281), .A2(n9557), .ZN(n5292) );
  NOR2_X1 U5121 ( .A1(n6914), .A2(n6906), .ZN(n4812) );
  OR2_X1 U5122 ( .A1(n7866), .A2(n4572), .ZN(n4571) );
  INV_X1 U5123 ( .A(n7867), .ZN(n4572) );
  NOR2_X1 U5124 ( .A1(n7882), .A2(n7881), .ZN(n4809) );
  OR2_X1 U5125 ( .A1(n5366), .A2(n9454), .ZN(n5377) );
  NAND2_X1 U5126 ( .A1(n4555), .A2(n7916), .ZN(n4554) );
  INV_X1 U5127 ( .A(n7971), .ZN(n4555) );
  AND2_X1 U5128 ( .A1(n8040), .A2(n4551), .ZN(n4550) );
  NAND2_X1 U5129 ( .A1(n4552), .A2(n4554), .ZN(n4551) );
  INV_X1 U5130 ( .A(n4556), .ZN(n4552) );
  INV_X1 U5131 ( .A(n4554), .ZN(n4553) );
  NAND2_X1 U5132 ( .A1(n7915), .A2(n7914), .ZN(n7917) );
  AND2_X1 U5133 ( .A1(n7910), .A2(n7909), .ZN(n7915) );
  OAI21_X1 U5134 ( .B1(n8156), .B2(n4702), .A(n4701), .ZN(n4700) );
  NAND2_X1 U5135 ( .A1(n4707), .A2(n7810), .ZN(n4702) );
  OAI21_X1 U5136 ( .B1(n4705), .B2(n4704), .A(n4395), .ZN(n4703) );
  NOR2_X1 U5137 ( .A1(n7815), .A2(n4522), .ZN(n4521) );
  INV_X1 U5138 ( .A(n7812), .ZN(n4522) );
  NAND2_X1 U5139 ( .A1(n7862), .A2(n9946), .ZN(n7850) );
  AOI21_X1 U5140 ( .B1(n4321), .B2(n4524), .A(n7851), .ZN(n4523) );
  AND2_X1 U5141 ( .A1(n8219), .A2(n4466), .ZN(n8147) );
  AND2_X1 U5142 ( .A1(n4468), .A2(n4467), .ZN(n4466) );
  NAND2_X1 U5143 ( .A1(n8219), .A2(n4468), .ZN(n8163) );
  NAND2_X1 U5144 ( .A1(n8156), .A2(n8155), .ZN(n8154) );
  OR2_X1 U5145 ( .A1(n8191), .A2(n8189), .ZN(n5444) );
  OR2_X1 U5146 ( .A1(n5416), .A2(n8005), .ZN(n5425) );
  OR2_X1 U5147 ( .A1(n8442), .A2(n8248), .ZN(n8214) );
  AND2_X1 U5148 ( .A1(n5403), .A2(n5402), .ZN(n8247) );
  NAND2_X1 U5149 ( .A1(n8310), .A2(n4444), .ZN(n4443) );
  NOR2_X1 U5150 ( .A1(n8292), .A2(n7759), .ZN(n4444) );
  INV_X1 U5151 ( .A(n8265), .ZN(n8273) );
  AND2_X1 U5152 ( .A1(n7768), .A2(n7769), .ZN(n8265) );
  NAND2_X1 U5153 ( .A1(n5388), .A2(n5387), .ZN(n8293) );
  AND3_X1 U5154 ( .A1(n5394), .A2(n5393), .A3(n5392), .ZN(n8308) );
  NAND2_X1 U5155 ( .A1(n5504), .A2(n4721), .ZN(n8310) );
  AND2_X1 U5156 ( .A1(n7841), .A2(n7750), .ZN(n4721) );
  INV_X1 U5157 ( .A(n5373), .ZN(n4739) );
  AND2_X1 U5158 ( .A1(n4737), .A2(n5374), .ZN(n4736) );
  NAND2_X1 U5159 ( .A1(n5373), .A2(n4738), .ZN(n4737) );
  INV_X1 U5160 ( .A(n5365), .ZN(n4738) );
  INV_X1 U5161 ( .A(n7838), .ZN(n8323) );
  NOR2_X1 U5162 ( .A1(n8334), .A2(n8471), .ZN(n8315) );
  NAND2_X1 U5163 ( .A1(n8348), .A2(n4356), .ZN(n8338) );
  INV_X1 U5164 ( .A(n7732), .ZN(n8352) );
  INV_X1 U5165 ( .A(n5334), .ZN(n5333) );
  NAND2_X1 U5166 ( .A1(n6781), .A2(n4751), .ZN(n6728) );
  NOR2_X1 U5167 ( .A1(n6787), .A2(n5308), .ZN(n6952) );
  OR2_X1 U5168 ( .A1(n5487), .A2(n5486), .ZN(n5488) );
  NAND2_X1 U5169 ( .A1(n9988), .A2(n6246), .ZN(n6615) );
  NAND2_X1 U5170 ( .A1(n6460), .A2(n5264), .ZN(n7646) );
  NAND2_X1 U5171 ( .A1(n6131), .A2(n6130), .ZN(n6129) );
  AND2_X1 U5172 ( .A1(n5822), .A2(n5507), .ZN(n8390) );
  INV_X1 U5173 ( .A(n8307), .ZN(n8392) );
  NAND2_X1 U5174 ( .A1(n5105), .A2(n5104), .ZN(n8484) );
  INV_X1 U5175 ( .A(n6206), .ZN(n9981) );
  AND2_X2 U5176 ( .A1(n9964), .A2(n7818), .ZN(n8499) );
  AND2_X1 U5177 ( .A1(n5218), .A2(n6543), .ZN(n9964) );
  XNOR2_X1 U5178 ( .A(n4981), .B(P2_IR_REG_30__SCAN_IN), .ZN(n5224) );
  OR2_X1 U5179 ( .A1(n4988), .A2(n4982), .ZN(n4981) );
  NOR2_X1 U5180 ( .A1(n4989), .A2(n4988), .ZN(n5223) );
  XNOR2_X1 U5181 ( .A(n4966), .B(n4965), .ZN(n4993) );
  NOR2_X1 U5182 ( .A1(n5019), .A2(n4576), .ZN(n4575) );
  NAND2_X1 U5183 ( .A1(n4577), .A2(n4959), .ZN(n4576) );
  AND2_X1 U5184 ( .A1(n5030), .A2(n5031), .ZN(n5039) );
  NOR2_X1 U5185 ( .A1(n5019), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n5030) );
  NOR2_X1 U5186 ( .A1(n7242), .A2(n4672), .ZN(n4671) );
  INV_X1 U5187 ( .A(n7166), .ZN(n4672) );
  INV_X1 U5188 ( .A(n4673), .ZN(n4669) );
  NAND2_X1 U5189 ( .A1(n8640), .A2(n8639), .ZN(n4665) );
  OR2_X1 U5190 ( .A1(n8640), .A2(n8639), .ZN(n4666) );
  OR2_X1 U5191 ( .A1(n8585), .A2(n8583), .ZN(n8582) );
  NAND2_X1 U5192 ( .A1(n7509), .A2(n7508), .ZN(n8548) );
  NAND2_X1 U5193 ( .A1(n4680), .A2(n4679), .ZN(n6828) );
  AND2_X1 U5194 ( .A1(n6762), .A2(n6761), .ZN(n4679) );
  OR2_X1 U5195 ( .A1(n7368), .A2(n8631), .ZN(n7385) );
  NAND2_X1 U5196 ( .A1(n4659), .A2(n4656), .ZN(n8594) );
  NOR2_X1 U5197 ( .A1(n4660), .A2(n4657), .ZN(n4656) );
  NOR2_X1 U5198 ( .A1(n4658), .A2(n7443), .ZN(n4657) );
  NAND2_X1 U5199 ( .A1(n4589), .A2(n4484), .ZN(n8884) );
  NAND2_X1 U5200 ( .A1(n4437), .A2(n8765), .ZN(n4589) );
  AOI21_X1 U5201 ( .B1(n4486), .B2(n4590), .A(n4485), .ZN(n4484) );
  OAI21_X1 U5202 ( .B1(n8766), .B2(n4438), .A(n8879), .ZN(n4437) );
  AND4_X1 U5203 ( .A1(n7413), .A2(n7412), .A3(n7411), .A4(n7410), .ZN(n8758)
         );
  NAND2_X1 U5204 ( .A1(n6167), .A2(n4347), .ZN(n9698) );
  NAND2_X1 U5205 ( .A1(n9722), .A2(n4474), .ZN(n9732) );
  NAND2_X1 U5206 ( .A1(n4475), .A2(n6083), .ZN(n4474) );
  OR2_X1 U5207 ( .A1(n9732), .A2(n9733), .ZN(n4473) );
  NOR2_X1 U5208 ( .A1(n9763), .A2(n4480), .ZN(n9777) );
  AND2_X1 U5209 ( .A1(n9757), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n4480) );
  OR2_X1 U5210 ( .A1(n9777), .A2(n9776), .ZN(n4479) );
  OR2_X1 U5211 ( .A1(n6538), .A2(n6539), .ZN(n4481) );
  AND2_X1 U5212 ( .A1(n6155), .A2(n6156), .ZN(n6707) );
  OR2_X1 U5213 ( .A1(n7148), .A2(n7147), .ZN(n4477) );
  NAND2_X1 U5214 ( .A1(n8764), .A2(n8763), .ZN(n8992) );
  NAND2_X1 U5215 ( .A1(n8770), .A2(n8769), .ZN(n9042) );
  AOI21_X1 U5216 ( .B1(n4630), .B2(n4325), .A(n9242), .ZN(n4627) );
  NAND2_X1 U5217 ( .A1(n4630), .A2(n4634), .ZN(n4629) );
  NAND2_X1 U5218 ( .A1(n9035), .A2(n9034), .ZN(n4634) );
  AND2_X1 U5219 ( .A1(n9034), .A2(n8809), .ZN(n9051) );
  INV_X1 U5220 ( .A(n4647), .ZN(n9074) );
  OAI21_X1 U5221 ( .B1(n9112), .B2(n4649), .A(n4648), .ZN(n4647) );
  AOI21_X1 U5222 ( .B1(n9032), .B2(n4651), .A(n9031), .ZN(n4648) );
  NAND2_X1 U5223 ( .A1(n9032), .A2(n4650), .ZN(n4649) );
  OR2_X1 U5224 ( .A1(n9095), .A2(n9278), .ZN(n9086) );
  NOR2_X1 U5225 ( .A1(n9086), .A2(n9271), .ZN(n9068) );
  AND2_X1 U5226 ( .A1(n9033), .A2(n8808), .ZN(n9073) );
  AOI21_X1 U5227 ( .B1(n4774), .B2(n4777), .A(n4772), .ZN(n4771) );
  INV_X1 U5228 ( .A(n9017), .ZN(n4772) );
  NAND2_X1 U5229 ( .A1(n9028), .A2(n9030), .ZN(n4651) );
  AND4_X1 U5230 ( .A1(n7586), .A2(n7585), .A3(n7584), .A4(n7583), .ZN(n9085)
         );
  AND2_X1 U5231 ( .A1(n4781), .A2(n9014), .ZN(n4780) );
  NAND2_X1 U5232 ( .A1(n4779), .A2(n4781), .ZN(n4778) );
  INV_X1 U5233 ( .A(n9101), .ZN(n4779) );
  AND2_X1 U5234 ( .A1(n9126), .A2(n9008), .ZN(n9009) );
  OR2_X1 U5235 ( .A1(n9306), .A2(n9179), .ZN(n9144) );
  INV_X1 U5236 ( .A(n4769), .ZN(n4768) );
  OAI21_X1 U5237 ( .B1(n4386), .B2(n7349), .A(n7361), .ZN(n4769) );
  OR2_X1 U5238 ( .A1(n9180), .A2(n9306), .ZN(n9160) );
  NAND2_X1 U5239 ( .A1(n9316), .A2(n7336), .ZN(n9173) );
  AOI21_X1 U5240 ( .B1(n9206), .B2(n7331), .A(n7330), .ZN(n9196) );
  NOR2_X1 U5241 ( .A1(n9222), .A2(n9325), .ZN(n9207) );
  NAND2_X1 U5242 ( .A1(n4639), .A2(n4640), .ZN(n9230) );
  NOR2_X1 U5243 ( .A1(n7307), .A2(n4798), .ZN(n4797) );
  INV_X1 U5244 ( .A(n4800), .ZN(n4798) );
  NOR2_X1 U5245 ( .A1(n7307), .A2(n4796), .ZN(n4795) );
  NAND2_X1 U5246 ( .A1(n4800), .A2(n7301), .ZN(n4796) );
  NAND2_X1 U5247 ( .A1(n7300), .A2(n9243), .ZN(n4800) );
  NOR2_X1 U5248 ( .A1(n7300), .A2(n9243), .ZN(n7301) );
  NAND2_X1 U5249 ( .A1(n7214), .A2(n4810), .ZN(n7256) );
  OR2_X1 U5250 ( .A1(n7213), .A2(n9641), .ZN(n4810) );
  NAND2_X1 U5251 ( .A1(n7068), .A2(n7067), .ZN(n9634) );
  NAND2_X1 U5252 ( .A1(n7094), .A2(n8850), .ZN(n9640) );
  NAND2_X1 U5253 ( .A1(n6933), .A2(n6937), .ZN(n7068) );
  NAND2_X1 U5254 ( .A1(n6508), .A2(n4762), .ZN(n6658) );
  NAND2_X1 U5255 ( .A1(n6567), .A2(n4763), .ZN(n4762) );
  INV_X1 U5256 ( .A(n9827), .ZN(n4763) );
  AND3_X1 U5257 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n6321) );
  AND2_X1 U5258 ( .A1(n6010), .A2(n8925), .ZN(n9825) );
  NAND2_X1 U5259 ( .A1(n6030), .A2(n4692), .ZN(n4693) );
  OAI22_X1 U5260 ( .A1(n5917), .A2(n5918), .B1(n5919), .B2(n4595), .ZN(n4692)
         );
  INV_X1 U5261 ( .A(n9825), .ZN(n9802) );
  OR2_X1 U5262 ( .A1(n8805), .A2(n8925), .ZN(n9800) );
  INV_X1 U5263 ( .A(n9800), .ZN(n9828) );
  NOR2_X1 U5264 ( .A1(n5558), .A2(n4498), .ZN(n5560) );
  NAND2_X1 U5265 ( .A1(n5556), .A2(n5559), .ZN(n4498) );
  OR2_X1 U5266 ( .A1(n5171), .A2(n9551), .ZN(n4942) );
  XNOR2_X1 U5267 ( .A(n5175), .B(n5174), .ZN(n8677) );
  NAND2_X1 U5268 ( .A1(n4605), .A2(n4936), .ZN(n5166) );
  XNOR2_X1 U5269 ( .A(n5162), .B(n5161), .ZN(n7575) );
  AND2_X1 U5270 ( .A1(n4932), .A2(n5155), .ZN(n5162) );
  XNOR2_X1 U5271 ( .A(n5158), .B(n5157), .ZN(n7547) );
  NAND2_X1 U5272 ( .A1(n5154), .A2(n5153), .ZN(n5158) );
  NAND2_X1 U5273 ( .A1(n4618), .A2(n4909), .ZN(n5138) );
  XNOR2_X1 U5274 ( .A(n5125), .B(n5124), .ZN(n7337) );
  XNOR2_X1 U5275 ( .A(n5113), .B(n5106), .ZN(n7318) );
  INV_X1 U5276 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5791) );
  NAND2_X1 U5277 ( .A1(n4609), .A2(n4860), .ZN(n5070) );
  NAND2_X1 U5278 ( .A1(n4857), .A2(n4610), .ZN(n4609) );
  NAND2_X1 U5279 ( .A1(n4311), .A2(n4334), .ZN(n4502) );
  NAND2_X1 U5280 ( .A1(n5092), .A2(n5091), .ZN(n8497) );
  NAND2_X1 U5281 ( .A1(n5144), .A2(n5143), .ZN(n8448) );
  NAND2_X1 U5282 ( .A1(n5136), .A2(n5135), .ZN(n8459) );
  INV_X1 U5283 ( .A(n8302), .ZN(n8464) );
  NAND2_X1 U5284 ( .A1(n5081), .A2(n5080), .ZN(n8505) );
  NAND2_X1 U5285 ( .A1(n5099), .A2(n5098), .ZN(n8492) );
  OAI21_X1 U5286 ( .B1(n9606), .B2(n5689), .A(n4405), .ZN(n9609) );
  NAND2_X1 U5287 ( .A1(n9606), .A2(n5689), .ZN(n4405) );
  XNOR2_X1 U5288 ( .A(n4406), .B(P2_IR_REG_1__SCAN_IN), .ZN(n9606) );
  NAND2_X1 U5289 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n4406) );
  NAND2_X1 U5290 ( .A1(n9622), .A2(n9621), .ZN(n9620) );
  NAND2_X1 U5291 ( .A1(n5747), .A2(n4387), .ZN(n5764) );
  NAND2_X1 U5292 ( .A1(n8081), .A2(n5767), .ZN(n8099) );
  NAND2_X1 U5293 ( .A1(n8099), .A2(n8098), .ZN(n8097) );
  NAND2_X1 U5294 ( .A1(n6112), .A2(n4389), .ZN(n6115) );
  NAND2_X1 U5295 ( .A1(n8110), .A2(n8109), .ZN(n8120) );
  NAND2_X1 U5296 ( .A1(n4970), .A2(n4969), .ZN(n7631) );
  NAND2_X1 U5297 ( .A1(n4724), .A2(n4723), .ZN(n5473) );
  AOI21_X1 U5298 ( .B1(n4727), .B2(n4323), .A(n4361), .ZN(n4723) );
  NAND2_X1 U5299 ( .A1(n8651), .A2(n7574), .ZN(n8540) );
  AND4_X1 U5300 ( .A1(n7093), .A2(n7092), .A3(n7091), .A4(n7090), .ZN(n7248)
         );
  NAND2_X1 U5301 ( .A1(n7529), .A2(n7528), .ZN(n9281) );
  INV_X1 U5302 ( .A(n9007), .ZN(n9296) );
  AND2_X1 U5303 ( .A1(n7537), .A2(n7536), .ZN(n9116) );
  NAND2_X1 U5304 ( .A1(n7306), .A2(n7305), .ZN(n9335) );
  OR2_X1 U5305 ( .A1(n4425), .A2(n4382), .ZN(n4422) );
  NOR2_X1 U5306 ( .A1(n8884), .A2(n4423), .ZN(n4421) );
  OR2_X1 U5307 ( .A1(n8805), .A2(n9154), .ZN(n4423) );
  INV_X1 U5308 ( .A(n8929), .ZN(n4424) );
  INV_X1 U5309 ( .A(n8928), .ZN(n4420) );
  INV_X1 U5310 ( .A(n8758), .ZN(n9075) );
  OR2_X1 U5311 ( .A1(n5933), .A2(n6264), .ZN(n5935) );
  NAND2_X1 U5312 ( .A1(n5931), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5937) );
  OR2_X1 U5313 ( .A1(n5933), .A2(n6176), .ZN(n5879) );
  OR2_X1 U5314 ( .A1(n7598), .A2(n5666), .ZN(n5667) );
  OR2_X1 U5315 ( .A1(n5933), .A2(n5665), .ZN(n5668) );
  INV_X1 U5316 ( .A(n6030), .ZN(n9688) );
  OAI21_X1 U5317 ( .B1(n6160), .B2(P1_REG2_REG_3__SCAN_IN), .A(n4471), .ZN(
        n6169) );
  NAND2_X1 U5318 ( .A1(n6168), .A2(n6169), .ZN(n6167) );
  NAND2_X1 U5319 ( .A1(n7661), .A2(n7660), .ZN(n7662) );
  NAND2_X1 U5320 ( .A1(n7643), .A2(n7642), .ZN(n7676) );
  NAND2_X1 U5321 ( .A1(n7640), .A2(n7639), .ZN(n7643) );
  MUX2_X1 U5322 ( .A(n7709), .B(n7708), .S(n7660), .Z(n7710) );
  NAND2_X1 U5323 ( .A1(n8700), .A2(n4494), .ZN(n8702) );
  OAI21_X1 U5324 ( .B1(n4496), .B2(n8826), .A(n4495), .ZN(n4494) );
  NOR2_X1 U5325 ( .A1(n8709), .A2(n4339), .ZN(n4495) );
  AOI21_X1 U5326 ( .B1(n4538), .B2(n4536), .A(n4359), .ZN(n7742) );
  NOR2_X1 U5327 ( .A1(n7833), .A2(n4537), .ZN(n4536) );
  NAND2_X1 U5328 ( .A1(n4540), .A2(n4539), .ZN(n4538) );
  OAI21_X1 U5329 ( .B1(n4427), .B2(n4426), .A(n8723), .ZN(n8727) );
  NAND2_X1 U5330 ( .A1(n8722), .A2(n9214), .ZN(n4426) );
  AOI21_X1 U5331 ( .B1(n8720), .B2(n4429), .A(n4428), .ZN(n4427) );
  INV_X1 U5332 ( .A(n7777), .ZN(n4534) );
  AOI21_X1 U5333 ( .B1(n4326), .B2(n7777), .A(n4369), .ZN(n4533) );
  AOI21_X1 U5334 ( .B1(n4527), .B2(n4530), .A(n4365), .ZN(n4526) );
  INV_X1 U5335 ( .A(n4531), .ZN(n4530) );
  AOI21_X1 U5336 ( .B1(n4499), .B2(n4432), .A(n8742), .ZN(n8752) );
  AOI21_X1 U5337 ( .B1(n4434), .B2(n4433), .A(n8741), .ZN(n4432) );
  NAND2_X1 U5338 ( .A1(n4501), .A2(n4500), .ZN(n4499) );
  NAND2_X1 U5339 ( .A1(n8695), .A2(n8716), .ZN(n8858) );
  AND2_X1 U5340 ( .A1(n8778), .A2(n9027), .ZN(n8740) );
  NOR2_X1 U5341 ( .A1(n4385), .A2(n4559), .ZN(n4558) );
  INV_X1 U5342 ( .A(n7893), .ZN(n4559) );
  OR2_X1 U5343 ( .A1(n7631), .A2(n7630), .ZN(n7814) );
  AND2_X1 U5344 ( .A1(n8474), .A2(n7956), .ZN(n7755) );
  NOR2_X1 U5345 ( .A1(n6975), .A2(n6682), .ZN(n7689) );
  OR2_X1 U5346 ( .A1(n7826), .A2(n7646), .ZN(n5485) );
  INV_X1 U5347 ( .A(n5141), .ZN(n4613) );
  INV_X1 U5348 ( .A(n5100), .ZN(n4597) );
  INV_X1 U5349 ( .A(n4860), .ZN(n4608) );
  NAND2_X1 U5350 ( .A1(n4861), .A2(n9469), .ZN(n4864) );
  NAND2_X1 U5351 ( .A1(n4842), .A2(n9562), .ZN(n4845) );
  INV_X1 U5352 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4440) );
  AOI21_X1 U5353 ( .B1(n4707), .B2(n4726), .A(n7796), .ZN(n4705) );
  AND2_X1 U5354 ( .A1(n7814), .A2(n7804), .ZN(n7809) );
  INV_X1 U5355 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n4954) );
  OR2_X1 U5356 ( .A1(n8416), .A2(n8158), .ZN(n7801) );
  AND2_X1 U5357 ( .A1(n4470), .A2(n4469), .ZN(n4468) );
  OR2_X1 U5358 ( .A1(n8433), .A2(n8181), .ZN(n7784) );
  AND2_X1 U5359 ( .A1(n4736), .A2(n4338), .ZN(n4735) );
  AND2_X1 U5360 ( .A1(n7751), .A2(n7761), .ZN(n7841) );
  AND2_X1 U5361 ( .A1(n7734), .A2(n7737), .ZN(n7732) );
  OR2_X1 U5362 ( .A1(n5302), .A2(n9540), .ZN(n5312) );
  NAND2_X1 U5363 ( .A1(n4742), .A2(n8065), .ZN(n4741) );
  INV_X1 U5364 ( .A(n7824), .ZN(n4742) );
  AND2_X1 U5365 ( .A1(n9981), .A2(n7670), .ZN(n4465) );
  INV_X1 U5366 ( .A(n6234), .ZN(n4464) );
  AND2_X1 U5367 ( .A1(n5483), .A2(n6615), .ZN(n7826) );
  NAND2_X1 U5368 ( .A1(n7672), .A2(n7674), .ZN(n7640) );
  AND2_X1 U5369 ( .A1(n8232), .A2(n8224), .ZN(n8219) );
  NAND2_X1 U5370 ( .A1(n4464), .A2(n4465), .ZN(n6691) );
  NOR2_X1 U5371 ( .A1(n6234), .A2(n6495), .ZN(n6236) );
  NOR2_X1 U5372 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_26__SCAN_IN), .ZN(
        n4963) );
  NAND2_X1 U5373 ( .A1(n4367), .A2(n4960), .ZN(n5190) );
  NAND2_X1 U5374 ( .A1(n4960), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4585) );
  AND2_X1 U5375 ( .A1(n4586), .A2(P2_IR_REG_21__SCAN_IN), .ZN(n4583) );
  AND2_X1 U5376 ( .A1(n4579), .A2(n4578), .ZN(n4577) );
  INV_X1 U5377 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n4579) );
  INV_X1 U5378 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n4578) );
  NAND2_X1 U5379 ( .A1(n4371), .A2(n4665), .ZN(n4664) );
  INV_X1 U5380 ( .A(n8596), .ZN(n4660) );
  INV_X1 U5381 ( .A(n7566), .ZN(n7590) );
  OR2_X1 U5382 ( .A1(n8875), .A2(n8777), .ZN(n4438) );
  NAND2_X1 U5383 ( .A1(n4491), .A2(n4490), .ZN(n4489) );
  OR2_X1 U5384 ( .A1(n8766), .A2(n4488), .ZN(n4487) );
  NAND2_X1 U5385 ( .A1(n4592), .A2(n8877), .ZN(n4485) );
  OR2_X1 U5386 ( .A1(n8771), .A2(n4593), .ZN(n4592) );
  OR2_X1 U5387 ( .A1(n9042), .A2(n8777), .ZN(n8874) );
  AND2_X1 U5388 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(n7581), .ZN(n7407) );
  INV_X1 U5389 ( .A(n9113), .ZN(n4650) );
  AOI21_X1 U5390 ( .B1(n4778), .B2(n4776), .A(n4775), .ZN(n4774) );
  INV_X1 U5391 ( .A(n4780), .ZN(n4776) );
  INV_X1 U5392 ( .A(n9016), .ZN(n4775) );
  INV_X1 U5393 ( .A(n4778), .ZN(n4777) );
  OR2_X1 U5394 ( .A1(n9291), .A2(n4690), .ZN(n4689) );
  NOR2_X1 U5395 ( .A1(n4386), .A2(n4766), .ZN(n4765) );
  INV_X1 U5396 ( .A(n7336), .ZN(n4766) );
  NAND2_X1 U5397 ( .A1(n9318), .A2(n9217), .ZN(n8825) );
  NAND2_X1 U5398 ( .A1(n9253), .A2(n4688), .ZN(n4687) );
  NOR2_X1 U5399 ( .A1(n9339), .A2(n7268), .ZN(n4688) );
  NAND2_X1 U5400 ( .A1(n7300), .A2(n4439), .ZN(n8716) );
  OAI21_X1 U5401 ( .B1(n6510), .B2(n4492), .A(n8838), .ZN(n8687) );
  NAND2_X1 U5402 ( .A1(n4493), .A2(n6513), .ZN(n4492) );
  AND2_X1 U5403 ( .A1(n6511), .A2(n9819), .ZN(n4493) );
  NOR2_X1 U5404 ( .A1(n6403), .A2(n6402), .ZN(n6425) );
  OR2_X1 U5405 ( .A1(n9637), .A2(n9665), .ZN(n7263) );
  NAND2_X1 U5406 ( .A1(n9834), .A2(n4318), .ZN(n6662) );
  NAND2_X1 U5407 ( .A1(n5154), .A2(n4929), .ZN(n4932) );
  NOR2_X1 U5408 ( .A1(n5132), .A2(n4620), .ZN(n4619) );
  INV_X1 U5409 ( .A(n4906), .ZN(n4620) );
  NAND2_X1 U5410 ( .A1(n4677), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4676) );
  INV_X1 U5411 ( .A(n5113), .ZN(n4891) );
  AND3_X1 U5412 ( .A1(n5586), .A2(n5527), .A3(n4682), .ZN(n5945) );
  NOR2_X1 U5413 ( .A1(n4683), .A2(n5540), .ZN(n4682) );
  NAND2_X1 U5414 ( .A1(n5791), .A2(n5661), .ZN(n5540) );
  INV_X1 U5415 ( .A(n4683), .ZN(n4681) );
  NOR2_X1 U5416 ( .A1(n4858), .A2(n4611), .ZN(n4610) );
  INV_X1 U5417 ( .A(n4856), .ZN(n4611) );
  AND2_X1 U5418 ( .A1(n4850), .A2(n4849), .ZN(n5052) );
  NAND2_X1 U5419 ( .A1(n4513), .A2(n4511), .ZN(n5049) );
  NAND2_X1 U5420 ( .A1(n5523), .A2(n4760), .ZN(n4759) );
  INV_X1 U5421 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n4760) );
  INV_X1 U5422 ( .A(SI_3_), .ZN(n9464) );
  INV_X1 U5423 ( .A(SI_4_), .ZN(n9533) );
  AND2_X1 U5424 ( .A1(n4812), .A2(n4566), .ZN(n4563) );
  NAND2_X1 U5425 ( .A1(n8017), .A2(n7906), .ZN(n7911) );
  OR2_X1 U5426 ( .A1(n6893), .A2(n6892), .ZN(n6898) );
  NAND2_X1 U5427 ( .A1(n7868), .A2(n4571), .ZN(n4567) );
  AND2_X1 U5428 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5256) );
  NAND2_X1 U5429 ( .A1(n5256), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5266) );
  NOR2_X1 U5430 ( .A1(n7911), .A2(n4805), .ZN(n7997) );
  NAND2_X1 U5431 ( .A1(n6219), .A2(n6218), .ZN(n4542) );
  NAND2_X1 U5432 ( .A1(n7954), .A2(n7953), .ZN(n7952) );
  NAND2_X1 U5433 ( .A1(n8019), .A2(n8018), .ZN(n8017) );
  OR2_X1 U5434 ( .A1(n5396), .A2(n8021), .ZN(n5407) );
  NAND2_X1 U5435 ( .A1(n6211), .A2(n4545), .ZN(n4544) );
  NAND2_X1 U5436 ( .A1(n5814), .A2(n5813), .ZN(n4546) );
  INV_X1 U5437 ( .A(n5359), .ZN(n5357) );
  NAND2_X1 U5438 ( .A1(n7971), .A2(n4557), .ZN(n4556) );
  AND2_X1 U5439 ( .A1(n7862), .A2(n7852), .ZN(n5822) );
  INV_X1 U5440 ( .A(n7809), .ZN(n7848) );
  INV_X1 U5441 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n9557) );
  OR2_X1 U5442 ( .A1(n5060), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n5065) );
  NOR2_X1 U5443 ( .A1(n6877), .A2(n6878), .ZN(n6882) );
  NAND2_X1 U5444 ( .A1(n6882), .A2(n6881), .ZN(n8105) );
  NAND2_X1 U5445 ( .A1(n8154), .A2(n4506), .ZN(n7625) );
  NAND2_X1 U5446 ( .A1(n7801), .A2(n7802), .ZN(n7846) );
  AND2_X1 U5447 ( .A1(n5464), .A2(n5456), .ZN(n8164) );
  AND2_X1 U5448 ( .A1(n5454), .A2(n5453), .ZN(n8157) );
  OR2_X1 U5449 ( .A1(n8175), .A2(n4312), .ZN(n5454) );
  NAND2_X1 U5450 ( .A1(n8197), .A2(n4349), .ZN(n8184) );
  NAND2_X1 U5451 ( .A1(n8197), .A2(n7785), .ZN(n8180) );
  NAND2_X1 U5452 ( .A1(n8219), .A2(n4470), .ZN(n8173) );
  NAND2_X1 U5453 ( .A1(n8219), .A2(n8204), .ZN(n8206) );
  OR2_X1 U5454 ( .A1(n5425), .A2(n9479), .ZN(n5433) );
  NAND2_X1 U5455 ( .A1(n8244), .A2(n4354), .ZN(n8215) );
  NOR2_X1 U5456 ( .A1(n8253), .A2(n8442), .ZN(n8232) );
  AND2_X1 U5457 ( .A1(n5423), .A2(n5422), .ZN(n8248) );
  AND2_X1 U5458 ( .A1(n8277), .A2(n7768), .ZN(n8245) );
  AND2_X1 U5459 ( .A1(n8285), .A2(n8291), .ZN(n8287) );
  INV_X1 U5460 ( .A(n7839), .ZN(n8292) );
  INV_X1 U5461 ( .A(n7756), .ZN(n7750) );
  AND2_X1 U5462 ( .A1(n7818), .A2(n7852), .ZN(n5810) );
  NAND2_X1 U5463 ( .A1(n4463), .A2(n4462), .ZN(n8334) );
  INV_X1 U5464 ( .A(n4463), .ZN(n8360) );
  AND2_X1 U5465 ( .A1(n8399), .A2(n8407), .ZN(n8400) );
  NAND2_X1 U5466 ( .A1(n5342), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5350) );
  NOR2_X1 U5467 ( .A1(n7035), .A2(n8497), .ZN(n8399) );
  OR2_X1 U5468 ( .A1(n7033), .A2(n8505), .ZN(n7035) );
  OR2_X1 U5469 ( .A1(n5327), .A2(n5326), .ZN(n5334) );
  NAND2_X1 U5470 ( .A1(n5310), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5320) );
  INV_X1 U5471 ( .A(n5312), .ZN(n5310) );
  OR2_X1 U5472 ( .A1(n5320), .A2(n9531), .ZN(n5327) );
  OAI21_X1 U5473 ( .B1(n6781), .B2(n4750), .A(n4748), .ZN(n5319) );
  INV_X1 U5474 ( .A(n4749), .ZN(n4748) );
  AND2_X1 U5475 ( .A1(n6952), .A2(n6986), .ZN(n6953) );
  AOI21_X1 U5476 ( .B1(n5491), .B2(n7696), .A(n5492), .ZN(n5495) );
  AND2_X1 U5477 ( .A1(n6781), .A2(n5300), .ZN(n6729) );
  NOR2_X1 U5478 ( .A1(n6975), .A2(n4459), .ZN(n4458) );
  INV_X1 U5479 ( .A(n4461), .ZN(n4459) );
  NAND2_X1 U5480 ( .A1(n4460), .A2(n4461), .ZN(n6812) );
  NOR2_X1 U5481 ( .A1(n6623), .A2(n6625), .ZN(n6810) );
  OR2_X1 U5482 ( .A1(n6692), .A2(n6472), .ZN(n6623) );
  AND2_X1 U5483 ( .A1(n7645), .A2(n7672), .ZN(n7822) );
  AOI21_X1 U5484 ( .B1(n6229), .B2(n7821), .A(n5482), .ZN(n6134) );
  NAND2_X1 U5485 ( .A1(n6226), .A2(n5249), .ZN(n6131) );
  NAND2_X1 U5486 ( .A1(n5808), .A2(n5234), .ZN(n7654) );
  OR2_X1 U5487 ( .A1(n5682), .A2(n5581), .ZN(n4450) );
  OR2_X1 U5488 ( .A1(n5035), .A2(n5917), .ZN(n4451) );
  NOR2_X1 U5489 ( .A1(n5233), .A2(n9963), .ZN(n5894) );
  NAND2_X1 U5490 ( .A1(n5140), .A2(n5139), .ZN(n8454) );
  AND3_X1 U5491 ( .A1(n5008), .A2(n5007), .A3(n5006), .ZN(n9975) );
  NAND2_X1 U5492 ( .A1(n5107), .A2(n4752), .ZN(n5193) );
  NAND2_X1 U5493 ( .A1(n5190), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5201) );
  INV_X1 U5494 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n4953) );
  NOR2_X2 U5495 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n4740) );
  NOR2_X2 U5496 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5003) );
  INV_X1 U5497 ( .A(n7552), .ZN(n7581) );
  INV_X1 U5498 ( .A(n8607), .ZN(n7522) );
  NAND2_X1 U5499 ( .A1(n6757), .A2(n6756), .ZN(n4680) );
  OR2_X1 U5500 ( .A1(n7485), .A2(n7500), .ZN(n7486) );
  NOR2_X1 U5501 ( .A1(n7178), .A2(n7177), .ZN(n7223) );
  NAND2_X1 U5502 ( .A1(n4678), .A2(n5848), .ZN(n4677) );
  INV_X1 U5503 ( .A(n5543), .ZN(n4678) );
  AND3_X1 U5504 ( .A1(n7373), .A2(n7372), .A3(n7371), .ZN(n8632) );
  AND4_X1 U5505 ( .A1(n6596), .A2(n6595), .A3(n6594), .A4(n6593), .ZN(n6936)
         );
  INV_X1 U5506 ( .A(n5933), .ZN(n7554) );
  OR2_X1 U5507 ( .A1(n4316), .A2(n5878), .ZN(n4756) );
  NOR2_X1 U5508 ( .A1(n6707), .A2(n4393), .ZN(n6963) );
  AND2_X1 U5509 ( .A1(n4477), .A2(n4476), .ZN(n8955) );
  NAND2_X1 U5510 ( .A1(n8952), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n4476) );
  NOR2_X1 U5511 ( .A1(n8955), .A2(n8954), .ZN(n8968) );
  NAND2_X1 U5512 ( .A1(n8679), .A2(n8678), .ZN(n8990) );
  NAND2_X1 U5513 ( .A1(n4696), .A2(n9258), .ZN(n4695) );
  NOR2_X1 U5514 ( .A1(n9095), .A2(n4694), .ZN(n9056) );
  INV_X1 U5515 ( .A(n4696), .ZN(n4694) );
  NOR3_X1 U5516 ( .A1(n9160), .A2(n9119), .A3(n4689), .ZN(n9117) );
  NAND2_X1 U5517 ( .A1(n9117), .A2(n9100), .ZN(n9095) );
  NOR2_X1 U5518 ( .A1(n7514), .A2(n8608), .ZN(n7530) );
  NOR2_X1 U5519 ( .A1(n9160), .A2(n4689), .ZN(n9129) );
  NOR2_X1 U5520 ( .A1(n9160), .A2(n4690), .ZN(n9128) );
  OR2_X1 U5521 ( .A1(n7375), .A2(n9142), .ZN(n9002) );
  NOR2_X1 U5522 ( .A1(n8817), .A2(n9024), .ZN(n8799) );
  NAND2_X1 U5523 ( .A1(n9198), .A2(n7348), .ZN(n9180) );
  AND2_X1 U5524 ( .A1(n9207), .A2(n9202), .ZN(n9198) );
  OR2_X1 U5525 ( .A1(n7323), .A2(n7322), .ZN(n7325) );
  INV_X1 U5526 ( .A(n4799), .ZN(n4788) );
  NAND2_X1 U5527 ( .A1(n4794), .A2(n4799), .ZN(n4789) );
  INV_X1 U5528 ( .A(n4792), .ZN(n4791) );
  AND2_X1 U5529 ( .A1(n7223), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n7311) );
  INV_X1 U5530 ( .A(n8793), .ZN(n4622) );
  NOR2_X1 U5531 ( .A1(n7263), .A2(n4686), .ZN(n9245) );
  INV_X1 U5532 ( .A(n4688), .ZN(n4686) );
  NOR2_X1 U5533 ( .A1(n7263), .A2(n7268), .ZN(n7264) );
  OR2_X1 U5534 ( .A1(n7088), .A2(n7087), .ZN(n7178) );
  OAI21_X1 U5535 ( .B1(n7094), .B2(n4624), .A(n4623), .ZN(n7257) );
  NOR2_X1 U5536 ( .A1(n9791), .A2(n7066), .ZN(n9635) );
  AND4_X1 U5537 ( .A1(n7085), .A2(n7084), .A3(n7083), .A4(n7082), .ZN(n9641)
         );
  NAND2_X1 U5538 ( .A1(n9834), .A2(n4319), .ZN(n9790) );
  AND4_X1 U5539 ( .A1(n6366), .A2(n6365), .A3(n6364), .A4(n6363), .ZN(n9803)
         );
  AND4_X1 U5540 ( .A1(n6773), .A2(n6772), .A3(n6771), .A4(n6770), .ZN(n9801)
         );
  NAND2_X1 U5541 ( .A1(n6659), .A2(n8785), .ZN(n6930) );
  AOI21_X1 U5542 ( .B1(n6658), .B2(n8784), .A(n4761), .ZN(n6659) );
  AND2_X1 U5543 ( .A1(n6657), .A2(n9892), .ZN(n4761) );
  OR2_X1 U5544 ( .A1(n8940), .A2(n9892), .ZN(n8703) );
  NOR2_X1 U5545 ( .A1(n6342), .A2(n6341), .ZN(n6361) );
  AND2_X1 U5546 ( .A1(n9834), .A2(n6567), .ZN(n6522) );
  OR2_X1 U5547 ( .A1(n6444), .A2(n6448), .ZN(n9831) );
  NOR2_X1 U5548 ( .A1(n9831), .A2(n9835), .ZN(n9834) );
  NAND2_X1 U5549 ( .A1(n6513), .A2(n6511), .ZN(n9821) );
  INV_X1 U5550 ( .A(n9821), .ZN(n9817) );
  NAND2_X1 U5551 ( .A1(n6407), .A2(n4637), .ZN(n4636) );
  INV_X1 U5552 ( .A(n6390), .ZN(n4637) );
  NAND2_X1 U5553 ( .A1(n6391), .A2(n6390), .ZN(n8893) );
  OR2_X1 U5554 ( .A1(n6388), .A2(n6302), .ZN(n6384) );
  AND2_X1 U5555 ( .A1(n6298), .A2(n6302), .ZN(n6009) );
  INV_X1 U5556 ( .A(n9042), .ZN(n9258) );
  NAND2_X1 U5557 ( .A1(n7320), .A2(n7319), .ZN(n9325) );
  AND3_X1 U5558 ( .A1(n6314), .A2(n6313), .A3(n6312), .ZN(n9876) );
  AND3_X1 U5559 ( .A1(n6072), .A2(n6071), .A3(n6070), .ZN(n9869) );
  AND2_X1 U5560 ( .A1(n6016), .A2(n5860), .ZN(n9906) );
  AND2_X1 U5561 ( .A1(n6994), .A2(n6993), .ZN(n7007) );
  XNOR2_X1 U5562 ( .A(n5171), .B(n5170), .ZN(n8768) );
  NAND2_X1 U5563 ( .A1(n4414), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5563) );
  NAND2_X1 U5564 ( .A1(n4337), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5557) );
  NAND2_X1 U5565 ( .A1(n5555), .A2(n4644), .ZN(n4643) );
  XNOR2_X1 U5566 ( .A(n5146), .B(n5145), .ZN(n7510) );
  INV_X1 U5567 ( .A(n4909), .ZN(n4617) );
  INV_X1 U5568 ( .A(n4616), .ZN(n4615) );
  OAI21_X1 U5569 ( .B1(n4619), .B2(n4331), .A(n4913), .ZN(n4616) );
  NAND2_X1 U5570 ( .A1(n6274), .A2(n5542), .ZN(n5543) );
  XNOR2_X1 U5571 ( .A(n5117), .B(n5116), .ZN(n7332) );
  NAND2_X1 U5572 ( .A1(n5115), .A2(n5114), .ZN(n5117) );
  OR2_X1 U5573 ( .A1(n5113), .A2(n5112), .ZN(n5115) );
  OAI21_X1 U5574 ( .B1(n4872), .B2(n4330), .A(n4599), .ZN(n5101) );
  NAND2_X1 U5575 ( .A1(n4602), .A2(n4875), .ZN(n5094) );
  NAND2_X1 U5576 ( .A1(n4872), .A2(n4603), .ZN(n4602) );
  XNOR2_X1 U5577 ( .A(n5064), .B(n4436), .ZN(n7069) );
  INV_X1 U5578 ( .A(n4858), .ZN(n4436) );
  XNOR2_X1 U5579 ( .A(n5058), .B(n5057), .ZN(n6829) );
  AND2_X1 U5580 ( .A1(n5607), .A2(n5606), .ZN(n6580) );
  NAND2_X1 U5581 ( .A1(n4715), .A2(n4839), .ZN(n5042) );
  XNOR2_X1 U5582 ( .A(n4833), .B(n9533), .ZN(n5022) );
  INV_X1 U5583 ( .A(n5577), .ZN(n4758) );
  XNOR2_X1 U5584 ( .A(n4830), .B(n9464), .ZN(n5013) );
  OR2_X1 U5585 ( .A1(n4828), .A2(n4448), .ZN(n5012) );
  NAND2_X1 U5586 ( .A1(n4827), .A2(n4826), .ZN(n5002) );
  NAND2_X1 U5587 ( .A1(n4999), .A2(n4998), .ZN(n4827) );
  XNOR2_X1 U5588 ( .A(n4824), .B(SI_1_), .ZN(n4999) );
  AOI21_X1 U5589 ( .B1(n4550), .B2(n4553), .A(n7920), .ZN(n4548) );
  NAND2_X1 U5590 ( .A1(n4562), .A2(n4561), .ZN(n7053) );
  XNOR2_X1 U5591 ( .A(n7911), .B(n4805), .ZN(n8000) );
  NAND2_X1 U5592 ( .A1(n7402), .A2(n5095), .ZN(n5168) );
  OAI21_X1 U5593 ( .B1(n6546), .B2(n6490), .A(n6489), .ZN(n6639) );
  NAND2_X1 U5594 ( .A1(n4543), .A2(n4546), .ZN(n6210) );
  INV_X1 U5595 ( .A(n4544), .ZN(n4543) );
  AND2_X1 U5596 ( .A1(n4546), .A2(n4545), .ZN(n6212) );
  NAND2_X1 U5597 ( .A1(n5075), .A2(n5074), .ZN(n6927) );
  INV_X1 U5598 ( .A(n7917), .ZN(n7973) );
  NAND2_X1 U5599 ( .A1(n5152), .A2(n5151), .ZN(n8439) );
  NAND2_X1 U5600 ( .A1(n6245), .A2(n6244), .ZN(n6546) );
  NAND2_X1 U5601 ( .A1(n4542), .A2(n6192), .ZN(n6201) );
  AND2_X1 U5602 ( .A1(n5287), .A2(n5286), .ZN(n6648) );
  AND3_X1 U5603 ( .A1(n5285), .A2(n5284), .A3(n5283), .ZN(n5287) );
  NAND2_X1 U5604 ( .A1(n7952), .A2(n7893), .ZN(n8012) );
  AND2_X1 U5605 ( .A1(n4565), .A2(n4564), .ZN(n7050) );
  NAND2_X1 U5606 ( .A1(n6907), .A2(n4812), .ZN(n4564) );
  AOI21_X1 U5607 ( .B1(n7868), .B2(n4346), .A(n4568), .ZN(n8028) );
  OR2_X1 U5608 ( .A1(n4809), .A2(n4374), .ZN(n4568) );
  INV_X1 U5609 ( .A(n8045), .ZN(n8033) );
  AND2_X1 U5610 ( .A1(n5038), .A2(n4445), .ZN(n9988) );
  AND2_X1 U5611 ( .A1(n5037), .A2(n4341), .ZN(n4445) );
  NAND2_X1 U5612 ( .A1(n4549), .A2(n4554), .ZN(n8041) );
  NAND2_X1 U5613 ( .A1(n7917), .A2(n4556), .ZN(n4549) );
  OAI21_X1 U5614 ( .B1(n7917), .B2(n4553), .A(n4550), .ZN(n8039) );
  INV_X1 U5615 ( .A(n8036), .ZN(n8038) );
  NAND2_X1 U5616 ( .A1(n7106), .A2(n7105), .ZN(n7868) );
  AND2_X1 U5617 ( .A1(n7636), .A2(n7856), .ZN(n4719) );
  AND2_X1 U5618 ( .A1(n4523), .A2(n7817), .ZN(n4519) );
  NAND2_X1 U5619 ( .A1(n4336), .A2(n7856), .ZN(n4716) );
  NAND2_X1 U5620 ( .A1(n4520), .A2(n4523), .ZN(n7855) );
  INV_X1 U5621 ( .A(n8181), .ZN(n8053) );
  INV_X1 U5622 ( .A(n6648), .ZN(n8062) );
  NAND4_X1 U5623 ( .A1(n5279), .A2(n5278), .A3(n5277), .A4(n5276), .ZN(n8063)
         );
  NAND2_X1 U5624 ( .A1(n5271), .A2(n4814), .ZN(n8064) );
  AND3_X1 U5625 ( .A1(n5270), .A2(n5269), .A3(n5268), .ZN(n4814) );
  NAND2_X1 U5626 ( .A1(n9608), .A2(n5690), .ZN(n9622) );
  NAND2_X1 U5627 ( .A1(n9620), .A2(n4398), .ZN(n5696) );
  NAND2_X1 U5628 ( .A1(n9618), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n4398) );
  NAND2_X1 U5629 ( .A1(n5696), .A2(n5695), .ZN(n5710) );
  NAND2_X1 U5630 ( .A1(n4404), .A2(n5765), .ZN(n8071) );
  NAND2_X1 U5631 ( .A1(n5764), .A2(n5763), .ZN(n4404) );
  NAND2_X1 U5632 ( .A1(n8071), .A2(n8070), .ZN(n8069) );
  NAND2_X1 U5633 ( .A1(n8097), .A2(n4390), .ZN(n5771) );
  NOR2_X1 U5634 ( .A1(n5771), .A2(n5770), .ZN(n5801) );
  NOR2_X1 U5635 ( .A1(n6282), .A2(n6283), .ZN(n6285) );
  NOR2_X1 U5636 ( .A1(n6285), .A2(n6284), .ZN(n6713) );
  AND2_X1 U5637 ( .A1(n5090), .A2(n5096), .ZN(n6718) );
  NAND2_X1 U5638 ( .A1(n8105), .A2(n8106), .ZN(n8110) );
  INV_X1 U5639 ( .A(n9933), .ZN(n9929) );
  NAND2_X1 U5640 ( .A1(n4408), .A2(n4407), .ZN(n8123) );
  OAI21_X1 U5641 ( .B1(n8141), .B2(n9933), .A(n4402), .ZN(n4401) );
  AOI21_X1 U5642 ( .B1(n8142), .B2(n9930), .A(n9619), .ZN(n4402) );
  AND2_X1 U5643 ( .A1(n5177), .A2(n5176), .ZN(n8415) );
  OAI21_X1 U5644 ( .B1(n8212), .B2(n4729), .A(n4727), .ZN(n8153) );
  NAND2_X1 U5645 ( .A1(n4730), .A2(n5445), .ZN(n8171) );
  NAND2_X1 U5646 ( .A1(n8259), .A2(n5415), .ZN(n8239) );
  NAND2_X1 U5647 ( .A1(n4443), .A2(n7762), .ZN(n8274) );
  AND2_X1 U5648 ( .A1(n5131), .A2(n5130), .ZN(n8302) );
  OAI21_X1 U5649 ( .B1(n8351), .B2(n4739), .A(n4736), .ZN(n8322) );
  NAND2_X1 U5650 ( .A1(n5127), .A2(n5126), .ZN(n8471) );
  AND2_X1 U5651 ( .A1(n8348), .A2(n7734), .ZN(n8340) );
  NAND2_X1 U5652 ( .A1(n8351), .A2(n5365), .ZN(n8333) );
  NAND2_X1 U5653 ( .A1(n5111), .A2(n5110), .ZN(n8480) );
  NAND2_X1 U5654 ( .A1(n8396), .A2(n5349), .ZN(n8369) );
  NAND2_X1 U5655 ( .A1(n5501), .A2(n5500), .ZN(n7017) );
  NAND2_X1 U5656 ( .A1(n6728), .A2(n5309), .ZN(n6949) );
  INV_X1 U5657 ( .A(n9988), .ZN(n6472) );
  NAND2_X1 U5658 ( .A1(n6129), .A2(n5255), .ZN(n6687) );
  OR2_X1 U5659 ( .A1(n9956), .A2(n5828), .ZN(n8356) );
  INV_X1 U5660 ( .A(n8406), .ZN(n8359) );
  INV_X1 U5661 ( .A(n8167), .ZN(n8402) );
  AND2_X1 U5662 ( .A1(n5180), .A2(n5179), .ZN(n9632) );
  NAND2_X1 U5663 ( .A1(n8418), .A2(n4446), .ZN(n8513) );
  NAND2_X1 U5664 ( .A1(n8417), .A2(n8499), .ZN(n4457) );
  INV_X1 U5665 ( .A(n4455), .ZN(n4454) );
  OR2_X1 U5666 ( .A1(n8453), .A2(n8452), .ZN(n8519) );
  INV_X1 U5667 ( .A(n9946), .ZN(n8325) );
  AND2_X1 U5668 ( .A1(P2_U3152), .A2(n4595), .ZN(n6279) );
  NAND2_X1 U5669 ( .A1(n7575), .A2(n8767), .ZN(n7578) );
  AOI21_X1 U5670 ( .B1(n4669), .B2(n4671), .A(n4364), .ZN(n4668) );
  INV_X1 U5671 ( .A(n4671), .ZN(n4670) );
  AND3_X1 U5672 ( .A1(n7299), .A2(n7298), .A3(n7297), .ZN(n9006) );
  NAND2_X1 U5673 ( .A1(n6101), .A2(n6043), .ZN(n7283) );
  NAND2_X1 U5674 ( .A1(n8642), .A2(n4666), .ZN(n4661) );
  NAND2_X1 U5675 ( .A1(n8582), .A2(n8586), .ZN(n8595) );
  NAND2_X1 U5676 ( .A1(n4680), .A2(n6761), .ZN(n6764) );
  NAND2_X1 U5677 ( .A1(n7353), .A2(n7352), .ZN(n9306) );
  NAND2_X1 U5678 ( .A1(n7167), .A2(n7166), .ZN(n7243) );
  CLKBUF_X1 U5679 ( .A(n7199), .Z(n7200) );
  AND2_X1 U5680 ( .A1(n6095), .A2(n5884), .ZN(n8612) );
  NAND4_X1 U5681 ( .A1(n6325), .A2(n6324), .A3(n6323), .A4(n6322), .ZN(n9827)
         );
  NAND4_X1 U5682 ( .A1(n6065), .A2(n6064), .A3(n6063), .A4(n6062), .ZN(n9826)
         );
  AND2_X1 U5683 ( .A1(n6167), .A2(n5956), .ZN(n9699) );
  INV_X1 U5684 ( .A(n4473), .ZN(n9731) );
  NAND2_X1 U5685 ( .A1(n5959), .A2(n5958), .ZN(n5983) );
  AND2_X1 U5686 ( .A1(n4473), .A2(n4472), .ZN(n5959) );
  NAND2_X1 U5687 ( .A1(n5973), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n4472) );
  INV_X1 U5688 ( .A(n4479), .ZN(n9775) );
  NAND2_X1 U5689 ( .A1(n5988), .A2(n5987), .ZN(n6152) );
  AND2_X1 U5690 ( .A1(n4479), .A2(n4478), .ZN(n5988) );
  NAND2_X1 U5691 ( .A1(n6830), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4478) );
  INV_X1 U5692 ( .A(n4481), .ZN(n6537) );
  NAND2_X1 U5693 ( .A1(n4481), .A2(n4394), .ZN(n6155) );
  NOR2_X1 U5694 ( .A1(n7144), .A2(n7145), .ZN(n7148) );
  INV_X1 U5695 ( .A(n4477), .ZN(n8951) );
  INV_X1 U5696 ( .A(n8992), .ZN(n9626) );
  INV_X1 U5697 ( .A(n8990), .ZN(n9652) );
  NAND2_X1 U5698 ( .A1(n4629), .A2(n9823), .ZN(n4628) );
  AND2_X1 U5699 ( .A1(n9049), .A2(n9048), .ZN(n9264) );
  NAND2_X1 U5700 ( .A1(n4757), .A2(n9020), .ZN(n9047) );
  AND2_X1 U5701 ( .A1(n9077), .A2(n9076), .ZN(n9274) );
  NAND2_X1 U5702 ( .A1(n7547), .A2(n8767), .ZN(n7550) );
  XNOR2_X1 U5703 ( .A(n4413), .B(n9083), .ZN(n9084) );
  OAI21_X1 U5704 ( .B1(n9111), .B2(n4651), .A(n9082), .ZN(n4413) );
  NAND2_X1 U5705 ( .A1(n4773), .A2(n4778), .ZN(n9081) );
  NAND2_X1 U5706 ( .A1(n9015), .A2(n4780), .ZN(n4773) );
  NOR2_X1 U5707 ( .A1(n9111), .A2(n9029), .ZN(n9102) );
  NAND2_X1 U5708 ( .A1(n9015), .A2(n9014), .ZN(n9094) );
  AND2_X1 U5709 ( .A1(n7294), .A2(n7293), .ZN(n9007) );
  NAND2_X1 U5710 ( .A1(n7365), .A2(n7364), .ZN(n9302) );
  INV_X1 U5711 ( .A(n4767), .ZN(n9159) );
  AOI21_X1 U5712 ( .B1(n9173), .B2(n7349), .A(n4386), .ZN(n4767) );
  NAND2_X1 U5713 ( .A1(n7340), .A2(n7339), .ZN(n9313) );
  AND2_X1 U5714 ( .A1(n4639), .A2(n4327), .ZN(n9215) );
  NAND2_X1 U5715 ( .A1(n9239), .A2(n8861), .ZN(n9231) );
  NAND2_X1 U5716 ( .A1(n4790), .A2(n4794), .ZN(n9221) );
  NAND2_X1 U5717 ( .A1(n7302), .A2(n4797), .ZN(n4790) );
  OAI21_X1 U5718 ( .B1(n7302), .B2(n7301), .A(n4800), .ZN(n9238) );
  NAND2_X1 U5719 ( .A1(n9640), .A2(n8698), .ZN(n7231) );
  AND2_X1 U5720 ( .A1(n4786), .A2(n4787), .ZN(n7086) );
  NAND2_X1 U5721 ( .A1(n9634), .A2(n9672), .ZN(n4787) );
  NAND2_X1 U5722 ( .A1(n4782), .A2(n7098), .ZN(n4786) );
  INV_X1 U5723 ( .A(n9876), .ZN(n9835) );
  OR2_X1 U5724 ( .A1(n9908), .A2(n6006), .ZN(n9809) );
  INV_X1 U5725 ( .A(n6014), .ZN(n6388) );
  INV_X1 U5726 ( .A(n9063), .ZN(n9794) );
  NOR2_X1 U5727 ( .A1(n4802), .A2(n5561), .ZN(n4804) );
  AND2_X1 U5728 ( .A1(n5625), .A2(n5627), .ZN(n4803) );
  XNOR2_X1 U5729 ( .A(n4952), .B(n4951), .ZN(n9363) );
  OAI21_X1 U5730 ( .B1(n5175), .B2(n5174), .A(n4948), .ZN(n4952) );
  NAND2_X1 U5731 ( .A1(n5533), .A2(n5625), .ZN(n4801) );
  NAND2_X1 U5732 ( .A1(n4415), .A2(n5641), .ZN(n4483) );
  XNOR2_X1 U5733 ( .A(n5536), .B(n5559), .ZN(n7010) );
  XNOR2_X1 U5734 ( .A(n5142), .B(n5141), .ZN(n7492) );
  OAI21_X1 U5735 ( .B1(n4907), .B2(n4331), .A(n4615), .ZN(n5142) );
  NOR2_X1 U5736 ( .A1(n4594), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7272) );
  INV_X1 U5737 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6027) );
  NOR2_X1 U5738 ( .A1(P1_ADDR_REG_19__SCAN_IN), .A2(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n9593) );
  NAND2_X1 U5739 ( .A1(n4403), .A2(n4399), .ZN(P2_U3264) );
  AOI21_X1 U5740 ( .B1(n4401), .B2(n9946), .A(n4400), .ZN(n4399) );
  OR2_X1 U5741 ( .A1(n8143), .A2(n9946), .ZN(n4403) );
  OAI21_X1 U5742 ( .B1(n9604), .B2(n8146), .A(n8145), .ZN(n4400) );
  NAND2_X1 U5743 ( .A1(n4453), .A2(n4452), .ZN(P2_U3517) );
  NAND2_X1 U5744 ( .A1(n10017), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n4452) );
  NAND2_X1 U5745 ( .A1(n8513), .A2(n10019), .ZN(n4453) );
  AOI21_X1 U5746 ( .B1(n4320), .B2(n4419), .A(n4418), .ZN(P1_U3240) );
  NOR2_X1 U5747 ( .A1(n4357), .A2(n4420), .ZN(n4418) );
  NOR3_X1 U5748 ( .A1(n4421), .A2(n4422), .A3(n4420), .ZN(n4419) );
  INV_X1 U5749 ( .A(n6996), .ZN(n5844) );
  XNOR2_X1 U5750 ( .A(n5547), .B(n5546), .ZN(n5859) );
  AND2_X1 U5751 ( .A1(n4310), .A2(n4575), .ZN(n4971) );
  INV_X1 U5752 ( .A(n5972), .ZN(n4475) );
  AND2_X1 U5753 ( .A1(n8874), .A2(n8915), .ZN(n9035) );
  NAND2_X1 U5754 ( .A1(n8862), .A2(n8822), .ZN(n9220) );
  XNOR2_X1 U5755 ( .A(n5201), .B(n5200), .ZN(n5218) );
  NAND2_X1 U5756 ( .A1(n5505), .A2(n8211), .ZN(n8193) );
  NAND2_X1 U5757 ( .A1(n4758), .A2(n5523), .ZN(n5579) );
  OR2_X1 U5758 ( .A1(n8427), .A2(n8052), .ZN(n4317) );
  AND2_X1 U5759 ( .A1(n9892), .A2(n6567), .ZN(n4318) );
  INV_X1 U5760 ( .A(n7795), .ZN(n4506) );
  INV_X1 U5761 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5625) );
  AND2_X1 U5762 ( .A1(n4318), .A2(n6931), .ZN(n4319) );
  INV_X1 U5763 ( .A(n6407), .ZN(n4638) );
  AND2_X1 U5764 ( .A1(n8885), .A2(n6996), .ZN(n4320) );
  AND2_X1 U5765 ( .A1(n4506), .A2(n5463), .ZN(n8155) );
  INV_X1 U5766 ( .A(n8155), .ZN(n4726) );
  AND2_X1 U5767 ( .A1(n7847), .A2(n7811), .ZN(n4321) );
  NOR2_X1 U5768 ( .A1(n4808), .A2(n4383), .ZN(n4322) );
  AND2_X1 U5769 ( .A1(n4729), .A2(n4726), .ZN(n4323) );
  AND2_X1 U5770 ( .A1(n4739), .A2(n4338), .ZN(n4324) );
  NAND2_X1 U5771 ( .A1(n4635), .A2(n9051), .ZN(n4325) );
  NOR2_X1 U5772 ( .A1(n7773), .A2(n7811), .ZN(n4326) );
  NAND2_X1 U5773 ( .A1(n7578), .A2(n7577), .ZN(n9271) );
  INV_X1 U5774 ( .A(n9271), .ZN(n4699) );
  INV_X1 U5775 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5944) );
  AND2_X1 U5776 ( .A1(n4640), .A2(n8822), .ZN(n4327) );
  NOR2_X1 U5777 ( .A1(n6453), .A2(n7678), .ZN(n4328) );
  INV_X1 U5778 ( .A(n7916), .ZN(n4557) );
  NAND2_X1 U5779 ( .A1(n7201), .A2(n4673), .ZN(n7167) );
  INV_X1 U5780 ( .A(n9243), .ZN(n4439) );
  INV_X1 U5781 ( .A(n7635), .ZN(n7902) );
  INV_X2 U5782 ( .A(n5035), .ZN(n5095) );
  INV_X2 U5783 ( .A(n6350), .ZN(n8767) );
  OAI211_X1 U5784 ( .C1(n5036), .C2(n5582), .A(n4451), .B(n4450), .ZN(n5233)
         );
  NAND2_X1 U5785 ( .A1(n6400), .A2(n7288), .ZN(n6429) );
  OR2_X1 U5786 ( .A1(n9095), .A2(n4695), .ZN(n4329) );
  NOR2_X1 U5787 ( .A1(n4984), .A2(P2_IR_REG_29__SCAN_IN), .ZN(n4988) );
  OR2_X1 U5788 ( .A1(n5093), .A2(n4601), .ZN(n4330) );
  OR2_X1 U5789 ( .A1(n5137), .A2(n4617), .ZN(n4331) );
  OR2_X1 U5790 ( .A1(n8260), .A2(n8261), .ZN(n8259) );
  OR2_X1 U5791 ( .A1(n5562), .A2(P1_IR_REG_23__SCAN_IN), .ZN(n4332) );
  AND2_X1 U5792 ( .A1(n9369), .A2(n9374), .ZN(n4333) );
  NAND2_X1 U5793 ( .A1(n5012), .A2(n4831), .ZN(n4334) );
  INV_X1 U5794 ( .A(n7623), .ZN(n5808) );
  NAND2_X1 U5795 ( .A1(n7465), .A2(n7464), .ZN(n4335) );
  NOR2_X1 U5796 ( .A1(n5577), .A2(n4759), .ZN(n5586) );
  OR2_X1 U5797 ( .A1(n5308), .A2(n6801), .ZN(n7705) );
  NAND2_X1 U5798 ( .A1(n5030), .A2(n4747), .ZN(n5045) );
  AND2_X1 U5799 ( .A1(n7855), .A2(n7854), .ZN(n4336) );
  OR2_X1 U5800 ( .A1(n5562), .A2(n4643), .ZN(n4337) );
  XNOR2_X1 U5801 ( .A(n6007), .B(n6014), .ZN(n6008) );
  OR2_X1 U5802 ( .A1(n8471), .A2(n8341), .ZN(n4338) );
  NAND4_X1 U5803 ( .A1(n5241), .A2(n5240), .A3(n5239), .A4(n5238), .ZN(n5818)
         );
  NAND2_X1 U5804 ( .A1(n8310), .A2(n7751), .ZN(n8282) );
  OR2_X1 U5805 ( .A1(n8694), .A2(n8773), .ZN(n4339) );
  OR2_X1 U5806 ( .A1(n8874), .A2(n8773), .ZN(n4340) );
  OR2_X1 U5807 ( .A1(n5682), .A2(n5748), .ZN(n4341) );
  OR2_X1 U5808 ( .A1(n8419), .A2(n8365), .ZN(n4342) );
  AND4_X1 U5809 ( .A1(n4964), .A2(n4963), .A3(n4962), .A4(n4961), .ZN(n4343)
         );
  OR2_X1 U5810 ( .A1(n6108), .A2(n5543), .ZN(n4344) );
  NAND2_X1 U5811 ( .A1(n8277), .A2(n4722), .ZN(n8244) );
  OR2_X1 U5812 ( .A1(n7066), .A2(n9801), .ZN(n8850) );
  AND2_X1 U5813 ( .A1(n7833), .A2(n7723), .ZN(n4345) );
  INV_X1 U5814 ( .A(n8879), .ZN(n4591) );
  NAND2_X1 U5815 ( .A1(n4740), .A2(n5003), .ZN(n5017) );
  AND2_X1 U5816 ( .A1(n7883), .A2(n4571), .ZN(n4346) );
  AND2_X1 U5817 ( .A1(n7212), .A2(n7211), .ZN(n7300) );
  INV_X1 U5818 ( .A(n7300), .ZN(n9339) );
  INV_X1 U5819 ( .A(n5918), .ZN(n4595) );
  NAND2_X1 U5820 ( .A1(n7405), .A2(n7404), .ZN(n9061) );
  AND2_X1 U5821 ( .A1(n5956), .A2(n9700), .ZN(n4347) );
  NAND2_X1 U5822 ( .A1(n4510), .A2(n5055), .ZN(n6975) );
  NAND4_X1 U5823 ( .A1(n5263), .A2(n5262), .A3(n5261), .A4(n5260), .ZN(n8065)
         );
  INV_X1 U5824 ( .A(n9907), .ZN(n6941) );
  AND2_X1 U5825 ( .A1(n6750), .A2(n6749), .ZN(n9907) );
  NAND2_X1 U5826 ( .A1(n5160), .A2(n5159), .ZN(n8433) );
  OR2_X1 U5827 ( .A1(n6030), .A2(n5963), .ZN(n4348) );
  INV_X1 U5828 ( .A(n5041), .ZN(n4840) );
  XNOR2_X1 U5829 ( .A(n4841), .B(SI_7_), .ZN(n5041) );
  INV_X1 U5830 ( .A(n7815), .ZN(n4524) );
  AND2_X1 U5831 ( .A1(n8172), .A2(n7785), .ZN(n4349) );
  NAND2_X1 U5832 ( .A1(n7780), .A2(n7781), .ZN(n8213) );
  NOR2_X1 U5833 ( .A1(n8422), .A2(n8182), .ZN(n7795) );
  AND2_X1 U5834 ( .A1(n7732), .A2(n7729), .ZN(n4350) );
  OR2_X1 U5835 ( .A1(n8065), .A2(n5264), .ZN(n4351) );
  AND2_X1 U5836 ( .A1(n4642), .A2(n8861), .ZN(n4352) );
  INV_X1 U5837 ( .A(n7724), .ZN(n4710) );
  AND2_X1 U5838 ( .A1(n8471), .A2(n8341), .ZN(n4353) );
  AND2_X1 U5839 ( .A1(n8240), .A2(n7775), .ZN(n4354) );
  NOR2_X1 U5840 ( .A1(n9253), .A2(n9235), .ZN(n4355) );
  AND2_X1 U5841 ( .A1(n8422), .A2(n8182), .ZN(n7794) );
  AND2_X1 U5842 ( .A1(n8339), .A2(n7734), .ZN(n4356) );
  AND2_X1 U5843 ( .A1(n5051), .A2(n5050), .ZN(n9995) );
  INV_X1 U5844 ( .A(n9995), .ZN(n6814) );
  INV_X1 U5845 ( .A(n4607), .ZN(n4606) );
  NOR2_X1 U5846 ( .A1(n5069), .A2(n4608), .ZN(n4607) );
  INV_X1 U5847 ( .A(n4570), .ZN(n4569) );
  NOR2_X1 U5848 ( .A1(n7869), .A2(n7867), .ZN(n4570) );
  AND2_X1 U5849 ( .A1(n8924), .A2(n4424), .ZN(n4357) );
  AND2_X1 U5850 ( .A1(n4520), .A2(n4519), .ZN(n4358) );
  INV_X1 U5851 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5542) );
  NAND2_X1 U5852 ( .A1(n5568), .A2(n4654), .ZN(n5577) );
  INV_X1 U5853 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n4959) );
  OR2_X1 U5854 ( .A1(n7727), .A2(n8397), .ZN(n4359) );
  INV_X1 U5855 ( .A(n7759), .ZN(n7751) );
  AND2_X1 U5856 ( .A1(n8302), .A2(n8319), .ZN(n7759) );
  AND2_X1 U5857 ( .A1(n4841), .A2(SI_7_), .ZN(n4360) );
  NOR2_X1 U5858 ( .A1(n8422), .A2(n8051), .ZN(n4361) );
  AND2_X1 U5859 ( .A1(n8889), .A2(n4636), .ZN(n4362) );
  NAND2_X1 U5860 ( .A1(n4971), .A2(n4972), .ZN(n4363) );
  INV_X1 U5861 ( .A(n4794), .ZN(n4793) );
  NOR2_X1 U5862 ( .A1(n4355), .A2(n4795), .ZN(n4794) );
  AND2_X1 U5863 ( .A1(n7241), .A2(n7240), .ZN(n4364) );
  NAND2_X1 U5864 ( .A1(n7786), .A2(n8172), .ZN(n4365) );
  AND2_X1 U5865 ( .A1(n6334), .A2(n6418), .ZN(n4366) );
  INV_X1 U5866 ( .A(n5561), .ZN(n4415) );
  INV_X1 U5867 ( .A(n4707), .ZN(n4706) );
  NOR2_X1 U5868 ( .A1(n7624), .A2(n7795), .ZN(n4707) );
  AND2_X1 U5869 ( .A1(n4971), .A2(n4586), .ZN(n4367) );
  INV_X1 U5870 ( .A(n7745), .ZN(n8375) );
  INV_X1 U5871 ( .A(n8228), .ZN(n8240) );
  NAND2_X1 U5872 ( .A1(n8214), .A2(n7777), .ZN(n8228) );
  INV_X1 U5873 ( .A(n7796), .ZN(n7802) );
  AND2_X1 U5874 ( .A1(n8416), .A2(n8158), .ZN(n7796) );
  OR2_X1 U5875 ( .A1(n5562), .A2(n4645), .ZN(n4368) );
  INV_X1 U5876 ( .A(n8172), .ZN(n8179) );
  AND2_X1 U5877 ( .A1(n7791), .A2(n7788), .ZN(n8172) );
  AND2_X1 U5878 ( .A1(n7776), .A2(n7811), .ZN(n4369) );
  INV_X1 U5879 ( .A(n9035), .ZN(n4635) );
  NAND2_X1 U5880 ( .A1(n8697), .A2(n4625), .ZN(n4370) );
  INV_X1 U5881 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n6274) );
  NAND2_X1 U5882 ( .A1(n4764), .A2(n4768), .ZN(n9005) );
  NAND2_X1 U5883 ( .A1(n8560), .A2(n8559), .ZN(n4371) );
  AND2_X1 U5884 ( .A1(n8244), .A2(n7775), .ZN(n8227) );
  NOR2_X1 U5885 ( .A1(n8134), .A2(n8133), .ZN(n4372) );
  NAND2_X1 U5886 ( .A1(n7495), .A2(n7494), .ZN(n9291) );
  NOR2_X1 U5887 ( .A1(n7048), .A2(n7047), .ZN(n4373) );
  AND2_X1 U5888 ( .A1(n7883), .A2(n4570), .ZN(n4374) );
  AND2_X1 U5889 ( .A1(n8211), .A2(n7779), .ZN(n4375) );
  AND2_X1 U5890 ( .A1(n4327), .A2(n8823), .ZN(n4376) );
  AND2_X1 U5891 ( .A1(n4752), .A2(n4967), .ZN(n4377) );
  AND2_X1 U5892 ( .A1(n8228), .A2(n5415), .ZN(n4378) );
  AND2_X1 U5893 ( .A1(n9021), .A2(n9020), .ZN(n4379) );
  AND2_X1 U5894 ( .A1(n7745), .A2(n5349), .ZN(n4380) );
  AND2_X1 U5895 ( .A1(n7569), .A2(n7545), .ZN(n4381) );
  AND2_X1 U5896 ( .A1(n8881), .A2(n9840), .ZN(n4382) );
  INV_X1 U5897 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5627) );
  AND2_X1 U5898 ( .A1(n7901), .A2(n7900), .ZN(n4383) );
  AND2_X1 U5899 ( .A1(n4319), .A2(n9907), .ZN(n4384) );
  AND2_X1 U5900 ( .A1(n5031), .A2(n4954), .ZN(n4747) );
  OR2_X1 U5901 ( .A1(n8011), .A2(n7898), .ZN(n4385) );
  INV_X1 U5902 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n4646) );
  NAND2_X1 U5903 ( .A1(n9239), .A2(n4352), .ZN(n4639) );
  NAND2_X1 U5904 ( .A1(n7072), .A2(n7071), .ZN(n8692) );
  INV_X1 U5905 ( .A(n8692), .ZN(n9672) );
  NOR2_X1 U5906 ( .A1(n7348), .A2(n7347), .ZN(n4386) );
  INV_X1 U5907 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n4509) );
  OR2_X1 U5908 ( .A1(n5748), .A2(n6462), .ZN(n4387) );
  OAI21_X1 U5909 ( .B1(n8389), .B2(n7741), .A(n7728), .ZN(n8374) );
  NAND2_X1 U5910 ( .A1(n4734), .A2(n4733), .ZN(n8297) );
  NAND2_X1 U5911 ( .A1(n7026), .A2(n7723), .ZN(n7014) );
  NAND2_X1 U5912 ( .A1(n7019), .A2(n7725), .ZN(n8389) );
  NAND2_X1 U5913 ( .A1(n4661), .A2(n4665), .ZN(n8558) );
  INV_X1 U5914 ( .A(n9229), .ZN(n4641) );
  INV_X1 U5915 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n4960) );
  AND2_X1 U5916 ( .A1(n5586), .A2(n5527), .ZN(n5639) );
  AND4_X1 U5917 ( .A1(n7604), .A2(n7603), .A3(n7602), .A4(n7601), .ZN(n8777)
         );
  NAND2_X1 U5918 ( .A1(n4720), .A2(n4350), .ZN(n8348) );
  NAND2_X1 U5919 ( .A1(n4567), .A2(n4569), .ZN(n7978) );
  NAND2_X1 U5920 ( .A1(n4720), .A2(n7729), .ZN(n8346) );
  NAND2_X1 U5921 ( .A1(n5504), .A2(n7750), .ZN(n8303) );
  NAND2_X1 U5922 ( .A1(n5168), .A2(n5167), .ZN(n8422) );
  INV_X1 U5923 ( .A(n8422), .ZN(n4469) );
  NAND2_X1 U5924 ( .A1(n5173), .A2(n5172), .ZN(n8416) );
  INV_X1 U5925 ( .A(n8416), .ZN(n4467) );
  NOR3_X1 U5926 ( .A1(n7263), .A2(n9330), .A3(n4687), .ZN(n4684) );
  NAND2_X1 U5927 ( .A1(n7550), .A2(n7549), .ZN(n9278) );
  INV_X1 U5928 ( .A(n9278), .ZN(n4698) );
  NAND2_X1 U5929 ( .A1(n4310), .A2(n5030), .ZN(n5102) );
  AND2_X1 U5930 ( .A1(n7201), .A2(n7134), .ZN(n7135) );
  OR2_X1 U5931 ( .A1(n6931), .A2(n9803), .ZN(n4388) );
  INV_X1 U5932 ( .A(n4691), .ZN(n9152) );
  NOR2_X1 U5933 ( .A1(n9160), .A2(n9302), .ZN(n4691) );
  INV_X1 U5934 ( .A(n4685), .ZN(n9246) );
  NOR2_X1 U5935 ( .A1(n7263), .A2(n4687), .ZN(n4685) );
  OR2_X1 U5936 ( .A1(n6113), .A2(n6114), .ZN(n4389) );
  OR2_X1 U5937 ( .A1(n5779), .A2(n5768), .ZN(n4390) );
  INV_X1 U5938 ( .A(n9318), .ZN(n9202) );
  NAND2_X1 U5939 ( .A1(n7334), .A2(n7333), .ZN(n9318) );
  AND2_X1 U5940 ( .A1(n8315), .A2(n8302), .ZN(n8285) );
  AND2_X1 U5941 ( .A1(n7513), .A2(n7512), .ZN(n9013) );
  INV_X1 U5942 ( .A(n9013), .ZN(n9119) );
  AND2_X1 U5943 ( .A1(n5161), .A2(n5155), .ZN(n4391) );
  OR2_X1 U5944 ( .A1(n9672), .A2(n7098), .ZN(n4392) );
  NAND4_X1 U5945 ( .A1(n5937), .A2(n5936), .A3(n5935), .A4(n5934), .ZN(n8944)
         );
  AND2_X1 U5946 ( .A1(n7169), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4393) );
  OAI22_X1 U5947 ( .A1(n6619), .A2(n5497), .B1(n5496), .B2(n5495), .ZN(n6950)
         );
  NAND2_X1 U5948 ( .A1(n5121), .A2(n5120), .ZN(n8474) );
  INV_X1 U5949 ( .A(n8474), .ZN(n4462) );
  OR2_X1 U5950 ( .A1(n7074), .A2(n7081), .ZN(n4394) );
  AND2_X1 U5951 ( .A1(n4573), .A2(n4310), .ZN(n5107) );
  AND2_X1 U5952 ( .A1(n7444), .A2(n7445), .ZN(n8583) );
  INV_X1 U5953 ( .A(n9242), .ZN(n9823) );
  NAND4_X1 U5954 ( .A1(n5228), .A2(n5227), .A3(n5226), .A4(n5225), .ZN(n5887)
         );
  NAND3_X1 U5955 ( .A1(n4584), .A2(n4582), .A3(n4580), .ZN(n7852) );
  INV_X1 U5956 ( .A(n7852), .ZN(n6543) );
  AND2_X1 U5957 ( .A1(n5237), .A2(n5236), .ZN(n5913) );
  OR2_X1 U5958 ( .A1(n5656), .A2(n6543), .ZN(n4395) );
  AND2_X1 U5959 ( .A1(n6026), .A2(n6025), .ZN(n4396) );
  INV_X1 U5960 ( .A(SI_2_), .ZN(n4448) );
  XNOR2_X1 U5961 ( .A(n4977), .B(n4976), .ZN(n7818) );
  INV_X1 U5962 ( .A(n5223), .ZN(n7400) );
  INV_X1 U5963 ( .A(n5224), .ZN(n7937) );
  AND2_X1 U5964 ( .A1(n5938), .A2(n6257), .ZN(n4397) );
  XNOR2_X1 U5965 ( .A(n5563), .B(n5625), .ZN(n6257) );
  INV_X2 U5966 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  AOI21_X1 U5967 ( .B1(n7631), .B2(n8498), .A(n7275), .ZN(n5180) );
  NAND2_X1 U5968 ( .A1(n8416), .A2(n8498), .ZN(n4456) );
  INV_X1 U5969 ( .A(n8498), .ZN(n10008) );
  NAND2_X1 U5970 ( .A1(n5515), .A2(n8395), .ZN(n4447) );
  NOR2_X1 U5971 ( .A1(n8123), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n8134) );
  NAND2_X1 U5972 ( .A1(n8122), .A2(n8135), .ZN(n4407) );
  INV_X1 U5973 ( .A(n8133), .ZN(n4408) );
  NAND3_X1 U5974 ( .A1(n8783), .A2(n9817), .A3(n4409), .ZN(n8787) );
  NOR2_X2 U5975 ( .A1(n9820), .A2(n8836), .ZN(n6519) );
  NAND2_X1 U5976 ( .A1(n6510), .A2(n8834), .ZN(n9820) );
  NAND2_X1 U5977 ( .A1(n8837), .A2(n6428), .ZN(n4410) );
  NOR2_X2 U5978 ( .A1(n7232), .A2(n8795), .ZN(n7381) );
  NAND3_X1 U5979 ( .A1(n4621), .A2(n8855), .A3(n4411), .ZN(n7232) );
  NAND3_X1 U5980 ( .A1(n7094), .A2(n4623), .A3(n4622), .ZN(n4411) );
  NAND4_X1 U5981 ( .A1(n5529), .A2(n4412), .A3(n6274), .A4(n5661), .ZN(n5532)
         );
  NOR2_X2 U5982 ( .A1(n9112), .A2(n9113), .ZN(n9111) );
  NAND3_X1 U5983 ( .A1(n5641), .A2(n5533), .A3(n4415), .ZN(n4414) );
  AND2_X1 U5984 ( .A1(n8882), .A2(n9154), .ZN(n4425) );
  NAND2_X1 U5985 ( .A1(n8338), .A2(n7749), .ZN(n8316) );
  OAI21_X1 U5986 ( .B1(n4829), .B2(P1_DATAO_REG_2__SCAN_IN), .A(n4449), .ZN(
        n4828) );
  NAND2_X1 U5987 ( .A1(n4829), .A2(n6027), .ZN(n4449) );
  NAND2_X2 U5988 ( .A1(n5682), .A2(n4595), .ZN(n5036) );
  NAND2_X2 U5989 ( .A1(n4994), .A2(n4993), .ZN(n5682) );
  NAND2_X1 U5990 ( .A1(n4460), .A2(n4458), .ZN(n6787) );
  NAND3_X1 U5991 ( .A1(n4464), .A2(n4465), .A3(n6248), .ZN(n6692) );
  NAND2_X1 U5992 ( .A1(n6160), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n4471) );
  NAND2_X1 U5993 ( .A1(n6267), .A2(n5954), .ZN(n6168) );
  NOR2_X2 U5994 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5568) );
  XNOR2_X2 U5995 ( .A(n4482), .B(n5627), .ZN(n9374) );
  NAND3_X1 U5996 ( .A1(n4489), .A2(n4487), .A3(n4340), .ZN(n4486) );
  NAND2_X1 U5997 ( .A1(n5002), .A2(n5001), .ZN(n4504) );
  NAND2_X1 U5998 ( .A1(n4503), .A2(n4502), .ZN(n5021) );
  NAND3_X1 U5999 ( .A1(n4311), .A2(n5002), .A3(n5001), .ZN(n4503) );
  NAND2_X1 U6000 ( .A1(n4504), .A2(n5012), .ZN(n5014) );
  NAND2_X1 U6001 ( .A1(n6748), .A2(n5095), .ZN(n4510) );
  XNOR2_X1 U6002 ( .A(n5053), .B(n5052), .ZN(n6748) );
  NAND2_X1 U6003 ( .A1(n5027), .A2(n4515), .ZN(n4513) );
  NAND2_X1 U6004 ( .A1(n5027), .A2(n5026), .ZN(n4514) );
  NAND2_X1 U6005 ( .A1(n7813), .A2(n4521), .ZN(n4520) );
  NAND2_X1 U6006 ( .A1(n7774), .A2(n4527), .ZN(n4525) );
  NAND2_X1 U6007 ( .A1(n4525), .A2(n4526), .ZN(n7793) );
  NAND2_X1 U6008 ( .A1(n5815), .A2(n5816), .ZN(n4545) );
  NAND2_X1 U6009 ( .A1(n4544), .A2(n4546), .ZN(n6188) );
  NAND2_X1 U6010 ( .A1(n7917), .A2(n4550), .ZN(n4547) );
  NAND2_X1 U6011 ( .A1(n4547), .A2(n4548), .ZN(n7942) );
  NAND2_X1 U6012 ( .A1(n7952), .A2(n4558), .ZN(n4560) );
  NAND3_X1 U6013 ( .A1(n4562), .A2(n4561), .A3(n7051), .ZN(n7106) );
  AOI21_X1 U6014 ( .B1(n4811), .B2(n4566), .A(n4373), .ZN(n4561) );
  NAND2_X1 U6015 ( .A1(n6907), .A2(n4563), .ZN(n4562) );
  INV_X1 U6016 ( .A(n4811), .ZN(n4565) );
  INV_X1 U6017 ( .A(n7049), .ZN(n4566) );
  OAI22_X1 U6018 ( .A1(n4586), .A2(n4585), .B1(P2_IR_REG_31__SCAN_IN), .B2(
        n4960), .ZN(n4581) );
  NAND2_X1 U6019 ( .A1(n4971), .A2(n4583), .ZN(n4582) );
  OR2_X1 U6020 ( .A1(n4971), .A2(n4585), .ZN(n4584) );
  OAI22_X1 U6021 ( .A1(n6188), .A2(n6187), .B1(n6186), .B2(n6185), .ZN(n6219)
         );
  NOR2_X1 U6022 ( .A1(n8875), .A2(n4591), .ZN(n4590) );
  INV_X1 U6023 ( .A(n8875), .ZN(n4593) );
  MUX2_X1 U6024 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(P1_DATAO_REG_4__SCAN_IN), 
        .S(n5918), .Z(n4833) );
  MUX2_X1 U6025 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n5918), .Z(n4841) );
  MUX2_X1 U6026 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n5918), .Z(n4838) );
  MUX2_X1 U6027 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n5918), .Z(n4836) );
  MUX2_X1 U6028 ( .A(n5609), .B(n5601), .S(n5918), .Z(n4842) );
  MUX2_X1 U6029 ( .A(n4846), .B(n5613), .S(n5918), .Z(n4847) );
  MUX2_X1 U6030 ( .A(n5619), .B(n5614), .S(n5918), .Z(n4853) );
  MUX2_X1 U6031 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(P1_DATAO_REG_11__SCAN_IN), 
        .S(n4594), .Z(n4859) );
  MUX2_X1 U6032 ( .A(n5644), .B(n5646), .S(n4594), .Z(n4861) );
  MUX2_X1 U6033 ( .A(n4865), .B(n4866), .S(n4594), .Z(n4868) );
  MUX2_X1 U6034 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(P1_DATAO_REG_14__SCAN_IN), 
        .S(n4594), .Z(n4874) );
  MUX2_X1 U6035 ( .A(n5793), .B(n5795), .S(n4594), .Z(n4877) );
  MUX2_X1 U6036 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(P1_DATAO_REG_18__SCAN_IN), 
        .S(n4594), .Z(n4888) );
  MUX2_X1 U6037 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(P1_DATAO_REG_17__SCAN_IN), 
        .S(n4594), .Z(n4892) );
  MUX2_X1 U6038 ( .A(n5947), .B(n6002), .S(n4594), .Z(n4882) );
  MUX2_X1 U6039 ( .A(n6373), .B(n6375), .S(n4594), .Z(n4896) );
  MUX2_X1 U6040 ( .A(n7351), .B(n6507), .S(n4594), .Z(n4903) );
  MUX2_X1 U6041 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n4594), .Z(n4908) );
  MUX2_X1 U6042 ( .A(n7292), .B(n7865), .S(n4594), .Z(n4910) );
  MUX2_X1 U6043 ( .A(n7493), .B(n6857), .S(n4594), .Z(n4915) );
  MUX2_X1 U6044 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n4594), .Z(n4922) );
  MUX2_X1 U6045 ( .A(n7527), .B(n7063), .S(n4594), .Z(n4925) );
  MUX2_X1 U6046 ( .A(n7548), .B(n7191), .S(n4594), .Z(n4930) );
  MUX2_X1 U6047 ( .A(n7576), .B(n7208), .S(n4594), .Z(n4933) );
  MUX2_X1 U6048 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(P1_DATAO_REG_28__SCAN_IN), 
        .S(n4594), .Z(n4937) );
  MUX2_X1 U6049 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(P1_DATAO_REG_29__SCAN_IN), 
        .S(n4594), .Z(n5169) );
  MUX2_X1 U6050 ( .A(n9371), .B(n7938), .S(n4594), .Z(n4945) );
  MUX2_X1 U6051 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n4594), .Z(n4950) );
  NAND2_X1 U6052 ( .A1(n4872), .A2(n4599), .ZN(n4598) );
  NAND2_X1 U6053 ( .A1(n4872), .A2(n4871), .ZN(n5083) );
  NAND2_X1 U6054 ( .A1(n4932), .A2(n4391), .ZN(n4605) );
  NAND2_X1 U6055 ( .A1(n4857), .A2(n4856), .ZN(n5064) );
  NAND2_X1 U6056 ( .A1(n4907), .A2(n4615), .ZN(n4614) );
  NAND2_X1 U6057 ( .A1(n4907), .A2(n4619), .ZN(n4618) );
  NAND2_X1 U6058 ( .A1(n4907), .A2(n4906), .ZN(n5134) );
  NAND3_X1 U6059 ( .A1(n4622), .A2(n4623), .A3(n4624), .ZN(n4621) );
  NAND2_X1 U6060 ( .A1(n9052), .A2(n4627), .ZN(n4626) );
  OAI211_X1 U6061 ( .C1(n9052), .C2(n4628), .A(n9038), .B(n4626), .ZN(n9261)
         );
  NAND2_X1 U6062 ( .A1(n9052), .A2(n9051), .ZN(n9050) );
  NAND2_X1 U6063 ( .A1(n4639), .A2(n4376), .ZN(n9190) );
  INV_X1 U6064 ( .A(n9220), .ZN(n4642) );
  INV_X1 U6065 ( .A(n4759), .ZN(n4653) );
  AND2_X2 U6066 ( .A1(n5527), .A2(n4652), .ZN(n5641) );
  NAND3_X1 U6067 ( .A1(n6102), .A2(n6026), .A3(n6025), .ZN(n6101) );
  OAI21_X2 U6068 ( .B1(n7283), .B2(n7279), .A(n7280), .ZN(n6307) );
  INV_X1 U6069 ( .A(n4655), .ZN(n6415) );
  NAND2_X1 U6070 ( .A1(n6565), .A2(n6558), .ZN(n6576) );
  OAI21_X2 U6071 ( .B1(n4655), .B2(n4366), .A(n6337), .ZN(n6565) );
  NAND2_X1 U6072 ( .A1(n6309), .A2(n6308), .ZN(n4655) );
  INV_X1 U6073 ( .A(n8586), .ZN(n4658) );
  NAND2_X1 U6074 ( .A1(n8585), .A2(n8586), .ZN(n4659) );
  OAI21_X1 U6075 ( .B1(n6108), .B2(n4677), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5843) );
  INV_X1 U6076 ( .A(n4674), .ZN(n5545) );
  NAND2_X1 U6077 ( .A1(n7546), .A2(n7545), .ZN(n8649) );
  NAND2_X1 U6078 ( .A1(n7546), .A2(n4381), .ZN(n8651) );
  NAND3_X1 U6079 ( .A1(n5586), .A2(n5527), .A3(n4681), .ZN(n5660) );
  INV_X1 U6080 ( .A(n4684), .ZN(n9222) );
  NAND2_X1 U6081 ( .A1(n4384), .A2(n9834), .ZN(n9791) );
  NAND2_X2 U6082 ( .A1(n6030), .A2(n5918), .ZN(n6067) );
  OAI21_X1 U6083 ( .B1(n8156), .B2(n4706), .A(n4705), .ZN(n7626) );
  INV_X1 U6084 ( .A(n4700), .ZN(n7627) );
  INV_X1 U6085 ( .A(n4703), .ZN(n4701) );
  INV_X1 U6086 ( .A(n7810), .ZN(n4704) );
  NAND2_X1 U6087 ( .A1(n5501), .A2(n4708), .ZN(n7019) );
  NAND2_X1 U6088 ( .A1(n7725), .A2(n7724), .ZN(n7833) );
  NAND2_X1 U6089 ( .A1(n5034), .A2(n5033), .ZN(n4715) );
  NAND2_X1 U6090 ( .A1(n4358), .A2(n7856), .ZN(n4717) );
  NAND2_X1 U6091 ( .A1(n7637), .A2(n4719), .ZN(n4718) );
  NAND4_X1 U6092 ( .A1(n4718), .A2(n7863), .A3(n4717), .A4(n4716), .ZN(
        P2_U3244) );
  NAND2_X1 U6093 ( .A1(n8212), .A2(n4725), .ZN(n4724) );
  NAND2_X1 U6094 ( .A1(n8212), .A2(n5442), .ZN(n4730) );
  NAND2_X1 U6095 ( .A1(n8351), .A2(n4735), .ZN(n4734) );
  NAND3_X1 U6096 ( .A1(n5003), .A2(n4740), .A3(n4953), .ZN(n5019) );
  NAND2_X1 U6097 ( .A1(n6226), .A2(n4744), .ZN(n4743) );
  OAI211_X1 U6098 ( .C1(n6130), .C2(n4746), .A(n4743), .B(n4741), .ZN(n6452)
         );
  NAND2_X1 U6099 ( .A1(n8396), .A2(n4380), .ZN(n8371) );
  NAND2_X1 U6100 ( .A1(n8259), .A2(n4378), .ZN(n8237) );
  NAND2_X1 U6101 ( .A1(n5107), .A2(n4377), .ZN(n4979) );
  INV_X1 U6102 ( .A(n4979), .ZN(n4980) );
  NAND2_X1 U6103 ( .A1(n9369), .A2(n4753), .ZN(n4754) );
  AND2_X1 U6104 ( .A1(n9374), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n4753) );
  NAND2_X2 U6105 ( .A1(n5631), .A2(n9374), .ZN(n7598) );
  NAND3_X1 U6106 ( .A1(n5631), .A2(n9374), .A3(P1_REG2_REG_1__SCAN_IN), .ZN(
        n4755) );
  NAND2_X1 U6107 ( .A1(n4757), .A2(n4379), .ZN(n9049) );
  NAND2_X1 U6108 ( .A1(n9316), .A2(n4765), .ZN(n4764) );
  NAND2_X1 U6109 ( .A1(n9015), .A2(n4774), .ZN(n4770) );
  NAND2_X1 U6110 ( .A1(n4770), .A2(n4771), .ZN(n9067) );
  NAND2_X1 U6111 ( .A1(n9634), .A2(n4392), .ZN(n4785) );
  OAI22_X1 U6112 ( .A1(n7302), .A2(n4789), .B1(n4788), .B2(n4791), .ZN(n9206)
         );
  NAND2_X1 U6113 ( .A1(n5533), .A2(n4803), .ZN(n4802) );
  NAND2_X1 U6114 ( .A1(n5641), .A2(n4804), .ZN(n9364) );
  NAND2_X1 U6115 ( .A1(n5178), .A2(n8499), .ZN(n5179) );
  NAND2_X1 U6116 ( .A1(n8147), .A2(n8415), .ZN(n8411) );
  NAND2_X1 U6117 ( .A1(n7623), .A2(n5233), .ZN(n7656) );
  NAND2_X1 U6118 ( .A1(n7623), .A2(n5234), .ZN(n5235) );
  NAND2_X1 U6119 ( .A1(n5435), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5285) );
  INV_X1 U6120 ( .A(n8000), .ZN(n7913) );
  OAI21_X2 U6121 ( .B1(n6519), .B2(n6517), .A(n6516), .ZN(n6935) );
  NAND2_X1 U6122 ( .A1(n7575), .A2(n5095), .ZN(n5164) );
  NAND2_X1 U6123 ( .A1(n5551), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5547) );
  NAND2_X1 U6124 ( .A1(n5549), .A2(n5548), .ZN(n5551) );
  NAND2_X1 U6125 ( .A1(n5545), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5549) );
  NAND2_X1 U6126 ( .A1(n4851), .A2(n4850), .ZN(n5058) );
  XNOR2_X1 U6127 ( .A(n4828), .B(SI_2_), .ZN(n5001) );
  NAND2_X1 U6128 ( .A1(n7656), .A2(n7617), .ZN(n7650) );
  NAND2_X1 U6129 ( .A1(n9593), .A2(n4821), .ZN(n4822) );
  OR2_X1 U6130 ( .A1(n5036), .A2(n5576), .ZN(n5023) );
  NAND2_X1 U6131 ( .A1(n5319), .A2(n5318), .ZN(n6864) );
  NAND2_X2 U6132 ( .A1(n8594), .A2(n7455), .ZN(n8642) );
  NAND2_X1 U6133 ( .A1(n4979), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4966) );
  XNOR2_X1 U6134 ( .A(n5921), .B(n7564), .ZN(n6019) );
  NAND2_X2 U6135 ( .A1(n5063), .A2(n5062), .ZN(n5308) );
  NAND2_X1 U6136 ( .A1(n4984), .A2(n4983), .ZN(n4987) );
  INV_X1 U6137 ( .A(n7302), .ZN(n7218) );
  AND2_X1 U6138 ( .A1(n7664), .A2(n7821), .ZN(n7665) );
  XNOR2_X1 U6139 ( .A(n5473), .B(n5472), .ZN(n8419) );
  NAND2_X1 U6140 ( .A1(n6378), .A2(n6377), .ZN(n6382) );
  NAND2_X1 U6141 ( .A1(n7651), .A2(n7655), .ZN(n7652) );
  NAND2_X1 U6142 ( .A1(n5906), .A2(n7655), .ZN(n6229) );
  NOR2_X1 U6143 ( .A1(n6382), .A2(n6407), .ZN(n6403) );
  INV_X1 U6144 ( .A(n5631), .ZN(n9369) );
  XOR2_X1 U6145 ( .A(n8448), .B(n7926), .Z(n4805) );
  OR2_X1 U6146 ( .A1(n9013), .A2(n9012), .ZN(n4806) );
  NAND2_X1 U6147 ( .A1(n8420), .A2(n10015), .ZN(n4807) );
  OR2_X1 U6148 ( .A1(n5675), .A2(n5832), .ZN(n8055) );
  NOR2_X1 U6149 ( .A1(n7898), .A2(n7962), .ZN(n4808) );
  NOR2_X1 U6150 ( .A1(n6906), .A2(n6916), .ZN(n4811) );
  NOR2_X1 U6151 ( .A1(n5112), .A2(n4895), .ZN(n4813) );
  INV_X1 U6152 ( .A(n5233), .ZN(n5234) );
  OR2_X1 U6153 ( .A1(n6030), .A2(n6029), .ZN(n4815) );
  AND2_X1 U6154 ( .A1(n5493), .A2(n7687), .ZN(n4816) );
  AND4_X1 U6155 ( .A1(n4958), .A2(n4957), .A3(n4956), .A4(n4955), .ZN(n4817)
         );
  INV_X1 U6156 ( .A(n7841), .ZN(n8304) );
  INV_X1 U6157 ( .A(n6975), .ZN(n5056) );
  INV_X1 U6158 ( .A(n8191), .ZN(n8194) );
  NOR2_X1 U6159 ( .A1(n9003), .A2(n9002), .ZN(n4818) );
  NOR2_X1 U6160 ( .A1(n7502), .A2(n7501), .ZN(n4819) );
  OR2_X1 U6161 ( .A1(n8474), .A2(n7956), .ZN(n4820) );
  INV_X1 U6162 ( .A(n9192), .ZN(n7347) );
  INV_X1 U6163 ( .A(n8942), .ZN(n6400) );
  INV_X1 U6164 ( .A(n7639), .ZN(n7660) );
  NAND2_X1 U6165 ( .A1(n7641), .A2(n7660), .ZN(n7642) );
  NAND2_X1 U6166 ( .A1(n7690), .A2(n7639), .ZN(n7691) );
  NAND2_X1 U6167 ( .A1(n7737), .A2(n7660), .ZN(n7738) );
  NOR3_X1 U6168 ( .A1(n7760), .A2(n7759), .A3(n7758), .ZN(n7765) );
  AND2_X1 U6169 ( .A1(n8261), .A2(n7770), .ZN(n7771) );
  NAND2_X1 U6170 ( .A1(n7778), .A2(n7811), .ZN(n7779) );
  OAI21_X1 U6171 ( .B1(n7798), .B2(n7660), .A(n7801), .ZN(n7799) );
  AND2_X1 U6172 ( .A1(n7804), .A2(n7810), .ZN(n7805) );
  NOR4_X1 U6173 ( .A1(n7848), .A2(n7847), .A3(n7846), .A4(n7845), .ZN(n7849)
         );
  INV_X1 U6174 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5524) );
  INV_X1 U6175 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n4982) );
  NAND2_X1 U6176 ( .A1(n6648), .A2(n6814), .ZN(n5493) );
  INV_X1 U6177 ( .A(n7820), .ZN(n5479) );
  INV_X1 U6178 ( .A(n8891), .ZN(n6380) );
  AOI21_X1 U6179 ( .B1(n8002), .B2(n8248), .A(n7999), .ZN(n7912) );
  INV_X1 U6180 ( .A(n5390), .ZN(n5389) );
  INV_X1 U6181 ( .A(n5407), .ZN(n5406) );
  INV_X1 U6182 ( .A(n5343), .ZN(n5342) );
  INV_X1 U6183 ( .A(n5377), .ZN(n5375) );
  AOI22_X1 U6184 ( .A1(n8051), .A2(n8390), .B1(n5513), .B2(n8050), .ZN(n5514)
         );
  NAND2_X1 U6185 ( .A1(n4985), .A2(n4982), .ZN(n4986) );
  INV_X1 U6186 ( .A(n8583), .ZN(n7443) );
  NAND2_X1 U6187 ( .A1(n7490), .A2(n7502), .ZN(n8627) );
  INV_X1 U6188 ( .A(n8877), .ZN(n8919) );
  INV_X1 U6189 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n6341) );
  OR2_X1 U6190 ( .A1(n7066), .A2(n8937), .ZN(n7067) );
  NAND2_X1 U6191 ( .A1(n5560), .A2(n4646), .ZN(n5561) );
  AND2_X1 U6192 ( .A1(n5122), .A2(n4899), .ZN(n4900) );
  OR2_X1 U6193 ( .A1(n5602), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n5603) );
  INV_X1 U6194 ( .A(n5274), .ZN(n5272) );
  OR2_X1 U6195 ( .A1(n7905), .A2(n7904), .ZN(n7906) );
  INV_X1 U6196 ( .A(n5292), .ZN(n5290) );
  NAND2_X1 U6197 ( .A1(n5389), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n5396) );
  INV_X1 U6198 ( .A(n5266), .ZN(n5265) );
  INV_X1 U6199 ( .A(n7054), .ZN(n7051) );
  NAND2_X1 U6200 ( .A1(n5406), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5416) );
  AND2_X1 U6201 ( .A1(n5444), .A2(n5443), .ZN(n5445) );
  NAND2_X1 U6202 ( .A1(n5375), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5383) );
  INV_X1 U6203 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n4974) );
  OR2_X1 U6204 ( .A1(n6767), .A2(n6843), .ZN(n6845) );
  NAND2_X1 U6205 ( .A1(n5924), .A2(n5923), .ZN(n5925) );
  NAND2_X1 U6206 ( .A1(n6039), .A2(n6038), .ZN(n6042) );
  AND2_X1 U6207 ( .A1(n7530), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n7551) );
  OR2_X1 U6208 ( .A1(n7385), .A2(n7384), .ZN(n7514) );
  AND2_X1 U6209 ( .A1(n7354), .A2(n7295), .ZN(n7366) );
  AND2_X1 U6210 ( .A1(n4806), .A2(n9108), .ZN(n9011) );
  INV_X1 U6211 ( .A(n9217), .ZN(n7335) );
  NAND2_X1 U6212 ( .A1(n7311), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n7323) );
  NOR2_X1 U6213 ( .A1(n6845), .A2(n6844), .ZN(n7079) );
  OR2_X1 U6214 ( .A1(n6591), .A2(n6590), .ZN(n6767) );
  NAND2_X2 U6215 ( .A1(n5845), .A2(n5844), .ZN(n5876) );
  NAND2_X1 U6216 ( .A1(n5123), .A2(n4900), .ZN(n4902) );
  NAND2_X1 U6217 ( .A1(n4847), .A2(n9574), .ZN(n4850) );
  NAND2_X1 U6218 ( .A1(n5272), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5281) );
  NAND2_X1 U6219 ( .A1(n5333), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5343) );
  INV_X1 U6220 ( .A(n8057), .ZN(n7055) );
  NAND2_X1 U6221 ( .A1(n5357), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n5366) );
  NAND2_X1 U6222 ( .A1(n5290), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5302) );
  INV_X1 U6223 ( .A(n5301), .ZN(n5469) );
  OR2_X1 U6224 ( .A1(n5383), .A2(n9481), .ZN(n5390) );
  OR2_X1 U6225 ( .A1(n5745), .A2(n5744), .ZN(n5772) );
  INV_X1 U6226 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n9540) );
  AND2_X1 U6227 ( .A1(n9964), .A2(n5825), .ZN(n8498) );
  OR3_X1 U6228 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .A3(
        P2_IR_REG_0__SCAN_IN), .ZN(n5009) );
  NOR2_X1 U6229 ( .A1(n7325), .A2(n8643), .ZN(n7354) );
  NAND2_X1 U6230 ( .A1(n8552), .A2(n7522), .ZN(n8604) );
  AND2_X1 U6231 ( .A1(n7174), .A2(n7173), .ZN(n7239) );
  INV_X1 U6232 ( .A(n8650), .ZN(n7569) );
  INV_X1 U6233 ( .A(n9281), .ZN(n9100) );
  NAND2_X1 U6234 ( .A1(n9318), .A2(n7335), .ZN(n7336) );
  NAND2_X1 U6235 ( .A1(n8684), .A2(n8825), .ZN(n9195) );
  INV_X1 U6236 ( .A(n9335), .ZN(n9253) );
  INV_X1 U6237 ( .A(n9906), .ZN(n9664) );
  INV_X1 U6238 ( .A(n6666), .ZN(n6931) );
  AND2_X1 U6239 ( .A1(n6012), .A2(n6011), .ZN(n9242) );
  NAND2_X1 U6240 ( .A1(n4845), .A2(n4844), .ZN(n5048) );
  INV_X1 U6241 ( .A(SI_5_), .ZN(n9568) );
  AND2_X1 U6242 ( .A1(n5462), .A2(n5461), .ZN(n8182) );
  AND4_X1 U6243 ( .A1(n5382), .A2(n5381), .A3(n5380), .A4(n5379), .ZN(n8306)
         );
  AND2_X1 U6244 ( .A1(n5684), .A2(n5683), .ZN(n9930) );
  INV_X1 U6245 ( .A(n8213), .ZN(n8211) );
  AND2_X1 U6246 ( .A1(n8379), .A2(n8487), .ZN(n8503) );
  AND2_X1 U6247 ( .A1(n5218), .A2(n5219), .ZN(n10006) );
  AND2_X1 U6248 ( .A1(n5209), .A2(n5208), .ZN(n9955) );
  NAND2_X1 U6249 ( .A1(n6321), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n6342) );
  AND2_X1 U6250 ( .A1(n8612), .A2(n9664), .ZN(n8670) );
  AND4_X1 U6251 ( .A1(n7317), .A2(n7316), .A3(n7315), .A4(n7314), .ZN(n9244)
         );
  AND4_X1 U6252 ( .A1(n7183), .A2(n7182), .A3(n7181), .A4(n7180), .ZN(n9243)
         );
  NAND2_X1 U6253 ( .A1(n9082), .A2(n9030), .ZN(n9101) );
  AND2_X1 U6254 ( .A1(n9189), .A2(n8823), .ZN(n9214) );
  AND2_X1 U6255 ( .A1(n9814), .A2(n9836), .ZN(n9174) );
  INV_X1 U6256 ( .A(n9895), .ZN(n9897) );
  AND3_X1 U6257 ( .A1(n7005), .A2(n9848), .A3(n6004), .ZN(n6995) );
  XNOR2_X1 U6258 ( .A(n4838), .B(n9458), .ZN(n5033) );
  INV_X1 U6259 ( .A(n9604), .ZN(n9935) );
  INV_X1 U6260 ( .A(n8047), .ZN(n8026) );
  NAND2_X1 U6261 ( .A1(n5824), .A2(n5823), .ZN(n8036) );
  INV_X1 U6262 ( .A(n8182), .ZN(n8051) );
  INV_X1 U6263 ( .A(n8308), .ZN(n8056) );
  INV_X1 U6264 ( .A(n9619), .ZN(n9932) );
  XNOR2_X1 U6265 ( .A(n8411), .B(n7631), .ZN(n7278) );
  AND3_X1 U6266 ( .A1(n7031), .A2(n7030), .A3(n7029), .ZN(n8511) );
  NAND2_X1 U6267 ( .A1(n5516), .A2(n8356), .ZN(n9953) );
  INV_X1 U6268 ( .A(n10033), .ZN(n10030) );
  INV_X1 U6269 ( .A(n10019), .ZN(n10017) );
  OR2_X1 U6270 ( .A1(n9956), .A2(n9955), .ZN(n9959) );
  INV_X1 U6271 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n5574) );
  AND2_X1 U6272 ( .A1(n6096), .A2(n6095), .ZN(n8668) );
  OR2_X1 U6273 ( .A1(n7360), .A2(n7359), .ZN(n9149) );
  AND4_X1 U6274 ( .A1(n5636), .A2(n5635), .A3(n5634), .A4(n5633), .ZN(n9217)
         );
  INV_X1 U6275 ( .A(n6936), .ZN(n8938) );
  OR2_X1 U6276 ( .A1(P1_U3083), .A2(n6256), .ZN(n9785) );
  INV_X1 U6277 ( .A(n9174), .ZN(n9808) );
  INV_X1 U6278 ( .A(n9928), .ZN(n9926) );
  INV_X1 U6279 ( .A(n9916), .ZN(n9914) );
  NAND2_X1 U6280 ( .A1(n4342), .A2(n5522), .ZN(P2_U3267) );
  AOI21_X1 U6281 ( .B1(n9632), .B2(n10019), .A(n5222), .ZN(P2_U3519) );
  NAND2_X2 U6282 ( .A1(n4823), .A2(n4822), .ZN(n4829) );
  MUX2_X1 U6283 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n4829), .Z(n4998) );
  INV_X1 U6284 ( .A(n4824), .ZN(n4825) );
  NAND2_X1 U6285 ( .A1(n4825), .A2(SI_1_), .ZN(n4826) );
  MUX2_X1 U6286 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .S(n4829), .Z(n4830) );
  NAND2_X1 U6287 ( .A1(n4830), .A2(SI_3_), .ZN(n4831) );
  INV_X1 U6288 ( .A(n4831), .ZN(n4832) );
  NAND2_X1 U6289 ( .A1(n5021), .A2(n5022), .ZN(n4835) );
  NAND2_X1 U6290 ( .A1(n4833), .A2(SI_4_), .ZN(n4834) );
  NAND2_X1 U6291 ( .A1(n4835), .A2(n4834), .ZN(n5027) );
  NAND2_X1 U6292 ( .A1(n4836), .A2(SI_5_), .ZN(n4837) );
  NAND2_X1 U6293 ( .A1(n4838), .A2(SI_6_), .ZN(n4839) );
  INV_X1 U6294 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n5601) );
  INV_X1 U6295 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n5609) );
  INV_X1 U6296 ( .A(SI_8_), .ZN(n9562) );
  INV_X1 U6297 ( .A(n4842), .ZN(n4843) );
  NAND2_X1 U6298 ( .A1(n4843), .A2(SI_8_), .ZN(n4844) );
  OAI21_X1 U6299 ( .B1(n5049), .B2(n5048), .A(n4845), .ZN(n5053) );
  INV_X1 U6300 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n5613) );
  INV_X1 U6301 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n4846) );
  INV_X1 U6302 ( .A(SI_9_), .ZN(n9574) );
  INV_X1 U6303 ( .A(n4847), .ZN(n4848) );
  NAND2_X1 U6304 ( .A1(n4848), .A2(SI_9_), .ZN(n4849) );
  NAND2_X1 U6305 ( .A1(n5053), .A2(n5052), .ZN(n4851) );
  INV_X1 U6306 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n5614) );
  INV_X1 U6307 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n5619) );
  INV_X1 U6308 ( .A(SI_10_), .ZN(n4852) );
  INV_X1 U6309 ( .A(n4853), .ZN(n4854) );
  NAND2_X1 U6310 ( .A1(n4854), .A2(SI_10_), .ZN(n4855) );
  NAND2_X1 U6311 ( .A1(n4859), .A2(SI_11_), .ZN(n4860) );
  INV_X1 U6312 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n5646) );
  INV_X1 U6313 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n5644) );
  INV_X1 U6314 ( .A(SI_12_), .ZN(n9469) );
  INV_X1 U6315 ( .A(n4861), .ZN(n4862) );
  NAND2_X1 U6316 ( .A1(n4862), .A2(SI_12_), .ZN(n4863) );
  INV_X1 U6317 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n4866) );
  INV_X1 U6318 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n4865) );
  INV_X1 U6319 ( .A(SI_13_), .ZN(n4867) );
  NAND2_X1 U6320 ( .A1(n4868), .A2(n4867), .ZN(n4871) );
  INV_X1 U6321 ( .A(n4868), .ZN(n4869) );
  NAND2_X1 U6322 ( .A1(n4869), .A2(SI_13_), .ZN(n4870) );
  INV_X1 U6323 ( .A(SI_14_), .ZN(n4873) );
  XNOR2_X1 U6324 ( .A(n4874), .B(n4873), .ZN(n5082) );
  INV_X1 U6325 ( .A(n5082), .ZN(n4876) );
  NAND2_X1 U6326 ( .A1(n4874), .A2(SI_14_), .ZN(n4875) );
  INV_X1 U6327 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n5795) );
  INV_X1 U6328 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n5793) );
  INV_X1 U6329 ( .A(SI_15_), .ZN(n9537) );
  NAND2_X1 U6330 ( .A1(n4877), .A2(n9537), .ZN(n4880) );
  INV_X1 U6331 ( .A(n4877), .ZN(n4878) );
  NAND2_X1 U6332 ( .A1(n4878), .A2(SI_15_), .ZN(n4879) );
  NAND2_X1 U6333 ( .A1(n4880), .A2(n4879), .ZN(n5093) );
  INV_X1 U6334 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n6002) );
  INV_X1 U6335 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n5947) );
  INV_X1 U6336 ( .A(SI_16_), .ZN(n4881) );
  NAND2_X1 U6337 ( .A1(n4882), .A2(n4881), .ZN(n4885) );
  INV_X1 U6338 ( .A(n4882), .ZN(n4883) );
  NAND2_X1 U6339 ( .A1(n4883), .A2(SI_16_), .ZN(n4884) );
  INV_X1 U6340 ( .A(SI_17_), .ZN(n4887) );
  XNOR2_X1 U6341 ( .A(n4892), .B(n4887), .ZN(n5106) );
  INV_X1 U6342 ( .A(n5106), .ZN(n5112) );
  NAND2_X1 U6343 ( .A1(n4888), .A2(SI_18_), .ZN(n4893) );
  INV_X1 U6344 ( .A(n4893), .ZN(n4890) );
  XNOR2_X1 U6345 ( .A(n4888), .B(SI_18_), .ZN(n5116) );
  INV_X1 U6346 ( .A(n5116), .ZN(n4889) );
  NOR2_X1 U6347 ( .A1(n4890), .A2(n4889), .ZN(n4895) );
  NAND2_X1 U6348 ( .A1(n4892), .A2(SI_17_), .ZN(n5114) );
  AND2_X1 U6349 ( .A1(n5114), .A2(n4893), .ZN(n4894) );
  OR2_X1 U6350 ( .A1(n4895), .A2(n4894), .ZN(n5122) );
  INV_X1 U6351 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n6375) );
  INV_X1 U6352 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n6373) );
  INV_X1 U6353 ( .A(SI_19_), .ZN(n9470) );
  NAND2_X1 U6354 ( .A1(n4896), .A2(n9470), .ZN(n4901) );
  INV_X1 U6355 ( .A(n4896), .ZN(n4897) );
  NAND2_X1 U6356 ( .A1(n4897), .A2(SI_19_), .ZN(n4898) );
  NAND2_X1 U6357 ( .A1(n4901), .A2(n4898), .ZN(n5124) );
  INV_X1 U6358 ( .A(n5124), .ZN(n4899) );
  INV_X1 U6359 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n6507) );
  INV_X1 U6360 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7351) );
  INV_X1 U6361 ( .A(SI_20_), .ZN(n9571) );
  NAND2_X1 U6362 ( .A1(n4903), .A2(n9571), .ZN(n4906) );
  INV_X1 U6363 ( .A(n4903), .ZN(n4904) );
  NAND2_X1 U6364 ( .A1(n4904), .A2(SI_20_), .ZN(n4905) );
  XNOR2_X1 U6365 ( .A(n4908), .B(SI_21_), .ZN(n5132) );
  NAND2_X1 U6366 ( .A1(n4908), .A2(SI_21_), .ZN(n4909) );
  INV_X1 U6367 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7865) );
  INV_X1 U6368 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7292) );
  INV_X1 U6369 ( .A(SI_22_), .ZN(n9441) );
  NAND2_X1 U6370 ( .A1(n4910), .A2(n9441), .ZN(n4913) );
  INV_X1 U6371 ( .A(n4910), .ZN(n4911) );
  NAND2_X1 U6372 ( .A1(n4911), .A2(SI_22_), .ZN(n4912) );
  NAND2_X1 U6373 ( .A1(n4913), .A2(n4912), .ZN(n5137) );
  INV_X1 U6374 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n6857) );
  INV_X1 U6375 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7493) );
  INV_X1 U6376 ( .A(SI_23_), .ZN(n4914) );
  NAND2_X1 U6377 ( .A1(n4915), .A2(n4914), .ZN(n4918) );
  INV_X1 U6378 ( .A(n4915), .ZN(n4916) );
  NAND2_X1 U6379 ( .A1(n4916), .A2(SI_23_), .ZN(n4917) );
  AND2_X1 U6380 ( .A1(n4918), .A2(n4917), .ZN(n5141) );
  INV_X1 U6381 ( .A(n5146), .ZN(n4921) );
  INV_X1 U6382 ( .A(SI_24_), .ZN(n4920) );
  XNOR2_X1 U6383 ( .A(n4922), .B(n4920), .ZN(n5145) );
  NAND2_X1 U6384 ( .A1(n4922), .A2(SI_24_), .ZN(n4923) );
  INV_X1 U6385 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7063) );
  INV_X1 U6386 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7527) );
  INV_X1 U6387 ( .A(SI_25_), .ZN(n4924) );
  NAND2_X1 U6388 ( .A1(n4925), .A2(n4924), .ZN(n5153) );
  INV_X1 U6389 ( .A(n4925), .ZN(n4926) );
  NAND2_X1 U6390 ( .A1(n4926), .A2(SI_25_), .ZN(n4927) );
  NAND2_X1 U6391 ( .A1(n5153), .A2(n4927), .ZN(n5149) );
  INV_X1 U6392 ( .A(n5149), .ZN(n4928) );
  INV_X1 U6393 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7191) );
  INV_X1 U6394 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7548) );
  INV_X1 U6395 ( .A(SI_26_), .ZN(n9569) );
  NAND2_X1 U6396 ( .A1(n4930), .A2(n9569), .ZN(n5156) );
  AND2_X1 U6397 ( .A1(n5153), .A2(n5156), .ZN(n4929) );
  INV_X1 U6398 ( .A(n4930), .ZN(n4931) );
  NAND2_X1 U6399 ( .A1(n4931), .A2(SI_26_), .ZN(n5155) );
  INV_X1 U6400 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n7208) );
  INV_X1 U6401 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n7576) );
  INV_X1 U6402 ( .A(SI_27_), .ZN(n9548) );
  NAND2_X1 U6403 ( .A1(n4933), .A2(n9548), .ZN(n4936) );
  INV_X1 U6404 ( .A(n4933), .ZN(n4934) );
  NAND2_X1 U6405 ( .A1(n4934), .A2(SI_27_), .ZN(n4935) );
  AND2_X1 U6406 ( .A1(n4936), .A2(n4935), .ZN(n5161) );
  INV_X1 U6407 ( .A(SI_28_), .ZN(n9452) );
  XNOR2_X1 U6408 ( .A(n4937), .B(n9452), .ZN(n5165) );
  INV_X1 U6409 ( .A(n4937), .ZN(n4938) );
  NAND2_X1 U6410 ( .A1(n4938), .A2(n9452), .ZN(n4939) );
  INV_X1 U6411 ( .A(SI_29_), .ZN(n9551) );
  NAND2_X1 U6412 ( .A1(n5171), .A2(n9551), .ZN(n4941) );
  NAND2_X1 U6413 ( .A1(n4941), .A2(n5169), .ZN(n4943) );
  NAND2_X1 U6414 ( .A1(n4943), .A2(n4942), .ZN(n5175) );
  INV_X1 U6415 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n7938) );
  INV_X1 U6416 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n9371) );
  INV_X1 U6417 ( .A(SI_30_), .ZN(n4944) );
  NAND2_X1 U6418 ( .A1(n4945), .A2(n4944), .ZN(n4948) );
  INV_X1 U6419 ( .A(n4945), .ZN(n4946) );
  NAND2_X1 U6420 ( .A1(n4946), .A2(SI_30_), .ZN(n4947) );
  NAND2_X1 U6421 ( .A1(n4948), .A2(n4947), .ZN(n5174) );
  INV_X1 U6422 ( .A(SI_31_), .ZN(n4949) );
  XNOR2_X1 U6423 ( .A(n4950), .B(n4949), .ZN(n4951) );
  NOR2_X1 U6424 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n4958) );
  NOR2_X1 U6425 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n4957) );
  NOR2_X1 U6426 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n4956) );
  NOR2_X1 U6427 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n4955) );
  NOR2_X1 U6428 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .ZN(
        n4962) );
  NOR2_X1 U6429 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .ZN(
        n4961) );
  INV_X1 U6430 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n4967) );
  INV_X1 U6431 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n4965) );
  XNOR2_X2 U6432 ( .A(n4968), .B(n4967), .ZN(n4994) );
  NAND2_X1 U6433 ( .A1(n9363), .A2(n5095), .ZN(n4970) );
  INV_X1 U6434 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n8535) );
  OR2_X1 U6435 ( .A1(n5036), .A2(n8535), .ZN(n4969) );
  INV_X1 U6436 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n4972) );
  NOR2_X1 U6437 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n4973) );
  NAND2_X1 U6438 ( .A1(n4363), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4978) );
  NAND2_X1 U6439 ( .A1(n4978), .A2(n4974), .ZN(n4975) );
  NAND2_X1 U6440 ( .A1(n4975), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4977) );
  INV_X1 U6441 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n4976) );
  AND2_X1 U6442 ( .A1(n7818), .A2(n8325), .ZN(n7857) );
  INV_X1 U6443 ( .A(n7857), .ZN(n5825) );
  NAND2_X1 U6444 ( .A1(n4980), .A2(n4965), .ZN(n4984) );
  INV_X1 U6445 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n8531) );
  INV_X1 U6446 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n4985) );
  NOR2_X1 U6447 ( .A1(n4985), .A2(n4982), .ZN(n4983) );
  NAND2_X1 U6448 ( .A1(n4987), .A2(n4986), .ZN(n4989) );
  NAND2_X1 U6449 ( .A1(n5301), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n4992) );
  NAND2_X1 U6450 ( .A1(n5465), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n4991) );
  NAND2_X1 U6451 ( .A1(n5508), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n4990) );
  AND3_X1 U6452 ( .A1(n4992), .A2(n4991), .A3(n4990), .ZN(n7630) );
  INV_X1 U6453 ( .A(n5218), .ZN(n7862) );
  NAND2_X1 U6454 ( .A1(n5822), .A2(n7397), .ZN(n8307) );
  INV_X1 U6455 ( .A(P2_B_REG_SCAN_IN), .ZN(n4995) );
  NOR2_X1 U6456 ( .A1(n4994), .A2(n4995), .ZN(n4996) );
  NOR2_X1 U6457 ( .A1(n8307), .A2(n4996), .ZN(n5513) );
  INV_X1 U6458 ( .A(n5513), .ZN(n4997) );
  NOR2_X1 U6459 ( .A1(n7630), .A2(n4997), .ZN(n7275) );
  INV_X1 U6460 ( .A(n9606), .ZN(n5581) );
  XNOR2_X1 U6461 ( .A(n4999), .B(n4998), .ZN(n5917) );
  INV_X1 U6462 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n5582) );
  NAND2_X1 U6463 ( .A1(n5918), .A2(SI_0_), .ZN(n5000) );
  XNOR2_X1 U6464 ( .A(n5000), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n8536) );
  MUX2_X1 U6465 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8536), .S(n5682), .Z(n9963) );
  XNOR2_X1 U6466 ( .A(n5002), .B(n5001), .ZN(n6028) );
  OR2_X1 U6467 ( .A1(n5035), .A2(n6028), .ZN(n5008) );
  OR2_X1 U6468 ( .A1(n5036), .A2(n5574), .ZN(n5007) );
  OR2_X1 U6469 ( .A1(n5003), .A2(n4982), .ZN(n5005) );
  INV_X1 U6470 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5004) );
  XNOR2_X1 U6471 ( .A(n5005), .B(n5004), .ZN(n5691) );
  OR2_X1 U6472 ( .A1(n5682), .A2(n5691), .ZN(n5006) );
  NAND2_X1 U6473 ( .A1(n5894), .A2(n9975), .ZN(n6234) );
  INV_X1 U6474 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5011) );
  NAND2_X1 U6475 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n5009), .ZN(n5010) );
  XNOR2_X1 U6476 ( .A(n5011), .B(n5010), .ZN(n5711) );
  XNOR2_X1 U6477 ( .A(n5014), .B(n5013), .ZN(n6050) );
  OR2_X1 U6478 ( .A1(n5035), .A2(n6050), .ZN(n5016) );
  INV_X1 U6479 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n5575) );
  OR2_X1 U6480 ( .A1(n5036), .A2(n5575), .ZN(n5015) );
  OAI211_X1 U6481 ( .C1(n5682), .C2(n5711), .A(n5016), .B(n5015), .ZN(n6495)
         );
  NAND2_X1 U6482 ( .A1(n5017), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5018) );
  MUX2_X1 U6483 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5018), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n5020) );
  NAND2_X1 U6484 ( .A1(n5020), .A2(n5019), .ZN(n5738) );
  XNOR2_X1 U6485 ( .A(n5021), .B(n5022), .ZN(n6066) );
  OR2_X1 U6486 ( .A1(n5035), .A2(n6066), .ZN(n5024) );
  INV_X1 U6487 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n5576) );
  OAI211_X1 U6488 ( .C1(n5682), .C2(n5738), .A(n5024), .B(n5023), .ZN(n6206)
         );
  NAND2_X1 U6489 ( .A1(n5019), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5025) );
  XNOR2_X1 U6490 ( .A(n5025), .B(P2_IR_REG_5__SCAN_IN), .ZN(n5708) );
  INV_X1 U6491 ( .A(n5708), .ZN(n5728) );
  XNOR2_X1 U6492 ( .A(n5027), .B(n5026), .ZN(n6310) );
  OR2_X1 U6493 ( .A1(n5035), .A2(n6310), .ZN(n5029) );
  INV_X1 U6494 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n5584) );
  OR2_X1 U6495 ( .A1(n5036), .A2(n5584), .ZN(n5028) );
  OAI211_X1 U6496 ( .C1(n5682), .C2(n5728), .A(n5029), .B(n5028), .ZN(n5264)
         );
  OR2_X1 U6497 ( .A1(n5030), .A2(n4982), .ZN(n5032) );
  XNOR2_X1 U6498 ( .A(n5032), .B(n5031), .ZN(n5748) );
  XNOR2_X1 U6499 ( .A(n5034), .B(n5033), .ZN(n6326) );
  OR2_X1 U6500 ( .A1(n5035), .A2(n6326), .ZN(n5038) );
  INV_X1 U6501 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n5585) );
  OR2_X1 U6502 ( .A1(n5036), .A2(n5585), .ZN(n5037) );
  OR2_X1 U6503 ( .A1(n5039), .A2(n4982), .ZN(n5040) );
  XNOR2_X1 U6504 ( .A(n5040), .B(P2_IR_REG_7__SCAN_IN), .ZN(n5761) );
  AOI22_X1 U6505 ( .A1(n5059), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n5647), .B2(
        n5761), .ZN(n5044) );
  XNOR2_X1 U6506 ( .A(n5042), .B(n5041), .ZN(n6351) );
  NAND2_X1 U6507 ( .A1(n6351), .A2(n5095), .ZN(n5043) );
  NAND2_X1 U6508 ( .A1(n5045), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5046) );
  MUX2_X1 U6509 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5046), .S(
        P2_IR_REG_8__SCAN_IN), .Z(n5047) );
  OR2_X1 U6510 ( .A1(n5045), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n5060) );
  AND2_X1 U6511 ( .A1(n5047), .A2(n5060), .ZN(n8073) );
  AOI22_X1 U6512 ( .A1(n5059), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n5647), .B2(
        n8073), .ZN(n5051) );
  XNOR2_X1 U6513 ( .A(n5049), .B(n5048), .ZN(n6579) );
  NAND2_X1 U6514 ( .A1(n6579), .A2(n5095), .ZN(n5050) );
  NAND2_X1 U6515 ( .A1(n5060), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5054) );
  XNOR2_X1 U6516 ( .A(n5054), .B(P2_IR_REG_9__SCAN_IN), .ZN(n8085) );
  AOI22_X1 U6517 ( .A1(n5059), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n5647), .B2(
        n8085), .ZN(n5055) );
  NAND2_X1 U6518 ( .A1(n6829), .A2(n5095), .ZN(n5063) );
  NAND2_X1 U6519 ( .A1(n5065), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5061) );
  XNOR2_X1 U6520 ( .A(n5061), .B(P2_IR_REG_10__SCAN_IN), .ZN(n8100) );
  AOI22_X1 U6521 ( .A1(n5059), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n5647), .B2(
        n8100), .ZN(n5062) );
  INV_X1 U6522 ( .A(n5308), .ZN(n10001) );
  NAND2_X1 U6523 ( .A1(n7069), .A2(n5095), .ZN(n5068) );
  NOR2_X1 U6524 ( .A1(n5065), .A2(P2_IR_REG_10__SCAN_IN), .ZN(n5072) );
  OR2_X1 U6525 ( .A1(n5072), .A2(n4982), .ZN(n5066) );
  XNOR2_X1 U6526 ( .A(n5066), .B(P2_IR_REG_11__SCAN_IN), .ZN(n5781) );
  AOI22_X1 U6527 ( .A1(n5059), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n5647), .B2(
        n5781), .ZN(n5067) );
  INV_X1 U6528 ( .A(n6955), .ZN(n6986) );
  XNOR2_X1 U6529 ( .A(n5070), .B(n5069), .ZN(n7073) );
  NAND2_X1 U6530 ( .A1(n7073), .A2(n5095), .ZN(n5075) );
  INV_X1 U6531 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5071) );
  NAND2_X1 U6532 ( .A1(n5072), .A2(n5071), .ZN(n5078) );
  NAND2_X1 U6533 ( .A1(n5078), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5073) );
  XNOR2_X1 U6534 ( .A(n5073), .B(P2_IR_REG_12__SCAN_IN), .ZN(n6120) );
  AOI22_X1 U6535 ( .A1(n5059), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n5647), .B2(
        n6120), .ZN(n5074) );
  INV_X1 U6536 ( .A(n6927), .ZN(n10009) );
  NAND2_X1 U6537 ( .A1(n6953), .A2(n10009), .ZN(n7033) );
  XNOR2_X1 U6538 ( .A(n5077), .B(n5076), .ZN(n7168) );
  NAND2_X1 U6539 ( .A1(n7168), .A2(n5095), .ZN(n5081) );
  OR2_X1 U6540 ( .A1(n5078), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n5079) );
  NAND2_X1 U6541 ( .A1(n5079), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5085) );
  XNOR2_X1 U6542 ( .A(n5085), .B(P2_IR_REG_13__SCAN_IN), .ZN(n6291) );
  AOI22_X1 U6543 ( .A1(n5059), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n5647), .B2(
        n6291), .ZN(n5080) );
  XNOR2_X1 U6544 ( .A(n5083), .B(n5082), .ZN(n7209) );
  NAND2_X1 U6545 ( .A1(n7209), .A2(n5095), .ZN(n5092) );
  INV_X1 U6546 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5084) );
  NAND2_X1 U6547 ( .A1(n5085), .A2(n5084), .ZN(n5086) );
  NAND2_X1 U6548 ( .A1(n5086), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5089) );
  INV_X1 U6549 ( .A(n5089), .ZN(n5087) );
  NAND2_X1 U6550 ( .A1(n5087), .A2(P2_IR_REG_14__SCAN_IN), .ZN(n5090) );
  INV_X1 U6551 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5088) );
  NAND2_X1 U6552 ( .A1(n5089), .A2(n5088), .ZN(n5096) );
  AOI22_X1 U6553 ( .A1(n5059), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6718), .B2(
        n5647), .ZN(n5091) );
  XNOR2_X1 U6554 ( .A(n5094), .B(n5093), .ZN(n7303) );
  NAND2_X1 U6555 ( .A1(n7303), .A2(n5095), .ZN(n5099) );
  NAND2_X1 U6556 ( .A1(n5096), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5097) );
  XNOR2_X1 U6557 ( .A(n5097), .B(P2_IR_REG_15__SCAN_IN), .ZN(n6876) );
  AOI22_X1 U6558 ( .A1(n6876), .A2(n5647), .B1(n5059), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n5098) );
  INV_X1 U6559 ( .A(n8492), .ZN(n8407) );
  XNOR2_X1 U6560 ( .A(n5101), .B(n5100), .ZN(n7308) );
  NAND2_X1 U6561 ( .A1(n7308), .A2(n5095), .ZN(n5105) );
  NAND2_X1 U6562 ( .A1(n5102), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5103) );
  XNOR2_X1 U6563 ( .A(n5103), .B(P2_IR_REG_16__SCAN_IN), .ZN(n8112) );
  AOI22_X1 U6564 ( .A1(n5059), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n5647), .B2(
        n8112), .ZN(n5104) );
  INV_X1 U6565 ( .A(n8484), .ZN(n8384) );
  NAND2_X1 U6566 ( .A1(n8400), .A2(n8384), .ZN(n8381) );
  NAND2_X1 U6567 ( .A1(n7318), .A2(n5095), .ZN(n5111) );
  INV_X1 U6568 ( .A(n5107), .ZN(n5108) );
  NAND2_X1 U6569 ( .A1(n5108), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5109) );
  XNOR2_X1 U6570 ( .A(n5109), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8125) );
  AOI22_X1 U6571 ( .A1(n5059), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n5647), .B2(
        n8125), .ZN(n5110) );
  NAND2_X1 U6572 ( .A1(n7332), .A2(n5095), .ZN(n5121) );
  INV_X1 U6573 ( .A(n4971), .ZN(n5118) );
  NAND2_X1 U6574 ( .A1(n5118), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5119) );
  XNOR2_X1 U6575 ( .A(n5119), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8135) );
  AOI22_X1 U6576 ( .A1(n5059), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n5647), .B2(
        n8135), .ZN(n5120) );
  NAND2_X1 U6577 ( .A1(n5123), .A2(n5122), .ZN(n5125) );
  NAND2_X1 U6578 ( .A1(n7337), .A2(n5095), .ZN(n5127) );
  AOI22_X1 U6579 ( .A1(n5059), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n9946), .B2(
        n5647), .ZN(n5126) );
  XNOR2_X1 U6580 ( .A(n5129), .B(n5128), .ZN(n7350) );
  NAND2_X1 U6581 ( .A1(n7350), .A2(n5095), .ZN(n5131) );
  OR2_X1 U6582 ( .A1(n5036), .A2(n6507), .ZN(n5130) );
  INV_X1 U6583 ( .A(n5132), .ZN(n5133) );
  XNOR2_X1 U6584 ( .A(n5134), .B(n5133), .ZN(n7362) );
  NAND2_X1 U6585 ( .A1(n7362), .A2(n5095), .ZN(n5136) );
  INV_X1 U6586 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n6544) );
  OR2_X1 U6587 ( .A1(n5036), .A2(n6544), .ZN(n5135) );
  INV_X1 U6588 ( .A(n8459), .ZN(n8291) );
  XNOR2_X1 U6589 ( .A(n5138), .B(n5137), .ZN(n7291) );
  NAND2_X1 U6590 ( .A1(n7291), .A2(n5095), .ZN(n5140) );
  OR2_X1 U6591 ( .A1(n5036), .A2(n7865), .ZN(n5139) );
  INV_X1 U6592 ( .A(n8454), .ZN(n8272) );
  NAND2_X1 U6593 ( .A1(n8287), .A2(n8272), .ZN(n8267) );
  NAND2_X1 U6594 ( .A1(n7492), .A2(n5095), .ZN(n5144) );
  OR2_X1 U6595 ( .A1(n5036), .A2(n6857), .ZN(n5143) );
  OR2_X2 U6596 ( .A1(n8267), .A2(n8448), .ZN(n8253) );
  NAND2_X1 U6597 ( .A1(n7510), .A2(n5095), .ZN(n5148) );
  INV_X1 U6598 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7011) );
  OR2_X1 U6599 ( .A1(n5036), .A2(n7011), .ZN(n5147) );
  XNOR2_X1 U6600 ( .A(n5150), .B(n5149), .ZN(n7526) );
  NAND2_X1 U6601 ( .A1(n7526), .A2(n5095), .ZN(n5152) );
  OR2_X1 U6602 ( .A1(n5036), .A2(n7063), .ZN(n5151) );
  INV_X1 U6603 ( .A(n8439), .ZN(n8224) );
  AND2_X1 U6604 ( .A1(n5156), .A2(n5155), .ZN(n5157) );
  NAND2_X1 U6605 ( .A1(n7547), .A2(n5095), .ZN(n5160) );
  OR2_X1 U6606 ( .A1(n5036), .A2(n7191), .ZN(n5159) );
  INV_X1 U6607 ( .A(n8433), .ZN(n8204) );
  OR2_X1 U6608 ( .A1(n5036), .A2(n7208), .ZN(n5163) );
  INV_X1 U6609 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n7399) );
  OR2_X1 U6610 ( .A1(n5036), .A2(n7399), .ZN(n5167) );
  XNOR2_X1 U6611 ( .A(n5169), .B(n9551), .ZN(n5170) );
  NAND2_X1 U6612 ( .A1(n8768), .A2(n5095), .ZN(n5173) );
  INV_X1 U6613 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n7401) );
  OR2_X1 U6614 ( .A1(n5036), .A2(n7401), .ZN(n5172) );
  NAND2_X1 U6615 ( .A1(n8677), .A2(n5095), .ZN(n5177) );
  OR2_X1 U6616 ( .A1(n5036), .A2(n7938), .ZN(n5176) );
  INV_X1 U6617 ( .A(n7278), .ZN(n5178) );
  NOR4_X1 U6618 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n5184) );
  NOR4_X1 U6619 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n5183) );
  NOR4_X1 U6620 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n5182) );
  NOR4_X1 U6621 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n5181) );
  NAND4_X1 U6622 ( .A1(n5184), .A2(n5183), .A3(n5182), .A4(n5181), .ZN(n5211)
         );
  NOR2_X1 U6623 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .ZN(
        n5188) );
  NOR4_X1 U6624 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n5187) );
  NOR4_X1 U6625 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n5186) );
  NOR4_X1 U6626 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n5185) );
  NAND4_X1 U6627 ( .A1(n5188), .A2(n5187), .A3(n5186), .A4(n5185), .ZN(n5210)
         );
  INV_X1 U6628 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5203) );
  INV_X1 U6629 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5205) );
  NAND3_X1 U6630 ( .A1(n5200), .A2(n5203), .A3(n5205), .ZN(n5189) );
  NOR2_X1 U6631 ( .A1(n5190), .A2(n5189), .ZN(n5195) );
  INV_X1 U6632 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5191) );
  NAND2_X1 U6633 ( .A1(n5195), .A2(n5191), .ZN(n5198) );
  NAND2_X1 U6634 ( .A1(n5198), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5192) );
  MUX2_X1 U6635 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5192), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n5194) );
  NAND2_X1 U6636 ( .A1(n5194), .A2(n5193), .ZN(n7193) );
  INV_X1 U6637 ( .A(n7193), .ZN(n5209) );
  INV_X1 U6638 ( .A(n5195), .ZN(n5196) );
  NAND2_X1 U6639 ( .A1(n5196), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5197) );
  MUX2_X1 U6640 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5197), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n5199) );
  NAND2_X1 U6641 ( .A1(n5199), .A2(n5198), .ZN(n7062) );
  NAND2_X1 U6642 ( .A1(n5201), .A2(n5200), .ZN(n5202) );
  NAND2_X1 U6643 ( .A1(n5202), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5214) );
  NAND2_X1 U6644 ( .A1(n5214), .A2(n5203), .ZN(n5204) );
  NAND2_X1 U6645 ( .A1(n5204), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5206) );
  XNOR2_X1 U6646 ( .A(n5206), .B(n5205), .ZN(n7013) );
  XNOR2_X1 U6647 ( .A(n7013), .B(P2_B_REG_SCAN_IN), .ZN(n5207) );
  NAND2_X1 U6648 ( .A1(n7062), .A2(n5207), .ZN(n5208) );
  OAI21_X1 U6649 ( .B1(n5211), .B2(n5210), .A(n9955), .ZN(n5821) );
  NOR2_X1 U6650 ( .A1(n7193), .A2(n7062), .ZN(n5213) );
  INV_X1 U6651 ( .A(n7013), .ZN(n5212) );
  NAND2_X1 U6652 ( .A1(n5213), .A2(n5212), .ZN(n5835) );
  XNOR2_X1 U6653 ( .A(n5214), .B(P2_IR_REG_23__SCAN_IN), .ZN(n5832) );
  NOR2_X1 U6654 ( .A1(n5832), .A2(P2_U3152), .ZN(n9961) );
  NAND2_X1 U6655 ( .A1(n5835), .A2(n9961), .ZN(n9956) );
  AND2_X1 U6656 ( .A1(n5822), .A2(n5825), .ZN(n5833) );
  NOR2_X1 U6657 ( .A1(n9956), .A2(n5833), .ZN(n5215) );
  NAND2_X1 U6658 ( .A1(n5821), .A2(n5215), .ZN(n5474) );
  INV_X1 U6659 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n9960) );
  NAND2_X1 U6660 ( .A1(n9955), .A2(n9960), .ZN(n5217) );
  AND2_X1 U6661 ( .A1(n7193), .A2(n7062), .ZN(n9962) );
  INV_X1 U6662 ( .A(n9962), .ZN(n5216) );
  NAND2_X1 U6663 ( .A1(n5217), .A2(n5216), .ZN(n5819) );
  AND2_X1 U6664 ( .A1(n7818), .A2(n9946), .ZN(n5219) );
  NAND2_X1 U6665 ( .A1(n10006), .A2(n6543), .ZN(n5828) );
  NAND2_X1 U6666 ( .A1(n5819), .A2(n5828), .ZN(n5220) );
  NOR2_X1 U6667 ( .A1(n5474), .A2(n5220), .ZN(n6503) );
  INV_X1 U6668 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n9957) );
  AND2_X1 U6669 ( .A1(n7013), .A2(n7193), .ZN(n9958) );
  AOI21_X1 U6670 ( .B1(n9955), .B2(n9957), .A(n9958), .ZN(n6502) );
  INV_X1 U6671 ( .A(n6502), .ZN(n5221) );
  AND2_X2 U6672 ( .A1(n6503), .A2(n5221), .ZN(n10019) );
  NOR2_X1 U6673 ( .A1(n10019), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n5222) );
  NAND2_X1 U6674 ( .A1(n5301), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5228) );
  NAND2_X1 U6675 ( .A1(n4314), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n5227) );
  NAND2_X1 U6676 ( .A1(n5435), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5226) );
  NAND2_X1 U6677 ( .A1(n5368), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5225) );
  AND2_X1 U6678 ( .A1(n5887), .A2(n9963), .ZN(n5893) );
  NAND2_X1 U6679 ( .A1(n5435), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5232) );
  NAND2_X1 U6680 ( .A1(n5368), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5231) );
  NAND2_X1 U6681 ( .A1(n5301), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5230) );
  NAND2_X1 U6682 ( .A1(n4313), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n5229) );
  NAND2_X1 U6683 ( .A1(n5893), .A2(n5235), .ZN(n5237) );
  NAND2_X1 U6684 ( .A1(n5808), .A2(n5233), .ZN(n5236) );
  NAND2_X1 U6685 ( .A1(n5435), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5241) );
  NAND2_X1 U6686 ( .A1(n4313), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n5240) );
  NAND2_X1 U6687 ( .A1(n5301), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5239) );
  NAND2_X1 U6688 ( .A1(n5368), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5238) );
  INV_X1 U6689 ( .A(n9975), .ZN(n5914) );
  NAND2_X1 U6690 ( .A1(n5818), .A2(n9975), .ZN(n7658) );
  NAND2_X1 U6691 ( .A1(n5913), .A2(n7820), .ZN(n5244) );
  NAND2_X1 U6692 ( .A1(n5242), .A2(n9975), .ZN(n5243) );
  NAND2_X1 U6693 ( .A1(n5244), .A2(n5243), .ZN(n6227) );
  NAND2_X1 U6694 ( .A1(n5301), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5248) );
  NAND2_X1 U6695 ( .A1(n4314), .A2(n9534), .ZN(n5247) );
  NAND2_X1 U6696 ( .A1(n5435), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5246) );
  NAND2_X1 U6697 ( .A1(n5368), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5245) );
  INV_X1 U6698 ( .A(n7821), .ZN(n6228) );
  NAND2_X1 U6699 ( .A1(n6227), .A2(n6228), .ZN(n6226) );
  INV_X1 U6700 ( .A(n8068), .ZN(n5481) );
  INV_X1 U6701 ( .A(n6495), .ZN(n7670) );
  NAND2_X1 U6702 ( .A1(n5481), .A2(n7670), .ZN(n5249) );
  NAND2_X1 U6703 ( .A1(n5301), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5254) );
  XNOR2_X1 U6704 ( .A(P2_REG3_REG_4__SCAN_IN), .B(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n6203) );
  INV_X1 U6705 ( .A(n6203), .ZN(n5250) );
  NAND2_X1 U6706 ( .A1(n4314), .A2(n5250), .ZN(n5253) );
  NAND2_X1 U6707 ( .A1(n5435), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5252) );
  NAND2_X1 U6708 ( .A1(n5368), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5251) );
  NAND4_X1 U6709 ( .A1(n5254), .A2(n5253), .A3(n5252), .A4(n5251), .ZN(n8067)
         );
  INV_X1 U6710 ( .A(n8067), .ZN(n6247) );
  NAND2_X1 U6711 ( .A1(n6247), .A2(n6206), .ZN(n7645) );
  NAND2_X1 U6712 ( .A1(n8067), .A2(n9981), .ZN(n7672) );
  INV_X1 U6713 ( .A(n7822), .ZN(n6130) );
  NAND2_X1 U6714 ( .A1(n6247), .A2(n9981), .ZN(n5255) );
  NAND2_X1 U6715 ( .A1(n5301), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5263) );
  INV_X1 U6716 ( .A(n5256), .ZN(n5258) );
  INV_X1 U6717 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5257) );
  NAND2_X1 U6718 ( .A1(n5258), .A2(n5257), .ZN(n5259) );
  AND2_X1 U6719 ( .A1(n5266), .A2(n5259), .ZN(n9943) );
  NAND2_X1 U6720 ( .A1(n4314), .A2(n9943), .ZN(n5262) );
  NAND2_X1 U6721 ( .A1(n5368), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5261) );
  NAND2_X1 U6722 ( .A1(n5435), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5260) );
  INV_X1 U6723 ( .A(n8065), .ZN(n6460) );
  INV_X1 U6724 ( .A(n5264), .ZN(n6248) );
  NAND2_X1 U6725 ( .A1(n8065), .A2(n6248), .ZN(n7674) );
  NAND2_X1 U6726 ( .A1(n7646), .A2(n7674), .ZN(n7824) );
  INV_X1 U6727 ( .A(n6452), .ZN(n5280) );
  NAND2_X1 U6728 ( .A1(n5465), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5271) );
  INV_X1 U6729 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n5699) );
  NAND2_X1 U6730 ( .A1(n5266), .A2(n5699), .ZN(n5267) );
  AND2_X1 U6731 ( .A1(n5274), .A2(n5267), .ZN(n6464) );
  NAND2_X1 U6732 ( .A1(n4314), .A2(n6464), .ZN(n5270) );
  NAND2_X1 U6733 ( .A1(n5435), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5269) );
  NAND2_X1 U6734 ( .A1(n5301), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5268) );
  NAND2_X1 U6735 ( .A1(n8064), .A2(n6472), .ZN(n5483) );
  INV_X1 U6736 ( .A(n5483), .ZN(n6453) );
  NAND2_X1 U6737 ( .A1(n5301), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5279) );
  INV_X1 U6738 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5273) );
  NAND2_X1 U6739 ( .A1(n5274), .A2(n5273), .ZN(n5275) );
  AND2_X1 U6740 ( .A1(n5281), .A2(n5275), .ZN(n6670) );
  NAND2_X1 U6741 ( .A1(n4314), .A2(n6670), .ZN(n5278) );
  NAND2_X1 U6742 ( .A1(n5368), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5277) );
  NAND2_X1 U6743 ( .A1(n5435), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5276) );
  INV_X1 U6744 ( .A(n8063), .ZN(n6459) );
  NAND2_X1 U6745 ( .A1(n6459), .A2(n6625), .ZN(n7702) );
  INV_X1 U6746 ( .A(n6625), .ZN(n6673) );
  NAND2_X1 U6747 ( .A1(n8063), .A2(n6673), .ZN(n7683) );
  NAND2_X1 U6748 ( .A1(n5280), .A2(n4328), .ZN(n6613) );
  NAND2_X1 U6749 ( .A1(n5301), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5284) );
  NAND2_X1 U6750 ( .A1(n5281), .A2(n9557), .ZN(n5282) );
  AND2_X1 U6751 ( .A1(n5292), .A2(n5282), .ZN(n6813) );
  NAND2_X1 U6752 ( .A1(n4314), .A2(n6813), .ZN(n5283) );
  NAND2_X1 U6753 ( .A1(n5465), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5286) );
  NAND2_X1 U6754 ( .A1(n8062), .A2(n9995), .ZN(n7687) );
  INV_X1 U6755 ( .A(n4816), .ZN(n7684) );
  OR2_X1 U6756 ( .A1(n7678), .A2(n6615), .ZN(n6614) );
  NAND2_X1 U6757 ( .A1(n6459), .A2(n6673), .ZN(n5288) );
  AND2_X1 U6758 ( .A1(n6614), .A2(n5288), .ZN(n6806) );
  AND2_X1 U6759 ( .A1(n7684), .A2(n6806), .ZN(n5289) );
  NAND2_X1 U6760 ( .A1(n6613), .A2(n5289), .ZN(n6809) );
  NAND2_X1 U6761 ( .A1(n6814), .A2(n8062), .ZN(n6780) );
  NAND2_X1 U6762 ( .A1(n5301), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5297) );
  INV_X1 U6763 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5291) );
  NAND2_X1 U6764 ( .A1(n5292), .A2(n5291), .ZN(n5293) );
  AND2_X1 U6765 ( .A1(n5302), .A2(n5293), .ZN(n6789) );
  NAND2_X1 U6766 ( .A1(n4314), .A2(n6789), .ZN(n5296) );
  NAND2_X1 U6767 ( .A1(n5368), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5295) );
  NAND2_X1 U6768 ( .A1(n5435), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5294) );
  NAND4_X1 U6769 ( .A1(n5297), .A2(n5296), .A3(n5295), .A4(n5294), .ZN(n8061)
         );
  INV_X1 U6770 ( .A(n8061), .ZN(n6682) );
  INV_X1 U6771 ( .A(n7689), .ZN(n7695) );
  NAND2_X1 U6772 ( .A1(n6975), .A2(n6682), .ZN(n7696) );
  INV_X1 U6773 ( .A(n7828), .ZN(n5298) );
  AND2_X1 U6774 ( .A1(n6780), .A2(n5298), .ZN(n5299) );
  NAND2_X1 U6775 ( .A1(n6809), .A2(n5299), .ZN(n6781) );
  OR2_X1 U6776 ( .A1(n6975), .A2(n8061), .ZN(n5300) );
  NAND2_X1 U6777 ( .A1(n5301), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5307) );
  NAND2_X1 U6778 ( .A1(n5302), .A2(n9540), .ZN(n5303) );
  AND2_X1 U6779 ( .A1(n5312), .A2(n5303), .ZN(n6742) );
  NAND2_X1 U6780 ( .A1(n4314), .A2(n6742), .ZN(n5306) );
  NAND2_X1 U6781 ( .A1(n5435), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5305) );
  NAND2_X1 U6782 ( .A1(n5368), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5304) );
  NAND4_X1 U6783 ( .A1(n5307), .A2(n5306), .A3(n5305), .A4(n5304), .ZN(n8060)
         );
  INV_X1 U6784 ( .A(n8060), .ZN(n6801) );
  AND2_X1 U6785 ( .A1(n5308), .A2(n6801), .ZN(n7699) );
  NAND2_X1 U6786 ( .A1(n5308), .A2(n8060), .ZN(n5309) );
  NAND2_X1 U6787 ( .A1(n5301), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5317) );
  INV_X1 U6788 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n5311) );
  NAND2_X1 U6789 ( .A1(n5312), .A2(n5311), .ZN(n5313) );
  AND2_X1 U6790 ( .A1(n5320), .A2(n5313), .ZN(n6984) );
  NAND2_X1 U6791 ( .A1(n4314), .A2(n6984), .ZN(n5316) );
  NAND2_X1 U6792 ( .A1(n5435), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5315) );
  NAND2_X1 U6793 ( .A1(n5465), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n5314) );
  NAND4_X1 U6794 ( .A1(n5317), .A2(n5316), .A3(n5315), .A4(n5314), .ZN(n8059)
         );
  INV_X1 U6795 ( .A(n8059), .ZN(n6924) );
  OR2_X1 U6796 ( .A1(n6955), .A2(n6924), .ZN(n7704) );
  NAND2_X1 U6797 ( .A1(n6955), .A2(n6924), .ZN(n7714) );
  NAND2_X1 U6798 ( .A1(n7704), .A2(n7714), .ZN(n7830) );
  NAND2_X1 U6799 ( .A1(n6955), .A2(n8059), .ZN(n5318) );
  NAND2_X1 U6800 ( .A1(n5301), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5325) );
  INV_X1 U6801 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n9531) );
  NAND2_X1 U6802 ( .A1(n5320), .A2(n9531), .ZN(n5321) );
  AND2_X1 U6803 ( .A1(n5327), .A2(n5321), .ZN(n6921) );
  NAND2_X1 U6804 ( .A1(n4314), .A2(n6921), .ZN(n5324) );
  NAND2_X1 U6805 ( .A1(n5435), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5323) );
  NAND2_X1 U6806 ( .A1(n5368), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5322) );
  NAND4_X1 U6807 ( .A1(n5325), .A2(n5324), .A3(n5323), .A4(n5322), .ZN(n8058)
         );
  INV_X1 U6808 ( .A(n8058), .ZN(n6908) );
  OR2_X1 U6809 ( .A1(n6927), .A2(n6908), .ZN(n7716) );
  NAND2_X1 U6810 ( .A1(n6927), .A2(n6908), .ZN(n7715) );
  NAND2_X1 U6811 ( .A1(n7716), .A2(n7715), .ZN(n7831) );
  INV_X1 U6812 ( .A(n7831), .ZN(n6863) );
  OAI22_X1 U6813 ( .A1(n6864), .A2(n6863), .B1(n6927), .B2(n8058), .ZN(n7024)
         );
  NAND2_X1 U6814 ( .A1(n5301), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n5332) );
  INV_X1 U6815 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5326) );
  NAND2_X1 U6816 ( .A1(n5327), .A2(n5326), .ZN(n5328) );
  AND2_X1 U6817 ( .A1(n5334), .A2(n5328), .ZN(n7036) );
  NAND2_X1 U6818 ( .A1(n4314), .A2(n7036), .ZN(n5331) );
  NAND2_X1 U6819 ( .A1(n5508), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5330) );
  NAND2_X1 U6820 ( .A1(n5465), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n5329) );
  NAND4_X1 U6821 ( .A1(n5332), .A2(n5331), .A3(n5330), .A4(n5329), .ZN(n8057)
         );
  XNOR2_X1 U6822 ( .A(n8505), .B(n7055), .ZN(n7721) );
  NAND2_X1 U6823 ( .A1(n8505), .A2(n8057), .ZN(n7723) );
  NAND2_X1 U6824 ( .A1(n5301), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n5339) );
  INV_X1 U6825 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n9465) );
  NAND2_X1 U6826 ( .A1(n5334), .A2(n9465), .ZN(n5335) );
  AND2_X1 U6827 ( .A1(n5343), .A2(n5335), .ZN(n7058) );
  NAND2_X1 U6828 ( .A1(n4314), .A2(n7058), .ZN(n5338) );
  NAND2_X1 U6829 ( .A1(n5435), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5337) );
  NAND2_X1 U6830 ( .A1(n5465), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n5336) );
  NAND4_X1 U6831 ( .A1(n5339), .A2(n5338), .A3(n5337), .A4(n5336), .ZN(n8391)
         );
  INV_X1 U6832 ( .A(n8391), .ZN(n7111) );
  NAND2_X1 U6833 ( .A1(n8497), .A2(n7111), .ZN(n7724) );
  OR2_X1 U6834 ( .A1(n8497), .A2(n8391), .ZN(n5340) );
  NAND2_X1 U6835 ( .A1(n5341), .A2(n5340), .ZN(n8398) );
  NAND2_X1 U6836 ( .A1(n5301), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n5348) );
  INV_X1 U6837 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n7108) );
  NAND2_X1 U6838 ( .A1(n5343), .A2(n7108), .ZN(n5344) );
  AND2_X1 U6839 ( .A1(n5350), .A2(n5344), .ZN(n8403) );
  NAND2_X1 U6840 ( .A1(n4314), .A2(n8403), .ZN(n5347) );
  NAND2_X1 U6841 ( .A1(n5508), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5346) );
  NAND2_X1 U6842 ( .A1(n5465), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n5345) );
  NAND4_X1 U6843 ( .A1(n5348), .A2(n5347), .A3(n5346), .A4(n5345), .ZN(n8373)
         );
  INV_X1 U6844 ( .A(n8373), .ZN(n7981) );
  OR2_X1 U6845 ( .A1(n8492), .A2(n7981), .ZN(n5502) );
  NAND2_X1 U6846 ( .A1(n8492), .A2(n7981), .ZN(n7728) );
  NAND2_X1 U6847 ( .A1(n5502), .A2(n7728), .ZN(n8397) );
  NAND2_X1 U6848 ( .A1(n8398), .A2(n8397), .ZN(n8396) );
  OR2_X1 U6849 ( .A1(n8492), .A2(n8373), .ZN(n5349) );
  NAND2_X1 U6850 ( .A1(n5301), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n5355) );
  INV_X1 U6851 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n9444) );
  NAND2_X1 U6852 ( .A1(n5350), .A2(n9444), .ZN(n5351) );
  AND2_X1 U6853 ( .A1(n5359), .A2(n5351), .ZN(n8382) );
  NAND2_X1 U6854 ( .A1(n4314), .A2(n8382), .ZN(n5354) );
  NAND2_X1 U6855 ( .A1(n5508), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5353) );
  NAND2_X1 U6856 ( .A1(n5465), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n5352) );
  NAND4_X1 U6857 ( .A1(n5355), .A2(n5354), .A3(n5353), .A4(n5352), .ZN(n8393)
         );
  INV_X1 U6858 ( .A(n8393), .ZN(n7110) );
  OR2_X1 U6859 ( .A1(n8484), .A2(n7110), .ZN(n7730) );
  NAND2_X1 U6860 ( .A1(n8484), .A2(n7110), .ZN(n7729) );
  NAND2_X1 U6861 ( .A1(n7730), .A2(n7729), .ZN(n7745) );
  NAND2_X1 U6862 ( .A1(n8484), .A2(n8393), .ZN(n5356) );
  NAND2_X1 U6863 ( .A1(n5301), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n5364) );
  INV_X1 U6864 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n5358) );
  NAND2_X1 U6865 ( .A1(n5359), .A2(n5358), .ZN(n5360) );
  AND2_X1 U6866 ( .A1(n5366), .A2(n5360), .ZN(n8355) );
  NAND2_X1 U6867 ( .A1(n4314), .A2(n8355), .ZN(n5363) );
  NAND2_X1 U6868 ( .A1(n5465), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n5362) );
  NAND2_X1 U6869 ( .A1(n5508), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5361) );
  NAND4_X1 U6870 ( .A1(n5364), .A2(n5363), .A3(n5362), .A4(n5361), .ZN(n8372)
         );
  INV_X1 U6871 ( .A(n8372), .ZN(n8031) );
  NAND2_X1 U6872 ( .A1(n8480), .A2(n8031), .ZN(n7737) );
  OR2_X1 U6873 ( .A1(n8480), .A2(n8372), .ZN(n5365) );
  NAND2_X1 U6874 ( .A1(n5301), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n5372) );
  INV_X1 U6875 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n9454) );
  NAND2_X1 U6876 ( .A1(n5366), .A2(n9454), .ZN(n5367) );
  AND2_X1 U6877 ( .A1(n5377), .A2(n5367), .ZN(n8336) );
  NAND2_X1 U6878 ( .A1(n4314), .A2(n8336), .ZN(n5371) );
  NAND2_X1 U6879 ( .A1(n5508), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n5370) );
  NAND2_X1 U6880 ( .A1(n5368), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n5369) );
  NAND4_X1 U6881 ( .A1(n5372), .A2(n5371), .A3(n5370), .A4(n5369), .ZN(n8318)
         );
  NAND2_X1 U6882 ( .A1(n8474), .A2(n8318), .ZN(n5373) );
  OR2_X1 U6883 ( .A1(n8474), .A2(n8318), .ZN(n5374) );
  INV_X1 U6884 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n5376) );
  NAND2_X1 U6885 ( .A1(n5377), .A2(n5376), .ZN(n5378) );
  NAND2_X1 U6886 ( .A1(n5383), .A2(n5378), .ZN(n8326) );
  OR2_X1 U6887 ( .A1(n4312), .A2(n8326), .ZN(n5382) );
  NAND2_X1 U6888 ( .A1(n5301), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n5381) );
  NAND2_X1 U6889 ( .A1(n5465), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n5380) );
  NAND2_X1 U6890 ( .A1(n5508), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n5379) );
  INV_X1 U6891 ( .A(n8306), .ZN(n8341) );
  INV_X1 U6892 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n9481) );
  NAND2_X1 U6893 ( .A1(n5383), .A2(n9481), .ZN(n5384) );
  NAND2_X1 U6894 ( .A1(n5390), .A2(n5384), .ZN(n8299) );
  AOI22_X1 U6895 ( .A1(n5301), .A2(P2_REG1_REG_20__SCAN_IN), .B1(n5508), .B2(
        P2_REG0_REG_20__SCAN_IN), .ZN(n5386) );
  NAND2_X1 U6896 ( .A1(n5465), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n5385) );
  OAI211_X1 U6897 ( .C1(n8299), .C2(n4312), .A(n5386), .B(n5385), .ZN(n8319)
         );
  INV_X1 U6898 ( .A(n8319), .ZN(n7966) );
  NAND2_X1 U6899 ( .A1(n8464), .A2(n7966), .ZN(n7761) );
  NAND2_X1 U6900 ( .A1(n8297), .A2(n8304), .ZN(n5388) );
  OR2_X1 U6901 ( .A1(n8302), .A2(n7966), .ZN(n5387) );
  INV_X1 U6902 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n9455) );
  NAND2_X1 U6903 ( .A1(n5390), .A2(n9455), .ZN(n5391) );
  NAND2_X1 U6904 ( .A1(n5396), .A2(n5391), .ZN(n8288) );
  OR2_X1 U6905 ( .A1(n8288), .A2(n4312), .ZN(n5394) );
  AOI22_X1 U6906 ( .A1(n5301), .A2(P2_REG1_REG_21__SCAN_IN), .B1(n5435), .B2(
        P2_REG0_REG_21__SCAN_IN), .ZN(n5393) );
  NAND2_X1 U6907 ( .A1(n5465), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n5392) );
  AND2_X1 U6908 ( .A1(n8459), .A2(n8056), .ZN(n5395) );
  INV_X1 U6909 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n8021) );
  NAND2_X1 U6910 ( .A1(n5396), .A2(n8021), .ZN(n5397) );
  AND2_X1 U6911 ( .A1(n5407), .A2(n5397), .ZN(n8270) );
  NAND2_X1 U6912 ( .A1(n8270), .A2(n4314), .ZN(n5403) );
  INV_X1 U6913 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n5400) );
  NAND2_X1 U6914 ( .A1(n5508), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n5399) );
  NAND2_X1 U6915 ( .A1(n5465), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n5398) );
  OAI211_X1 U6916 ( .C1(n5469), .C2(n5400), .A(n5399), .B(n5398), .ZN(n5401)
         );
  INV_X1 U6917 ( .A(n5401), .ZN(n5402) );
  NAND2_X1 U6918 ( .A1(n8454), .A2(n8247), .ZN(n7769) );
  NAND2_X1 U6919 ( .A1(n8266), .A2(n8273), .ZN(n5405) );
  INV_X1 U6920 ( .A(n8247), .ZN(n8283) );
  OR2_X1 U6921 ( .A1(n8454), .A2(n8283), .ZN(n5404) );
  NAND2_X1 U6922 ( .A1(n5405), .A2(n5404), .ZN(n8260) );
  INV_X1 U6923 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n7947) );
  NAND2_X1 U6924 ( .A1(n5407), .A2(n7947), .ZN(n5408) );
  NAND2_X1 U6925 ( .A1(n5416), .A2(n5408), .ZN(n8254) );
  OR2_X1 U6926 ( .A1(n8254), .A2(n4312), .ZN(n5414) );
  INV_X1 U6927 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n5411) );
  NAND2_X1 U6928 ( .A1(n5465), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n5410) );
  NAND2_X1 U6929 ( .A1(n5435), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n5409) );
  OAI211_X1 U6930 ( .C1(n5469), .C2(n5411), .A(n5410), .B(n5409), .ZN(n5412)
         );
  INV_X1 U6931 ( .A(n5412), .ZN(n5413) );
  NAND2_X1 U6932 ( .A1(n5414), .A2(n5413), .ZN(n8229) );
  NAND2_X1 U6933 ( .A1(n8448), .A2(n8229), .ZN(n5415) );
  INV_X1 U6934 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n8005) );
  NAND2_X1 U6935 ( .A1(n5416), .A2(n8005), .ZN(n5417) );
  NAND2_X1 U6936 ( .A1(n5425), .A2(n5417), .ZN(n8233) );
  OR2_X1 U6937 ( .A1(n8233), .A2(n4312), .ZN(n5423) );
  INV_X1 U6938 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n5420) );
  NAND2_X1 U6939 ( .A1(n5465), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n5419) );
  NAND2_X1 U6940 ( .A1(n5508), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n5418) );
  OAI211_X1 U6941 ( .C1(n5469), .C2(n5420), .A(n5419), .B(n5418), .ZN(n5421)
         );
  INV_X1 U6942 ( .A(n5421), .ZN(n5422) );
  NAND2_X1 U6943 ( .A1(n8442), .A2(n8248), .ZN(n7777) );
  INV_X1 U6944 ( .A(n8248), .ZN(n8054) );
  OR2_X1 U6945 ( .A1(n8442), .A2(n8054), .ZN(n5424) );
  NAND2_X2 U6946 ( .A1(n8237), .A2(n5424), .ZN(n8212) );
  INV_X1 U6947 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n9479) );
  NAND2_X1 U6948 ( .A1(n5425), .A2(n9479), .ZN(n5426) );
  AND2_X1 U6949 ( .A1(n5433), .A2(n5426), .ZN(n8221) );
  INV_X1 U6950 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n5429) );
  NAND2_X1 U6951 ( .A1(n5508), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n5428) );
  NAND2_X1 U6952 ( .A1(n5465), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n5427) );
  OAI211_X1 U6953 ( .C1(n5469), .C2(n5429), .A(n5428), .B(n5427), .ZN(n5430)
         );
  AOI21_X1 U6954 ( .B1(n8221), .B2(n4314), .A(n5430), .ZN(n8042) );
  NAND2_X1 U6955 ( .A1(n8439), .A2(n8042), .ZN(n7781) );
  INV_X1 U6956 ( .A(n5433), .ZN(n5431) );
  NAND2_X1 U6957 ( .A1(n5431), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5447) );
  INV_X1 U6958 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n5432) );
  NAND2_X1 U6959 ( .A1(n5433), .A2(n5432), .ZN(n5434) );
  NAND2_X1 U6960 ( .A1(n5447), .A2(n5434), .ZN(n8202) );
  INV_X1 U6961 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n5438) );
  NAND2_X1 U6962 ( .A1(n5435), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n5437) );
  NAND2_X1 U6963 ( .A1(n5465), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n5436) );
  OAI211_X1 U6964 ( .C1(n5469), .C2(n5438), .A(n5437), .B(n5436), .ZN(n5439)
         );
  INV_X1 U6965 ( .A(n5439), .ZN(n5440) );
  NAND2_X1 U6966 ( .A1(n8433), .A2(n8181), .ZN(n7785) );
  AND2_X1 U6967 ( .A1(n8213), .A2(n8194), .ZN(n5442) );
  INV_X1 U6968 ( .A(n8042), .ZN(n8230) );
  OR2_X1 U6969 ( .A1(n8439), .A2(n8230), .ZN(n8189) );
  OR2_X1 U6970 ( .A1(n8433), .A2(n8053), .ZN(n5443) );
  INV_X1 U6971 ( .A(n5447), .ZN(n5446) );
  NAND2_X1 U6972 ( .A1(n5446), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n5455) );
  INV_X1 U6973 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n9536) );
  NAND2_X1 U6974 ( .A1(n5447), .A2(n9536), .ZN(n5448) );
  NAND2_X1 U6975 ( .A1(n5455), .A2(n5448), .ZN(n8175) );
  INV_X1 U6976 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n5451) );
  NAND2_X1 U6977 ( .A1(n5465), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n5450) );
  NAND2_X1 U6978 ( .A1(n5508), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n5449) );
  OAI211_X1 U6979 ( .C1(n5469), .C2(n5451), .A(n5450), .B(n5449), .ZN(n5452)
         );
  INV_X1 U6980 ( .A(n5452), .ZN(n5453) );
  NAND2_X1 U6981 ( .A1(n8427), .A2(n8157), .ZN(n7788) );
  INV_X1 U6982 ( .A(n8157), .ZN(n8052) );
  INV_X1 U6983 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n7931) );
  NAND2_X1 U6984 ( .A1(n5455), .A2(n7931), .ZN(n5456) );
  NAND2_X1 U6985 ( .A1(n8164), .A2(n4314), .ZN(n5462) );
  INV_X1 U6986 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n5459) );
  NAND2_X1 U6987 ( .A1(n5508), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n5458) );
  NAND2_X1 U6988 ( .A1(n5465), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n5457) );
  OAI211_X1 U6989 ( .C1(n5469), .C2(n5459), .A(n5458), .B(n5457), .ZN(n5460)
         );
  INV_X1 U6990 ( .A(n5460), .ZN(n5461) );
  INV_X1 U6991 ( .A(n7794), .ZN(n5463) );
  INV_X1 U6992 ( .A(n5464), .ZN(n5517) );
  INV_X1 U6993 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n5468) );
  NAND2_X1 U6994 ( .A1(n5508), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n5467) );
  NAND2_X1 U6995 ( .A1(n5465), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n5466) );
  OAI211_X1 U6996 ( .C1(n5469), .C2(n5468), .A(n5467), .B(n5466), .ZN(n5470)
         );
  AOI21_X1 U6997 ( .B1(n5517), .B2(n4314), .A(n5470), .ZN(n8158) );
  INV_X1 U6998 ( .A(n7846), .ZN(n5472) );
  INV_X1 U6999 ( .A(n5474), .ZN(n5476) );
  NOR2_X1 U7000 ( .A1(n6502), .A2(n5819), .ZN(n5475) );
  NAND2_X1 U7001 ( .A1(n5476), .A2(n5475), .ZN(n5516) );
  XNOR2_X1 U7002 ( .A(n5218), .B(n5810), .ZN(n5477) );
  NAND2_X1 U7003 ( .A1(n5477), .A2(n8325), .ZN(n8379) );
  NAND2_X1 U7004 ( .A1(n5810), .A2(n9946), .ZN(n6239) );
  NAND2_X1 U7005 ( .A1(n8379), .A2(n6239), .ZN(n9952) );
  NAND2_X1 U7006 ( .A1(n9953), .A2(n9952), .ZN(n8365) );
  INV_X1 U7007 ( .A(n5887), .ZN(n5478) );
  NAND2_X1 U7008 ( .A1(n5478), .A2(n9963), .ZN(n7617) );
  NAND2_X1 U7009 ( .A1(n7650), .A2(n7654), .ZN(n5904) );
  INV_X1 U7010 ( .A(n5904), .ZN(n5480) );
  NAND2_X1 U7011 ( .A1(n5480), .A2(n5479), .ZN(n5906) );
  NAND2_X1 U7012 ( .A1(n5481), .A2(n6495), .ZN(n7644) );
  INV_X1 U7013 ( .A(n7644), .ZN(n5482) );
  AND2_X1 U7014 ( .A1(n7822), .A2(n5485), .ZN(n5484) );
  NAND2_X1 U7015 ( .A1(n6134), .A2(n5484), .ZN(n5489) );
  INV_X1 U7016 ( .A(n5485), .ZN(n5487) );
  INV_X1 U7017 ( .A(n7640), .ZN(n6455) );
  INV_X1 U7018 ( .A(n7826), .ZN(n6457) );
  AND2_X1 U7019 ( .A1(n6455), .A2(n6457), .ZN(n5486) );
  NAND2_X1 U7020 ( .A1(n5489), .A2(n5488), .ZN(n5490) );
  NAND2_X1 U7021 ( .A1(n6246), .A2(n6472), .ZN(n7679) );
  NAND2_X1 U7022 ( .A1(n5490), .A2(n7679), .ZN(n6619) );
  INV_X1 U7023 ( .A(n7705), .ZN(n5492) );
  INV_X1 U7024 ( .A(n7678), .ZN(n7825) );
  INV_X1 U7025 ( .A(n5493), .ZN(n7686) );
  OR2_X1 U7026 ( .A1(n7825), .A2(n7686), .ZN(n6730) );
  OR2_X1 U7027 ( .A1(n5495), .A2(n6730), .ZN(n5497) );
  AND2_X1 U7028 ( .A1(n7828), .A2(n7705), .ZN(n5494) );
  OR2_X1 U7029 ( .A1(n7686), .A2(n6816), .ZN(n6731) );
  AND2_X1 U7030 ( .A1(n5494), .A2(n6731), .ZN(n5496) );
  NAND2_X1 U7031 ( .A1(n6950), .A2(n7714), .ZN(n6860) );
  NAND2_X1 U7032 ( .A1(n7716), .A2(n7704), .ZN(n7713) );
  INV_X1 U7033 ( .A(n7713), .ZN(n5498) );
  NAND2_X1 U7034 ( .A1(n6860), .A2(n5498), .ZN(n5499) );
  NAND2_X1 U7035 ( .A1(n5499), .A2(n7715), .ZN(n7027) );
  NAND2_X1 U7036 ( .A1(n7027), .A2(n7834), .ZN(n5501) );
  NAND2_X1 U7037 ( .A1(n8505), .A2(n7055), .ZN(n5500) );
  INV_X1 U7038 ( .A(n5502), .ZN(n7741) );
  INV_X1 U7039 ( .A(n8318), .ZN(n7956) );
  NAND2_X1 U7040 ( .A1(n4820), .A2(n7749), .ZN(n8332) );
  INV_X1 U7041 ( .A(n8332), .ZN(n8339) );
  NOR2_X1 U7042 ( .A1(n8471), .A2(n8306), .ZN(n7758) );
  INV_X1 U7043 ( .A(n7758), .ZN(n5503) );
  AND2_X1 U7044 ( .A1(n8471), .A2(n8306), .ZN(n7756) );
  NAND2_X1 U7045 ( .A1(n5503), .A2(n7750), .ZN(n7838) );
  NAND2_X1 U7046 ( .A1(n8316), .A2(n8323), .ZN(n5504) );
  XNOR2_X1 U7047 ( .A(n8459), .B(n8056), .ZN(n7839) );
  NAND2_X1 U7048 ( .A1(n8459), .A2(n8308), .ZN(n7762) );
  INV_X1 U7049 ( .A(n8229), .ZN(n8006) );
  NAND2_X1 U7050 ( .A1(n8448), .A2(n8006), .ZN(n7775) );
  NAND2_X1 U7051 ( .A1(n8215), .A2(n8214), .ZN(n5505) );
  INV_X1 U7052 ( .A(n7780), .ZN(n8195) );
  NOR2_X1 U7053 ( .A1(n8194), .A2(n8195), .ZN(n5506) );
  XNOR2_X1 U7054 ( .A(n7625), .B(n7846), .ZN(n5515) );
  INV_X1 U7055 ( .A(n7818), .ZN(n7851) );
  NAND2_X1 U7056 ( .A1(n7851), .A2(n7852), .ZN(n7634) );
  NAND2_X1 U7057 ( .A1(n7850), .A2(n7634), .ZN(n8395) );
  INV_X1 U7058 ( .A(n7397), .ZN(n5507) );
  INV_X1 U7059 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n5511) );
  NAND2_X1 U7060 ( .A1(n5301), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n5510) );
  NAND2_X1 U7061 ( .A1(n5508), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n5509) );
  OAI211_X1 U7062 ( .C1(n5512), .C2(n5511), .A(n5510), .B(n5509), .ZN(n8050)
         );
  INV_X2 U7063 ( .A(n9953), .ZN(n8368) );
  AOI21_X1 U7064 ( .B1(n8416), .B2(n8163), .A(n8147), .ZN(n8417) );
  NAND2_X2 U7065 ( .A1(n8499), .A2(n8325), .ZN(n7635) );
  OR2_X1 U7066 ( .A1(n5516), .A2(n7635), .ZN(n8167) );
  AND2_X1 U7067 ( .A1(n9964), .A2(n7851), .ZN(n9942) );
  NAND2_X1 U7068 ( .A1(n9953), .A2(n9942), .ZN(n8406) );
  INV_X1 U7069 ( .A(n8356), .ZN(n9944) );
  AOI22_X1 U7070 ( .A1(n5517), .A2(n9944), .B1(P2_REG2_REG_29__SCAN_IN), .B2(
        n8368), .ZN(n5518) );
  OAI21_X1 U7071 ( .B1(n4467), .B2(n8406), .A(n5518), .ZN(n5519) );
  AOI21_X1 U7072 ( .B1(n8417), .B2(n8402), .A(n5519), .ZN(n5520) );
  OAI21_X1 U7073 ( .B1(n8418), .B2(n8368), .A(n5520), .ZN(n5521) );
  INV_X1 U7074 ( .A(n5521), .ZN(n5522) );
  OR2_X1 U7075 ( .A1(n5835), .A2(P2_U3152), .ZN(n5675) );
  NOR2_X1 U7076 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n5526) );
  NOR2_X1 U7077 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n5525) );
  NOR2_X1 U7078 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), .ZN(
        n5529) );
  INV_X1 U7079 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5530) );
  NAND4_X1 U7080 ( .A1(n5541), .A2(n5530), .A3(n5542), .A4(n5546), .ZN(n5531)
         );
  NOR2_X2 U7081 ( .A1(n5532), .A2(n5531), .ZN(n5533) );
  INV_X1 U7082 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5559) );
  NAND2_X1 U7083 ( .A1(n5537), .A2(n5554), .ZN(n5534) );
  NAND2_X1 U7084 ( .A1(n5534), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5535) );
  NAND2_X1 U7085 ( .A1(n4332), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5536) );
  XNOR2_X1 U7086 ( .A(n5537), .B(n5554), .ZN(n7064) );
  NAND2_X1 U7087 ( .A1(n5562), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5538) );
  MUX2_X1 U7088 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5538), .S(
        P1_IR_REG_23__SCAN_IN), .Z(n5539) );
  NAND2_X1 U7089 ( .A1(n5539), .A2(n4332), .ZN(n6089) );
  INV_X1 U7090 ( .A(n6089), .ZN(n6858) );
  NOR2_X1 U7091 ( .A1(n6090), .A2(n6858), .ZN(n6256) );
  NAND2_X1 U7092 ( .A1(n5945), .A2(n5541), .ZN(n6108) );
  INV_X1 U7093 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5544) );
  INV_X1 U7094 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5548) );
  OR2_X1 U7095 ( .A1(n5549), .A2(n5548), .ZN(n5550) );
  NAND2_X1 U7096 ( .A1(n5551), .A2(n5550), .ZN(n5842) );
  NAND2_X1 U7097 ( .A1(n5875), .A2(n5845), .ZN(n8805) );
  NAND2_X1 U7098 ( .A1(n8805), .A2(n6090), .ZN(n5552) );
  NAND2_X1 U7099 ( .A1(n5552), .A2(n6089), .ZN(n9695) );
  INV_X1 U7100 ( .A(n5558), .ZN(n5555) );
  INV_X1 U7101 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5556) );
  NAND2_X1 U7102 ( .A1(n9695), .A2(n6030), .ZN(n5564) );
  NAND2_X1 U7103 ( .A1(n5564), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  XNOR2_X1 U7104 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  AND2_X1 U7105 ( .A1(n5918), .A2(P1_U3084), .ZN(n9366) );
  INV_X1 U7106 ( .A(n9366), .ZN(n9376) );
  INV_X1 U7107 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n5919) );
  INV_X1 U7108 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n5566) );
  NAND2_X1 U7109 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5565) );
  XNOR2_X1 U7110 ( .A(n5566), .B(n5565), .ZN(n5963) );
  INV_X2 U7111 ( .A(n7272), .ZN(n9373) );
  OAI222_X1 U7112 ( .A1(n9376), .A2(n5919), .B1(n5963), .B2(P1_U3084), .C1(
        n9373), .C2(n5917), .ZN(P1_U3352) );
  OR2_X1 U7113 ( .A1(n5568), .A2(n5944), .ZN(n5570) );
  INV_X1 U7114 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5569) );
  NAND2_X1 U7115 ( .A1(n5570), .A2(n5569), .ZN(n5571) );
  OAI21_X1 U7116 ( .B1(n5570), .B2(n5569), .A(n5571), .ZN(n6029) );
  OAI222_X1 U7117 ( .A1(n9376), .A2(n6027), .B1(n9373), .B2(n6028), .C1(
        P1_U3084), .C2(n6029), .ZN(P1_U3351) );
  INV_X1 U7118 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6051) );
  NAND2_X1 U7119 ( .A1(n5571), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5573) );
  INV_X1 U7120 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5572) );
  XNOR2_X1 U7121 ( .A(n5573), .B(n5572), .ZN(n6160) );
  OAI222_X1 U7122 ( .A1(n9376), .A2(n6051), .B1(n9373), .B2(n6050), .C1(
        P1_U3084), .C2(n6160), .ZN(P1_U3350) );
  INV_X2 U7123 ( .A(n6279), .ZN(n8534) );
  AND2_X1 U7124 ( .A1(n5918), .A2(P2_U3152), .ZN(n8530) );
  OAI222_X1 U7125 ( .A1(n8534), .A2(n5574), .B1(n7939), .B2(n6028), .C1(
        P2_U3152), .C2(n5691), .ZN(P2_U3356) );
  OAI222_X1 U7126 ( .A1(n8534), .A2(n5575), .B1(n7939), .B2(n6050), .C1(
        P2_U3152), .C2(n5711), .ZN(P2_U3355) );
  OAI222_X1 U7127 ( .A1(n8534), .A2(n5576), .B1(n7939), .B2(n6066), .C1(
        P2_U3152), .C2(n5738), .ZN(P2_U3354) );
  INV_X1 U7128 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6068) );
  NAND2_X1 U7129 ( .A1(n5577), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5578) );
  MUX2_X1 U7130 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5578), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n5580) );
  NAND2_X1 U7131 ( .A1(n5580), .A2(n5579), .ZN(n6069) );
  OAI222_X1 U7132 ( .A1(n9376), .A2(n6068), .B1(n9373), .B2(n6066), .C1(
        P1_U3084), .C2(n6069), .ZN(P1_U3349) );
  OAI222_X1 U7133 ( .A1(n8534), .A2(n5582), .B1(n7939), .B2(n5917), .C1(n5581), 
        .C2(P2_U3152), .ZN(P2_U3357) );
  INV_X1 U7134 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6311) );
  NAND2_X1 U7135 ( .A1(n5579), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5583) );
  XNOR2_X1 U7136 ( .A(n5583), .B(P1_IR_REG_5__SCAN_IN), .ZN(n5972) );
  OAI222_X1 U7137 ( .A1(n9376), .A2(n6311), .B1(n9373), .B2(n6310), .C1(
        P1_U3084), .C2(n4475), .ZN(P1_U3348) );
  OAI222_X1 U7138 ( .A1(n8534), .A2(n5584), .B1(n7939), .B2(n6310), .C1(
        P2_U3152), .C2(n5728), .ZN(P2_U3353) );
  OAI222_X1 U7139 ( .A1(n8534), .A2(n5585), .B1(n7939), .B2(n6326), .C1(
        P2_U3152), .C2(n5748), .ZN(P2_U3352) );
  INV_X1 U7140 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6327) );
  OR2_X1 U7141 ( .A1(n5586), .A2(n5944), .ZN(n5587) );
  INV_X1 U7142 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5589) );
  XNOR2_X1 U7143 ( .A(n5587), .B(n5589), .ZN(n9737) );
  OAI222_X1 U7144 ( .A1(n9376), .A2(n6327), .B1(n9373), .B2(n6326), .C1(
        P1_U3084), .C2(n9737), .ZN(P1_U3347) );
  INV_X1 U7145 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n5588) );
  INV_X1 U7146 ( .A(n6351), .ZN(n5591) );
  INV_X1 U7147 ( .A(n5761), .ZN(n5773) );
  OAI222_X1 U7148 ( .A1(n8534), .A2(n5588), .B1(n7939), .B2(n5591), .C1(
        P2_U3152), .C2(n5773), .ZN(P2_U3351) );
  INV_X1 U7149 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n5592) );
  NAND2_X1 U7150 ( .A1(n5586), .A2(n5589), .ZN(n5602) );
  NAND2_X1 U7151 ( .A1(n5602), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5590) );
  XNOR2_X1 U7152 ( .A(n5590), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6349) );
  INV_X1 U7153 ( .A(n6349), .ZN(n5978) );
  OAI222_X1 U7154 ( .A1(n9376), .A2(n5592), .B1(n9373), .B2(n5591), .C1(
        P1_U3084), .C2(n5978), .ZN(P1_U3346) );
  AND2_X1 U7155 ( .A1(n6089), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5593) );
  NAND2_X1 U7156 ( .A1(n6090), .A2(n5593), .ZN(n9850) );
  INV_X1 U7157 ( .A(n9850), .ZN(n9846) );
  INV_X1 U7158 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n5600) );
  INV_X1 U7159 ( .A(n7064), .ZN(n5595) );
  NAND2_X1 U7160 ( .A1(n7010), .A2(P1_B_REG_SCAN_IN), .ZN(n5594) );
  OAI22_X1 U7161 ( .A1(n5595), .A2(n5594), .B1(P1_B_REG_SCAN_IN), .B2(n7010), 
        .ZN(n5596) );
  OR2_X1 U7162 ( .A1(n5596), .A2(n7162), .ZN(n9845) );
  OR2_X1 U7163 ( .A1(n9845), .A2(P1_D_REG_1__SCAN_IN), .ZN(n5598) );
  NAND2_X1 U7164 ( .A1(n7162), .A2(n7064), .ZN(n5597) );
  NAND2_X1 U7165 ( .A1(n5598), .A2(n5597), .ZN(n6993) );
  INV_X1 U7166 ( .A(n6993), .ZN(n6005) );
  NAND2_X1 U7167 ( .A1(n6005), .A2(n9846), .ZN(n5599) );
  OAI21_X1 U7168 ( .B1(n9846), .B2(n5600), .A(n5599), .ZN(P1_U3441) );
  INV_X1 U7169 ( .A(n6579), .ZN(n5608) );
  INV_X1 U7170 ( .A(n8073), .ZN(n5775) );
  OAI222_X1 U7171 ( .A1(n8534), .A2(n5601), .B1(n7939), .B2(n5608), .C1(
        P2_U3152), .C2(n5775), .ZN(P2_U3350) );
  NOR2_X1 U7172 ( .A1(n5603), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n5616) );
  INV_X1 U7173 ( .A(n5616), .ZN(n5607) );
  NAND2_X1 U7174 ( .A1(n5603), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5605) );
  MUX2_X1 U7175 ( .A(n5605), .B(P1_IR_REG_31__SCAN_IN), .S(n5604), .Z(n5606)
         );
  INV_X1 U7176 ( .A(n6580), .ZN(n9752) );
  OAI222_X1 U7177 ( .A1(n9376), .A2(n5609), .B1(n9373), .B2(n5608), .C1(
        P1_U3084), .C2(n9752), .ZN(P1_U3345) );
  INV_X1 U7178 ( .A(n6748), .ZN(n5612) );
  OR2_X1 U7179 ( .A1(n5616), .A2(n5944), .ZN(n5610) );
  XNOR2_X1 U7180 ( .A(n5610), .B(P1_IR_REG_9__SCAN_IN), .ZN(n9757) );
  AOI22_X1 U7181 ( .A1(n9757), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n9366), .ZN(n5611) );
  OAI21_X1 U7182 ( .B1(n5612), .B2(n9373), .A(n5611), .ZN(P1_U3344) );
  INV_X1 U7183 ( .A(n8085), .ZN(n5777) );
  OAI222_X1 U7184 ( .A1(n8534), .A2(n5613), .B1(n7939), .B2(n5612), .C1(n5777), 
        .C2(P2_U3152), .ZN(P2_U3349) );
  INV_X1 U7185 ( .A(n6829), .ZN(n5618) );
  INV_X1 U7186 ( .A(n8100), .ZN(n5779) );
  OAI222_X1 U7187 ( .A1(n8534), .A2(n5614), .B1(n7939), .B2(n5618), .C1(n5779), 
        .C2(P2_U3152), .ZN(P2_U3348) );
  INV_X1 U7188 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n5615) );
  NAND2_X1 U7189 ( .A1(n5616), .A2(n5615), .ZN(n5620) );
  NAND2_X1 U7190 ( .A1(n5620), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5617) );
  XNOR2_X1 U7191 ( .A(n5617), .B(P1_IR_REG_10__SCAN_IN), .ZN(n6830) );
  INV_X1 U7192 ( .A(n6830), .ZN(n9782) );
  OAI222_X1 U7193 ( .A1(n9376), .A2(n5619), .B1(n9782), .B2(P1_U3084), .C1(
        n9373), .C2(n5618), .ZN(P1_U3343) );
  INV_X1 U7194 ( .A(n7069), .ZN(n5623) );
  OAI21_X1 U7195 ( .B1(n5620), .B2(P1_IR_REG_10__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5621) );
  XNOR2_X1 U7196 ( .A(n5621), .B(P1_IR_REG_11__SCAN_IN), .ZN(n7070) );
  INV_X1 U7197 ( .A(n7070), .ZN(n5996) );
  INV_X1 U7198 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n5622) );
  OAI222_X1 U7199 ( .A1(n9373), .A2(n5623), .B1(n5996), .B2(P1_U3084), .C1(
        n5622), .C2(n9376), .ZN(P1_U3342) );
  INV_X1 U7200 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n5624) );
  INV_X1 U7201 ( .A(n5781), .ZN(n5802) );
  OAI222_X1 U7202 ( .A1(n8534), .A2(n5624), .B1(n7939), .B2(n5623), .C1(n5802), 
        .C2(P2_U3152), .ZN(P2_U3347) );
  NAND2_X1 U7203 ( .A1(n6361), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n6591) );
  INV_X1 U7204 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n6590) );
  INV_X1 U7205 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n6843) );
  INV_X1 U7206 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n6844) );
  NAND2_X1 U7207 ( .A1(n7079), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n7088) );
  INV_X1 U7208 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n7087) );
  INV_X1 U7209 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n7177) );
  INV_X1 U7210 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n7322) );
  INV_X1 U7211 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n8643) );
  AND2_X1 U7212 ( .A1(n7325), .A2(n8643), .ZN(n5628) );
  NOR2_X1 U7213 ( .A1(n7354), .A2(n5628), .ZN(n9200) );
  NAND2_X1 U7214 ( .A1(n7554), .A2(n9200), .ZN(n5636) );
  INV_X1 U7215 ( .A(n7555), .ZN(n7600) );
  INV_X1 U7216 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n5629) );
  OR2_X1 U7217 ( .A1(n7600), .A2(n5629), .ZN(n5635) );
  INV_X1 U7218 ( .A(n6044), .ZN(n6081) );
  INV_X1 U7219 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n8960) );
  OR2_X1 U7220 ( .A1(n6044), .A2(n8960), .ZN(n5634) );
  INV_X1 U7221 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n5632) );
  OR2_X1 U7222 ( .A1(n7598), .A2(n5632), .ZN(n5633) );
  INV_X1 U7223 ( .A(P1_U4006), .ZN(n5638) );
  NAND2_X1 U7224 ( .A1(n5638), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n5637) );
  OAI21_X1 U7225 ( .B1(n9217), .B2(n5638), .A(n5637), .ZN(P1_U3573) );
  INV_X1 U7226 ( .A(n7073), .ZN(n5645) );
  NOR2_X1 U7227 ( .A1(n5639), .A2(n5944), .ZN(n5640) );
  MUX2_X1 U7228 ( .A(n5944), .B(n5640), .S(P1_IR_REG_12__SCAN_IN), .Z(n5643)
         );
  INV_X1 U7229 ( .A(n5641), .ZN(n5642) );
  OR2_X1 U7230 ( .A1(n5643), .A2(n5641), .ZN(n7074) );
  OAI222_X1 U7231 ( .A1(n9376), .A2(n5644), .B1(n9373), .B2(n5645), .C1(
        P1_U3084), .C2(n7074), .ZN(P1_U3341) );
  INV_X1 U7232 ( .A(n6120), .ZN(n6113) );
  OAI222_X1 U7233 ( .A1(n8534), .A2(n5646), .B1(n7939), .B2(n5645), .C1(
        P2_U3152), .C2(n6113), .ZN(P2_U3346) );
  AND2_X1 U7234 ( .A1(n5832), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7856) );
  INV_X1 U7235 ( .A(n7856), .ZN(n7861) );
  NAND2_X1 U7236 ( .A1(n9956), .A2(n7861), .ZN(n5648) );
  NAND2_X1 U7237 ( .A1(n5648), .A2(n5647), .ZN(n5651) );
  INV_X1 U7238 ( .A(n5822), .ZN(n5649) );
  OR2_X1 U7239 ( .A1(n9956), .A2(n5649), .ZN(n5650) );
  AND2_X1 U7240 ( .A1(n5651), .A2(n5650), .ZN(n9604) );
  NOR2_X1 U7241 ( .A1(n9935), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U7242 ( .A(n7168), .ZN(n5655) );
  NAND2_X1 U7243 ( .A1(n5642), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5652) );
  XNOR2_X1 U7244 ( .A(n5652), .B(P1_IR_REG_13__SCAN_IN), .ZN(n7169) );
  AOI22_X1 U7245 ( .A1(n7169), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n9366), .ZN(n5653) );
  OAI21_X1 U7246 ( .B1(n5655), .B2(n9373), .A(n5653), .ZN(P1_U3340) );
  AOI22_X1 U7247 ( .A1(n6291), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_13__SCAN_IN), .B2(n6279), .ZN(n5654) );
  OAI21_X1 U7248 ( .B1(n5655), .B2(n7939), .A(n5654), .ZN(P2_U3345) );
  INV_X1 U7249 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n5658) );
  INV_X1 U7250 ( .A(n7630), .ZN(n5656) );
  NAND2_X1 U7251 ( .A1(P2_U3966), .A2(n5656), .ZN(n5657) );
  OAI21_X1 U7252 ( .B1(P2_U3966), .B2(n5658), .A(n5657), .ZN(P2_U3583) );
  NAND2_X1 U7253 ( .A1(P2_U3966), .A2(n5887), .ZN(n5659) );
  OAI21_X1 U7254 ( .B1(P2_U3966), .B2(n4509), .A(n5659), .ZN(P2_U3552) );
  INV_X1 U7255 ( .A(n7209), .ZN(n5673) );
  NAND2_X1 U7256 ( .A1(n5660), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5662) );
  OR2_X1 U7257 ( .A1(n5662), .A2(n5661), .ZN(n5663) );
  NAND2_X1 U7258 ( .A1(n5662), .A2(n5661), .ZN(n5790) );
  AND2_X1 U7259 ( .A1(n5663), .A2(n5790), .ZN(n7210) );
  INV_X1 U7260 ( .A(n7210), .ZN(n6962) );
  INV_X1 U7261 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n5664) );
  OAI222_X1 U7262 ( .A1(n9373), .A2(n5673), .B1(n6962), .B2(P1_U3084), .C1(
        n5664), .C2(n9376), .ZN(P1_U3339) );
  INV_X1 U7263 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5672) );
  NAND2_X1 U7264 ( .A1(n4333), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5670) );
  INV_X1 U7265 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n5854) );
  OR2_X1 U7266 ( .A1(n4316), .A2(n5854), .ZN(n5669) );
  INV_X1 U7267 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n5665) );
  INV_X1 U7268 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n5666) );
  NAND2_X1 U7269 ( .A1(n6298), .A2(P1_U4006), .ZN(n5671) );
  OAI21_X1 U7270 ( .B1(P1_U4006), .B2(n5672), .A(n5671), .ZN(P1_U3555) );
  INV_X1 U7271 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n5674) );
  INV_X1 U7272 ( .A(n6718), .ZN(n6715) );
  OAI222_X1 U7273 ( .A1(n8534), .A2(n5674), .B1(n7939), .B2(n5673), .C1(n6715), 
        .C2(P2_U3152), .ZN(P2_U3344) );
  OAI211_X1 U7274 ( .C1(n9956), .C2(n5822), .A(n7861), .B(n5675), .ZN(n5684)
         );
  NAND2_X1 U7275 ( .A1(n5684), .A2(n5682), .ZN(n5676) );
  NAND2_X1 U7276 ( .A1(n8055), .A2(n5676), .ZN(n5694) );
  AND2_X1 U7277 ( .A1(n5694), .A2(n7397), .ZN(n9619) );
  INV_X1 U7278 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n9534) );
  NOR2_X1 U7279 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9534), .ZN(n5688) );
  INV_X1 U7280 ( .A(n5691), .ZN(n9618) );
  INV_X1 U7281 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n9938) );
  INV_X1 U7282 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10020) );
  OR2_X1 U7283 ( .A1(n9606), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5678) );
  NAND2_X1 U7284 ( .A1(n9606), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5677) );
  NAND2_X1 U7285 ( .A1(n5678), .A2(n5677), .ZN(n9598) );
  NOR3_X1 U7286 ( .A1(n9938), .A2(n10020), .A3(n9598), .ZN(n9596) );
  AND2_X1 U7287 ( .A1(n9606), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5679) );
  NOR2_X1 U7288 ( .A1(n9596), .A2(n5679), .ZN(n9616) );
  INV_X1 U7289 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n5680) );
  MUX2_X1 U7290 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n5680), .S(n5691), .Z(n9615)
         );
  NOR2_X1 U7291 ( .A1(n9616), .A2(n9615), .ZN(n9614) );
  AOI21_X1 U7292 ( .B1(n9618), .B2(P2_REG1_REG_2__SCAN_IN), .A(n9614), .ZN(
        n5686) );
  INV_X1 U7293 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n5681) );
  MUX2_X1 U7294 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n5681), .S(n5711), .Z(n5685)
         );
  NOR2_X1 U7295 ( .A1(n5686), .A2(n5685), .ZN(n5700) );
  AND2_X1 U7296 ( .A1(n5682), .A2(n4994), .ZN(n5683) );
  INV_X1 U7297 ( .A(n9930), .ZN(n9613) );
  AOI211_X1 U7298 ( .C1(n5686), .C2(n5685), .A(n5700), .B(n9613), .ZN(n5687)
         );
  AOI211_X1 U7299 ( .C1(P2_ADDR_REG_3__SCAN_IN), .C2(n9935), .A(n5688), .B(
        n5687), .ZN(n5698) );
  INV_X1 U7300 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n5910) );
  MUX2_X1 U7301 ( .A(n5910), .B(P2_REG2_REG_2__SCAN_IN), .S(n5691), .Z(n9621)
         );
  NAND2_X1 U7302 ( .A1(n9606), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5690) );
  INV_X1 U7303 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n5689) );
  NAND3_X1 U7304 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .A3(n9609), .ZN(n9608) );
  INV_X1 U7305 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n5692) );
  MUX2_X1 U7306 ( .A(n5692), .B(P2_REG2_REG_3__SCAN_IN), .S(n5711), .Z(n5695)
         );
  NOR2_X1 U7307 ( .A1(n7397), .A2(n4994), .ZN(n5693) );
  NAND2_X1 U7308 ( .A1(n5694), .A2(n5693), .ZN(n9933) );
  OAI211_X1 U7309 ( .C1(n5696), .C2(n5695), .A(n9929), .B(n5710), .ZN(n5697)
         );
  OAI211_X1 U7310 ( .C1(n9932), .C2(n5711), .A(n5698), .B(n5697), .ZN(P2_U3248) );
  NOR2_X1 U7311 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5699), .ZN(n6553) );
  INV_X1 U7312 ( .A(n5738), .ZN(n5702) );
  XOR2_X1 U7313 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n5738), .Z(n5730) );
  INV_X1 U7314 ( .A(n5711), .ZN(n5701) );
  AOI21_X1 U7315 ( .B1(n5701), .B2(P2_REG1_REG_3__SCAN_IN), .A(n5700), .ZN(
        n5731) );
  NOR2_X1 U7316 ( .A1(n5730), .A2(n5731), .ZN(n5729) );
  AOI21_X1 U7317 ( .B1(P2_REG1_REG_4__SCAN_IN), .B2(n5702), .A(n5729), .ZN(
        n5720) );
  NAND2_X1 U7318 ( .A1(n5708), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5703) );
  OAI21_X1 U7319 ( .B1(n5708), .B2(P2_REG1_REG_5__SCAN_IN), .A(n5703), .ZN(
        n5719) );
  NOR2_X1 U7320 ( .A1(n5720), .A2(n5719), .ZN(n5718) );
  AOI21_X1 U7321 ( .B1(P2_REG1_REG_5__SCAN_IN), .B2(n5708), .A(n5718), .ZN(
        n5706) );
  INV_X1 U7322 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n5704) );
  MUX2_X1 U7323 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n5704), .S(n5748), .Z(n5705)
         );
  NOR2_X1 U7324 ( .A1(n5706), .A2(n5705), .ZN(n5739) );
  AOI211_X1 U7325 ( .C1(n5706), .C2(n5705), .A(n5739), .B(n9613), .ZN(n5707)
         );
  AOI211_X1 U7326 ( .C1(P2_ADDR_REG_6__SCAN_IN), .C2(n9935), .A(n6553), .B(
        n5707), .ZN(n5717) );
  NAND2_X1 U7327 ( .A1(n5708), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5713) );
  INV_X1 U7328 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n5709) );
  MUX2_X1 U7329 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n5709), .S(n5708), .Z(n5725)
         );
  INV_X1 U7330 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n5712) );
  MUX2_X1 U7331 ( .A(n5712), .B(P2_REG2_REG_4__SCAN_IN), .S(n5738), .Z(n5735)
         );
  OAI21_X1 U7332 ( .B1(n5711), .B2(n5692), .A(n5710), .ZN(n5734) );
  NAND2_X1 U7333 ( .A1(n5735), .A2(n5734), .ZN(n5733) );
  OAI21_X1 U7334 ( .B1(n5712), .B2(n5738), .A(n5733), .ZN(n5724) );
  NAND2_X1 U7335 ( .A1(n5725), .A2(n5724), .ZN(n5723) );
  NAND2_X1 U7336 ( .A1(n5713), .A2(n5723), .ZN(n5715) );
  INV_X1 U7337 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6462) );
  MUX2_X1 U7338 ( .A(n6462), .B(P2_REG2_REG_6__SCAN_IN), .S(n5748), .Z(n5714)
         );
  NAND2_X1 U7339 ( .A1(n5715), .A2(n5714), .ZN(n5747) );
  OAI211_X1 U7340 ( .C1(n5715), .C2(n5714), .A(n9929), .B(n5747), .ZN(n5716)
         );
  OAI211_X1 U7341 ( .C1(n9932), .C2(n5748), .A(n5717), .B(n5716), .ZN(P2_U3251) );
  NOR2_X1 U7342 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5257), .ZN(n5722) );
  AOI211_X1 U7343 ( .C1(n5720), .C2(n5719), .A(n5718), .B(n9613), .ZN(n5721)
         );
  AOI211_X1 U7344 ( .C1(P2_ADDR_REG_5__SCAN_IN), .C2(n9935), .A(n5722), .B(
        n5721), .ZN(n5727) );
  OAI211_X1 U7345 ( .C1(n5725), .C2(n5724), .A(n9929), .B(n5723), .ZN(n5726)
         );
  OAI211_X1 U7346 ( .C1(n9932), .C2(n5728), .A(n5727), .B(n5726), .ZN(P2_U3250) );
  INV_X1 U7347 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n9572) );
  NOR2_X1 U7348 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9572), .ZN(n6205) );
  AOI211_X1 U7349 ( .C1(n5731), .C2(n5730), .A(n5729), .B(n9613), .ZN(n5732)
         );
  AOI211_X1 U7350 ( .C1(P2_ADDR_REG_4__SCAN_IN), .C2(n9935), .A(n6205), .B(
        n5732), .ZN(n5737) );
  OAI211_X1 U7351 ( .C1(n5735), .C2(n5734), .A(n9929), .B(n5733), .ZN(n5736)
         );
  OAI211_X1 U7352 ( .C1(n9932), .C2(n5738), .A(n5737), .B(n5736), .ZN(P2_U3249) );
  NOR2_X1 U7353 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5273), .ZN(n6607) );
  INV_X1 U7354 ( .A(n5748), .ZN(n5740) );
  AOI21_X1 U7355 ( .B1(P2_REG1_REG_6__SCAN_IN), .B2(n5740), .A(n5739), .ZN(
        n5745) );
  OR2_X1 U7356 ( .A1(n5761), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5742) );
  NAND2_X1 U7357 ( .A1(n5761), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5741) );
  NAND2_X1 U7358 ( .A1(n5742), .A2(n5741), .ZN(n5744) );
  INV_X1 U7359 ( .A(n5772), .ZN(n5743) );
  AOI211_X1 U7360 ( .C1(n5745), .C2(n5744), .A(n5743), .B(n9613), .ZN(n5746)
         );
  AOI211_X1 U7361 ( .C1(P2_ADDR_REG_7__SCAN_IN), .C2(n9935), .A(n6607), .B(
        n5746), .ZN(n5752) );
  INV_X1 U7362 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n5749) );
  MUX2_X1 U7363 ( .A(n5749), .B(P2_REG2_REG_7__SCAN_IN), .S(n5761), .Z(n5762)
         );
  XNOR2_X1 U7364 ( .A(n5764), .B(n5762), .ZN(n5750) );
  NAND2_X1 U7365 ( .A1(n9929), .A2(n5750), .ZN(n5751) );
  OAI211_X1 U7366 ( .C1(n9932), .C2(n5773), .A(n5752), .B(n5751), .ZN(P2_U3252) );
  NAND2_X1 U7367 ( .A1(n7555), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n5757) );
  INV_X1 U7368 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n5753) );
  OR2_X1 U7369 ( .A1(n6044), .A2(n5753), .ZN(n5756) );
  INV_X1 U7370 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n5754) );
  OR2_X1 U7371 ( .A1(n7598), .A2(n5754), .ZN(n5755) );
  AND3_X1 U7372 ( .A1(n5757), .A2(n5756), .A3(n5755), .ZN(n8772) );
  INV_X1 U7373 ( .A(n8772), .ZN(n8994) );
  NAND2_X1 U7374 ( .A1(n8994), .A2(P1_U4006), .ZN(n5758) );
  OAI21_X1 U7375 ( .B1(P1_U4006), .B2(n8535), .A(n5758), .ZN(P1_U3586) );
  INV_X1 U7376 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n5768) );
  NAND2_X1 U7377 ( .A1(n8085), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5767) );
  INV_X1 U7378 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n5759) );
  MUX2_X1 U7379 ( .A(n5759), .B(P2_REG2_REG_9__SCAN_IN), .S(n8085), .Z(n5760)
         );
  INV_X1 U7380 ( .A(n5760), .ZN(n8083) );
  INV_X1 U7381 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n5766) );
  NAND2_X1 U7382 ( .A1(n5761), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5765) );
  INV_X1 U7383 ( .A(n5762), .ZN(n5763) );
  MUX2_X1 U7384 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n5766), .S(n8073), .Z(n8070)
         );
  OAI21_X1 U7385 ( .B1(n5766), .B2(n5775), .A(n8069), .ZN(n8082) );
  NAND2_X1 U7386 ( .A1(n8083), .A2(n8082), .ZN(n8081) );
  MUX2_X1 U7387 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n5768), .S(n8100), .Z(n8098)
         );
  INV_X1 U7388 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n5769) );
  MUX2_X1 U7389 ( .A(n5769), .B(P2_REG2_REG_11__SCAN_IN), .S(n5781), .Z(n5770)
         );
  AOI21_X1 U7390 ( .B1(n5771), .B2(n5770), .A(n5801), .ZN(n5789) );
  INV_X1 U7391 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n5780) );
  INV_X1 U7392 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n5778) );
  INV_X1 U7393 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n5776) );
  INV_X1 U7394 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n5774) );
  OAI21_X1 U7395 ( .B1(n5774), .B2(n5773), .A(n5772), .ZN(n8075) );
  MUX2_X1 U7396 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n5776), .S(n8073), .Z(n8076)
         );
  NAND2_X1 U7397 ( .A1(n8075), .A2(n8076), .ZN(n8074) );
  OAI21_X1 U7398 ( .B1(n5776), .B2(n5775), .A(n8074), .ZN(n8088) );
  MUX2_X1 U7399 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n5778), .S(n8085), .Z(n8087)
         );
  NAND2_X1 U7400 ( .A1(n8088), .A2(n8087), .ZN(n8086) );
  OAI21_X1 U7401 ( .B1(n5778), .B2(n5777), .A(n8086), .ZN(n8095) );
  MUX2_X1 U7402 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n5780), .S(n8100), .Z(n8094)
         );
  NAND2_X1 U7403 ( .A1(n8095), .A2(n8094), .ZN(n8093) );
  OAI21_X1 U7404 ( .B1(n5780), .B2(n5779), .A(n8093), .ZN(n5783) );
  INV_X1 U7405 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n6961) );
  MUX2_X1 U7406 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n6961), .S(n5781), .Z(n5782)
         );
  NAND2_X1 U7407 ( .A1(n5783), .A2(n5782), .ZN(n5796) );
  OAI211_X1 U7408 ( .C1(n5783), .C2(n5782), .A(n5796), .B(n9930), .ZN(n5786)
         );
  NOR2_X1 U7409 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5311), .ZN(n5784) );
  AOI21_X1 U7410 ( .B1(n9935), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n5784), .ZN(
        n5785) );
  OAI211_X1 U7411 ( .C1(n9932), .C2(n5802), .A(n5786), .B(n5785), .ZN(n5787)
         );
  INV_X1 U7412 ( .A(n5787), .ZN(n5788) );
  OAI21_X1 U7413 ( .B1(n5789), .B2(n9933), .A(n5788), .ZN(P2_U3256) );
  INV_X1 U7414 ( .A(n7303), .ZN(n5794) );
  NAND2_X1 U7415 ( .A1(n5790), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5792) );
  XNOR2_X1 U7416 ( .A(n5792), .B(n5791), .ZN(n7150) );
  OAI222_X1 U7417 ( .A1(n9376), .A2(n5793), .B1(n9373), .B2(n5794), .C1(
        P1_U3084), .C2(n7150), .ZN(P1_U3338) );
  INV_X1 U7418 ( .A(n6876), .ZN(n6870) );
  OAI222_X1 U7419 ( .A1(n8534), .A2(n5795), .B1(n7939), .B2(n5794), .C1(
        P2_U3152), .C2(n6870), .ZN(P2_U3343) );
  INV_X1 U7420 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n10031) );
  MUX2_X1 U7421 ( .A(n10031), .B(P2_REG1_REG_12__SCAN_IN), .S(n6120), .Z(n5798) );
  OAI21_X1 U7422 ( .B1(n6961), .B2(n5802), .A(n5796), .ZN(n5797) );
  NOR2_X1 U7423 ( .A1(n5797), .A2(n5798), .ZN(n6118) );
  AOI21_X1 U7424 ( .B1(n5798), .B2(n5797), .A(n6118), .ZN(n5807) );
  NAND2_X1 U7425 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3152), .ZN(n6922) );
  INV_X1 U7426 ( .A(n6922), .ZN(n5800) );
  NOR2_X1 U7427 ( .A1(n9932), .A2(n6113), .ZN(n5799) );
  AOI211_X1 U7428 ( .C1(P2_ADDR_REG_12__SCAN_IN), .C2(n9935), .A(n5800), .B(
        n5799), .ZN(n5806) );
  AOI21_X1 U7429 ( .B1(n5802), .B2(n5769), .A(n5801), .ZN(n5804) );
  INV_X1 U7430 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n6114) );
  MUX2_X1 U7431 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n6114), .S(n6120), .Z(n5803)
         );
  NAND2_X1 U7432 ( .A1(n5803), .A2(n5804), .ZN(n6112) );
  OAI211_X1 U7433 ( .C1(n5804), .C2(n5803), .A(n9929), .B(n6112), .ZN(n5805)
         );
  OAI211_X1 U7434 ( .C1(n5807), .C2(n9613), .A(n5806), .B(n5805), .ZN(P2_U3257) );
  INV_X1 U7435 ( .A(n5816), .ZN(n5814) );
  INV_X1 U7436 ( .A(n9964), .ZN(n5809) );
  NAND3_X1 U7437 ( .A1(n5809), .A2(n6543), .A3(n7850), .ZN(n5812) );
  INV_X1 U7438 ( .A(n5810), .ZN(n5811) );
  INV_X1 U7439 ( .A(n5815), .ZN(n5813) );
  NOR2_X1 U7440 ( .A1(n7926), .A2(n9963), .ZN(n5817) );
  AOI21_X1 U7441 ( .B1(n5893), .B2(n7635), .A(n5817), .ZN(n6211) );
  XNOR2_X1 U7442 ( .A(n7926), .B(n9975), .ZN(n6186) );
  NAND2_X1 U7443 ( .A1(n5818), .A2(n7635), .ZN(n6185) );
  XNOR2_X1 U7444 ( .A(n6186), .B(n6185), .ZN(n6187) );
  XNOR2_X1 U7445 ( .A(n6188), .B(n6187), .ZN(n5840) );
  INV_X1 U7446 ( .A(n5819), .ZN(n5820) );
  AND3_X1 U7447 ( .A1(n5821), .A2(n5820), .A3(n6502), .ZN(n5827) );
  INV_X1 U7448 ( .A(n9956), .ZN(n7859) );
  NAND2_X1 U7449 ( .A1(n5827), .A2(n7859), .ZN(n5826) );
  INV_X1 U7450 ( .A(n5826), .ZN(n5824) );
  NOR2_X1 U7451 ( .A1(n8498), .A2(n5822), .ZN(n5823) );
  NOR2_X1 U7452 ( .A1(n5826), .A2(n5825), .ZN(n8043) );
  NAND2_X1 U7453 ( .A1(n8043), .A2(n8390), .ZN(n8030) );
  INV_X1 U7454 ( .A(n8030), .ZN(n6609) );
  NAND2_X1 U7455 ( .A1(n8043), .A2(n8392), .ZN(n8029) );
  INV_X1 U7456 ( .A(n8029), .ZN(n6608) );
  AOI22_X1 U7457 ( .A1(n6609), .A2(n5808), .B1(n6608), .B2(n8068), .ZN(n5839)
         );
  INV_X1 U7458 ( .A(n5827), .ZN(n5829) );
  NAND2_X1 U7459 ( .A1(n5829), .A2(n5828), .ZN(n5837) );
  INV_X1 U7460 ( .A(n5837), .ZN(n5830) );
  NOR3_X1 U7461 ( .A1(n5830), .A2(n10008), .A3(n9956), .ZN(n5831) );
  NOR2_X1 U7462 ( .A1(n5833), .A2(n5832), .ZN(n5834) );
  AND2_X1 U7463 ( .A1(n5835), .A2(n5834), .ZN(n5836) );
  NAND2_X1 U7464 ( .A1(n5837), .A2(n5836), .ZN(n6202) );
  OR2_X1 U7465 ( .A1(n6202), .A2(P2_U3152), .ZN(n7621) );
  AOI22_X1 U7466 ( .A1(n8047), .A2(n5914), .B1(P2_REG3_REG_2__SCAN_IN), .B2(
        n7621), .ZN(n5838) );
  OAI211_X1 U7467 ( .C1(n5840), .C2(n8036), .A(n5839), .B(n5838), .ZN(P2_U3239) );
  INV_X1 U7468 ( .A(SI_0_), .ZN(n9539) );
  NOR2_X1 U7469 ( .A1(n5918), .A2(n9539), .ZN(n5841) );
  XNOR2_X1 U7470 ( .A(n5841), .B(n4509), .ZN(n9377) );
  MUX2_X1 U7471 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9377), .S(n6030), .Z(n6302) );
  INV_X1 U7472 ( .A(n5842), .ZN(n5845) );
  XNOR2_X1 U7473 ( .A(n5843), .B(P1_IR_REG_20__SCAN_IN), .ZN(n6996) );
  NOR2_X2 U7474 ( .A1(n5876), .A2(n5846), .ZN(n6036) );
  AOI22_X1 U7475 ( .A1(n6302), .A2(n6036), .B1(n5846), .B2(
        P1_IR_REG_0__SCAN_IN), .ZN(n5847) );
  INV_X1 U7476 ( .A(n5847), .ZN(n5853) );
  NAND2_X1 U7477 ( .A1(n4344), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5849) );
  XNOR2_X2 U7478 ( .A(n5849), .B(n5848), .ZN(n9154) );
  NAND2_X1 U7479 ( .A1(n5883), .A2(n5859), .ZN(n5850) );
  AND2_X4 U7480 ( .A1(n5876), .A2(n6090), .ZN(n7579) );
  NAND2_X1 U7481 ( .A1(n6298), .A2(n6036), .ZN(n5857) );
  NOR2_X1 U7482 ( .A1(n6090), .A2(n5854), .ZN(n5855) );
  AOI21_X1 U7483 ( .B1(n6302), .B2(n7579), .A(n5855), .ZN(n5856) );
  NAND2_X1 U7484 ( .A1(n5857), .A2(n5856), .ZN(n5922) );
  NAND2_X1 U7485 ( .A1(n5858), .A2(n5922), .ZN(n5926) );
  OAI21_X1 U7486 ( .B1(n5858), .B2(n5922), .A(n5926), .ZN(n6253) );
  NAND2_X1 U7487 ( .A1(n5859), .A2(n5842), .ZN(n9344) );
  OR2_X1 U7488 ( .A1(n9344), .A2(n5844), .ZN(n6016) );
  OR2_X1 U7489 ( .A1(n9344), .A2(n9154), .ZN(n5860) );
  NAND2_X1 U7490 ( .A1(n9906), .A2(n8805), .ZN(n6093) );
  OR2_X1 U7491 ( .A1(n9845), .A2(P1_D_REG_0__SCAN_IN), .ZN(n5862) );
  NAND2_X1 U7492 ( .A1(n7162), .A2(n7010), .ZN(n5861) );
  AND2_X1 U7493 ( .A1(n5862), .A2(n5861), .ZN(n6003) );
  NOR4_X1 U7494 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n5866) );
  NOR4_X1 U7495 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n5865) );
  NOR4_X1 U7496 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5864) );
  NOR4_X1 U7497 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n5863) );
  NAND4_X1 U7498 ( .A1(n5866), .A2(n5865), .A3(n5864), .A4(n5863), .ZN(n5872)
         );
  NOR2_X1 U7499 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .ZN(
        n5870) );
  NOR4_X1 U7500 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n5869) );
  NOR4_X1 U7501 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n5868) );
  NOR4_X1 U7502 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n5867) );
  NAND4_X1 U7503 ( .A1(n5870), .A2(n5869), .A3(n5868), .A4(n5867), .ZN(n5871)
         );
  NOR2_X1 U7504 ( .A1(n5872), .A2(n5871), .ZN(n5873) );
  OR2_X1 U7505 ( .A1(n9845), .A2(n5873), .ZN(n6004) );
  NAND2_X1 U7506 ( .A1(n6003), .A2(n6004), .ZN(n7003) );
  NOR2_X1 U7507 ( .A1(n7003), .A2(n6993), .ZN(n6092) );
  AND2_X1 U7508 ( .A1(n6092), .A2(n9846), .ZN(n5877) );
  INV_X1 U7509 ( .A(n5877), .ZN(n5874) );
  OR2_X2 U7510 ( .A1(n6093), .A2(n5874), .ZN(n8672) );
  INV_X1 U7511 ( .A(n8672), .ZN(n8597) );
  NAND2_X1 U7512 ( .A1(n5875), .A2(n9154), .ZN(n6392) );
  NOR2_X1 U7513 ( .A1(n6392), .A2(n5876), .ZN(n8926) );
  AND2_X1 U7514 ( .A1(n5877), .A2(n8926), .ZN(n5938) );
  AND2_X1 U7515 ( .A1(n5938), .A2(n6257), .ZN(n8666) );
  INV_X1 U7516 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n5878) );
  INV_X1 U7517 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n6176) );
  AOI22_X1 U7518 ( .A1(n6253), .A2(n8597), .B1(n4397), .B2(n6007), .ZN(n5886)
         );
  INV_X1 U7519 ( .A(n8926), .ZN(n5880) );
  NAND2_X1 U7520 ( .A1(n6016), .A2(n5880), .ZN(n5882) );
  INV_X1 U7521 ( .A(n6092), .ZN(n5881) );
  NAND3_X1 U7522 ( .A1(n5882), .A2(n9846), .A3(n5881), .ZN(n6095) );
  OR2_X1 U7523 ( .A1(n8805), .A2(n5883), .ZN(n7005) );
  AND2_X1 U7524 ( .A1(n7005), .A2(n9846), .ZN(n5884) );
  OAI21_X1 U7525 ( .B1(n9664), .B2(n6092), .A(n8612), .ZN(n6105) );
  AOI22_X1 U7526 ( .A1(n6302), .A2(n8670), .B1(n6105), .B2(
        P1_REG3_REG_0__SCAN_IN), .ZN(n5885) );
  NAND2_X1 U7527 ( .A1(n5886), .A2(n5885), .ZN(P1_U3230) );
  INV_X1 U7528 ( .A(n9963), .ZN(n7618) );
  NAND2_X1 U7529 ( .A1(n5887), .A2(n7618), .ZN(n7653) );
  NAND2_X1 U7530 ( .A1(n7617), .A2(n7653), .ZN(n9965) );
  INV_X1 U7531 ( .A(n9965), .ZN(n5892) );
  INV_X1 U7532 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n9467) );
  AOI22_X1 U7533 ( .A1(n9965), .A2(n8395), .B1(n8392), .B2(n5808), .ZN(n9967)
         );
  OAI21_X1 U7534 ( .B1(n9467), .B2(n8356), .A(n9967), .ZN(n5889) );
  INV_X1 U7535 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n9607) );
  NOR2_X1 U7536 ( .A1(n9953), .A2(n9607), .ZN(n5888) );
  AOI21_X1 U7537 ( .B1(n9953), .B2(n5889), .A(n5888), .ZN(n5891) );
  OAI21_X1 U7538 ( .B1(n8359), .B2(n8402), .A(n9963), .ZN(n5890) );
  OAI211_X1 U7539 ( .C1(n5892), .C2(n8365), .A(n5891), .B(n5890), .ZN(P2_U3296) );
  INV_X1 U7540 ( .A(n8365), .ZN(n8409) );
  NAND2_X1 U7541 ( .A1(n7656), .A2(n7654), .ZN(n7819) );
  XOR2_X1 U7542 ( .A(n5893), .B(n7819), .Z(n9973) );
  AOI21_X1 U7543 ( .B1(n9963), .B2(n5233), .A(n5894), .ZN(n9969) );
  AOI22_X1 U7544 ( .A1(n8409), .A2(n9973), .B1(n8402), .B2(n9969), .ZN(n5903)
         );
  INV_X1 U7545 ( .A(n7654), .ZN(n5897) );
  INV_X1 U7546 ( .A(n7617), .ZN(n5895) );
  NAND2_X1 U7547 ( .A1(n7819), .A2(n5895), .ZN(n5896) );
  OAI211_X1 U7548 ( .C1(n7650), .C2(n5897), .A(n5896), .B(n8395), .ZN(n5900)
         );
  NAND2_X1 U7549 ( .A1(n5887), .A2(n8390), .ZN(n5899) );
  NAND2_X1 U7550 ( .A1(n5818), .A2(n8392), .ZN(n5898) );
  AND2_X1 U7551 ( .A1(n5899), .A2(n5898), .ZN(n6213) );
  NAND2_X1 U7552 ( .A1(n5900), .A2(n6213), .ZN(n9971) );
  AOI21_X1 U7553 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(n9944), .A(n9971), .ZN(
        n5901) );
  MUX2_X1 U7554 ( .A(n5689), .B(n5901), .S(n9953), .Z(n5902) );
  OAI211_X1 U7555 ( .C1(n5234), .C2(n8406), .A(n5903), .B(n5902), .ZN(P2_U3295) );
  NAND2_X1 U7556 ( .A1(n5904), .A2(n7820), .ZN(n5905) );
  NAND2_X1 U7557 ( .A1(n5906), .A2(n5905), .ZN(n5907) );
  NAND2_X1 U7558 ( .A1(n5907), .A2(n8395), .ZN(n5909) );
  AOI22_X1 U7559 ( .A1(n8390), .A2(n5808), .B1(n8068), .B2(n8392), .ZN(n5908)
         );
  NAND2_X1 U7560 ( .A1(n5909), .A2(n5908), .ZN(n9977) );
  INV_X1 U7561 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n9446) );
  OAI22_X1 U7562 ( .A1(n9446), .A2(n8356), .B1(n5910), .B2(n9953), .ZN(n5912)
         );
  OAI21_X1 U7563 ( .B1(n5894), .B2(n9975), .A(n6234), .ZN(n9976) );
  NOR2_X1 U7564 ( .A1(n8167), .A2(n9976), .ZN(n5911) );
  AOI211_X1 U7565 ( .C1(n9953), .C2(n9977), .A(n5912), .B(n5911), .ZN(n5916)
         );
  XNOR2_X1 U7566 ( .A(n5913), .B(n7820), .ZN(n9979) );
  AOI22_X1 U7567 ( .A1(n9979), .A2(n8409), .B1(n8359), .B2(n5914), .ZN(n5915)
         );
  NAND2_X1 U7568 ( .A1(n5916), .A2(n5915), .ZN(P2_U3294) );
  NAND2_X1 U7569 ( .A1(n6007), .A2(n6036), .ZN(n5920) );
  AND2_X4 U7570 ( .A1(n6392), .A2(n5876), .ZN(n7564) );
  INV_X1 U7571 ( .A(n6019), .ZN(n6023) );
  INV_X1 U7572 ( .A(n5922), .ZN(n5924) );
  NAND2_X1 U7573 ( .A1(n5926), .A2(n5925), .ZN(n6022) );
  INV_X4 U7574 ( .A(n5927), .ZN(n7566) );
  NAND2_X1 U7575 ( .A1(n6007), .A2(n7566), .ZN(n5929) );
  INV_X2 U7576 ( .A(n6036), .ZN(n6049) );
  OR2_X1 U7577 ( .A1(n6014), .A2(n6049), .ZN(n5928) );
  NAND2_X1 U7578 ( .A1(n5929), .A2(n5928), .ZN(n6020) );
  XNOR2_X1 U7579 ( .A(n6022), .B(n6020), .ZN(n5930) );
  XNOR2_X1 U7580 ( .A(n6023), .B(n5930), .ZN(n5943) );
  NOR2_X1 U7581 ( .A1(n9906), .A2(n6014), .ZN(n9851) );
  INV_X1 U7582 ( .A(n8666), .ZN(n8599) );
  INV_X1 U7583 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n5932) );
  OR2_X1 U7584 ( .A1(n4315), .A2(n5932), .ZN(n5936) );
  INV_X1 U7585 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n6264) );
  NAND2_X1 U7586 ( .A1(n4333), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5934) );
  INV_X1 U7587 ( .A(n5938), .ZN(n5939) );
  OR2_X1 U7588 ( .A1(n5939), .A2(n6257), .ZN(n8663) );
  OAI22_X1 U7589 ( .A1(n8599), .A2(n6379), .B1(n5851), .B2(n8663), .ZN(n5940)
         );
  AOI21_X1 U7590 ( .B1(n8612), .B2(n9851), .A(n5940), .ZN(n5942) );
  NAND2_X1 U7591 ( .A1(n6105), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5941) );
  OAI211_X1 U7592 ( .C1(n5943), .C2(n8672), .A(n5942), .B(n5941), .ZN(P1_U3220) );
  INV_X1 U7593 ( .A(n7308), .ZN(n6001) );
  OR2_X1 U7594 ( .A1(n5945), .A2(n5944), .ZN(n5946) );
  XNOR2_X1 U7595 ( .A(n5946), .B(P1_IR_REG_16__SCAN_IN), .ZN(n8952) );
  INV_X1 U7596 ( .A(n8952), .ZN(n7158) );
  OAI222_X1 U7597 ( .A1(n9373), .A2(n6001), .B1(n7158), .B2(P1_U3084), .C1(
        n5947), .C2(n9376), .ZN(P1_U3337) );
  INV_X1 U7598 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n5982) );
  NOR2_X1 U7599 ( .A1(n5948), .A2(P1_U3084), .ZN(n7194) );
  NAND2_X1 U7600 ( .A1(n9695), .A2(n7194), .ZN(n5960) );
  NOR2_X2 U7601 ( .A1(n5960), .A2(n6257), .ZN(n9751) );
  INV_X1 U7602 ( .A(n9737), .ZN(n5973) );
  INV_X1 U7603 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n5949) );
  MUX2_X1 U7604 ( .A(n5949), .B(P1_REG2_REG_6__SCAN_IN), .S(n9737), .Z(n5950)
         );
  INV_X1 U7605 ( .A(n5950), .ZN(n9733) );
  NOR2_X1 U7606 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(n5972), .ZN(n5951) );
  AOI21_X1 U7607 ( .B1(n5972), .B2(P1_REG2_REG_5__SCAN_IN), .A(n5951), .ZN(
        n9723) );
  INV_X1 U7608 ( .A(n6069), .ZN(n9701) );
  INV_X1 U7609 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n5952) );
  MUX2_X1 U7610 ( .A(n5952), .B(P1_REG2_REG_2__SCAN_IN), .S(n6029), .Z(n6269)
         );
  XNOR2_X1 U7611 ( .A(n5963), .B(P1_REG2_REG_1__SCAN_IN), .ZN(n6181) );
  AND2_X1 U7612 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n6255) );
  NAND2_X1 U7613 ( .A1(n6181), .A2(n6255), .ZN(n6180) );
  INV_X1 U7614 ( .A(n5963), .ZN(n6179) );
  NAND2_X1 U7615 ( .A1(n6179), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5953) );
  NAND2_X1 U7616 ( .A1(n6180), .A2(n5953), .ZN(n6268) );
  NAND2_X1 U7617 ( .A1(n6269), .A2(n6268), .ZN(n6267) );
  INV_X1 U7618 ( .A(n6029), .ZN(n6266) );
  NAND2_X1 U7619 ( .A1(n6266), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5954) );
  INV_X1 U7620 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n5955) );
  OR2_X1 U7621 ( .A1(n6160), .A2(n5955), .ZN(n5956) );
  XNOR2_X1 U7622 ( .A(n6069), .B(P1_REG2_REG_4__SCAN_IN), .ZN(n9700) );
  OAI21_X1 U7623 ( .B1(P1_REG2_REG_4__SCAN_IN), .B2(n9701), .A(n9698), .ZN(
        n9724) );
  NAND2_X1 U7624 ( .A1(n9723), .A2(n9724), .ZN(n9722) );
  NOR2_X1 U7625 ( .A1(P1_REG2_REG_7__SCAN_IN), .A2(n6349), .ZN(n5957) );
  AOI21_X1 U7626 ( .B1(n6349), .B2(P1_REG2_REG_7__SCAN_IN), .A(n5957), .ZN(
        n5958) );
  OAI21_X1 U7627 ( .B1(n5959), .B2(n5958), .A(n5983), .ZN(n5980) );
  INV_X1 U7628 ( .A(n6257), .ZN(n8925) );
  OR2_X1 U7629 ( .A1(n5960), .A2(n8925), .ZN(n9783) );
  OR2_X1 U7630 ( .A1(n6257), .A2(P1_U3084), .ZN(n7273) );
  INV_X1 U7631 ( .A(n5948), .ZN(n9686) );
  NOR2_X1 U7632 ( .A1(n7273), .A2(n9686), .ZN(n5961) );
  NAND2_X1 U7633 ( .A1(n9695), .A2(n5961), .ZN(n9744) );
  INV_X1 U7634 ( .A(n9744), .ZN(n9781) );
  NOR2_X1 U7635 ( .A1(P1_REG1_REG_7__SCAN_IN), .A2(n6349), .ZN(n5962) );
  AOI21_X1 U7636 ( .B1(n6349), .B2(P1_REG1_REG_7__SCAN_IN), .A(n5962), .ZN(
        n5975) );
  INV_X1 U7637 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6320) );
  MUX2_X1 U7638 ( .A(n6320), .B(P1_REG1_REG_6__SCAN_IN), .S(n9737), .Z(n9729)
         );
  MUX2_X1 U7639 ( .A(n5932), .B(P1_REG1_REG_2__SCAN_IN), .S(n6029), .Z(n6262)
         );
  XNOR2_X1 U7640 ( .A(n5963), .B(P1_REG1_REG_1__SCAN_IN), .ZN(n6175) );
  AND2_X1 U7641 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n6174) );
  NAND2_X1 U7642 ( .A1(n6175), .A2(n6174), .ZN(n6173) );
  NAND2_X1 U7643 ( .A1(n6179), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5964) );
  NAND2_X1 U7644 ( .A1(n6173), .A2(n5964), .ZN(n6261) );
  NAND2_X1 U7645 ( .A1(n6262), .A2(n6261), .ZN(n6260) );
  NAND2_X1 U7646 ( .A1(n6266), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5965) );
  NAND2_X1 U7647 ( .A1(n6260), .A2(n5965), .ZN(n6162) );
  INV_X1 U7648 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n9919) );
  MUX2_X1 U7649 ( .A(n9919), .B(P1_REG1_REG_3__SCAN_IN), .S(n6160), .Z(n6163)
         );
  AND2_X1 U7650 ( .A1(n6162), .A2(n6163), .ZN(n9705) );
  INV_X1 U7651 ( .A(n9705), .ZN(n6161) );
  INV_X1 U7652 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6061) );
  XNOR2_X1 U7653 ( .A(n6069), .B(n6061), .ZN(n9703) );
  INV_X1 U7654 ( .A(n9703), .ZN(n5967) );
  NOR2_X1 U7655 ( .A1(n6160), .A2(n9919), .ZN(n9704) );
  INV_X1 U7656 ( .A(n9704), .ZN(n5966) );
  AND2_X1 U7657 ( .A1(n5967), .A2(n5966), .ZN(n5968) );
  NAND2_X1 U7658 ( .A1(n6161), .A2(n5968), .ZN(n9707) );
  NAND2_X1 U7659 ( .A1(n6069), .A2(n6061), .ZN(n5969) );
  NAND2_X1 U7660 ( .A1(n9707), .A2(n5969), .ZN(n9716) );
  OR2_X1 U7661 ( .A1(n5972), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5971) );
  NAND2_X1 U7662 ( .A1(P1_REG1_REG_5__SCAN_IN), .A2(n5972), .ZN(n5970) );
  NAND2_X1 U7663 ( .A1(n5971), .A2(n5970), .ZN(n9715) );
  NOR2_X1 U7664 ( .A1(n9716), .A2(n9715), .ZN(n9718) );
  AOI21_X1 U7665 ( .B1(n5972), .B2(P1_REG1_REG_5__SCAN_IN), .A(n9718), .ZN(
        n9730) );
  NAND2_X1 U7666 ( .A1(n9729), .A2(n9730), .ZN(n9728) );
  OAI21_X1 U7667 ( .B1(P1_REG1_REG_6__SCAN_IN), .B2(n5973), .A(n9728), .ZN(
        n5974) );
  NAND2_X1 U7668 ( .A1(n5975), .A2(n5974), .ZN(n5989) );
  OAI21_X1 U7669 ( .B1(n5975), .B2(n5974), .A(n5989), .ZN(n5976) );
  AND2_X1 U7670 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n6367) );
  AOI21_X1 U7671 ( .B1(n9781), .B2(n5976), .A(n6367), .ZN(n5977) );
  OAI21_X1 U7672 ( .B1(n5978), .B2(n9783), .A(n5977), .ZN(n5979) );
  AOI21_X1 U7673 ( .B1(n9751), .B2(n5980), .A(n5979), .ZN(n5981) );
  OAI21_X1 U7674 ( .B1(n9785), .B2(n5982), .A(n5981), .ZN(P1_U3248) );
  INV_X1 U7675 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n6000) );
  XNOR2_X1 U7676 ( .A(n6580), .B(P1_REG2_REG_8__SCAN_IN), .ZN(n9743) );
  OAI21_X1 U7677 ( .B1(P1_REG2_REG_7__SCAN_IN), .B2(n6349), .A(n5983), .ZN(
        n5984) );
  INV_X1 U7678 ( .A(n5984), .ZN(n9742) );
  OAI22_X1 U7679 ( .A1(n9743), .A2(n9742), .B1(n6580), .B2(
        P1_REG2_REG_8__SCAN_IN), .ZN(n9765) );
  NAND2_X1 U7680 ( .A1(n9757), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5985) );
  OAI21_X1 U7681 ( .B1(n9757), .B2(P1_REG2_REG_9__SCAN_IN), .A(n5985), .ZN(
        n9764) );
  NOR2_X1 U7682 ( .A1(n9765), .A2(n9764), .ZN(n9763) );
  XNOR2_X1 U7683 ( .A(n6830), .B(P1_REG2_REG_10__SCAN_IN), .ZN(n9776) );
  INV_X1 U7684 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n5986) );
  AOI22_X1 U7685 ( .A1(P1_REG2_REG_11__SCAN_IN), .A2(n7070), .B1(n5996), .B2(
        n5986), .ZN(n5987) );
  OAI21_X1 U7686 ( .B1(n5988), .B2(n5987), .A(n6152), .ZN(n5998) );
  INV_X1 U7687 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n9677) );
  AOI22_X1 U7688 ( .A1(P1_REG1_REG_11__SCAN_IN), .A2(n7070), .B1(n5996), .B2(
        n9677), .ZN(n5993) );
  INV_X1 U7689 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6766) );
  MUX2_X1 U7690 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n6766), .S(n6830), .Z(n9772)
         );
  XNOR2_X1 U7691 ( .A(n6580), .B(P1_REG1_REG_8__SCAN_IN), .ZN(n9747) );
  OR2_X1 U7692 ( .A1(n6349), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5990) );
  NAND2_X1 U7693 ( .A1(n5990), .A2(n5989), .ZN(n9746) );
  NOR2_X1 U7694 ( .A1(n9747), .A2(n9746), .ZN(n9745) );
  AOI21_X1 U7695 ( .B1(P1_REG1_REG_8__SCAN_IN), .B2(n6580), .A(n9745), .ZN(
        n9762) );
  NOR2_X1 U7696 ( .A1(n9757), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5991) );
  AOI21_X1 U7697 ( .B1(P1_REG1_REG_9__SCAN_IN), .B2(n9757), .A(n5991), .ZN(
        n9761) );
  NAND2_X1 U7698 ( .A1(n9762), .A2(n9761), .ZN(n9760) );
  OAI21_X1 U7699 ( .B1(n9757), .B2(P1_REG1_REG_9__SCAN_IN), .A(n9760), .ZN(
        n9773) );
  NAND2_X1 U7700 ( .A1(n9772), .A2(n9773), .ZN(n9771) );
  OAI21_X1 U7701 ( .B1(P1_REG1_REG_10__SCAN_IN), .B2(n6830), .A(n9771), .ZN(
        n5992) );
  NAND2_X1 U7702 ( .A1(n5993), .A2(n5992), .ZN(n6141) );
  OAI21_X1 U7703 ( .B1(n5993), .B2(n5992), .A(n6141), .ZN(n5994) );
  AND2_X1 U7704 ( .A1(P1_U3084), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n7196) );
  AOI21_X1 U7705 ( .B1(n9781), .B2(n5994), .A(n7196), .ZN(n5995) );
  OAI21_X1 U7706 ( .B1(n5996), .B2(n9783), .A(n5995), .ZN(n5997) );
  AOI21_X1 U7707 ( .B1(n9751), .B2(n5998), .A(n5997), .ZN(n5999) );
  OAI21_X1 U7708 ( .B1(n9785), .B2(n6000), .A(n5999), .ZN(P1_U3252) );
  INV_X1 U7709 ( .A(n8112), .ZN(n6885) );
  OAI222_X1 U7710 ( .A1(n8534), .A2(n6002), .B1(n7939), .B2(n6001), .C1(n6885), 
        .C2(P2_U3152), .ZN(P2_U3342) );
  NOR2_X1 U7711 ( .A1(n6003), .A2(n9850), .ZN(n9848) );
  NAND2_X1 U7712 ( .A1(n6995), .A2(n6005), .ZN(n6523) );
  OR2_X1 U7713 ( .A1(n9344), .A2(n6996), .ZN(n9908) );
  OR2_X1 U7714 ( .A1(n9850), .A2(n9154), .ZN(n6006) );
  AND2_X2 U7715 ( .A1(n6523), .A2(n9809), .ZN(n9844) );
  INV_X2 U7716 ( .A(n9844), .ZN(n9814) );
  NOR2_X1 U7717 ( .A1(n8926), .A2(n7564), .ZN(n9842) );
  NAND2_X1 U7718 ( .A1(n9814), .A2(n9842), .ZN(n9256) );
  NAND2_X1 U7719 ( .A1(n6009), .A2(n6008), .ZN(n6378) );
  OAI21_X1 U7720 ( .B1(n6008), .B2(n6009), .A(n6378), .ZN(n9854) );
  INV_X1 U7721 ( .A(n8805), .ZN(n6010) );
  INV_X1 U7722 ( .A(n6302), .ZN(n9345) );
  NOR2_X1 U7723 ( .A1(n6298), .A2(n9345), .ZN(n6387) );
  XNOR2_X1 U7724 ( .A(n6008), .B(n6387), .ZN(n6013) );
  INV_X1 U7725 ( .A(n9154), .ZN(n9840) );
  NAND2_X1 U7726 ( .A1(n5875), .A2(n9840), .ZN(n6012) );
  OR2_X1 U7727 ( .A1(n5842), .A2(n5844), .ZN(n6011) );
  OAI222_X1 U7728 ( .A1(n9802), .A2(n5851), .B1(n9800), .B2(n6379), .C1(n6013), 
        .C2(n9242), .ZN(n9856) );
  INV_X1 U7729 ( .A(n9908), .ZN(n9881) );
  OAI211_X1 U7730 ( .C1(n9345), .C2(n6014), .A(n9881), .B(n6384), .ZN(n9853)
         );
  OAI22_X1 U7731 ( .A1(n9853), .A2(n9840), .B1(n9809), .B2(n6176), .ZN(n6015)
         );
  OAI21_X1 U7732 ( .B1(n9856), .B2(n6015), .A(n9814), .ZN(n6018) );
  INV_X1 U7733 ( .A(n6016), .ZN(n9836) );
  AOI22_X1 U7734 ( .A1(n9174), .A2(n6388), .B1(n9844), .B2(
        P1_REG2_REG_1__SCAN_IN), .ZN(n6017) );
  OAI211_X1 U7735 ( .C1(n9256), .C2(n9854), .A(n6018), .B(n6017), .ZN(P1_U3290) );
  NAND2_X1 U7736 ( .A1(n6022), .A2(n6019), .ZN(n6021) );
  NAND2_X1 U7737 ( .A1(n6021), .A2(n6020), .ZN(n6026) );
  INV_X1 U7738 ( .A(n6022), .ZN(n6024) );
  NAND2_X1 U7739 ( .A1(n6024), .A2(n6023), .ZN(n6025) );
  NAND2_X1 U7740 ( .A1(n8944), .A2(n6036), .ZN(n6034) );
  OR2_X1 U7741 ( .A1(n6067), .A2(n6027), .ZN(n6032) );
  OR2_X1 U7742 ( .A1(n6350), .A2(n6028), .ZN(n6031) );
  NAND2_X1 U7743 ( .A1(n8891), .A2(n7579), .ZN(n6033) );
  NAND2_X1 U7744 ( .A1(n6034), .A2(n6033), .ZN(n6035) );
  XNOR2_X1 U7745 ( .A(n6035), .B(n7564), .ZN(n6041) );
  INV_X1 U7746 ( .A(n6041), .ZN(n6039) );
  AND2_X1 U7747 ( .A1(n8891), .A2(n6036), .ZN(n6037) );
  AOI21_X1 U7748 ( .B1(n8944), .B2(n7566), .A(n6037), .ZN(n6040) );
  INV_X1 U7749 ( .A(n6040), .ZN(n6038) );
  NAND2_X1 U7750 ( .A1(n6041), .A2(n6040), .ZN(n6043) );
  NAND2_X1 U7751 ( .A1(n4333), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n6048) );
  OR2_X1 U7752 ( .A1(n4316), .A2(n9919), .ZN(n6047) );
  OR2_X1 U7753 ( .A1(n5933), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n6046) );
  OR2_X1 U7754 ( .A1(n7598), .A2(n5955), .ZN(n6045) );
  NAND2_X1 U7755 ( .A1(n8942), .A2(n6036), .ZN(n6057) );
  OR2_X1 U7756 ( .A1(n6350), .A2(n6050), .ZN(n6054) );
  OR2_X1 U7757 ( .A1(n6067), .A2(n6051), .ZN(n6053) );
  OR2_X1 U7758 ( .A1(n6030), .A2(n6160), .ZN(n6052) );
  OR2_X1 U7759 ( .A1(n9863), .A2(n6055), .ZN(n6056) );
  NAND2_X1 U7760 ( .A1(n6057), .A2(n6056), .ZN(n6058) );
  XNOR2_X1 U7761 ( .A(n6058), .B(n7564), .ZN(n6060) );
  INV_X1 U7762 ( .A(n9863), .ZN(n7288) );
  AOI22_X1 U7763 ( .A1(n8942), .A2(n7566), .B1(n7288), .B2(n7592), .ZN(n6059)
         );
  AND2_X1 U7764 ( .A1(n6060), .A2(n6059), .ZN(n7279) );
  OR2_X1 U7765 ( .A1(n6060), .A2(n6059), .ZN(n7280) );
  NAND2_X1 U7766 ( .A1(n7555), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n6065) );
  OR2_X1 U7767 ( .A1(n4316), .A2(n6061), .ZN(n6064) );
  XNOR2_X1 U7768 ( .A(P1_REG3_REG_3__SCAN_IN), .B(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n6442) );
  OR2_X1 U7769 ( .A1(n5933), .A2(n6442), .ZN(n6063) );
  INV_X1 U7770 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6443) );
  OR2_X1 U7771 ( .A1(n7598), .A2(n6443), .ZN(n6062) );
  NAND2_X1 U7772 ( .A1(n9826), .A2(n7566), .ZN(n6074) );
  OR2_X1 U7773 ( .A1(n6350), .A2(n6066), .ZN(n6072) );
  OR2_X1 U7774 ( .A1(n6067), .A2(n6068), .ZN(n6071) );
  OR2_X1 U7775 ( .A1(n6030), .A2(n6069), .ZN(n6070) );
  OR2_X1 U7776 ( .A1(n9869), .A2(n6049), .ZN(n6073) );
  NAND2_X1 U7777 ( .A1(n6074), .A2(n6073), .ZN(n6305) );
  NAND2_X1 U7778 ( .A1(n9826), .A2(n7568), .ZN(n6076) );
  OR2_X1 U7779 ( .A1(n9869), .A2(n6055), .ZN(n6075) );
  NAND2_X1 U7780 ( .A1(n6076), .A2(n6075), .ZN(n6077) );
  XNOR2_X1 U7781 ( .A(n6077), .B(n5923), .ZN(n6306) );
  XOR2_X1 U7782 ( .A(n6305), .B(n6306), .Z(n6078) );
  XNOR2_X1 U7783 ( .A(n6307), .B(n6078), .ZN(n6100) );
  INV_X1 U7784 ( .A(n9869), .ZN(n6448) );
  AOI21_X1 U7785 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(P1_REG3_REG_5__SCAN_IN), .ZN(n6079) );
  NOR2_X1 U7786 ( .A1(n6079), .A2(n6321), .ZN(n9837) );
  NAND2_X1 U7787 ( .A1(n7554), .A2(n9837), .ZN(n6087) );
  INV_X1 U7788 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n6080) );
  OR2_X1 U7789 ( .A1(n7600), .A2(n6080), .ZN(n6086) );
  INV_X1 U7790 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6082) );
  OR2_X1 U7791 ( .A1(n4316), .A2(n6082), .ZN(n6085) );
  INV_X1 U7792 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n6083) );
  OR2_X1 U7793 ( .A1(n7598), .A2(n6083), .ZN(n6084) );
  NAND4_X1 U7794 ( .A1(n6087), .A2(n6086), .A3(n6085), .A4(n6084), .ZN(n8941)
         );
  INV_X1 U7795 ( .A(n8941), .ZN(n6432) );
  INV_X1 U7796 ( .A(n8663), .ZN(n8621) );
  AND2_X1 U7797 ( .A1(P1_U3084), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n9709) );
  AOI21_X1 U7798 ( .B1(n8621), .B2(n8942), .A(n9709), .ZN(n6088) );
  OAI21_X1 U7799 ( .B1(n8599), .B2(n6432), .A(n6088), .ZN(n6098) );
  AND3_X1 U7800 ( .A1(n7005), .A2(n6090), .A3(n6089), .ZN(n6091) );
  OAI21_X1 U7801 ( .B1(n6093), .B2(n6092), .A(n6091), .ZN(n6094) );
  NAND2_X1 U7802 ( .A1(n6094), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6096) );
  NOR2_X1 U7803 ( .A1(n8668), .A2(n6442), .ZN(n6097) );
  AOI211_X1 U7804 ( .C1(n8670), .C2(n6448), .A(n6098), .B(n6097), .ZN(n6099)
         );
  OAI21_X1 U7805 ( .B1(n6100), .B2(n8672), .A(n6099), .ZN(P1_U3228) );
  INV_X1 U7806 ( .A(n8670), .ZN(n8658) );
  OAI21_X1 U7807 ( .B1(n6102), .B2(n4396), .A(n6101), .ZN(n6103) );
  NAND2_X1 U7808 ( .A1(n6103), .A2(n8597), .ZN(n6107) );
  INV_X1 U7809 ( .A(n6007), .ZN(n6389) );
  OAI22_X1 U7810 ( .A1(n8599), .A2(n6400), .B1(n6389), .B2(n8663), .ZN(n6104)
         );
  AOI21_X1 U7811 ( .B1(P1_REG3_REG_2__SCAN_IN), .B2(n6105), .A(n6104), .ZN(
        n6106) );
  OAI211_X1 U7812 ( .C1(n6380), .C2(n8658), .A(n6107), .B(n6106), .ZN(P1_U3235) );
  INV_X1 U7813 ( .A(n7318), .ZN(n6224) );
  NAND2_X1 U7814 ( .A1(n6108), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6275) );
  XNOR2_X1 U7815 ( .A(n6275), .B(P1_IR_REG_17__SCAN_IN), .ZN(n8969) );
  AOI22_X1 U7816 ( .A1(n8969), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n9366), .ZN(n6109) );
  OAI21_X1 U7817 ( .B1(n6224), .B2(n9373), .A(n6109), .ZN(P1_U3336) );
  INV_X1 U7818 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n6110) );
  MUX2_X1 U7819 ( .A(P2_REG2_REG_13__SCAN_IN), .B(n6110), .S(n6291), .Z(n6111)
         );
  INV_X1 U7820 ( .A(n6111), .ZN(n6116) );
  AOI21_X1 U7821 ( .B1(n6116), .B2(n6115), .A(n6282), .ZN(n6128) );
  INV_X1 U7822 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n6117) );
  MUX2_X1 U7823 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n6117), .S(n6291), .Z(n6122)
         );
  INV_X1 U7824 ( .A(n6118), .ZN(n6119) );
  OAI21_X1 U7825 ( .B1(n6120), .B2(P2_REG1_REG_12__SCAN_IN), .A(n6119), .ZN(
        n6121) );
  NAND2_X1 U7826 ( .A1(n6121), .A2(n6122), .ZN(n6290) );
  OAI21_X1 U7827 ( .B1(n6122), .B2(n6121), .A(n6290), .ZN(n6123) );
  NAND2_X1 U7828 ( .A1(n6123), .A2(n9930), .ZN(n6127) );
  NOR2_X1 U7829 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5326), .ZN(n6910) );
  INV_X1 U7830 ( .A(n6291), .ZN(n6124) );
  NOR2_X1 U7831 ( .A1(n9932), .A2(n6124), .ZN(n6125) );
  AOI211_X1 U7832 ( .C1(P2_ADDR_REG_13__SCAN_IN), .C2(n9935), .A(n6910), .B(
        n6125), .ZN(n6126) );
  OAI211_X1 U7833 ( .C1(n6128), .C2(n9933), .A(n6127), .B(n6126), .ZN(P2_U3258) );
  OAI21_X1 U7834 ( .B1(n6131), .B2(n6130), .A(n6129), .ZN(n9985) );
  INV_X1 U7835 ( .A(n9985), .ZN(n6139) );
  OAI22_X1 U7836 ( .A1(n6203), .A2(n8356), .B1(n5712), .B2(n9953), .ZN(n6133)
         );
  OAI21_X1 U7837 ( .B1(n6236), .B2(n9981), .A(n6691), .ZN(n9982) );
  NOR2_X1 U7838 ( .A1(n8167), .A2(n9982), .ZN(n6132) );
  AOI211_X1 U7839 ( .C1(n8359), .C2(n6206), .A(n6133), .B(n6132), .ZN(n6138)
         );
  NAND2_X1 U7840 ( .A1(n6134), .A2(n7822), .ZN(n6688) );
  OAI211_X1 U7841 ( .C1(n6134), .C2(n7822), .A(n6688), .B(n8395), .ZN(n6136)
         );
  AOI22_X1 U7842 ( .A1(n8390), .A2(n8068), .B1(n8065), .B2(n8392), .ZN(n6135)
         );
  NAND2_X1 U7843 ( .A1(n6136), .A2(n6135), .ZN(n9983) );
  NAND2_X1 U7844 ( .A1(n9983), .A2(n9953), .ZN(n6137) );
  OAI211_X1 U7845 ( .C1(n6139), .C2(n8365), .A(n6138), .B(n6137), .ZN(P2_U3292) );
  NAND2_X1 U7846 ( .A1(n8055), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n6140) );
  OAI21_X1 U7847 ( .B1(n8158), .B2(n8055), .A(n6140), .ZN(P2_U3581) );
  INV_X1 U7848 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n6159) );
  INV_X1 U7849 ( .A(n9783), .ZN(n9758) );
  INV_X1 U7850 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n7078) );
  OR2_X1 U7851 ( .A1(n7070), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n6142) );
  NAND2_X1 U7852 ( .A1(n6142), .A2(n6141), .ZN(n6532) );
  NAND2_X1 U7853 ( .A1(n7074), .A2(n7078), .ZN(n6143) );
  OAI21_X1 U7854 ( .B1(n7074), .B2(n7078), .A(n6143), .ZN(n6144) );
  INV_X1 U7855 ( .A(n6144), .ZN(n6533) );
  NAND2_X1 U7856 ( .A1(n6532), .A2(n6533), .ZN(n6531) );
  INV_X1 U7857 ( .A(n6531), .ZN(n6145) );
  AOI21_X1 U7858 ( .B1(n7074), .B2(n7078), .A(n6145), .ZN(n6147) );
  INV_X1 U7859 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n9661) );
  MUX2_X1 U7860 ( .A(n9661), .B(P1_REG1_REG_13__SCAN_IN), .S(n7169), .Z(n6146)
         );
  NOR2_X1 U7861 ( .A1(n6147), .A2(n6146), .ZN(n6700) );
  AOI21_X1 U7862 ( .B1(n6147), .B2(n6146), .A(n6700), .ZN(n6148) );
  NAND2_X1 U7863 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n7184) );
  OAI21_X1 U7864 ( .B1(n6148), .B2(n9744), .A(n7184), .ZN(n6149) );
  AOI21_X1 U7865 ( .B1(n7169), .B2(n9758), .A(n6149), .ZN(n6158) );
  OR2_X1 U7866 ( .A1(n7169), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n6151) );
  NAND2_X1 U7867 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n7169), .ZN(n6150) );
  AND2_X1 U7868 ( .A1(n6151), .A2(n6150), .ZN(n6156) );
  OR2_X1 U7869 ( .A1(n7070), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6153) );
  NAND2_X1 U7870 ( .A1(n6153), .A2(n6152), .ZN(n6538) );
  INV_X1 U7871 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7081) );
  XNOR2_X1 U7872 ( .A(n7074), .B(n7081), .ZN(n6539) );
  INV_X1 U7873 ( .A(n6707), .ZN(n6154) );
  OAI211_X1 U7874 ( .C1(n6156), .C2(n6155), .A(n9751), .B(n6154), .ZN(n6157)
         );
  OAI211_X1 U7875 ( .C1(n6159), .C2(n9785), .A(n6158), .B(n6157), .ZN(P1_U3254) );
  INV_X1 U7876 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n6172) );
  INV_X1 U7877 ( .A(n6160), .ZN(n6166) );
  OAI21_X1 U7878 ( .B1(n6163), .B2(n6162), .A(n6161), .ZN(n6164) );
  INV_X1 U7879 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n6405) );
  OR2_X1 U7880 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6405), .ZN(n7284) );
  OAI21_X1 U7881 ( .B1(n9744), .B2(n6164), .A(n7284), .ZN(n6165) );
  AOI21_X1 U7882 ( .B1(n9758), .B2(n6166), .A(n6165), .ZN(n6171) );
  OAI211_X1 U7883 ( .C1(n6169), .C2(n6168), .A(n9751), .B(n6167), .ZN(n6170)
         );
  OAI211_X1 U7884 ( .C1(n6172), .C2(n9785), .A(n6171), .B(n6170), .ZN(P1_U3244) );
  INV_X1 U7885 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n6184) );
  OAI21_X1 U7886 ( .B1(n6175), .B2(n6174), .A(n6173), .ZN(n6177) );
  OAI22_X1 U7887 ( .A1(n9744), .A2(n6177), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6176), .ZN(n6178) );
  AOI21_X1 U7888 ( .B1(n6179), .B2(n9758), .A(n6178), .ZN(n6183) );
  OAI211_X1 U7889 ( .C1(n6181), .C2(n6255), .A(n9751), .B(n6180), .ZN(n6182)
         );
  OAI211_X1 U7890 ( .C1(n6184), .C2(n9785), .A(n6183), .B(n6182), .ZN(P1_U3242) );
  XNOR2_X1 U7891 ( .A(n7926), .B(n6495), .ZN(n6190) );
  NAND2_X1 U7892 ( .A1(n8068), .A2(n7635), .ZN(n6189) );
  XNOR2_X1 U7893 ( .A(n6190), .B(n6189), .ZN(n6218) );
  INV_X1 U7894 ( .A(n6189), .ZN(n6191) );
  NAND2_X1 U7895 ( .A1(n6191), .A2(n6190), .ZN(n6192) );
  AND2_X1 U7896 ( .A1(n8067), .A2(n7635), .ZN(n6194) );
  XNOR2_X1 U7897 ( .A(n7926), .B(n6206), .ZN(n6193) );
  NAND2_X1 U7898 ( .A1(n6194), .A2(n6193), .ZN(n6197) );
  INV_X1 U7899 ( .A(n6193), .ZN(n6196) );
  INV_X1 U7900 ( .A(n6194), .ZN(n6195) );
  NAND2_X1 U7901 ( .A1(n6196), .A2(n6195), .ZN(n6244) );
  NAND2_X1 U7902 ( .A1(n6197), .A2(n6244), .ZN(n6200) );
  INV_X1 U7903 ( .A(n6200), .ZN(n6198) );
  INV_X1 U7904 ( .A(n6245), .ZN(n6199) );
  AOI21_X1 U7905 ( .B1(n6201), .B2(n6200), .A(n6199), .ZN(n6209) );
  NAND2_X1 U7906 ( .A1(n6202), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8045) );
  NOR2_X1 U7907 ( .A1(n8045), .A2(n6203), .ZN(n6204) );
  AOI211_X1 U7908 ( .C1(n8047), .C2(n6206), .A(n6205), .B(n6204), .ZN(n6208)
         );
  AOI22_X1 U7909 ( .A1(n6609), .A2(n8068), .B1(n6608), .B2(n8065), .ZN(n6207)
         );
  OAI211_X1 U7910 ( .C1(n6209), .C2(n8036), .A(n6208), .B(n6207), .ZN(P2_U3232) );
  INV_X1 U7911 ( .A(n7621), .ZN(n6217) );
  INV_X1 U7912 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n9560) );
  OAI21_X1 U7913 ( .B1(n6212), .B2(n6211), .A(n6210), .ZN(n6215) );
  INV_X1 U7914 ( .A(n8043), .ZN(n8022) );
  OAI22_X1 U7915 ( .A1(n8026), .A2(n5234), .B1(n6213), .B2(n8022), .ZN(n6214)
         );
  AOI21_X1 U7916 ( .B1(n8038), .B2(n6215), .A(n6214), .ZN(n6216) );
  OAI21_X1 U7917 ( .B1(n6217), .B2(n9560), .A(n6216), .ZN(P2_U3224) );
  XNOR2_X1 U7918 ( .A(n6219), .B(n6218), .ZN(n6223) );
  OAI22_X1 U7919 ( .A1(n5242), .A2(n8030), .B1(n8029), .B2(n6247), .ZN(n6221)
         );
  OAI22_X1 U7920 ( .A1(n8026), .A2(n7670), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9534), .ZN(n6220) );
  AOI211_X1 U7921 ( .C1(n8033), .C2(n9534), .A(n6221), .B(n6220), .ZN(n6222)
         );
  OAI21_X1 U7922 ( .B1(n8036), .B2(n6223), .A(n6222), .ZN(P2_U3220) );
  INV_X1 U7923 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n6225) );
  INV_X1 U7924 ( .A(n8125), .ZN(n8119) );
  OAI222_X1 U7925 ( .A1(n8534), .A2(n6225), .B1(n7939), .B2(n6224), .C1(n8119), 
        .C2(P2_U3152), .ZN(P2_U3341) );
  INV_X1 U7926 ( .A(n8379), .ZN(n6233) );
  OAI21_X1 U7927 ( .B1(n6227), .B2(n6228), .A(n6226), .ZN(n6238) );
  INV_X1 U7928 ( .A(n8390), .ZN(n8305) );
  OAI22_X1 U7929 ( .A1(n5242), .A2(n8305), .B1(n6247), .B2(n8307), .ZN(n6232)
         );
  XNOR2_X1 U7930 ( .A(n6229), .B(n6228), .ZN(n6230) );
  INV_X1 U7931 ( .A(n8395), .ZN(n8347) );
  NOR2_X1 U7932 ( .A1(n6230), .A2(n8347), .ZN(n6231) );
  AOI211_X1 U7933 ( .C1(n6233), .C2(n6238), .A(n6232), .B(n6231), .ZN(n6498)
         );
  AND2_X1 U7934 ( .A1(n6234), .A2(n6495), .ZN(n6235) );
  NOR2_X1 U7935 ( .A1(n6236), .A2(n6235), .ZN(n6496) );
  INV_X1 U7936 ( .A(n6496), .ZN(n6237) );
  OAI22_X1 U7937 ( .A1(n8167), .A2(n6237), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n8356), .ZN(n6242) );
  INV_X1 U7938 ( .A(n6238), .ZN(n6499) );
  INV_X1 U7939 ( .A(n6239), .ZN(n6240) );
  NAND2_X1 U7940 ( .A1(n9953), .A2(n6240), .ZN(n8388) );
  OAI22_X1 U7941 ( .A1(n6499), .A2(n8388), .B1(n7670), .B2(n8406), .ZN(n6241)
         );
  AOI211_X1 U7942 ( .C1(n8368), .C2(P2_REG2_REG_3__SCAN_IN), .A(n6242), .B(
        n6241), .ZN(n6243) );
  OAI21_X1 U7943 ( .B1(n6498), .B2(n8368), .A(n6243), .ZN(P2_U3293) );
  XNOR2_X1 U7944 ( .A(n7926), .B(n6248), .ZN(n6483) );
  NAND2_X1 U7945 ( .A1(n8065), .A2(n7635), .ZN(n6482) );
  XNOR2_X1 U7946 ( .A(n6483), .B(n6482), .ZN(n6545) );
  XNOR2_X1 U7947 ( .A(n6546), .B(n6545), .ZN(n6252) );
  OAI22_X1 U7948 ( .A1(n6247), .A2(n8030), .B1(n8029), .B2(n6246), .ZN(n6250)
         );
  OAI22_X1 U7949 ( .A1(n8026), .A2(n6248), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5257), .ZN(n6249) );
  AOI211_X1 U7950 ( .C1(n9943), .C2(n8033), .A(n6250), .B(n6249), .ZN(n6251)
         );
  OAI21_X1 U7951 ( .B1(n6252), .B2(n8036), .A(n6251), .ZN(P2_U3229) );
  INV_X1 U7952 ( .A(n6253), .ZN(n6254) );
  MUX2_X1 U7953 ( .A(n6255), .B(n6254), .S(n5948), .Z(n6259) );
  INV_X1 U7954 ( .A(n6256), .ZN(n6258) );
  AOI21_X1 U7955 ( .B1(n9686), .B2(n5666), .A(n6257), .ZN(n9690) );
  OAI21_X1 U7956 ( .B1(n9690), .B2(P1_IR_REG_0__SCAN_IN), .A(
        P1_STATE_REG_SCAN_IN), .ZN(n9687) );
  AOI211_X1 U7957 ( .C1(n6259), .C2(n8925), .A(n6258), .B(n9687), .ZN(n9710)
         );
  INV_X1 U7958 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n6272) );
  OAI211_X1 U7959 ( .C1(n6262), .C2(n6261), .A(n9781), .B(n6260), .ZN(n6263)
         );
  OAI21_X1 U7960 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n6264), .A(n6263), .ZN(n6265) );
  AOI21_X1 U7961 ( .B1(n6266), .B2(n9758), .A(n6265), .ZN(n6271) );
  OAI211_X1 U7962 ( .C1(n6269), .C2(n6268), .A(n9751), .B(n6267), .ZN(n6270)
         );
  OAI211_X1 U7963 ( .C1(n6272), .C2(n9785), .A(n6271), .B(n6270), .ZN(n6273)
         );
  OR2_X1 U7964 ( .A1(n9710), .A2(n6273), .ZN(P1_U3243) );
  INV_X1 U7965 ( .A(n7332), .ZN(n6281) );
  NAND2_X1 U7966 ( .A1(n6275), .A2(n6274), .ZN(n6276) );
  NAND2_X1 U7967 ( .A1(n6276), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6277) );
  XNOR2_X1 U7968 ( .A(n6277), .B(P1_IR_REG_18__SCAN_IN), .ZN(n8979) );
  AOI22_X1 U7969 ( .A1(n8979), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n9366), .ZN(n6278) );
  OAI21_X1 U7970 ( .B1(n6281), .B2(n9373), .A(n6278), .ZN(P1_U3335) );
  AOI22_X1 U7971 ( .A1(n8135), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n6279), .ZN(n6280) );
  OAI21_X1 U7972 ( .B1(n6281), .B2(n7939), .A(n6280), .ZN(P2_U3340) );
  NOR2_X1 U7973 ( .A1(n6291), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n6283) );
  INV_X1 U7974 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n6714) );
  AOI22_X1 U7975 ( .A1(n6718), .A2(n6714), .B1(P2_REG2_REG_14__SCAN_IN), .B2(
        n6715), .ZN(n6284) );
  AOI21_X1 U7976 ( .B1(n6285), .B2(n6284), .A(n6713), .ZN(n6297) );
  INV_X1 U7977 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n6287) );
  AND2_X1 U7978 ( .A1(P2_U3152), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n7057) );
  INV_X1 U7979 ( .A(n7057), .ZN(n6286) );
  OAI21_X1 U7980 ( .B1(n9604), .B2(n6287), .A(n6286), .ZN(n6288) );
  AOI21_X1 U7981 ( .B1(n9619), .B2(n6718), .A(n6288), .ZN(n6296) );
  INV_X1 U7982 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n6289) );
  AOI22_X1 U7983 ( .A1(n6718), .A2(P2_REG1_REG_14__SCAN_IN), .B1(n6289), .B2(
        n6715), .ZN(n6293) );
  OAI21_X1 U7984 ( .B1(n6291), .B2(P2_REG1_REG_13__SCAN_IN), .A(n6290), .ZN(
        n6292) );
  NAND2_X1 U7985 ( .A1(n6293), .A2(n6292), .ZN(n6717) );
  OAI21_X1 U7986 ( .B1(n6293), .B2(n6292), .A(n6717), .ZN(n6294) );
  NAND2_X1 U7987 ( .A1(n6294), .A2(n9930), .ZN(n6295) );
  OAI211_X1 U7988 ( .C1(n6297), .C2(n9933), .A(n6296), .B(n6295), .ZN(P2_U3259) );
  INV_X1 U7989 ( .A(n6387), .ZN(n6299) );
  NAND2_X1 U7990 ( .A1(n6298), .A2(n9345), .ZN(n8888) );
  NAND2_X1 U7991 ( .A1(n6299), .A2(n8888), .ZN(n8782) );
  INV_X1 U7992 ( .A(n9344), .ZN(n6300) );
  NOR2_X1 U7993 ( .A1(n8926), .A2(n6300), .ZN(n6301) );
  AOI22_X1 U7994 ( .A1(n8782), .A2(n6301), .B1(n9828), .B2(n6007), .ZN(n9343)
         );
  NAND2_X1 U7995 ( .A1(n9814), .A2(n9154), .ZN(n9208) );
  OR2_X1 U7996 ( .A1(n9208), .A2(n9908), .ZN(n9063) );
  OAI21_X1 U7997 ( .B1(n9794), .B2(n9174), .A(n6302), .ZN(n6304) );
  INV_X1 U7998 ( .A(n9809), .ZN(n9838) );
  AOI22_X1 U7999 ( .A1(n9844), .A2(P1_REG2_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(n9838), .ZN(n6303) );
  OAI211_X1 U8000 ( .C1(n9844), .C2(n9343), .A(n6304), .B(n6303), .ZN(P1_U3291) );
  OAI21_X1 U8001 ( .B1(n6307), .B2(n6306), .A(n6305), .ZN(n6309) );
  NAND2_X1 U8002 ( .A1(n6307), .A2(n6306), .ZN(n6308) );
  NAND2_X1 U8003 ( .A1(n8941), .A2(n7568), .ZN(n6316) );
  OR2_X1 U8004 ( .A1(n6350), .A2(n6310), .ZN(n6314) );
  OR2_X1 U8005 ( .A1(n6067), .A2(n6311), .ZN(n6313) );
  OR2_X1 U8006 ( .A1(n6030), .A2(n4475), .ZN(n6312) );
  OR2_X1 U8007 ( .A1(n9876), .A2(n6055), .ZN(n6315) );
  NAND2_X1 U8008 ( .A1(n6316), .A2(n6315), .ZN(n6317) );
  XNOR2_X1 U8009 ( .A(n6317), .B(n5923), .ZN(n6334) );
  NAND2_X1 U8010 ( .A1(n8941), .A2(n7566), .ZN(n6319) );
  OR2_X1 U8011 ( .A1(n9876), .A2(n6049), .ZN(n6318) );
  NAND2_X1 U8012 ( .A1(n6319), .A2(n6318), .ZN(n6418) );
  NAND2_X1 U8013 ( .A1(n7555), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n6325) );
  OR2_X1 U8014 ( .A1(n4316), .A2(n6320), .ZN(n6324) );
  OAI21_X1 U8015 ( .B1(n6321), .B2(P1_REG3_REG_6__SCAN_IN), .A(n6342), .ZN(
        n6573) );
  OR2_X1 U8016 ( .A1(n5933), .A2(n6573), .ZN(n6323) );
  OR2_X1 U8017 ( .A1(n7598), .A2(n5949), .ZN(n6322) );
  NAND2_X1 U8018 ( .A1(n9827), .A2(n7592), .ZN(n6332) );
  OR2_X1 U8019 ( .A1(n6350), .A2(n6326), .ZN(n6330) );
  OR2_X1 U8020 ( .A1(n6067), .A2(n6327), .ZN(n6329) );
  OR2_X1 U8021 ( .A1(n6030), .A2(n9737), .ZN(n6328) );
  AND3_X2 U8022 ( .A1(n6330), .A2(n6329), .A3(n6328), .ZN(n6567) );
  OR2_X1 U8023 ( .A1(n6567), .A2(n6055), .ZN(n6331) );
  NAND2_X1 U8024 ( .A1(n6332), .A2(n6331), .ZN(n6333) );
  XNOR2_X1 U8025 ( .A(n6333), .B(n7564), .ZN(n6339) );
  INV_X1 U8026 ( .A(n6567), .ZN(n6509) );
  AOI22_X1 U8027 ( .A1(n9827), .A2(n7566), .B1(n6509), .B2(n7592), .ZN(n6338)
         );
  NAND2_X1 U8028 ( .A1(n6339), .A2(n6338), .ZN(n6560) );
  INV_X1 U8029 ( .A(n6334), .ZN(n6416) );
  INV_X1 U8030 ( .A(n6418), .ZN(n6335) );
  NAND2_X1 U8031 ( .A1(n6416), .A2(n6335), .ZN(n6336) );
  AND2_X1 U8032 ( .A1(n6560), .A2(n6336), .ZN(n6337) );
  OR2_X1 U8033 ( .A1(n6339), .A2(n6338), .ZN(n6558) );
  NAND2_X1 U8034 ( .A1(n7555), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n6348) );
  INV_X1 U8035 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n6340) );
  OR2_X1 U8036 ( .A1(n4316), .A2(n6340), .ZN(n6347) );
  AND2_X1 U8037 ( .A1(n6342), .A2(n6341), .ZN(n6343) );
  OR2_X1 U8038 ( .A1(n6343), .A2(n6361), .ZN(n6521) );
  OR2_X1 U8039 ( .A1(n5933), .A2(n6521), .ZN(n6346) );
  INV_X1 U8040 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n6344) );
  OR2_X1 U8041 ( .A1(n7598), .A2(n6344), .ZN(n6345) );
  NAND4_X1 U8042 ( .A1(n6348), .A2(n6347), .A3(n6346), .A4(n6345), .ZN(n8940)
         );
  NAND2_X1 U8043 ( .A1(n8940), .A2(n7566), .ZN(n6355) );
  AOI22_X1 U8044 ( .A1(n7338), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n9688), .B2(
        n6349), .ZN(n6353) );
  NAND2_X1 U8045 ( .A1(n6351), .A2(n8767), .ZN(n6352) );
  OR2_X1 U8046 ( .A1(n9892), .A2(n6049), .ZN(n6354) );
  NAND2_X1 U8047 ( .A1(n6355), .A2(n6354), .ZN(n6575) );
  NAND2_X1 U8048 ( .A1(n8940), .A2(n7592), .ZN(n6357) );
  OR2_X1 U8049 ( .A1(n9892), .A2(n6055), .ZN(n6356) );
  NAND2_X1 U8050 ( .A1(n6357), .A2(n6356), .ZN(n6358) );
  XNOR2_X1 U8051 ( .A(n6358), .B(n5923), .ZN(n6574) );
  XOR2_X1 U8052 ( .A(n6575), .B(n6574), .Z(n6359) );
  XNOR2_X1 U8053 ( .A(n6576), .B(n6359), .ZN(n6372) );
  INV_X1 U8054 ( .A(n9892), .ZN(n6524) );
  NAND2_X1 U8055 ( .A1(n7555), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n6366) );
  INV_X1 U8056 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6360) );
  OR2_X1 U8057 ( .A1(n4315), .A2(n6360), .ZN(n6365) );
  OR2_X1 U8058 ( .A1(n6361), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n6362) );
  NAND2_X1 U8059 ( .A1(n6591), .A2(n6362), .ZN(n6660) );
  OR2_X1 U8060 ( .A1(n5933), .A2(n6660), .ZN(n6364) );
  INV_X1 U8061 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n6661) );
  OR2_X1 U8062 ( .A1(n7598), .A2(n6661), .ZN(n6363) );
  INV_X1 U8063 ( .A(n9803), .ZN(n8939) );
  AOI21_X1 U8064 ( .B1(n4397), .B2(n8939), .A(n6367), .ZN(n6369) );
  NAND2_X1 U8065 ( .A1(n8621), .A2(n9827), .ZN(n6368) );
  OAI211_X1 U8066 ( .C1(n8668), .C2(n6521), .A(n6369), .B(n6368), .ZN(n6370)
         );
  AOI21_X1 U8067 ( .B1(n8670), .B2(n6524), .A(n6370), .ZN(n6371) );
  OAI21_X1 U8068 ( .B1(n6372), .B2(n8672), .A(n6371), .ZN(P1_U3211) );
  INV_X1 U8069 ( .A(n7337), .ZN(n6374) );
  OAI222_X1 U8070 ( .A1(n9376), .A2(n6373), .B1(n9373), .B2(n6374), .C1(n9154), 
        .C2(P1_U3084), .ZN(P1_U3334) );
  OAI222_X1 U8071 ( .A1(n8534), .A2(n6375), .B1(n7939), .B2(n6374), .C1(
        P2_U3152), .C2(n8325), .ZN(P2_U3339) );
  NOR2_X1 U8072 ( .A1(n5876), .A2(n9154), .ZN(n6376) );
  NAND2_X1 U8073 ( .A1(n9814), .A2(n6376), .ZN(n7271) );
  INV_X1 U8074 ( .A(n7271), .ZN(n9795) );
  NAND2_X1 U8075 ( .A1(n6007), .A2(n6388), .ZN(n6377) );
  NAND2_X1 U8076 ( .A1(n6380), .A2(n6379), .ZN(n6401) );
  NAND2_X1 U8077 ( .A1(n8944), .A2(n8891), .ZN(n6381) );
  NAND2_X1 U8078 ( .A1(n6401), .A2(n6381), .ZN(n6407) );
  AND2_X1 U8079 ( .A1(n6382), .A2(n6407), .ZN(n6383) );
  OR2_X1 U8080 ( .A1(n6403), .A2(n6383), .ZN(n9861) );
  AND2_X1 U8081 ( .A1(n6384), .A2(n8891), .ZN(n6385) );
  NOR2_X1 U8082 ( .A1(n6384), .A2(n8891), .ZN(n6404) );
  OR2_X1 U8083 ( .A1(n6385), .A2(n6404), .ZN(n9858) );
  AOI22_X1 U8084 ( .A1(n9174), .A2(n8891), .B1(P1_REG3_REG_2__SCAN_IN), .B2(
        n9838), .ZN(n6386) );
  OAI21_X1 U8085 ( .B1(n9063), .B2(n9858), .A(n6386), .ZN(n6398) );
  NAND2_X1 U8086 ( .A1(n6389), .A2(n6388), .ZN(n6390) );
  XNOR2_X1 U8087 ( .A(n8893), .B(n4638), .ZN(n6396) );
  NAND2_X1 U8088 ( .A1(n5859), .A2(n9154), .ZN(n6393) );
  MUX2_X1 U8089 ( .A(n6393), .B(n6392), .S(n5876), .Z(n9884) );
  INV_X1 U8090 ( .A(n9884), .ZN(n9671) );
  NAND2_X1 U8091 ( .A1(n9861), .A2(n9671), .ZN(n6395) );
  AOI22_X1 U8092 ( .A1(n9828), .A2(n8942), .B1(n6007), .B2(n9825), .ZN(n6394)
         );
  OAI211_X1 U8093 ( .C1(n9242), .C2(n6396), .A(n6395), .B(n6394), .ZN(n9859)
         );
  MUX2_X1 U8094 ( .A(n9859), .B(P1_REG2_REG_2__SCAN_IN), .S(n9844), .Z(n6397)
         );
  AOI211_X1 U8095 ( .C1(n9795), .C2(n9861), .A(n6398), .B(n6397), .ZN(n6399)
         );
  INV_X1 U8096 ( .A(n6399), .ZN(P1_U3289) );
  NAND2_X1 U8097 ( .A1(n8942), .A2(n9863), .ZN(n8833) );
  NAND2_X1 U8098 ( .A1(n6429), .A2(n8833), .ZN(n8780) );
  INV_X1 U8099 ( .A(n6401), .ZN(n6402) );
  XNOR2_X1 U8100 ( .A(n8780), .B(n6425), .ZN(n6411) );
  INV_X1 U8101 ( .A(n6411), .ZN(n9867) );
  NAND2_X1 U8102 ( .A1(n6404), .A2(n9863), .ZN(n6444) );
  OAI21_X1 U8103 ( .B1(n6404), .B2(n9863), .A(n6444), .ZN(n9864) );
  AOI22_X1 U8104 ( .A1(n9174), .A2(n7288), .B1(n6405), .B2(n9838), .ZN(n6406)
         );
  OAI21_X1 U8105 ( .B1(n9063), .B2(n9864), .A(n6406), .ZN(n6413) );
  OR2_X1 U8106 ( .A1(n8944), .A2(n6380), .ZN(n8889) );
  INV_X1 U8107 ( .A(n8780), .ZN(n6428) );
  XNOR2_X1 U8108 ( .A(n8837), .B(n6428), .ZN(n6409) );
  INV_X1 U8109 ( .A(n9826), .ZN(n6426) );
  OAI22_X1 U8110 ( .A1(n6379), .A2(n9802), .B1(n6426), .B2(n9800), .ZN(n6408)
         );
  AOI21_X1 U8111 ( .B1(n6409), .B2(n9823), .A(n6408), .ZN(n6410) );
  OAI21_X1 U8112 ( .B1(n6411), .B2(n9884), .A(n6410), .ZN(n9865) );
  MUX2_X1 U8113 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n9865), .S(n9814), .Z(n6412)
         );
  AOI211_X1 U8114 ( .C1(n9795), .C2(n9867), .A(n6413), .B(n6412), .ZN(n6414)
         );
  INV_X1 U8115 ( .A(n6414), .ZN(P1_U3288) );
  NAND2_X1 U8116 ( .A1(n6415), .A2(n6416), .ZN(n6559) );
  OAI21_X1 U8117 ( .B1(n6415), .B2(n6416), .A(n6559), .ZN(n6417) );
  NOR2_X1 U8118 ( .A1(n6417), .A2(n6418), .ZN(n6563) );
  AOI21_X1 U8119 ( .B1(n6418), .B2(n6417), .A(n6563), .ZN(n6424) );
  INV_X1 U8120 ( .A(n8668), .ZN(n8655) );
  AND2_X1 U8121 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n9714) );
  AOI21_X1 U8122 ( .B1(n8621), .B2(n9826), .A(n9714), .ZN(n6421) );
  NAND2_X1 U8123 ( .A1(n8670), .A2(n9835), .ZN(n6420) );
  NAND2_X1 U8124 ( .A1(n4397), .A2(n9827), .ZN(n6419) );
  NAND3_X1 U8125 ( .A1(n6421), .A2(n6420), .A3(n6419), .ZN(n6422) );
  AOI21_X1 U8126 ( .B1(n9837), .B2(n8655), .A(n6422), .ZN(n6423) );
  OAI21_X1 U8127 ( .B1(n6424), .B2(n8672), .A(n6423), .ZN(P1_U3225) );
  OAI22_X1 U8128 ( .A1(n6425), .A2(n6428), .B1(n8942), .B2(n7288), .ZN(n6438)
         );
  OR2_X1 U8129 ( .A1(n9826), .A2(n9869), .ZN(n9819) );
  NAND2_X1 U8130 ( .A1(n9826), .A2(n9869), .ZN(n8834) );
  NAND2_X1 U8131 ( .A1(n9819), .A2(n8834), .ZN(n8781) );
  AOI22_X1 U8132 ( .A1(n6438), .A2(n8781), .B1(n6426), .B2(n9869), .ZN(n9818)
         );
  OR2_X1 U8133 ( .A1(n8941), .A2(n9876), .ZN(n6513) );
  NAND2_X1 U8134 ( .A1(n8941), .A2(n9876), .ZN(n6511) );
  AOI22_X1 U8135 ( .A1(n9818), .A2(n9821), .B1(n8941), .B2(n9835), .ZN(n6427)
         );
  NAND2_X1 U8136 ( .A1(n9827), .A2(n6567), .ZN(n8842) );
  NAND2_X1 U8137 ( .A1(n8839), .A2(n8842), .ZN(n8786) );
  NAND2_X1 U8138 ( .A1(n6427), .A2(n8786), .ZN(n6508) );
  OAI21_X1 U8139 ( .B1(n6427), .B2(n8786), .A(n6508), .ZN(n9888) );
  INV_X1 U8140 ( .A(n9888), .ZN(n9885) );
  INV_X1 U8141 ( .A(n8940), .ZN(n6657) );
  NAND2_X1 U8142 ( .A1(n6511), .A2(n8834), .ZN(n6430) );
  NAND2_X1 U8143 ( .A1(n6430), .A2(n6513), .ZN(n8838) );
  INV_X1 U8144 ( .A(n8687), .ZN(n8686) );
  XNOR2_X1 U8145 ( .A(n8686), .B(n8786), .ZN(n6431) );
  OAI222_X1 U8146 ( .A1(n9800), .A2(n6657), .B1(n9802), .B2(n6432), .C1(n6431), 
        .C2(n9242), .ZN(n9887) );
  INV_X1 U8147 ( .A(n9887), .ZN(n6433) );
  MUX2_X1 U8148 ( .A(n5949), .B(n6433), .S(n9814), .Z(n6437) );
  INV_X1 U8149 ( .A(n9834), .ZN(n6434) );
  AOI21_X1 U8150 ( .B1(n6509), .B2(n6434), .A(n6522), .ZN(n9882) );
  OAI22_X1 U8151 ( .A1(n9808), .A2(n6567), .B1(n6573), .B2(n9809), .ZN(n6435)
         );
  AOI21_X1 U8152 ( .B1(n9882), .B2(n9794), .A(n6435), .ZN(n6436) );
  OAI211_X1 U8153 ( .C1(n9885), .C2(n9256), .A(n6437), .B(n6436), .ZN(P1_U3285) );
  XNOR2_X1 U8154 ( .A(n6438), .B(n8781), .ZN(n9873) );
  INV_X1 U8155 ( .A(n9873), .ZN(n6451) );
  XNOR2_X1 U8156 ( .A(n6510), .B(n8781), .ZN(n6441) );
  NAND2_X1 U8157 ( .A1(n9873), .A2(n9671), .ZN(n6440) );
  AOI22_X1 U8158 ( .A1(n9828), .A2(n8941), .B1(n8942), .B2(n9825), .ZN(n6439)
         );
  OAI211_X1 U8159 ( .C1(n9242), .C2(n6441), .A(n6440), .B(n6439), .ZN(n9871)
         );
  NAND2_X1 U8160 ( .A1(n9871), .A2(n9814), .ZN(n6450) );
  OAI22_X1 U8161 ( .A1(n9814), .A2(n6443), .B1(n6442), .B2(n9809), .ZN(n6447)
         );
  NAND2_X1 U8162 ( .A1(n6444), .A2(n6448), .ZN(n6445) );
  NAND2_X1 U8163 ( .A1(n9831), .A2(n6445), .ZN(n9870) );
  NOR2_X1 U8164 ( .A1(n9063), .A2(n9870), .ZN(n6446) );
  AOI211_X1 U8165 ( .C1(n9174), .C2(n6448), .A(n6447), .B(n6446), .ZN(n6449)
         );
  OAI211_X1 U8166 ( .C1(n6451), .C2(n7271), .A(n6450), .B(n6449), .ZN(P1_U3287) );
  OR2_X1 U8167 ( .A1(n6452), .A2(n6453), .ZN(n6616) );
  INV_X1 U8168 ( .A(n6616), .ZN(n6454) );
  AOI22_X1 U8169 ( .A1(n6454), .A2(n6615), .B1(n6457), .B2(n6452), .ZN(n9987)
         );
  NAND2_X1 U8170 ( .A1(n6688), .A2(n6455), .ZN(n6456) );
  NAND2_X1 U8171 ( .A1(n6456), .A2(n7646), .ZN(n6458) );
  XNOR2_X1 U8172 ( .A(n6458), .B(n6457), .ZN(n6461) );
  OAI22_X1 U8173 ( .A1(n6460), .A2(n8305), .B1(n6459), .B2(n8307), .ZN(n6554)
         );
  AOI21_X1 U8174 ( .B1(n6461), .B2(n8395), .A(n6554), .ZN(n9990) );
  MUX2_X1 U8175 ( .A(n6462), .B(n9990), .S(n9953), .Z(n6467) );
  INV_X1 U8176 ( .A(n6692), .ZN(n6463) );
  OAI21_X1 U8177 ( .B1(n6463), .B2(n9988), .A(n6623), .ZN(n9989) );
  INV_X1 U8178 ( .A(n6464), .ZN(n6557) );
  OAI22_X1 U8179 ( .A1(n9989), .A2(n8167), .B1(n6557), .B2(n8356), .ZN(n6465)
         );
  AOI21_X1 U8180 ( .B1(n8359), .B2(n6472), .A(n6465), .ZN(n6466) );
  OAI211_X1 U8181 ( .C1(n9987), .C2(n8365), .A(n6467), .B(n6466), .ZN(P2_U3290) );
  NAND2_X1 U8182 ( .A1(n8063), .A2(n7635), .ZN(n6470) );
  INV_X1 U8183 ( .A(n6470), .ZN(n6469) );
  XNOR2_X1 U8184 ( .A(n7921), .B(n6625), .ZN(n6471) );
  INV_X1 U8185 ( .A(n6471), .ZN(n6468) );
  NAND2_X1 U8186 ( .A1(n6469), .A2(n6468), .ZN(n6481) );
  INV_X1 U8187 ( .A(n6481), .ZN(n6477) );
  XNOR2_X1 U8188 ( .A(n6471), .B(n6470), .ZN(n6604) );
  INV_X1 U8189 ( .A(n6604), .ZN(n6475) );
  XNOR2_X1 U8190 ( .A(n7926), .B(n6472), .ZN(n6478) );
  INV_X1 U8191 ( .A(n6478), .ZN(n6474) );
  AND2_X1 U8192 ( .A1(n8064), .A2(n7635), .ZN(n6479) );
  INV_X1 U8193 ( .A(n6479), .ZN(n6473) );
  NAND2_X1 U8194 ( .A1(n6474), .A2(n6473), .ZN(n6602) );
  AND2_X1 U8195 ( .A1(n6475), .A2(n6602), .ZN(n6476) );
  NOR2_X1 U8196 ( .A1(n6477), .A2(n6476), .ZN(n6488) );
  OR2_X1 U8197 ( .A1(n6545), .A2(n6488), .ZN(n6490) );
  NAND2_X1 U8198 ( .A1(n6479), .A2(n6478), .ZN(n6480) );
  AND2_X1 U8199 ( .A1(n6480), .A2(n6602), .ZN(n6550) );
  AND2_X1 U8200 ( .A1(n6550), .A2(n6481), .ZN(n6486) );
  INV_X1 U8201 ( .A(n6482), .ZN(n6485) );
  INV_X1 U8202 ( .A(n6483), .ZN(n6484) );
  NAND2_X1 U8203 ( .A1(n6485), .A2(n6484), .ZN(n6547) );
  AND2_X1 U8204 ( .A1(n6486), .A2(n6547), .ZN(n6487) );
  OR2_X1 U8205 ( .A1(n6488), .A2(n6487), .ZN(n6489) );
  XNOR2_X1 U8206 ( .A(n6814), .B(n7926), .ZN(n6636) );
  NAND2_X1 U8207 ( .A1(n8062), .A2(n7635), .ZN(n6634) );
  XNOR2_X1 U8208 ( .A(n6636), .B(n6634), .ZN(n6638) );
  XNOR2_X1 U8209 ( .A(n6639), .B(n6638), .ZN(n6494) );
  AOI22_X1 U8210 ( .A1(n6608), .A2(n8061), .B1(n8033), .B2(n6813), .ZN(n6493)
         );
  OAI22_X1 U8211 ( .A1(n8026), .A2(n9995), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9557), .ZN(n6491) );
  AOI21_X1 U8212 ( .B1(n6609), .B2(n8063), .A(n6491), .ZN(n6492) );
  OAI211_X1 U8213 ( .C1(n6494), .C2(n8036), .A(n6493), .B(n6492), .ZN(P2_U3223) );
  INV_X1 U8214 ( .A(n7350), .ZN(n6506) );
  OAI222_X1 U8215 ( .A1(n9373), .A2(n6506), .B1(P1_U3084), .B2(n5844), .C1(
        n7351), .C2(n9376), .ZN(P1_U3333) );
  INV_X1 U8216 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n6501) );
  INV_X1 U8217 ( .A(n10006), .ZN(n8487) );
  AOI22_X1 U8218 ( .A1(n6496), .A2(n8499), .B1(n8498), .B2(n6495), .ZN(n6497)
         );
  OAI211_X1 U8219 ( .C1(n6499), .C2(n8487), .A(n6498), .B(n6497), .ZN(n6504)
         );
  NAND2_X1 U8220 ( .A1(n6504), .A2(n10019), .ZN(n6500) );
  OAI21_X1 U8221 ( .B1(n10019), .B2(n6501), .A(n6500), .ZN(P2_U3460) );
  AND2_X2 U8222 ( .A1(n6503), .A2(n6502), .ZN(n10033) );
  NAND2_X1 U8223 ( .A1(n6504), .A2(n10033), .ZN(n6505) );
  OAI21_X1 U8224 ( .B1(n10033), .B2(n5681), .A(n6505), .ZN(P2_U3523) );
  OAI222_X1 U8225 ( .A1(n8534), .A2(n6507), .B1(n7939), .B2(n6506), .C1(n7818), 
        .C2(P2_U3152), .ZN(P2_U3338) );
  NAND2_X1 U8226 ( .A1(n8940), .A2(n9892), .ZN(n8845) );
  NAND2_X1 U8227 ( .A1(n8703), .A2(n8845), .ZN(n8784) );
  XNOR2_X1 U8228 ( .A(n6658), .B(n8784), .ZN(n9894) );
  INV_X1 U8229 ( .A(n9894), .ZN(n6530) );
  NAND2_X1 U8230 ( .A1(n8842), .A2(n6511), .ZN(n6512) );
  AND2_X1 U8231 ( .A1(n6513), .A2(n9819), .ZN(n6514) );
  NAND2_X1 U8232 ( .A1(n6514), .A2(n8839), .ZN(n8844) );
  INV_X1 U8233 ( .A(n8836), .ZN(n6515) );
  AND2_X1 U8234 ( .A1(n8844), .A2(n6515), .ZN(n6517) );
  INV_X1 U8235 ( .A(n6517), .ZN(n8898) );
  NAND2_X1 U8236 ( .A1(n8898), .A2(n8784), .ZN(n6518) );
  INV_X1 U8237 ( .A(n8784), .ZN(n6516) );
  OAI21_X1 U8238 ( .B1(n6519), .B2(n6518), .A(n6935), .ZN(n6520) );
  AOI222_X1 U8239 ( .A1(n9823), .A2(n6520), .B1(n8939), .B2(n9828), .C1(n9827), 
        .C2(n9825), .ZN(n9891) );
  OAI21_X1 U8240 ( .B1(n6521), .B2(n9809), .A(n9891), .ZN(n6528) );
  OAI211_X1 U8241 ( .C1(n6522), .C2(n9892), .A(n9881), .B(n6662), .ZN(n9890)
         );
  NOR2_X1 U8242 ( .A1(n6523), .A2(n9840), .ZN(n9228) );
  INV_X1 U8243 ( .A(n9228), .ZN(n6526) );
  AOI22_X1 U8244 ( .A1(n9174), .A2(n6524), .B1(n9844), .B2(
        P1_REG2_REG_7__SCAN_IN), .ZN(n6525) );
  OAI21_X1 U8245 ( .B1(n9890), .B2(n6526), .A(n6525), .ZN(n6527) );
  AOI21_X1 U8246 ( .B1(n6528), .B2(n9814), .A(n6527), .ZN(n6529) );
  OAI21_X1 U8247 ( .B1(n6530), .B2(n9256), .A(n6529), .ZN(P1_U3284) );
  INV_X1 U8248 ( .A(n9785), .ZN(n9759) );
  NAND2_X1 U8249 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_U3084), .ZN(n6536) );
  OAI21_X1 U8250 ( .B1(n6533), .B2(n6532), .A(n6531), .ZN(n6534) );
  NAND2_X1 U8251 ( .A1(n9781), .A2(n6534), .ZN(n6535) );
  OAI211_X1 U8252 ( .C1(n9783), .C2(n7074), .A(n6536), .B(n6535), .ZN(n6541)
         );
  INV_X1 U8253 ( .A(n9751), .ZN(n9774) );
  AOI211_X1 U8254 ( .C1(n6539), .C2(n6538), .A(n6537), .B(n9774), .ZN(n6540)
         );
  AOI211_X1 U8255 ( .C1(P1_ADDR_REG_12__SCAN_IN), .C2(n9759), .A(n6541), .B(
        n6540), .ZN(n6542) );
  INV_X1 U8256 ( .A(n6542), .ZN(P1_U3253) );
  INV_X1 U8257 ( .A(n7362), .ZN(n6633) );
  OAI222_X1 U8258 ( .A1(n8534), .A2(n6544), .B1(n7939), .B2(n6633), .C1(n6543), 
        .C2(P2_U3152), .ZN(P2_U3337) );
  OR2_X1 U8259 ( .A1(n6546), .A2(n6545), .ZN(n6548) );
  AND2_X1 U8260 ( .A1(n6548), .A2(n6547), .ZN(n6549) );
  NAND2_X1 U8261 ( .A1(n6549), .A2(n6550), .ZN(n6603) );
  OAI21_X1 U8262 ( .B1(n6550), .B2(n6549), .A(n6603), .ZN(n6551) );
  NAND2_X1 U8263 ( .A1(n6551), .A2(n8038), .ZN(n6556) );
  NOR2_X1 U8264 ( .A1(n8026), .A2(n9988), .ZN(n6552) );
  AOI211_X1 U8265 ( .C1(n8043), .C2(n6554), .A(n6553), .B(n6552), .ZN(n6555)
         );
  OAI211_X1 U8266 ( .C1(n8045), .C2(n6557), .A(n6556), .B(n6555), .ZN(P2_U3241) );
  INV_X1 U8267 ( .A(n6558), .ZN(n6566) );
  INV_X1 U8268 ( .A(n6559), .ZN(n6562) );
  INV_X1 U8269 ( .A(n6560), .ZN(n6561) );
  OAI22_X1 U8270 ( .A1(n6563), .A2(n6562), .B1(n6566), .B2(n6561), .ZN(n6564)
         );
  OAI211_X1 U8271 ( .C1(n6566), .C2(n6565), .A(n6564), .B(n8597), .ZN(n6572)
         );
  NOR2_X1 U8272 ( .A1(n9906), .A2(n6567), .ZN(n9880) );
  INV_X1 U8273 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6568) );
  NOR2_X1 U8274 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6568), .ZN(n9735) );
  AOI21_X1 U8275 ( .B1(n8621), .B2(n8941), .A(n9735), .ZN(n6569) );
  OAI21_X1 U8276 ( .B1(n8599), .B2(n6657), .A(n6569), .ZN(n6570) );
  AOI21_X1 U8277 ( .B1(n8612), .B2(n9880), .A(n6570), .ZN(n6571) );
  OAI211_X1 U8278 ( .C1(n8668), .C2(n6573), .A(n6572), .B(n6571), .ZN(P1_U3237) );
  OAI21_X1 U8279 ( .B1(n6576), .B2(n6575), .A(n6574), .ZN(n6578) );
  NAND2_X1 U8280 ( .A1(n6576), .A2(n6575), .ZN(n6577) );
  NAND2_X1 U8281 ( .A1(n6578), .A2(n6577), .ZN(n6757) );
  NAND2_X1 U8282 ( .A1(n6579), .A2(n8767), .ZN(n6582) );
  AOI22_X1 U8283 ( .A1(n7338), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n9688), .B2(
        n6580), .ZN(n6581) );
  NAND2_X1 U8284 ( .A1(n6582), .A2(n6581), .ZN(n6666) );
  NAND2_X1 U8285 ( .A1(n6666), .A2(n7579), .ZN(n6583) );
  OAI21_X1 U8286 ( .B1(n9803), .B2(n6049), .A(n6583), .ZN(n6584) );
  XNOR2_X1 U8287 ( .A(n6584), .B(n7564), .ZN(n6758) );
  OR2_X1 U8288 ( .A1(n9803), .A2(n7590), .ZN(n6586) );
  NAND2_X1 U8289 ( .A1(n6666), .A2(n7592), .ZN(n6585) );
  AND2_X1 U8290 ( .A1(n6586), .A2(n6585), .ZN(n6755) );
  INV_X1 U8291 ( .A(n6755), .ZN(n6759) );
  XNOR2_X1 U8292 ( .A(n6758), .B(n6759), .ZN(n6587) );
  XNOR2_X1 U8293 ( .A(n6757), .B(n6587), .ZN(n6601) );
  NOR2_X1 U8294 ( .A1(n6931), .A2(n9906), .ZN(n9903) );
  INV_X1 U8295 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n6588) );
  NOR2_X1 U8296 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6588), .ZN(n9749) );
  AOI21_X1 U8297 ( .B1(n8621), .B2(n8940), .A(n9749), .ZN(n6598) );
  NAND2_X1 U8298 ( .A1(n7555), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n6596) );
  INV_X1 U8299 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n6589) );
  OR2_X1 U8300 ( .A1(n4315), .A2(n6589), .ZN(n6595) );
  NAND2_X1 U8301 ( .A1(n6591), .A2(n6590), .ZN(n6592) );
  NAND2_X1 U8302 ( .A1(n6767), .A2(n6592), .ZN(n9810) );
  OR2_X1 U8303 ( .A1(n5933), .A2(n9810), .ZN(n6594) );
  INV_X1 U8304 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n9811) );
  OR2_X1 U8305 ( .A1(n7598), .A2(n9811), .ZN(n6593) );
  NAND2_X1 U8306 ( .A1(n4397), .A2(n8938), .ZN(n6597) );
  OAI211_X1 U8307 ( .C1(n8668), .C2(n6660), .A(n6598), .B(n6597), .ZN(n6599)
         );
  AOI21_X1 U8308 ( .B1(n8612), .B2(n9903), .A(n6599), .ZN(n6600) );
  OAI21_X1 U8309 ( .B1(n6601), .B2(n8672), .A(n6600), .ZN(P1_U3219) );
  NAND2_X1 U8310 ( .A1(n6603), .A2(n6602), .ZN(n6605) );
  XNOR2_X1 U8311 ( .A(n6605), .B(n6604), .ZN(n6612) );
  NOR2_X1 U8312 ( .A1(n8026), .A2(n6673), .ZN(n6606) );
  AOI211_X1 U8313 ( .C1(n8033), .C2(n6670), .A(n6607), .B(n6606), .ZN(n6611)
         );
  AOI22_X1 U8314 ( .A1(n6609), .A2(n8064), .B1(n6608), .B2(n8062), .ZN(n6610)
         );
  OAI211_X1 U8315 ( .C1(n6612), .C2(n8036), .A(n6611), .B(n6610), .ZN(P2_U3215) );
  INV_X1 U8316 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n6630) );
  AND2_X1 U8317 ( .A1(n6613), .A2(n6614), .ZN(n6618) );
  NAND3_X1 U8318 ( .A1(n6616), .A2(n7678), .A3(n6615), .ZN(n6617) );
  NAND2_X1 U8319 ( .A1(n6618), .A2(n6617), .ZN(n6677) );
  INV_X1 U8320 ( .A(n6677), .ZN(n6628) );
  OR2_X1 U8321 ( .A1(n6619), .A2(n7825), .ZN(n6817) );
  NAND2_X1 U8322 ( .A1(n6619), .A2(n7825), .ZN(n6620) );
  NAND3_X1 U8323 ( .A1(n6817), .A2(n8395), .A3(n6620), .ZN(n6622) );
  AOI22_X1 U8324 ( .A1(n8390), .A2(n8064), .B1(n8062), .B2(n8392), .ZN(n6621)
         );
  NAND2_X1 U8325 ( .A1(n6622), .A2(n6621), .ZN(n6674) );
  INV_X1 U8326 ( .A(n6674), .ZN(n6627) );
  AND2_X1 U8327 ( .A1(n6623), .A2(n6625), .ZN(n6624) );
  NOR2_X1 U8328 ( .A1(n6810), .A2(n6624), .ZN(n6671) );
  AOI22_X1 U8329 ( .A1(n6671), .A2(n8499), .B1(n8498), .B2(n6625), .ZN(n6626)
         );
  OAI211_X1 U8330 ( .C1(n8503), .C2(n6628), .A(n6627), .B(n6626), .ZN(n6631)
         );
  NAND2_X1 U8331 ( .A1(n6631), .A2(n10019), .ZN(n6629) );
  OAI21_X1 U8332 ( .B1(n10019), .B2(n6630), .A(n6629), .ZN(P2_U3472) );
  NAND2_X1 U8333 ( .A1(n6631), .A2(n10033), .ZN(n6632) );
  OAI21_X1 U8334 ( .B1(n10033), .B2(n5774), .A(n6632), .ZN(P2_U3527) );
  INV_X1 U8335 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7363) );
  OAI222_X1 U8336 ( .A1(n9373), .A2(n6633), .B1(P1_U3084), .B2(n5842), .C1(
        n7363), .C2(n9376), .ZN(P1_U3332) );
  INV_X1 U8337 ( .A(n6634), .ZN(n6635) );
  AND2_X1 U8338 ( .A1(n6636), .A2(n6635), .ZN(n6637) );
  XNOR2_X1 U8339 ( .A(n6975), .B(n7921), .ZN(n6640) );
  NAND2_X1 U8340 ( .A1(n8061), .A2(n7635), .ZN(n6641) );
  NAND2_X1 U8341 ( .A1(n6640), .A2(n6641), .ZN(n6679) );
  INV_X1 U8342 ( .A(n6640), .ZN(n6643) );
  INV_X1 U8343 ( .A(n6641), .ZN(n6642) );
  NAND2_X1 U8344 ( .A1(n6643), .A2(n6642), .ZN(n6644) );
  AND2_X1 U8345 ( .A1(n6679), .A2(n6644), .ZN(n6645) );
  NAND2_X1 U8346 ( .A1(n6646), .A2(n6645), .ZN(n6680) );
  OAI21_X1 U8347 ( .B1(n6646), .B2(n6645), .A(n6680), .ZN(n6647) );
  NAND2_X1 U8348 ( .A1(n6647), .A2(n8038), .ZN(n6651) );
  AND2_X1 U8349 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3152), .ZN(n8084) );
  OAI22_X1 U8350 ( .A1(n6648), .A2(n8030), .B1(n8029), .B2(n6801), .ZN(n6649)
         );
  AOI211_X1 U8351 ( .C1(n6789), .C2(n8033), .A(n8084), .B(n6649), .ZN(n6650)
         );
  OAI211_X1 U8352 ( .C1(n5056), .C2(n8026), .A(n6651), .B(n6650), .ZN(P2_U3233) );
  NAND2_X1 U8353 ( .A1(n9803), .A2(n6666), .ZN(n8706) );
  NAND2_X1 U8354 ( .A1(n6931), .A2(n8939), .ZN(n9796) );
  NAND2_X1 U8355 ( .A1(n8706), .A2(n9796), .ZN(n8785) );
  INV_X1 U8356 ( .A(n8785), .ZN(n6652) );
  AOI21_X1 U8357 ( .B1(n6935), .B2(n8703), .A(n6652), .ZN(n6656) );
  AND2_X1 U8358 ( .A1(n8706), .A2(n8703), .ZN(n8830) );
  NAND3_X1 U8359 ( .A1(n6935), .A2(n8830), .A3(n9796), .ZN(n6653) );
  NAND2_X1 U8360 ( .A1(n6653), .A2(n9823), .ZN(n6655) );
  AOI22_X1 U8361 ( .A1(n8938), .A2(n9828), .B1(n9825), .B2(n8940), .ZN(n6654)
         );
  OAI21_X1 U8362 ( .B1(n6656), .B2(n6655), .A(n6654), .ZN(n9901) );
  INV_X1 U8363 ( .A(n9901), .ZN(n6669) );
  NOR2_X1 U8364 ( .A1(n6659), .A2(n8785), .ZN(n9899) );
  INV_X1 U8365 ( .A(n6930), .ZN(n9898) );
  OR3_X1 U8366 ( .A1(n9899), .A2(n9898), .A3(n9256), .ZN(n6668) );
  OAI22_X1 U8367 ( .A1(n9814), .A2(n6661), .B1(n6660), .B2(n9809), .ZN(n6665)
         );
  INV_X1 U8368 ( .A(n6662), .ZN(n6663) );
  OAI21_X1 U8369 ( .B1(n6663), .B2(n6931), .A(n9790), .ZN(n9900) );
  NOR2_X1 U8370 ( .A1(n9900), .A2(n9063), .ZN(n6664) );
  AOI211_X1 U8371 ( .C1(n9174), .C2(n6666), .A(n6665), .B(n6664), .ZN(n6667)
         );
  OAI211_X1 U8372 ( .C1(n9844), .C2(n6669), .A(n6668), .B(n6667), .ZN(P1_U3283) );
  AOI22_X1 U8373 ( .A1(n6671), .A2(n8402), .B1(n6670), .B2(n9944), .ZN(n6672)
         );
  OAI21_X1 U8374 ( .B1(n6673), .B2(n8406), .A(n6672), .ZN(n6676) );
  MUX2_X1 U8375 ( .A(n6674), .B(P2_REG2_REG_7__SCAN_IN), .S(n8368), .Z(n6675)
         );
  AOI211_X1 U8376 ( .C1(n8409), .C2(n6677), .A(n6676), .B(n6675), .ZN(n6678)
         );
  INV_X1 U8377 ( .A(n6678), .ZN(P2_U3289) );
  NAND2_X1 U8378 ( .A1(n6680), .A2(n6679), .ZN(n6889) );
  XNOR2_X1 U8379 ( .A(n5308), .B(n7921), .ZN(n6794) );
  NAND2_X1 U8380 ( .A1(n8060), .A2(n7635), .ZN(n6795) );
  XNOR2_X1 U8381 ( .A(n6794), .B(n6795), .ZN(n6891) );
  XNOR2_X1 U8382 ( .A(n6889), .B(n6891), .ZN(n6686) );
  INV_X1 U8383 ( .A(n6742), .ZN(n6681) );
  OAI22_X1 U8384 ( .A1(n8045), .A2(n6681), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9540), .ZN(n6684) );
  OAI22_X1 U8385 ( .A1(n6682), .A2(n8030), .B1(n8029), .B2(n6924), .ZN(n6683)
         );
  AOI211_X1 U8386 ( .C1(n8047), .C2(n5308), .A(n6684), .B(n6683), .ZN(n6685)
         );
  OAI21_X1 U8387 ( .B1(n6686), .B2(n8036), .A(n6685), .ZN(P2_U3219) );
  INV_X1 U8388 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6696) );
  XOR2_X1 U8389 ( .A(n6687), .B(n7824), .Z(n9940) );
  NAND2_X1 U8390 ( .A1(n6688), .A2(n7672), .ZN(n6689) );
  XNOR2_X1 U8391 ( .A(n6689), .B(n7824), .ZN(n6690) );
  AOI222_X1 U8392 ( .A1(n8395), .A2(n6690), .B1(n8064), .B2(n8392), .C1(n8067), 
        .C2(n8390), .ZN(n9948) );
  INV_X1 U8393 ( .A(n8499), .ZN(n10010) );
  AOI21_X1 U8394 ( .B1(n6691), .B2(n5264), .A(n10010), .ZN(n6693) );
  AND2_X1 U8395 ( .A1(n6693), .A2(n6692), .ZN(n9941) );
  AOI21_X1 U8396 ( .B1(n8498), .B2(n5264), .A(n9941), .ZN(n6694) );
  OAI211_X1 U8397 ( .C1(n8503), .C2(n9940), .A(n9948), .B(n6694), .ZN(n6697)
         );
  NAND2_X1 U8398 ( .A1(n6697), .A2(n10033), .ZN(n6695) );
  OAI21_X1 U8399 ( .B1(n10033), .B2(n6696), .A(n6695), .ZN(P2_U3525) );
  INV_X1 U8400 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n6699) );
  NAND2_X1 U8401 ( .A1(n6697), .A2(n10019), .ZN(n6698) );
  OAI21_X1 U8402 ( .B1(n10019), .B2(n6699), .A(n6698), .ZN(P2_U3466) );
  INV_X1 U8403 ( .A(n6700), .ZN(n6701) );
  OAI21_X1 U8404 ( .B1(n7169), .B2(P1_REG1_REG_13__SCAN_IN), .A(n6701), .ZN(
        n6703) );
  INV_X1 U8405 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n7176) );
  MUX2_X1 U8406 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n7176), .S(n7210), .Z(n6702)
         );
  NAND2_X1 U8407 ( .A1(n6702), .A2(n6703), .ZN(n6969) );
  OAI21_X1 U8408 ( .B1(n6703), .B2(n6702), .A(n6969), .ZN(n6704) );
  NAND2_X1 U8409 ( .A1(n6704), .A2(n9781), .ZN(n6706) );
  NOR2_X1 U8410 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7177), .ZN(n7250) );
  INV_X1 U8411 ( .A(n7250), .ZN(n6705) );
  OAI211_X1 U8412 ( .C1(n9783), .C2(n6962), .A(n6706), .B(n6705), .ZN(n6711)
         );
  XNOR2_X1 U8413 ( .A(n6962), .B(n6963), .ZN(n6709) );
  INV_X1 U8414 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n6708) );
  NOR2_X1 U8415 ( .A1(n6708), .A2(n6709), .ZN(n6964) );
  AOI211_X1 U8416 ( .C1(n6709), .C2(n6708), .A(n6964), .B(n9774), .ZN(n6710)
         );
  AOI211_X1 U8417 ( .C1(P1_ADDR_REG_14__SCAN_IN), .C2(n9759), .A(n6711), .B(
        n6710), .ZN(n6712) );
  INV_X1 U8418 ( .A(n6712), .ZN(P1_U3255) );
  AOI21_X1 U8419 ( .B1(n6715), .B2(n6714), .A(n6713), .ZN(n6875) );
  XNOR2_X1 U8420 ( .A(n6875), .B(n6876), .ZN(n6716) );
  NOR2_X1 U8421 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n6716), .ZN(n6877) );
  AOI21_X1 U8422 ( .B1(n6716), .B2(P2_REG2_REG_15__SCAN_IN), .A(n6877), .ZN(
        n6727) );
  OAI21_X1 U8423 ( .B1(n6718), .B2(P2_REG1_REG_14__SCAN_IN), .A(n6717), .ZN(
        n6869) );
  XNOR2_X1 U8424 ( .A(n6869), .B(n6870), .ZN(n6719) );
  INV_X1 U8425 ( .A(n6719), .ZN(n6722) );
  INV_X1 U8426 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n6720) );
  NOR2_X1 U8427 ( .A1(n6720), .A2(n6719), .ZN(n6871) );
  INV_X1 U8428 ( .A(n6871), .ZN(n6721) );
  OAI211_X1 U8429 ( .C1(n6722), .C2(P2_REG1_REG_15__SCAN_IN), .A(n9930), .B(
        n6721), .ZN(n6726) );
  NOR2_X1 U8430 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7108), .ZN(n6724) );
  NOR2_X1 U8431 ( .A1(n9932), .A2(n6870), .ZN(n6723) );
  AOI211_X1 U8432 ( .C1(P2_ADDR_REG_15__SCAN_IN), .C2(n9935), .A(n6724), .B(
        n6723), .ZN(n6725) );
  OAI211_X1 U8433 ( .C1(n6727), .C2(n9933), .A(n6726), .B(n6725), .ZN(P2_U3260) );
  OAI21_X1 U8434 ( .B1(n6729), .B2(n6734), .A(n6728), .ZN(n6740) );
  AOI22_X1 U8435 ( .A1(n8390), .A2(n8061), .B1(n8059), .B2(n8392), .ZN(n6739)
         );
  OR2_X1 U8436 ( .A1(n6619), .A2(n6730), .ZN(n6732) );
  AND2_X1 U8437 ( .A1(n6732), .A2(n6731), .ZN(n6779) );
  NAND2_X1 U8438 ( .A1(n6779), .A2(n7828), .ZN(n6733) );
  NAND2_X1 U8439 ( .A1(n6733), .A2(n7696), .ZN(n6735) );
  INV_X1 U8440 ( .A(n6735), .ZN(n6737) );
  OR2_X1 U8441 ( .A1(n6735), .A2(n6734), .ZN(n6736) );
  OAI211_X1 U8442 ( .C1(n6737), .C2(n5491), .A(n8395), .B(n6736), .ZN(n6738)
         );
  OAI211_X1 U8443 ( .C1(n6740), .C2(n8379), .A(n6739), .B(n6738), .ZN(n10003)
         );
  INV_X1 U8444 ( .A(n10003), .ZN(n6747) );
  INV_X1 U8445 ( .A(n6740), .ZN(n10005) );
  INV_X1 U8446 ( .A(n8388), .ZN(n7040) );
  AND2_X1 U8447 ( .A1(n6787), .A2(n5308), .ZN(n6741) );
  OR2_X1 U8448 ( .A1(n6741), .A2(n6952), .ZN(n10002) );
  AOI22_X1 U8449 ( .A1(n8368), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n6742), .B2(
        n9944), .ZN(n6744) );
  NAND2_X1 U8450 ( .A1(n8359), .A2(n5308), .ZN(n6743) );
  OAI211_X1 U8451 ( .C1(n10002), .C2(n8167), .A(n6744), .B(n6743), .ZN(n6745)
         );
  AOI21_X1 U8452 ( .B1(n10005), .B2(n7040), .A(n6745), .ZN(n6746) );
  OAI21_X1 U8453 ( .B1(n6747), .B2(n8368), .A(n6746), .ZN(P2_U3286) );
  INV_X1 U8454 ( .A(n7291), .ZN(n7864) );
  OAI222_X1 U8455 ( .A1(n9376), .A2(n7292), .B1(n9373), .B2(n7864), .C1(n5859), 
        .C2(P1_U3084), .ZN(P1_U3331) );
  NAND2_X1 U8456 ( .A1(n6748), .A2(n8767), .ZN(n6750) );
  AOI22_X1 U8457 ( .A1(n7338), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n9688), .B2(
        n9757), .ZN(n6749) );
  OAI22_X1 U8458 ( .A1(n9907), .A2(n6055), .B1(n6936), .B2(n6049), .ZN(n6751)
         );
  XNOR2_X1 U8459 ( .A(n6751), .B(n5923), .ZN(n6753) );
  OAI22_X1 U8460 ( .A1(n9907), .A2(n6049), .B1(n6936), .B2(n7590), .ZN(n6752)
         );
  OR2_X1 U8461 ( .A1(n6753), .A2(n6752), .ZN(n6827) );
  NAND2_X1 U8462 ( .A1(n6753), .A2(n6752), .ZN(n6754) );
  NAND2_X1 U8463 ( .A1(n6827), .A2(n6754), .ZN(n6765) );
  NAND2_X1 U8464 ( .A1(n6758), .A2(n6755), .ZN(n6756) );
  INV_X1 U8465 ( .A(n6758), .ZN(n6760) );
  NAND2_X1 U8466 ( .A1(n6760), .A2(n6759), .ZN(n6761) );
  INV_X1 U8467 ( .A(n6765), .ZN(n6762) );
  INV_X1 U8468 ( .A(n6828), .ZN(n6763) );
  AOI21_X1 U8469 ( .B1(n6765), .B2(n6764), .A(n6763), .ZN(n6778) );
  NAND2_X1 U8470 ( .A1(n7555), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n6773) );
  OR2_X1 U8471 ( .A1(n4316), .A2(n6766), .ZN(n6772) );
  NAND2_X1 U8472 ( .A1(n6767), .A2(n6843), .ZN(n6768) );
  NAND2_X1 U8473 ( .A1(n6845), .A2(n6768), .ZN(n6942) );
  OR2_X1 U8474 ( .A1(n5933), .A2(n6942), .ZN(n6771) );
  INV_X1 U8475 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n6769) );
  OR2_X1 U8476 ( .A1(n7598), .A2(n6769), .ZN(n6770) );
  INV_X1 U8477 ( .A(n9801), .ZN(n8937) );
  AND2_X1 U8478 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n9767) );
  NOR2_X1 U8479 ( .A1(n8663), .A2(n9803), .ZN(n6774) );
  AOI211_X1 U8480 ( .C1(n4397), .C2(n8937), .A(n9767), .B(n6774), .ZN(n6775)
         );
  OAI21_X1 U8481 ( .B1(n8668), .B2(n9810), .A(n6775), .ZN(n6776) );
  AOI21_X1 U8482 ( .B1(n8670), .B2(n6941), .A(n6776), .ZN(n6777) );
  OAI21_X1 U8483 ( .B1(n6778), .B2(n8672), .A(n6777), .ZN(P1_U3229) );
  XNOR2_X1 U8484 ( .A(n6779), .B(n7828), .ZN(n6786) );
  NAND2_X1 U8485 ( .A1(n6809), .A2(n6780), .ZN(n6783) );
  INV_X1 U8486 ( .A(n6781), .ZN(n6782) );
  AOI21_X1 U8487 ( .B1(n7828), .B2(n6783), .A(n6782), .ZN(n6979) );
  AOI22_X1 U8488 ( .A1(n8390), .A2(n8062), .B1(n8060), .B2(n8392), .ZN(n6784)
         );
  OAI21_X1 U8489 ( .B1(n6979), .B2(n8379), .A(n6784), .ZN(n6785) );
  AOI21_X1 U8490 ( .B1(n6786), .B2(n8395), .A(n6785), .ZN(n6978) );
  INV_X1 U8491 ( .A(n6787), .ZN(n6788) );
  AOI21_X1 U8492 ( .B1(n6975), .B2(n6812), .A(n6788), .ZN(n6976) );
  AOI22_X1 U8493 ( .A1(n8368), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n6789), .B2(
        n9944), .ZN(n6790) );
  OAI21_X1 U8494 ( .B1(n5056), .B2(n8406), .A(n6790), .ZN(n6792) );
  NOR2_X1 U8495 ( .A1(n6979), .A2(n8388), .ZN(n6791) );
  AOI211_X1 U8496 ( .C1(n6976), .C2(n8402), .A(n6792), .B(n6791), .ZN(n6793)
         );
  OAI21_X1 U8497 ( .B1(n8368), .B2(n6978), .A(n6793), .ZN(P2_U3287) );
  OR2_X1 U8498 ( .A1(n6889), .A2(n6891), .ZN(n6798) );
  INV_X1 U8499 ( .A(n6794), .ZN(n6797) );
  INV_X1 U8500 ( .A(n6795), .ZN(n6796) );
  NAND2_X1 U8501 ( .A1(n6797), .A2(n6796), .ZN(n6892) );
  NAND2_X1 U8502 ( .A1(n6798), .A2(n6892), .ZN(n6799) );
  XNOR2_X1 U8503 ( .A(n6955), .B(n7926), .ZN(n6896) );
  NAND2_X1 U8504 ( .A1(n8059), .A2(n7635), .ZN(n6894) );
  XNOR2_X1 U8505 ( .A(n6896), .B(n6894), .ZN(n6890) );
  XNOR2_X1 U8506 ( .A(n6799), .B(n6890), .ZN(n6805) );
  INV_X1 U8507 ( .A(n6984), .ZN(n6800) );
  OAI22_X1 U8508 ( .A1(n8045), .A2(n6800), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5311), .ZN(n6803) );
  OAI22_X1 U8509 ( .A1(n6801), .A2(n8030), .B1(n8029), .B2(n6908), .ZN(n6802)
         );
  AOI211_X1 U8510 ( .C1(n8047), .C2(n6955), .A(n6803), .B(n6802), .ZN(n6804)
         );
  OAI21_X1 U8511 ( .B1(n6805), .B2(n8036), .A(n6804), .ZN(P2_U3238) );
  NAND2_X1 U8512 ( .A1(n6613), .A2(n6806), .ZN(n6807) );
  NAND2_X1 U8513 ( .A1(n6807), .A2(n4816), .ZN(n6808) );
  NAND2_X1 U8514 ( .A1(n6809), .A2(n6808), .ZN(n6823) );
  INV_X1 U8515 ( .A(n6823), .ZN(n9999) );
  OR2_X1 U8516 ( .A1(n6810), .A2(n9995), .ZN(n6811) );
  NAND2_X1 U8517 ( .A1(n6812), .A2(n6811), .ZN(n9996) );
  AOI22_X1 U8518 ( .A1(n8359), .A2(n6814), .B1(n9944), .B2(n6813), .ZN(n6815)
         );
  OAI21_X1 U8519 ( .B1(n9996), .B2(n8167), .A(n6815), .ZN(n6825) );
  AND2_X1 U8520 ( .A1(n6817), .A2(n7683), .ZN(n6819) );
  NAND2_X1 U8521 ( .A1(n6817), .A2(n6816), .ZN(n6818) );
  OAI21_X1 U8522 ( .B1(n6819), .B2(n4816), .A(n6818), .ZN(n6820) );
  NAND2_X1 U8523 ( .A1(n6820), .A2(n8395), .ZN(n6822) );
  AOI22_X1 U8524 ( .A1(n8390), .A2(n8063), .B1(n8061), .B2(n8392), .ZN(n6821)
         );
  OAI211_X1 U8525 ( .C1(n8379), .C2(n6823), .A(n6822), .B(n6821), .ZN(n9997)
         );
  MUX2_X1 U8526 ( .A(n9997), .B(P2_REG2_REG_8__SCAN_IN), .S(n8368), .Z(n6824)
         );
  AOI211_X1 U8527 ( .C1(n9999), .C2(n7040), .A(n6825), .B(n6824), .ZN(n6826)
         );
  INV_X1 U8528 ( .A(n6826), .ZN(P2_U3288) );
  NAND2_X1 U8529 ( .A1(n6828), .A2(n6827), .ZN(n7121) );
  NAND2_X1 U8530 ( .A1(n6829), .A2(n8767), .ZN(n6832) );
  AOI22_X1 U8531 ( .A1(n7338), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n9688), .B2(
        n6830), .ZN(n6831) );
  NAND2_X1 U8532 ( .A1(n7066), .A2(n7579), .ZN(n6834) );
  OR2_X1 U8533 ( .A1(n9801), .A2(n6049), .ZN(n6833) );
  NAND2_X1 U8534 ( .A1(n6834), .A2(n6833), .ZN(n6835) );
  XNOR2_X1 U8535 ( .A(n6835), .B(n5923), .ZN(n6838) );
  NAND2_X1 U8536 ( .A1(n7066), .A2(n7592), .ZN(n6837) );
  OR2_X1 U8537 ( .A1(n9801), .A2(n7590), .ZN(n6836) );
  NAND2_X1 U8538 ( .A1(n6837), .A2(n6836), .ZN(n6839) );
  NAND2_X1 U8539 ( .A1(n6838), .A2(n6839), .ZN(n7120) );
  INV_X1 U8540 ( .A(n6838), .ZN(n6841) );
  INV_X1 U8541 ( .A(n6839), .ZN(n6840) );
  NAND2_X1 U8542 ( .A1(n6841), .A2(n6840), .ZN(n7122) );
  NAND2_X1 U8543 ( .A1(n7120), .A2(n7122), .ZN(n6842) );
  XNOR2_X1 U8544 ( .A(n7121), .B(n6842), .ZN(n6855) );
  NOR2_X1 U8545 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6843), .ZN(n9779) );
  AOI21_X1 U8546 ( .B1(n8621), .B2(n8938), .A(n9779), .ZN(n6852) );
  NAND2_X1 U8547 ( .A1(n7555), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n6850) );
  OR2_X1 U8548 ( .A1(n4316), .A2(n9677), .ZN(n6849) );
  AND2_X1 U8549 ( .A1(n6845), .A2(n6844), .ZN(n6846) );
  OR2_X1 U8550 ( .A1(n6846), .A2(n7079), .ZN(n9646) );
  OR2_X1 U8551 ( .A1(n5933), .A2(n9646), .ZN(n6848) );
  OR2_X1 U8552 ( .A1(n7598), .A2(n5986), .ZN(n6847) );
  NAND4_X1 U8553 ( .A1(n6850), .A2(n6849), .A3(n6848), .A4(n6847), .ZN(n8936)
         );
  NAND2_X1 U8554 ( .A1(n4397), .A2(n8936), .ZN(n6851) );
  OAI211_X1 U8555 ( .C1(n8668), .C2(n6942), .A(n6852), .B(n6851), .ZN(n6853)
         );
  AOI21_X1 U8556 ( .B1(n8670), .B2(n7066), .A(n6853), .ZN(n6854) );
  OAI21_X1 U8557 ( .B1(n6855), .B2(n8672), .A(n6854), .ZN(P1_U3215) );
  NAND2_X1 U8558 ( .A1(n7492), .A2(n8530), .ZN(n6856) );
  OAI211_X1 U8559 ( .C1(n6857), .C2(n8534), .A(n6856), .B(n7861), .ZN(P2_U3335) );
  NAND2_X1 U8560 ( .A1(n7492), .A2(n7272), .ZN(n6859) );
  NAND2_X1 U8561 ( .A1(n6858), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8929) );
  OAI211_X1 U8562 ( .C1(n7493), .C2(n9376), .A(n6859), .B(n8929), .ZN(P1_U3330) );
  NAND2_X1 U8563 ( .A1(n6860), .A2(n7704), .ZN(n6861) );
  XNOR2_X1 U8564 ( .A(n6861), .B(n7831), .ZN(n6862) );
  AOI222_X1 U8565 ( .A1(n8395), .A2(n6862), .B1(n8057), .B2(n8392), .C1(n8059), 
        .C2(n8390), .ZN(n10012) );
  XNOR2_X1 U8566 ( .A(n6864), .B(n6863), .ZN(n10016) );
  OAI21_X1 U8567 ( .B1(n6953), .B2(n10009), .A(n7033), .ZN(n10011) );
  AOI22_X1 U8568 ( .A1(n8368), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n6921), .B2(
        n9944), .ZN(n6866) );
  NAND2_X1 U8569 ( .A1(n8359), .A2(n6927), .ZN(n6865) );
  OAI211_X1 U8570 ( .C1(n10011), .C2(n8167), .A(n6866), .B(n6865), .ZN(n6867)
         );
  AOI21_X1 U8571 ( .B1(n10016), .B2(n8409), .A(n6867), .ZN(n6868) );
  OAI21_X1 U8572 ( .B1(n10012), .B2(n8368), .A(n6868), .ZN(P2_U3284) );
  NOR2_X1 U8573 ( .A1(n6870), .A2(n6869), .ZN(n6872) );
  NOR2_X1 U8574 ( .A1(n6872), .A2(n6871), .ZN(n6874) );
  XOR2_X1 U8575 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n8112), .Z(n6873) );
  NAND2_X1 U8576 ( .A1(n6873), .A2(n6874), .ZN(n8111) );
  OAI21_X1 U8577 ( .B1(n6874), .B2(n6873), .A(n8111), .ZN(n6887) );
  NOR2_X1 U8578 ( .A1(n6876), .A2(n6875), .ZN(n6878) );
  INV_X1 U8579 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n6880) );
  NAND2_X1 U8580 ( .A1(n8112), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n8106) );
  INV_X1 U8581 ( .A(n8106), .ZN(n6879) );
  AOI21_X1 U8582 ( .B1(n6880), .B2(n6885), .A(n6879), .ZN(n6881) );
  OAI211_X1 U8583 ( .C1(n6882), .C2(n6881), .A(n9929), .B(n8105), .ZN(n6884)
         );
  AND2_X1 U8584 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3152), .ZN(n7983) );
  AOI21_X1 U8585 ( .B1(n9935), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n7983), .ZN(
        n6883) );
  OAI211_X1 U8586 ( .C1(n9932), .C2(n6885), .A(n6884), .B(n6883), .ZN(n6886)
         );
  AOI21_X1 U8587 ( .B1(n9930), .B2(n6887), .A(n6886), .ZN(n6888) );
  INV_X1 U8588 ( .A(n6888), .ZN(P2_U3261) );
  INV_X1 U8589 ( .A(n6889), .ZN(n6907) );
  INV_X1 U8590 ( .A(n6890), .ZN(n6893) );
  OR2_X1 U8591 ( .A1(n6891), .A2(n6893), .ZN(n6914) );
  XNOR2_X1 U8592 ( .A(n6927), .B(n7921), .ZN(n6899) );
  NAND2_X1 U8593 ( .A1(n8058), .A2(n7635), .ZN(n6900) );
  NAND2_X1 U8594 ( .A1(n6899), .A2(n6900), .ZN(n6904) );
  INV_X1 U8595 ( .A(n6904), .ZN(n6906) );
  INV_X1 U8596 ( .A(n6894), .ZN(n6895) );
  NAND2_X1 U8597 ( .A1(n6896), .A2(n6895), .ZN(n6897) );
  AND2_X1 U8598 ( .A1(n6898), .A2(n6897), .ZN(n6915) );
  INV_X1 U8599 ( .A(n6899), .ZN(n6902) );
  INV_X1 U8600 ( .A(n6900), .ZN(n6901) );
  NAND2_X1 U8601 ( .A1(n6902), .A2(n6901), .ZN(n6903) );
  NAND2_X1 U8602 ( .A1(n6904), .A2(n6903), .ZN(n6920) );
  INV_X1 U8603 ( .A(n6920), .ZN(n6905) );
  AND2_X1 U8604 ( .A1(n6915), .A2(n6905), .ZN(n6916) );
  XNOR2_X1 U8605 ( .A(n8505), .B(n7921), .ZN(n7048) );
  NAND2_X1 U8606 ( .A1(n8057), .A2(n7635), .ZN(n7047) );
  XNOR2_X1 U8607 ( .A(n7048), .B(n7047), .ZN(n7049) );
  XNOR2_X1 U8608 ( .A(n7050), .B(n7049), .ZN(n6913) );
  OAI22_X1 U8609 ( .A1(n6908), .A2(n8030), .B1(n8029), .B2(n7111), .ZN(n6909)
         );
  AOI211_X1 U8610 ( .C1(n8033), .C2(n7036), .A(n6910), .B(n6909), .ZN(n6912)
         );
  NAND2_X1 U8611 ( .A1(n8047), .A2(n8505), .ZN(n6911) );
  OAI211_X1 U8612 ( .C1(n6913), .C2(n8036), .A(n6912), .B(n6911), .ZN(P2_U3236) );
  OR2_X1 U8613 ( .A1(n6889), .A2(n6914), .ZN(n6917) );
  NAND2_X1 U8614 ( .A1(n6917), .A2(n6915), .ZN(n6919) );
  AND2_X1 U8615 ( .A1(n6917), .A2(n6916), .ZN(n6918) );
  AOI21_X1 U8616 ( .B1(n6920), .B2(n6919), .A(n6918), .ZN(n6929) );
  INV_X1 U8617 ( .A(n6921), .ZN(n6923) );
  OAI21_X1 U8618 ( .B1(n8045), .B2(n6923), .A(n6922), .ZN(n6926) );
  OAI22_X1 U8619 ( .A1(n6924), .A2(n8030), .B1(n8029), .B2(n7055), .ZN(n6925)
         );
  AOI211_X1 U8620 ( .C1(n8047), .C2(n6927), .A(n6926), .B(n6925), .ZN(n6928)
         );
  OAI21_X1 U8621 ( .B1(n6929), .B2(n8036), .A(n6928), .ZN(P2_U3226) );
  NAND2_X1 U8622 ( .A1(n9907), .A2(n6936), .ZN(n6932) );
  NAND2_X1 U8623 ( .A1(n7066), .A2(n9801), .ZN(n8693) );
  NAND2_X1 U8624 ( .A1(n8850), .A2(n8693), .ZN(n6937) );
  OAI21_X1 U8625 ( .B1(n6933), .B2(n6937), .A(n7068), .ZN(n6934) );
  INV_X1 U8626 ( .A(n6934), .ZN(n7000) );
  NAND2_X1 U8627 ( .A1(n6935), .A2(n8830), .ZN(n9797) );
  OR2_X1 U8628 ( .A1(n6941), .A2(n6936), .ZN(n8788) );
  AND2_X1 U8629 ( .A1(n8788), .A2(n9796), .ZN(n8849) );
  AND2_X1 U8630 ( .A1(n6941), .A2(n6936), .ZN(n8691) );
  AOI21_X1 U8631 ( .B1(n9797), .B2(n8849), .A(n8691), .ZN(n6938) );
  INV_X1 U8632 ( .A(n6937), .ZN(n8790) );
  OAI211_X1 U8633 ( .C1(n6938), .C2(n8790), .A(n7094), .B(n9823), .ZN(n6940)
         );
  AOI22_X1 U8634 ( .A1(n8938), .A2(n9825), .B1(n9828), .B2(n8936), .ZN(n6939)
         );
  NAND2_X1 U8635 ( .A1(n6940), .A2(n6939), .ZN(n6997) );
  INV_X1 U8636 ( .A(n7066), .ZN(n6946) );
  AOI211_X1 U8637 ( .C1(n7066), .C2(n9791), .A(n9908), .B(n9635), .ZN(n6998)
         );
  NAND2_X1 U8638 ( .A1(n6998), .A2(n9228), .ZN(n6945) );
  INV_X1 U8639 ( .A(n6942), .ZN(n6943) );
  AOI22_X1 U8640 ( .A1(n9844), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n6943), .B2(
        n9838), .ZN(n6944) );
  OAI211_X1 U8641 ( .C1(n6946), .C2(n9808), .A(n6945), .B(n6944), .ZN(n6947)
         );
  AOI21_X1 U8642 ( .B1(n9814), .B2(n6997), .A(n6947), .ZN(n6948) );
  OAI21_X1 U8643 ( .B1(n7000), .B2(n9256), .A(n6948), .ZN(P1_U3281) );
  INV_X1 U8644 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n6958) );
  XNOR2_X1 U8645 ( .A(n6949), .B(n7830), .ZN(n6987) );
  XNOR2_X1 U8646 ( .A(n6950), .B(n7830), .ZN(n6951) );
  AOI222_X1 U8647 ( .A1(n8395), .A2(n6951), .B1(n8058), .B2(n8392), .C1(n8060), 
        .C2(n8390), .ZN(n6992) );
  INV_X1 U8648 ( .A(n6952), .ZN(n6954) );
  AOI21_X1 U8649 ( .B1(n6955), .B2(n6954), .A(n6953), .ZN(n6990) );
  AOI22_X1 U8650 ( .A1(n6990), .A2(n8499), .B1(n8498), .B2(n6955), .ZN(n6956)
         );
  OAI211_X1 U8651 ( .C1(n8503), .C2(n6987), .A(n6992), .B(n6956), .ZN(n6959)
         );
  NAND2_X1 U8652 ( .A1(n6959), .A2(n10019), .ZN(n6957) );
  OAI21_X1 U8653 ( .B1(n10019), .B2(n6958), .A(n6957), .ZN(P2_U3484) );
  NAND2_X1 U8654 ( .A1(n6959), .A2(n10033), .ZN(n6960) );
  OAI21_X1 U8655 ( .B1(n10033), .B2(n6961), .A(n6960), .ZN(P2_U3531) );
  INV_X1 U8656 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n6974) );
  NOR2_X1 U8657 ( .A1(n6963), .A2(n6962), .ZN(n6965) );
  NOR2_X1 U8658 ( .A1(n6965), .A2(n6964), .ZN(n7143) );
  XNOR2_X1 U8659 ( .A(n7143), .B(n7150), .ZN(n6966) );
  INV_X1 U8660 ( .A(n6966), .ZN(n6968) );
  INV_X1 U8661 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n7225) );
  NOR2_X1 U8662 ( .A1(n7225), .A2(n6966), .ZN(n7144) );
  INV_X1 U8663 ( .A(n7144), .ZN(n6967) );
  OAI211_X1 U8664 ( .C1(n6968), .C2(P1_REG2_REG_15__SCAN_IN), .A(n9751), .B(
        n6967), .ZN(n6973) );
  INV_X1 U8665 ( .A(n7150), .ZN(n7304) );
  AND2_X1 U8666 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n8665) );
  OAI21_X1 U8667 ( .B1(n7210), .B2(P1_REG1_REG_14__SCAN_IN), .A(n6969), .ZN(
        n7149) );
  XNOR2_X1 U8668 ( .A(n7150), .B(n7149), .ZN(n6970) );
  INV_X1 U8669 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n7222) );
  NOR2_X1 U8670 ( .A1(n7222), .A2(n6970), .ZN(n7151) );
  AOI211_X1 U8671 ( .C1(n6970), .C2(n7222), .A(n7151), .B(n9744), .ZN(n6971)
         );
  AOI211_X1 U8672 ( .C1(n9758), .C2(n7304), .A(n8665), .B(n6971), .ZN(n6972)
         );
  OAI211_X1 U8673 ( .C1(n9785), .C2(n6974), .A(n6973), .B(n6972), .ZN(P1_U3256) );
  AOI22_X1 U8674 ( .A1(n6976), .A2(n8499), .B1(n8498), .B2(n6975), .ZN(n6977)
         );
  OAI211_X1 U8675 ( .C1(n6979), .C2(n8487), .A(n6978), .B(n6977), .ZN(n6981)
         );
  NAND2_X1 U8676 ( .A1(n6981), .A2(n10033), .ZN(n6980) );
  OAI21_X1 U8677 ( .B1(n10033), .B2(n5778), .A(n6980), .ZN(P2_U3529) );
  INV_X1 U8678 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n6983) );
  NAND2_X1 U8679 ( .A1(n6981), .A2(n10019), .ZN(n6982) );
  OAI21_X1 U8680 ( .B1(n10019), .B2(n6983), .A(n6982), .ZN(P2_U3478) );
  AOI22_X1 U8681 ( .A1(n8368), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n6984), .B2(
        n9944), .ZN(n6985) );
  OAI21_X1 U8682 ( .B1(n6986), .B2(n8406), .A(n6985), .ZN(n6989) );
  NOR2_X1 U8683 ( .A1(n6987), .A2(n8365), .ZN(n6988) );
  AOI211_X1 U8684 ( .C1(n6990), .C2(n8402), .A(n6989), .B(n6988), .ZN(n6991)
         );
  OAI21_X1 U8685 ( .B1(n8368), .B2(n6992), .A(n6991), .ZN(P2_U3285) );
  OR2_X1 U8686 ( .A1(n9908), .A2(n9154), .ZN(n6994) );
  AND2_X2 U8687 ( .A1(n7007), .A2(n6995), .ZN(n9916) );
  INV_X1 U8688 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n7002) );
  NAND2_X1 U8689 ( .A1(n5859), .A2(n9840), .ZN(n8773) );
  OR2_X1 U8690 ( .A1(n8773), .A2(n6996), .ZN(n9667) );
  NAND2_X1 U8691 ( .A1(n9884), .A2(n9667), .ZN(n9895) );
  AOI211_X1 U8692 ( .C1(n7066), .C2(n9664), .A(n6998), .B(n6997), .ZN(n6999)
         );
  OAI21_X1 U8693 ( .B1(n7000), .B2(n9897), .A(n6999), .ZN(n7008) );
  NAND2_X1 U8694 ( .A1(n7008), .A2(n9916), .ZN(n7001) );
  OAI21_X1 U8695 ( .B1(n9916), .B2(n7002), .A(n7001), .ZN(P1_U3484) );
  NOR2_X1 U8696 ( .A1(n7003), .A2(n9850), .ZN(n7004) );
  AND2_X1 U8697 ( .A1(n7005), .A2(n7004), .ZN(n7006) );
  AND2_X2 U8698 ( .A1(n7007), .A2(n7006), .ZN(n9928) );
  NAND2_X1 U8699 ( .A1(n7008), .A2(n9928), .ZN(n7009) );
  OAI21_X1 U8700 ( .B1(n9928), .B2(n6766), .A(n7009), .ZN(P1_U3533) );
  INV_X1 U8701 ( .A(n7510), .ZN(n7012) );
  INV_X1 U8702 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7511) );
  OAI222_X1 U8703 ( .A1(n9373), .A2(n7012), .B1(P1_U3084), .B2(n7010), .C1(
        n7511), .C2(n9376), .ZN(P1_U3329) );
  OAI222_X1 U8704 ( .A1(P2_U3152), .A2(n7013), .B1(n7939), .B2(n7012), .C1(
        n7011), .C2(n8534), .ZN(P2_U3334) );
  XNOR2_X1 U8705 ( .A(n7014), .B(n7833), .ZN(n8504) );
  AOI21_X1 U8706 ( .B1(n8497), .B2(n7035), .A(n8399), .ZN(n8500) );
  INV_X1 U8707 ( .A(n8497), .ZN(n7016) );
  AOI22_X1 U8708 ( .A1(n8368), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n7058), .B2(
        n9944), .ZN(n7015) );
  OAI21_X1 U8709 ( .B1(n7016), .B2(n8406), .A(n7015), .ZN(n7022) );
  AOI21_X1 U8710 ( .B1(n7017), .B2(n7833), .A(n8347), .ZN(n7020) );
  OAI22_X1 U8711 ( .A1(n7981), .A2(n8307), .B1(n7055), .B2(n8305), .ZN(n7018)
         );
  AOI21_X1 U8712 ( .B1(n7020), .B2(n7019), .A(n7018), .ZN(n8502) );
  NOR2_X1 U8713 ( .A1(n8502), .A2(n8368), .ZN(n7021) );
  AOI211_X1 U8714 ( .C1(n8500), .C2(n8402), .A(n7022), .B(n7021), .ZN(n7023)
         );
  OAI21_X1 U8715 ( .B1(n8365), .B2(n8504), .A(n7023), .ZN(P2_U3282) );
  NAND2_X1 U8716 ( .A1(n7024), .A2(n7834), .ZN(n7025) );
  NAND2_X1 U8717 ( .A1(n7026), .A2(n7025), .ZN(n7032) );
  OR2_X1 U8718 ( .A1(n7032), .A2(n8379), .ZN(n7031) );
  AOI22_X1 U8719 ( .A1(n8390), .A2(n8058), .B1(n8391), .B2(n8392), .ZN(n7030)
         );
  XNOR2_X1 U8720 ( .A(n7027), .B(n7834), .ZN(n7028) );
  NAND2_X1 U8721 ( .A1(n7028), .A2(n8395), .ZN(n7029) );
  INV_X1 U8722 ( .A(n7032), .ZN(n8509) );
  NAND2_X1 U8723 ( .A1(n7033), .A2(n8505), .ZN(n7034) );
  NAND2_X1 U8724 ( .A1(n7035), .A2(n7034), .ZN(n8507) );
  AOI22_X1 U8725 ( .A1(n8368), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n7036), .B2(
        n9944), .ZN(n7038) );
  NAND2_X1 U8726 ( .A1(n8505), .A2(n8359), .ZN(n7037) );
  OAI211_X1 U8727 ( .C1(n8507), .C2(n8167), .A(n7038), .B(n7037), .ZN(n7039)
         );
  AOI21_X1 U8728 ( .B1(n8509), .B2(n7040), .A(n7039), .ZN(n7041) );
  OAI21_X1 U8729 ( .B1(n8511), .B2(n8368), .A(n7041), .ZN(P2_U3283) );
  XNOR2_X1 U8730 ( .A(n8497), .B(n7921), .ZN(n7042) );
  NAND2_X1 U8731 ( .A1(n8391), .A2(n7635), .ZN(n7043) );
  NAND2_X1 U8732 ( .A1(n7042), .A2(n7043), .ZN(n7105) );
  INV_X1 U8733 ( .A(n7042), .ZN(n7045) );
  INV_X1 U8734 ( .A(n7043), .ZN(n7044) );
  NAND2_X1 U8735 ( .A1(n7045), .A2(n7044), .ZN(n7046) );
  NAND2_X1 U8736 ( .A1(n7105), .A2(n7046), .ZN(n7054) );
  INV_X1 U8737 ( .A(n7106), .ZN(n7052) );
  AOI21_X1 U8738 ( .B1(n7054), .B2(n7053), .A(n7052), .ZN(n7061) );
  OAI22_X1 U8739 ( .A1(n7981), .A2(n8029), .B1(n8030), .B2(n7055), .ZN(n7056)
         );
  AOI211_X1 U8740 ( .C1(n8033), .C2(n7058), .A(n7057), .B(n7056), .ZN(n7060)
         );
  NAND2_X1 U8741 ( .A1(n8497), .A2(n8047), .ZN(n7059) );
  OAI211_X1 U8742 ( .C1(n7061), .C2(n8036), .A(n7060), .B(n7059), .ZN(P2_U3217) );
  INV_X1 U8743 ( .A(n7526), .ZN(n7065) );
  OAI222_X1 U8744 ( .A1(n8534), .A2(n7063), .B1(n7939), .B2(n7065), .C1(
        P2_U3152), .C2(n7062), .ZN(P2_U3333) );
  OAI222_X1 U8745 ( .A1(n9376), .A2(n7527), .B1(n9373), .B2(n7065), .C1(n7064), 
        .C2(P1_U3084), .ZN(P1_U3328) );
  NAND2_X1 U8746 ( .A1(n7069), .A2(n8767), .ZN(n7072) );
  AOI22_X1 U8747 ( .A1(n7338), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n9688), .B2(
        n7070), .ZN(n7071) );
  NAND2_X1 U8748 ( .A1(n7073), .A2(n8767), .ZN(n7077) );
  INV_X1 U8749 ( .A(n7074), .ZN(n7075) );
  AOI22_X1 U8750 ( .A1(n7338), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n9688), .B2(
        n7075), .ZN(n7076) );
  NAND2_X1 U8751 ( .A1(n7555), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n7085) );
  OR2_X1 U8752 ( .A1(n4315), .A2(n7078), .ZN(n7084) );
  OR2_X1 U8753 ( .A1(n7079), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n7080) );
  NAND2_X1 U8754 ( .A1(n7088), .A2(n7080), .ZN(n7100) );
  OR2_X1 U8755 ( .A1(n5933), .A2(n7100), .ZN(n7083) );
  OR2_X1 U8756 ( .A1(n7598), .A2(n7081), .ZN(n7082) );
  NAND2_X1 U8757 ( .A1(n9665), .A2(n9641), .ZN(n8699) );
  NAND2_X1 U8758 ( .A1(n8701), .A2(n8699), .ZN(n7095) );
  OAI21_X1 U8759 ( .B1(n7086), .B2(n7095), .A(n7214), .ZN(n9668) );
  NAND2_X1 U8760 ( .A1(n7555), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n7093) );
  OR2_X1 U8761 ( .A1(n4316), .A2(n9661), .ZN(n7092) );
  NAND2_X1 U8762 ( .A1(n7088), .A2(n7087), .ZN(n7089) );
  NAND2_X1 U8763 ( .A1(n7178), .A2(n7089), .ZN(n7261) );
  OR2_X1 U8764 ( .A1(n5933), .A2(n7261), .ZN(n7091) );
  INV_X1 U8765 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7262) );
  OR2_X1 U8766 ( .A1(n7598), .A2(n7262), .ZN(n7090) );
  INV_X1 U8767 ( .A(n8936), .ZN(n7098) );
  NAND2_X1 U8768 ( .A1(n8692), .A2(n7098), .ZN(n8698) );
  OR2_X1 U8769 ( .A1(n8692), .A2(n7098), .ZN(n7230) );
  NAND2_X1 U8770 ( .A1(n7231), .A2(n7230), .ZN(n7096) );
  INV_X1 U8771 ( .A(n7095), .ZN(n8791) );
  XNOR2_X1 U8772 ( .A(n7096), .B(n8791), .ZN(n7097) );
  OAI222_X1 U8773 ( .A1(n9800), .A2(n7248), .B1(n9802), .B2(n7098), .C1(n9242), 
        .C2(n7097), .ZN(n9662) );
  INV_X1 U8774 ( .A(n9665), .ZN(n7213) );
  NAND2_X1 U8775 ( .A1(n9635), .A2(n9672), .ZN(n9637) );
  INV_X1 U8776 ( .A(n7263), .ZN(n7099) );
  AOI211_X1 U8777 ( .C1(n9665), .C2(n9637), .A(n9908), .B(n7099), .ZN(n9663)
         );
  NAND2_X1 U8778 ( .A1(n9663), .A2(n9228), .ZN(n7102) );
  INV_X1 U8779 ( .A(n7100), .ZN(n7140) );
  AOI22_X1 U8780 ( .A1(n9844), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n7140), .B2(
        n9838), .ZN(n7101) );
  OAI211_X1 U8781 ( .C1(n7213), .C2(n9808), .A(n7102), .B(n7101), .ZN(n7103)
         );
  AOI21_X1 U8782 ( .B1(n9662), .B2(n9814), .A(n7103), .ZN(n7104) );
  OAI21_X1 U8783 ( .B1(n9668), .B2(n9256), .A(n7104), .ZN(P1_U3279) );
  XNOR2_X1 U8784 ( .A(n8492), .B(n7921), .ZN(n7866) );
  INV_X1 U8785 ( .A(n7866), .ZN(n7869) );
  AND2_X1 U8786 ( .A1(n8373), .A2(n7635), .ZN(n7867) );
  XNOR2_X1 U8787 ( .A(n7869), .B(n7867), .ZN(n7107) );
  XNOR2_X1 U8788 ( .A(n7868), .B(n7107), .ZN(n7115) );
  INV_X1 U8789 ( .A(n8403), .ZN(n7109) );
  OAI22_X1 U8790 ( .A1(n8045), .A2(n7109), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7108), .ZN(n7113) );
  OAI22_X1 U8791 ( .A1(n7111), .A2(n8030), .B1(n8029), .B2(n7110), .ZN(n7112)
         );
  AOI211_X1 U8792 ( .C1(n8047), .C2(n8492), .A(n7113), .B(n7112), .ZN(n7114)
         );
  OAI21_X1 U8793 ( .B1(n7115), .B2(n8036), .A(n7114), .ZN(P2_U3243) );
  NAND2_X1 U8794 ( .A1(n9665), .A2(n7579), .ZN(n7117) );
  OR2_X1 U8795 ( .A1(n9641), .A2(n6049), .ZN(n7116) );
  NAND2_X1 U8796 ( .A1(n7117), .A2(n7116), .ZN(n7118) );
  XNOR2_X1 U8797 ( .A(n7118), .B(n5923), .ZN(n7163) );
  NOR2_X1 U8798 ( .A1(n9641), .A2(n7590), .ZN(n7119) );
  AOI21_X1 U8799 ( .B1(n9665), .B2(n7592), .A(n7119), .ZN(n7164) );
  XNOR2_X1 U8800 ( .A(n7163), .B(n7164), .ZN(n7136) );
  NAND2_X1 U8801 ( .A1(n7121), .A2(n7120), .ZN(n7123) );
  NAND2_X1 U8802 ( .A1(n7123), .A2(n7122), .ZN(n7199) );
  INV_X1 U8803 ( .A(n7199), .ZN(n7129) );
  NAND2_X1 U8804 ( .A1(n8692), .A2(n7579), .ZN(n7125) );
  NAND2_X1 U8805 ( .A1(n8936), .A2(n7592), .ZN(n7124) );
  NAND2_X1 U8806 ( .A1(n7125), .A2(n7124), .ZN(n7126) );
  XNOR2_X1 U8807 ( .A(n7126), .B(n7564), .ZN(n7130) );
  AND2_X1 U8808 ( .A1(n8936), .A2(n7566), .ZN(n7127) );
  AOI21_X1 U8809 ( .B1(n8692), .B2(n7592), .A(n7127), .ZN(n7131) );
  XNOR2_X1 U8810 ( .A(n7130), .B(n7131), .ZN(n7203) );
  INV_X1 U8811 ( .A(n7203), .ZN(n7128) );
  NAND2_X1 U8812 ( .A1(n7129), .A2(n7128), .ZN(n7201) );
  INV_X1 U8813 ( .A(n7130), .ZN(n7133) );
  INV_X1 U8814 ( .A(n7131), .ZN(n7132) );
  NAND2_X1 U8815 ( .A1(n7133), .A2(n7132), .ZN(n7134) );
  OAI21_X1 U8816 ( .B1(n7136), .B2(n7135), .A(n7167), .ZN(n7137) );
  NAND2_X1 U8817 ( .A1(n7137), .A2(n8597), .ZN(n7142) );
  AOI22_X1 U8818 ( .A1(n8621), .A2(n8936), .B1(P1_REG3_REG_12__SCAN_IN), .B2(
        P1_U3084), .ZN(n7138) );
  OAI21_X1 U8819 ( .B1(n7248), .B2(n8599), .A(n7138), .ZN(n7139) );
  AOI21_X1 U8820 ( .B1(n7140), .B2(n8655), .A(n7139), .ZN(n7141) );
  OAI211_X1 U8821 ( .C1(n7213), .C2(n8658), .A(n7142), .B(n7141), .ZN(P1_U3222) );
  NOR2_X1 U8822 ( .A1(n7143), .A2(n7150), .ZN(n7145) );
  NAND2_X1 U8823 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n8952), .ZN(n7146) );
  OAI21_X1 U8824 ( .B1(n8952), .B2(P1_REG2_REG_16__SCAN_IN), .A(n7146), .ZN(
        n7147) );
  AOI211_X1 U8825 ( .C1(n7148), .C2(n7147), .A(n8951), .B(n9774), .ZN(n7161)
         );
  NOR2_X1 U8826 ( .A1(n7150), .A2(n7149), .ZN(n7152) );
  NOR2_X1 U8827 ( .A1(n7152), .A2(n7151), .ZN(n7154) );
  XNOR2_X1 U8828 ( .A(n8952), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n7153) );
  NOR2_X1 U8829 ( .A1(n7154), .A2(n7153), .ZN(n8946) );
  AOI211_X1 U8830 ( .C1(n7154), .C2(n7153), .A(n8946), .B(n9744), .ZN(n7160)
         );
  NAND2_X1 U8831 ( .A1(n9759), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n7157) );
  INV_X1 U8832 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n7155) );
  NOR2_X1 U8833 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7155), .ZN(n8589) );
  INV_X1 U8834 ( .A(n8589), .ZN(n7156) );
  OAI211_X1 U8835 ( .C1(n9783), .C2(n7158), .A(n7157), .B(n7156), .ZN(n7159)
         );
  OR3_X1 U8836 ( .A1(n7161), .A2(n7160), .A3(n7159), .ZN(P1_U3257) );
  INV_X1 U8837 ( .A(n7547), .ZN(n7192) );
  OAI222_X1 U8838 ( .A1(n9373), .A2(n7192), .B1(P1_U3084), .B2(n7162), .C1(
        n7548), .C2(n9376), .ZN(P1_U3327) );
  INV_X1 U8839 ( .A(n7163), .ZN(n7165) );
  NAND2_X1 U8840 ( .A1(n7165), .A2(n7164), .ZN(n7166) );
  NAND2_X1 U8841 ( .A1(n7168), .A2(n8767), .ZN(n7171) );
  AOI22_X1 U8842 ( .A1(n7338), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n9688), .B2(
        n7169), .ZN(n7170) );
  OAI22_X1 U8843 ( .A1(n9656), .A2(n6055), .B1(n7248), .B2(n6049), .ZN(n7172)
         );
  XNOR2_X1 U8844 ( .A(n7172), .B(n7564), .ZN(n7238) );
  OR2_X1 U8845 ( .A1(n9656), .A2(n6049), .ZN(n7174) );
  OR2_X1 U8846 ( .A1(n7248), .A2(n7590), .ZN(n7173) );
  XNOR2_X1 U8847 ( .A(n7238), .B(n7239), .ZN(n7175) );
  XNOR2_X1 U8848 ( .A(n7243), .B(n7175), .ZN(n7190) );
  NAND2_X1 U8849 ( .A1(n7555), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n7183) );
  OR2_X1 U8850 ( .A1(n4316), .A2(n7176), .ZN(n7182) );
  AND2_X1 U8851 ( .A1(n7178), .A2(n7177), .ZN(n7179) );
  OR2_X1 U8852 ( .A1(n7179), .A2(n7223), .ZN(n7252) );
  OR2_X1 U8853 ( .A1(n5933), .A2(n7252), .ZN(n7181) );
  OR2_X1 U8854 ( .A1(n7598), .A2(n6708), .ZN(n7180) );
  INV_X1 U8855 ( .A(n7184), .ZN(n7186) );
  NOR2_X1 U8856 ( .A1(n8663), .A2(n9641), .ZN(n7185) );
  AOI211_X1 U8857 ( .C1(n4397), .C2(n4439), .A(n7186), .B(n7185), .ZN(n7187)
         );
  OAI21_X1 U8858 ( .B1(n8668), .B2(n7261), .A(n7187), .ZN(n7188) );
  AOI21_X1 U8859 ( .B1(n7268), .B2(n8670), .A(n7188), .ZN(n7189) );
  OAI21_X1 U8860 ( .B1(n7190), .B2(n8672), .A(n7189), .ZN(P1_U3232) );
  OAI222_X1 U8861 ( .A1(P2_U3152), .A2(n7193), .B1(n7939), .B2(n7192), .C1(
        n7191), .C2(n8534), .ZN(P2_U3332) );
  INV_X1 U8862 ( .A(n7575), .ZN(n7207) );
  AOI21_X1 U8863 ( .B1(n9366), .B2(P2_DATAO_REG_27__SCAN_IN), .A(n7194), .ZN(
        n7195) );
  OAI21_X1 U8864 ( .B1(n7207), .B2(n9373), .A(n7195), .ZN(P1_U3326) );
  INV_X1 U8865 ( .A(n9641), .ZN(n8935) );
  AOI21_X1 U8866 ( .B1(n8666), .B2(n8935), .A(n7196), .ZN(n7198) );
  NAND2_X1 U8867 ( .A1(n8621), .A2(n8937), .ZN(n7197) );
  OAI211_X1 U8868 ( .C1(n8668), .C2(n9646), .A(n7198), .B(n7197), .ZN(n7205)
         );
  INV_X1 U8869 ( .A(n7201), .ZN(n7202) );
  AOI211_X1 U8870 ( .C1(n7203), .C2(n7200), .A(n8672), .B(n7202), .ZN(n7204)
         );
  AOI211_X1 U8871 ( .C1(n8670), .C2(n8692), .A(n7205), .B(n7204), .ZN(n7206)
         );
  INV_X1 U8872 ( .A(n7206), .ZN(P1_U3234) );
  OAI222_X1 U8873 ( .A1(n8534), .A2(n7208), .B1(n7939), .B2(n7207), .C1(n4994), 
        .C2(P2_U3152), .ZN(P2_U3331) );
  NAND2_X1 U8874 ( .A1(n7209), .A2(n8767), .ZN(n7212) );
  AOI22_X1 U8875 ( .A1(n7338), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n9688), .B2(
        n7210), .ZN(n7211) );
  NAND2_X1 U8876 ( .A1(n9339), .A2(n9243), .ZN(n8857) );
  NAND2_X1 U8877 ( .A1(n8716), .A2(n8857), .ZN(n8795) );
  NAND2_X1 U8878 ( .A1(n9656), .A2(n7248), .ZN(n7215) );
  NAND2_X1 U8879 ( .A1(n7256), .A2(n7215), .ZN(n7217) );
  INV_X1 U8880 ( .A(n7248), .ZN(n8934) );
  XOR2_X1 U8881 ( .A(n8795), .B(n7218), .Z(n9342) );
  INV_X1 U8882 ( .A(n7264), .ZN(n7219) );
  AOI211_X1 U8883 ( .C1(n9339), .C2(n7219), .A(n9908), .B(n9245), .ZN(n9338)
         );
  INV_X1 U8884 ( .A(n7252), .ZN(n7220) );
  AOI22_X1 U8885 ( .A1(n9844), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n7220), .B2(
        n9838), .ZN(n7221) );
  OAI21_X1 U8886 ( .B1(n7300), .B2(n9808), .A(n7221), .ZN(n7236) );
  NAND2_X1 U8887 ( .A1(n7555), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n7229) );
  OR2_X1 U8888 ( .A1(n4315), .A2(n7222), .ZN(n7228) );
  NOR2_X1 U8889 ( .A1(n7223), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n7224) );
  OR2_X1 U8890 ( .A1(n7311), .A2(n7224), .ZN(n9249) );
  OR2_X1 U8891 ( .A1(n5933), .A2(n9249), .ZN(n7227) );
  OR2_X1 U8892 ( .A1(n7598), .A2(n7225), .ZN(n7226) );
  NAND4_X1 U8893 ( .A1(n7229), .A2(n7228), .A3(n7227), .A4(n7226), .ZN(n8933)
         );
  NOR2_X1 U8894 ( .A1(n7248), .A2(n9802), .ZN(n7234) );
  AND2_X1 U8895 ( .A1(n8701), .A2(n7230), .ZN(n8697) );
  INV_X1 U8896 ( .A(n8699), .ZN(n8696) );
  OR2_X1 U8897 ( .A1(n7268), .A2(n7248), .ZN(n8695) );
  NAND2_X1 U8898 ( .A1(n7268), .A2(n7248), .ZN(n8855) );
  NAND2_X1 U8899 ( .A1(n8695), .A2(n8855), .ZN(n8793) );
  AOI211_X1 U8900 ( .C1(n8795), .C2(n7232), .A(n9242), .B(n7381), .ZN(n7233)
         );
  AOI211_X1 U8901 ( .C1(n9828), .C2(n8933), .A(n7234), .B(n7233), .ZN(n9341)
         );
  NOR2_X1 U8902 ( .A1(n9341), .A2(n9844), .ZN(n7235) );
  AOI211_X1 U8903 ( .C1(n9228), .C2(n9338), .A(n7236), .B(n7235), .ZN(n7237)
         );
  OAI21_X1 U8904 ( .B1(n9342), .B2(n9256), .A(n7237), .ZN(P1_U3277) );
  AND2_X1 U8905 ( .A1(n7238), .A2(n7239), .ZN(n7242) );
  INV_X1 U8906 ( .A(n7238), .ZN(n7241) );
  INV_X1 U8907 ( .A(n7239), .ZN(n7240) );
  OAI22_X1 U8908 ( .A1(n7300), .A2(n6055), .B1(n9243), .B2(n6049), .ZN(n7244)
         );
  XNOR2_X1 U8909 ( .A(n7244), .B(n5923), .ZN(n7423) );
  OR2_X1 U8910 ( .A1(n7300), .A2(n6049), .ZN(n7246) );
  OR2_X1 U8911 ( .A1(n9243), .A2(n7590), .ZN(n7245) );
  NAND2_X1 U8912 ( .A1(n7246), .A2(n7245), .ZN(n7422) );
  INV_X1 U8913 ( .A(n7422), .ZN(n7420) );
  XNOR2_X1 U8914 ( .A(n7423), .B(n7420), .ZN(n7247) );
  XNOR2_X1 U8915 ( .A(n7436), .B(n7247), .ZN(n7255) );
  NOR2_X1 U8916 ( .A1(n8663), .A2(n7248), .ZN(n7249) );
  AOI211_X1 U8917 ( .C1(n4397), .C2(n8933), .A(n7250), .B(n7249), .ZN(n7251)
         );
  OAI21_X1 U8918 ( .B1(n8668), .B2(n7252), .A(n7251), .ZN(n7253) );
  AOI21_X1 U8919 ( .B1(n9339), .B2(n8670), .A(n7253), .ZN(n7254) );
  OAI21_X1 U8920 ( .B1(n7255), .B2(n8672), .A(n7254), .ZN(P1_U3213) );
  XNOR2_X1 U8921 ( .A(n7256), .B(n8793), .ZN(n9655) );
  XNOR2_X1 U8922 ( .A(n7257), .B(n8793), .ZN(n7259) );
  OAI22_X1 U8923 ( .A1(n9243), .A2(n9800), .B1(n9641), .B2(n9802), .ZN(n7258)
         );
  AOI21_X1 U8924 ( .B1(n7259), .B2(n9823), .A(n7258), .ZN(n7260) );
  OAI21_X1 U8925 ( .B1(n9655), .B2(n9884), .A(n7260), .ZN(n9658) );
  NAND2_X1 U8926 ( .A1(n9658), .A2(n9814), .ZN(n7270) );
  OAI22_X1 U8927 ( .A1(n9814), .A2(n7262), .B1(n7261), .B2(n9809), .ZN(n7267)
         );
  AND2_X1 U8928 ( .A1(n7263), .A2(n7268), .ZN(n7265) );
  OR2_X1 U8929 ( .A1(n7265), .A2(n7264), .ZN(n9657) );
  NOR2_X1 U8930 ( .A1(n9657), .A2(n9063), .ZN(n7266) );
  AOI211_X1 U8931 ( .C1(n9174), .C2(n7268), .A(n7267), .B(n7266), .ZN(n7269)
         );
  OAI211_X1 U8932 ( .C1(n9655), .C2(n7271), .A(n7270), .B(n7269), .ZN(P1_U3278) );
  INV_X1 U8933 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n7403) );
  NAND2_X1 U8934 ( .A1(n7402), .A2(n7272), .ZN(n7274) );
  OAI211_X1 U8935 ( .C1(n9376), .C2(n7403), .A(n7274), .B(n7273), .ZN(P1_U3325) );
  INV_X1 U8936 ( .A(n7275), .ZN(n8413) );
  NOR2_X1 U8937 ( .A1(n8368), .A2(n8413), .ZN(n8150) );
  AOI21_X1 U8938 ( .B1(n8368), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8150), .ZN(
        n7277) );
  NAND2_X1 U8939 ( .A1(n7631), .A2(n8359), .ZN(n7276) );
  OAI211_X1 U8940 ( .C1(n7278), .C2(n8167), .A(n7277), .B(n7276), .ZN(P2_U3265) );
  INV_X1 U8941 ( .A(n7279), .ZN(n7281) );
  NAND2_X1 U8942 ( .A1(n7281), .A2(n7280), .ZN(n7282) );
  XNOR2_X1 U8943 ( .A(n7283), .B(n7282), .ZN(n7290) );
  NAND2_X1 U8944 ( .A1(n8666), .A2(n9826), .ZN(n7285) );
  OAI211_X1 U8945 ( .C1(n6379), .C2(n8663), .A(n7285), .B(n7284), .ZN(n7287)
         );
  NOR2_X1 U8946 ( .A1(n8668), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n7286) );
  AOI211_X1 U8947 ( .C1(n8670), .C2(n7288), .A(n7287), .B(n7286), .ZN(n7289)
         );
  OAI21_X1 U8948 ( .B1(n7290), .B2(n8672), .A(n7289), .ZN(P1_U3216) );
  NAND2_X1 U8949 ( .A1(n7291), .A2(n8767), .ZN(n7294) );
  OR2_X1 U8950 ( .A1(n6067), .A2(n7292), .ZN(n7293) );
  AND2_X1 U8951 ( .A1(P1_REG3_REG_20__SCAN_IN), .A2(P1_REG3_REG_19__SCAN_IN), 
        .ZN(n7295) );
  NAND2_X1 U8952 ( .A1(n7366), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n7368) );
  INV_X1 U8953 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n8631) );
  NAND2_X1 U8954 ( .A1(n7368), .A2(n8631), .ZN(n7296) );
  NAND2_X1 U8955 ( .A1(n7385), .A2(n7296), .ZN(n8635) );
  OR2_X1 U8956 ( .A1(n8635), .A2(n5933), .ZN(n7299) );
  AOI22_X1 U8957 ( .A1(n6081), .A2(P1_REG1_REG_22__SCAN_IN), .B1(n7555), .B2(
        P1_REG0_REG_22__SCAN_IN), .ZN(n7298) );
  NAND2_X1 U8958 ( .A1(n5931), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n7297) );
  INV_X1 U8959 ( .A(n9006), .ZN(n9150) );
  AND2_X1 U8960 ( .A1(n9007), .A2(n9150), .ZN(n8817) );
  NAND2_X1 U8961 ( .A1(n7303), .A2(n8767), .ZN(n7306) );
  AOI22_X1 U8962 ( .A1(n7338), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n9688), .B2(
        n7304), .ZN(n7305) );
  NOR2_X1 U8963 ( .A1(n9335), .A2(n8933), .ZN(n7307) );
  INV_X1 U8964 ( .A(n8933), .ZN(n9235) );
  NAND2_X1 U8965 ( .A1(n7308), .A2(n8767), .ZN(n7310) );
  AOI22_X1 U8966 ( .A1(n7338), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n9688), .B2(
        n8952), .ZN(n7309) );
  NAND2_X1 U8967 ( .A1(n6081), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n7317) );
  INV_X1 U8968 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n9225) );
  OR2_X1 U8969 ( .A1(n7598), .A2(n9225), .ZN(n7316) );
  OR2_X1 U8970 ( .A1(n7311), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n7312) );
  NAND2_X1 U8971 ( .A1(n7323), .A2(n7312), .ZN(n9224) );
  OR2_X1 U8972 ( .A1(n5933), .A2(n9224), .ZN(n7315) );
  INV_X1 U8973 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n7313) );
  OR2_X1 U8974 ( .A1(n7600), .A2(n7313), .ZN(n7314) );
  OR2_X1 U8975 ( .A1(n9330), .A2(n9244), .ZN(n8862) );
  NAND2_X1 U8976 ( .A1(n9330), .A2(n9244), .ZN(n8822) );
  INV_X1 U8977 ( .A(n9244), .ZN(n8932) );
  NAND2_X1 U8978 ( .A1(n7318), .A2(n8767), .ZN(n7320) );
  AOI22_X1 U8979 ( .A1(n7338), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n9688), .B2(
        n8969), .ZN(n7319) );
  NAND2_X1 U8980 ( .A1(n7555), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n7329) );
  INV_X1 U8981 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n7321) );
  OR2_X1 U8982 ( .A1(n4315), .A2(n7321), .ZN(n7328) );
  NAND2_X1 U8983 ( .A1(n7323), .A2(n7322), .ZN(n7324) );
  NAND2_X1 U8984 ( .A1(n7325), .A2(n7324), .ZN(n9210) );
  OR2_X1 U8985 ( .A1(n5933), .A2(n9210), .ZN(n7327) );
  INV_X1 U8986 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n9211) );
  OR2_X1 U8987 ( .A1(n7598), .A2(n9211), .ZN(n7326) );
  NAND4_X1 U8988 ( .A1(n7329), .A2(n7328), .A3(n7327), .A4(n7326), .ZN(n9193)
         );
  NAND2_X1 U8989 ( .A1(n9325), .A2(n9193), .ZN(n7331) );
  NOR2_X1 U8990 ( .A1(n9325), .A2(n9193), .ZN(n7330) );
  NAND2_X1 U8991 ( .A1(n7332), .A2(n8767), .ZN(n7334) );
  AOI22_X1 U8992 ( .A1(n7338), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n9688), .B2(
        n8979), .ZN(n7333) );
  OR2_X1 U8993 ( .A1(n9318), .A2(n9217), .ZN(n8684) );
  NAND2_X1 U8994 ( .A1(n9196), .A2(n9195), .ZN(n9316) );
  NAND2_X1 U8995 ( .A1(n7337), .A2(n8767), .ZN(n7340) );
  AOI22_X1 U8996 ( .A1(n7338), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9840), .B2(
        n9688), .ZN(n7339) );
  INV_X1 U8997 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n7341) );
  XNOR2_X1 U8998 ( .A(n7354), .B(n7341), .ZN(n9183) );
  NAND2_X1 U8999 ( .A1(n9183), .A2(n7554), .ZN(n7346) );
  NAND2_X1 U9000 ( .A1(n6081), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n7345) );
  NAND2_X1 U9001 ( .A1(n7555), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n7344) );
  INV_X1 U9002 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n7342) );
  OR2_X1 U9003 ( .A1(n7598), .A2(n7342), .ZN(n7343) );
  NAND4_X1 U9004 ( .A1(n7346), .A2(n7345), .A3(n7344), .A4(n7343), .ZN(n9192)
         );
  NAND2_X1 U9005 ( .A1(n7348), .A2(n7347), .ZN(n7349) );
  NAND2_X1 U9006 ( .A1(n7350), .A2(n8767), .ZN(n7353) );
  OR2_X1 U9007 ( .A1(n6067), .A2(n7351), .ZN(n7352) );
  AOI21_X1 U9008 ( .B1(n7354), .B2(P1_REG3_REG_19__SCAN_IN), .A(
        P1_REG3_REG_20__SCAN_IN), .ZN(n7355) );
  OR2_X1 U9009 ( .A1(n7366), .A2(n7355), .ZN(n9162) );
  INV_X1 U9010 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n7356) );
  OAI22_X1 U9011 ( .A1(n9162), .A2(n5933), .B1(n7598), .B2(n7356), .ZN(n7360)
         );
  INV_X1 U9012 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n7358) );
  NAND2_X1 U9013 ( .A1(n7555), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n7357) );
  OAI21_X1 U9014 ( .B1(n6044), .B2(n7358), .A(n7357), .ZN(n7359) );
  NAND2_X1 U9015 ( .A1(n9306), .A2(n9149), .ZN(n9141) );
  NAND2_X1 U9016 ( .A1(n7362), .A2(n8767), .ZN(n7365) );
  OR2_X1 U9017 ( .A1(n6067), .A2(n7363), .ZN(n7364) );
  OR2_X1 U9018 ( .A1(n7366), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n7367) );
  AND2_X1 U9019 ( .A1(n7368), .A2(n7367), .ZN(n9153) );
  NAND2_X1 U9020 ( .A1(n9153), .A2(n7554), .ZN(n7373) );
  NAND2_X1 U9021 ( .A1(n6081), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n7370) );
  NAND2_X1 U9022 ( .A1(n5931), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n7369) );
  AND2_X1 U9023 ( .A1(n7370), .A2(n7369), .ZN(n7372) );
  NAND2_X1 U9024 ( .A1(n7555), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n7371) );
  INV_X1 U9025 ( .A(n8632), .ZN(n9168) );
  NAND2_X1 U9026 ( .A1(n9302), .A2(n9168), .ZN(n7374) );
  AND2_X1 U9027 ( .A1(n9141), .A2(n7374), .ZN(n9001) );
  NAND2_X1 U9028 ( .A1(n9005), .A2(n9001), .ZN(n7376) );
  INV_X1 U9029 ( .A(n7374), .ZN(n7375) );
  NAND2_X1 U9030 ( .A1(n9302), .A2(n8632), .ZN(n8736) );
  NAND2_X1 U9031 ( .A1(n8816), .A2(n8736), .ZN(n9142) );
  AND2_X1 U9032 ( .A1(n7376), .A2(n9002), .ZN(n7377) );
  XOR2_X1 U9033 ( .A(n8799), .B(n7377), .Z(n9300) );
  AOI21_X1 U9034 ( .B1(n9296), .B2(n9152), .A(n9128), .ZN(n9297) );
  INV_X1 U9035 ( .A(n8635), .ZN(n7378) );
  AOI22_X1 U9036 ( .A1(n9844), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n7378), .B2(
        n9838), .ZN(n7379) );
  OAI21_X1 U9037 ( .B1(n9007), .B2(n9808), .A(n7379), .ZN(n7395) );
  INV_X1 U9038 ( .A(n8716), .ZN(n7380) );
  NOR2_X2 U9039 ( .A1(n7381), .A2(n7380), .ZN(n9239) );
  OR2_X1 U9040 ( .A1(n9335), .A2(n9235), .ZN(n8861) );
  NAND2_X1 U9041 ( .A1(n9335), .A2(n9235), .ZN(n9229) );
  INV_X1 U9042 ( .A(n9193), .ZN(n9234) );
  NAND2_X1 U9043 ( .A1(n9325), .A2(n9234), .ZN(n8823) );
  OR2_X1 U9044 ( .A1(n9325), .A2(n9234), .ZN(n9189) );
  AND2_X1 U9045 ( .A1(n8684), .A2(n9189), .ZN(n8811) );
  INV_X1 U9046 ( .A(n8825), .ZN(n7382) );
  AOI21_X1 U9047 ( .B1(n9190), .B2(n8811), .A(n7382), .ZN(n9177) );
  OR2_X1 U9048 ( .A1(n9313), .A2(n7347), .ZN(n8726) );
  NAND2_X1 U9049 ( .A1(n9313), .A2(n7347), .ZN(n8812) );
  NAND2_X1 U9050 ( .A1(n8726), .A2(n8812), .ZN(n9176) );
  NOR2_X1 U9051 ( .A1(n9177), .A2(n9176), .ZN(n9175) );
  INV_X1 U9052 ( .A(n8812), .ZN(n8820) );
  NOR2_X2 U9053 ( .A1(n9175), .A2(n8820), .ZN(n9167) );
  INV_X1 U9054 ( .A(n9149), .ZN(n9179) );
  NAND2_X1 U9055 ( .A1(n9306), .A2(n9179), .ZN(n8779) );
  NAND2_X1 U9056 ( .A1(n9167), .A2(n8779), .ZN(n9145) );
  INV_X1 U9057 ( .A(n9142), .ZN(n9147) );
  NAND3_X1 U9058 ( .A1(n9145), .A2(n9147), .A3(n9144), .ZN(n9146) );
  NAND2_X1 U9059 ( .A1(n9146), .A2(n8736), .ZN(n7383) );
  NAND2_X1 U9060 ( .A1(n7383), .A2(n8799), .ZN(n9026) );
  OAI21_X1 U9061 ( .B1(n8799), .B2(n7383), .A(n9026), .ZN(n7393) );
  INV_X1 U9062 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n7384) );
  NAND2_X1 U9063 ( .A1(n7385), .A2(n7384), .ZN(n7386) );
  AND2_X1 U9064 ( .A1(n7514), .A2(n7386), .ZN(n9131) );
  NAND2_X1 U9065 ( .A1(n9131), .A2(n7554), .ZN(n7392) );
  INV_X1 U9066 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n7389) );
  NAND2_X1 U9067 ( .A1(n7555), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n7388) );
  NAND2_X1 U9068 ( .A1(n5931), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n7387) );
  OAI211_X1 U9069 ( .C1(n6044), .C2(n7389), .A(n7388), .B(n7387), .ZN(n7390)
         );
  INV_X1 U9070 ( .A(n7390), .ZN(n7391) );
  NAND2_X1 U9071 ( .A1(n7392), .A2(n7391), .ZN(n9010) );
  AOI222_X1 U9072 ( .A1(n9823), .A2(n7393), .B1(n9010), .B2(n9828), .C1(n9168), 
        .C2(n9825), .ZN(n9299) );
  NOR2_X1 U9073 ( .A1(n9299), .A2(n9844), .ZN(n7394) );
  AOI211_X1 U9074 ( .C1(n9297), .C2(n9794), .A(n7395), .B(n7394), .ZN(n7396)
         );
  OAI21_X1 U9075 ( .B1(n9300), .B2(n9256), .A(n7396), .ZN(P1_U3269) );
  INV_X1 U9076 ( .A(n7402), .ZN(n7398) );
  OAI222_X1 U9077 ( .A1(n8534), .A2(n7399), .B1(n7939), .B2(n7398), .C1(n7397), 
        .C2(P2_U3152), .ZN(P2_U3330) );
  INV_X1 U9078 ( .A(n8768), .ZN(n9372) );
  OAI222_X1 U9079 ( .A1(n7400), .A2(P2_U3152), .B1(n7939), .B2(n9372), .C1(
        n7401), .C2(n8534), .ZN(P2_U3329) );
  NAND2_X1 U9080 ( .A1(n7402), .A2(n8767), .ZN(n7405) );
  OR2_X1 U9081 ( .A1(n6067), .A2(n7403), .ZN(n7404) );
  NAND2_X1 U9082 ( .A1(n9061), .A2(n7579), .ZN(n7415) );
  NAND2_X1 U9083 ( .A1(n7555), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n7413) );
  INV_X1 U9084 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n7406) );
  OR2_X1 U9085 ( .A1(n6044), .A2(n7406), .ZN(n7412) );
  INV_X1 U9086 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n8608) );
  NAND2_X1 U9087 ( .A1(n7551), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n7552) );
  NAND2_X1 U9088 ( .A1(n7407), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n9039) );
  INV_X1 U9089 ( .A(n7407), .ZN(n7408) );
  INV_X1 U9090 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n7605) );
  NAND2_X1 U9091 ( .A1(n7408), .A2(n7605), .ZN(n7409) );
  NAND2_X1 U9092 ( .A1(n9039), .A2(n7409), .ZN(n9058) );
  OR2_X1 U9093 ( .A1(n5933), .A2(n9058), .ZN(n7411) );
  INV_X1 U9094 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n9059) );
  OR2_X1 U9095 ( .A1(n7598), .A2(n9059), .ZN(n7410) );
  OR2_X1 U9096 ( .A1(n8758), .A2(n6049), .ZN(n7414) );
  NAND2_X1 U9097 ( .A1(n7415), .A2(n7414), .ZN(n7416) );
  XNOR2_X1 U9098 ( .A(n7416), .B(n5923), .ZN(n7418) );
  AOI22_X1 U9099 ( .A1(n9061), .A2(n7568), .B1(n7566), .B2(n9075), .ZN(n7417)
         );
  XNOR2_X1 U9100 ( .A(n7418), .B(n7417), .ZN(n7609) );
  INV_X1 U9101 ( .A(n7609), .ZN(n7419) );
  NAND2_X1 U9102 ( .A1(n7419), .A2(n8597), .ZN(n7615) );
  INV_X1 U9103 ( .A(n7423), .ZN(n7421) );
  NAND2_X1 U9104 ( .A1(n7421), .A2(n7420), .ZN(n7434) );
  NAND2_X1 U9105 ( .A1(n7436), .A2(n7434), .ZN(n7430) );
  AND2_X1 U9106 ( .A1(n7423), .A2(n7422), .ZN(n7435) );
  INV_X1 U9107 ( .A(n7435), .ZN(n7428) );
  NAND2_X1 U9108 ( .A1(n9335), .A2(n7579), .ZN(n7425) );
  NAND2_X1 U9109 ( .A1(n8933), .A2(n7568), .ZN(n7424) );
  NAND2_X1 U9110 ( .A1(n7425), .A2(n7424), .ZN(n7426) );
  XNOR2_X1 U9111 ( .A(n7426), .B(n5923), .ZN(n7433) );
  INV_X1 U9112 ( .A(n7433), .ZN(n7427) );
  AND2_X1 U9113 ( .A1(n7428), .A2(n7427), .ZN(n7429) );
  NAND2_X1 U9114 ( .A1(n7430), .A2(n7429), .ZN(n8659) );
  NAND2_X1 U9115 ( .A1(n9335), .A2(n7592), .ZN(n7432) );
  NAND2_X1 U9116 ( .A1(n8933), .A2(n7566), .ZN(n7431) );
  NAND2_X1 U9117 ( .A1(n7432), .A2(n7431), .ZN(n8662) );
  NAND2_X1 U9118 ( .A1(n8659), .A2(n8662), .ZN(n7437) );
  NAND2_X1 U9119 ( .A1(n7437), .A2(n8660), .ZN(n8585) );
  NAND2_X1 U9120 ( .A1(n9330), .A2(n7579), .ZN(n7439) );
  OR2_X1 U9121 ( .A1(n9244), .A2(n6049), .ZN(n7438) );
  NAND2_X1 U9122 ( .A1(n7439), .A2(n7438), .ZN(n7440) );
  XNOR2_X1 U9123 ( .A(n7440), .B(n5923), .ZN(n7444) );
  NAND2_X1 U9124 ( .A1(n9330), .A2(n7592), .ZN(n7442) );
  OR2_X1 U9125 ( .A1(n9244), .A2(n7590), .ZN(n7441) );
  NAND2_X1 U9126 ( .A1(n7442), .A2(n7441), .ZN(n7445) );
  INV_X1 U9127 ( .A(n7444), .ZN(n7447) );
  INV_X1 U9128 ( .A(n7445), .ZN(n7446) );
  NAND2_X1 U9129 ( .A1(n7447), .A2(n7446), .ZN(n8586) );
  NAND2_X1 U9130 ( .A1(n9325), .A2(n7579), .ZN(n7449) );
  NAND2_X1 U9131 ( .A1(n9193), .A2(n7592), .ZN(n7448) );
  NAND2_X1 U9132 ( .A1(n7449), .A2(n7448), .ZN(n7450) );
  XNOR2_X1 U9133 ( .A(n7450), .B(n5923), .ZN(n7452) );
  AND2_X1 U9134 ( .A1(n9193), .A2(n7566), .ZN(n7451) );
  AOI21_X1 U9135 ( .B1(n9325), .B2(n7568), .A(n7451), .ZN(n7453) );
  XNOR2_X1 U9136 ( .A(n7452), .B(n7453), .ZN(n8596) );
  INV_X1 U9137 ( .A(n7452), .ZN(n7454) );
  NAND2_X1 U9138 ( .A1(n7454), .A2(n7453), .ZN(n7455) );
  NAND2_X1 U9139 ( .A1(n9318), .A2(n7579), .ZN(n7457) );
  OR2_X1 U9140 ( .A1(n9217), .A2(n6049), .ZN(n7456) );
  NAND2_X1 U9141 ( .A1(n7457), .A2(n7456), .ZN(n7458) );
  XNOR2_X1 U9142 ( .A(n7458), .B(n7564), .ZN(n8640) );
  NOR2_X1 U9143 ( .A1(n9217), .A2(n7590), .ZN(n7459) );
  AOI21_X1 U9144 ( .B1(n9318), .B2(n7592), .A(n7459), .ZN(n8639) );
  NAND2_X1 U9145 ( .A1(n9313), .A2(n7579), .ZN(n7461) );
  NAND2_X1 U9146 ( .A1(n9192), .A2(n7592), .ZN(n7460) );
  NAND2_X1 U9147 ( .A1(n7461), .A2(n7460), .ZN(n7462) );
  XNOR2_X1 U9148 ( .A(n7462), .B(n7564), .ZN(n8560) );
  AND2_X1 U9149 ( .A1(n9192), .A2(n7566), .ZN(n7463) );
  AOI21_X1 U9150 ( .B1(n9313), .B2(n7568), .A(n7463), .ZN(n8559) );
  INV_X1 U9151 ( .A(n8560), .ZN(n7465) );
  INV_X1 U9152 ( .A(n8559), .ZN(n7464) );
  NAND2_X1 U9153 ( .A1(n9306), .A2(n7579), .ZN(n7467) );
  NAND2_X1 U9154 ( .A1(n9149), .A2(n7592), .ZN(n7466) );
  NAND2_X1 U9155 ( .A1(n7467), .A2(n7466), .ZN(n7468) );
  XNOR2_X1 U9156 ( .A(n7468), .B(n5923), .ZN(n7480) );
  NAND2_X1 U9157 ( .A1(n9306), .A2(n7568), .ZN(n7470) );
  NAND2_X1 U9158 ( .A1(n9149), .A2(n7566), .ZN(n7469) );
  NAND2_X1 U9159 ( .A1(n7470), .A2(n7469), .ZN(n7481) );
  NAND2_X1 U9160 ( .A1(n7480), .A2(n7481), .ZN(n8617) );
  NAND2_X1 U9161 ( .A1(n9302), .A2(n7579), .ZN(n7472) );
  OR2_X1 U9162 ( .A1(n8632), .A2(n6049), .ZN(n7471) );
  NAND2_X1 U9163 ( .A1(n7472), .A2(n7471), .ZN(n7473) );
  XNOR2_X1 U9164 ( .A(n7473), .B(n5923), .ZN(n7477) );
  INV_X1 U9165 ( .A(n7477), .ZN(n7475) );
  NOR2_X1 U9166 ( .A1(n8632), .A2(n7590), .ZN(n7474) );
  AOI21_X1 U9167 ( .B1(n9302), .B2(n7568), .A(n7474), .ZN(n7476) );
  NAND2_X1 U9168 ( .A1(n7475), .A2(n7476), .ZN(n7484) );
  INV_X1 U9169 ( .A(n7484), .ZN(n7478) );
  XNOR2_X1 U9170 ( .A(n7477), .B(n7476), .ZN(n8568) );
  AND2_X1 U9171 ( .A1(n8617), .A2(n7501), .ZN(n7479) );
  NAND2_X1 U9172 ( .A1(n8616), .A2(n7479), .ZN(n7487) );
  INV_X1 U9173 ( .A(n7501), .ZN(n7485) );
  INV_X1 U9174 ( .A(n7480), .ZN(n7483) );
  INV_X1 U9175 ( .A(n7481), .ZN(n7482) );
  NAND2_X1 U9176 ( .A1(n7483), .A2(n7482), .ZN(n8619) );
  AND2_X1 U9177 ( .A1(n8619), .A2(n7484), .ZN(n7500) );
  NAND2_X1 U9178 ( .A1(n7487), .A2(n7486), .ZN(n7490) );
  OR2_X1 U9179 ( .A1(n9007), .A2(n6049), .ZN(n7489) );
  NAND2_X1 U9180 ( .A1(n9150), .A2(n7566), .ZN(n7488) );
  OAI22_X1 U9181 ( .A1(n9007), .A2(n6055), .B1(n9006), .B2(n6049), .ZN(n7491)
         );
  XNOR2_X1 U9182 ( .A(n7491), .B(n5923), .ZN(n8630) );
  NAND2_X1 U9183 ( .A1(n8627), .A2(n8630), .ZN(n7506) );
  NAND2_X1 U9184 ( .A1(n7492), .A2(n8767), .ZN(n7495) );
  OR2_X1 U9185 ( .A1(n6067), .A2(n7493), .ZN(n7494) );
  NAND2_X1 U9186 ( .A1(n9291), .A2(n7579), .ZN(n7497) );
  NAND2_X1 U9187 ( .A1(n9010), .A2(n7592), .ZN(n7496) );
  NAND2_X1 U9188 ( .A1(n7497), .A2(n7496), .ZN(n7498) );
  XNOR2_X1 U9189 ( .A(n7498), .B(n7564), .ZN(n7507) );
  NAND2_X1 U9190 ( .A1(n8616), .A2(n8617), .ZN(n8615) );
  INV_X1 U9191 ( .A(n7502), .ZN(n7499) );
  AND2_X1 U9192 ( .A1(n7500), .A2(n7499), .ZN(n7503) );
  AOI21_X2 U9193 ( .B1(n8615), .B2(n7503), .A(n4819), .ZN(n8628) );
  NAND3_X1 U9194 ( .A1(n7506), .A2(n7507), .A3(n8628), .ZN(n8546) );
  NAND2_X1 U9195 ( .A1(n9291), .A2(n7568), .ZN(n7505) );
  NAND2_X1 U9196 ( .A1(n9010), .A2(n7566), .ZN(n7504) );
  NAND2_X1 U9197 ( .A1(n7505), .A2(n7504), .ZN(n8550) );
  NAND2_X1 U9198 ( .A1(n8546), .A2(n8550), .ZN(n8547) );
  NAND2_X1 U9199 ( .A1(n7506), .A2(n8628), .ZN(n7509) );
  INV_X1 U9200 ( .A(n7507), .ZN(n7508) );
  NAND2_X1 U9201 ( .A1(n8547), .A2(n8548), .ZN(n8606) );
  INV_X1 U9202 ( .A(n8606), .ZN(n8552) );
  NAND2_X1 U9203 ( .A1(n7510), .A2(n8767), .ZN(n7513) );
  OR2_X1 U9204 ( .A1(n6067), .A2(n7511), .ZN(n7512) );
  AND2_X1 U9205 ( .A1(n7514), .A2(n8608), .ZN(n7515) );
  OR2_X1 U9206 ( .A1(n7515), .A2(n7530), .ZN(n9120) );
  INV_X1 U9207 ( .A(n9120), .ZN(n7520) );
  INV_X1 U9208 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n7518) );
  NAND2_X1 U9209 ( .A1(n7555), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n7517) );
  NAND2_X1 U9210 ( .A1(n5931), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n7516) );
  OAI211_X1 U9211 ( .C1(n6044), .C2(n7518), .A(n7517), .B(n7516), .ZN(n7519)
         );
  AOI21_X1 U9212 ( .B1(n7520), .B2(n7554), .A(n7519), .ZN(n9012) );
  OAI22_X1 U9213 ( .A1(n9013), .A2(n6055), .B1(n9012), .B2(n6049), .ZN(n7521)
         );
  XNOR2_X1 U9214 ( .A(n7521), .B(n5923), .ZN(n7524) );
  OAI22_X1 U9215 ( .A1(n9013), .A2(n6049), .B1(n9012), .B2(n7590), .ZN(n7523)
         );
  XNOR2_X1 U9216 ( .A(n7524), .B(n7523), .ZN(n8607) );
  OR2_X1 U9217 ( .A1(n7524), .A2(n7523), .ZN(n7525) );
  NAND2_X1 U9218 ( .A1(n8604), .A2(n7525), .ZN(n8574) );
  NAND2_X1 U9219 ( .A1(n7526), .A2(n8767), .ZN(n7529) );
  OR2_X1 U9220 ( .A1(n6067), .A2(n7527), .ZN(n7528) );
  NAND2_X1 U9221 ( .A1(n9281), .A2(n7579), .ZN(n7539) );
  NOR2_X1 U9222 ( .A1(n7530), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n7531) );
  OR2_X1 U9223 ( .A1(n7551), .A2(n7531), .ZN(n8578) );
  INV_X1 U9224 ( .A(n8578), .ZN(n9098) );
  NAND2_X1 U9225 ( .A1(n9098), .A2(n7554), .ZN(n7537) );
  INV_X1 U9226 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n7534) );
  NAND2_X1 U9227 ( .A1(n7555), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n7533) );
  NAND2_X1 U9228 ( .A1(n5931), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n7532) );
  OAI211_X1 U9229 ( .C1(n6044), .C2(n7534), .A(n7533), .B(n7532), .ZN(n7535)
         );
  INV_X1 U9230 ( .A(n7535), .ZN(n7536) );
  INV_X1 U9231 ( .A(n9116), .ZN(n8931) );
  NAND2_X1 U9232 ( .A1(n8931), .A2(n7592), .ZN(n7538) );
  NAND2_X1 U9233 ( .A1(n7539), .A2(n7538), .ZN(n7540) );
  XNOR2_X1 U9234 ( .A(n7540), .B(n5923), .ZN(n7542) );
  NOR2_X1 U9235 ( .A1(n9116), .A2(n7590), .ZN(n7541) );
  AOI21_X1 U9236 ( .B1(n9281), .B2(n7592), .A(n7541), .ZN(n7543) );
  XNOR2_X1 U9237 ( .A(n7542), .B(n7543), .ZN(n8575) );
  NAND2_X1 U9238 ( .A1(n8574), .A2(n8575), .ZN(n7546) );
  INV_X1 U9239 ( .A(n7542), .ZN(n7544) );
  NAND2_X1 U9240 ( .A1(n7544), .A2(n7543), .ZN(n7545) );
  OR2_X1 U9241 ( .A1(n6067), .A2(n7548), .ZN(n7549) );
  NAND2_X1 U9242 ( .A1(n9278), .A2(n7579), .ZN(n7563) );
  OR2_X1 U9243 ( .A1(n7551), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n7553) );
  AND2_X1 U9244 ( .A1(n7553), .A2(n7552), .ZN(n9088) );
  NAND2_X1 U9245 ( .A1(n9088), .A2(n7554), .ZN(n7561) );
  INV_X1 U9246 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n7558) );
  NAND2_X1 U9247 ( .A1(n7555), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n7557) );
  NAND2_X1 U9248 ( .A1(n5931), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n7556) );
  OAI211_X1 U9249 ( .C1(n6044), .C2(n7558), .A(n7557), .B(n7556), .ZN(n7559)
         );
  INV_X1 U9250 ( .A(n7559), .ZN(n7560) );
  NAND2_X1 U9251 ( .A1(n7561), .A2(n7560), .ZN(n9103) );
  NAND2_X1 U9252 ( .A1(n9103), .A2(n7568), .ZN(n7562) );
  NAND2_X1 U9253 ( .A1(n7563), .A2(n7562), .ZN(n7565) );
  XNOR2_X1 U9254 ( .A(n7565), .B(n7564), .ZN(n7570) );
  AND2_X1 U9255 ( .A1(n9103), .A2(n7566), .ZN(n7567) );
  AOI21_X1 U9256 ( .B1(n9278), .B2(n7568), .A(n7567), .ZN(n7571) );
  XNOR2_X1 U9257 ( .A(n7570), .B(n7571), .ZN(n8650) );
  INV_X1 U9258 ( .A(n7570), .ZN(n7573) );
  INV_X1 U9259 ( .A(n7571), .ZN(n7572) );
  NAND2_X1 U9260 ( .A1(n7573), .A2(n7572), .ZN(n7574) );
  OR2_X1 U9261 ( .A1(n6067), .A2(n7576), .ZN(n7577) );
  NAND2_X1 U9262 ( .A1(n9271), .A2(n7579), .ZN(n7588) );
  NAND2_X1 U9263 ( .A1(n6081), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n7586) );
  INV_X1 U9264 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n7580) );
  OR2_X1 U9265 ( .A1(n7600), .A2(n7580), .ZN(n7585) );
  XNOR2_X1 U9266 ( .A(P1_REG3_REG_27__SCAN_IN), .B(n7581), .ZN(n9069) );
  OR2_X1 U9267 ( .A1(n5933), .A2(n9069), .ZN(n7584) );
  INV_X1 U9268 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n7582) );
  OR2_X1 U9269 ( .A1(n7598), .A2(n7582), .ZN(n7583) );
  OR2_X1 U9270 ( .A1(n9085), .A2(n6049), .ZN(n7587) );
  NAND2_X1 U9271 ( .A1(n7588), .A2(n7587), .ZN(n7589) );
  XNOR2_X1 U9272 ( .A(n7589), .B(n5923), .ZN(n8538) );
  NOR2_X1 U9273 ( .A1(n9085), .A2(n7590), .ZN(n7591) );
  AOI21_X1 U9274 ( .B1(n9271), .B2(n7592), .A(n7591), .ZN(n8537) );
  INV_X1 U9275 ( .A(n8537), .ZN(n7594) );
  OR2_X1 U9276 ( .A1(n8538), .A2(n7594), .ZN(n7593) );
  NAND2_X1 U9277 ( .A1(n8540), .A2(n7593), .ZN(n7614) );
  NAND2_X1 U9278 ( .A1(n8538), .A2(n7594), .ZN(n7608) );
  INV_X1 U9279 ( .A(n7608), .ZN(n7595) );
  NOR2_X1 U9280 ( .A1(n7595), .A2(n8672), .ZN(n7596) );
  AND2_X1 U9281 ( .A1(n7609), .A2(n7596), .ZN(n7597) );
  NAND2_X1 U9282 ( .A1(n7614), .A2(n7597), .ZN(n7613) );
  NAND2_X1 U9283 ( .A1(n6081), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n7604) );
  INV_X1 U9284 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n9040) );
  OR2_X1 U9285 ( .A1(n7598), .A2(n9040), .ZN(n7603) );
  OR2_X1 U9286 ( .A1(n5933), .A2(n9039), .ZN(n7602) );
  INV_X1 U9287 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n7599) );
  OR2_X1 U9288 ( .A1(n7600), .A2(n7599), .ZN(n7601) );
  INV_X1 U9289 ( .A(n8777), .ZN(n9053) );
  OAI22_X1 U9290 ( .A1(n8663), .A2(n9085), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7605), .ZN(n7606) );
  AOI21_X1 U9291 ( .B1(n8666), .B2(n9053), .A(n7606), .ZN(n7607) );
  OAI21_X1 U9292 ( .B1(n8668), .B2(n9058), .A(n7607), .ZN(n7611) );
  NOR3_X1 U9293 ( .A1(n7609), .A2(n8672), .A3(n7608), .ZN(n7610) );
  AOI211_X1 U9294 ( .C1(n8670), .C2(n9061), .A(n7611), .B(n7610), .ZN(n7612)
         );
  OAI211_X1 U9295 ( .C1(n7615), .C2(n7614), .A(n7613), .B(n7612), .ZN(P1_U3218) );
  MUX2_X1 U9296 ( .A(n7653), .B(n7618), .S(n7902), .Z(n7616) );
  AOI21_X1 U9297 ( .B1(n7617), .B2(n7616), .A(n8036), .ZN(n7620) );
  NOR2_X1 U9298 ( .A1(n8026), .A2(n7618), .ZN(n7619) );
  AOI211_X1 U9299 ( .C1(P2_REG3_REG_0__SCAN_IN), .C2(n7621), .A(n7620), .B(
        n7619), .ZN(n7622) );
  OAI21_X1 U9300 ( .B1(n7623), .B2(n8029), .A(n7622), .ZN(P2_U3234) );
  INV_X1 U9301 ( .A(n7801), .ZN(n7624) );
  INV_X1 U9302 ( .A(n7626), .ZN(n7628) );
  NAND2_X1 U9303 ( .A1(n8415), .A2(n8050), .ZN(n7810) );
  AOI21_X1 U9304 ( .B1(n8415), .B2(n7628), .A(n7627), .ZN(n7632) );
  INV_X1 U9305 ( .A(n8415), .ZN(n8149) );
  INV_X1 U9306 ( .A(n8050), .ZN(n7629) );
  NAND2_X1 U9307 ( .A1(n8149), .A2(n7629), .ZN(n7804) );
  NAND2_X1 U9308 ( .A1(n7631), .A2(n7630), .ZN(n7812) );
  OAI21_X1 U9309 ( .B1(n7632), .B2(n7848), .A(n7812), .ZN(n7633) );
  XNOR2_X1 U9310 ( .A(n7633), .B(n9946), .ZN(n7637) );
  NAND2_X1 U9311 ( .A1(n7635), .A2(n7634), .ZN(n7636) );
  AND2_X1 U9312 ( .A1(n7852), .A2(n9946), .ZN(n7638) );
  NAND2_X1 U9313 ( .A1(n5218), .A2(n7638), .ZN(n7639) );
  INV_X1 U9314 ( .A(n7660), .ZN(n7811) );
  MUX2_X1 U9315 ( .A(n8057), .B(n8505), .S(n7639), .Z(n7722) );
  NAND2_X1 U9316 ( .A1(n7646), .A2(n7645), .ZN(n7641) );
  AND2_X1 U9317 ( .A1(n7645), .A2(n7644), .ZN(n7647) );
  OAI211_X1 U9318 ( .C1(n7676), .C2(n7647), .A(n7646), .B(n7679), .ZN(n7648)
         );
  NAND2_X1 U9319 ( .A1(n7648), .A2(n7811), .ZN(n7668) );
  AND2_X1 U9320 ( .A1(n7653), .A2(n7852), .ZN(n7649) );
  OAI211_X1 U9321 ( .C1(n7650), .C2(n7649), .A(n7658), .B(n7654), .ZN(n7651)
         );
  NAND2_X1 U9322 ( .A1(n7652), .A2(n7639), .ZN(n7663) );
  NAND2_X1 U9323 ( .A1(n7654), .A2(n7653), .ZN(n7657) );
  NAND3_X1 U9324 ( .A1(n7657), .A2(n7656), .A3(n7655), .ZN(n7659) );
  NAND2_X1 U9325 ( .A1(n7659), .A2(n7658), .ZN(n7661) );
  NAND2_X1 U9326 ( .A1(n7663), .A2(n7662), .ZN(n7666) );
  INV_X1 U9327 ( .A(n7676), .ZN(n7664) );
  NAND2_X1 U9328 ( .A1(n7666), .A2(n7665), .ZN(n7667) );
  NAND2_X1 U9329 ( .A1(n7668), .A2(n7667), .ZN(n7669) );
  NAND2_X1 U9330 ( .A1(n8064), .A2(n9988), .ZN(n7673) );
  NAND2_X1 U9331 ( .A1(n7669), .A2(n7673), .ZN(n7682) );
  NAND2_X1 U9332 ( .A1(n8068), .A2(n7670), .ZN(n7671) );
  AND2_X1 U9333 ( .A1(n7672), .A2(n7671), .ZN(n7675) );
  OAI211_X1 U9334 ( .C1(n7676), .C2(n7675), .A(n7674), .B(n7673), .ZN(n7677)
         );
  NAND2_X1 U9335 ( .A1(n7677), .A2(n7660), .ZN(n7681) );
  OAI21_X1 U9336 ( .B1(n7679), .B2(n7639), .A(n7678), .ZN(n7680) );
  INV_X1 U9337 ( .A(n7683), .ZN(n7685) );
  NOR3_X1 U9338 ( .A1(n7701), .A2(n7685), .A3(n7684), .ZN(n7693) );
  INV_X1 U9339 ( .A(n7687), .ZN(n7688) );
  NOR2_X1 U9340 ( .A1(n7689), .A2(n7688), .ZN(n7690) );
  OAI21_X1 U9341 ( .B1(n7693), .B2(n7692), .A(n7691), .ZN(n7694) );
  NAND2_X1 U9342 ( .A1(n7694), .A2(n7696), .ZN(n7712) );
  NAND2_X1 U9343 ( .A1(n7705), .A2(n7695), .ZN(n7698) );
  INV_X1 U9344 ( .A(n7696), .ZN(n7697) );
  MUX2_X1 U9345 ( .A(n7698), .B(n7697), .S(n7811), .Z(n7700) );
  NOR2_X1 U9346 ( .A1(n7700), .A2(n7699), .ZN(n7711) );
  INV_X1 U9347 ( .A(n7701), .ZN(n7703) );
  NAND4_X1 U9348 ( .A1(n7703), .A2(n4816), .A3(n7711), .A4(n7702), .ZN(n7706)
         );
  NAND3_X1 U9349 ( .A1(n7706), .A2(n7705), .A3(n7704), .ZN(n7709) );
  NAND2_X1 U9350 ( .A1(n7714), .A2(n7707), .ZN(n7708) );
  AOI21_X1 U9351 ( .B1(n7712), .B2(n7711), .A(n7710), .ZN(n7718) );
  OAI21_X1 U9352 ( .B1(n7718), .B2(n7713), .A(n7715), .ZN(n7720) );
  NAND2_X1 U9353 ( .A1(n7715), .A2(n7714), .ZN(n7717) );
  OAI21_X1 U9354 ( .B1(n7718), .B2(n7717), .A(n7716), .ZN(n7719) );
  INV_X1 U9355 ( .A(n7725), .ZN(n7726) );
  MUX2_X1 U9356 ( .A(n4710), .B(n7726), .S(n7811), .Z(n7727) );
  INV_X1 U9357 ( .A(n7728), .ZN(n7733) );
  MUX2_X1 U9358 ( .A(n7730), .B(n7729), .S(n7639), .Z(n7731) );
  NAND2_X1 U9359 ( .A1(n7732), .A2(n7731), .ZN(n7743) );
  NOR3_X1 U9360 ( .A1(n7742), .A2(n7733), .A3(n7743), .ZN(n7740) );
  INV_X1 U9361 ( .A(n7734), .ZN(n7735) );
  NOR2_X1 U9362 ( .A1(n7735), .A2(n7660), .ZN(n7736) );
  NAND2_X1 U9363 ( .A1(n4820), .A2(n7736), .ZN(n7739) );
  OAI21_X1 U9364 ( .B1(n7740), .B2(n7739), .A(n7738), .ZN(n7748) );
  NOR3_X1 U9365 ( .A1(n7742), .A2(n7741), .A3(n7811), .ZN(n7746) );
  INV_X1 U9366 ( .A(n7743), .ZN(n7744) );
  OAI21_X1 U9367 ( .B1(n7746), .B2(n7745), .A(n7744), .ZN(n7747) );
  NAND2_X1 U9368 ( .A1(n7748), .A2(n7747), .ZN(n7757) );
  AOI21_X1 U9369 ( .B1(n7757), .B2(n7749), .A(n7758), .ZN(n7753) );
  NAND2_X1 U9370 ( .A1(n7761), .A2(n7750), .ZN(n7752) );
  NAND2_X1 U9371 ( .A1(n8291), .A2(n8056), .ZN(n7763) );
  OAI211_X1 U9372 ( .C1(n7753), .C2(n7752), .A(n7751), .B(n7763), .ZN(n7754)
         );
  NAND3_X1 U9373 ( .A1(n7754), .A2(n7762), .A3(n7769), .ZN(n7767) );
  AOI211_X1 U9374 ( .C1(n7757), .C2(n4820), .A(n7756), .B(n7755), .ZN(n7760)
         );
  NAND2_X1 U9375 ( .A1(n7762), .A2(n7761), .ZN(n7764) );
  OAI211_X1 U9376 ( .C1(n7765), .C2(n7764), .A(n7768), .B(n7763), .ZN(n7766)
         );
  MUX2_X1 U9377 ( .A(n7767), .B(n7766), .S(n7660), .Z(n7772) );
  MUX2_X1 U9378 ( .A(n7769), .B(n7768), .S(n7811), .Z(n7770) );
  NAND2_X1 U9379 ( .A1(n7772), .A2(n7771), .ZN(n7774) );
  INV_X1 U9380 ( .A(n8448), .ZN(n8257) );
  AOI21_X1 U9381 ( .B1(n8257), .B2(n8229), .A(n8228), .ZN(n7773) );
  NAND2_X1 U9382 ( .A1(n7777), .A2(n7775), .ZN(n7776) );
  INV_X1 U9383 ( .A(n8214), .ZN(n7778) );
  NAND2_X1 U9384 ( .A1(n7784), .A2(n7780), .ZN(n7783) );
  NAND2_X1 U9385 ( .A1(n8191), .A2(n7781), .ZN(n7782) );
  MUX2_X1 U9386 ( .A(n7783), .B(n7782), .S(n7639), .Z(n7787) );
  MUX2_X1 U9387 ( .A(n7785), .B(n7784), .S(n7811), .Z(n7786) );
  INV_X1 U9388 ( .A(n7788), .ZN(n7789) );
  NOR2_X1 U9389 ( .A1(n7794), .A2(n7789), .ZN(n7790) );
  MUX2_X1 U9390 ( .A(n7791), .B(n7790), .S(n7639), .Z(n7792) );
  NAND2_X1 U9391 ( .A1(n7793), .A2(n7792), .ZN(n7797) );
  AOI21_X1 U9392 ( .B1(n7797), .B2(n8182), .A(n7796), .ZN(n7798) );
  NOR2_X1 U9393 ( .A1(n7800), .A2(n7799), .ZN(n7807) );
  MUX2_X1 U9394 ( .A(n7802), .B(n7801), .S(n7639), .Z(n7803) );
  INV_X1 U9395 ( .A(n7803), .ZN(n7806) );
  OAI21_X1 U9396 ( .B1(n7807), .B2(n7806), .A(n7805), .ZN(n7808) );
  OAI21_X1 U9397 ( .B1(n7809), .B2(n7811), .A(n7808), .ZN(n7813) );
  NAND2_X1 U9398 ( .A1(n7812), .A2(n7810), .ZN(n7847) );
  NOR2_X1 U9399 ( .A1(n7814), .A2(n7660), .ZN(n7815) );
  INV_X1 U9400 ( .A(n7850), .ZN(n7816) );
  NOR2_X1 U9401 ( .A1(n7816), .A2(n9964), .ZN(n7817) );
  INV_X1 U9402 ( .A(n8261), .ZN(n7843) );
  INV_X1 U9403 ( .A(n8397), .ZN(n7836) );
  NOR4_X1 U9404 ( .A1(n7820), .A2(n9965), .A3(n7819), .A4(n7818), .ZN(n7823)
         );
  NAND3_X1 U9405 ( .A1(n7823), .A2(n7822), .A3(n7821), .ZN(n7827) );
  NOR4_X1 U9406 ( .A1(n7827), .A2(n7826), .A3(n7825), .A4(n7824), .ZN(n7829)
         );
  NAND4_X1 U9407 ( .A1(n7829), .A2(n4816), .A3(n7828), .A4(n5491), .ZN(n7832)
         );
  NOR4_X1 U9408 ( .A1(n7833), .A2(n7832), .A3(n7831), .A4(n7830), .ZN(n7835)
         );
  NAND4_X1 U9409 ( .A1(n8375), .A2(n7836), .A3(n7835), .A4(n7834), .ZN(n7837)
         );
  NOR4_X1 U9410 ( .A1(n7838), .A2(n8332), .A3(n8352), .A4(n7837), .ZN(n7840)
         );
  NAND4_X1 U9411 ( .A1(n8265), .A2(n7841), .A3(n7840), .A4(n7839), .ZN(n7842)
         );
  NOR4_X1 U9412 ( .A1(n8213), .A2(n8228), .A3(n7843), .A4(n7842), .ZN(n7844)
         );
  NAND4_X1 U9413 ( .A1(n8155), .A2(n8191), .A3(n8172), .A4(n7844), .ZN(n7845)
         );
  XNOR2_X1 U9414 ( .A(n7849), .B(n9946), .ZN(n7853) );
  OAI22_X1 U9415 ( .A1(n7853), .A2(n7852), .B1(n7851), .B2(n7850), .ZN(n7854)
         );
  INV_X1 U9416 ( .A(n4994), .ZN(n7858) );
  NAND4_X1 U9417 ( .A1(n7859), .A2(n7858), .A3(n7857), .A4(n8390), .ZN(n7860)
         );
  OAI211_X1 U9418 ( .C1(n7862), .C2(n7861), .A(n7860), .B(P2_B_REG_SCAN_IN), 
        .ZN(n7863) );
  OAI222_X1 U9419 ( .A1(n8534), .A2(n7865), .B1(n7939), .B2(n7864), .C1(
        P2_U3152), .C2(n5218), .ZN(P2_U3336) );
  NOR2_X1 U9420 ( .A1(n8248), .A2(n7902), .ZN(n8001) );
  XOR2_X1 U9421 ( .A(n7926), .B(n8442), .Z(n8002) );
  INV_X1 U9422 ( .A(n8002), .ZN(n7907) );
  XNOR2_X1 U9423 ( .A(n8484), .B(n7921), .ZN(n7870) );
  NAND2_X1 U9424 ( .A1(n8393), .A2(n7635), .ZN(n7871) );
  NAND2_X1 U9425 ( .A1(n7870), .A2(n7871), .ZN(n7986) );
  INV_X1 U9426 ( .A(n7870), .ZN(n7873) );
  INV_X1 U9427 ( .A(n7871), .ZN(n7872) );
  NAND2_X1 U9428 ( .A1(n7873), .A2(n7872), .ZN(n7874) );
  XNOR2_X1 U9429 ( .A(n8480), .B(n7921), .ZN(n7879) );
  INV_X1 U9430 ( .A(n7879), .ZN(n7876) );
  NAND2_X1 U9431 ( .A1(n8372), .A2(n7635), .ZN(n7878) );
  INV_X1 U9432 ( .A(n7878), .ZN(n7875) );
  NAND2_X1 U9433 ( .A1(n7876), .A2(n7875), .ZN(n7877) );
  AND2_X1 U9434 ( .A1(n7979), .A2(n7877), .ZN(n7883) );
  INV_X1 U9435 ( .A(n7877), .ZN(n7882) );
  XNOR2_X1 U9436 ( .A(n7879), .B(n7878), .ZN(n7988) );
  INV_X1 U9437 ( .A(n7988), .ZN(n7880) );
  AND2_X1 U9438 ( .A1(n7880), .A2(n7986), .ZN(n7881) );
  XNOR2_X1 U9439 ( .A(n8474), .B(n7926), .ZN(n7886) );
  NAND2_X1 U9440 ( .A1(n8318), .A2(n7635), .ZN(n7884) );
  XNOR2_X1 U9441 ( .A(n7886), .B(n7884), .ZN(n8027) );
  INV_X1 U9442 ( .A(n7884), .ZN(n7885) );
  AND2_X1 U9443 ( .A1(n7886), .A2(n7885), .ZN(n7887) );
  XNOR2_X1 U9444 ( .A(n8471), .B(n7921), .ZN(n7888) );
  NAND2_X1 U9445 ( .A1(n8341), .A2(n7635), .ZN(n7889) );
  NAND2_X1 U9446 ( .A1(n7888), .A2(n7889), .ZN(n7893) );
  INV_X1 U9447 ( .A(n7888), .ZN(n7891) );
  INV_X1 U9448 ( .A(n7889), .ZN(n7890) );
  NAND2_X1 U9449 ( .A1(n7891), .A2(n7890), .ZN(n7892) );
  AND2_X1 U9450 ( .A1(n7893), .A2(n7892), .ZN(n7953) );
  XNOR2_X1 U9451 ( .A(n8302), .B(n7926), .ZN(n7894) );
  NAND2_X1 U9452 ( .A1(n8319), .A2(n7635), .ZN(n7895) );
  XNOR2_X1 U9453 ( .A(n7894), .B(n7895), .ZN(n8011) );
  XNOR2_X1 U9454 ( .A(n8459), .B(n7921), .ZN(n7899) );
  NOR2_X1 U9455 ( .A1(n8308), .A2(n7902), .ZN(n7900) );
  XNOR2_X1 U9456 ( .A(n7899), .B(n7900), .ZN(n7964) );
  INV_X1 U9457 ( .A(n7964), .ZN(n7898) );
  INV_X1 U9458 ( .A(n7894), .ZN(n7897) );
  INV_X1 U9459 ( .A(n7895), .ZN(n7896) );
  NAND2_X1 U9460 ( .A1(n7897), .A2(n7896), .ZN(n7962) );
  INV_X1 U9461 ( .A(n7899), .ZN(n7901) );
  XNOR2_X1 U9462 ( .A(n8454), .B(n7921), .ZN(n7903) );
  XNOR2_X1 U9463 ( .A(n7905), .B(n7903), .ZN(n8019) );
  OR2_X1 U9464 ( .A1(n8247), .A2(n7902), .ZN(n8018) );
  INV_X1 U9465 ( .A(n7903), .ZN(n7904) );
  OAI21_X1 U9466 ( .B1(n8001), .B2(n7907), .A(n7997), .ZN(n7910) );
  INV_X1 U9467 ( .A(n8001), .ZN(n7908) );
  OR2_X1 U9468 ( .A1(n8002), .A2(n7908), .ZN(n7909) );
  NAND2_X1 U9469 ( .A1(n8229), .A2(n7635), .ZN(n7999) );
  NAND2_X1 U9470 ( .A1(n7913), .A2(n7912), .ZN(n7914) );
  XNOR2_X1 U9471 ( .A(n8439), .B(n7926), .ZN(n7916) );
  NAND2_X1 U9472 ( .A1(n8230), .A2(n7635), .ZN(n7971) );
  XNOR2_X1 U9473 ( .A(n8433), .B(n7921), .ZN(n7919) );
  NAND2_X1 U9474 ( .A1(n8053), .A2(n7635), .ZN(n7918) );
  NOR2_X1 U9475 ( .A1(n7919), .A2(n7918), .ZN(n7920) );
  AOI21_X1 U9476 ( .B1(n7919), .B2(n7918), .A(n7920), .ZN(n8040) );
  XNOR2_X1 U9477 ( .A(n8427), .B(n7921), .ZN(n7923) );
  NAND2_X1 U9478 ( .A1(n8052), .A2(n7635), .ZN(n7922) );
  NOR2_X1 U9479 ( .A1(n7923), .A2(n7922), .ZN(n7924) );
  AOI21_X1 U9480 ( .B1(n7923), .B2(n7922), .A(n7924), .ZN(n7941) );
  NAND2_X1 U9481 ( .A1(n7942), .A2(n7941), .ZN(n7940) );
  INV_X1 U9482 ( .A(n7924), .ZN(n7925) );
  NAND2_X1 U9483 ( .A1(n7940), .A2(n7925), .ZN(n7930) );
  NAND2_X1 U9484 ( .A1(n8051), .A2(n7635), .ZN(n7927) );
  XNOR2_X1 U9485 ( .A(n7927), .B(n7926), .ZN(n7928) );
  XNOR2_X1 U9486 ( .A(n8422), .B(n7928), .ZN(n7929) );
  XNOR2_X1 U9487 ( .A(n7930), .B(n7929), .ZN(n7936) );
  INV_X1 U9488 ( .A(n8164), .ZN(n7932) );
  OAI22_X1 U9489 ( .A1(n7932), .A2(n8045), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7931), .ZN(n7934) );
  OAI22_X1 U9490 ( .A1(n8158), .A2(n8029), .B1(n8157), .B2(n8030), .ZN(n7933)
         );
  AOI211_X1 U9491 ( .C1(n8422), .C2(n8047), .A(n7934), .B(n7933), .ZN(n7935)
         );
  OAI21_X1 U9492 ( .B1(n7936), .B2(n8036), .A(n7935), .ZN(P2_U3222) );
  INV_X1 U9493 ( .A(n8677), .ZN(n9370) );
  OAI222_X1 U9494 ( .A1(P2_U3152), .A2(n7937), .B1(n7939), .B2(n9370), .C1(
        n7938), .C2(n8534), .ZN(P2_U3328) );
  OAI211_X1 U9495 ( .C1(n7942), .C2(n7941), .A(n7940), .B(n8038), .ZN(n7946)
         );
  OAI22_X1 U9496 ( .A1(n8175), .A2(n8045), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9536), .ZN(n7944) );
  OAI22_X1 U9497 ( .A1(n8182), .A2(n8029), .B1(n8181), .B2(n8030), .ZN(n7943)
         );
  AOI211_X1 U9498 ( .C1(n8427), .C2(n8047), .A(n7944), .B(n7943), .ZN(n7945)
         );
  NAND2_X1 U9499 ( .A1(n7946), .A2(n7945), .ZN(P2_U3216) );
  XNOR2_X1 U9500 ( .A(n8000), .B(n7999), .ZN(n7951) );
  OAI22_X1 U9501 ( .A1(n8045), .A2(n8254), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7947), .ZN(n7949) );
  OAI22_X1 U9502 ( .A1(n8248), .A2(n8029), .B1(n8030), .B2(n8247), .ZN(n7948)
         );
  AOI211_X1 U9503 ( .C1(n8448), .C2(n8047), .A(n7949), .B(n7948), .ZN(n7950)
         );
  OAI21_X1 U9504 ( .B1(n7951), .B2(n8036), .A(n7950), .ZN(P2_U3218) );
  INV_X1 U9505 ( .A(n8471), .ZN(n7961) );
  OAI21_X1 U9506 ( .B1(n7954), .B2(n7953), .A(n7952), .ZN(n7955) );
  NAND2_X1 U9507 ( .A1(n7955), .A2(n8038), .ZN(n7960) );
  INV_X1 U9508 ( .A(n8326), .ZN(n7958) );
  AND2_X1 U9509 ( .A1(P2_U3152), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8144) );
  OAI22_X1 U9510 ( .A1(n7956), .A2(n8030), .B1(n8029), .B2(n7966), .ZN(n7957)
         );
  AOI211_X1 U9511 ( .C1(n8033), .C2(n7958), .A(n8144), .B(n7957), .ZN(n7959)
         );
  OAI211_X1 U9512 ( .C1(n7961), .C2(n8026), .A(n7960), .B(n7959), .ZN(P2_U3221) );
  OR2_X1 U9513 ( .A1(n8012), .A2(n8011), .ZN(n7963) );
  NAND2_X1 U9514 ( .A1(n7963), .A2(n7962), .ZN(n7965) );
  XNOR2_X1 U9515 ( .A(n7965), .B(n7964), .ZN(n7970) );
  OAI22_X1 U9516 ( .A1(n8045), .A2(n8288), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9455), .ZN(n7968) );
  OAI22_X1 U9517 ( .A1(n7966), .A2(n8030), .B1(n8029), .B2(n8247), .ZN(n7967)
         );
  AOI211_X1 U9518 ( .C1(n8459), .C2(n8047), .A(n7968), .B(n7967), .ZN(n7969)
         );
  OAI21_X1 U9519 ( .B1(n7970), .B2(n8036), .A(n7969), .ZN(P2_U3225) );
  XNOR2_X1 U9520 ( .A(n4557), .B(n7971), .ZN(n7972) );
  XNOR2_X1 U9521 ( .A(n7973), .B(n7972), .ZN(n7977) );
  AOI22_X1 U9522 ( .A1(n8053), .A2(n8392), .B1(n8390), .B2(n8054), .ZN(n8217)
         );
  OAI22_X1 U9523 ( .A1(n8217), .A2(n8022), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9479), .ZN(n7974) );
  AOI21_X1 U9524 ( .B1(n8221), .B2(n8033), .A(n7974), .ZN(n7976) );
  NAND2_X1 U9525 ( .A1(n8439), .A2(n8047), .ZN(n7975) );
  OAI211_X1 U9526 ( .C1(n7977), .C2(n8036), .A(n7976), .B(n7975), .ZN(P2_U3227) );
  NAND2_X1 U9527 ( .A1(n7978), .A2(n7979), .ZN(n7987) );
  OAI21_X1 U9528 ( .B1(n7979), .B2(n7978), .A(n7987), .ZN(n7980) );
  NAND2_X1 U9529 ( .A1(n7980), .A2(n8038), .ZN(n7985) );
  OAI22_X1 U9530 ( .A1(n7981), .A2(n8030), .B1(n8029), .B2(n8031), .ZN(n7982)
         );
  AOI211_X1 U9531 ( .C1(n8382), .C2(n8033), .A(n7983), .B(n7982), .ZN(n7984)
         );
  OAI211_X1 U9532 ( .C1(n8384), .C2(n8026), .A(n7985), .B(n7984), .ZN(P2_U3228) );
  NAND2_X1 U9533 ( .A1(n7987), .A2(n7986), .ZN(n7989) );
  XNOR2_X1 U9534 ( .A(n7989), .B(n7988), .ZN(n7996) );
  NAND2_X1 U9535 ( .A1(n8393), .A2(n8390), .ZN(n7991) );
  NAND2_X1 U9536 ( .A1(n8318), .A2(n8392), .ZN(n7990) );
  NAND2_X1 U9537 ( .A1(n7991), .A2(n7990), .ZN(n8349) );
  INV_X1 U9538 ( .A(n8349), .ZN(n7992) );
  OAI22_X1 U9539 ( .A1(n8022), .A2(n7992), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5358), .ZN(n7993) );
  AOI21_X1 U9540 ( .B1(n8355), .B2(n8033), .A(n7993), .ZN(n7995) );
  NAND2_X1 U9541 ( .A1(n8480), .A2(n8047), .ZN(n7994) );
  OAI211_X1 U9542 ( .C1(n7996), .C2(n8036), .A(n7995), .B(n7994), .ZN(P2_U3230) );
  INV_X1 U9543 ( .A(n7997), .ZN(n7998) );
  OAI21_X1 U9544 ( .B1(n8000), .B2(n7999), .A(n7998), .ZN(n8004) );
  XNOR2_X1 U9545 ( .A(n8002), .B(n8001), .ZN(n8003) );
  XNOR2_X1 U9546 ( .A(n8004), .B(n8003), .ZN(n8010) );
  OAI22_X1 U9547 ( .A1(n8045), .A2(n8233), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8005), .ZN(n8008) );
  OAI22_X1 U9548 ( .A1(n8006), .A2(n8030), .B1(n8029), .B2(n8042), .ZN(n8007)
         );
  AOI211_X1 U9549 ( .C1(n8442), .C2(n8047), .A(n8008), .B(n8007), .ZN(n8009)
         );
  OAI21_X1 U9550 ( .B1(n8010), .B2(n8036), .A(n8009), .ZN(P2_U3231) );
  XNOR2_X1 U9551 ( .A(n8012), .B(n8011), .ZN(n8016) );
  OAI22_X1 U9552 ( .A1(n8045), .A2(n8299), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9481), .ZN(n8014) );
  OAI22_X1 U9553 ( .A1(n8306), .A2(n8030), .B1(n8029), .B2(n8308), .ZN(n8013)
         );
  AOI211_X1 U9554 ( .C1(n8464), .C2(n8047), .A(n8014), .B(n8013), .ZN(n8015)
         );
  OAI21_X1 U9555 ( .B1(n8016), .B2(n8036), .A(n8015), .ZN(P2_U3235) );
  OAI21_X1 U9556 ( .B1(n8019), .B2(n8018), .A(n8017), .ZN(n8020) );
  NAND2_X1 U9557 ( .A1(n8020), .A2(n8038), .ZN(n8025) );
  AOI22_X1 U9558 ( .A1(n8229), .A2(n8392), .B1(n8056), .B2(n8390), .ZN(n8275)
         );
  OAI22_X1 U9559 ( .A1(n8022), .A2(n8275), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8021), .ZN(n8023) );
  AOI21_X1 U9560 ( .B1(n8270), .B2(n8033), .A(n8023), .ZN(n8024) );
  OAI211_X1 U9561 ( .C1(n8272), .C2(n8026), .A(n8025), .B(n8024), .ZN(P2_U3237) );
  XNOR2_X1 U9562 ( .A(n8028), .B(n8027), .ZN(n8037) );
  NOR2_X1 U9563 ( .A1(n9454), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8127) );
  OAI22_X1 U9564 ( .A1(n8031), .A2(n8030), .B1(n8029), .B2(n8306), .ZN(n8032)
         );
  AOI211_X1 U9565 ( .C1(n8033), .C2(n8336), .A(n8127), .B(n8032), .ZN(n8035)
         );
  NAND2_X1 U9566 ( .A1(n8474), .A2(n8047), .ZN(n8034) );
  OAI211_X1 U9567 ( .C1(n8037), .C2(n8036), .A(n8035), .B(n8034), .ZN(P2_U3240) );
  OAI211_X1 U9568 ( .C1(n8041), .C2(n8040), .A(n8039), .B(n8038), .ZN(n8049)
         );
  OAI22_X1 U9569 ( .A1(n8157), .A2(n8307), .B1(n8042), .B2(n8305), .ZN(n8199)
         );
  AOI22_X1 U9570 ( .A1(n8199), .A2(n8043), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3152), .ZN(n8044) );
  OAI21_X1 U9571 ( .B1(n8202), .B2(n8045), .A(n8044), .ZN(n8046) );
  AOI21_X1 U9572 ( .B1(n8433), .B2(n8047), .A(n8046), .ZN(n8048) );
  NAND2_X1 U9573 ( .A1(n8049), .A2(n8048), .ZN(P2_U3242) );
  MUX2_X1 U9574 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8050), .S(P2_U3966), .Z(
        P2_U3582) );
  MUX2_X1 U9575 ( .A(n8051), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8055), .Z(
        P2_U3580) );
  MUX2_X1 U9576 ( .A(n8052), .B(P2_DATAO_REG_27__SCAN_IN), .S(n8055), .Z(
        P2_U3579) );
  MUX2_X1 U9577 ( .A(n8053), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8055), .Z(
        P2_U3578) );
  MUX2_X1 U9578 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8230), .S(P2_U3966), .Z(
        P2_U3577) );
  MUX2_X1 U9579 ( .A(n8054), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8055), .Z(
        P2_U3576) );
  MUX2_X1 U9580 ( .A(n8229), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8055), .Z(
        P2_U3575) );
  MUX2_X1 U9581 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8283), .S(P2_U3966), .Z(
        P2_U3574) );
  INV_X2 U9582 ( .A(n8055), .ZN(P2_U3966) );
  MUX2_X1 U9583 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8056), .S(P2_U3966), .Z(
        P2_U3573) );
  MUX2_X1 U9584 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8319), .S(P2_U3966), .Z(
        P2_U3572) );
  MUX2_X1 U9585 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8341), .S(P2_U3966), .Z(
        P2_U3571) );
  MUX2_X1 U9586 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8318), .S(P2_U3966), .Z(
        P2_U3570) );
  MUX2_X1 U9587 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8372), .S(P2_U3966), .Z(
        P2_U3569) );
  MUX2_X1 U9588 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8393), .S(P2_U3966), .Z(
        P2_U3568) );
  MUX2_X1 U9589 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8373), .S(P2_U3966), .Z(
        P2_U3567) );
  MUX2_X1 U9590 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8391), .S(P2_U3966), .Z(
        P2_U3566) );
  MUX2_X1 U9591 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n8057), .S(P2_U3966), .Z(
        P2_U3565) );
  MUX2_X1 U9592 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n8058), .S(P2_U3966), .Z(
        P2_U3564) );
  MUX2_X1 U9593 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n8059), .S(P2_U3966), .Z(
        P2_U3563) );
  MUX2_X1 U9594 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n8060), .S(P2_U3966), .Z(
        P2_U3562) );
  MUX2_X1 U9595 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n8061), .S(P2_U3966), .Z(
        P2_U3561) );
  MUX2_X1 U9596 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n8062), .S(P2_U3966), .Z(
        P2_U3560) );
  MUX2_X1 U9597 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n8063), .S(P2_U3966), .Z(
        P2_U3559) );
  MUX2_X1 U9598 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n8064), .S(P2_U3966), .Z(
        P2_U3558) );
  MUX2_X1 U9599 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n8065), .S(P2_U3966), .Z(
        P2_U3557) );
  MUX2_X1 U9600 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n8067), .S(P2_U3966), .Z(
        P2_U3556) );
  MUX2_X1 U9601 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n8068), .S(P2_U3966), .Z(
        P2_U3555) );
  MUX2_X1 U9602 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n5818), .S(P2_U3966), .Z(
        P2_U3554) );
  MUX2_X1 U9603 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n5808), .S(P2_U3966), .Z(
        P2_U3553) );
  OAI211_X1 U9604 ( .C1(n8071), .C2(n8070), .A(n9929), .B(n8069), .ZN(n8080)
         );
  NOR2_X1 U9605 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9557), .ZN(n8072) );
  AOI21_X1 U9606 ( .B1(n9935), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n8072), .ZN(
        n8079) );
  NAND2_X1 U9607 ( .A1(n9619), .A2(n8073), .ZN(n8078) );
  OAI211_X1 U9608 ( .C1(n8076), .C2(n8075), .A(n9930), .B(n8074), .ZN(n8077)
         );
  NAND4_X1 U9609 ( .A1(n8080), .A2(n8079), .A3(n8078), .A4(n8077), .ZN(
        P2_U3253) );
  OAI211_X1 U9610 ( .C1(n8083), .C2(n8082), .A(n9929), .B(n8081), .ZN(n8092)
         );
  AOI21_X1 U9611 ( .B1(n9935), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n8084), .ZN(
        n8091) );
  NAND2_X1 U9612 ( .A1(n9619), .A2(n8085), .ZN(n8090) );
  OAI211_X1 U9613 ( .C1(n8088), .C2(n8087), .A(n8086), .B(n9930), .ZN(n8089)
         );
  NAND4_X1 U9614 ( .A1(n8092), .A2(n8091), .A3(n8090), .A4(n8089), .ZN(
        P2_U3254) );
  OAI211_X1 U9615 ( .C1(n8095), .C2(n8094), .A(n8093), .B(n9930), .ZN(n8104)
         );
  NOR2_X1 U9616 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9540), .ZN(n8096) );
  AOI21_X1 U9617 ( .B1(n9935), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n8096), .ZN(
        n8103) );
  OAI211_X1 U9618 ( .C1(n8099), .C2(n8098), .A(n9929), .B(n8097), .ZN(n8102)
         );
  NAND2_X1 U9619 ( .A1(n9619), .A2(n8100), .ZN(n8101) );
  NAND4_X1 U9620 ( .A1(n8104), .A2(n8103), .A3(n8102), .A4(n8101), .ZN(
        P2_U3255) );
  INV_X1 U9621 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8108) );
  NAND2_X1 U9622 ( .A1(n8125), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8121) );
  INV_X1 U9623 ( .A(n8121), .ZN(n8107) );
  AOI21_X1 U9624 ( .B1(n8108), .B2(n8119), .A(n8107), .ZN(n8109) );
  OAI211_X1 U9625 ( .C1(n8110), .C2(n8109), .A(n9929), .B(n8120), .ZN(n8118)
         );
  NOR2_X1 U9626 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5358), .ZN(n8116) );
  OAI21_X1 U9627 ( .B1(n8112), .B2(P2_REG1_REG_16__SCAN_IN), .A(n8111), .ZN(
        n8114) );
  XNOR2_X1 U9628 ( .A(n8125), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n8113) );
  NOR2_X1 U9629 ( .A1(n8113), .A2(n8114), .ZN(n8124) );
  AOI211_X1 U9630 ( .C1(n8114), .C2(n8113), .A(n8124), .B(n9613), .ZN(n8115)
         );
  AOI211_X1 U9631 ( .C1(P2_ADDR_REG_17__SCAN_IN), .C2(n9935), .A(n8116), .B(
        n8115), .ZN(n8117) );
  OAI211_X1 U9632 ( .C1(n9932), .C2(n8119), .A(n8118), .B(n8117), .ZN(P2_U3262) );
  NAND2_X1 U9633 ( .A1(n8121), .A2(n8120), .ZN(n8122) );
  NOR2_X1 U9634 ( .A1(n8122), .A2(n8135), .ZN(n8133) );
  AOI21_X1 U9635 ( .B1(n8123), .B2(P2_REG2_REG_18__SCAN_IN), .A(n8134), .ZN(
        n8132) );
  AOI21_X1 U9636 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(n8125), .A(n8124), .ZN(
        n8137) );
  INV_X1 U9637 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8126) );
  XNOR2_X1 U9638 ( .A(n8135), .B(n8126), .ZN(n8138) );
  XOR2_X1 U9639 ( .A(n8137), .B(n8138), .Z(n8129) );
  AOI21_X1 U9640 ( .B1(n9935), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n8127), .ZN(
        n8128) );
  OAI21_X1 U9641 ( .B1(n9613), .B2(n8129), .A(n8128), .ZN(n8130) );
  AOI21_X1 U9642 ( .B1(n8135), .B2(n9619), .A(n8130), .ZN(n8131) );
  OAI21_X1 U9643 ( .B1(n8132), .B2(n9933), .A(n8131), .ZN(P2_U3263) );
  INV_X1 U9644 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n8146) );
  XOR2_X1 U9645 ( .A(n4372), .B(P2_REG2_REG_19__SCAN_IN), .Z(n8141) );
  NOR2_X1 U9646 ( .A1(n8135), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8136) );
  AOI21_X1 U9647 ( .B1(n8138), .B2(n8137), .A(n8136), .ZN(n8139) );
  XNOR2_X1 U9648 ( .A(n8139), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8142) );
  INV_X1 U9649 ( .A(n8142), .ZN(n8140) );
  AOI22_X1 U9650 ( .A1(n8141), .A2(n9929), .B1(n8140), .B2(n9930), .ZN(n8143)
         );
  INV_X1 U9651 ( .A(n8144), .ZN(n8145) );
  INV_X1 U9652 ( .A(n8147), .ZN(n8148) );
  NAND2_X1 U9653 ( .A1(n8149), .A2(n8148), .ZN(n8412) );
  NAND3_X1 U9654 ( .A1(n8412), .A2(n8402), .A3(n8411), .ZN(n8152) );
  AOI21_X1 U9655 ( .B1(n8368), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8150), .ZN(
        n8151) );
  OAI211_X1 U9656 ( .C1(n8415), .C2(n8406), .A(n8152), .B(n8151), .ZN(P2_U3266) );
  XNOR2_X1 U9657 ( .A(n8153), .B(n8155), .ZN(n8420) );
  INV_X1 U9658 ( .A(n8420), .ZN(n8170) );
  OAI211_X1 U9659 ( .C1(n8156), .C2(n8155), .A(n8154), .B(n8395), .ZN(n8161)
         );
  OAI22_X1 U9660 ( .A1(n8158), .A2(n8307), .B1(n8157), .B2(n8305), .ZN(n8159)
         );
  INV_X1 U9661 ( .A(n8159), .ZN(n8160) );
  NAND2_X1 U9662 ( .A1(n8161), .A2(n8160), .ZN(n8421) );
  NAND2_X1 U9663 ( .A1(n8422), .A2(n8173), .ZN(n8162) );
  NAND2_X1 U9664 ( .A1(n8163), .A2(n8162), .ZN(n8423) );
  AOI22_X1 U9665 ( .A1(n8164), .A2(n9944), .B1(P2_REG2_REG_28__SCAN_IN), .B2(
        n8368), .ZN(n8166) );
  NAND2_X1 U9666 ( .A1(n8422), .A2(n8359), .ZN(n8165) );
  OAI211_X1 U9667 ( .C1(n8423), .C2(n8167), .A(n8166), .B(n8165), .ZN(n8168)
         );
  AOI21_X1 U9668 ( .B1(n8421), .B2(n9953), .A(n8168), .ZN(n8169) );
  OAI21_X1 U9669 ( .B1(n8170), .B2(n8365), .A(n8169), .ZN(P2_U3268) );
  XNOR2_X1 U9670 ( .A(n8171), .B(n8172), .ZN(n8431) );
  INV_X1 U9671 ( .A(n8173), .ZN(n8174) );
  AOI21_X1 U9672 ( .B1(n8427), .B2(n8206), .A(n8174), .ZN(n8428) );
  INV_X1 U9673 ( .A(n8427), .ZN(n8178) );
  INV_X1 U9674 ( .A(n8175), .ZN(n8176) );
  AOI22_X1 U9675 ( .A1(n8176), .A2(n9944), .B1(P2_REG2_REG_27__SCAN_IN), .B2(
        n8368), .ZN(n8177) );
  OAI21_X1 U9676 ( .B1(n8178), .B2(n8406), .A(n8177), .ZN(n8187) );
  AOI21_X1 U9677 ( .B1(n8180), .B2(n8179), .A(n8347), .ZN(n8185) );
  OAI22_X1 U9678 ( .A1(n8182), .A2(n8307), .B1(n8181), .B2(n8305), .ZN(n8183)
         );
  AOI21_X1 U9679 ( .B1(n8185), .B2(n8184), .A(n8183), .ZN(n8430) );
  NOR2_X1 U9680 ( .A1(n8430), .A2(n8368), .ZN(n8186) );
  AOI211_X1 U9681 ( .C1(n8428), .C2(n8402), .A(n8187), .B(n8186), .ZN(n8188)
         );
  OAI21_X1 U9682 ( .B1(n8431), .B2(n8365), .A(n8188), .ZN(P2_U3269) );
  NAND2_X1 U9683 ( .A1(n8212), .A2(n8213), .ZN(n8190) );
  NAND2_X1 U9684 ( .A1(n8190), .A2(n8189), .ZN(n8192) );
  XNOR2_X1 U9685 ( .A(n8192), .B(n8191), .ZN(n8436) );
  INV_X1 U9686 ( .A(n8193), .ZN(n8196) );
  OAI21_X1 U9687 ( .B1(n8196), .B2(n8195), .A(n8194), .ZN(n8198) );
  AOI21_X1 U9688 ( .B1(n8198), .B2(n8197), .A(n8347), .ZN(n8200) );
  NOR2_X1 U9689 ( .A1(n8200), .A2(n8199), .ZN(n8435) );
  INV_X1 U9690 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8201) );
  OAI22_X1 U9691 ( .A1(n8202), .A2(n8356), .B1(n8201), .B2(n9953), .ZN(n8203)
         );
  AOI21_X1 U9692 ( .B1(n8433), .B2(n8359), .A(n8203), .ZN(n8208) );
  OR2_X1 U9693 ( .A1(n8204), .A2(n8219), .ZN(n8205) );
  AND3_X1 U9694 ( .A1(n8206), .A2(n8205), .A3(n8499), .ZN(n8432) );
  AND2_X1 U9695 ( .A1(n9953), .A2(n8325), .ZN(n8362) );
  NAND2_X1 U9696 ( .A1(n8432), .A2(n8362), .ZN(n8207) );
  OAI211_X1 U9697 ( .C1(n8435), .C2(n8368), .A(n8208), .B(n8207), .ZN(n8209)
         );
  INV_X1 U9698 ( .A(n8209), .ZN(n8210) );
  OAI21_X1 U9699 ( .B1(n8436), .B2(n8365), .A(n8210), .ZN(P2_U3270) );
  XNOR2_X1 U9700 ( .A(n8212), .B(n8211), .ZN(n8441) );
  NAND3_X1 U9701 ( .A1(n8215), .A2(n8214), .A3(n8213), .ZN(n8216) );
  NAND3_X1 U9702 ( .A1(n8193), .A2(n8395), .A3(n8216), .ZN(n8218) );
  NAND2_X1 U9703 ( .A1(n8218), .A2(n8217), .ZN(n8437) );
  OAI21_X1 U9704 ( .B1(n8232), .B2(n8224), .A(n8499), .ZN(n8220) );
  NOR2_X1 U9705 ( .A1(n8220), .A2(n8219), .ZN(n8438) );
  NAND2_X1 U9706 ( .A1(n8438), .A2(n8362), .ZN(n8223) );
  AOI22_X1 U9707 ( .A1(n8368), .A2(P2_REG2_REG_25__SCAN_IN), .B1(n8221), .B2(
        n9944), .ZN(n8222) );
  OAI211_X1 U9708 ( .C1(n8224), .C2(n8406), .A(n8223), .B(n8222), .ZN(n8225)
         );
  AOI21_X1 U9709 ( .B1(n8437), .B2(n9953), .A(n8225), .ZN(n8226) );
  OAI21_X1 U9710 ( .B1(n8441), .B2(n8365), .A(n8226), .ZN(P2_U3271) );
  XNOR2_X1 U9711 ( .A(n8227), .B(n8228), .ZN(n8231) );
  AOI222_X1 U9712 ( .A1(n8395), .A2(n8231), .B1(n8230), .B2(n8392), .C1(n8229), 
        .C2(n8390), .ZN(n8445) );
  AOI21_X1 U9713 ( .B1(n8442), .B2(n8253), .A(n8232), .ZN(n8443) );
  INV_X1 U9714 ( .A(n8442), .ZN(n8236) );
  INV_X1 U9715 ( .A(n8233), .ZN(n8234) );
  AOI22_X1 U9716 ( .A1(n8368), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n8234), .B2(
        n9944), .ZN(n8235) );
  OAI21_X1 U9717 ( .B1(n8236), .B2(n8406), .A(n8235), .ZN(n8242) );
  INV_X1 U9718 ( .A(n8237), .ZN(n8238) );
  AOI21_X1 U9719 ( .B1(n8240), .B2(n8239), .A(n8238), .ZN(n8446) );
  NOR2_X1 U9720 ( .A1(n8446), .A2(n8365), .ZN(n8241) );
  AOI211_X1 U9721 ( .C1(n8443), .C2(n8402), .A(n8242), .B(n8241), .ZN(n8243)
         );
  OAI21_X1 U9722 ( .B1(n8368), .B2(n8445), .A(n8243), .ZN(P2_U3272) );
  OAI21_X1 U9723 ( .B1(n8245), .B2(n8261), .A(n8244), .ZN(n8246) );
  NAND2_X1 U9724 ( .A1(n8246), .A2(n8395), .ZN(n8251) );
  OAI22_X1 U9725 ( .A1(n8248), .A2(n8307), .B1(n8247), .B2(n8305), .ZN(n8249)
         );
  INV_X1 U9726 ( .A(n8249), .ZN(n8250) );
  NAND2_X1 U9727 ( .A1(n8251), .A2(n8250), .ZN(n8453) );
  INV_X1 U9728 ( .A(n8453), .ZN(n8264) );
  NAND2_X1 U9729 ( .A1(n8267), .A2(n8448), .ZN(n8252) );
  AND2_X1 U9730 ( .A1(n8253), .A2(n8252), .ZN(n8449) );
  INV_X1 U9731 ( .A(n8254), .ZN(n8255) );
  AOI22_X1 U9732 ( .A1(n8368), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n8255), .B2(
        n9944), .ZN(n8256) );
  OAI21_X1 U9733 ( .B1(n8257), .B2(n8406), .A(n8256), .ZN(n8258) );
  AOI21_X1 U9734 ( .B1(n8449), .B2(n8402), .A(n8258), .ZN(n8263) );
  NAND2_X1 U9735 ( .A1(n8260), .A2(n8261), .ZN(n8447) );
  NAND3_X1 U9736 ( .A1(n8259), .A2(n8447), .A3(n8409), .ZN(n8262) );
  OAI211_X1 U9737 ( .C1(n8264), .C2(n8368), .A(n8263), .B(n8262), .ZN(P2_U3273) );
  XNOR2_X1 U9738 ( .A(n8266), .B(n8265), .ZN(n8458) );
  INV_X1 U9739 ( .A(n8287), .ZN(n8269) );
  INV_X1 U9740 ( .A(n8267), .ZN(n8268) );
  AOI21_X1 U9741 ( .B1(n8454), .B2(n8269), .A(n8268), .ZN(n8455) );
  AOI22_X1 U9742 ( .A1(n8368), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8270), .B2(
        n9944), .ZN(n8271) );
  OAI21_X1 U9743 ( .B1(n8272), .B2(n8406), .A(n8271), .ZN(n8280) );
  AOI21_X1 U9744 ( .B1(n8274), .B2(n8273), .A(n8347), .ZN(n8278) );
  INV_X1 U9745 ( .A(n8275), .ZN(n8276) );
  AOI21_X1 U9746 ( .B1(n8278), .B2(n8277), .A(n8276), .ZN(n8457) );
  NOR2_X1 U9747 ( .A1(n8457), .A2(n8368), .ZN(n8279) );
  AOI211_X1 U9748 ( .C1(n8455), .C2(n8402), .A(n8280), .B(n8279), .ZN(n8281)
         );
  OAI21_X1 U9749 ( .B1(n8458), .B2(n8365), .A(n8281), .ZN(P2_U3274) );
  XNOR2_X1 U9750 ( .A(n8282), .B(n8292), .ZN(n8284) );
  AOI222_X1 U9751 ( .A1(n8395), .A2(n8284), .B1(n8283), .B2(n8392), .C1(n8319), 
        .C2(n8390), .ZN(n8462) );
  NOR2_X1 U9752 ( .A1(n8285), .A2(n8291), .ZN(n8286) );
  NOR2_X1 U9753 ( .A1(n8287), .A2(n8286), .ZN(n8460) );
  INV_X1 U9754 ( .A(n8288), .ZN(n8289) );
  AOI22_X1 U9755 ( .A1(n8368), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8289), .B2(
        n9944), .ZN(n8290) );
  OAI21_X1 U9756 ( .B1(n8291), .B2(n8406), .A(n8290), .ZN(n8295) );
  XNOR2_X1 U9757 ( .A(n8293), .B(n8292), .ZN(n8463) );
  NOR2_X1 U9758 ( .A1(n8463), .A2(n8365), .ZN(n8294) );
  AOI211_X1 U9759 ( .C1(n8460), .C2(n8402), .A(n8295), .B(n8294), .ZN(n8296)
         );
  OAI21_X1 U9760 ( .B1(n8368), .B2(n8462), .A(n8296), .ZN(P2_U3275) );
  XNOR2_X1 U9761 ( .A(n8297), .B(n8304), .ZN(n8468) );
  INV_X1 U9762 ( .A(n8315), .ZN(n8298) );
  AOI21_X1 U9763 ( .B1(n8464), .B2(n8298), .A(n8285), .ZN(n8465) );
  INV_X1 U9764 ( .A(n8299), .ZN(n8300) );
  AOI22_X1 U9765 ( .A1(n8368), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8300), .B2(
        n9944), .ZN(n8301) );
  OAI21_X1 U9766 ( .B1(n8302), .B2(n8406), .A(n8301), .ZN(n8313) );
  AOI21_X1 U9767 ( .B1(n8303), .B2(n8304), .A(n8347), .ZN(n8311) );
  OAI22_X1 U9768 ( .A1(n8308), .A2(n8307), .B1(n8306), .B2(n8305), .ZN(n8309)
         );
  AOI21_X1 U9769 ( .B1(n8311), .B2(n8310), .A(n8309), .ZN(n8467) );
  NOR2_X1 U9770 ( .A1(n8467), .A2(n8368), .ZN(n8312) );
  AOI211_X1 U9771 ( .C1(n8465), .C2(n8402), .A(n8313), .B(n8312), .ZN(n8314)
         );
  OAI21_X1 U9772 ( .B1(n8365), .B2(n8468), .A(n8314), .ZN(P2_U3276) );
  AOI211_X1 U9773 ( .C1(n8471), .C2(n8334), .A(n10010), .B(n8315), .ZN(n8470)
         );
  XNOR2_X1 U9774 ( .A(n8316), .B(n8323), .ZN(n8317) );
  NAND2_X1 U9775 ( .A1(n8317), .A2(n8395), .ZN(n8321) );
  AOI22_X1 U9776 ( .A1(n8319), .A2(n8392), .B1(n8390), .B2(n8318), .ZN(n8320)
         );
  NAND2_X1 U9777 ( .A1(n8321), .A2(n8320), .ZN(n8469) );
  XNOR2_X1 U9778 ( .A(n8322), .B(n8323), .ZN(n8473) );
  NOR2_X1 U9779 ( .A1(n8473), .A2(n8379), .ZN(n8324) );
  AOI211_X1 U9780 ( .C1(n8470), .C2(n8325), .A(n8469), .B(n8324), .ZN(n8331)
         );
  INV_X1 U9781 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8327) );
  OAI22_X1 U9782 ( .A1(n9953), .A2(n8327), .B1(n8326), .B2(n8356), .ZN(n8329)
         );
  NOR2_X1 U9783 ( .A1(n8473), .A2(n8388), .ZN(n8328) );
  AOI211_X1 U9784 ( .C1(n8359), .C2(n8471), .A(n8329), .B(n8328), .ZN(n8330)
         );
  OAI21_X1 U9785 ( .B1(n8331), .B2(n8368), .A(n8330), .ZN(P2_U3277) );
  XOR2_X1 U9786 ( .A(n8333), .B(n8332), .Z(n8478) );
  INV_X1 U9787 ( .A(n8334), .ZN(n8335) );
  AOI21_X1 U9788 ( .B1(n8474), .B2(n8360), .A(n8335), .ZN(n8475) );
  AOI22_X1 U9789 ( .A1(n8368), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8336), .B2(
        n9944), .ZN(n8337) );
  OAI21_X1 U9790 ( .B1(n4462), .B2(n8406), .A(n8337), .ZN(n8344) );
  OAI21_X1 U9791 ( .B1(n8340), .B2(n8339), .A(n8338), .ZN(n8342) );
  AOI222_X1 U9792 ( .A1(n8395), .A2(n8342), .B1(n8341), .B2(n8392), .C1(n8372), 
        .C2(n8390), .ZN(n8477) );
  NOR2_X1 U9793 ( .A1(n8477), .A2(n8368), .ZN(n8343) );
  AOI211_X1 U9794 ( .C1(n8475), .C2(n8402), .A(n8344), .B(n8343), .ZN(n8345)
         );
  OAI21_X1 U9795 ( .B1(n8478), .B2(n8365), .A(n8345), .ZN(P2_U3278) );
  AOI21_X1 U9796 ( .B1(n8346), .B2(n8352), .A(n8347), .ZN(n8350) );
  AOI21_X1 U9797 ( .B1(n8350), .B2(n8348), .A(n8349), .ZN(n8482) );
  OAI21_X1 U9798 ( .B1(n8353), .B2(n8352), .A(n8351), .ZN(n8354) );
  INV_X1 U9799 ( .A(n8354), .ZN(n8483) );
  INV_X1 U9800 ( .A(n8355), .ZN(n8357) );
  OAI22_X1 U9801 ( .A1(n9953), .A2(n8108), .B1(n8357), .B2(n8356), .ZN(n8358)
         );
  AOI21_X1 U9802 ( .B1(n8480), .B2(n8359), .A(n8358), .ZN(n8364) );
  AOI21_X1 U9803 ( .B1(n8381), .B2(n8480), .A(n10010), .ZN(n8361) );
  AND2_X1 U9804 ( .A1(n8361), .A2(n8360), .ZN(n8479) );
  NAND2_X1 U9805 ( .A1(n8479), .A2(n8362), .ZN(n8363) );
  OAI211_X1 U9806 ( .C1(n8483), .C2(n8365), .A(n8364), .B(n8363), .ZN(n8366)
         );
  INV_X1 U9807 ( .A(n8366), .ZN(n8367) );
  OAI21_X1 U9808 ( .B1(n8368), .B2(n8482), .A(n8367), .ZN(P2_U3279) );
  NAND2_X1 U9809 ( .A1(n8369), .A2(n8375), .ZN(n8370) );
  NAND2_X1 U9810 ( .A1(n8371), .A2(n8370), .ZN(n8488) );
  AOI22_X1 U9811 ( .A1(n8390), .A2(n8373), .B1(n8372), .B2(n8392), .ZN(n8378)
         );
  XNOR2_X1 U9812 ( .A(n8374), .B(n8375), .ZN(n8376) );
  NAND2_X1 U9813 ( .A1(n8376), .A2(n8395), .ZN(n8377) );
  OAI211_X1 U9814 ( .C1(n8488), .C2(n8379), .A(n8378), .B(n8377), .ZN(n8490)
         );
  NAND2_X1 U9815 ( .A1(n8490), .A2(n9953), .ZN(n8387) );
  OR2_X1 U9816 ( .A1(n8400), .A2(n8384), .ZN(n8380) );
  AND2_X1 U9817 ( .A1(n8381), .A2(n8380), .ZN(n8485) );
  AOI22_X1 U9818 ( .A1(n8368), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n8382), .B2(
        n9944), .ZN(n8383) );
  OAI21_X1 U9819 ( .B1(n8384), .B2(n8406), .A(n8383), .ZN(n8385) );
  AOI21_X1 U9820 ( .B1(n8485), .B2(n8402), .A(n8385), .ZN(n8386) );
  OAI211_X1 U9821 ( .C1(n8488), .C2(n8388), .A(n8387), .B(n8386), .ZN(P2_U3280) );
  XNOR2_X1 U9822 ( .A(n8389), .B(n8397), .ZN(n8394) );
  AOI222_X1 U9823 ( .A1(n8395), .A2(n8394), .B1(n8393), .B2(n8392), .C1(n8391), 
        .C2(n8390), .ZN(n8495) );
  OAI21_X1 U9824 ( .B1(n8398), .B2(n8397), .A(n8396), .ZN(n8491) );
  INV_X1 U9825 ( .A(n8399), .ZN(n8401) );
  AOI21_X1 U9826 ( .B1(n8492), .B2(n8401), .A(n8400), .ZN(n8493) );
  NAND2_X1 U9827 ( .A1(n8493), .A2(n8402), .ZN(n8405) );
  AOI22_X1 U9828 ( .A1(n8368), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n8403), .B2(
        n9944), .ZN(n8404) );
  OAI211_X1 U9829 ( .C1(n8407), .C2(n8406), .A(n8405), .B(n8404), .ZN(n8408)
         );
  AOI21_X1 U9830 ( .B1(n8491), .B2(n8409), .A(n8408), .ZN(n8410) );
  OAI21_X1 U9831 ( .B1(n8495), .B2(n8368), .A(n8410), .ZN(P2_U3281) );
  NAND3_X1 U9832 ( .A1(n8412), .A2(n8499), .A3(n8411), .ZN(n8414) );
  OAI211_X1 U9833 ( .C1(n8415), .C2(n10008), .A(n8414), .B(n8413), .ZN(n8512)
         );
  MUX2_X1 U9834 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n8512), .S(n10033), .Z(
        P2_U3550) );
  MUX2_X1 U9835 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n8513), .S(n10033), .Z(
        P2_U3549) );
  INV_X1 U9836 ( .A(n8503), .ZN(n10015) );
  INV_X1 U9837 ( .A(n8421), .ZN(n8426) );
  OAI22_X1 U9838 ( .A1(n8423), .A2(n10010), .B1(n4469), .B2(n10008), .ZN(n8424) );
  INV_X1 U9839 ( .A(n8424), .ZN(n8425) );
  NAND3_X1 U9840 ( .A1(n4807), .A2(n8426), .A3(n8425), .ZN(n8514) );
  MUX2_X1 U9841 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n8514), .S(n10033), .Z(
        P2_U3548) );
  AOI22_X1 U9842 ( .A1(n8428), .A2(n8499), .B1(n8498), .B2(n8427), .ZN(n8429)
         );
  OAI211_X1 U9843 ( .C1(n8431), .C2(n8503), .A(n8430), .B(n8429), .ZN(n8515)
         );
  MUX2_X1 U9844 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n8515), .S(n10033), .Z(
        P2_U3547) );
  AOI21_X1 U9845 ( .B1(n8498), .B2(n8433), .A(n8432), .ZN(n8434) );
  OAI211_X1 U9846 ( .C1(n8503), .C2(n8436), .A(n8435), .B(n8434), .ZN(n8516)
         );
  MUX2_X1 U9847 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n8516), .S(n10033), .Z(
        P2_U3546) );
  AOI211_X1 U9848 ( .C1(n8498), .C2(n8439), .A(n8438), .B(n8437), .ZN(n8440)
         );
  OAI21_X1 U9849 ( .B1(n8503), .B2(n8441), .A(n8440), .ZN(n8517) );
  MUX2_X1 U9850 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n8517), .S(n10033), .Z(
        P2_U3545) );
  AOI22_X1 U9851 ( .A1(n8443), .A2(n8499), .B1(n8498), .B2(n8442), .ZN(n8444)
         );
  OAI211_X1 U9852 ( .C1(n8503), .C2(n8446), .A(n8445), .B(n8444), .ZN(n8518)
         );
  MUX2_X1 U9853 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8518), .S(n10033), .Z(
        P2_U3544) );
  NAND3_X1 U9854 ( .A1(n8259), .A2(n8447), .A3(n10015), .ZN(n8451) );
  AOI22_X1 U9855 ( .A1(n8449), .A2(n8499), .B1(n8498), .B2(n8448), .ZN(n8450)
         );
  NAND2_X1 U9856 ( .A1(n8451), .A2(n8450), .ZN(n8452) );
  MUX2_X1 U9857 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n8519), .S(n10033), .Z(
        P2_U3543) );
  AOI22_X1 U9858 ( .A1(n8455), .A2(n8499), .B1(n8498), .B2(n8454), .ZN(n8456)
         );
  OAI211_X1 U9859 ( .C1(n8458), .C2(n8503), .A(n8457), .B(n8456), .ZN(n8520)
         );
  MUX2_X1 U9860 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n8520), .S(n10033), .Z(
        P2_U3542) );
  AOI22_X1 U9861 ( .A1(n8460), .A2(n8499), .B1(n8498), .B2(n8459), .ZN(n8461)
         );
  OAI211_X1 U9862 ( .C1(n8503), .C2(n8463), .A(n8462), .B(n8461), .ZN(n8521)
         );
  MUX2_X1 U9863 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n8521), .S(n10033), .Z(
        P2_U3541) );
  AOI22_X1 U9864 ( .A1(n8465), .A2(n8499), .B1(n8498), .B2(n8464), .ZN(n8466)
         );
  OAI211_X1 U9865 ( .C1(n8468), .C2(n8503), .A(n8467), .B(n8466), .ZN(n8522)
         );
  MUX2_X1 U9866 ( .A(n8522), .B(P2_REG1_REG_20__SCAN_IN), .S(n10030), .Z(
        P2_U3540) );
  AOI211_X1 U9867 ( .C1(n8498), .C2(n8471), .A(n8470), .B(n8469), .ZN(n8472)
         );
  OAI21_X1 U9868 ( .B1(n8503), .B2(n8473), .A(n8472), .ZN(n8523) );
  MUX2_X1 U9869 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8523), .S(n10033), .Z(
        P2_U3539) );
  AOI22_X1 U9870 ( .A1(n8475), .A2(n8499), .B1(n8498), .B2(n8474), .ZN(n8476)
         );
  OAI211_X1 U9871 ( .C1(n8503), .C2(n8478), .A(n8477), .B(n8476), .ZN(n8524)
         );
  MUX2_X1 U9872 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n8524), .S(n10033), .Z(
        P2_U3538) );
  AOI21_X1 U9873 ( .B1(n8498), .B2(n8480), .A(n8479), .ZN(n8481) );
  OAI211_X1 U9874 ( .C1(n8483), .C2(n8503), .A(n8482), .B(n8481), .ZN(n8525)
         );
  MUX2_X1 U9875 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n8525), .S(n10033), .Z(
        P2_U3537) );
  AOI22_X1 U9876 ( .A1(n8485), .A2(n8499), .B1(n8498), .B2(n8484), .ZN(n8486)
         );
  OAI21_X1 U9877 ( .B1(n8488), .B2(n8487), .A(n8486), .ZN(n8489) );
  OR2_X1 U9878 ( .A1(n8490), .A2(n8489), .ZN(n8526) );
  MUX2_X1 U9879 ( .A(n8526), .B(P2_REG1_REG_16__SCAN_IN), .S(n10030), .Z(
        P2_U3536) );
  INV_X1 U9880 ( .A(n8491), .ZN(n8496) );
  AOI22_X1 U9881 ( .A1(n8493), .A2(n8499), .B1(n8498), .B2(n8492), .ZN(n8494)
         );
  OAI211_X1 U9882 ( .C1(n8503), .C2(n8496), .A(n8495), .B(n8494), .ZN(n8527)
         );
  MUX2_X1 U9883 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n8527), .S(n10033), .Z(
        P2_U3535) );
  AOI22_X1 U9884 ( .A1(n8500), .A2(n8499), .B1(n8498), .B2(n8497), .ZN(n8501)
         );
  OAI211_X1 U9885 ( .C1(n8504), .C2(n8503), .A(n8502), .B(n8501), .ZN(n8528)
         );
  MUX2_X1 U9886 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n8528), .S(n10033), .Z(
        P2_U3534) );
  INV_X1 U9887 ( .A(n8505), .ZN(n8506) );
  OAI22_X1 U9888 ( .A1(n8507), .A2(n10010), .B1(n8506), .B2(n10008), .ZN(n8508) );
  AOI21_X1 U9889 ( .B1(n8509), .B2(n10006), .A(n8508), .ZN(n8510) );
  NAND2_X1 U9890 ( .A1(n8511), .A2(n8510), .ZN(n8529) );
  MUX2_X1 U9891 ( .A(n8529), .B(P2_REG1_REG_13__SCAN_IN), .S(n10030), .Z(
        P2_U3533) );
  MUX2_X1 U9892 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n8512), .S(n10019), .Z(
        P2_U3518) );
  MUX2_X1 U9893 ( .A(n8514), .B(P2_REG0_REG_28__SCAN_IN), .S(n10017), .Z(
        P2_U3516) );
  MUX2_X1 U9894 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n8515), .S(n10019), .Z(
        P2_U3515) );
  MUX2_X1 U9895 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n8516), .S(n10019), .Z(
        P2_U3514) );
  MUX2_X1 U9896 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n8517), .S(n10019), .Z(
        P2_U3513) );
  MUX2_X1 U9897 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n8518), .S(n10019), .Z(
        P2_U3512) );
  MUX2_X1 U9898 ( .A(n8519), .B(P2_REG0_REG_23__SCAN_IN), .S(n10017), .Z(
        P2_U3511) );
  MUX2_X1 U9899 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n8520), .S(n10019), .Z(
        P2_U3510) );
  MUX2_X1 U9900 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n8521), .S(n10019), .Z(
        P2_U3509) );
  MUX2_X1 U9901 ( .A(n8522), .B(P2_REG0_REG_20__SCAN_IN), .S(n10017), .Z(
        P2_U3508) );
  MUX2_X1 U9902 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n8523), .S(n10019), .Z(
        P2_U3507) );
  MUX2_X1 U9903 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n8524), .S(n10019), .Z(
        P2_U3505) );
  MUX2_X1 U9904 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n8525), .S(n10019), .Z(
        P2_U3502) );
  MUX2_X1 U9905 ( .A(n8526), .B(P2_REG0_REG_16__SCAN_IN), .S(n10017), .Z(
        P2_U3499) );
  MUX2_X1 U9906 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n8527), .S(n10019), .Z(
        P2_U3496) );
  MUX2_X1 U9907 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n8528), .S(n10019), .Z(
        P2_U3493) );
  MUX2_X1 U9908 ( .A(n8529), .B(P2_REG0_REG_13__SCAN_IN), .S(n10017), .Z(
        P2_U3490) );
  NAND2_X1 U9909 ( .A1(n9363), .A2(n8530), .ZN(n8533) );
  NAND4_X1 U9910 ( .A1(n4988), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .A4(n8531), .ZN(n8532) );
  OAI211_X1 U9911 ( .C1(n8535), .C2(n8534), .A(n8533), .B(n8532), .ZN(P2_U3327) );
  MUX2_X1 U9912 ( .A(n8536), .B(P2_IR_REG_0__SCAN_IN), .S(P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  XNOR2_X1 U9913 ( .A(n8538), .B(n8537), .ZN(n8539) );
  XNOR2_X1 U9914 ( .A(n8540), .B(n8539), .ZN(n8545) );
  NOR2_X1 U9915 ( .A1(n8668), .A2(n9069), .ZN(n8543) );
  INV_X1 U9916 ( .A(n9103), .ZN(n8869) );
  AOI22_X1 U9917 ( .A1(n8666), .A2(n9075), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3084), .ZN(n8541) );
  OAI21_X1 U9918 ( .B1(n8869), .B2(n8663), .A(n8541), .ZN(n8542) );
  AOI211_X1 U9919 ( .C1(n9271), .C2(n8670), .A(n8543), .B(n8542), .ZN(n8544)
         );
  OAI21_X1 U9920 ( .B1(n8545), .B2(n8672), .A(n8544), .ZN(P1_U3212) );
  INV_X1 U9921 ( .A(n8547), .ZN(n8549) );
  NAND2_X1 U9922 ( .A1(n8549), .A2(n8548), .ZN(n8551) );
  AOI22_X1 U9923 ( .A1(n8552), .A2(n8546), .B1(n8551), .B2(n8550), .ZN(n8557)
         );
  INV_X1 U9924 ( .A(n9012), .ZN(n9136) );
  AOI22_X1 U9925 ( .A1(n9136), .A2(n8666), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3084), .ZN(n8554) );
  NAND2_X1 U9926 ( .A1(n8655), .A2(n9131), .ZN(n8553) );
  OAI211_X1 U9927 ( .C1(n9006), .C2(n8663), .A(n8554), .B(n8553), .ZN(n8555)
         );
  AOI21_X1 U9928 ( .B1(n9291), .B2(n8670), .A(n8555), .ZN(n8556) );
  OAI21_X1 U9929 ( .B1(n8557), .B2(n8672), .A(n8556), .ZN(P1_U3214) );
  XNOR2_X1 U9930 ( .A(n8560), .B(n8559), .ZN(n8561) );
  XNOR2_X1 U9931 ( .A(n8558), .B(n8561), .ZN(n8566) );
  NAND2_X1 U9932 ( .A1(n8666), .A2(n9149), .ZN(n8562) );
  NAND2_X1 U9933 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n8987) );
  OAI211_X1 U9934 ( .C1(n9217), .C2(n8663), .A(n8562), .B(n8987), .ZN(n8564)
         );
  NOR2_X1 U9935 ( .A1(n7348), .A2(n8658), .ZN(n8563) );
  AOI211_X1 U9936 ( .C1(n9183), .C2(n8655), .A(n8564), .B(n8563), .ZN(n8565)
         );
  OAI21_X1 U9937 ( .B1(n8566), .B2(n8672), .A(n8565), .ZN(P1_U3217) );
  NAND2_X1 U9938 ( .A1(n8615), .A2(n8619), .ZN(n8567) );
  XOR2_X1 U9939 ( .A(n8568), .B(n8567), .Z(n8573) );
  NAND2_X1 U9940 ( .A1(n8655), .A2(n9153), .ZN(n8570) );
  AOI22_X1 U9941 ( .A1(n9150), .A2(n8666), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3084), .ZN(n8569) );
  OAI211_X1 U9942 ( .C1(n9179), .C2(n8663), .A(n8570), .B(n8569), .ZN(n8571)
         );
  AOI21_X1 U9943 ( .B1(n9302), .B2(n8670), .A(n8571), .ZN(n8572) );
  OAI21_X1 U9944 ( .B1(n8573), .B2(n8672), .A(n8572), .ZN(P1_U3221) );
  XOR2_X1 U9945 ( .A(n8575), .B(n8574), .Z(n8581) );
  AOI22_X1 U9946 ( .A1(n9136), .A2(n8621), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3084), .ZN(n8577) );
  NAND2_X1 U9947 ( .A1(n9103), .A2(n4397), .ZN(n8576) );
  OAI211_X1 U9948 ( .C1(n8668), .C2(n8578), .A(n8577), .B(n8576), .ZN(n8579)
         );
  AOI21_X1 U9949 ( .B1(n9281), .B2(n8670), .A(n8579), .ZN(n8580) );
  OAI21_X1 U9950 ( .B1(n8581), .B2(n8672), .A(n8580), .ZN(P1_U3223) );
  INV_X1 U9951 ( .A(n8582), .ZN(n8587) );
  NAND2_X1 U9952 ( .A1(n7443), .A2(n8586), .ZN(n8584) );
  AOI22_X1 U9953 ( .A1(n8587), .A2(n8586), .B1(n8585), .B2(n8584), .ZN(n8593)
         );
  NOR2_X1 U9954 ( .A1(n8663), .A2(n9235), .ZN(n8588) );
  AOI211_X1 U9955 ( .C1(n8666), .C2(n9193), .A(n8589), .B(n8588), .ZN(n8590)
         );
  OAI21_X1 U9956 ( .B1(n8668), .B2(n9224), .A(n8590), .ZN(n8591) );
  AOI21_X1 U9957 ( .B1(n9330), .B2(n8670), .A(n8591), .ZN(n8592) );
  OAI21_X1 U9958 ( .B1(n8593), .B2(n8672), .A(n8592), .ZN(P1_U3224) );
  INV_X1 U9959 ( .A(n9325), .ZN(n9209) );
  OAI21_X1 U9960 ( .B1(n8596), .B2(n8595), .A(n8594), .ZN(n8598) );
  NAND2_X1 U9961 ( .A1(n8598), .A2(n8597), .ZN(n8603) );
  NAND2_X1 U9962 ( .A1(P1_U3084), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n8945) );
  OAI21_X1 U9963 ( .B1(n8599), .B2(n9217), .A(n8945), .ZN(n8601) );
  NOR2_X1 U9964 ( .A1(n8668), .A2(n9210), .ZN(n8600) );
  AOI211_X1 U9965 ( .C1(n8621), .C2(n8932), .A(n8601), .B(n8600), .ZN(n8602)
         );
  OAI211_X1 U9966 ( .C1(n9209), .C2(n8658), .A(n8603), .B(n8602), .ZN(P1_U3226) );
  INV_X1 U9967 ( .A(n8604), .ZN(n8605) );
  AOI21_X1 U9968 ( .B1(n8607), .B2(n8606), .A(n8605), .ZN(n8614) );
  NOR2_X1 U9969 ( .A1(n9013), .A2(n9906), .ZN(n9287) );
  INV_X1 U9970 ( .A(n9010), .ZN(n9115) );
  OAI22_X1 U9971 ( .A1(n9115), .A2(n8663), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8608), .ZN(n8609) );
  AOI21_X1 U9972 ( .B1(n8931), .B2(n4397), .A(n8609), .ZN(n8610) );
  OAI21_X1 U9973 ( .B1(n8668), .B2(n9120), .A(n8610), .ZN(n8611) );
  AOI21_X1 U9974 ( .B1(n9287), .B2(n8612), .A(n8611), .ZN(n8613) );
  OAI21_X1 U9975 ( .B1(n8614), .B2(n8672), .A(n8613), .ZN(P1_U3227) );
  INV_X1 U9976 ( .A(n8615), .ZN(n8620) );
  AOI21_X1 U9977 ( .B1(n8617), .B2(n8619), .A(n8616), .ZN(n8618) );
  AOI21_X1 U9978 ( .B1(n8620), .B2(n8619), .A(n8618), .ZN(n8626) );
  AOI22_X1 U9979 ( .A1(n4397), .A2(n9168), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3084), .ZN(n8623) );
  NAND2_X1 U9980 ( .A1(n8621), .A2(n9192), .ZN(n8622) );
  OAI211_X1 U9981 ( .C1(n8668), .C2(n9162), .A(n8623), .B(n8622), .ZN(n8624)
         );
  AOI21_X1 U9982 ( .B1(n9306), .B2(n8670), .A(n8624), .ZN(n8625) );
  OAI21_X1 U9983 ( .B1(n8626), .B2(n8672), .A(n8625), .ZN(P1_U3231) );
  NAND2_X1 U9984 ( .A1(n8628), .A2(n8627), .ZN(n8629) );
  XOR2_X1 U9985 ( .A(n8630), .B(n8629), .Z(n8638) );
  OAI22_X1 U9986 ( .A1(n8663), .A2(n8632), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8631), .ZN(n8633) );
  AOI21_X1 U9987 ( .B1(n4397), .B2(n9010), .A(n8633), .ZN(n8634) );
  OAI21_X1 U9988 ( .B1(n8668), .B2(n8635), .A(n8634), .ZN(n8636) );
  AOI21_X1 U9989 ( .B1(n9296), .B2(n8670), .A(n8636), .ZN(n8637) );
  OAI21_X1 U9990 ( .B1(n8638), .B2(n8672), .A(n8637), .ZN(P1_U3233) );
  XNOR2_X1 U9991 ( .A(n8640), .B(n8639), .ZN(n8641) );
  XNOR2_X1 U9992 ( .A(n8642), .B(n8641), .ZN(n8648) );
  NAND2_X1 U9993 ( .A1(n8655), .A2(n9200), .ZN(n8645) );
  NOR2_X1 U9994 ( .A1(n8643), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8964) );
  AOI21_X1 U9995 ( .B1(n4397), .B2(n9192), .A(n8964), .ZN(n8644) );
  OAI211_X1 U9996 ( .C1(n9234), .C2(n8663), .A(n8645), .B(n8644), .ZN(n8646)
         );
  AOI21_X1 U9997 ( .B1(n9318), .B2(n8670), .A(n8646), .ZN(n8647) );
  OAI21_X1 U9998 ( .B1(n8648), .B2(n8672), .A(n8647), .ZN(P1_U3236) );
  AOI21_X1 U9999 ( .B1(n8649), .B2(n8650), .A(n8672), .ZN(n8652) );
  NAND2_X1 U10000 ( .A1(n8652), .A2(n8651), .ZN(n8657) );
  INV_X1 U10001 ( .A(n9085), .ZN(n8930) );
  AOI22_X1 U10002 ( .A1(n4397), .A2(n8930), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3084), .ZN(n8653) );
  OAI21_X1 U10003 ( .B1(n9116), .B2(n8663), .A(n8653), .ZN(n8654) );
  AOI21_X1 U10004 ( .B1(n9088), .B2(n8655), .A(n8654), .ZN(n8656) );
  OAI211_X1 U10005 ( .C1(n4698), .C2(n8658), .A(n8657), .B(n8656), .ZN(
        P1_U3238) );
  NAND2_X1 U10006 ( .A1(n8660), .A2(n8659), .ZN(n8661) );
  XOR2_X1 U10007 ( .A(n8662), .B(n8661), .Z(n8673) );
  NOR2_X1 U10008 ( .A1(n8663), .A2(n9243), .ZN(n8664) );
  AOI211_X1 U10009 ( .C1(n4397), .C2(n8932), .A(n8665), .B(n8664), .ZN(n8667)
         );
  OAI21_X1 U10010 ( .B1(n8668), .B2(n9249), .A(n8667), .ZN(n8669) );
  AOI21_X1 U10011 ( .B1(n9335), .B2(n8670), .A(n8669), .ZN(n8671) );
  OAI21_X1 U10012 ( .B1(n8673), .B2(n8672), .A(n8671), .ZN(P1_U3239) );
  INV_X1 U10013 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n8676) );
  NAND2_X1 U10014 ( .A1(n5931), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n8675) );
  NAND2_X1 U10015 ( .A1(n7555), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n8674) );
  OAI211_X1 U10016 ( .C1(n6044), .C2(n8676), .A(n8675), .B(n8674), .ZN(n9036)
         );
  NAND2_X1 U10017 ( .A1(n8677), .A2(n8767), .ZN(n8679) );
  OR2_X1 U10018 ( .A1(n6067), .A2(n9371), .ZN(n8678) );
  AOI21_X1 U10019 ( .B1(n8994), .B2(n9036), .A(n9652), .ZN(n8875) );
  OR2_X1 U10020 ( .A1(n9119), .A2(n9012), .ZN(n8778) );
  OR2_X1 U10021 ( .A1(n9291), .A2(n9115), .ZN(n9027) );
  INV_X1 U10022 ( .A(n8740), .ZN(n8909) );
  NAND2_X1 U10023 ( .A1(n9119), .A2(n9012), .ZN(n9028) );
  NAND2_X1 U10024 ( .A1(n8909), .A2(n9028), .ZN(n8680) );
  NAND2_X1 U10025 ( .A1(n9082), .A2(n8680), .ZN(n8683) );
  NAND2_X1 U10026 ( .A1(n9291), .A2(n9115), .ZN(n8905) );
  AND2_X1 U10027 ( .A1(n9028), .A2(n8905), .ZN(n8739) );
  INV_X1 U10028 ( .A(n8739), .ZN(n8681) );
  NAND2_X1 U10029 ( .A1(n8681), .A2(n8778), .ZN(n8682) );
  NAND2_X1 U10030 ( .A1(n9030), .A2(n8682), .ZN(n8871) );
  INV_X1 U10031 ( .A(n8773), .ZN(n8765) );
  MUX2_X1 U10032 ( .A(n8683), .B(n8871), .S(n8765), .Z(n8742) );
  AND2_X1 U10033 ( .A1(n8726), .A2(n8684), .ZN(n8725) );
  AND2_X1 U10034 ( .A1(n8825), .A2(n8823), .ZN(n8685) );
  MUX2_X1 U10035 ( .A(n8811), .B(n8685), .S(n8765), .Z(n8723) );
  MUX2_X1 U10036 ( .A(n8687), .B(n8686), .S(n8773), .Z(n8689) );
  INV_X1 U10037 ( .A(n8786), .ZN(n8688) );
  NAND2_X1 U10038 ( .A1(n8689), .A2(n8688), .ZN(n8704) );
  NAND3_X1 U10039 ( .A1(n8704), .A2(n8845), .A3(n8842), .ZN(n8690) );
  INV_X1 U10040 ( .A(n8691), .ZN(n8789) );
  NAND2_X1 U10041 ( .A1(n8693), .A2(n8789), .ZN(n8826) );
  INV_X1 U10042 ( .A(n8850), .ZN(n8694) );
  XNOR2_X1 U10043 ( .A(n8692), .B(n8936), .ZN(n9633) );
  OAI211_X1 U10044 ( .C1(n8765), .C2(n8693), .A(n8699), .B(n9633), .ZN(n8709)
         );
  NOR2_X1 U10045 ( .A1(n8697), .A2(n8696), .ZN(n8851) );
  OR3_X1 U10046 ( .A1(n8858), .A2(n8851), .A3(n8765), .ZN(n8711) );
  NAND2_X1 U10047 ( .A1(n8699), .A2(n8698), .ZN(n8828) );
  NAND2_X1 U10048 ( .A1(n8711), .A2(n8828), .ZN(n8700) );
  NAND2_X1 U10049 ( .A1(n8702), .A2(n8701), .ZN(n8715) );
  NAND3_X1 U10050 ( .A1(n8704), .A2(n8839), .A3(n8703), .ZN(n8705) );
  NAND3_X1 U10051 ( .A1(n8705), .A2(n9796), .A3(n8845), .ZN(n8707) );
  NAND3_X1 U10052 ( .A1(n8707), .A2(n8789), .A3(n8706), .ZN(n8708) );
  NAND3_X1 U10053 ( .A1(n8708), .A2(n8850), .A3(n8788), .ZN(n8713) );
  NOR2_X1 U10054 ( .A1(n8709), .A2(n8765), .ZN(n8712) );
  NAND3_X1 U10055 ( .A1(n8857), .A2(n8765), .A3(n8855), .ZN(n8710) );
  AOI22_X1 U10056 ( .A1(n8713), .A2(n8712), .B1(n8711), .B2(n8710), .ZN(n8714)
         );
  NAND2_X1 U10057 ( .A1(n8715), .A2(n8714), .ZN(n8720) );
  AND2_X1 U10058 ( .A1(n8861), .A2(n9229), .ZN(n9240) );
  NAND2_X1 U10059 ( .A1(n8857), .A2(n8855), .ZN(n8829) );
  NAND2_X1 U10060 ( .A1(n8829), .A2(n8716), .ZN(n8718) );
  NAND2_X1 U10061 ( .A1(n8858), .A2(n8857), .ZN(n8717) );
  MUX2_X1 U10062 ( .A(n8718), .B(n8717), .S(n8765), .Z(n8719) );
  MUX2_X1 U10063 ( .A(n8861), .B(n9229), .S(n8765), .Z(n8721) );
  MUX2_X1 U10064 ( .A(n8862), .B(n8822), .S(n8773), .Z(n8722) );
  NAND2_X1 U10065 ( .A1(n8779), .A2(n8812), .ZN(n8724) );
  AOI21_X1 U10066 ( .B1(n8725), .B2(n8727), .A(n8724), .ZN(n8730) );
  AND2_X1 U10067 ( .A1(n8812), .A2(n8825), .ZN(n8728) );
  NAND2_X1 U10068 ( .A1(n9144), .A2(n8726), .ZN(n8810) );
  AOI21_X1 U10069 ( .B1(n8728), .B2(n8727), .A(n8810), .ZN(n8729) );
  MUX2_X1 U10070 ( .A(n8730), .B(n8729), .S(n8773), .Z(n8734) );
  NAND2_X1 U10071 ( .A1(n8816), .A2(n9144), .ZN(n8731) );
  OAI21_X1 U10072 ( .B1(n8734), .B2(n8731), .A(n8736), .ZN(n8733) );
  INV_X1 U10073 ( .A(n8817), .ZN(n8732) );
  INV_X1 U10074 ( .A(n8779), .ZN(n8735) );
  AND2_X1 U10075 ( .A1(n8816), .A2(n8735), .ZN(n8738) );
  INV_X1 U10076 ( .A(n8736), .ZN(n8737) );
  OR3_X1 U10077 ( .A1(n9024), .A2(n8738), .A3(n8737), .ZN(n8821) );
  INV_X1 U10078 ( .A(n8821), .ZN(n8819) );
  NAND2_X1 U10079 ( .A1(n8740), .A2(n8739), .ZN(n8741) );
  INV_X1 U10080 ( .A(n8752), .ZN(n8743) );
  NOR2_X1 U10081 ( .A1(n8743), .A2(n9016), .ZN(n8757) );
  NOR2_X1 U10082 ( .A1(n9030), .A2(n9103), .ZN(n8744) );
  OR2_X1 U10083 ( .A1(n8744), .A2(n9278), .ZN(n8747) );
  AND2_X1 U10084 ( .A1(n9082), .A2(n8869), .ZN(n8745) );
  NOR2_X1 U10085 ( .A1(n9031), .A2(n8745), .ZN(n8746) );
  MUX2_X1 U10086 ( .A(n8747), .B(n8746), .S(n8765), .Z(n8756) );
  NAND2_X1 U10087 ( .A1(n9271), .A2(n9085), .ZN(n8808) );
  NAND2_X1 U10088 ( .A1(n9278), .A2(n9082), .ZN(n8748) );
  NAND2_X1 U10089 ( .A1(n8808), .A2(n8748), .ZN(n8751) );
  NAND2_X1 U10090 ( .A1(n9030), .A2(n9103), .ZN(n8749) );
  NAND2_X1 U10091 ( .A1(n9033), .A2(n8749), .ZN(n8750) );
  MUX2_X1 U10092 ( .A(n8751), .B(n8750), .S(n8773), .Z(n8754) );
  NAND2_X1 U10093 ( .A1(n9073), .A2(n8752), .ZN(n8753) );
  NAND2_X1 U10094 ( .A1(n8754), .A2(n8753), .ZN(n8755) );
  OAI21_X1 U10095 ( .B1(n8757), .B2(n8756), .A(n8755), .ZN(n8760) );
  NAND2_X1 U10096 ( .A1(n9061), .A2(n8758), .ZN(n8809) );
  MUX2_X1 U10097 ( .A(n9033), .B(n8808), .S(n8773), .Z(n8759) );
  NAND3_X1 U10098 ( .A1(n8760), .A2(n9051), .A3(n8759), .ZN(n8762) );
  MUX2_X1 U10099 ( .A(n8809), .B(n9034), .S(n8773), .Z(n8761) );
  NAND2_X1 U10100 ( .A1(n8762), .A2(n8761), .ZN(n8766) );
  INV_X1 U10101 ( .A(n9036), .ZN(n8802) );
  NOR2_X1 U10102 ( .A1(n8990), .A2(n8802), .ZN(n8774) );
  NAND2_X1 U10103 ( .A1(n9363), .A2(n8767), .ZN(n8764) );
  OR2_X1 U10104 ( .A1(n6067), .A2(n5658), .ZN(n8763) );
  OAI21_X1 U10105 ( .B1(n8774), .B2(n8772), .A(n8992), .ZN(n8879) );
  NAND2_X1 U10106 ( .A1(n8768), .A2(n8767), .ZN(n8770) );
  INV_X1 U10107 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n9375) );
  OR2_X1 U10108 ( .A1(n6067), .A2(n9375), .ZN(n8769) );
  NAND2_X1 U10109 ( .A1(n8776), .A2(n8773), .ZN(n8771) );
  INV_X1 U10110 ( .A(n8774), .ZN(n8775) );
  NAND2_X1 U10111 ( .A1(n8776), .A2(n8775), .ZN(n8886) );
  NAND2_X1 U10112 ( .A1(n9042), .A2(n8777), .ZN(n8915) );
  XNOR2_X1 U10113 ( .A(n9291), .B(n9115), .ZN(n9135) );
  NAND2_X1 U10114 ( .A1(n8778), .A2(n9028), .ZN(n9113) );
  NAND2_X1 U10115 ( .A1(n9144), .A2(n8779), .ZN(n9166) );
  NOR4_X1 U10116 ( .A1(n8782), .A2(n4638), .A3(n8781), .A4(n8780), .ZN(n8783)
         );
  NOR4_X1 U10117 ( .A1(n8787), .A2(n8786), .A3(n8785), .A4(n8784), .ZN(n8792)
         );
  AND2_X1 U10118 ( .A1(n8789), .A2(n8788), .ZN(n9799) );
  NAND4_X1 U10119 ( .A1(n8792), .A2(n8791), .A3(n8790), .A4(n9799), .ZN(n8794)
         );
  INV_X1 U10120 ( .A(n9633), .ZN(n9639) );
  NOR4_X1 U10121 ( .A1(n8795), .A2(n8794), .A3(n8793), .A4(n9639), .ZN(n8796)
         );
  NAND4_X1 U10122 ( .A1(n9214), .A2(n9240), .A3(n4642), .A4(n8796), .ZN(n8797)
         );
  NOR4_X1 U10123 ( .A1(n9166), .A2(n9176), .A3(n9195), .A4(n8797), .ZN(n8798)
         );
  NAND3_X1 U10124 ( .A1(n8799), .A2(n9147), .A3(n8798), .ZN(n8800) );
  NOR4_X1 U10125 ( .A1(n9101), .A2(n9135), .A3(n9113), .A4(n8800), .ZN(n8801)
         );
  NAND2_X1 U10126 ( .A1(n9278), .A2(n9103), .ZN(n9017) );
  NAND2_X1 U10127 ( .A1(n9016), .A2(n9017), .ZN(n9083) );
  AND4_X1 U10128 ( .A1(n9051), .A2(n9073), .A3(n8801), .A4(n9083), .ZN(n8803)
         );
  NAND2_X1 U10129 ( .A1(n8990), .A2(n8802), .ZN(n8916) );
  NAND4_X1 U10130 ( .A1(n8877), .A2(n9035), .A3(n8803), .A4(n8916), .ZN(n8804)
         );
  OAI21_X1 U10131 ( .B1(n8886), .B2(n8804), .A(n5842), .ZN(n8806) );
  INV_X1 U10132 ( .A(n8806), .ZN(n8881) );
  NAND2_X1 U10133 ( .A1(n9033), .A2(n9031), .ZN(n8807) );
  AND3_X1 U10134 ( .A1(n8809), .A2(n8808), .A3(n8807), .ZN(n8912) );
  INV_X1 U10135 ( .A(n8810), .ZN(n8815) );
  INV_X1 U10136 ( .A(n8811), .ZN(n8813) );
  NAND3_X1 U10137 ( .A1(n8813), .A2(n8825), .A3(n8812), .ZN(n8814) );
  NAND3_X1 U10138 ( .A1(n8816), .A2(n8815), .A3(n8814), .ZN(n8818) );
  AOI21_X1 U10139 ( .B1(n8819), .B2(n8818), .A(n8817), .ZN(n8908) );
  NOR2_X1 U10140 ( .A1(n8821), .A2(n8820), .ZN(n8904) );
  AND2_X1 U10141 ( .A1(n8823), .A2(n8822), .ZN(n8824) );
  NAND2_X1 U10142 ( .A1(n8825), .A2(n8824), .ZN(n8864) );
  AND2_X1 U10143 ( .A1(n8826), .A2(n8850), .ZN(n8827) );
  NOR2_X1 U10144 ( .A1(n8828), .A2(n8827), .ZN(n8848) );
  INV_X1 U10145 ( .A(n8829), .ZN(n8831) );
  NAND4_X1 U10146 ( .A1(n9229), .A2(n8848), .A3(n8831), .A4(n8830), .ZN(n8832)
         );
  OR2_X1 U10147 ( .A1(n8864), .A2(n8832), .ZN(n8902) );
  NAND2_X1 U10148 ( .A1(n8834), .A2(n8833), .ZN(n8835) );
  NOR2_X1 U10149 ( .A1(n8836), .A2(n8835), .ZN(n8895) );
  NAND2_X1 U10150 ( .A1(n8837), .A2(n8895), .ZN(n8847) );
  INV_X1 U10151 ( .A(n6429), .ZN(n8843) );
  INV_X1 U10152 ( .A(n8838), .ZN(n8840) );
  NAND2_X1 U10153 ( .A1(n8840), .A2(n8839), .ZN(n8841) );
  OAI211_X1 U10154 ( .C1(n8844), .C2(n8843), .A(n8842), .B(n8841), .ZN(n8846)
         );
  INV_X1 U10155 ( .A(n8845), .ZN(n8897) );
  AOI21_X1 U10156 ( .B1(n8847), .B2(n8846), .A(n8897), .ZN(n8865) );
  INV_X1 U10157 ( .A(n8848), .ZN(n8854) );
  AND2_X1 U10158 ( .A1(n8850), .A2(n8849), .ZN(n8853) );
  INV_X1 U10159 ( .A(n8851), .ZN(n8852) );
  OAI21_X1 U10160 ( .B1(n8854), .B2(n8853), .A(n8852), .ZN(n8856) );
  AND2_X1 U10161 ( .A1(n8856), .A2(n8855), .ZN(n8859) );
  OAI211_X1 U10162 ( .C1(n8859), .C2(n8858), .A(n8857), .B(n9229), .ZN(n8860)
         );
  AND3_X1 U10163 ( .A1(n8862), .A2(n8861), .A3(n8860), .ZN(n8863) );
  OR2_X1 U10164 ( .A1(n8864), .A2(n8863), .ZN(n8900) );
  OAI21_X1 U10165 ( .B1(n8902), .B2(n8865), .A(n8900), .ZN(n8866) );
  NAND2_X1 U10166 ( .A1(n8904), .A2(n8866), .ZN(n8867) );
  NAND2_X1 U10167 ( .A1(n8908), .A2(n8867), .ZN(n8868) );
  NOR2_X1 U10168 ( .A1(n8868), .A2(n8909), .ZN(n8872) );
  OR2_X1 U10169 ( .A1(n9278), .A2(n8869), .ZN(n8870) );
  OAI211_X1 U10170 ( .C1(n8872), .C2(n8871), .A(n9033), .B(n9032), .ZN(n8873)
         );
  AND2_X1 U10171 ( .A1(n8912), .A2(n8873), .ZN(n8876) );
  NAND2_X1 U10172 ( .A1(n8874), .A2(n9034), .ZN(n8917) );
  OAI211_X1 U10173 ( .C1(n8876), .C2(n8917), .A(n4593), .B(n8915), .ZN(n8878)
         );
  AOI211_X1 U10174 ( .C1(n8879), .C2(n8878), .A(n5842), .B(n8919), .ZN(n8880)
         );
  NOR2_X1 U10175 ( .A1(n8881), .A2(n8880), .ZN(n8882) );
  NOR3_X1 U10176 ( .A1(n8919), .A2(n5875), .A3(n5842), .ZN(n8883) );
  NAND2_X1 U10177 ( .A1(n8884), .A2(n8883), .ZN(n8885) );
  INV_X1 U10178 ( .A(n8886), .ZN(n8921) );
  NAND2_X1 U10179 ( .A1(n6007), .A2(n6014), .ZN(n8887) );
  NAND3_X1 U10180 ( .A1(n8888), .A2(n5845), .A3(n8887), .ZN(n8890) );
  NAND2_X1 U10181 ( .A1(n8890), .A2(n8889), .ZN(n8892) );
  OAI22_X1 U10182 ( .A1(n8893), .A2(n8892), .B1(n6379), .B2(n8891), .ZN(n8894)
         );
  NAND2_X1 U10183 ( .A1(n8894), .A2(n6429), .ZN(n8896) );
  NAND2_X1 U10184 ( .A1(n8896), .A2(n8895), .ZN(n8899) );
  AOI21_X1 U10185 ( .B1(n8899), .B2(n8898), .A(n8897), .ZN(n8901) );
  OAI21_X1 U10186 ( .B1(n8902), .B2(n8901), .A(n8900), .ZN(n8903) );
  NAND2_X1 U10187 ( .A1(n8904), .A2(n8903), .ZN(n8907) );
  INV_X1 U10188 ( .A(n8905), .ZN(n8906) );
  AOI21_X1 U10189 ( .B1(n8908), .B2(n8907), .A(n8906), .ZN(n8910) );
  OAI211_X1 U10190 ( .C1(n8910), .C2(n8909), .A(n9028), .B(n9030), .ZN(n8911)
         );
  AND3_X1 U10191 ( .A1(n9073), .A2(n9032), .A3(n8911), .ZN(n8914) );
  INV_X1 U10192 ( .A(n8912), .ZN(n8913) );
  NOR2_X1 U10193 ( .A1(n8914), .A2(n8913), .ZN(n8918) );
  OAI211_X1 U10194 ( .C1(n8918), .C2(n8917), .A(n8916), .B(n8915), .ZN(n8920)
         );
  AOI21_X1 U10195 ( .B1(n8921), .B2(n8920), .A(n8919), .ZN(n8922) );
  XNOR2_X1 U10196 ( .A(n8922), .B(n9154), .ZN(n8923) );
  NAND2_X1 U10197 ( .A1(n8923), .A2(n5844), .ZN(n8924) );
  NAND4_X1 U10198 ( .A1(n8926), .A2(n9846), .A3(n9686), .A4(n8925), .ZN(n8927)
         );
  OAI211_X1 U10199 ( .C1(n5875), .C2(n8929), .A(n8927), .B(P1_B_REG_SCAN_IN), 
        .ZN(n8928) );
  MUX2_X1 U10200 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9036), .S(P1_U4006), .Z(
        P1_U3585) );
  MUX2_X1 U10201 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9053), .S(P1_U4006), .Z(
        P1_U3584) );
  MUX2_X1 U10202 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9075), .S(P1_U4006), .Z(
        P1_U3583) );
  MUX2_X1 U10203 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n8930), .S(P1_U4006), .Z(
        P1_U3582) );
  MUX2_X1 U10204 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9103), .S(P1_U4006), .Z(
        P1_U3581) );
  MUX2_X1 U10205 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n8931), .S(P1_U4006), .Z(
        P1_U3580) );
  MUX2_X1 U10206 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9136), .S(P1_U4006), .Z(
        P1_U3579) );
  MUX2_X1 U10207 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9010), .S(P1_U4006), .Z(
        P1_U3578) );
  MUX2_X1 U10208 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9150), .S(P1_U4006), .Z(
        P1_U3577) );
  MUX2_X1 U10209 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9168), .S(P1_U4006), .Z(
        P1_U3576) );
  MUX2_X1 U10210 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9149), .S(P1_U4006), .Z(
        P1_U3575) );
  MUX2_X1 U10211 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9192), .S(P1_U4006), .Z(
        P1_U3574) );
  MUX2_X1 U10212 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9193), .S(P1_U4006), .Z(
        P1_U3572) );
  MUX2_X1 U10213 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n8932), .S(P1_U4006), .Z(
        P1_U3571) );
  MUX2_X1 U10214 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n8933), .S(P1_U4006), .Z(
        P1_U3570) );
  MUX2_X1 U10215 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n4439), .S(P1_U4006), .Z(
        P1_U3569) );
  MUX2_X1 U10216 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n8934), .S(P1_U4006), .Z(
        P1_U3568) );
  MUX2_X1 U10217 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n8935), .S(P1_U4006), .Z(
        P1_U3567) );
  MUX2_X1 U10218 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n8936), .S(P1_U4006), .Z(
        P1_U3566) );
  MUX2_X1 U10219 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n8937), .S(P1_U4006), .Z(
        P1_U3565) );
  MUX2_X1 U10220 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n8938), .S(P1_U4006), .Z(
        P1_U3564) );
  MUX2_X1 U10221 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n8939), .S(P1_U4006), .Z(
        P1_U3563) );
  MUX2_X1 U10222 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n8940), .S(P1_U4006), .Z(
        P1_U3562) );
  MUX2_X1 U10223 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9827), .S(P1_U4006), .Z(
        P1_U3561) );
  MUX2_X1 U10224 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n8941), .S(P1_U4006), .Z(
        P1_U3560) );
  MUX2_X1 U10225 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9826), .S(P1_U4006), .Z(
        P1_U3559) );
  MUX2_X1 U10226 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n8942), .S(P1_U4006), .Z(
        P1_U3558) );
  MUX2_X1 U10227 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n8944), .S(P1_U4006), .Z(
        P1_U3557) );
  MUX2_X1 U10228 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n6007), .S(P1_U4006), .Z(
        P1_U3556) );
  INV_X1 U10229 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n8959) );
  INV_X1 U10230 ( .A(n8945), .ZN(n8950) );
  AOI21_X1 U10231 ( .B1(n8952), .B2(P1_REG1_REG_16__SCAN_IN), .A(n8946), .ZN(
        n8948) );
  XNOR2_X1 U10232 ( .A(n8969), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n8947) );
  NOR2_X1 U10233 ( .A1(n8948), .A2(n8947), .ZN(n8961) );
  AOI211_X1 U10234 ( .C1(n8948), .C2(n8947), .A(n8961), .B(n9744), .ZN(n8949)
         );
  AOI211_X1 U10235 ( .C1(n8969), .C2(n9758), .A(n8950), .B(n8949), .ZN(n8958)
         );
  NAND2_X1 U10236 ( .A1(n8969), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n8953) );
  OAI21_X1 U10237 ( .B1(n8969), .B2(P1_REG2_REG_17__SCAN_IN), .A(n8953), .ZN(
        n8954) );
  AOI211_X1 U10238 ( .C1(n8955), .C2(n8954), .A(n8968), .B(n9774), .ZN(n8956)
         );
  INV_X1 U10239 ( .A(n8956), .ZN(n8957) );
  OAI211_X1 U10240 ( .C1(n8959), .C2(n9785), .A(n8958), .B(n8957), .ZN(
        P1_U3258) );
  INV_X1 U10241 ( .A(n8979), .ZN(n8967) );
  XNOR2_X1 U10242 ( .A(n8979), .B(n8960), .ZN(n8963) );
  AOI21_X1 U10243 ( .B1(n8969), .B2(P1_REG1_REG_17__SCAN_IN), .A(n8961), .ZN(
        n8962) );
  NAND2_X1 U10244 ( .A1(n8963), .A2(n8962), .ZN(n8978) );
  OAI21_X1 U10245 ( .B1(n8963), .B2(n8962), .A(n8978), .ZN(n8965) );
  AOI21_X1 U10246 ( .B1(n9781), .B2(n8965), .A(n8964), .ZN(n8966) );
  OAI21_X1 U10247 ( .B1(n8967), .B2(n9783), .A(n8966), .ZN(n8974) );
  AOI21_X1 U10248 ( .B1(n8969), .B2(P1_REG2_REG_17__SCAN_IN), .A(n8968), .ZN(
        n8972) );
  NAND2_X1 U10249 ( .A1(n8979), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n8970) );
  OAI21_X1 U10250 ( .B1(n8979), .B2(P1_REG2_REG_18__SCAN_IN), .A(n8970), .ZN(
        n8971) );
  NOR2_X1 U10251 ( .A1(n8972), .A2(n8971), .ZN(n8976) );
  AOI211_X1 U10252 ( .C1(n8972), .C2(n8971), .A(n8976), .B(n9774), .ZN(n8973)
         );
  AOI211_X1 U10253 ( .C1(P1_ADDR_REG_18__SCAN_IN), .C2(n9759), .A(n8974), .B(
        n8973), .ZN(n8975) );
  INV_X1 U10254 ( .A(n8975), .ZN(P1_U3259) );
  INV_X1 U10255 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n8989) );
  AOI21_X1 U10256 ( .B1(P1_REG2_REG_18__SCAN_IN), .B2(n8979), .A(n8976), .ZN(
        n8977) );
  XNOR2_X1 U10257 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n8977), .ZN(n8984) );
  INV_X1 U10258 ( .A(n8984), .ZN(n8982) );
  OAI21_X1 U10259 ( .B1(n8979), .B2(P1_REG1_REG_18__SCAN_IN), .A(n8978), .ZN(
        n8980) );
  XNOR2_X1 U10260 ( .A(n8980), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n8983) );
  OAI21_X1 U10261 ( .B1(n8983), .B2(n9744), .A(n9783), .ZN(n8981) );
  AOI21_X1 U10262 ( .B1(n8982), .B2(n9751), .A(n8981), .ZN(n8986) );
  AOI22_X1 U10263 ( .A1(n8984), .A2(n9751), .B1(n9781), .B2(n8983), .ZN(n8985)
         );
  MUX2_X1 U10264 ( .A(n8986), .B(n8985), .S(n9154), .Z(n8988) );
  OAI211_X1 U10265 ( .C1(n8989), .C2(n9785), .A(n8988), .B(n8987), .ZN(
        P1_U3260) );
  INV_X1 U10266 ( .A(n9061), .ZN(n9265) );
  INV_X1 U10267 ( .A(n9291), .ZN(n9133) );
  NOR2_X1 U10268 ( .A1(n8990), .A2(n4329), .ZN(n8991) );
  XNOR2_X1 U10269 ( .A(n8992), .B(n8991), .ZN(n9628) );
  NAND2_X1 U10270 ( .A1(n9628), .A2(n9794), .ZN(n8996) );
  AND2_X1 U10271 ( .A1(n9686), .A2(P1_B_REG_SCAN_IN), .ZN(n8993) );
  NOR2_X1 U10272 ( .A1(n9800), .A2(n8993), .ZN(n9037) );
  NAND2_X1 U10273 ( .A1(n8994), .A2(n9037), .ZN(n9651) );
  NOR2_X1 U10274 ( .A1(n9844), .A2(n9651), .ZN(n8997) );
  AOI21_X1 U10275 ( .B1(n9844), .B2(P1_REG2_REG_31__SCAN_IN), .A(n8997), .ZN(
        n8995) );
  OAI211_X1 U10276 ( .C1(n9626), .C2(n9808), .A(n8996), .B(n8995), .ZN(
        P1_U3261) );
  XNOR2_X1 U10277 ( .A(n9652), .B(n4329), .ZN(n9654) );
  NAND2_X1 U10278 ( .A1(n9654), .A2(n9794), .ZN(n8999) );
  AOI21_X1 U10279 ( .B1(n9844), .B2(P1_REG2_REG_30__SCAN_IN), .A(n8997), .ZN(
        n8998) );
  OAI211_X1 U10280 ( .C1(n9652), .C2(n9808), .A(n8999), .B(n8998), .ZN(
        P1_U3262) );
  NOR2_X1 U10281 ( .A1(n9007), .A2(n9006), .ZN(n9003) );
  INV_X1 U10282 ( .A(n9003), .ZN(n9000) );
  AOI21_X1 U10283 ( .B1(n9005), .B2(n9004), .A(n4818), .ZN(n9125) );
  NAND2_X1 U10284 ( .A1(n9007), .A2(n9006), .ZN(n9126) );
  OR2_X1 U10285 ( .A1(n9291), .A2(n9010), .ZN(n9008) );
  NAND2_X1 U10286 ( .A1(n9125), .A2(n9009), .ZN(n9109) );
  NAND2_X1 U10287 ( .A1(n9291), .A2(n9010), .ZN(n9108) );
  NAND2_X1 U10288 ( .A1(n9109), .A2(n9011), .ZN(n9015) );
  NAND2_X1 U10289 ( .A1(n9013), .A2(n9012), .ZN(n9014) );
  INV_X1 U10290 ( .A(n9067), .ZN(n9019) );
  INV_X1 U10291 ( .A(n9073), .ZN(n9018) );
  NAND2_X1 U10292 ( .A1(n4699), .A2(n9085), .ZN(n9020) );
  INV_X1 U10293 ( .A(n9051), .ZN(n9021) );
  NAND2_X1 U10294 ( .A1(n9061), .A2(n9075), .ZN(n9022) );
  NAND2_X1 U10295 ( .A1(n9049), .A2(n9022), .ZN(n9023) );
  XNOR2_X1 U10296 ( .A(n9023), .B(n9035), .ZN(n9257) );
  INV_X1 U10297 ( .A(n9257), .ZN(n9046) );
  INV_X1 U10298 ( .A(n9024), .ZN(n9025) );
  NAND2_X1 U10299 ( .A1(n9026), .A2(n9025), .ZN(n9134) );
  OAI21_X2 U10300 ( .B1(n9134), .B2(n9135), .A(n9027), .ZN(n9112) );
  INV_X1 U10301 ( .A(n9028), .ZN(n9029) );
  NAND2_X1 U10302 ( .A1(n9074), .A2(n9073), .ZN(n9072) );
  NAND2_X1 U10303 ( .A1(n9072), .A2(n9033), .ZN(n9052) );
  AOI22_X1 U10304 ( .A1(n9037), .A2(n9036), .B1(n9075), .B2(n9825), .ZN(n9038)
         );
  OAI21_X1 U10305 ( .B1(n9258), .B2(n9056), .A(n4329), .ZN(n9259) );
  OAI22_X1 U10306 ( .A1(n9814), .A2(n9040), .B1(n9039), .B2(n9809), .ZN(n9041)
         );
  AOI21_X1 U10307 ( .B1(n9042), .B2(n9174), .A(n9041), .ZN(n9043) );
  OAI21_X1 U10308 ( .B1(n9259), .B2(n9063), .A(n9043), .ZN(n9044) );
  AOI21_X1 U10309 ( .B1(n9261), .B2(n9814), .A(n9044), .ZN(n9045) );
  OAI21_X1 U10310 ( .B1(n9046), .B2(n9256), .A(n9045), .ZN(P1_U3355) );
  NAND2_X1 U10311 ( .A1(n9047), .A2(n9051), .ZN(n9048) );
  INV_X1 U10312 ( .A(n9264), .ZN(n9066) );
  OAI211_X1 U10313 ( .C1(n9052), .C2(n9051), .A(n9050), .B(n9823), .ZN(n9055)
         );
  NAND2_X1 U10314 ( .A1(n9053), .A2(n9828), .ZN(n9054) );
  OAI211_X1 U10315 ( .C1(n9085), .C2(n9802), .A(n9055), .B(n9054), .ZN(n9268)
         );
  INV_X1 U10316 ( .A(n9056), .ZN(n9057) );
  OAI21_X1 U10317 ( .B1(n9265), .B2(n9068), .A(n9057), .ZN(n9266) );
  OAI22_X1 U10318 ( .A1(n9814), .A2(n9059), .B1(n9058), .B2(n9809), .ZN(n9060)
         );
  AOI21_X1 U10319 ( .B1(n9061), .B2(n9174), .A(n9060), .ZN(n9062) );
  OAI21_X1 U10320 ( .B1(n9266), .B2(n9063), .A(n9062), .ZN(n9064) );
  AOI21_X1 U10321 ( .B1(n9268), .B2(n9814), .A(n9064), .ZN(n9065) );
  OAI21_X1 U10322 ( .B1(n9066), .B2(n9256), .A(n9065), .ZN(P1_U3263) );
  XOR2_X1 U10323 ( .A(n9067), .B(n9073), .Z(n9275) );
  AOI21_X1 U10324 ( .B1(n9271), .B2(n9086), .A(n9068), .ZN(n9272) );
  INV_X1 U10325 ( .A(n9069), .ZN(n9070) );
  AOI22_X1 U10326 ( .A1(n9844), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n9838), .B2(
        n9070), .ZN(n9071) );
  OAI21_X1 U10327 ( .B1(n4699), .B2(n9808), .A(n9071), .ZN(n9079) );
  OAI211_X1 U10328 ( .C1(n9074), .C2(n9073), .A(n9072), .B(n9823), .ZN(n9077)
         );
  AOI22_X1 U10329 ( .A1(n9103), .A2(n9825), .B1(n9828), .B2(n9075), .ZN(n9076)
         );
  NOR2_X1 U10330 ( .A1(n9274), .A2(n9844), .ZN(n9078) );
  AOI211_X1 U10331 ( .C1(n9794), .C2(n9272), .A(n9079), .B(n9078), .ZN(n9080)
         );
  OAI21_X1 U10332 ( .B1(n9275), .B2(n9256), .A(n9080), .ZN(P1_U3264) );
  XOR2_X1 U10333 ( .A(n9083), .B(n9081), .Z(n9280) );
  AOI22_X1 U10334 ( .A1(n9278), .A2(n9174), .B1(P1_REG2_REG_26__SCAN_IN), .B2(
        n9844), .ZN(n9093) );
  OAI222_X1 U10335 ( .A1(n9800), .A2(n9085), .B1(n9802), .B2(n9116), .C1(n9084), .C2(n9242), .ZN(n9276) );
  INV_X1 U10336 ( .A(n9086), .ZN(n9087) );
  AOI211_X1 U10337 ( .C1(n9278), .C2(n9095), .A(n9908), .B(n9087), .ZN(n9277)
         );
  INV_X1 U10338 ( .A(n9277), .ZN(n9090) );
  INV_X1 U10339 ( .A(n9088), .ZN(n9089) );
  OAI22_X1 U10340 ( .A1(n9090), .A2(n9840), .B1(n9809), .B2(n9089), .ZN(n9091)
         );
  OAI21_X1 U10341 ( .B1(n9276), .B2(n9091), .A(n9814), .ZN(n9092) );
  OAI211_X1 U10342 ( .C1(n9280), .C2(n9256), .A(n9093), .B(n9092), .ZN(
        P1_U3265) );
  XOR2_X1 U10343 ( .A(n9101), .B(n9094), .Z(n9285) );
  INV_X1 U10344 ( .A(n9117), .ZN(n9097) );
  INV_X1 U10345 ( .A(n9095), .ZN(n9096) );
  AOI21_X1 U10346 ( .B1(n9281), .B2(n9097), .A(n9096), .ZN(n9282) );
  AOI22_X1 U10347 ( .A1(n9098), .A2(n9838), .B1(P1_REG2_REG_25__SCAN_IN), .B2(
        n9844), .ZN(n9099) );
  OAI21_X1 U10348 ( .B1(n9100), .B2(n9808), .A(n9099), .ZN(n9106) );
  XNOR2_X1 U10349 ( .A(n9102), .B(n9101), .ZN(n9104) );
  AOI222_X1 U10350 ( .A1(n9823), .A2(n9104), .B1(n9103), .B2(n9828), .C1(n9136), .C2(n9825), .ZN(n9284) );
  NOR2_X1 U10351 ( .A1(n9284), .A2(n9844), .ZN(n9105) );
  AOI211_X1 U10352 ( .C1(n9282), .C2(n9794), .A(n9106), .B(n9105), .ZN(n9107)
         );
  OAI21_X1 U10353 ( .B1(n9285), .B2(n9256), .A(n9107), .ZN(P1_U3266) );
  NAND2_X1 U10354 ( .A1(n9109), .A2(n9108), .ZN(n9110) );
  XNOR2_X1 U10355 ( .A(n9110), .B(n9113), .ZN(n9290) );
  AOI22_X1 U10356 ( .A1(n9119), .A2(n9174), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n9844), .ZN(n9124) );
  AOI21_X1 U10357 ( .B1(n9113), .B2(n9112), .A(n9111), .ZN(n9114) );
  OAI222_X1 U10358 ( .A1(n9800), .A2(n9116), .B1(n9802), .B2(n9115), .C1(n9242), .C2(n9114), .ZN(n9288) );
  INV_X1 U10359 ( .A(n9129), .ZN(n9118) );
  AOI211_X1 U10360 ( .C1(n9119), .C2(n9118), .A(n9908), .B(n9117), .ZN(n9286)
         );
  INV_X1 U10361 ( .A(n9286), .ZN(n9121) );
  OAI22_X1 U10362 ( .A1(n9121), .A2(n9840), .B1(n9809), .B2(n9120), .ZN(n9122)
         );
  OAI21_X1 U10363 ( .B1(n9288), .B2(n9122), .A(n9814), .ZN(n9123) );
  OAI211_X1 U10364 ( .C1(n9290), .C2(n9256), .A(n9124), .B(n9123), .ZN(
        P1_U3267) );
  NAND2_X1 U10365 ( .A1(n9125), .A2(n9126), .ZN(n9127) );
  XOR2_X1 U10366 ( .A(n9135), .B(n9127), .Z(n9295) );
  INV_X1 U10367 ( .A(n9128), .ZN(n9130) );
  AOI21_X1 U10368 ( .B1(n9291), .B2(n9130), .A(n9129), .ZN(n9292) );
  AOI22_X1 U10369 ( .A1(n9844), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n9131), .B2(
        n9838), .ZN(n9132) );
  OAI21_X1 U10370 ( .B1(n9133), .B2(n9808), .A(n9132), .ZN(n9139) );
  XOR2_X1 U10371 ( .A(n9135), .B(n9134), .Z(n9137) );
  AOI222_X1 U10372 ( .A1(n9823), .A2(n9137), .B1(n9150), .B2(n9825), .C1(n9136), .C2(n9828), .ZN(n9294) );
  NOR2_X1 U10373 ( .A1(n9294), .A2(n9844), .ZN(n9138) );
  AOI211_X1 U10374 ( .C1(n9292), .C2(n9794), .A(n9139), .B(n9138), .ZN(n9140)
         );
  OAI21_X1 U10375 ( .B1(n9295), .B2(n9256), .A(n9140), .ZN(P1_U3268) );
  NAND2_X1 U10376 ( .A1(n9005), .A2(n9141), .ZN(n9143) );
  XNOR2_X1 U10377 ( .A(n9143), .B(n9142), .ZN(n9305) );
  AOI22_X1 U10378 ( .A1(n9302), .A2(n9174), .B1(P1_REG2_REG_21__SCAN_IN), .B2(
        n9844), .ZN(n9158) );
  AND2_X1 U10379 ( .A1(n9145), .A2(n9144), .ZN(n9148) );
  OAI21_X1 U10380 ( .B1(n9148), .B2(n9147), .A(n9146), .ZN(n9151) );
  AOI222_X1 U10381 ( .A1(n9823), .A2(n9151), .B1(n9150), .B2(n9828), .C1(n9149), .C2(n9825), .ZN(n9304) );
  AOI211_X1 U10382 ( .C1(n9302), .C2(n9160), .A(n9908), .B(n4691), .ZN(n9301)
         );
  AOI22_X1 U10383 ( .A1(n9301), .A2(n9154), .B1(n9838), .B2(n9153), .ZN(n9155)
         );
  AOI21_X1 U10384 ( .B1(n9304), .B2(n9155), .A(n9844), .ZN(n9156) );
  INV_X1 U10385 ( .A(n9156), .ZN(n9157) );
  OAI211_X1 U10386 ( .C1(n9305), .C2(n9256), .A(n9158), .B(n9157), .ZN(
        P1_U3270) );
  XNOR2_X1 U10387 ( .A(n9159), .B(n9166), .ZN(n9310) );
  INV_X1 U10388 ( .A(n9160), .ZN(n9161) );
  AOI21_X1 U10389 ( .B1(n9306), .B2(n9180), .A(n9161), .ZN(n9307) );
  INV_X1 U10390 ( .A(n9306), .ZN(n9165) );
  INV_X1 U10391 ( .A(n9162), .ZN(n9163) );
  AOI22_X1 U10392 ( .A1(n9844), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9163), .B2(
        n9838), .ZN(n9164) );
  OAI21_X1 U10393 ( .B1(n9165), .B2(n9808), .A(n9164), .ZN(n9171) );
  XNOR2_X1 U10394 ( .A(n9167), .B(n9166), .ZN(n9169) );
  AOI222_X1 U10395 ( .A1(n9823), .A2(n9169), .B1(n9192), .B2(n9825), .C1(n9168), .C2(n9828), .ZN(n9309) );
  NOR2_X1 U10396 ( .A1(n9309), .A2(n9844), .ZN(n9170) );
  AOI211_X1 U10397 ( .C1(n9307), .C2(n9794), .A(n9171), .B(n9170), .ZN(n9172)
         );
  OAI21_X1 U10398 ( .B1(n9310), .B2(n9256), .A(n9172), .ZN(P1_U3271) );
  XNOR2_X1 U10399 ( .A(n9173), .B(n9176), .ZN(n9315) );
  AOI22_X1 U10400 ( .A1(n9313), .A2(n9174), .B1(P1_REG2_REG_19__SCAN_IN), .B2(
        n9844), .ZN(n9188) );
  AOI21_X1 U10401 ( .B1(n9177), .B2(n9176), .A(n9175), .ZN(n9178) );
  OAI222_X1 U10402 ( .A1(n9802), .A2(n9217), .B1(n9800), .B2(n9179), .C1(n9242), .C2(n9178), .ZN(n9311) );
  INV_X1 U10403 ( .A(n9198), .ZN(n9182) );
  INV_X1 U10404 ( .A(n9180), .ZN(n9181) );
  AOI211_X1 U10405 ( .C1(n9313), .C2(n9182), .A(n9908), .B(n9181), .ZN(n9312)
         );
  INV_X1 U10406 ( .A(n9312), .ZN(n9185) );
  INV_X1 U10407 ( .A(n9183), .ZN(n9184) );
  OAI22_X1 U10408 ( .A1(n9185), .A2(n9840), .B1(n9809), .B2(n9184), .ZN(n9186)
         );
  OAI21_X1 U10409 ( .B1(n9311), .B2(n9186), .A(n9814), .ZN(n9187) );
  OAI211_X1 U10410 ( .C1(n9315), .C2(n9256), .A(n9188), .B(n9187), .ZN(
        P1_U3272) );
  NAND2_X1 U10411 ( .A1(n9190), .A2(n9189), .ZN(n9191) );
  XNOR2_X1 U10412 ( .A(n9191), .B(n9195), .ZN(n9194) );
  AOI222_X1 U10413 ( .A1(n9823), .A2(n9194), .B1(n9193), .B2(n9825), .C1(n9192), .C2(n9828), .ZN(n9321) );
  OR2_X1 U10414 ( .A1(n9196), .A2(n9195), .ZN(n9317) );
  INV_X1 U10415 ( .A(n9256), .ZN(n9197) );
  NAND3_X1 U10416 ( .A1(n9317), .A2(n9316), .A3(n9197), .ZN(n9205) );
  INV_X1 U10417 ( .A(n9207), .ZN(n9199) );
  AOI21_X1 U10418 ( .B1(n9318), .B2(n9199), .A(n9198), .ZN(n9319) );
  AOI22_X1 U10419 ( .A1(n9844), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9200), .B2(
        n9838), .ZN(n9201) );
  OAI21_X1 U10420 ( .B1(n9202), .B2(n9808), .A(n9201), .ZN(n9203) );
  AOI21_X1 U10421 ( .B1(n9319), .B2(n9794), .A(n9203), .ZN(n9204) );
  OAI211_X1 U10422 ( .C1(n9844), .C2(n9321), .A(n9205), .B(n9204), .ZN(
        P1_U3273) );
  XNOR2_X1 U10423 ( .A(n9206), .B(n9214), .ZN(n9327) );
  AOI211_X1 U10424 ( .C1(n9325), .C2(n9222), .A(n9908), .B(n9207), .ZN(n9324)
         );
  INV_X1 U10425 ( .A(n9208), .ZN(n9248) );
  NOR2_X1 U10426 ( .A1(n9209), .A2(n9808), .ZN(n9213) );
  OAI22_X1 U10427 ( .A1(n9814), .A2(n9211), .B1(n9210), .B2(n9809), .ZN(n9212)
         );
  AOI211_X1 U10428 ( .C1(n9324), .C2(n9248), .A(n9213), .B(n9212), .ZN(n9219)
         );
  XNOR2_X1 U10429 ( .A(n9215), .B(n9214), .ZN(n9216) );
  OAI222_X1 U10430 ( .A1(n9802), .A2(n9244), .B1(n9800), .B2(n9217), .C1(n9216), .C2(n9242), .ZN(n9323) );
  NAND2_X1 U10431 ( .A1(n9323), .A2(n9814), .ZN(n9218) );
  OAI211_X1 U10432 ( .C1(n9327), .C2(n9256), .A(n9219), .B(n9218), .ZN(
        P1_U3274) );
  XNOR2_X1 U10433 ( .A(n9221), .B(n9220), .ZN(n9332) );
  AOI211_X1 U10434 ( .C1(n9330), .C2(n9246), .A(n9908), .B(n4684), .ZN(n9329)
         );
  INV_X1 U10435 ( .A(n9330), .ZN(n9223) );
  NOR2_X1 U10436 ( .A1(n9223), .A2(n9808), .ZN(n9227) );
  OAI22_X1 U10437 ( .A1(n9814), .A2(n9225), .B1(n9224), .B2(n9809), .ZN(n9226)
         );
  AOI211_X1 U10438 ( .C1(n9329), .C2(n9228), .A(n9227), .B(n9226), .ZN(n9237)
         );
  NOR2_X1 U10439 ( .A1(n4642), .A2(n4641), .ZN(n9232) );
  AOI21_X1 U10440 ( .B1(n9232), .B2(n9231), .A(n9230), .ZN(n9233) );
  OAI222_X1 U10441 ( .A1(n9802), .A2(n9235), .B1(n9800), .B2(n9234), .C1(n9242), .C2(n9233), .ZN(n9328) );
  NAND2_X1 U10442 ( .A1(n9328), .A2(n9814), .ZN(n9236) );
  OAI211_X1 U10443 ( .C1(n9332), .C2(n9256), .A(n9237), .B(n9236), .ZN(
        P1_U3275) );
  XNOR2_X1 U10444 ( .A(n9238), .B(n9240), .ZN(n9337) );
  XOR2_X1 U10445 ( .A(n9240), .B(n9239), .Z(n9241) );
  OAI222_X1 U10446 ( .A1(n9800), .A2(n9244), .B1(n9802), .B2(n9243), .C1(n9242), .C2(n9241), .ZN(n9333) );
  INV_X1 U10447 ( .A(n9245), .ZN(n9247) );
  AOI211_X1 U10448 ( .C1(n9335), .C2(n9247), .A(n9908), .B(n4685), .ZN(n9334)
         );
  NAND2_X1 U10449 ( .A1(n9334), .A2(n9248), .ZN(n9252) );
  INV_X1 U10450 ( .A(n9249), .ZN(n9250) );
  AOI22_X1 U10451 ( .A1(n9844), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n9250), .B2(
        n9838), .ZN(n9251) );
  OAI211_X1 U10452 ( .C1(n9253), .C2(n9808), .A(n9252), .B(n9251), .ZN(n9254)
         );
  AOI21_X1 U10453 ( .B1(n9333), .B2(n9814), .A(n9254), .ZN(n9255) );
  OAI21_X1 U10454 ( .B1(n9337), .B2(n9256), .A(n9255), .ZN(P1_U3276) );
  NAND2_X1 U10455 ( .A1(n9257), .A2(n9895), .ZN(n9263) );
  OAI22_X1 U10456 ( .A1(n9259), .A2(n9908), .B1(n9258), .B2(n9906), .ZN(n9260)
         );
  NOR2_X1 U10457 ( .A1(n9261), .A2(n9260), .ZN(n9262) );
  NAND2_X1 U10458 ( .A1(n9263), .A2(n9262), .ZN(n9346) );
  MUX2_X1 U10459 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9346), .S(n9928), .Z(
        P1_U3552) );
  NAND2_X1 U10460 ( .A1(n9264), .A2(n9895), .ZN(n9270) );
  OAI22_X1 U10461 ( .A1(n9266), .A2(n9908), .B1(n9265), .B2(n9906), .ZN(n9267)
         );
  NOR2_X1 U10462 ( .A1(n9268), .A2(n9267), .ZN(n9269) );
  NAND2_X1 U10463 ( .A1(n9270), .A2(n9269), .ZN(n9347) );
  MUX2_X1 U10464 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9347), .S(n9928), .Z(
        P1_U3551) );
  AOI22_X1 U10465 ( .A1(n9272), .A2(n9881), .B1(n9271), .B2(n9664), .ZN(n9273)
         );
  OAI211_X1 U10466 ( .C1(n9275), .C2(n9897), .A(n9274), .B(n9273), .ZN(n9348)
         );
  MUX2_X1 U10467 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9348), .S(n9928), .Z(
        P1_U3550) );
  OAI21_X1 U10468 ( .B1(n9280), .B2(n9897), .A(n9279), .ZN(n9349) );
  MUX2_X1 U10469 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9349), .S(n9928), .Z(
        P1_U3549) );
  AOI22_X1 U10470 ( .A1(n9282), .A2(n9881), .B1(n9281), .B2(n9664), .ZN(n9283)
         );
  OAI211_X1 U10471 ( .C1(n9285), .C2(n9897), .A(n9284), .B(n9283), .ZN(n9350)
         );
  MUX2_X1 U10472 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9350), .S(n9928), .Z(
        P1_U3548) );
  NOR3_X1 U10473 ( .A1(n9288), .A2(n9287), .A3(n9286), .ZN(n9289) );
  OAI21_X1 U10474 ( .B1(n9290), .B2(n9897), .A(n9289), .ZN(n9351) );
  MUX2_X1 U10475 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9351), .S(n9928), .Z(
        P1_U3547) );
  AOI22_X1 U10476 ( .A1(n9292), .A2(n9881), .B1(n9291), .B2(n9664), .ZN(n9293)
         );
  OAI211_X1 U10477 ( .C1(n9295), .C2(n9897), .A(n9294), .B(n9293), .ZN(n9352)
         );
  MUX2_X1 U10478 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9352), .S(n9928), .Z(
        P1_U3546) );
  AOI22_X1 U10479 ( .A1(n9297), .A2(n9881), .B1(n9296), .B2(n9664), .ZN(n9298)
         );
  OAI211_X1 U10480 ( .C1(n9300), .C2(n9897), .A(n9299), .B(n9298), .ZN(n9353)
         );
  MUX2_X1 U10481 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9353), .S(n9928), .Z(
        P1_U3545) );
  AOI21_X1 U10482 ( .B1(n9302), .B2(n9664), .A(n9301), .ZN(n9303) );
  OAI211_X1 U10483 ( .C1(n9305), .C2(n9897), .A(n9304), .B(n9303), .ZN(n9354)
         );
  MUX2_X1 U10484 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9354), .S(n9928), .Z(
        P1_U3544) );
  AOI22_X1 U10485 ( .A1(n9307), .A2(n9881), .B1(n9306), .B2(n9664), .ZN(n9308)
         );
  OAI211_X1 U10486 ( .C1(n9310), .C2(n9897), .A(n9309), .B(n9308), .ZN(n9355)
         );
  MUX2_X1 U10487 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9355), .S(n9928), .Z(
        P1_U3543) );
  AOI211_X1 U10488 ( .C1(n9313), .C2(n9664), .A(n9312), .B(n9311), .ZN(n9314)
         );
  OAI21_X1 U10489 ( .B1(n9315), .B2(n9897), .A(n9314), .ZN(n9356) );
  MUX2_X1 U10490 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9356), .S(n9928), .Z(
        P1_U3542) );
  NAND3_X1 U10491 ( .A1(n9317), .A2(n9316), .A3(n9895), .ZN(n9322) );
  AOI22_X1 U10492 ( .A1(n9319), .A2(n9881), .B1(n9318), .B2(n9664), .ZN(n9320)
         );
  NAND3_X1 U10493 ( .A1(n9322), .A2(n9321), .A3(n9320), .ZN(n9357) );
  MUX2_X1 U10494 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9357), .S(n9928), .Z(
        P1_U3541) );
  AOI211_X1 U10495 ( .C1(n9325), .C2(n9664), .A(n9324), .B(n9323), .ZN(n9326)
         );
  OAI21_X1 U10496 ( .B1(n9327), .B2(n9897), .A(n9326), .ZN(n9358) );
  MUX2_X1 U10497 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9358), .S(n9928), .Z(
        P1_U3540) );
  AOI211_X1 U10498 ( .C1(n9330), .C2(n9664), .A(n9329), .B(n9328), .ZN(n9331)
         );
  OAI21_X1 U10499 ( .B1(n9332), .B2(n9897), .A(n9331), .ZN(n9359) );
  MUX2_X1 U10500 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9359), .S(n9928), .Z(
        P1_U3539) );
  AOI211_X1 U10501 ( .C1(n9335), .C2(n9664), .A(n9334), .B(n9333), .ZN(n9336)
         );
  OAI21_X1 U10502 ( .B1(n9337), .B2(n9897), .A(n9336), .ZN(n9360) );
  MUX2_X1 U10503 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n9360), .S(n9928), .Z(
        P1_U3538) );
  AOI21_X1 U10504 ( .B1(n9339), .B2(n9664), .A(n9338), .ZN(n9340) );
  OAI211_X1 U10505 ( .C1(n9342), .C2(n9897), .A(n9341), .B(n9340), .ZN(n9361)
         );
  MUX2_X1 U10506 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n9361), .S(n9928), .Z(
        P1_U3537) );
  OAI21_X1 U10507 ( .B1(n9345), .B2(n9344), .A(n9343), .ZN(n9362) );
  MUX2_X1 U10508 ( .A(P1_REG1_REG_0__SCAN_IN), .B(n9362), .S(n9928), .Z(
        P1_U3523) );
  MUX2_X1 U10509 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9346), .S(n9916), .Z(
        P1_U3520) );
  MUX2_X1 U10510 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9347), .S(n9916), .Z(
        P1_U3519) );
  MUX2_X1 U10511 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9348), .S(n9916), .Z(
        P1_U3518) );
  MUX2_X1 U10512 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9349), .S(n9916), .Z(
        P1_U3517) );
  MUX2_X1 U10513 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9350), .S(n9916), .Z(
        P1_U3516) );
  MUX2_X1 U10514 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9351), .S(n9916), .Z(
        P1_U3515) );
  MUX2_X1 U10515 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9352), .S(n9916), .Z(
        P1_U3514) );
  MUX2_X1 U10516 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9353), .S(n9916), .Z(
        P1_U3513) );
  MUX2_X1 U10517 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9354), .S(n9916), .Z(
        P1_U3512) );
  MUX2_X1 U10518 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9355), .S(n9916), .Z(
        P1_U3511) );
  MUX2_X1 U10519 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9356), .S(n9916), .Z(
        P1_U3510) );
  MUX2_X1 U10520 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9357), .S(n9916), .Z(
        P1_U3508) );
  MUX2_X1 U10521 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9358), .S(n9916), .Z(
        P1_U3505) );
  MUX2_X1 U10522 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9359), .S(n9916), .Z(
        P1_U3502) );
  MUX2_X1 U10523 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n9360), .S(n9916), .Z(
        P1_U3499) );
  MUX2_X1 U10524 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n9361), .S(n9916), .Z(
        P1_U3496) );
  MUX2_X1 U10525 ( .A(P1_REG0_REG_0__SCAN_IN), .B(n9362), .S(n9916), .Z(
        P1_U3454) );
  INV_X1 U10526 ( .A(n9363), .ZN(n9368) );
  NOR4_X1 U10527 ( .A1(n9364), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3084), .A4(
        n5944), .ZN(n9365) );
  AOI21_X1 U10528 ( .B1(n9366), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9365), .ZN(
        n9367) );
  OAI21_X1 U10529 ( .B1(n9368), .B2(n9373), .A(n9367), .ZN(P1_U3322) );
  OAI222_X1 U10530 ( .A1(n9376), .A2(n9371), .B1(n9373), .B2(n9370), .C1(
        P1_U3084), .C2(n9369), .ZN(P1_U3323) );
  OAI222_X1 U10531 ( .A1(n9376), .A2(n9375), .B1(n9374), .B2(P1_U3084), .C1(
        n9373), .C2(n9372), .ZN(P1_U3324) );
  MUX2_X1 U10532 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9377), .S(P1_U3084), .Z(
        P1_U3353) );
  INV_X1 U10533 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10070) );
  NOR2_X1 U10534 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n9378) );
  AOI21_X1 U10535 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n9378), .ZN(n10040) );
  NOR2_X1 U10536 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n9379) );
  AOI21_X1 U10537 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n9379), .ZN(n10043) );
  NOR2_X1 U10538 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n9380) );
  AOI21_X1 U10539 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n9380), .ZN(n10046) );
  NOR2_X1 U10540 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n9381) );
  AOI21_X1 U10541 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n9381), .ZN(n10049) );
  NOR2_X1 U10542 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n9382) );
  AOI21_X1 U10543 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n9382), .ZN(n10052) );
  INV_X1 U10544 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n10076) );
  NOR2_X1 U10545 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n9388) );
  XNOR2_X1 U10546 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10081) );
  NAND2_X1 U10547 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n9386) );
  XOR2_X1 U10548 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10079) );
  NAND2_X1 U10549 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n9384) );
  XOR2_X1 U10550 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(P1_ADDR_REG_2__SCAN_IN), .Z(
        n10066) );
  AOI21_X1 U10551 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10034) );
  INV_X1 U10552 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n9603) );
  NAND3_X1 U10553 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n10036) );
  OAI21_X1 U10554 ( .B1(n10034), .B2(n9603), .A(n10036), .ZN(n10065) );
  NAND2_X1 U10555 ( .A1(n10066), .A2(n10065), .ZN(n9383) );
  NAND2_X1 U10556 ( .A1(n9384), .A2(n9383), .ZN(n10078) );
  NAND2_X1 U10557 ( .A1(n10079), .A2(n10078), .ZN(n9385) );
  NAND2_X1 U10558 ( .A1(n9386), .A2(n9385), .ZN(n10080) );
  NOR2_X1 U10559 ( .A1(n10081), .A2(n10080), .ZN(n9387) );
  NOR2_X1 U10560 ( .A1(n9388), .A2(n9387), .ZN(n10075) );
  NAND2_X1 U10561 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n10075), .ZN(n9389) );
  NOR2_X1 U10562 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n10075), .ZN(n10074) );
  AOI21_X1 U10563 ( .B1(n10076), .B2(n9389), .A(n10074), .ZN(n9390) );
  NAND2_X1 U10564 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(n9390), .ZN(n9392) );
  XOR2_X1 U10565 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(n9390), .Z(n10073) );
  NAND2_X1 U10566 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(n10073), .ZN(n9391) );
  NAND2_X1 U10567 ( .A1(n9392), .A2(n9391), .ZN(n9393) );
  NAND2_X1 U10568 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n9393), .ZN(n9395) );
  XOR2_X1 U10569 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n9393), .Z(n10072) );
  NAND2_X1 U10570 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n10072), .ZN(n9394) );
  NAND2_X1 U10571 ( .A1(n9395), .A2(n9394), .ZN(n9396) );
  NAND2_X1 U10572 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n9396), .ZN(n9398) );
  XOR2_X1 U10573 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n9396), .Z(n10067) );
  NAND2_X1 U10574 ( .A1(n10067), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n9397) );
  NAND2_X1 U10575 ( .A1(n9398), .A2(n9397), .ZN(n9399) );
  AND2_X1 U10576 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n9399), .ZN(n9400) );
  XNOR2_X1 U10577 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n9399), .ZN(n10064) );
  INV_X1 U10578 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10063) );
  NOR2_X1 U10579 ( .A1(n10064), .A2(n10063), .ZN(n10062) );
  NOR2_X1 U10580 ( .A1(n9400), .A2(n10062), .ZN(n10061) );
  NAND2_X1 U10581 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n9401) );
  OAI21_X1 U10582 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n9401), .ZN(n10060) );
  NOR2_X1 U10583 ( .A1(n10061), .A2(n10060), .ZN(n10059) );
  AOI21_X1 U10584 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10059), .ZN(n10058) );
  NAND2_X1 U10585 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n9402) );
  OAI21_X1 U10586 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n9402), .ZN(n10057) );
  NOR2_X1 U10587 ( .A1(n10058), .A2(n10057), .ZN(n10056) );
  AOI21_X1 U10588 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10056), .ZN(n10055) );
  NOR2_X1 U10589 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n9403) );
  AOI21_X1 U10590 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n9403), .ZN(n10054) );
  NAND2_X1 U10591 ( .A1(n10055), .A2(n10054), .ZN(n10053) );
  OAI21_X1 U10592 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10053), .ZN(n10051) );
  NAND2_X1 U10593 ( .A1(n10052), .A2(n10051), .ZN(n10050) );
  OAI21_X1 U10594 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10050), .ZN(n10048) );
  NAND2_X1 U10595 ( .A1(n10049), .A2(n10048), .ZN(n10047) );
  OAI21_X1 U10596 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10047), .ZN(n10045) );
  NAND2_X1 U10597 ( .A1(n10046), .A2(n10045), .ZN(n10044) );
  OAI21_X1 U10598 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10044), .ZN(n10042) );
  NAND2_X1 U10599 ( .A1(n10043), .A2(n10042), .ZN(n10041) );
  OAI21_X1 U10600 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10041), .ZN(n10039) );
  NAND2_X1 U10601 ( .A1(n10040), .A2(n10039), .ZN(n10038) );
  OAI21_X1 U10602 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10038), .ZN(n10069) );
  NOR2_X1 U10603 ( .A1(n10070), .A2(n10069), .ZN(n9404) );
  NAND2_X1 U10604 ( .A1(n10070), .A2(n10069), .ZN(n10068) );
  OAI21_X1 U10605 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n9404), .A(n10068), .ZN(
        n9591) );
  AOI22_X1 U10606 ( .A1(P2_REG3_REG_24__SCAN_IN), .A2(keyinput_f51), .B1(
        SI_14_), .B2(keyinput_f18), .ZN(n9405) );
  OAI221_X1 U10607 ( .B1(P2_REG3_REG_24__SCAN_IN), .B2(keyinput_f51), .C1(
        SI_14_), .C2(keyinput_f18), .A(n9405), .ZN(n9412) );
  AOI22_X1 U10608 ( .A1(SI_31_), .A2(keyinput_f1), .B1(P2_REG3_REG_12__SCAN_IN), .B2(keyinput_f46), .ZN(n9406) );
  OAI221_X1 U10609 ( .B1(SI_31_), .B2(keyinput_f1), .C1(
        P2_REG3_REG_12__SCAN_IN), .C2(keyinput_f46), .A(n9406), .ZN(n9411) );
  AOI22_X1 U10610 ( .A1(SI_15_), .A2(keyinput_f17), .B1(SI_26_), .B2(
        keyinput_f6), .ZN(n9407) );
  OAI221_X1 U10611 ( .B1(SI_15_), .B2(keyinput_f17), .C1(SI_26_), .C2(
        keyinput_f6), .A(n9407), .ZN(n9410) );
  AOI22_X1 U10612 ( .A1(SI_24_), .A2(keyinput_f8), .B1(SI_25_), .B2(
        keyinput_f7), .ZN(n9408) );
  OAI221_X1 U10613 ( .B1(SI_24_), .B2(keyinput_f8), .C1(SI_25_), .C2(
        keyinput_f7), .A(n9408), .ZN(n9409) );
  NOR4_X1 U10614 ( .A1(n9412), .A2(n9411), .A3(n9410), .A4(n9409), .ZN(n9439)
         );
  XOR2_X1 U10615 ( .A(SI_20_), .B(keyinput_f12), .Z(n9419) );
  AOI22_X1 U10616 ( .A1(P2_REG3_REG_23__SCAN_IN), .A2(keyinput_f38), .B1(
        P2_REG3_REG_28__SCAN_IN), .B2(keyinput_f42), .ZN(n9413) );
  OAI221_X1 U10617 ( .B1(P2_REG3_REG_23__SCAN_IN), .B2(keyinput_f38), .C1(
        P2_REG3_REG_28__SCAN_IN), .C2(keyinput_f42), .A(n9413), .ZN(n9418) );
  AOI22_X1 U10618 ( .A1(P2_REG3_REG_1__SCAN_IN), .A2(keyinput_f44), .B1(SI_16_), .B2(keyinput_f16), .ZN(n9414) );
  OAI221_X1 U10619 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(keyinput_f44), .C1(
        SI_16_), .C2(keyinput_f16), .A(n9414), .ZN(n9417) );
  AOI22_X1 U10620 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(keyinput_f56), .B1(
        P2_REG3_REG_22__SCAN_IN), .B2(keyinput_f57), .ZN(n9415) );
  OAI221_X1 U10621 ( .B1(P2_REG3_REG_13__SCAN_IN), .B2(keyinput_f56), .C1(
        P2_REG3_REG_22__SCAN_IN), .C2(keyinput_f57), .A(n9415), .ZN(n9416) );
  NOR4_X1 U10622 ( .A1(n9419), .A2(n9418), .A3(n9417), .A4(n9416), .ZN(n9438)
         );
  AOI22_X1 U10623 ( .A1(P2_WR_REG_SCAN_IN), .A2(keyinput_f0), .B1(
        P2_REG3_REG_15__SCAN_IN), .B2(keyinput_f63), .ZN(n9420) );
  OAI221_X1 U10624 ( .B1(P2_WR_REG_SCAN_IN), .B2(keyinput_f0), .C1(
        P2_REG3_REG_15__SCAN_IN), .C2(keyinput_f63), .A(n9420), .ZN(n9427) );
  AOI22_X1 U10625 ( .A1(SI_30_), .A2(keyinput_f2), .B1(SI_13_), .B2(
        keyinput_f19), .ZN(n9421) );
  OAI221_X1 U10626 ( .B1(SI_30_), .B2(keyinput_f2), .C1(SI_13_), .C2(
        keyinput_f19), .A(n9421), .ZN(n9426) );
  INV_X1 U10627 ( .A(SI_18_), .ZN(n9577) );
  AOI22_X1 U10628 ( .A1(SI_9_), .A2(keyinput_f23), .B1(n9577), .B2(
        keyinput_f14), .ZN(n9422) );
  OAI221_X1 U10629 ( .B1(SI_9_), .B2(keyinput_f23), .C1(n9577), .C2(
        keyinput_f14), .A(n9422), .ZN(n9425) );
  AOI22_X1 U10630 ( .A1(SI_10_), .A2(keyinput_f22), .B1(P2_RD_REG_SCAN_IN), 
        .B2(keyinput_f33), .ZN(n9423) );
  OAI221_X1 U10631 ( .B1(SI_10_), .B2(keyinput_f22), .C1(P2_RD_REG_SCAN_IN), 
        .C2(keyinput_f33), .A(n9423), .ZN(n9424) );
  NOR4_X1 U10632 ( .A1(n9427), .A2(n9426), .A3(n9425), .A4(n9424), .ZN(n9437)
         );
  AOI22_X1 U10633 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(keyinput_f40), .B1(SI_4_), 
        .B2(keyinput_f28), .ZN(n9428) );
  OAI221_X1 U10634 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(keyinput_f40), .C1(SI_4_), .C2(keyinput_f28), .A(n9428), .ZN(n9435) );
  AOI22_X1 U10635 ( .A1(P2_REG3_REG_26__SCAN_IN), .A2(keyinput_f62), .B1(
        SI_23_), .B2(keyinput_f9), .ZN(n9429) );
  OAI221_X1 U10636 ( .B1(P2_REG3_REG_26__SCAN_IN), .B2(keyinput_f62), .C1(
        SI_23_), .C2(keyinput_f9), .A(n9429), .ZN(n9434) );
  AOI22_X1 U10637 ( .A1(SI_5_), .A2(keyinput_f27), .B1(SI_8_), .B2(
        keyinput_f24), .ZN(n9430) );
  OAI221_X1 U10638 ( .B1(SI_5_), .B2(keyinput_f27), .C1(SI_8_), .C2(
        keyinput_f24), .A(n9430), .ZN(n9433) );
  AOI22_X1 U10639 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(keyinput_f61), .B1(
        P2_REG3_REG_27__SCAN_IN), .B2(keyinput_f36), .ZN(n9431) );
  OAI221_X1 U10640 ( .B1(P2_REG3_REG_6__SCAN_IN), .B2(keyinput_f61), .C1(
        P2_REG3_REG_27__SCAN_IN), .C2(keyinput_f36), .A(n9431), .ZN(n9432) );
  NOR4_X1 U10641 ( .A1(n9435), .A2(n9434), .A3(n9433), .A4(n9432), .ZN(n9436)
         );
  NAND4_X1 U10642 ( .A1(n9439), .A2(n9438), .A3(n9437), .A4(n9436), .ZN(n9493)
         );
  AOI22_X1 U10643 ( .A1(n9441), .A2(keyinput_f10), .B1(keyinput_f39), .B2(
        n9540), .ZN(n9440) );
  OAI221_X1 U10644 ( .B1(n9441), .B2(keyinput_f10), .C1(n9540), .C2(
        keyinput_f39), .A(n9440), .ZN(n9450) );
  AOI22_X1 U10645 ( .A1(n9557), .A2(keyinput_f43), .B1(P2_U3152), .B2(
        keyinput_f34), .ZN(n9442) );
  OAI221_X1 U10646 ( .B1(n9557), .B2(keyinput_f43), .C1(P2_U3152), .C2(
        keyinput_f34), .A(n9442), .ZN(n9449) );
  AOI22_X1 U10647 ( .A1(n9444), .A2(keyinput_f48), .B1(keyinput_f53), .B2(
        n5291), .ZN(n9443) );
  OAI221_X1 U10648 ( .B1(n9444), .B2(keyinput_f48), .C1(n5291), .C2(
        keyinput_f53), .A(n9443), .ZN(n9448) );
  AOI22_X1 U10649 ( .A1(n9446), .A2(keyinput_f59), .B1(n5311), .B2(
        keyinput_f58), .ZN(n9445) );
  OAI221_X1 U10650 ( .B1(n9446), .B2(keyinput_f59), .C1(n5311), .C2(
        keyinput_f58), .A(n9445), .ZN(n9447) );
  NOR4_X1 U10651 ( .A1(n9450), .A2(n9449), .A3(n9448), .A4(n9447), .ZN(n9491)
         );
  AOI22_X1 U10652 ( .A1(n9452), .A2(keyinput_f4), .B1(keyinput_f49), .B2(n5257), .ZN(n9451) );
  OAI221_X1 U10653 ( .B1(n9452), .B2(keyinput_f4), .C1(n5257), .C2(
        keyinput_f49), .A(n9451), .ZN(n9462) );
  AOI22_X1 U10654 ( .A1(n9455), .A2(keyinput_f45), .B1(keyinput_f60), .B2(
        n9454), .ZN(n9453) );
  OAI221_X1 U10655 ( .B1(n9455), .B2(keyinput_f45), .C1(n9454), .C2(
        keyinput_f60), .A(n9453), .ZN(n9461) );
  INV_X1 U10656 ( .A(SI_21_), .ZN(n9549) );
  AOI22_X1 U10657 ( .A1(n9572), .A2(keyinput_f52), .B1(n9549), .B2(
        keyinput_f11), .ZN(n9456) );
  OAI221_X1 U10658 ( .B1(n9572), .B2(keyinput_f52), .C1(n9549), .C2(
        keyinput_f11), .A(n9456), .ZN(n9460) );
  AOI22_X1 U10659 ( .A1(n5273), .A2(keyinput_f35), .B1(n9458), .B2(
        keyinput_f26), .ZN(n9457) );
  OAI221_X1 U10660 ( .B1(n5273), .B2(keyinput_f35), .C1(n9458), .C2(
        keyinput_f26), .A(n9457), .ZN(n9459) );
  NOR4_X1 U10661 ( .A1(n9462), .A2(n9461), .A3(n9460), .A4(n9459), .ZN(n9490)
         );
  AOI22_X1 U10662 ( .A1(n9465), .A2(keyinput_f37), .B1(n9464), .B2(
        keyinput_f29), .ZN(n9463) );
  OAI221_X1 U10663 ( .B1(n9465), .B2(keyinput_f37), .C1(n9464), .C2(
        keyinput_f29), .A(n9463), .ZN(n9476) );
  AOI22_X1 U10664 ( .A1(n4448), .A2(keyinput_f30), .B1(keyinput_f54), .B2(
        n9467), .ZN(n9466) );
  OAI221_X1 U10665 ( .B1(n4448), .B2(keyinput_f30), .C1(n9467), .C2(
        keyinput_f54), .A(n9466), .ZN(n9475) );
  AOI22_X1 U10666 ( .A1(n9470), .A2(keyinput_f13), .B1(keyinput_f20), .B2(
        n9469), .ZN(n9468) );
  OAI221_X1 U10667 ( .B1(n9470), .B2(keyinput_f13), .C1(n9469), .C2(
        keyinput_f20), .A(n9468), .ZN(n9474) );
  INV_X1 U10668 ( .A(SI_7_), .ZN(n9472) );
  AOI22_X1 U10669 ( .A1(n5358), .A2(keyinput_f50), .B1(n9472), .B2(
        keyinput_f25), .ZN(n9471) );
  OAI221_X1 U10670 ( .B1(n5358), .B2(keyinput_f50), .C1(n9472), .C2(
        keyinput_f25), .A(n9471), .ZN(n9473) );
  NOR4_X1 U10671 ( .A1(n9476), .A2(n9475), .A3(n9474), .A4(n9473), .ZN(n9489)
         );
  AOI22_X1 U10672 ( .A1(n4887), .A2(keyinput_f15), .B1(n9548), .B2(keyinput_f5), .ZN(n9477) );
  OAI221_X1 U10673 ( .B1(n4887), .B2(keyinput_f15), .C1(n9548), .C2(
        keyinput_f5), .A(n9477), .ZN(n9487) );
  AOI22_X1 U10674 ( .A1(n5376), .A2(keyinput_f41), .B1(n9479), .B2(
        keyinput_f47), .ZN(n9478) );
  OAI221_X1 U10675 ( .B1(n5376), .B2(keyinput_f41), .C1(n9479), .C2(
        keyinput_f47), .A(n9478), .ZN(n9486) );
  AOI22_X1 U10676 ( .A1(n9481), .A2(keyinput_f55), .B1(n9539), .B2(
        keyinput_f32), .ZN(n9480) );
  OAI221_X1 U10677 ( .B1(n9481), .B2(keyinput_f55), .C1(n9539), .C2(
        keyinput_f32), .A(n9480), .ZN(n9485) );
  XNOR2_X1 U10678 ( .A(SI_1_), .B(keyinput_f31), .ZN(n9483) );
  XNOR2_X1 U10679 ( .A(SI_29_), .B(keyinput_f3), .ZN(n9482) );
  NAND2_X1 U10680 ( .A1(n9483), .A2(n9482), .ZN(n9484) );
  NOR4_X1 U10681 ( .A1(n9487), .A2(n9486), .A3(n9485), .A4(n9484), .ZN(n9488)
         );
  NAND4_X1 U10682 ( .A1(n9491), .A2(n9490), .A3(n9489), .A4(n9488), .ZN(n9492)
         );
  OAI22_X1 U10683 ( .A1(n9493), .A2(n9492), .B1(keyinput_f21), .B2(SI_11_), 
        .ZN(n9494) );
  AOI21_X1 U10684 ( .B1(keyinput_f21), .B2(SI_11_), .A(n9494), .ZN(n9589) );
  AOI22_X1 U10685 ( .A1(P2_REG3_REG_25__SCAN_IN), .A2(keyinput_g47), .B1(
        SI_10_), .B2(keyinput_g22), .ZN(n9495) );
  OAI221_X1 U10686 ( .B1(P2_REG3_REG_25__SCAN_IN), .B2(keyinput_g47), .C1(
        SI_10_), .C2(keyinput_g22), .A(n9495), .ZN(n9502) );
  AOI22_X1 U10687 ( .A1(P2_REG3_REG_26__SCAN_IN), .A2(keyinput_g62), .B1(SI_6_), .B2(keyinput_g26), .ZN(n9496) );
  OAI221_X1 U10688 ( .B1(P2_REG3_REG_26__SCAN_IN), .B2(keyinput_g62), .C1(
        SI_6_), .C2(keyinput_g26), .A(n9496), .ZN(n9501) );
  AOI22_X1 U10689 ( .A1(SI_13_), .A2(keyinput_g19), .B1(SI_24_), .B2(
        keyinput_g8), .ZN(n9497) );
  OAI221_X1 U10690 ( .B1(SI_13_), .B2(keyinput_g19), .C1(SI_24_), .C2(
        keyinput_g8), .A(n9497), .ZN(n9500) );
  AOI22_X1 U10691 ( .A1(SI_30_), .A2(keyinput_g2), .B1(SI_7_), .B2(
        keyinput_g25), .ZN(n9498) );
  OAI221_X1 U10692 ( .B1(SI_30_), .B2(keyinput_g2), .C1(SI_7_), .C2(
        keyinput_g25), .A(n9498), .ZN(n9499) );
  NOR4_X1 U10693 ( .A1(n9502), .A2(n9501), .A3(n9500), .A4(n9499), .ZN(n9529)
         );
  XOR2_X1 U10694 ( .A(SI_16_), .B(keyinput_g16), .Z(n9509) );
  AOI22_X1 U10695 ( .A1(P2_REG3_REG_22__SCAN_IN), .A2(keyinput_g57), .B1(
        P2_STATE_REG_SCAN_IN), .B2(keyinput_g34), .ZN(n9503) );
  OAI221_X1 U10696 ( .B1(P2_REG3_REG_22__SCAN_IN), .B2(keyinput_g57), .C1(
        P2_STATE_REG_SCAN_IN), .C2(keyinput_g34), .A(n9503), .ZN(n9508) );
  AOI22_X1 U10697 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(keyinput_g60), .B1(
        P2_RD_REG_SCAN_IN), .B2(keyinput_g33), .ZN(n9504) );
  OAI221_X1 U10698 ( .B1(P2_REG3_REG_18__SCAN_IN), .B2(keyinput_g60), .C1(
        P2_RD_REG_SCAN_IN), .C2(keyinput_g33), .A(n9504), .ZN(n9507) );
  AOI22_X1 U10699 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(keyinput_g49), .B1(
        P2_REG3_REG_23__SCAN_IN), .B2(keyinput_g38), .ZN(n9505) );
  OAI221_X1 U10700 ( .B1(P2_REG3_REG_5__SCAN_IN), .B2(keyinput_g49), .C1(
        P2_REG3_REG_23__SCAN_IN), .C2(keyinput_g38), .A(n9505), .ZN(n9506) );
  NOR4_X1 U10701 ( .A1(n9509), .A2(n9508), .A3(n9507), .A4(n9506), .ZN(n9528)
         );
  AOI22_X1 U10702 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(keyinput_g37), .B1(SI_1_), .B2(keyinput_g31), .ZN(n9510) );
  OAI221_X1 U10703 ( .B1(P2_REG3_REG_14__SCAN_IN), .B2(keyinput_g37), .C1(
        SI_1_), .C2(keyinput_g31), .A(n9510), .ZN(n9517) );
  AOI22_X1 U10704 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(keyinput_g53), .B1(
        P2_REG3_REG_28__SCAN_IN), .B2(keyinput_g42), .ZN(n9511) );
  OAI221_X1 U10705 ( .B1(P2_REG3_REG_9__SCAN_IN), .B2(keyinput_g53), .C1(
        P2_REG3_REG_28__SCAN_IN), .C2(keyinput_g42), .A(n9511), .ZN(n9516) );
  AOI22_X1 U10706 ( .A1(P2_REG3_REG_21__SCAN_IN), .A2(keyinput_g45), .B1(
        SI_23_), .B2(keyinput_g9), .ZN(n9512) );
  OAI221_X1 U10707 ( .B1(P2_REG3_REG_21__SCAN_IN), .B2(keyinput_g45), .C1(
        SI_23_), .C2(keyinput_g9), .A(n9512), .ZN(n9515) );
  AOI22_X1 U10708 ( .A1(SI_28_), .A2(keyinput_g4), .B1(SI_22_), .B2(
        keyinput_g10), .ZN(n9513) );
  OAI221_X1 U10709 ( .B1(SI_28_), .B2(keyinput_g4), .C1(SI_22_), .C2(
        keyinput_g10), .A(n9513), .ZN(n9514) );
  NOR4_X1 U10710 ( .A1(n9517), .A2(n9516), .A3(n9515), .A4(n9514), .ZN(n9527)
         );
  AOI22_X1 U10711 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(keyinput_g61), .B1(
        P2_REG3_REG_19__SCAN_IN), .B2(keyinput_g41), .ZN(n9518) );
  OAI221_X1 U10712 ( .B1(P2_REG3_REG_6__SCAN_IN), .B2(keyinput_g61), .C1(
        P2_REG3_REG_19__SCAN_IN), .C2(keyinput_g41), .A(n9518), .ZN(n9525) );
  AOI22_X1 U10713 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(keyinput_g48), .B1(
        SI_12_), .B2(keyinput_g20), .ZN(n9519) );
  OAI221_X1 U10714 ( .B1(P2_REG3_REG_16__SCAN_IN), .B2(keyinput_g48), .C1(
        SI_12_), .C2(keyinput_g20), .A(n9519), .ZN(n9524) );
  AOI22_X1 U10715 ( .A1(P2_REG3_REG_0__SCAN_IN), .A2(keyinput_g54), .B1(
        P2_REG3_REG_20__SCAN_IN), .B2(keyinput_g55), .ZN(n9520) );
  OAI221_X1 U10716 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(keyinput_g54), .C1(
        P2_REG3_REG_20__SCAN_IN), .C2(keyinput_g55), .A(n9520), .ZN(n9523) );
  AOI22_X1 U10717 ( .A1(SI_3_), .A2(keyinput_g29), .B1(SI_17_), .B2(
        keyinput_g15), .ZN(n9521) );
  OAI221_X1 U10718 ( .B1(SI_3_), .B2(keyinput_g29), .C1(SI_17_), .C2(
        keyinput_g15), .A(n9521), .ZN(n9522) );
  NOR4_X1 U10719 ( .A1(n9525), .A2(n9524), .A3(n9523), .A4(n9522), .ZN(n9526)
         );
  NAND4_X1 U10720 ( .A1(n9529), .A2(n9528), .A3(n9527), .A4(n9526), .ZN(n9587)
         );
  AOI22_X1 U10721 ( .A1(n9531), .A2(keyinput_g46), .B1(n4448), .B2(
        keyinput_g30), .ZN(n9530) );
  OAI221_X1 U10722 ( .B1(n9531), .B2(keyinput_g46), .C1(n4448), .C2(
        keyinput_g30), .A(n9530), .ZN(n9544) );
  AOI22_X1 U10723 ( .A1(n9534), .A2(keyinput_g40), .B1(n9533), .B2(
        keyinput_g28), .ZN(n9532) );
  OAI221_X1 U10724 ( .B1(n9534), .B2(keyinput_g40), .C1(n9533), .C2(
        keyinput_g28), .A(n9532), .ZN(n9543) );
  AOI22_X1 U10725 ( .A1(n9537), .A2(keyinput_g17), .B1(keyinput_g36), .B2(
        n9536), .ZN(n9535) );
  OAI221_X1 U10726 ( .B1(n9537), .B2(keyinput_g17), .C1(n9536), .C2(
        keyinput_g36), .A(n9535), .ZN(n9542) );
  AOI22_X1 U10727 ( .A1(n9540), .A2(keyinput_g39), .B1(n9539), .B2(
        keyinput_g32), .ZN(n9538) );
  OAI221_X1 U10728 ( .B1(n9540), .B2(keyinput_g39), .C1(n9539), .C2(
        keyinput_g32), .A(n9538), .ZN(n9541) );
  NOR4_X1 U10729 ( .A1(n9544), .A2(n9543), .A3(n9542), .A4(n9541), .ZN(n9585)
         );
  AOI22_X1 U10730 ( .A1(P2_REG3_REG_24__SCAN_IN), .A2(keyinput_g51), .B1(
        SI_19_), .B2(keyinput_g13), .ZN(n9545) );
  OAI221_X1 U10731 ( .B1(P2_REG3_REG_24__SCAN_IN), .B2(keyinput_g51), .C1(
        SI_19_), .C2(keyinput_g13), .A(n9545), .ZN(n9555) );
  AOI22_X1 U10732 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(keyinput_g50), .B1(
        SI_25_), .B2(keyinput_g7), .ZN(n9546) );
  OAI221_X1 U10733 ( .B1(P2_REG3_REG_17__SCAN_IN), .B2(keyinput_g50), .C1(
        SI_25_), .C2(keyinput_g7), .A(n9546), .ZN(n9554) );
  AOI22_X1 U10734 ( .A1(n9549), .A2(keyinput_g11), .B1(n9548), .B2(keyinput_g5), .ZN(n9547) );
  OAI221_X1 U10735 ( .B1(n9549), .B2(keyinput_g11), .C1(n9548), .C2(
        keyinput_g5), .A(n9547), .ZN(n9553) );
  AOI22_X1 U10736 ( .A1(P2_REG3_REG_2__SCAN_IN), .A2(keyinput_g59), .B1(n9551), 
        .B2(keyinput_g3), .ZN(n9550) );
  OAI221_X1 U10737 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(keyinput_g59), .C1(n9551), .C2(keyinput_g3), .A(n9550), .ZN(n9552) );
  NOR4_X1 U10738 ( .A1(n9555), .A2(n9554), .A3(n9553), .A4(n9552), .ZN(n9584)
         );
  AOI22_X1 U10739 ( .A1(n9557), .A2(keyinput_g43), .B1(n4873), .B2(
        keyinput_g18), .ZN(n9556) );
  OAI221_X1 U10740 ( .B1(n9557), .B2(keyinput_g43), .C1(n4873), .C2(
        keyinput_g18), .A(n9556), .ZN(n9566) );
  AOI22_X1 U10741 ( .A1(n5326), .A2(keyinput_g56), .B1(keyinput_g1), .B2(n4949), .ZN(n9558) );
  OAI221_X1 U10742 ( .B1(n5326), .B2(keyinput_g56), .C1(n4949), .C2(
        keyinput_g1), .A(n9558), .ZN(n9565) );
  AOI22_X1 U10743 ( .A1(n5311), .A2(keyinput_g58), .B1(keyinput_g44), .B2(
        n9560), .ZN(n9559) );
  OAI221_X1 U10744 ( .B1(n5311), .B2(keyinput_g58), .C1(n9560), .C2(
        keyinput_g44), .A(n9559), .ZN(n9564) );
  AOI22_X1 U10745 ( .A1(n9562), .A2(keyinput_g24), .B1(keyinput_g35), .B2(
        n5273), .ZN(n9561) );
  OAI221_X1 U10746 ( .B1(n9562), .B2(keyinput_g24), .C1(n5273), .C2(
        keyinput_g35), .A(n9561), .ZN(n9563) );
  NOR4_X1 U10747 ( .A1(n9566), .A2(n9565), .A3(n9564), .A4(n9563), .ZN(n9583)
         );
  AOI22_X1 U10748 ( .A1(n9569), .A2(keyinput_g6), .B1(keyinput_g27), .B2(n9568), .ZN(n9567) );
  OAI221_X1 U10749 ( .B1(n9569), .B2(keyinput_g6), .C1(n9568), .C2(
        keyinput_g27), .A(n9567), .ZN(n9581) );
  AOI22_X1 U10750 ( .A1(n9572), .A2(keyinput_g52), .B1(n9571), .B2(
        keyinput_g12), .ZN(n9570) );
  OAI221_X1 U10751 ( .B1(n9572), .B2(keyinput_g52), .C1(n9571), .C2(
        keyinput_g12), .A(n9570), .ZN(n9580) );
  AOI22_X1 U10752 ( .A1(n7108), .A2(keyinput_g63), .B1(n9574), .B2(
        keyinput_g23), .ZN(n9573) );
  OAI221_X1 U10753 ( .B1(n7108), .B2(keyinput_g63), .C1(n9574), .C2(
        keyinput_g23), .A(n9573), .ZN(n9579) );
  INV_X1 U10754 ( .A(P2_WR_REG_SCAN_IN), .ZN(n9576) );
  AOI22_X1 U10755 ( .A1(n9577), .A2(keyinput_g14), .B1(keyinput_g0), .B2(n9576), .ZN(n9575) );
  OAI221_X1 U10756 ( .B1(n9577), .B2(keyinput_g14), .C1(n9576), .C2(
        keyinput_g0), .A(n9575), .ZN(n9578) );
  NOR4_X1 U10757 ( .A1(n9581), .A2(n9580), .A3(n9579), .A4(n9578), .ZN(n9582)
         );
  NAND4_X1 U10758 ( .A1(n9585), .A2(n9584), .A3(n9583), .A4(n9582), .ZN(n9586)
         );
  OAI22_X1 U10759 ( .A1(SI_11_), .A2(keyinput_g21), .B1(n9587), .B2(n9586), 
        .ZN(n9588) );
  AOI211_X1 U10760 ( .C1(SI_11_), .C2(keyinput_g21), .A(n9589), .B(n9588), 
        .ZN(n9590) );
  XNOR2_X1 U10761 ( .A(n9591), .B(n9590), .ZN(n9595) );
  NOR2_X1 U10762 ( .A1(n9593), .A2(n9592), .ZN(n9594) );
  XOR2_X1 U10763 ( .A(n9595), .B(n9594), .Z(ADD_1071_U4) );
  INV_X1 U10764 ( .A(n9596), .ZN(n9600) );
  NAND2_X1 U10765 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n9597) );
  NAND2_X1 U10766 ( .A1(n9598), .A2(n9597), .ZN(n9599) );
  NAND3_X1 U10767 ( .A1(n9930), .A2(n9600), .A3(n9599), .ZN(n9602) );
  NAND2_X1 U10768 ( .A1(P2_U3152), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n9601) );
  OAI211_X1 U10769 ( .C1(n9604), .C2(n9603), .A(n9602), .B(n9601), .ZN(n9605)
         );
  AOI21_X1 U10770 ( .B1(n9606), .B2(n9619), .A(n9605), .ZN(n9612) );
  NOR2_X1 U10771 ( .A1(n9938), .A2(n9607), .ZN(n9610) );
  OAI211_X1 U10772 ( .C1(n9610), .C2(n9609), .A(n9929), .B(n9608), .ZN(n9611)
         );
  NAND2_X1 U10773 ( .A1(n9612), .A2(n9611), .ZN(P2_U3246) );
  AOI22_X1 U10774 ( .A1(n9935), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n9625) );
  AOI211_X1 U10775 ( .C1(n9616), .C2(n9615), .A(n9614), .B(n9613), .ZN(n9617)
         );
  AOI21_X1 U10776 ( .B1(n9619), .B2(n9618), .A(n9617), .ZN(n9624) );
  OAI211_X1 U10777 ( .C1(n9622), .C2(n9621), .A(n9929), .B(n9620), .ZN(n9623)
         );
  NAND3_X1 U10778 ( .A1(n9625), .A2(n9624), .A3(n9623), .ZN(P2_U3247) );
  OAI21_X1 U10779 ( .B1(n9626), .B2(n9906), .A(n9651), .ZN(n9627) );
  AOI21_X1 U10780 ( .B1(n9881), .B2(n9628), .A(n9627), .ZN(n9630) );
  AOI22_X1 U10781 ( .A1(n9928), .A2(n9630), .B1(n5753), .B2(n9926), .ZN(
        P1_U3554) );
  INV_X1 U10782 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n9629) );
  AOI22_X1 U10783 ( .A1(n9916), .A2(n9630), .B1(n9629), .B2(n9914), .ZN(
        P1_U3522) );
  INV_X1 U10784 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n9631) );
  AOI22_X1 U10785 ( .A1(n10033), .A2(n9632), .B1(n9631), .B2(n10030), .ZN(
        P2_U3551) );
  XNOR2_X1 U10786 ( .A(n9634), .B(n9633), .ZN(n9645) );
  INV_X1 U10787 ( .A(n9645), .ZN(n9676) );
  OR2_X1 U10788 ( .A1(n9635), .A2(n9672), .ZN(n9636) );
  NAND2_X1 U10789 ( .A1(n9637), .A2(n9636), .ZN(n9673) );
  INV_X1 U10790 ( .A(n9673), .ZN(n9638) );
  AOI22_X1 U10791 ( .A1(n9676), .A2(n9795), .B1(n9794), .B2(n9638), .ZN(n9650)
         );
  XNOR2_X1 U10792 ( .A(n9640), .B(n9639), .ZN(n9643) );
  OAI22_X1 U10793 ( .A1(n9801), .A2(n9802), .B1(n9641), .B2(n9800), .ZN(n9642)
         );
  AOI21_X1 U10794 ( .B1(n9643), .B2(n9823), .A(n9642), .ZN(n9644) );
  OAI21_X1 U10795 ( .B1(n9645), .B2(n9884), .A(n9644), .ZN(n9674) );
  NOR2_X1 U10796 ( .A1(n9672), .A2(n9808), .ZN(n9648) );
  OAI22_X1 U10797 ( .A1(n9814), .A2(n5986), .B1(n9646), .B2(n9809), .ZN(n9647)
         );
  AOI211_X1 U10798 ( .C1(n9674), .C2(n9814), .A(n9648), .B(n9647), .ZN(n9649)
         );
  NAND2_X1 U10799 ( .A1(n9650), .A2(n9649), .ZN(P1_U3280) );
  OAI21_X1 U10800 ( .B1(n9652), .B2(n9906), .A(n9651), .ZN(n9653) );
  AOI21_X1 U10801 ( .B1(n9654), .B2(n9881), .A(n9653), .ZN(n9679) );
  AOI22_X1 U10802 ( .A1(n9928), .A2(n9679), .B1(n8676), .B2(n9926), .ZN(
        P1_U3553) );
  INV_X1 U10803 ( .A(n9667), .ZN(n9913) );
  INV_X1 U10804 ( .A(n9655), .ZN(n9660) );
  OAI22_X1 U10805 ( .A1(n9657), .A2(n9908), .B1(n9656), .B2(n9906), .ZN(n9659)
         );
  AOI211_X1 U10806 ( .C1(n9913), .C2(n9660), .A(n9659), .B(n9658), .ZN(n9681)
         );
  AOI22_X1 U10807 ( .A1(n9928), .A2(n9681), .B1(n9661), .B2(n9926), .ZN(
        P1_U3536) );
  INV_X1 U10808 ( .A(n9668), .ZN(n9670) );
  AOI211_X1 U10809 ( .C1(n9665), .C2(n9664), .A(n9663), .B(n9662), .ZN(n9666)
         );
  OAI21_X1 U10810 ( .B1(n9668), .B2(n9667), .A(n9666), .ZN(n9669) );
  AOI21_X1 U10811 ( .B1(n9671), .B2(n9670), .A(n9669), .ZN(n9683) );
  AOI22_X1 U10812 ( .A1(n9928), .A2(n9683), .B1(n7078), .B2(n9926), .ZN(
        P1_U3535) );
  OAI22_X1 U10813 ( .A1(n9673), .A2(n9908), .B1(n9672), .B2(n9906), .ZN(n9675)
         );
  AOI211_X1 U10814 ( .C1(n9913), .C2(n9676), .A(n9675), .B(n9674), .ZN(n9685)
         );
  AOI22_X1 U10815 ( .A1(n9928), .A2(n9685), .B1(n9677), .B2(n9926), .ZN(
        P1_U3534) );
  INV_X1 U10816 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9678) );
  AOI22_X1 U10817 ( .A1(n9916), .A2(n9679), .B1(n9678), .B2(n9914), .ZN(
        P1_U3521) );
  INV_X1 U10818 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n9680) );
  AOI22_X1 U10819 ( .A1(n9916), .A2(n9681), .B1(n9680), .B2(n9914), .ZN(
        P1_U3493) );
  INV_X1 U10820 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n9682) );
  AOI22_X1 U10821 ( .A1(n9916), .A2(n9683), .B1(n9682), .B2(n9914), .ZN(
        P1_U3490) );
  INV_X1 U10822 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n9684) );
  AOI22_X1 U10823 ( .A1(n9916), .A2(n9685), .B1(n9684), .B2(n9914), .ZN(
        P1_U3487) );
  XNOR2_X1 U10824 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  INV_X1 U10825 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n9691) );
  OAI21_X1 U10826 ( .B1(n9686), .B2(P1_REG1_REG_0__SCAN_IN), .A(n9691), .ZN(
        n9689) );
  AOI211_X1 U10827 ( .C1(n9690), .C2(n9689), .A(n9688), .B(n9687), .ZN(n9696)
         );
  NOR3_X1 U10828 ( .A1(n9744), .A2(P1_REG1_REG_0__SCAN_IN), .A3(n9691), .ZN(
        n9694) );
  INV_X1 U10829 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n9692) );
  NOR2_X1 U10830 ( .A1(n9785), .A2(n9692), .ZN(n9693) );
  AOI211_X1 U10831 ( .C1(n9696), .C2(n9695), .A(n9694), .B(n9693), .ZN(n9697)
         );
  OAI21_X1 U10832 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n5665), .A(n9697), .ZN(
        P1_U3241) );
  INV_X1 U10833 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9713) );
  OAI21_X1 U10834 ( .B1(n9700), .B2(n9699), .A(n9698), .ZN(n9702) );
  AOI22_X1 U10835 ( .A1(n9751), .A2(n9702), .B1(n9758), .B2(n9701), .ZN(n9712)
         );
  OAI21_X1 U10836 ( .B1(n9705), .B2(n9704), .A(n9703), .ZN(n9706) );
  AOI21_X1 U10837 ( .B1(n9707), .B2(n9706), .A(n9744), .ZN(n9708) );
  NOR3_X1 U10838 ( .A1(n9710), .A2(n9709), .A3(n9708), .ZN(n9711) );
  OAI211_X1 U10839 ( .C1(n9785), .C2(n9713), .A(n9712), .B(n9711), .ZN(
        P1_U3245) );
  INV_X1 U10840 ( .A(n9714), .ZN(n9720) );
  AND2_X1 U10841 ( .A1(n9716), .A2(n9715), .ZN(n9717) );
  OR3_X1 U10842 ( .A1(n9744), .A2(n9718), .A3(n9717), .ZN(n9719) );
  OAI211_X1 U10843 ( .C1(n9783), .C2(n4475), .A(n9720), .B(n9719), .ZN(n9721)
         );
  INV_X1 U10844 ( .A(n9721), .ZN(n9727) );
  OAI21_X1 U10845 ( .B1(n9724), .B2(n9723), .A(n9722), .ZN(n9725) );
  NAND2_X1 U10846 ( .A1(n9751), .A2(n9725), .ZN(n9726) );
  OAI211_X1 U10847 ( .C1(n10076), .C2(n9785), .A(n9727), .B(n9726), .ZN(
        P1_U3246) );
  OAI21_X1 U10848 ( .B1(n9730), .B2(n9729), .A(n9728), .ZN(n9736) );
  AOI211_X1 U10849 ( .C1(n9733), .C2(n9732), .A(n9731), .B(n9774), .ZN(n9734)
         );
  AOI211_X1 U10850 ( .C1(n9781), .C2(n9736), .A(n9735), .B(n9734), .ZN(n9741)
         );
  INV_X1 U10851 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n9738) );
  OAI22_X1 U10852 ( .A1(n9785), .A2(n9738), .B1(n9783), .B2(n9737), .ZN(n9739)
         );
  INV_X1 U10853 ( .A(n9739), .ZN(n9740) );
  NAND2_X1 U10854 ( .A1(n9741), .A2(n9740), .ZN(P1_U3247) );
  XNOR2_X1 U10855 ( .A(n9743), .B(n9742), .ZN(n9750) );
  AOI211_X1 U10856 ( .C1(n9747), .C2(n9746), .A(n9745), .B(n9744), .ZN(n9748)
         );
  AOI211_X1 U10857 ( .C1(n9751), .C2(n9750), .A(n9749), .B(n9748), .ZN(n9756)
         );
  INV_X1 U10858 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n9753) );
  OAI22_X1 U10859 ( .A1(n9785), .A2(n9753), .B1(n9783), .B2(n9752), .ZN(n9754)
         );
  INV_X1 U10860 ( .A(n9754), .ZN(n9755) );
  NAND2_X1 U10861 ( .A1(n9756), .A2(n9755), .ZN(P1_U3249) );
  AOI22_X1 U10862 ( .A1(n9759), .A2(P1_ADDR_REG_9__SCAN_IN), .B1(n9758), .B2(
        n9757), .ZN(n9770) );
  OAI21_X1 U10863 ( .B1(n9762), .B2(n9761), .A(n9760), .ZN(n9768) );
  AOI211_X1 U10864 ( .C1(n9765), .C2(n9764), .A(n9763), .B(n9774), .ZN(n9766)
         );
  AOI211_X1 U10865 ( .C1(n9781), .C2(n9768), .A(n9767), .B(n9766), .ZN(n9769)
         );
  NAND2_X1 U10866 ( .A1(n9770), .A2(n9769), .ZN(P1_U3250) );
  OAI21_X1 U10867 ( .B1(n9773), .B2(n9772), .A(n9771), .ZN(n9780) );
  AOI211_X1 U10868 ( .C1(n9777), .C2(n9776), .A(n9775), .B(n9774), .ZN(n9778)
         );
  AOI211_X1 U10869 ( .C1(n9781), .C2(n9780), .A(n9779), .B(n9778), .ZN(n9788)
         );
  INV_X1 U10870 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n9784) );
  OAI22_X1 U10871 ( .A1(n9785), .A2(n9784), .B1(n9783), .B2(n9782), .ZN(n9786)
         );
  INV_X1 U10872 ( .A(n9786), .ZN(n9787) );
  NAND2_X1 U10873 ( .A1(n9788), .A2(n9787), .ZN(P1_U3251) );
  XOR2_X1 U10874 ( .A(n9799), .B(n9789), .Z(n9807) );
  INV_X1 U10875 ( .A(n9807), .ZN(n9912) );
  INV_X1 U10876 ( .A(n9790), .ZN(n9792) );
  OAI21_X1 U10877 ( .B1(n9792), .B2(n9907), .A(n9791), .ZN(n9909) );
  INV_X1 U10878 ( .A(n9909), .ZN(n9793) );
  AOI22_X1 U10879 ( .A1(n9912), .A2(n9795), .B1(n9794), .B2(n9793), .ZN(n9816)
         );
  NAND2_X1 U10880 ( .A1(n9797), .A2(n9796), .ZN(n9798) );
  XOR2_X1 U10881 ( .A(n9799), .B(n9798), .Z(n9805) );
  OAI22_X1 U10882 ( .A1(n9803), .A2(n9802), .B1(n9801), .B2(n9800), .ZN(n9804)
         );
  AOI21_X1 U10883 ( .B1(n9805), .B2(n9823), .A(n9804), .ZN(n9806) );
  OAI21_X1 U10884 ( .B1(n9807), .B2(n9884), .A(n9806), .ZN(n9910) );
  NOR2_X1 U10885 ( .A1(n9808), .A2(n9907), .ZN(n9813) );
  OAI22_X1 U10886 ( .A1(n9814), .A2(n9811), .B1(n9810), .B2(n9809), .ZN(n9812)
         );
  AOI211_X1 U10887 ( .C1(n9910), .C2(n9814), .A(n9813), .B(n9812), .ZN(n9815)
         );
  NAND2_X1 U10888 ( .A1(n9816), .A2(n9815), .ZN(P1_U3282) );
  XNOR2_X1 U10889 ( .A(n9818), .B(n9817), .ZN(n9879) );
  AND2_X1 U10890 ( .A1(n9820), .A2(n9819), .ZN(n9822) );
  XNOR2_X1 U10891 ( .A(n9822), .B(n9821), .ZN(n9824) );
  NAND2_X1 U10892 ( .A1(n9824), .A2(n9823), .ZN(n9830) );
  AOI22_X1 U10893 ( .A1(n9828), .A2(n9827), .B1(n9826), .B2(n9825), .ZN(n9829)
         );
  NAND2_X1 U10894 ( .A1(n9830), .A2(n9829), .ZN(n9878) );
  NAND2_X1 U10895 ( .A1(n9831), .A2(n9835), .ZN(n9832) );
  NAND2_X1 U10896 ( .A1(n9832), .A2(n9881), .ZN(n9833) );
  OR2_X1 U10897 ( .A1(n9834), .A2(n9833), .ZN(n9875) );
  AOI22_X1 U10898 ( .A1(n9838), .A2(n9837), .B1(n9836), .B2(n9835), .ZN(n9839)
         );
  OAI21_X1 U10899 ( .B1(n9875), .B2(n9840), .A(n9839), .ZN(n9841) );
  AOI211_X1 U10900 ( .C1(n9879), .C2(n9842), .A(n9878), .B(n9841), .ZN(n9843)
         );
  AOI22_X1 U10901 ( .A1(n9844), .A2(n6083), .B1(n9843), .B2(n9814), .ZN(
        P1_U3286) );
  NAND2_X1 U10902 ( .A1(n9846), .A2(n9845), .ZN(n9847) );
  AND2_X1 U10903 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9847), .ZN(P1_U3292) );
  AND2_X1 U10904 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9847), .ZN(P1_U3293) );
  AND2_X1 U10905 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9847), .ZN(P1_U3294) );
  AND2_X1 U10906 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9847), .ZN(P1_U3295) );
  AND2_X1 U10907 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9847), .ZN(P1_U3296) );
  AND2_X1 U10908 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9847), .ZN(P1_U3297) );
  AND2_X1 U10909 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9847), .ZN(P1_U3298) );
  AND2_X1 U10910 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9847), .ZN(P1_U3299) );
  AND2_X1 U10911 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9847), .ZN(P1_U3300) );
  AND2_X1 U10912 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9847), .ZN(P1_U3301) );
  AND2_X1 U10913 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9847), .ZN(P1_U3302) );
  AND2_X1 U10914 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9847), .ZN(P1_U3303) );
  AND2_X1 U10915 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9847), .ZN(P1_U3304) );
  AND2_X1 U10916 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9847), .ZN(P1_U3305) );
  AND2_X1 U10917 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9847), .ZN(P1_U3306) );
  AND2_X1 U10918 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9847), .ZN(P1_U3307) );
  AND2_X1 U10919 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9847), .ZN(P1_U3308) );
  AND2_X1 U10920 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9847), .ZN(P1_U3309) );
  AND2_X1 U10921 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9847), .ZN(P1_U3310) );
  AND2_X1 U10922 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9847), .ZN(P1_U3311) );
  AND2_X1 U10923 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9847), .ZN(P1_U3312) );
  AND2_X1 U10924 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9847), .ZN(P1_U3313) );
  AND2_X1 U10925 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9847), .ZN(P1_U3314) );
  AND2_X1 U10926 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9847), .ZN(P1_U3315) );
  AND2_X1 U10927 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9847), .ZN(P1_U3316) );
  AND2_X1 U10928 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9847), .ZN(P1_U3317) );
  AND2_X1 U10929 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9847), .ZN(P1_U3318) );
  AND2_X1 U10930 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n9847), .ZN(P1_U3319) );
  AND2_X1 U10931 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9847), .ZN(P1_U3320) );
  AND2_X1 U10932 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9847), .ZN(P1_U3321) );
  INV_X1 U10933 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n9849) );
  AOI21_X1 U10934 ( .B1(n9850), .B2(n9849), .A(n9848), .ZN(P1_U3440) );
  INV_X1 U10935 ( .A(n9851), .ZN(n9852) );
  OAI211_X1 U10936 ( .C1(n9854), .C2(n9897), .A(n9853), .B(n9852), .ZN(n9855)
         );
  NOR2_X1 U10937 ( .A1(n9856), .A2(n9855), .ZN(n9917) );
  INV_X1 U10938 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9857) );
  AOI22_X1 U10939 ( .A1(n9916), .A2(n9917), .B1(n9857), .B2(n9914), .ZN(
        P1_U3457) );
  OAI22_X1 U10940 ( .A1(n9858), .A2(n9908), .B1(n6380), .B2(n9906), .ZN(n9860)
         );
  AOI211_X1 U10941 ( .C1(n9913), .C2(n9861), .A(n9860), .B(n9859), .ZN(n9918)
         );
  INV_X1 U10942 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9862) );
  AOI22_X1 U10943 ( .A1(n9916), .A2(n9918), .B1(n9862), .B2(n9914), .ZN(
        P1_U3460) );
  OAI22_X1 U10944 ( .A1(n9864), .A2(n9908), .B1(n9863), .B2(n9906), .ZN(n9866)
         );
  AOI211_X1 U10945 ( .C1(n9913), .C2(n9867), .A(n9866), .B(n9865), .ZN(n9920)
         );
  INV_X1 U10946 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n9868) );
  AOI22_X1 U10947 ( .A1(n9916), .A2(n9920), .B1(n9868), .B2(n9914), .ZN(
        P1_U3463) );
  OAI22_X1 U10948 ( .A1(n9870), .A2(n9908), .B1(n9869), .B2(n9906), .ZN(n9872)
         );
  AOI211_X1 U10949 ( .C1(n9913), .C2(n9873), .A(n9872), .B(n9871), .ZN(n9921)
         );
  INV_X1 U10950 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n9874) );
  AOI22_X1 U10951 ( .A1(n9916), .A2(n9921), .B1(n9874), .B2(n9914), .ZN(
        P1_U3466) );
  OAI21_X1 U10952 ( .B1(n9876), .B2(n9906), .A(n9875), .ZN(n9877) );
  AOI211_X1 U10953 ( .C1(n9879), .C2(n9895), .A(n9878), .B(n9877), .ZN(n9922)
         );
  AOI22_X1 U10954 ( .A1(n9916), .A2(n9922), .B1(n6080), .B2(n9914), .ZN(
        P1_U3469) );
  AOI21_X1 U10955 ( .B1(n9882), .B2(n9881), .A(n9880), .ZN(n9883) );
  OAI21_X1 U10956 ( .B1(n9885), .B2(n9884), .A(n9883), .ZN(n9886) );
  AOI211_X1 U10957 ( .C1(n9913), .C2(n9888), .A(n9887), .B(n9886), .ZN(n9923)
         );
  INV_X1 U10958 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9889) );
  AOI22_X1 U10959 ( .A1(n9916), .A2(n9923), .B1(n9889), .B2(n9914), .ZN(
        P1_U3472) );
  OAI211_X1 U10960 ( .C1(n9892), .C2(n9906), .A(n9891), .B(n9890), .ZN(n9893)
         );
  AOI21_X1 U10961 ( .B1(n9895), .B2(n9894), .A(n9893), .ZN(n9924) );
  INV_X1 U10962 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9896) );
  AOI22_X1 U10963 ( .A1(n9916), .A2(n9924), .B1(n9896), .B2(n9914), .ZN(
        P1_U3475) );
  NOR3_X1 U10964 ( .A1(n9899), .A2(n9898), .A3(n9897), .ZN(n9904) );
  NOR2_X1 U10965 ( .A1(n9900), .A2(n9908), .ZN(n9902) );
  NOR4_X1 U10966 ( .A1(n9904), .A2(n9903), .A3(n9902), .A4(n9901), .ZN(n9925)
         );
  INV_X1 U10967 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n9905) );
  AOI22_X1 U10968 ( .A1(n9916), .A2(n9925), .B1(n9905), .B2(n9914), .ZN(
        P1_U3478) );
  OAI22_X1 U10969 ( .A1(n9909), .A2(n9908), .B1(n9907), .B2(n9906), .ZN(n9911)
         );
  AOI211_X1 U10970 ( .C1(n9913), .C2(n9912), .A(n9911), .B(n9910), .ZN(n9927)
         );
  INV_X1 U10971 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9915) );
  AOI22_X1 U10972 ( .A1(n9916), .A2(n9927), .B1(n9915), .B2(n9914), .ZN(
        P1_U3481) );
  AOI22_X1 U10973 ( .A1(n9928), .A2(n9917), .B1(n5878), .B2(n9926), .ZN(
        P1_U3524) );
  AOI22_X1 U10974 ( .A1(n9928), .A2(n9918), .B1(n5932), .B2(n9926), .ZN(
        P1_U3525) );
  AOI22_X1 U10975 ( .A1(n9928), .A2(n9920), .B1(n9919), .B2(n9926), .ZN(
        P1_U3526) );
  AOI22_X1 U10976 ( .A1(n9928), .A2(n9921), .B1(n6061), .B2(n9926), .ZN(
        P1_U3527) );
  AOI22_X1 U10977 ( .A1(n9928), .A2(n9922), .B1(n6082), .B2(n9926), .ZN(
        P1_U3528) );
  AOI22_X1 U10978 ( .A1(n9928), .A2(n9923), .B1(n6320), .B2(n9926), .ZN(
        P1_U3529) );
  AOI22_X1 U10979 ( .A1(n9928), .A2(n9924), .B1(n6340), .B2(n9926), .ZN(
        P1_U3530) );
  AOI22_X1 U10980 ( .A1(n9928), .A2(n9925), .B1(n6360), .B2(n9926), .ZN(
        P1_U3531) );
  AOI22_X1 U10981 ( .A1(n9928), .A2(n9927), .B1(n6589), .B2(n9926), .ZN(
        P1_U3532) );
  AOI22_X1 U10982 ( .A1(n9929), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n9930), .ZN(n9939) );
  NAND2_X1 U10983 ( .A1(n9930), .A2(n10020), .ZN(n9931) );
  OAI211_X1 U10984 ( .C1(P2_REG2_REG_0__SCAN_IN), .C2(n9933), .A(n9932), .B(
        n9931), .ZN(n9934) );
  INV_X1 U10985 ( .A(n9934), .ZN(n9937) );
  AOI22_X1 U10986 ( .A1(n9935), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n9936) );
  OAI221_X1 U10987 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n9939), .C1(n9938), .C2(
        n9937), .A(n9936), .ZN(P2_U3245) );
  INV_X1 U10988 ( .A(n9940), .ZN(n9951) );
  INV_X1 U10989 ( .A(n9941), .ZN(n9947) );
  AOI22_X1 U10990 ( .A1(n9944), .A2(n9943), .B1(n9942), .B2(n5264), .ZN(n9945)
         );
  OAI21_X1 U10991 ( .B1(n9947), .B2(n9946), .A(n9945), .ZN(n9950) );
  INV_X1 U10992 ( .A(n9948), .ZN(n9949) );
  AOI211_X1 U10993 ( .C1(n9952), .C2(n9951), .A(n9950), .B(n9949), .ZN(n9954)
         );
  AOI22_X1 U10994 ( .A1(n8368), .A2(n5709), .B1(n9954), .B2(n9953), .ZN(
        P2_U3291) );
  AND2_X1 U10995 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n9959), .ZN(P2_U3297) );
  AND2_X1 U10996 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n9959), .ZN(P2_U3298) );
  AND2_X1 U10997 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n9959), .ZN(P2_U3299) );
  AND2_X1 U10998 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n9959), .ZN(P2_U3300) );
  AND2_X1 U10999 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n9959), .ZN(P2_U3301) );
  AND2_X1 U11000 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n9959), .ZN(P2_U3302) );
  AND2_X1 U11001 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n9959), .ZN(P2_U3303) );
  AND2_X1 U11002 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n9959), .ZN(P2_U3304) );
  AND2_X1 U11003 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n9959), .ZN(P2_U3305) );
  AND2_X1 U11004 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n9959), .ZN(P2_U3306) );
  AND2_X1 U11005 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n9959), .ZN(P2_U3307) );
  AND2_X1 U11006 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n9959), .ZN(P2_U3308) );
  AND2_X1 U11007 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n9959), .ZN(P2_U3309) );
  AND2_X1 U11008 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n9959), .ZN(P2_U3310) );
  AND2_X1 U11009 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n9959), .ZN(P2_U3311) );
  AND2_X1 U11010 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n9959), .ZN(P2_U3312) );
  AND2_X1 U11011 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n9959), .ZN(P2_U3313) );
  AND2_X1 U11012 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n9959), .ZN(P2_U3314) );
  AND2_X1 U11013 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n9959), .ZN(P2_U3315) );
  AND2_X1 U11014 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n9959), .ZN(P2_U3316) );
  AND2_X1 U11015 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n9959), .ZN(P2_U3317) );
  AND2_X1 U11016 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n9959), .ZN(P2_U3318) );
  AND2_X1 U11017 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n9959), .ZN(P2_U3319) );
  AND2_X1 U11018 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n9959), .ZN(P2_U3320) );
  AND2_X1 U11019 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n9959), .ZN(P2_U3321) );
  AND2_X1 U11020 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n9959), .ZN(P2_U3322) );
  AND2_X1 U11021 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n9959), .ZN(P2_U3323) );
  AND2_X1 U11022 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n9959), .ZN(P2_U3324) );
  AND2_X1 U11023 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n9959), .ZN(P2_U3325) );
  AND2_X1 U11024 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n9959), .ZN(P2_U3326) );
  AOI22_X1 U11025 ( .A1(n9958), .A2(n9961), .B1(n9957), .B2(n9959), .ZN(
        P2_U3437) );
  AOI22_X1 U11026 ( .A1(n9962), .A2(n9961), .B1(n9960), .B2(n9959), .ZN(
        P2_U3438) );
  AOI22_X1 U11027 ( .A1(n9965), .A2(n10015), .B1(n9964), .B2(n9963), .ZN(n9966) );
  AND2_X1 U11028 ( .A1(n9967), .A2(n9966), .ZN(n10021) );
  INV_X1 U11029 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n9968) );
  AOI22_X1 U11030 ( .A1(n10019), .A2(n10021), .B1(n9968), .B2(n10017), .ZN(
        P2_U3451) );
  INV_X1 U11031 ( .A(n9969), .ZN(n9970) );
  OAI22_X1 U11032 ( .A1(n9970), .A2(n10010), .B1(n5234), .B2(n10008), .ZN(
        n9972) );
  AOI211_X1 U11033 ( .C1(n10015), .C2(n9973), .A(n9972), .B(n9971), .ZN(n10023) );
  INV_X1 U11034 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n9974) );
  AOI22_X1 U11035 ( .A1(n10019), .A2(n10023), .B1(n9974), .B2(n10017), .ZN(
        P2_U3454) );
  OAI22_X1 U11036 ( .A1(n9976), .A2(n10010), .B1(n9975), .B2(n10008), .ZN(
        n9978) );
  AOI211_X1 U11037 ( .C1(n9979), .C2(n10015), .A(n9978), .B(n9977), .ZN(n10024) );
  INV_X1 U11038 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n9980) );
  AOI22_X1 U11039 ( .A1(n10019), .A2(n10024), .B1(n9980), .B2(n10017), .ZN(
        P2_U3457) );
  OAI22_X1 U11040 ( .A1(n9982), .A2(n10010), .B1(n9981), .B2(n10008), .ZN(
        n9984) );
  AOI211_X1 U11041 ( .C1(n10015), .C2(n9985), .A(n9984), .B(n9983), .ZN(n10026) );
  INV_X1 U11042 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n9986) );
  AOI22_X1 U11043 ( .A1(n10019), .A2(n10026), .B1(n9986), .B2(n10017), .ZN(
        P2_U3463) );
  INV_X1 U11044 ( .A(n9987), .ZN(n9993) );
  OAI22_X1 U11045 ( .A1(n9989), .A2(n10010), .B1(n9988), .B2(n10008), .ZN(
        n9992) );
  INV_X1 U11046 ( .A(n9990), .ZN(n9991) );
  AOI211_X1 U11047 ( .C1(n10015), .C2(n9993), .A(n9992), .B(n9991), .ZN(n10027) );
  INV_X1 U11048 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n9994) );
  AOI22_X1 U11049 ( .A1(n10019), .A2(n10027), .B1(n9994), .B2(n10017), .ZN(
        P2_U3469) );
  OAI22_X1 U11050 ( .A1(n9996), .A2(n10010), .B1(n9995), .B2(n10008), .ZN(
        n9998) );
  AOI211_X1 U11051 ( .C1(n10006), .C2(n9999), .A(n9998), .B(n9997), .ZN(n10028) );
  INV_X1 U11052 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10000) );
  AOI22_X1 U11053 ( .A1(n10019), .A2(n10028), .B1(n10000), .B2(n10017), .ZN(
        P2_U3475) );
  OAI22_X1 U11054 ( .A1(n10002), .A2(n10010), .B1(n10001), .B2(n10008), .ZN(
        n10004) );
  AOI211_X1 U11055 ( .C1(n10006), .C2(n10005), .A(n10004), .B(n10003), .ZN(
        n10029) );
  INV_X1 U11056 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10007) );
  AOI22_X1 U11057 ( .A1(n10019), .A2(n10029), .B1(n10007), .B2(n10017), .ZN(
        P2_U3481) );
  OAI22_X1 U11058 ( .A1(n10011), .A2(n10010), .B1(n10009), .B2(n10008), .ZN(
        n10014) );
  INV_X1 U11059 ( .A(n10012), .ZN(n10013) );
  AOI211_X1 U11060 ( .C1(n10016), .C2(n10015), .A(n10014), .B(n10013), .ZN(
        n10032) );
  INV_X1 U11061 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10018) );
  AOI22_X1 U11062 ( .A1(n10019), .A2(n10032), .B1(n10018), .B2(n10017), .ZN(
        P2_U3487) );
  AOI22_X1 U11063 ( .A1(n10033), .A2(n10021), .B1(n10020), .B2(n10030), .ZN(
        P2_U3520) );
  INV_X1 U11064 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10022) );
  AOI22_X1 U11065 ( .A1(n10033), .A2(n10023), .B1(n10022), .B2(n10030), .ZN(
        P2_U3521) );
  AOI22_X1 U11066 ( .A1(n10033), .A2(n10024), .B1(n5680), .B2(n10030), .ZN(
        P2_U3522) );
  INV_X1 U11067 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10025) );
  AOI22_X1 U11068 ( .A1(n10033), .A2(n10026), .B1(n10025), .B2(n10030), .ZN(
        P2_U3524) );
  AOI22_X1 U11069 ( .A1(n10033), .A2(n10027), .B1(n5704), .B2(n10030), .ZN(
        P2_U3526) );
  AOI22_X1 U11070 ( .A1(n10033), .A2(n10028), .B1(n5776), .B2(n10030), .ZN(
        P2_U3528) );
  AOI22_X1 U11071 ( .A1(n10033), .A2(n10029), .B1(n5780), .B2(n10030), .ZN(
        P2_U3530) );
  AOI22_X1 U11072 ( .A1(n10033), .A2(n10032), .B1(n10031), .B2(n10030), .ZN(
        P2_U3532) );
  INV_X1 U11073 ( .A(n10034), .ZN(n10035) );
  NAND2_X1 U11074 ( .A1(n10036), .A2(n10035), .ZN(n10037) );
  XNOR2_X1 U11075 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n10037), .ZN(ADD_1071_U5)
         );
  XOR2_X1 U11076 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  OAI21_X1 U11077 ( .B1(n10040), .B2(n10039), .A(n10038), .ZN(ADD_1071_U56) );
  OAI21_X1 U11078 ( .B1(n10043), .B2(n10042), .A(n10041), .ZN(ADD_1071_U57) );
  OAI21_X1 U11079 ( .B1(n10046), .B2(n10045), .A(n10044), .ZN(ADD_1071_U58) );
  OAI21_X1 U11080 ( .B1(n10049), .B2(n10048), .A(n10047), .ZN(ADD_1071_U59) );
  OAI21_X1 U11081 ( .B1(n10052), .B2(n10051), .A(n10050), .ZN(ADD_1071_U60) );
  OAI21_X1 U11082 ( .B1(n10055), .B2(n10054), .A(n10053), .ZN(ADD_1071_U61) );
  AOI21_X1 U11083 ( .B1(n10058), .B2(n10057), .A(n10056), .ZN(ADD_1071_U62) );
  AOI21_X1 U11084 ( .B1(n10061), .B2(n10060), .A(n10059), .ZN(ADD_1071_U63) );
  AOI21_X1 U11085 ( .B1(n10064), .B2(n10063), .A(n10062), .ZN(ADD_1071_U47) );
  XOR2_X1 U11086 ( .A(n10066), .B(n10065), .Z(ADD_1071_U54) );
  XOR2_X1 U11087 ( .A(n10067), .B(P2_ADDR_REG_8__SCAN_IN), .Z(ADD_1071_U48) );
  OAI21_X1 U11088 ( .B1(n10070), .B2(n10069), .A(n10068), .ZN(n10071) );
  XNOR2_X1 U11089 ( .A(n10071), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  XOR2_X1 U11090 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(n10072), .Z(ADD_1071_U49) );
  XOR2_X1 U11091 ( .A(P2_ADDR_REG_6__SCAN_IN), .B(n10073), .Z(ADD_1071_U50) );
  AOI21_X1 U11092 ( .B1(n10075), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n10074), .ZN(
        n10077) );
  XNOR2_X1 U11093 ( .A(n10077), .B(n10076), .ZN(ADD_1071_U51) );
  XOR2_X1 U11094 ( .A(n10079), .B(n10078), .Z(ADD_1071_U53) );
  XNOR2_X1 U11095 ( .A(n10081), .B(n10080), .ZN(ADD_1071_U52) );
  INV_X1 U4817 ( .A(n7598), .ZN(n5931) );
endmodule

