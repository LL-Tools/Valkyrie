

module b22_C_2inp_gates_syn ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, SUB_1596_U4, 
        SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, 
        SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, 
        SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, 
        SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, U29, U28, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, 
        P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, 
        P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, P1_U3515, 
        P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, 
        P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, 
        P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, 
        P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, 
        P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, 
        P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, P1_U3557, 
        P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, P1_U3561, 
        P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, 
        P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, 
        P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, 
        P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, P1_U3589, 
        P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U4016, 
        P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, 
        P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, 
        P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, 
        P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, 
        P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, P2_U3295, 
        P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, 
        P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, 
        P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, 
        P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, 
        P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, P2_U3445, 
        P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, 
        P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3486, 
        P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, P2_U3493, 
        P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, 
        P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, 
        P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, 
        P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, 
        P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, 
        P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, 
        P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, P2_U3532, 
        P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, 
        P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, 
        P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, P2_U3553, 
        P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, 
        P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, P2_U3210, 
        P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, 
        P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, 
        P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, 
        P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, P2_U3947, 
        P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, P3_U3289, 
        P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, P3_U3282, 
        P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, P3_U3275, 
        P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, P3_U3268, 
        P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, P3_U3263, 
        P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, P3_U3256, 
        P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, P3_U3249, 
        P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, P3_U3242, 
        P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, P3_U3235, 
        P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, P3_U3405, 
        P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, P3_U3426, 
        P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, P3_U3446, 
        P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, P3_U3453, 
        P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, P3_U3460, 
        P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, P3_U3467, 
        P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, P3_U3474, 
        P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, P3_U3481, 
        P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, P3_U3488, 
        P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, P3_U3229, 
        P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, P3_U3222, 
        P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, P3_U3215, 
        P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, P3_U3208, 
        P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, P3_U3201, 
        P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, P3_U3194, 
        P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, P3_U3187, 
        P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, P3_U3492, 
        P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, P3_U3499, 
        P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, P3_U3506, 
        P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, P3_U3513, 
        P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, P3_U3520, 
        P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, P3_U3178, 
        P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, P3_U3171, 
        P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, P3_U3164, 
        P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, P3_U3157, 
        P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, P3_U3897, 
        keyinput127, keyinput126, keyinput125, keyinput124, keyinput123, 
        keyinput122, keyinput121, keyinput120, keyinput119, keyinput118, 
        keyinput117, keyinput116, keyinput115, keyinput114, keyinput113, 
        keyinput112, keyinput111, keyinput110, keyinput109, keyinput108, 
        keyinput107, keyinput106, keyinput105, keyinput104, keyinput103, 
        keyinput102, keyinput101, keyinput100, keyinput99, keyinput98, 
        keyinput97, keyinput96, keyinput95, keyinput94, keyinput93, keyinput92, 
        keyinput91, keyinput90, keyinput89, keyinput88, keyinput87, keyinput86, 
        keyinput85, keyinput84, keyinput83, keyinput82, keyinput81, keyinput80, 
        keyinput79, keyinput78, keyinput77, keyinput76, keyinput75, keyinput74, 
        keyinput73, keyinput72, keyinput71, keyinput70, keyinput69, keyinput68, 
        keyinput67, keyinput66, keyinput65, keyinput64, keyinput63, keyinput62, 
        keyinput61, keyinput60, keyinput59, keyinput58, keyinput57, keyinput56, 
        keyinput55, keyinput54, keyinput53, keyinput52, keyinput51, keyinput50, 
        keyinput49, keyinput48, keyinput47, keyinput46, keyinput45, keyinput44, 
        keyinput43, keyinput42, keyinput41, keyinput40, keyinput39, keyinput38, 
        keyinput37, keyinput36, keyinput35, keyinput34, keyinput33, keyinput32, 
        keyinput31, keyinput30, keyinput29, keyinput28, keyinput27, keyinput26, 
        keyinput25, keyinput24, keyinput23, keyinput22, keyinput21, keyinput20, 
        keyinput19, keyinput18, keyinput17, keyinput16, keyinput15, keyinput14, 
        keyinput13, keyinput12, keyinput11, keyinput10, keyinput9, keyinput8, 
        keyinput7, keyinput6, keyinput5, keyinput4, keyinput3, keyinput2, 
        keyinput1, keyinput0 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput127,
         keyinput126, keyinput125, keyinput124, keyinput123, keyinput122,
         keyinput121, keyinput120, keyinput119, keyinput118, keyinput117,
         keyinput116, keyinput115, keyinput114, keyinput113, keyinput112,
         keyinput111, keyinput110, keyinput109, keyinput108, keyinput107,
         keyinput106, keyinput105, keyinput104, keyinput103, keyinput102,
         keyinput101, keyinput100, keyinput99, keyinput98, keyinput97,
         keyinput96, keyinput95, keyinput94, keyinput93, keyinput92,
         keyinput91, keyinput90, keyinput89, keyinput88, keyinput87,
         keyinput86, keyinput85, keyinput84, keyinput83, keyinput82,
         keyinput81, keyinput80, keyinput79, keyinput78, keyinput77,
         keyinput76, keyinput75, keyinput74, keyinput73, keyinput72,
         keyinput71, keyinput70, keyinput69, keyinput68, keyinput67,
         keyinput66, keyinput65, keyinput64, keyinput63, keyinput62,
         keyinput61, keyinput60, keyinput59, keyinput58, keyinput57,
         keyinput56, keyinput55, keyinput54, keyinput53, keyinput52,
         keyinput51, keyinput50, keyinput49, keyinput48, keyinput47,
         keyinput46, keyinput45, keyinput44, keyinput43, keyinput42,
         keyinput41, keyinput40, keyinput39, keyinput38, keyinput37,
         keyinput36, keyinput35, keyinput34, keyinput33, keyinput32,
         keyinput31, keyinput30, keyinput29, keyinput28, keyinput27,
         keyinput26, keyinput25, keyinput24, keyinput23, keyinput22,
         keyinput21, keyinput20, keyinput19, keyinput18, keyinput17,
         keyinput16, keyinput15, keyinput14, keyinput13, keyinput12,
         keyinput11, keyinput10, keyinput9, keyinput8, keyinput7, keyinput6,
         keyinput5, keyinput4, keyinput3, keyinput2, keyinput1, keyinput0;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554,
         n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564,
         n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574,
         n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584,
         n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594,
         n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
         n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614,
         n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624,
         n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634,
         n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644,
         n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654,
         n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664,
         n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674,
         n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684,
         n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694,
         n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704,
         n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714,
         n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724,
         n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734,
         n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744,
         n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754,
         n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764,
         n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774,
         n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784,
         n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794,
         n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804,
         n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814,
         n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824,
         n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834,
         n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844,
         n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854,
         n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864,
         n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874,
         n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884,
         n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894,
         n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904,
         n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914,
         n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924,
         n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934,
         n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944,
         n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954,
         n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964,
         n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974,
         n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984,
         n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994,
         n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004,
         n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014,
         n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024,
         n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034,
         n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044,
         n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054,
         n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064,
         n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074,
         n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084,
         n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094,
         n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104,
         n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114,
         n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124,
         n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134,
         n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144,
         n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154,
         n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164,
         n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174,
         n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184,
         n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194,
         n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204,
         n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214,
         n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224,
         n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234,
         n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244,
         n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254,
         n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264,
         n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274,
         n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284,
         n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294,
         n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304,
         n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314,
         n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324,
         n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334,
         n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344,
         n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354,
         n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364,
         n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374,
         n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384,
         n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394,
         n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404,
         n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414,
         n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424,
         n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434,
         n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444,
         n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454,
         n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464,
         n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474,
         n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484,
         n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494,
         n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504,
         n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514,
         n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524,
         n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534,
         n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544,
         n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554,
         n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564,
         n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574,
         n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584,
         n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594,
         n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604,
         n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614,
         n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624,
         n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634,
         n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644,
         n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654,
         n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664,
         n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674,
         n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684,
         n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694,
         n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704,
         n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714,
         n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724,
         n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734,
         n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744,
         n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754,
         n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764,
         n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774,
         n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784,
         n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794,
         n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804,
         n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814,
         n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824,
         n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834,
         n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844,
         n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854,
         n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864,
         n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874,
         n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884,
         n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894,
         n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904,
         n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914,
         n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924,
         n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934,
         n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944,
         n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954,
         n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964,
         n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974,
         n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984,
         n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994,
         n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004,
         n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014,
         n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024,
         n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034,
         n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044,
         n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054,
         n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064,
         n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074,
         n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084,
         n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094,
         n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104,
         n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114,
         n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124,
         n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134,
         n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144,
         n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154,
         n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164,
         n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174,
         n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184,
         n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194,
         n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204,
         n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214,
         n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224,
         n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234,
         n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244,
         n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254,
         n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264,
         n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274,
         n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284,
         n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294,
         n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304,
         n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314,
         n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324,
         n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334,
         n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344,
         n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354,
         n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364,
         n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374,
         n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384,
         n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394,
         n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404,
         n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414,
         n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424,
         n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434,
         n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444,
         n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454,
         n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464,
         n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474,
         n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484,
         n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494,
         n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504,
         n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514,
         n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524,
         n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534,
         n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544,
         n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554,
         n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564,
         n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574,
         n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584,
         n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594,
         n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604,
         n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614,
         n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624,
         n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634,
         n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644,
         n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654,
         n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664,
         n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674,
         n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684,
         n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694,
         n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704,
         n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714,
         n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724,
         n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734,
         n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744,
         n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754,
         n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764,
         n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774,
         n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784,
         n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794,
         n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804,
         n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814,
         n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824,
         n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834,
         n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844,
         n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854,
         n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864,
         n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874,
         n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884,
         n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894,
         n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904,
         n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914,
         n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924,
         n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934,
         n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944,
         n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954,
         n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964,
         n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974,
         n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984,
         n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994,
         n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004,
         n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014,
         n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024,
         n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034,
         n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044,
         n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054,
         n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064,
         n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074,
         n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084,
         n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094,
         n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104,
         n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114,
         n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124,
         n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134,
         n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144,
         n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154,
         n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164,
         n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174,
         n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184,
         n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194,
         n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204,
         n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214,
         n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224,
         n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234,
         n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244,
         n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254,
         n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264,
         n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274,
         n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284,
         n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294,
         n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304,
         n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314,
         n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324,
         n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334,
         n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344,
         n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354,
         n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364,
         n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374,
         n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384,
         n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394,
         n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404,
         n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414,
         n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424,
         n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434,
         n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444,
         n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454,
         n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464,
         n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474,
         n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484,
         n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494,
         n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504,
         n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514,
         n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524,
         n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534,
         n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544,
         n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554,
         n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564,
         n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574,
         n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584,
         n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594,
         n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604,
         n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614,
         n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624,
         n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634,
         n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644,
         n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654,
         n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664,
         n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674,
         n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684,
         n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694,
         n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704,
         n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714,
         n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724,
         n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734,
         n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744,
         n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754,
         n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764,
         n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774,
         n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784,
         n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794,
         n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804,
         n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814,
         n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824,
         n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834,
         n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844,
         n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854,
         n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864,
         n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874,
         n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884,
         n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894,
         n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904,
         n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914,
         n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924,
         n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934,
         n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944,
         n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954,
         n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964,
         n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974,
         n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984,
         n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994,
         n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003,
         n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011,
         n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019,
         n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027,
         n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035,
         n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043,
         n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051,
         n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059,
         n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067,
         n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075,
         n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083,
         n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091,
         n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099,
         n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107,
         n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115,
         n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123,
         n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131,
         n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139,
         n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147,
         n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155,
         n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163,
         n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171,
         n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179,
         n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187,
         n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195,
         n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203,
         n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211,
         n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219,
         n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227,
         n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235,
         n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243,
         n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251,
         n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259,
         n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267,
         n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275,
         n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283,
         n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291,
         n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299,
         n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307,
         n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315,
         n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323,
         n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331,
         n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339,
         n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347,
         n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355,
         n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363,
         n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371,
         n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379,
         n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387,
         n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395,
         n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403,
         n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411,
         n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419,
         n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427,
         n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435,
         n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443,
         n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451,
         n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459,
         n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467,
         n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475,
         n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483,
         n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491,
         n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499,
         n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507,
         n10508, n10509, n10510, n10511, n10512, n10513, n10514, n10515,
         n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523,
         n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531,
         n10532, n10533, n10534, n10535, n10536, n10537, n10538, n10539,
         n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547,
         n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555,
         n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563,
         n10564, n10565, n10566, n10567, n10568, n10569, n10570, n10571,
         n10572, n10573, n10574, n10575, n10576, n10577, n10578, n10579,
         n10580, n10581, n10582, n10583, n10584, n10585, n10586, n10587,
         n10588, n10589, n10590, n10591, n10592, n10593, n10594, n10595,
         n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603,
         n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10611,
         n10612, n10613, n10614, n10615, n10616, n10617, n10618, n10619,
         n10620, n10621, n10622, n10623, n10624, n10625, n10626, n10627,
         n10628, n10629, n10630, n10631, n10632, n10633, n10634, n10635,
         n10636, n10637, n10638, n10639, n10640, n10641, n10642, n10643,
         n10644, n10645, n10646, n10647, n10648, n10649, n10650, n10651,
         n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659,
         n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667,
         n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675,
         n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10683,
         n10684, n10685, n10686, n10687, n10688, n10689, n10690, n10691,
         n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699,
         n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707,
         n10708, n10709, n10710, n10711, n10712, n10713, n10714, n10715,
         n10716, n10717, n10718, n10719, n10720, n10721, n10722, n10723,
         n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731,
         n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739,
         n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747,
         n10748, n10749, n10750, n10751, n10752, n10753, n10754, n10755,
         n10756, n10757, n10758, n10759, n10760, n10761, n10762, n10763,
         n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771,
         n10772, n10773, n10774, n10775, n10776, n10777, n10778, n10779,
         n10780, n10781, n10782, n10783, n10784, n10785, n10786, n10787,
         n10788, n10789, n10790, n10791, n10792, n10793, n10794, n10795,
         n10796, n10797, n10798, n10799, n10800, n10801, n10802, n10803,
         n10804, n10805, n10806, n10807, n10808, n10809, n10810, n10811,
         n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819,
         n10820, n10821, n10822, n10823, n10824, n10825, n10826, n10827,
         n10828, n10829, n10830, n10831, n10832, n10833, n10834, n10835,
         n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843,
         n10844, n10845, n10846, n10847, n10848, n10849, n10850, n10851,
         n10852, n10853, n10854, n10855, n10856, n10857, n10858, n10859,
         n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867,
         n10868, n10869, n10870, n10871, n10872, n10873, n10874, n10875,
         n10876, n10877, n10878, n10879, n10880, n10881, n10882, n10883,
         n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891,
         n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899,
         n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907,
         n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915,
         n10916, n10917, n10918, n10919, n10920, n10921, n10922, n10923,
         n10924, n10925, n10926, n10927, n10928, n10929, n10930, n10931,
         n10932, n10933, n10934, n10935, n10936, n10937, n10938, n10939,
         n10940, n10941, n10942, n10943, n10944, n10945, n10946, n10947,
         n10948, n10949, n10950, n10951, n10952, n10953, n10954, n10955,
         n10956, n10957, n10958, n10959, n10960, n10961, n10962, n10963,
         n10964, n10965, n10966, n10967, n10968, n10969, n10970, n10971,
         n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979,
         n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987,
         n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995,
         n10996, n10997, n10998, n10999, n11000, n11001, n11002, n11003,
         n11004, n11005, n11006, n11007, n11008, n11009, n11010, n11011,
         n11012, n11013, n11014, n11015, n11016, n11017, n11018, n11019,
         n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027,
         n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035,
         n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11043,
         n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051,
         n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059,
         n11060, n11061, n11062, n11063, n11064, n11065, n11066, n11067,
         n11068, n11069, n11070, n11071, n11072, n11073, n11074, n11075,
         n11076, n11077, n11078, n11079, n11080, n11081, n11082, n11083,
         n11084, n11085, n11086, n11087, n11088, n11089, n11090, n11091,
         n11092, n11093, n11094, n11095, n11096, n11097, n11098, n11099,
         n11100, n11101, n11102, n11103, n11104, n11105, n11106, n11107,
         n11108, n11109, n11110, n11111, n11112, n11113, n11114, n11115,
         n11116, n11117, n11118, n11119, n11120, n11121, n11122, n11123,
         n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131,
         n11132, n11133, n11134, n11135, n11136, n11137, n11138, n11139,
         n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147,
         n11148, n11149, n11150, n11151, n11152, n11153, n11154, n11155,
         n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163,
         n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171,
         n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179,
         n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187,
         n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195,
         n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203,
         n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211,
         n11212, n11213, n11214, n11215, n11216, n11217, n11218, n11219,
         n11220, n11221, n11222, n11223, n11224, n11225, n11226, n11227,
         n11228, n11229, n11230, n11231, n11232, n11233, n11234, n11235,
         n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243,
         n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251,
         n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259,
         n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267,
         n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275,
         n11276, n11277, n11278, n11279, n11280, n11281, n11282, n11283,
         n11284, n11285, n11286, n11287, n11288, n11289, n11290, n11291,
         n11292, n11293, n11294, n11295, n11296, n11297, n11298, n11299,
         n11300, n11301, n11302, n11303, n11304, n11305, n11306, n11307,
         n11308, n11309, n11310, n11311, n11312, n11313, n11314, n11315,
         n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323,
         n11324, n11325, n11326, n11327, n11328, n11329, n11330, n11331,
         n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339,
         n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347,
         n11348, n11349, n11350, n11351, n11352, n11353, n11354, n11355,
         n11356, n11357, n11358, n11359, n11360, n11361, n11362, n11363,
         n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371,
         n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379,
         n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387,
         n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395,
         n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403,
         n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411,
         n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419,
         n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427,
         n11428, n11429, n11430, n11431, n11432, n11433, n11434, n11435,
         n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443,
         n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451,
         n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459,
         n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467,
         n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475,
         n11476, n11477, n11478, n11479, n11480, n11481, n11482, n11483,
         n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491,
         n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499,
         n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507,
         n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515,
         n11516, n11517, n11518, n11519, n11520, n11521, n11522, n11523,
         n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531,
         n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539,
         n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547,
         n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555,
         n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563,
         n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571,
         n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11579,
         n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587,
         n11588, n11589, n11590, n11591, n11592, n11593, n11594, n11595,
         n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603,
         n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611,
         n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619,
         n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627,
         n11628, n11629, n11630, n11631, n11632, n11633, n11634, n11635,
         n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643,
         n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651,
         n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659,
         n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667,
         n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675,
         n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683,
         n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691,
         n11692, n11693, n11694, n11695, n11696, n11697, n11698, n11699,
         n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707,
         n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715,
         n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723,
         n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11731,
         n11732, n11733, n11734, n11735, n11736, n11737, n11738, n11739,
         n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747,
         n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755,
         n11756, n11757, n11758, n11759, n11760, n11761, n11762, n11763,
         n11764, n11765, n11766, n11767, n11768, n11769, n11770, n11771,
         n11772, n11773, n11774, n11775, n11776, n11777, n11778, n11779,
         n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787,
         n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795,
         n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803,
         n11804, n11805, n11806, n11807, n11808, n11809, n11810, n11811,
         n11812, n11813, n11814, n11815, n11816, n11817, n11818, n11819,
         n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827,
         n11828, n11829, n11830, n11831, n11832, n11833, n11834, n11835,
         n11836, n11837, n11838, n11839, n11840, n11841, n11842, n11843,
         n11844, n11845, n11846, n11847, n11848, n11849, n11850, n11851,
         n11852, n11853, n11854, n11855, n11856, n11857, n11858, n11859,
         n11860, n11861, n11862, n11863, n11864, n11865, n11866, n11867,
         n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875,
         n11876, n11877, n11878, n11879, n11880, n11881, n11882, n11883,
         n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891,
         n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899,
         n11900, n11901, n11902, n11903, n11904, n11905, n11906, n11907,
         n11908, n11909, n11910, n11911, n11912, n11913, n11914, n11915,
         n11916, n11917, n11918, n11919, n11920, n11921, n11922, n11923,
         n11924, n11925, n11926, n11927, n11928, n11929, n11930, n11931,
         n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939,
         n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947,
         n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955,
         n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963,
         n11964, n11965, n11966, n11967, n11968, n11969, n11970, n11971,
         n11972, n11973, n11974, n11975, n11976, n11977, n11978, n11979,
         n11980, n11981, n11982, n11983, n11984, n11985, n11986, n11987,
         n11988, n11989, n11990, n11991, n11992, n11993, n11994, n11995,
         n11996, n11997, n11998, n11999, n12000, n12001, n12002, n12003,
         n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011,
         n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019,
         n12020, n12021, n12022, n12023, n12024, n12025, n12026, n12027,
         n12028, n12029, n12030, n12031, n12032, n12033, n12034, n12035,
         n12036, n12037, n12038, n12039, n12040, n12041, n12042, n12043,
         n12044, n12045, n12046, n12047, n12048, n12049, n12050, n12051,
         n12052, n12053, n12054, n12055, n12056, n12057, n12058, n12059,
         n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067,
         n12068, n12069, n12070, n12071, n12072, n12073, n12074, n12075,
         n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083,
         n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091,
         n12092, n12093, n12094, n12095, n12096, n12097, n12098, n12099,
         n12100, n12101, n12102, n12103, n12104, n12105, n12106, n12107,
         n12108, n12109, n12110, n12111, n12112, n12113, n12114, n12115,
         n12116, n12117, n12118, n12119, n12120, n12121, n12122, n12123,
         n12124, n12125, n12126, n12127, n12128, n12129, n12130, n12131,
         n12132, n12133, n12134, n12135, n12136, n12137, n12138, n12139,
         n12140, n12141, n12142, n12143, n12144, n12145, n12146, n12147,
         n12148, n12149, n12150, n12151, n12152, n12153, n12154, n12155,
         n12156, n12157, n12158, n12159, n12160, n12161, n12162, n12163,
         n12164, n12165, n12166, n12167, n12168, n12169, n12170, n12171,
         n12172, n12173, n12174, n12175, n12176, n12177, n12178, n12179,
         n12180, n12181, n12182, n12183, n12184, n12185, n12186, n12187,
         n12188, n12189, n12190, n12191, n12192, n12193, n12194, n12195,
         n12196, n12197, n12198, n12199, n12200, n12201, n12202, n12203,
         n12204, n12205, n12206, n12207, n12208, n12209, n12210, n12211,
         n12212, n12213, n12214, n12215, n12216, n12217, n12218, n12219,
         n12220, n12221, n12222, n12223, n12224, n12225, n12226, n12227,
         n12228, n12229, n12230, n12231, n12232, n12233, n12234, n12235,
         n12236, n12237, n12238, n12239, n12240, n12241, n12242, n12243,
         n12244, n12245, n12246, n12247, n12248, n12249, n12250, n12251,
         n12252, n12253, n12254, n12255, n12256, n12257, n12258, n12259,
         n12260, n12261, n12262, n12263, n12264, n12265, n12266, n12267,
         n12268, n12269, n12270, n12271, n12272, n12273, n12274, n12275,
         n12276, n12277, n12278, n12279, n12280, n12281, n12282, n12283,
         n12284, n12285, n12286, n12287, n12288, n12289, n12290, n12291,
         n12292, n12293, n12294, n12295, n12296, n12297, n12298, n12299,
         n12300, n12301, n12302, n12303, n12304, n12305, n12306, n12307,
         n12308, n12309, n12310, n12311, n12312, n12313, n12314, n12315,
         n12316, n12317, n12318, n12319, n12320, n12321, n12322, n12323,
         n12324, n12325, n12326, n12327, n12328, n12329, n12330, n12331,
         n12332, n12333, n12334, n12335, n12336, n12337, n12338, n12339,
         n12340, n12341, n12342, n12343, n12344, n12345, n12346, n12347,
         n12348, n12349, n12350, n12351, n12352, n12353, n12354, n12355,
         n12356, n12357, n12358, n12359, n12360, n12361, n12362, n12363,
         n12364, n12365, n12366, n12367, n12368, n12369, n12370, n12371,
         n12372, n12373, n12374, n12375, n12376, n12377, n12378, n12379,
         n12380, n12381, n12382, n12383, n12384, n12385, n12386, n12387,
         n12388, n12389, n12390, n12391, n12392, n12393, n12394, n12395,
         n12396, n12397, n12398, n12399, n12400, n12401, n12402, n12403,
         n12404, n12405, n12406, n12407, n12408, n12409, n12410, n12411,
         n12412, n12413, n12414, n12415, n12416, n12417, n12418, n12419,
         n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427,
         n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435,
         n12436, n12437, n12438, n12439, n12440, n12441, n12442, n12443,
         n12444, n12445, n12446, n12447, n12448, n12449, n12450, n12451,
         n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459,
         n12460, n12461, n12462, n12463, n12464, n12465, n12466, n12467,
         n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475,
         n12476, n12477, n12478, n12479, n12480, n12481, n12482, n12483,
         n12484, n12485, n12486, n12487, n12488, n12489, n12490, n12491,
         n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499,
         n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507,
         n12508, n12509, n12510, n12511, n12512, n12513, n12514, n12515,
         n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523,
         n12524, n12525, n12526, n12527, n12528, n12529, n12530, n12531,
         n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12539,
         n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547,
         n12548, n12549, n12550, n12551, n12552, n12553, n12554, n12555,
         n12556, n12557, n12558, n12559, n12560, n12561, n12562, n12563,
         n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571,
         n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579,
         n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12587,
         n12588, n12589, n12590, n12591, n12592, n12593, n12594, n12595,
         n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603,
         n12604, n12605, n12606, n12607, n12608, n12609, n12610, n12611,
         n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619,
         n12620, n12621, n12622, n12623, n12624, n12625, n12626, n12627,
         n12628, n12629, n12630, n12631, n12632, n12633, n12634, n12635,
         n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643,
         n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651,
         n12652, n12653, n12654, n12655, n12656, n12657, n12658, n12659,
         n12660, n12661, n12662, n12663, n12664, n12665, n12666, n12667,
         n12668, n12669, n12670, n12671, n12672, n12673, n12674, n12675,
         n12676, n12677, n12678, n12679, n12680, n12681, n12682, n12683,
         n12684, n12685, n12686, n12687, n12688, n12689, n12690, n12691,
         n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699,
         n12700, n12701, n12702, n12703, n12704, n12705, n12706, n12707,
         n12708, n12709, n12710, n12711, n12712, n12713, n12714, n12715,
         n12716, n12717, n12718, n12719, n12720, n12721, n12722, n12723,
         n12724, n12725, n12726, n12727, n12728, n12729, n12730, n12731,
         n12732, n12733, n12734, n12735, n12736, n12737, n12738, n12739,
         n12740, n12741, n12742, n12743, n12744, n12745, n12746, n12747,
         n12748, n12749, n12750, n12751, n12752, n12753, n12754, n12755,
         n12756, n12757, n12758, n12759, n12760, n12761, n12762, n12763,
         n12764, n12765, n12766, n12767, n12768, n12769, n12770, n12771,
         n12772, n12773, n12774, n12775, n12776, n12777, n12778, n12779,
         n12780, n12781, n12782, n12783, n12784, n12785, n12786, n12787,
         n12788, n12789, n12790, n12791, n12792, n12793, n12794, n12795,
         n12796, n12797, n12798, n12799, n12800, n12801, n12802, n12803,
         n12804, n12805, n12806, n12807, n12808, n12809, n12810, n12811,
         n12812, n12813, n12814, n12815, n12816, n12817, n12818, n12819,
         n12820, n12821, n12822, n12823, n12824, n12825, n12826, n12827,
         n12828, n12829, n12830, n12831, n12832, n12833, n12834, n12835,
         n12836, n12837, n12838, n12839, n12840, n12841, n12842, n12843,
         n12844, n12845, n12846, n12847, n12848, n12849, n12850, n12851,
         n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859,
         n12860, n12861, n12862, n12863, n12864, n12865, n12866, n12867,
         n12868, n12869, n12870, n12871, n12872, n12873, n12874, n12875,
         n12876, n12877, n12878, n12879, n12880, n12881, n12882, n12883,
         n12884, n12885, n12886, n12887, n12888, n12889, n12890, n12891,
         n12892, n12893, n12894, n12895, n12896, n12897, n12898, n12899,
         n12900, n12901, n12902, n12903, n12904, n12905, n12906, n12907,
         n12908, n12909, n12910, n12911, n12912, n12913, n12914, n12915,
         n12916, n12917, n12918, n12919, n12920, n12921, n12922, n12923,
         n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931,
         n12932, n12933, n12934, n12935, n12936, n12937, n12938, n12939,
         n12940, n12941, n12942, n12943, n12944, n12945, n12946, n12947,
         n12948, n12949, n12950, n12951, n12952, n12953, n12954, n12955,
         n12956, n12957, n12958, n12959, n12960, n12961, n12962, n12963,
         n12964, n12965, n12966, n12967, n12968, n12969, n12970, n12971,
         n12972, n12973, n12974, n12975, n12976, n12977, n12978, n12979,
         n12980, n12981, n12982, n12983, n12984, n12985, n12986, n12987,
         n12988, n12989, n12990, n12991, n12992, n12993, n12994, n12995,
         n12996, n12997, n12998, n12999, n13000, n13001, n13002, n13003,
         n13004, n13005, n13006, n13007, n13008, n13009, n13010, n13011,
         n13012, n13013, n13014, n13015, n13016, n13017, n13018, n13019,
         n13020, n13021, n13022, n13023, n13024, n13025, n13026, n13027,
         n13028, n13029, n13030, n13031, n13032, n13033, n13034, n13035,
         n13036, n13037, n13038, n13039, n13040, n13041, n13042, n13043,
         n13044, n13045, n13046, n13047, n13048, n13049, n13050, n13051,
         n13052, n13053, n13054, n13055, n13056, n13057, n13058, n13059,
         n13060, n13061, n13062, n13063, n13064, n13065, n13066, n13067,
         n13068, n13069, n13070, n13071, n13072, n13073, n13074, n13075,
         n13076, n13077, n13078, n13079, n13080, n13081, n13082, n13083,
         n13084, n13085, n13086, n13087, n13088, n13089, n13090, n13091,
         n13092, n13093, n13094, n13095, n13096, n13097, n13098, n13099,
         n13100, n13101, n13102, n13103, n13104, n13105, n13106, n13107,
         n13108, n13109, n13110, n13111, n13112, n13113, n13114, n13115,
         n13116, n13117, n13118, n13119, n13120, n13121, n13122, n13123,
         n13124, n13125, n13126, n13127, n13128, n13129, n13130, n13131,
         n13132, n13133, n13134, n13135, n13136, n13137, n13138, n13139,
         n13140, n13141, n13142, n13143, n13144, n13145, n13146, n13147,
         n13148, n13149, n13150, n13151, n13152, n13153, n13154, n13155,
         n13156, n13157, n13158, n13159, n13160, n13161, n13162, n13163,
         n13164, n13165, n13166, n13167, n13168, n13169, n13170, n13171,
         n13172, n13173, n13174, n13175, n13176, n13177, n13178, n13179,
         n13180, n13181, n13182, n13183, n13184, n13185, n13186, n13187,
         n13188, n13189, n13190, n13191, n13192, n13193, n13194, n13195,
         n13196, n13197, n13198, n13199, n13200, n13201, n13202, n13203,
         n13204, n13205, n13206, n13207, n13208, n13209, n13211, n13212,
         n13213, n13214, n13215, n13216, n13217, n13218, n13219, n13220,
         n13221, n13222, n13223, n13224, n13225, n13226, n13227, n13228,
         n13229, n13230, n13231, n13232, n13233, n13234, n13235, n13236,
         n13237, n13238, n13239, n13240, n13241, n13242, n13243, n13244,
         n13245, n13246, n13247, n13248, n13249, n13250, n13251, n13252,
         n13253, n13254, n13255, n13256, n13257, n13258, n13259, n13260,
         n13261, n13262, n13263, n13264, n13265, n13266, n13267, n13268,
         n13269, n13270, n13271, n13272, n13273, n13274, n13275, n13276,
         n13277, n13278, n13279, n13280, n13281, n13282, n13283, n13284,
         n13285, n13286, n13287, n13288, n13289, n13290, n13291, n13292,
         n13293, n13294, n13295, n13296, n13297, n13298, n13299, n13300,
         n13301, n13302, n13303, n13304, n13305, n13306, n13307, n13308,
         n13309, n13310, n13311, n13312, n13313, n13314, n13315, n13316,
         n13317, n13318, n13319, n13320, n13321, n13322, n13323, n13324,
         n13325, n13326, n13327, n13328, n13329, n13330, n13331, n13332,
         n13333, n13334, n13335, n13336, n13337, n13338, n13339, n13340,
         n13341, n13342, n13343, n13344, n13345, n13346, n13347, n13348,
         n13349, n13350, n13351, n13352, n13353, n13354, n13355, n13356,
         n13357, n13358, n13359, n13360, n13361, n13362, n13363, n13364,
         n13365, n13366, n13367, n13368, n13369, n13370, n13371, n13372,
         n13373, n13374, n13375, n13376, n13377, n13378, n13379, n13380,
         n13381, n13382, n13383, n13384, n13385, n13386, n13387, n13388,
         n13389, n13390, n13391, n13392, n13393, n13394, n13395, n13396,
         n13397, n13398, n13399, n13400, n13401, n13402, n13403, n13404,
         n13405, n13406, n13407, n13408, n13409, n13410, n13411, n13412,
         n13413, n13414, n13415, n13416, n13417, n13418, n13419, n13420,
         n13421, n13422, n13423, n13424, n13425, n13426, n13427, n13428,
         n13429, n13430, n13431, n13432, n13433, n13434, n13435, n13436,
         n13437, n13438, n13439, n13440, n13441, n13442, n13443, n13444,
         n13445, n13446, n13447, n13448, n13449, n13450, n13451, n13452,
         n13453, n13454, n13455, n13456, n13457, n13458, n13459, n13460,
         n13461, n13462, n13463, n13464, n13465, n13466, n13467, n13468,
         n13469, n13470, n13471, n13472, n13473, n13474, n13475, n13476,
         n13477, n13478, n13479, n13480, n13481, n13482, n13483, n13484,
         n13485, n13486, n13487, n13488, n13489, n13490, n13491, n13492,
         n13493, n13494, n13495, n13496, n13497, n13498, n13499, n13500,
         n13501, n13502, n13503, n13504, n13505, n13506, n13507, n13508,
         n13509, n13510, n13511, n13512, n13513, n13514, n13515, n13516,
         n13517, n13518, n13519, n13520, n13521, n13522, n13523, n13524,
         n13525, n13526, n13527, n13528, n13529, n13530, n13531, n13532,
         n13533, n13534, n13535, n13536, n13537, n13538, n13539, n13540,
         n13541, n13542, n13543, n13544, n13545, n13546, n13547, n13548,
         n13549, n13550, n13551, n13552, n13553, n13554, n13555, n13556,
         n13557, n13558, n13559, n13560, n13561, n13562, n13563, n13564,
         n13565, n13566, n13567, n13568, n13569, n13570, n13571, n13572,
         n13573, n13574, n13575, n13576, n13577, n13578, n13579, n13580,
         n13581, n13582, n13583, n13584, n13585, n13586, n13587, n13588,
         n13589, n13590, n13591, n13592, n13593, n13594, n13595, n13596,
         n13597, n13598, n13599, n13600, n13601, n13602, n13603, n13604,
         n13605, n13606, n13607, n13608, n13609, n13610, n13611, n13612,
         n13613, n13614, n13615, n13616, n13617, n13618, n13619, n13620,
         n13621, n13622, n13623, n13624, n13625, n13626, n13627, n13628,
         n13629, n13630, n13631, n13632, n13633, n13634, n13635, n13636,
         n13637, n13638, n13639, n13640, n13641, n13642, n13643, n13644,
         n13645, n13646, n13647, n13648, n13649, n13650, n13651, n13652,
         n13653, n13654, n13655, n13656, n13657, n13658, n13659, n13660,
         n13661, n13662, n13663, n13664, n13665, n13666, n13667, n13668,
         n13669, n13670, n13671, n13672, n13673, n13674, n13675, n13676,
         n13677, n13678, n13679, n13680, n13681, n13682, n13683, n13684,
         n13685, n13686, n13687, n13688, n13689, n13690, n13691, n13692,
         n13693, n13694, n13695, n13696, n13697, n13698, n13699, n13700,
         n13701, n13702, n13703, n13704, n13705, n13706, n13707, n13708,
         n13709, n13710, n13711, n13712, n13713, n13714, n13715, n13716,
         n13717, n13718, n13719, n13720, n13721, n13722, n13723, n13724,
         n13725, n13726, n13727, n13728, n13729, n13730, n13731, n13732,
         n13733, n13734, n13735, n13736, n13737, n13738, n13739, n13740,
         n13741, n13742, n13743, n13744, n13745, n13746, n13747, n13748,
         n13749, n13750, n13751, n13752, n13753, n13754, n13755, n13756,
         n13757, n13758, n13759, n13760, n13761, n13762, n13763, n13764,
         n13765, n13766, n13767, n13768, n13769, n13770, n13771, n13772,
         n13773, n13774, n13775, n13776, n13777, n13778, n13779, n13780,
         n13781, n13782, n13783, n13784, n13785, n13786, n13787, n13788,
         n13789, n13790, n13791, n13792, n13793, n13794, n13795, n13796,
         n13797, n13798, n13799, n13800, n13801, n13802, n13803, n13804,
         n13805, n13806, n13807, n13808, n13809, n13810, n13811, n13812,
         n13813, n13814, n13815, n13816, n13817, n13818, n13819, n13820,
         n13821, n13822, n13823, n13824, n13825, n13826, n13827, n13828,
         n13829, n13830, n13831, n13832, n13833, n13834, n13835, n13836,
         n13837, n13838, n13839, n13840, n13841, n13842, n13843, n13844,
         n13845, n13846, n13847, n13848, n13849, n13850, n13851, n13852,
         n13853, n13854, n13855, n13856, n13857, n13858, n13859, n13860,
         n13861, n13862, n13863, n13864, n13865, n13866, n13867, n13868,
         n13869, n13870, n13871, n13872, n13873, n13874, n13875, n13876,
         n13877, n13878, n13879, n13880, n13881, n13882, n13883, n13884,
         n13885, n13886, n13887, n13888, n13889, n13890, n13891, n13892,
         n13893, n13894, n13895, n13896, n13897, n13898, n13900, n13901,
         n13902, n13903, n13904, n13905, n13906, n13907, n13908, n13909,
         n13910, n13911, n13912, n13913, n13914, n13915, n13916, n13917,
         n13918, n13919, n13920, n13921, n13922, n13923, n13924, n13925,
         n13926, n13927, n13928, n13929, n13930, n13931, n13932, n13933,
         n13934, n13935, n13936, n13937, n13938, n13939, n13940, n13941,
         n13942, n13943, n13944, n13945, n13946, n13947, n13948, n13949,
         n13950, n13951, n13952, n13953, n13954, n13955, n13956, n13957,
         n13958, n13959, n13960, n13961, n13962, n13963, n13964, n13965,
         n13966, n13967, n13968, n13969, n13970, n13971, n13972, n13973,
         n13974, n13975, n13976, n13977, n13978, n13979, n13980, n13981,
         n13982, n13983, n13984, n13985, n13986, n13987, n13988, n13989,
         n13990, n13991, n13992, n13993, n13994, n13995, n13996, n13997,
         n13998, n13999, n14000, n14001, n14002, n14003, n14004, n14005,
         n14006, n14007, n14008, n14009, n14010, n14011, n14012, n14013,
         n14014, n14015, n14016, n14017, n14018, n14019, n14020, n14021,
         n14022, n14023, n14024, n14025, n14026, n14027, n14028, n14029,
         n14030, n14031, n14032, n14033, n14034, n14035, n14036, n14037,
         n14038, n14039, n14040, n14041, n14042, n14043, n14044, n14045,
         n14046, n14047, n14048, n14049, n14050, n14051, n14052, n14053,
         n14054, n14055, n14056, n14057, n14058, n14059, n14060, n14061,
         n14062, n14063, n14064, n14065, n14066, n14067, n14068, n14069,
         n14070, n14071, n14072, n14073, n14074, n14075, n14076, n14077,
         n14078, n14079, n14080, n14081, n14082, n14083, n14084, n14085,
         n14086, n14087, n14088, n14089, n14090, n14091, n14092, n14093,
         n14094, n14095, n14096, n14097, n14098, n14099, n14100, n14101,
         n14102, n14103, n14104, n14105, n14106, n14107, n14108, n14109,
         n14110, n14111, n14112, n14113, n14114, n14115, n14116, n14117,
         n14118, n14119, n14120, n14121, n14122, n14123, n14124, n14125,
         n14126, n14127, n14128, n14129, n14130, n14131, n14132, n14133,
         n14134, n14135, n14136, n14137, n14138, n14139, n14140, n14141,
         n14142, n14143, n14144, n14145, n14146, n14147, n14148, n14149,
         n14150, n14151, n14152, n14153, n14154, n14155, n14156, n14157,
         n14158, n14159, n14160, n14161, n14162, n14163, n14164, n14165,
         n14166, n14167, n14168, n14169, n14170, n14171, n14172, n14173,
         n14174, n14175, n14176, n14177, n14178, n14179, n14180, n14181,
         n14182, n14183, n14184, n14185, n14186, n14187, n14188, n14189,
         n14190, n14191, n14192, n14193, n14194, n14195, n14196, n14197,
         n14198, n14199, n14200, n14201, n14202, n14203, n14204, n14205,
         n14206, n14207, n14208, n14209, n14210, n14211, n14212, n14213,
         n14214, n14215, n14216, n14217, n14218, n14219, n14220, n14221,
         n14222, n14223, n14224, n14225, n14226, n14227, n14228, n14229,
         n14230, n14231, n14232, n14233, n14234, n14235, n14236, n14237,
         n14238, n14239, n14240, n14241, n14242, n14243, n14244, n14245,
         n14246, n14247, n14248, n14249, n14250, n14251, n14252, n14253,
         n14254, n14255, n14256, n14257, n14258, n14259, n14260, n14261,
         n14262, n14263, n14264, n14265, n14266, n14267, n14268, n14269,
         n14270, n14271, n14272, n14273, n14274, n14275, n14276, n14277,
         n14278, n14279, n14280, n14281, n14282, n14283, n14284, n14285,
         n14286, n14287, n14288, n14289, n14290, n14291, n14292, n14293,
         n14294, n14295, n14296, n14297, n14298, n14299, n14300, n14301,
         n14302, n14303, n14304, n14305, n14306, n14307, n14308, n14309,
         n14310, n14311, n14312, n14313, n14314, n14315, n14316, n14317,
         n14318, n14319, n14320, n14321, n14322, n14323, n14324, n14325,
         n14326, n14327, n14328, n14329, n14330, n14331, n14332, n14333,
         n14334, n14335, n14336, n14337, n14338, n14339, n14340, n14341,
         n14342, n14343, n14344, n14345, n14346, n14347, n14348, n14349,
         n14350, n14351, n14352, n14353, n14354, n14355, n14356, n14357,
         n14358, n14359, n14360, n14361, n14362, n14363, n14364, n14365,
         n14366, n14367, n14368, n14369, n14370, n14371, n14372, n14373,
         n14374, n14375, n14376, n14377, n14378, n14379, n14380, n14381,
         n14382, n14383, n14384, n14385, n14386, n14387, n14388, n14389,
         n14390, n14391, n14392, n14393, n14394, n14395, n14396, n14397,
         n14398, n14399, n14400, n14401, n14402, n14403, n14404, n14405,
         n14406, n14407, n14408, n14409, n14410, n14411, n14412, n14413,
         n14414, n14415, n14416, n14417, n14418, n14419, n14420, n14421,
         n14422, n14423, n14424, n14425, n14426, n14427, n14428, n14429,
         n14430, n14431, n14432, n14433, n14434, n14435, n14437, n14438,
         n14439, n14440, n14441, n14442, n14443, n14444, n14445, n14446,
         n14447, n14448, n14449, n14450, n14451, n14452, n14453, n14454,
         n14455, n14456, n14457, n14458, n14459, n14460, n14461, n14462,
         n14463, n14464, n14465, n14466, n14467, n14468, n14469, n14470,
         n14471, n14472, n14473, n14474, n14475, n14476, n14477, n14478,
         n14479, n14480, n14481, n14482, n14483, n14484, n14485, n14486,
         n14487, n14488, n14489, n14490, n14491, n14492, n14493, n14494,
         n14495, n14496, n14497, n14498, n14499, n14500, n14501, n14502,
         n14503, n14504, n14505, n14506, n14507, n14508, n14509, n14510,
         n14511, n14512, n14513, n14514, n14515, n14516, n14517, n14518,
         n14519, n14520, n14521, n14522, n14523, n14524, n14525, n14526,
         n14527, n14528, n14529, n14530, n14531, n14532, n14533, n14534,
         n14535, n14536, n14537, n14538, n14539, n14540, n14541, n14542,
         n14543, n14544, n14545, n14546, n14547, n14548, n14549, n14550,
         n14551, n14552, n14553, n14554, n14555, n14556, n14557, n14558,
         n14559, n14560, n14561, n14562, n14563, n14564, n14565, n14566,
         n14567, n14568, n14569, n14570, n14571, n14572, n14573, n14574,
         n14575, n14576, n14577, n14578, n14579, n14580, n14581, n14582,
         n14583, n14584, n14585, n14586, n14587, n14588, n14589, n14590,
         n14591, n14592, n14593, n14594, n14595, n14596, n14597, n14598,
         n14599, n14600, n14601, n14602, n14603, n14604, n14605, n14606,
         n14607, n14608, n14609, n14610, n14611, n14612, n14613, n14614,
         n14615, n14616, n14617, n14618, n14619, n14620, n14621, n14622,
         n14623, n14624, n14625, n14626, n14627, n14628, n14629, n14630,
         n14631, n14632, n14633, n14634, n14635, n14636, n14637, n14638,
         n14639, n14640, n14641, n14642, n14643, n14644, n14645, n14646,
         n14647, n14648, n14649, n14650, n14651, n14652, n14653, n14654,
         n14655, n14656, n14657, n14658, n14659, n14660, n14661, n14662,
         n14663, n14664, n14665, n14666, n14667, n14668, n14669, n14670,
         n14671, n14672, n14673, n14674, n14675, n14676, n14677, n14678,
         n14679, n14680, n14681, n14682, n14683, n14684, n14685, n14686,
         n14687, n14688, n14689, n14690, n14691, n14692, n14693, n14694,
         n14695, n14696, n14697, n14698, n14699, n14700, n14701, n14702,
         n14703, n14704, n14705, n14706, n14707, n14708, n14709, n14710,
         n14711, n14712, n14713, n14714, n14715, n14716, n14717, n14718,
         n14719, n14720, n14721, n14722, n14723, n14724, n14725, n14726,
         n14727, n14728, n14729, n14730, n14731, n14732, n14733, n14734,
         n14735, n14736, n14737, n14738, n14739, n14740, n14741, n14742,
         n14743, n14744, n14745, n14746, n14747, n14748, n14749, n14750,
         n14751, n14752, n14753, n14754, n14755, n14756, n14757, n14758,
         n14759, n14760, n14761, n14762, n14763, n14764, n14765, n14766,
         n14767, n14768, n14769, n14770, n14771, n14772, n14773, n14774,
         n14775, n14776, n14777, n14778, n14779, n14780, n14781, n14782,
         n14783, n14784, n14785, n14786, n14787, n14788, n14789, n14790,
         n14791, n14792, n14793, n14794, n14795, n14796, n14797, n14798,
         n14799, n14800, n14801, n14802, n14803, n14804, n14805, n14806,
         n14807, n14808, n14809, n14810, n14811, n14812, n14813, n14814,
         n14815, n14816, n14817, n14818, n14819, n14820, n14821, n14822,
         n14823, n14824, n14825, n14826, n14827, n14828, n14829, n14830,
         n14831, n14832, n14833, n14834, n14835, n14836, n14837, n14838,
         n14839, n14840, n14841, n14842, n14843, n14844, n14845, n14846,
         n14847, n14848, n14849, n14850, n14851, n14852, n14853, n14854,
         n14855, n14856, n14857, n14858, n14859, n14860, n14861, n14862,
         n14863, n14864, n14865, n14866, n14867, n14868, n14869, n14870,
         n14871, n14872, n14873, n14874, n14875, n14876, n14877, n14878,
         n14879, n14880, n14881, n14882, n14883, n14884, n14885, n14886,
         n14887, n14888, n14889, n14890, n14891, n14892, n14893, n14894,
         n14895, n14896, n14897, n14898, n14899, n14900, n14901, n14902,
         n14903, n14904, n14905, n14906, n14907, n14908, n14909, n14910,
         n14911, n14912, n14913, n14914, n14915, n14916, n14917, n14918,
         n14919, n14920, n14921, n14922, n14923, n14924, n14925, n14926,
         n14927, n14928, n14929, n14930, n14931, n14932, n14933, n14934,
         n14935, n14936, n14937, n14938, n14939, n14940, n14941, n14942,
         n14943, n14944, n14945, n14946, n14947, n14948, n14949, n14950,
         n14951, n14952, n14953, n14954, n14955, n14956, n14957, n14958,
         n14959, n14960, n14961, n14962, n14963, n14964, n14965, n14966,
         n14967, n14968, n14969, n14970, n14971, n14972, n14973, n14974,
         n14975, n14976, n14977, n14978, n14979, n14980, n14981, n14982,
         n14983, n14984, n14985, n14986, n14987, n14988, n14989, n14990,
         n14991, n14992, n14993, n14994, n14995, n14996, n14997, n14998,
         n14999, n15000, n15001, n15002, n15003, n15004, n15005, n15006,
         n15007, n15008, n15009, n15010, n15011, n15012, n15013, n15014,
         n15015, n15016, n15017, n15018, n15019, n15020, n15021, n15022,
         n15023, n15024, n15025, n15026, n15027, n15028, n15029, n15030,
         n15031, n15032, n15033, n15034, n15035, n15036, n15037, n15038,
         n15039, n15040, n15041, n15042, n15043, n15044, n15045, n15046,
         n15047, n15048, n15049, n15050, n15051, n15052, n15053, n15054,
         n15055, n15056, n15057, n15058, n15059, n15060, n15061, n15062,
         n15063, n15064, n15065, n15066, n15067, n15068, n15069, n15070,
         n15071, n15072, n15073, n15074, n15075, n15076, n15077, n15078,
         n15079, n15080, n15081, n15082, n15083, n15084, n15085, n15086,
         n15087, n15088, n15089, n15090, n15091, n15092, n15093, n15094,
         n15095, n15096, n15097, n15098, n15099, n15100, n15101, n15102,
         n15103, n15104, n15105, n15106, n15107, n15108, n15109, n15110,
         n15111, n15112, n15113, n15114, n15115, n15116, n15117, n15118,
         n15119, n15120, n15121, n15122, n15123, n15124, n15125, n15126,
         n15127, n15128, n15129, n15130, n15131, n15132, n15133, n15134,
         n15135, n15136, n15137, n15138, n15139, n15140, n15141, n15142,
         n15143, n15144, n15145, n15146, n15147, n15148, n15149, n15150,
         n15151, n15152, n15153, n15154, n15155, n15156, n15157, n15158,
         n15159, n15160, n15161, n15162, n15163, n15164, n15165, n15166,
         n15167, n15168, n15169, n15170, n15171, n15172, n15173, n15174,
         n15175, n15176, n15177, n15178, n15179, n15180, n15181, n15182,
         n15183, n15184, n15185, n15186, n15187, n15188, n15189, n15190,
         n15191, n15192, n15193, n15194, n15195, n15196, n15197, n15198,
         n15199, n15200, n15201, n15202, n15203, n15204, n15205, n15206,
         n15207, n15208, n15209, n15210, n15211, n15212, n15213, n15214,
         n15215, n15216, n15217, n15218, n15219, n15220, n15221, n15222,
         n15223, n15224, n15225, n15226, n15227, n15228, n15229, n15230,
         n15231, n15232, n15233, n15234, n15235, n15236, n15237, n15238,
         n15239, n15240, n15241, n15242, n15243, n15244, n15245, n15246,
         n15247, n15248, n15249, n15250, n15251, n15252, n15253, n15254,
         n15255, n15256, n15257, n15258, n15259, n15260, n15261, n15262,
         n15263, n15264, n15265, n15266, n15267, n15268, n15269, n15270,
         n15271, n15272, n15273, n15274, n15275, n15276, n15277, n15278,
         n15279, n15280, n15281, n15282, n15283, n15284, n15285, n15286,
         n15287, n15288, n15289, n15290, n15291, n15292, n15293, n15294,
         n15295, n15296, n15297, n15298, n15299, n15300, n15301, n15302,
         n15303, n15304, n15305, n15306, n15307, n15308, n15309, n15310,
         n15311, n15312, n15313, n15314, n15315, n15316, n15317, n15318,
         n15319, n15320, n15321, n15322, n15323, n15324, n15325, n15326,
         n15327, n15328, n15329, n15330, n15331, n15332, n15333, n15334,
         n15335, n15336, n15337, n15338, n15339, n15340, n15341, n15342,
         n15343, n15344, n15345, n15346, n15347, n15348, n15349, n15350,
         n15351, n15352, n15353, n15354, n15355, n15356, n15357, n15358,
         n15359, n15360, n15361, n15362, n15363, n15364, n15365, n15366,
         n15367, n15368, n15369, n15370, n15371, n15372, n15373, n15374,
         n15375, n15376, n15377, n15378, n15379, n15380, n15381, n15382,
         n15383, n15384, n15385, n15386, n15387, n15388, n15389, n15390,
         n15391, n15392, n15393, n15394, n15395, n15396, n15397, n15398,
         n15399, n15400, n15401, n15402, n15403, n15404, n15405, n15406,
         n15407, n15408, n15409, n15410, n15411, n15412, n15413, n15414,
         n15415, n15416, n15417, n15418, n15419, n15420, n15421, n15422,
         n15423, n15424, n15425, n15426, n15427, n15428, n15429, n15430,
         n15431, n15432, n15433, n15434, n15435, n15436, n15437, n15438,
         n15439, n15440, n15441, n15442, n15443, n15444, n15445, n15446,
         n15447, n15448, n15449, n15450, n15451, n15452, n15453, n15454,
         n15455, n15456, n15457, n15458, n15459, n15460, n15461, n15462,
         n15463, n15464, n15465, n15466, n15467, n15468, n15469, n15470,
         n15471, n15472, n15473, n15474, n15475, n15476, n15477, n15478,
         n15479, n15480, n15481, n15482, n15483, n15484, n15485, n15486,
         n15487, n15488, n15489, n15490, n15491, n15492, n15493, n15494,
         n15495, n15496, n15497, n15498, n15499, n15500, n15501, n15502,
         n15503, n15504, n15505, n15506, n15507, n15508, n15509, n15510,
         n15511, n15512, n15513, n15514, n15515, n15516, n15517, n15518,
         n15519, n15520, n15521, n15522, n15523, n15524, n15525, n15526,
         n15527, n15528, n15529, n15530, n15531, n15532;

  INV_X4 U7293 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  XNOR2_X1 U7294 ( .A(n13244), .B(n6649), .ZN(n13262) );
  AND2_X1 U7295 ( .A1(n9019), .A2(n9018), .ZN(n12375) );
  CLKBUF_X2 U7296 ( .A(n10626), .Z(n11975) );
  NAND2_X1 U7298 ( .A1(n7800), .A2(n7799), .ZN(n7802) );
  NAND4_X1 U7299 ( .A1(n8534), .A2(n8533), .A3(n8532), .A4(n8531), .ZN(n15121)
         );
  INV_X1 U7300 ( .A(n6546), .ZN(n9524) );
  INV_X1 U7301 ( .A(n8385), .ZN(n8133) );
  BUF_X2 U7302 ( .A(n9172), .Z(n6546) );
  CLKBUF_X1 U7303 ( .A(n11034), .Z(n6549) );
  INV_X2 U7305 ( .A(n7602), .ZN(n9769) );
  CLKBUF_X2 U7306 ( .A(n12293), .Z(n12215) );
  INV_X1 U7307 ( .A(n8403), .ZN(n8376) );
  NAND2_X1 U7308 ( .A1(n9579), .A2(n10529), .ZN(n12289) );
  NAND3_X1 U7309 ( .A1(n7544), .A2(n7689), .A3(n10178), .ZN(n14766) );
  NAND2_X1 U7310 ( .A1(n10804), .A2(n12859), .ZN(n9740) );
  INV_X1 U7311 ( .A(n11938), .ZN(n11979) );
  NAND2_X1 U7312 ( .A1(n14439), .A2(n14061), .ZN(n8149) );
  XNOR2_X1 U7313 ( .A(n10862), .B(n10900), .ZN(n12331) );
  INV_X1 U7314 ( .A(n12381), .ZN(n9065) );
  INV_X1 U7315 ( .A(n12560), .ZN(n12881) );
  OAI21_X1 U7316 ( .B1(n11717), .B2(n12490), .A(n12489), .ZN(n11794) );
  OAI21_X1 U7317 ( .B1(n8775), .B2(n8774), .A(n8776), .ZN(n8796) );
  AND2_X2 U7318 ( .A1(n6552), .A2(n12612), .ZN(n12162) );
  CLKBUF_X2 U7319 ( .A(n7699), .Z(n8385) );
  NAND2_X1 U7320 ( .A1(n8984), .A2(n8983), .ZN(n13084) );
  AOI21_X2 U7321 ( .B1(n13789), .B2(n13790), .A(n6904), .ZN(n13848) );
  NOR2_X1 U7322 ( .A1(n14067), .A2(n14793), .ZN(n14288) );
  NOR2_X1 U7323 ( .A1(n15027), .A2(P1_ADDR_REG_0__SCAN_IN), .ZN(n14490) );
  AND2_X1 U7324 ( .A1(n8933), .A2(n8932), .ZN(n13159) );
  INV_X1 U7325 ( .A(n13884), .ZN(n10519) );
  XNOR2_X1 U7326 ( .A(n8144), .B(n8143), .ZN(n12608) );
  AND3_X1 U7327 ( .A1(n7445), .A2(n9084), .A3(n8519), .ZN(n6545) );
  NAND2_X2 U7328 ( .A1(n8158), .A2(n13962), .ZN(n7716) );
  NAND2_X2 U7329 ( .A1(n11352), .A2(n7513), .ZN(n11631) );
  NAND4_X2 U7330 ( .A1(n7739), .A2(n7738), .A3(n7737), .A4(n7736), .ZN(n13938)
         );
  INV_X1 U7331 ( .A(n8601), .ZN(n8602) );
  NAND2_X2 U7332 ( .A1(n11184), .A2(n11186), .ZN(n11183) );
  OR2_X2 U7333 ( .A1(n15093), .A2(n7208), .ZN(n7206) );
  NAND2_X2 U7334 ( .A1(n7717), .A2(n6947), .ZN(n13884) );
  INV_X1 U7335 ( .A(n10379), .ZN(n7734) );
  XNOR2_X2 U7336 ( .A(n10691), .B(n10692), .ZN(n10690) );
  NAND2_X2 U7337 ( .A1(n10625), .A2(n10624), .ZN(n10691) );
  NAND2_X2 U7338 ( .A1(n13196), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8525) );
  AND2_X4 U7339 ( .A1(n7726), .A2(n7049), .ZN(n7733) );
  OR2_X2 U7340 ( .A1(n7727), .A2(n6713), .ZN(n7230) );
  OAI22_X2 U7341 ( .A1(n8649), .A2(n8648), .B1(P1_DATAO_REG_6__SCAN_IN), .B2(
        n9773), .ZN(n8652) );
  NAND2_X2 U7342 ( .A1(n11469), .A2(n7879), .ZN(n11354) );
  NAND2_X2 U7343 ( .A1(n7508), .A2(n6645), .ZN(n11469) );
  OAI21_X2 U7346 ( .B1(n8831), .B2(n8830), .A(n8833), .ZN(n8853) );
  NAND2_X2 U7347 ( .A1(n8814), .A2(n8813), .ZN(n8831) );
  BUF_X8 U7348 ( .A(n8637), .Z(n8988) );
  XNOR2_X2 U7349 ( .A(n12766), .B(n12783), .ZN(n12749) );
  NAND2_X1 U7350 ( .A1(n12612), .A2(n9149), .ZN(n9172) );
  NAND2_X2 U7351 ( .A1(n10278), .A2(n8437), .ZN(n10497) );
  NAND2_X2 U7352 ( .A1(n10298), .A2(n7735), .ZN(n10278) );
  XNOR2_X2 U7353 ( .A(n10577), .B(n10578), .ZN(n10576) );
  INV_X1 U7354 ( .A(n11940), .ZN(n6547) );
  XNOR2_X2 U7355 ( .A(n8148), .B(n8147), .ZN(n8152) );
  MUX2_X2 U7356 ( .A(P2_IR_REG_0__SCAN_IN), .B(n13781), .S(n9841), .Z(n12002)
         );
  NAND4_X2 U7357 ( .A1(n7649), .A2(n7743), .A3(n7648), .A4(n7506), .ZN(n7959)
         );
  OAI222_X1 U7358 ( .A1(n6551), .A2(n14437), .B1(P2_U3088), .B2(n9149), .C1(
        n15332), .C2(n13780), .ZN(P2_U3298) );
  INV_X1 U7359 ( .A(n9149), .ZN(n6552) );
  NAND2_X2 U7360 ( .A1(n7273), .A2(n8759), .ZN(n8775) );
  NAND2_X2 U7361 ( .A1(n6581), .A2(n7073), .ZN(n12016) );
  BUF_X1 U7362 ( .A(n11034), .Z(n6548) );
  OAI22_X2 U7363 ( .A1(n8576), .A2(n8575), .B1(P2_DATAO_REG_2__SCAN_IN), .B2(
        n10028), .ZN(n8589) );
  NAND2_X2 U7364 ( .A1(n7233), .A2(n8561), .ZN(n8576) );
  NOR4_X2 U7365 ( .A1(n12568), .A2(n12573), .A3(n12574), .A4(n12404), .ZN(
        n12405) );
  XOR2_X2 U7366 ( .A(n14520), .B(n14519), .Z(n14559) );
  NOR2_X4 U7367 ( .A1(n7276), .A2(n14516), .ZN(n14519) );
  OR2_X1 U7368 ( .A1(n8398), .A2(n8397), .ZN(n8413) );
  OR2_X1 U7369 ( .A1(n14146), .A2(n14400), .ZN(n14109) );
  NAND2_X1 U7370 ( .A1(n9493), .A2(n9492), .ZN(n13661) );
  NAND2_X1 U7371 ( .A1(n8081), .A2(n8080), .ZN(n14400) );
  AND2_X1 U7372 ( .A1(n8314), .A2(n8308), .ZN(n11633) );
  INV_X1 U7373 ( .A(n10631), .ZN(n10642) );
  INV_X4 U7374 ( .A(n8367), .ZN(n8403) );
  CLKBUF_X2 U7375 ( .A(P2_U3947), .Z(n6550) );
  BUF_X2 U7376 ( .A(n10354), .Z(n11938) );
  INV_X4 U7377 ( .A(n9115), .ZN(n12549) );
  BUF_X2 U7378 ( .A(n9032), .Z(n10792) );
  INV_X2 U7379 ( .A(n11939), .ZN(n10626) );
  NAND2_X1 U7380 ( .A1(n14792), .A2(n10352), .ZN(n10178) );
  CLKBUF_X1 U7381 ( .A(n10363), .Z(n13808) );
  INV_X1 U7382 ( .A(n14780), .ZN(n14760) );
  CLKBUF_X2 U7383 ( .A(n10428), .Z(n13282) );
  CLKBUF_X2 U7384 ( .A(n9476), .Z(n9525) );
  BUF_X2 U7385 ( .A(n7723), .Z(n8384) );
  NAND2_X2 U7386 ( .A1(n9148), .A2(n6552), .ZN(n9476) );
  INV_X2 U7387 ( .A(n7711), .ZN(n8418) );
  XNOR2_X1 U7388 ( .A(n8145), .B(n8141), .ZN(n11034) );
  XNOR2_X1 U7389 ( .A(n7663), .B(P1_IR_REG_29__SCAN_IN), .ZN(n6828) );
  INV_X2 U7390 ( .A(n7658), .ZN(n7388) );
  INV_X1 U7391 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n7849) );
  INV_X2 U7392 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  NOR2_X1 U7393 ( .A1(P3_IR_REG_12__SCAN_IN), .A2(P3_IR_REG_14__SCAN_IN), .ZN(
        n8513) );
  OR2_X1 U7394 ( .A1(n9619), .A2(n14809), .ZN(n9624) );
  OR2_X1 U7395 ( .A1(n9619), .A2(n14804), .ZN(n8507) );
  OAI21_X1 U7396 ( .B1(n14081), .B2(n14755), .A(n14087), .ZN(n8503) );
  AND2_X1 U7397 ( .A1(n8484), .A2(n8483), .ZN(n14099) );
  NOR2_X1 U7398 ( .A1(n12580), .A2(n12579), .ZN(n12587) );
  OR2_X1 U7399 ( .A1(n9127), .A2(n15206), .ZN(n9114) );
  OR2_X1 U7400 ( .A1(n9127), .A2(n9126), .ZN(n9134) );
  AND2_X1 U7401 ( .A1(n6692), .A2(n13081), .ZN(n13145) );
  NOR2_X1 U7402 ( .A1(n6700), .A2(n8167), .ZN(n6699) );
  NAND2_X1 U7403 ( .A1(n9064), .A2(n9063), .ZN(n12379) );
  NAND2_X1 U7404 ( .A1(n13857), .A2(n13856), .ZN(n13855) );
  AND2_X1 U7405 ( .A1(n14073), .A2(n8154), .ZN(n12593) );
  NAND2_X1 U7406 ( .A1(n8401), .A2(n8400), .ZN(n14291) );
  CLKBUF_X1 U7407 ( .A(n12160), .Z(n8417) );
  OR2_X1 U7408 ( .A1(n14432), .A2(n7711), .ZN(n8401) );
  NAND2_X1 U7409 ( .A1(n8413), .A2(n8399), .ZN(n14432) );
  NAND2_X1 U7410 ( .A1(n12688), .A2(n12985), .ZN(n12687) );
  NAND2_X2 U7411 ( .A1(n8113), .A2(n8112), .ZN(n14095) );
  AND2_X1 U7412 ( .A1(n9703), .A2(n9702), .ZN(n12688) );
  OR2_X1 U7413 ( .A1(n9701), .A2(n9700), .ZN(n9702) );
  NAND2_X2 U7414 ( .A1(n8095), .A2(n8094), .ZN(n14396) );
  OAI21_X1 U7415 ( .B1(n12678), .B2(n7318), .A(n7315), .ZN(n9701) );
  NAND2_X1 U7416 ( .A1(n11862), .A2(n11861), .ZN(n11863) );
  NAND2_X1 U7417 ( .A1(n7232), .A2(n8966), .ZN(n8979) );
  AND2_X1 U7418 ( .A1(n14190), .A2(n8021), .ZN(n7514) );
  NAND2_X1 U7419 ( .A1(n8945), .A2(n8946), .ZN(n8964) );
  NAND2_X1 U7420 ( .A1(n9411), .A2(n9410), .ZN(n13708) );
  OR2_X1 U7421 ( .A1(n11781), .A2(n9683), .ZN(n9686) );
  NAND2_X1 U7422 ( .A1(n11544), .A2(n6600), .ZN(n11593) );
  AND2_X1 U7423 ( .A1(n7296), .A2(n7294), .ZN(n14706) );
  NAND2_X1 U7424 ( .A1(n6886), .A2(n6602), .ZN(n11544) );
  NAND2_X1 U7425 ( .A1(n7974), .A2(n7973), .ZN(n14350) );
  NAND2_X1 U7426 ( .A1(n9394), .A2(n9393), .ZN(n13711) );
  OAI21_X1 U7427 ( .B1(n8042), .B2(n7407), .A(n7621), .ZN(n7622) );
  NAND2_X1 U7428 ( .A1(n11156), .A2(n6604), .ZN(n6886) );
  NAND2_X1 U7429 ( .A1(n8902), .A2(n8901), .ZN(n8917) );
  NAND2_X1 U7430 ( .A1(n10964), .A2(n10963), .ZN(n11156) );
  NAND2_X1 U7431 ( .A1(n10957), .A2(n10956), .ZN(n10964) );
  INV_X1 U7432 ( .A(n7265), .ZN(n8899) );
  NAND2_X1 U7433 ( .A1(n7408), .A2(n7409), .ZN(n7940) );
  NAND2_X1 U7434 ( .A1(n9316), .A2(n9315), .ZN(n12087) );
  AND3_X1 U7435 ( .A1(n7207), .A2(n7206), .A3(n6672), .ZN(n11483) );
  OR2_X1 U7436 ( .A1(n6571), .A2(n10867), .ZN(n7207) );
  NAND2_X1 U7437 ( .A1(n9286), .A2(n9285), .ZN(n12075) );
  AOI21_X1 U7438 ( .B1(n6998), .B2(n7002), .A(n6996), .ZN(n6995) );
  NAND2_X1 U7439 ( .A1(n9260), .A2(n9259), .ZN(n12060) );
  NAND2_X1 U7440 ( .A1(n7802), .A2(n7581), .ZN(n7816) );
  AND2_X1 U7441 ( .A1(n12446), .A2(n12436), .ZN(n12437) );
  AND2_X2 U7442 ( .A1(n7340), .A2(n10359), .ZN(n13803) );
  AND2_X1 U7443 ( .A1(n12440), .A2(n12439), .ZN(n12433) );
  NAND2_X1 U7444 ( .A1(n7283), .A2(n14509), .ZN(n14511) );
  NAND2_X2 U7445 ( .A1(n10392), .A2(n15118), .ZN(n15132) );
  NAND4_X1 U7446 ( .A1(n8626), .A2(n8625), .A3(n8624), .A4(n8623), .ZN(n12742)
         );
  AND3_X1 U7447 ( .A1(n8542), .A2(n8541), .A3(n8540), .ZN(n8551) );
  AND2_X2 U7448 ( .A1(n12596), .A2(n14777), .ZN(n14281) );
  BUF_X2 U7449 ( .A(n9017), .Z(n12362) );
  NAND2_X1 U7450 ( .A1(n9205), .A2(n9204), .ZN(n12025) );
  INV_X2 U7451 ( .A(n10218), .ZN(n13209) );
  INV_X2 U7452 ( .A(n8602), .ZN(n8861) );
  XNOR2_X1 U7453 ( .A(n14501), .B(P1_ADDR_REG_5__SCAN_IN), .ZN(n14502) );
  NAND2_X1 U7454 ( .A1(n7741), .A2(n7567), .ZN(n7569) );
  OR2_X1 U7455 ( .A1(n10352), .A2(n14792), .ZN(n7689) );
  NAND2_X1 U7456 ( .A1(n9024), .A2(n6572), .ZN(n12416) );
  AND2_X1 U7457 ( .A1(n8530), .A2(n8528), .ZN(n8637) );
  AND2_X1 U7458 ( .A1(n12591), .A2(n8529), .ZN(n8601) );
  INV_X4 U7459 ( .A(n11149), .ZN(n8150) );
  AND3_X2 U7460 ( .A1(n7677), .A2(n7678), .A3(n7504), .ZN(n10352) );
  AND3_X1 U7461 ( .A1(n7694), .A2(n7693), .A3(n6830), .ZN(n14763) );
  OR2_X1 U7462 ( .A1(n14485), .A2(P1_ADDR_REG_4__SCAN_IN), .ZN(n7277) );
  INV_X2 U7463 ( .A(n12293), .ZN(n12153) );
  MUX2_X1 U7464 ( .A(P1_IR_REG_0__SCAN_IN), .B(n14440), .S(n7716), .Z(n14780)
         );
  INV_X1 U7465 ( .A(n12608), .ZN(n8157) );
  NAND2_X2 U7466 ( .A1(n11997), .A2(n12000), .ZN(n12293) );
  AOI21_X1 U7467 ( .B1(n7749), .B2(n7382), .A(n7381), .ZN(n7380) );
  NAND2_X1 U7468 ( .A1(n8535), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7009) );
  OR2_X1 U7469 ( .A1(n8526), .A2(n13195), .ZN(n8527) );
  INV_X2 U7470 ( .A(n14425), .ZN(n12610) );
  AND2_X1 U7471 ( .A1(n14497), .A2(n14496), .ZN(n15528) );
  NAND2_X1 U7472 ( .A1(n8146), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8144) );
  INV_X2 U7473 ( .A(n13775), .ZN(n6551) );
  NAND2_X2 U7474 ( .A1(n8538), .A2(P3_U3151), .ZN(n13217) );
  NAND2_X2 U7475 ( .A1(n7502), .A2(n6828), .ZN(n8115) );
  OAI21_X1 U7476 ( .B1(n8146), .B2(P1_IR_REG_21__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8148) );
  OAI21_X1 U7477 ( .B1(n7566), .B2(SI_4_), .A(n7568), .ZN(n7740) );
  NAND2_X1 U7478 ( .A1(n7566), .A2(SI_4_), .ZN(n7568) );
  NAND2_X2 U7479 ( .A1(n9769), .A2(P3_U3151), .ZN(n13213) );
  AOI21_X1 U7480 ( .B1(n9907), .B2(n14494), .A(n14552), .ZN(n14496) );
  OAI21_X1 U7481 ( .B1(n7602), .B2(n9757), .A(n6710), .ZN(n7562) );
  XNOR2_X1 U7482 ( .A(n9517), .B(P2_IR_REG_22__SCAN_IN), .ZN(n9578) );
  NOR2_X1 U7483 ( .A1(n14443), .A2(n7278), .ZN(n14445) );
  XNOR2_X1 U7484 ( .A(n7662), .B(P1_IR_REG_30__SCAN_IN), .ZN(n7664) );
  MUX2_X1 U7485 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8206), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n8208) );
  NAND2_X1 U7486 ( .A1(n14427), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7662) );
  NAND2_X1 U7487 ( .A1(n7066), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7663) );
  OAI21_X1 U7488 ( .B1(n9518), .B2(P2_IR_REG_21__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9517) );
  NOR2_X1 U7489 ( .A1(n14487), .A2(n14488), .ZN(n14443) );
  NAND2_X1 U7490 ( .A1(n6880), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6882) );
  NAND2_X1 U7491 ( .A1(n7076), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7075) );
  AND3_X1 U7492 ( .A1(n6580), .A2(n7541), .A3(n7472), .ZN(n7474) );
  NOR2_X1 U7493 ( .A1(n7475), .A2(P2_IR_REG_29__SCAN_IN), .ZN(n7472) );
  INV_X1 U7494 ( .A(n8514), .ZN(n7445) );
  AND3_X2 U7495 ( .A1(n9311), .A2(n9201), .A3(n9140), .ZN(n9144) );
  AND2_X1 U7496 ( .A1(n15479), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n8560) );
  NAND2_X1 U7497 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n8965), .ZN(n8966) );
  AND4_X1 U7498 ( .A1(n8518), .A2(n8517), .A3(n8516), .A4(n8515), .ZN(n8519)
         );
  AND3_X1 U7499 ( .A1(n9139), .A2(n9138), .A3(n9180), .ZN(n9201) );
  XNOR2_X1 U7500 ( .A(n15386), .B(P1_ADDR_REG_1__SCAN_IN), .ZN(n14489) );
  NAND4_X1 U7501 ( .A1(n8513), .A2(n15498), .A3(n8744), .A4(n8709), .ZN(n8514)
         );
  AND2_X1 U7502 ( .A1(n14444), .A2(P3_ADDR_REG_2__SCAN_IN), .ZN(n7278) );
  NOR2_X1 U7503 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n7642) );
  NOR2_X1 U7504 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n6834) );
  NOR2_X1 U7505 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n6833) );
  NOR2_X1 U7506 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n6835) );
  INV_X1 U7507 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n8216) );
  NOR2_X1 U7508 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n7643) );
  INV_X1 U7509 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n9589) );
  INV_X1 U7510 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n15479) );
  NOR2_X1 U7511 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n9136) );
  NOR2_X1 U7512 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n9135) );
  INV_X1 U7513 ( .A(P2_RD_REG_SCAN_IN), .ZN(n15481) );
  INV_X1 U7514 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n9600) );
  INV_X1 U7515 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n13415) );
  NOR2_X1 U7516 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n9515) );
  INV_X1 U7517 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n15027) );
  INV_X1 U7518 ( .A(P3_ADDR_REG_1__SCAN_IN), .ZN(n15386) );
  NOR2_X2 U7519 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .ZN(
        n10204) );
  INV_X4 U7520 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  NOR2_X1 U7521 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n9138) );
  INV_X1 U7522 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n9180) );
  INV_X1 U7523 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n15498) );
  NOR2_X1 U7524 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n9139) );
  XNOR2_X1 U7525 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n8559) );
  INV_X1 U7526 ( .A(P3_IR_REG_8__SCAN_IN), .ZN(n15350) );
  NOR2_X1 U7527 ( .A1(P3_IR_REG_7__SCAN_IN), .A2(P3_IR_REG_9__SCAN_IN), .ZN(
        n8508) );
  NOR2_X1 U7528 ( .A1(P3_IR_REG_4__SCAN_IN), .A2(P3_IR_REG_3__SCAN_IN), .ZN(
        n8509) );
  BUF_X2 U7529 ( .A(P3_IR_REG_0__SCAN_IN), .Z(n15507) );
  INV_X1 U7530 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n8744) );
  AND2_X1 U7531 ( .A1(n14525), .A2(n14524), .ZN(n14692) );
  OR2_X1 U7532 ( .A1(n14525), .A2(n14524), .ZN(n6697) );
  NAND2_X2 U7533 ( .A1(n13864), .A2(n11946), .ZN(n13789) );
  INV_X1 U7534 ( .A(n7727), .ZN(n6553) );
  OAI21_X2 U7535 ( .B1(n11794), .B2(n12492), .A(n12496), .ZN(n13072) );
  NAND2_X2 U7536 ( .A1(n7716), .A2(n9769), .ZN(n7711) );
  OAI222_X1 U7537 ( .A1(n6551), .A2(n14432), .B1(P2_U3088), .B2(n12612), .C1(
        n12611), .C2(n13780), .ZN(P2_U3297) );
  XNOR2_X2 U7538 ( .A(n9147), .B(n13767), .ZN(n12612) );
  NOR2_X1 U7539 ( .A1(n9442), .A2(n7162), .ZN(n7161) );
  INV_X1 U7540 ( .A(n9431), .ZN(n7162) );
  NAND2_X1 U7541 ( .A1(n10036), .A2(n10035), .ZN(n11940) );
  NAND2_X1 U7542 ( .A1(n8454), .A2(n8376), .ZN(n8457) );
  NAND2_X1 U7543 ( .A1(n8199), .A2(n8127), .ZN(n8449) );
  OR2_X1 U7544 ( .A1(n14085), .A2(n8128), .ZN(n8127) );
  NAND2_X1 U7545 ( .A1(n7570), .A2(SI_5_), .ZN(n7572) );
  BUF_X1 U7546 ( .A(n9177), .Z(n6790) );
  INV_X4 U7547 ( .A(n6790), .ZN(n12168) );
  NOR2_X1 U7548 ( .A1(n8295), .A2(n8298), .ZN(n7060) );
  NAND2_X1 U7549 ( .A1(n8295), .A2(n8298), .ZN(n7059) );
  INV_X1 U7550 ( .A(n8354), .ZN(n6817) );
  OAI21_X1 U7551 ( .B1(n8346), .B2(n8345), .A(n8344), .ZN(n8348) );
  NOR2_X1 U7552 ( .A1(n6815), .A2(n6817), .ZN(n6816) );
  NAND2_X1 U7553 ( .A1(n6815), .A2(n6817), .ZN(n6814) );
  INV_X1 U7554 ( .A(n8357), .ZN(n6809) );
  INV_X1 U7555 ( .A(n12146), .ZN(n7497) );
  OAI22_X1 U7556 ( .A1(n8364), .A2(n6837), .B1(n6836), .B2(n8365), .ZN(n7033)
         );
  INV_X1 U7557 ( .A(n8363), .ZN(n6836) );
  NOR2_X1 U7558 ( .A1(n8366), .A2(n8363), .ZN(n6837) );
  NOR2_X1 U7559 ( .A1(n7616), .A2(n7419), .ZN(n7418) );
  INV_X1 U7560 ( .A(n7609), .ZN(n7419) );
  OR2_X1 U7561 ( .A1(n12742), .A2(n15178), .ZN(n12447) );
  AND2_X1 U7562 ( .A1(n12149), .A2(n12150), .ZN(n12152) );
  AOI21_X1 U7563 ( .B1(n7156), .B2(n6788), .A(n6608), .ZN(n6787) );
  INV_X1 U7564 ( .A(n7159), .ZN(n6788) );
  OR2_X1 U7565 ( .A1(n7788), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n7853) );
  AOI21_X1 U7566 ( .B1(n6847), .B2(n6846), .A(n6857), .ZN(n6845) );
  INV_X1 U7567 ( .A(n6851), .ZN(n6846) );
  NAND2_X1 U7568 ( .A1(n6868), .A2(n6867), .ZN(n6866) );
  INV_X1 U7569 ( .A(n11255), .ZN(n6867) );
  NOR2_X1 U7570 ( .A1(n8915), .A2(n7440), .ZN(n7439) );
  INV_X1 U7571 ( .A(n8896), .ZN(n7440) );
  INV_X1 U7572 ( .A(n12960), .ZN(n12953) );
  NAND2_X1 U7573 ( .A1(n8897), .A2(n7439), .ZN(n7438) );
  OR2_X1 U7574 ( .A1(n12686), .A2(n12985), .ZN(n12410) );
  AND2_X1 U7575 ( .A1(n13175), .A2(n12995), .ZN(n12523) );
  INV_X1 U7576 ( .A(n8773), .ZN(n7431) );
  AND2_X1 U7577 ( .A1(n12473), .A2(n12479), .ZN(n12476) );
  OR2_X1 U7578 ( .A1(n12741), .A2(n15183), .ZN(n12454) );
  NAND2_X1 U7579 ( .A1(n6841), .A2(n6624), .ZN(n9076) );
  INV_X1 U7580 ( .A(n9078), .ZN(n6841) );
  NOR2_X1 U7581 ( .A1(n8694), .A2(n7261), .ZN(n7260) );
  AND2_X1 U7582 ( .A1(n9840), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n8694) );
  INV_X1 U7583 ( .A(n8682), .ZN(n7261) );
  INV_X1 U7584 ( .A(n11874), .ZN(n7136) );
  AND2_X1 U7585 ( .A1(n12234), .A2(n12191), .ZN(n12192) );
  NOR2_X1 U7586 ( .A1(n13287), .A2(n6977), .ZN(n6976) );
  INV_X1 U7587 ( .A(n6978), .ZN(n6977) );
  XNOR2_X1 U7588 ( .A(n13373), .B(n12016), .ZN(n12248) );
  OAI21_X1 U7589 ( .B1(n9796), .B2(n6790), .A(n9216), .ZN(n14964) );
  XNOR2_X1 U7590 ( .A(n6906), .B(n8150), .ZN(n10356) );
  OAI21_X1 U7591 ( .B1(n14792), .B2(n11940), .A(n10353), .ZN(n6906) );
  NAND2_X1 U7592 ( .A1(n6547), .A2(n10823), .ZN(n10354) );
  MUX2_X1 U7593 ( .A(n8402), .B(n14291), .S(n8376), .Z(n8409) );
  XNOR2_X1 U7594 ( .A(n8454), .B(n8428), .ZN(n8468) );
  NAND2_X1 U7595 ( .A1(n7664), .A2(n6828), .ZN(n7703) );
  AND2_X1 U7596 ( .A1(n8197), .A2(n8089), .ZN(n8446) );
  NAND2_X1 U7597 ( .A1(n7222), .A2(n6930), .ZN(n6929) );
  INV_X1 U7598 ( .A(n7224), .ZN(n6930) );
  INV_X1 U7599 ( .A(n8182), .ZN(n7226) );
  OR2_X1 U7600 ( .A1(n14680), .A2(n13906), .ZN(n8314) );
  INV_X1 U7601 ( .A(n9443), .ZN(n7407) );
  OAI21_X1 U7602 ( .B1(n7958), .B2(n7607), .A(n7609), .ZN(n7986) );
  AOI21_X1 U7603 ( .B1(n7412), .B2(n7414), .A(n7410), .ZN(n7409) );
  INV_X1 U7604 ( .A(n7413), .ZN(n7412) );
  XNOR2_X1 U7605 ( .A(n7914), .B(SI_14_), .ZN(n7913) );
  OAI21_X1 U7606 ( .B1(n7562), .B2(SI_3_), .A(n7564), .ZN(n7729) );
  OAI21_X1 U7607 ( .B1(n7658), .B2(n6713), .A(n6712), .ZN(n7557) );
  NAND2_X1 U7608 ( .A1(n7658), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n6712) );
  NAND2_X1 U7609 ( .A1(n7385), .A2(n7679), .ZN(n7384) );
  NOR2_X1 U7610 ( .A1(n12573), .A2(n12378), .ZN(n7263) );
  NAND2_X1 U7611 ( .A1(n12379), .A2(n12569), .ZN(n7007) );
  OR2_X1 U7612 ( .A1(n12913), .A2(n12657), .ZN(n8977) );
  NAND2_X1 U7613 ( .A1(n6984), .A2(n6983), .ZN(n12901) );
  AOI21_X1 U7614 ( .B1(n6985), .B2(n6986), .A(n12899), .ZN(n6983) );
  XNOR2_X1 U7615 ( .A(n12548), .B(n12905), .ZN(n12923) );
  NAND2_X1 U7616 ( .A1(n7438), .A2(n7436), .ZN(n12917) );
  XNOR2_X1 U7617 ( .A(n13000), .B(n13009), .ZN(n13004) );
  NOR2_X1 U7618 ( .A1(n13013), .A2(n7451), .ZN(n7450) );
  INV_X1 U7619 ( .A(n8849), .ZN(n7451) );
  NOR2_X1 U7620 ( .A1(n13029), .A2(n12520), .ZN(n7006) );
  NAND2_X1 U7621 ( .A1(n11207), .A2(n12389), .ZN(n7005) );
  INV_X1 U7622 ( .A(n15143), .ZN(n13064) );
  AND2_X1 U7623 ( .A1(n15312), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n7272) );
  NAND2_X1 U7624 ( .A1(n7333), .A2(n7332), .ZN(n9028) );
  AND2_X1 U7625 ( .A1(n8839), .A2(n8856), .ZN(n7332) );
  INV_X1 U7626 ( .A(n8838), .ZN(n7333) );
  NAND2_X1 U7627 ( .A1(n7255), .A2(n7251), .ZN(n8723) );
  INV_X1 U7628 ( .A(n7252), .ZN(n7251) );
  OAI21_X1 U7629 ( .B1(n7254), .B2(n7253), .A(n8703), .ZN(n7252) );
  OAI21_X1 U7630 ( .B1(n7238), .B2(n6557), .A(n8612), .ZN(n7235) );
  NAND2_X1 U7631 ( .A1(n7240), .A2(n6557), .ZN(n7239) );
  NAND2_X1 U7632 ( .A1(n10930), .A2(n10931), .ZN(n10993) );
  XNOR2_X1 U7633 ( .A(n12060), .B(n13236), .ZN(n10777) );
  NAND2_X1 U7634 ( .A1(n10777), .A2(n10778), .ZN(n10935) );
  AND2_X1 U7635 ( .A1(n13250), .A2(n13251), .ZN(n6702) );
  INV_X1 U7636 ( .A(n6911), .ZN(n13398) );
  OAI21_X1 U7637 ( .B1(n9573), .B2(n7096), .A(n7095), .ZN(n9577) );
  INV_X1 U7638 ( .A(n7097), .ZN(n7096) );
  AOI21_X1 U7639 ( .B1(n7097), .B2(n7101), .A(n6563), .ZN(n7095) );
  NAND2_X1 U7640 ( .A1(n7077), .A2(n7079), .ZN(n13560) );
  AOI21_X1 U7641 ( .B1(n7080), .B2(n7083), .A(n12275), .ZN(n7079) );
  NOR2_X1 U7642 ( .A1(n13571), .A2(n13690), .ZN(n13555) );
  AND2_X1 U7643 ( .A1(n11264), .A2(n9309), .ZN(n11306) );
  NAND2_X1 U7644 ( .A1(n9282), .A2(n9281), .ZN(n11005) );
  NAND2_X1 U7645 ( .A1(n10982), .A2(n12256), .ZN(n7091) );
  AND2_X1 U7646 ( .A1(n9535), .A2(n9534), .ZN(n13450) );
  NAND2_X1 U7647 ( .A1(n6795), .A2(n6793), .ZN(n9535) );
  AOI21_X1 U7648 ( .B1(n6796), .B2(n7185), .A(n13600), .ZN(n6795) );
  CLKBUF_X1 U7649 ( .A(n9403), .Z(n9502) );
  NAND2_X1 U7650 ( .A1(n9354), .A2(n9353), .ZN(n12110) );
  NAND2_X1 U7651 ( .A1(n9841), .A2(n9769), .ZN(n9403) );
  NAND2_X1 U7652 ( .A1(n9841), .A2(n8538), .ZN(n9177) );
  AND2_X1 U7653 ( .A1(n13624), .A2(n14970), .ZN(n13730) );
  OR2_X1 U7654 ( .A1(n10360), .A2(n8150), .ZN(n10361) );
  NAND2_X1 U7655 ( .A1(n7889), .A2(n7888), .ZN(n11736) );
  AOI211_X1 U7656 ( .C1(n8459), .C2(n14068), .A(n8455), .B(n8426), .ZN(n8427)
         );
  AND2_X1 U7657 ( .A1(n6585), .A2(n8449), .ZN(n7517) );
  NAND2_X1 U7658 ( .A1(n8481), .A2(n8480), .ZN(n8482) );
  OR2_X1 U7659 ( .A1(n8478), .A2(n14755), .ZN(n8481) );
  NAND2_X1 U7660 ( .A1(n7021), .A2(n7020), .ZN(n8494) );
  INV_X1 U7661 ( .A(n14095), .ZN(n7020) );
  NAND2_X1 U7662 ( .A1(n14211), .A2(n7022), .ZN(n14146) );
  NOR2_X1 U7663 ( .A1(n14148), .A2(n7023), .ZN(n7022) );
  INV_X1 U7664 ( .A(n7024), .ZN(n7023) );
  INV_X1 U7665 ( .A(n8011), .ZN(n7516) );
  NAND2_X1 U7666 ( .A1(n8187), .A2(n6945), .ZN(n6944) );
  NOR2_X1 U7667 ( .A1(n7229), .A2(n6946), .ZN(n6945) );
  INV_X1 U7668 ( .A(n8186), .ZN(n6946) );
  NAND2_X1 U7669 ( .A1(n14264), .A2(n14272), .ZN(n14265) );
  INV_X1 U7670 ( .A(n7525), .ZN(n7524) );
  OAI21_X1 U7671 ( .B1(n7937), .B2(n7526), .A(n7955), .ZN(n7525) );
  AND2_X1 U7672 ( .A1(n11351), .A2(n7225), .ZN(n7224) );
  OR2_X1 U7673 ( .A1(n11464), .A2(n7226), .ZN(n7225) );
  NAND2_X1 U7674 ( .A1(n7822), .A2(n7821), .ZN(n11232) );
  AND2_X1 U7675 ( .A1(n8439), .A2(n8175), .ZN(n7227) );
  NAND2_X1 U7676 ( .A1(n7716), .A2(n8538), .ZN(n7727) );
  INV_X1 U7677 ( .A(n14085), .ZN(n9620) );
  CLKBUF_X1 U7678 ( .A(n7727), .Z(n8419) );
  INV_X1 U7679 ( .A(n14783), .ZN(n14761) );
  INV_X1 U7680 ( .A(n7638), .ZN(n7636) );
  XNOR2_X1 U7681 ( .A(n8111), .B(n8110), .ZN(n11872) );
  NAND2_X1 U7682 ( .A1(n7402), .A2(n7403), .ZN(n8111) );
  XNOR2_X1 U7683 ( .A(n7622), .B(n7623), .ZN(n8052) );
  XNOR2_X1 U7684 ( .A(n7620), .B(SI_22_), .ZN(n8042) );
  AOI21_X1 U7685 ( .B1(n7380), .B2(n7571), .A(n7574), .ZN(n7379) );
  OAI21_X1 U7686 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(n14462), .A(n14461), .ZN(
        n14482) );
  AND2_X1 U7687 ( .A1(n8976), .A2(n8975), .ZN(n12926) );
  AOI21_X1 U7688 ( .B1(n8258), .B2(n8257), .A(n10300), .ZN(n6679) );
  NOR2_X1 U7689 ( .A1(n7464), .A2(n7463), .ZN(n7462) );
  OR2_X1 U7690 ( .A1(n12022), .A2(n12023), .ZN(n7461) );
  NAND2_X1 U7691 ( .A1(n6615), .A2(n7467), .ZN(n7466) );
  INV_X1 U7692 ( .A(n8277), .ZN(n6801) );
  INV_X1 U7693 ( .A(n12069), .ZN(n7483) );
  NAND2_X1 U7694 ( .A1(n12063), .A2(n7487), .ZN(n7486) );
  INV_X1 U7695 ( .A(n12064), .ZN(n7487) );
  NAND2_X1 U7696 ( .A1(n6825), .A2(n8292), .ZN(n6824) );
  INV_X1 U7697 ( .A(n8293), .ZN(n6825) );
  NOR2_X1 U7698 ( .A1(n7060), .A2(n6822), .ZN(n6821) );
  INV_X1 U7699 ( .A(n6824), .ZN(n6822) );
  INV_X1 U7700 ( .A(n7059), .ZN(n6819) );
  AND2_X1 U7701 ( .A1(n6827), .A2(n8293), .ZN(n6826) );
  INV_X1 U7702 ( .A(n8292), .ZN(n6827) );
  NAND2_X1 U7703 ( .A1(n12084), .A2(n6775), .ZN(n7460) );
  NAND2_X1 U7704 ( .A1(n7479), .A2(n7477), .ZN(n12084) );
  AOI21_X1 U7705 ( .B1(n7478), .B2(n12083), .A(n12082), .ZN(n7477) );
  AOI21_X1 U7706 ( .B1(n7060), .B2(n7059), .A(n7057), .ZN(n7056) );
  INV_X1 U7707 ( .A(n12088), .ZN(n7458) );
  NAND2_X1 U7708 ( .A1(n6816), .A2(n6814), .ZN(n6813) );
  INV_X1 U7709 ( .A(n6814), .ZN(n6810) );
  OAI22_X1 U7710 ( .A1(n8350), .A2(n7051), .B1(n8351), .B2(n7050), .ZN(n8356)
         );
  INV_X1 U7711 ( .A(n8349), .ZN(n7050) );
  NOR2_X1 U7712 ( .A1(n8352), .A2(n8349), .ZN(n7051) );
  NAND2_X1 U7713 ( .A1(n12135), .A2(n6641), .ZN(n6748) );
  AND2_X1 U7714 ( .A1(n6751), .A2(n6750), .ZN(n6749) );
  NAND2_X1 U7715 ( .A1(n12144), .A2(n12145), .ZN(n7500) );
  NAND2_X1 U7716 ( .A1(n7501), .A2(n12147), .ZN(n7499) );
  INV_X1 U7717 ( .A(n12679), .ZN(n7317) );
  NAND2_X1 U7718 ( .A1(n9076), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n6840) );
  INV_X1 U7719 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n7449) );
  NOR2_X1 U7720 ( .A1(n13287), .A2(n7188), .ZN(n7187) );
  INV_X1 U7721 ( .A(n7167), .ZN(n6786) );
  AND2_X1 U7722 ( .A1(n13509), .A2(n7171), .ZN(n7170) );
  NAND2_X1 U7723 ( .A1(n7172), .A2(n9462), .ZN(n7171) );
  NOR2_X1 U7724 ( .A1(n13661), .A2(n13670), .ZN(n6978) );
  INV_X1 U7725 ( .A(n9540), .ZN(n7069) );
  NAND2_X1 U7726 ( .A1(n7029), .A2(n8370), .ZN(n7028) );
  INV_X1 U7727 ( .A(n7596), .ZN(n7414) );
  INV_X1 U7728 ( .A(n7846), .ZN(n7391) );
  NOR2_X1 U7729 ( .A1(n7586), .A2(n7396), .ZN(n7395) );
  INV_X1 U7730 ( .A(n7584), .ZN(n7396) );
  INV_X1 U7731 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n7553) );
  INV_X1 U7732 ( .A(P1_RD_REG_SCAN_IN), .ZN(n7374) );
  INV_X1 U7733 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n14446) );
  NOR2_X1 U7734 ( .A1(n11513), .A2(n11518), .ZN(n7327) );
  INV_X1 U7735 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n15485) );
  INV_X1 U7736 ( .A(n8529), .ZN(n8528) );
  NAND2_X1 U7737 ( .A1(n10897), .A2(n15083), .ZN(n6742) );
  OAI21_X1 U7738 ( .B1(n6741), .B2(n15087), .A(n6739), .ZN(n10898) );
  AOI21_X1 U7739 ( .B1(n6742), .B2(n6740), .A(n12350), .ZN(n6739) );
  INV_X1 U7740 ( .A(n12314), .ZN(n6849) );
  NAND2_X1 U7741 ( .A1(n12317), .A2(n6744), .ZN(n10904) );
  OR2_X1 U7742 ( .A1(n10903), .A2(n15217), .ZN(n6744) );
  NAND2_X1 U7743 ( .A1(n11248), .A2(n6667), .ZN(n11490) );
  NAND2_X1 U7744 ( .A1(n12559), .A2(n12879), .ZN(n12382) );
  OR2_X1 U7745 ( .A1(n12913), .A2(n12926), .ZN(n12554) );
  INV_X1 U7746 ( .A(n13159), .ZN(n9057) );
  NOR2_X1 U7747 ( .A1(n12953), .A2(n7437), .ZN(n7436) );
  INV_X1 U7748 ( .A(n8914), .ZN(n7437) );
  OR2_X1 U7749 ( .A1(n13122), .A2(n13037), .ZN(n12513) );
  OAI21_X1 U7750 ( .B1(n7432), .B2(n7431), .A(n8791), .ZN(n7430) );
  NOR2_X1 U7751 ( .A1(n9050), .A2(n7433), .ZN(n7432) );
  INV_X1 U7752 ( .A(n8755), .ZN(n7433) );
  INV_X1 U7753 ( .A(n8702), .ZN(n7425) );
  NOR2_X1 U7754 ( .A1(n6576), .A2(n7422), .ZN(n7421) );
  INV_X1 U7755 ( .A(n12471), .ZN(n7422) );
  OR2_X1 U7756 ( .A1(n15121), .A2(n8551), .ZN(n12422) );
  INV_X1 U7757 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n9084) );
  NAND2_X1 U7758 ( .A1(n6624), .A2(n8522), .ZN(n7448) );
  INV_X1 U7759 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n8520) );
  INV_X1 U7760 ( .A(n9080), .ZN(n6981) );
  NAND2_X1 U7761 ( .A1(n8667), .A2(n8666), .ZN(n8681) );
  NAND2_X1 U7762 ( .A1(n9794), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n8666) );
  NAND2_X1 U7763 ( .A1(n7241), .A2(n8588), .ZN(n7238) );
  NAND2_X1 U7764 ( .A1(n10204), .A2(n15485), .ZN(n8586) );
  XNOR2_X1 U7765 ( .A(n12068), .B(n13236), .ZN(n10930) );
  XNOR2_X1 U7766 ( .A(n14964), .B(n13236), .ZN(n10430) );
  NOR2_X1 U7767 ( .A1(n6767), .A2(n12159), .ZN(n6766) );
  NOR2_X1 U7768 ( .A1(n12156), .A2(n12157), .ZN(n6761) );
  NAND2_X1 U7769 ( .A1(n12159), .A2(n6767), .ZN(n6765) );
  NOR2_X1 U7770 ( .A1(n12231), .A2(n12186), .ZN(n12234) );
  NAND2_X1 U7771 ( .A1(n7406), .A2(n6665), .ZN(n12291) );
  NAND2_X1 U7772 ( .A1(n7149), .A2(n9375), .ZN(n7148) );
  AND2_X1 U7773 ( .A1(n9388), .A2(n7150), .ZN(n7149) );
  AOI21_X1 U7774 ( .B1(n7167), .B2(n7168), .A(n7166), .ZN(n7165) );
  INV_X1 U7775 ( .A(n13493), .ZN(n7166) );
  AOI21_X1 U7776 ( .B1(n7161), .B2(n13584), .A(n6595), .ZN(n7159) );
  NOR2_X1 U7777 ( .A1(n6971), .A2(n13708), .ZN(n6970) );
  INV_X1 U7778 ( .A(n6972), .ZN(n6971) );
  NAND2_X1 U7779 ( .A1(n11846), .A2(n9386), .ZN(n7176) );
  AND2_X1 U7780 ( .A1(n6783), .A2(n11430), .ZN(n6782) );
  OR2_X1 U7781 ( .A1(n12105), .A2(n9334), .ZN(n6783) );
  INV_X1 U7782 ( .A(n6782), .ZN(n6781) );
  OR2_X1 U7783 ( .A1(n9578), .A2(n10529), .ZN(n10019) );
  OAI21_X1 U7784 ( .B1(n13585), .B2(n6789), .A(n6787), .ZN(n13531) );
  INV_X1 U7785 ( .A(n13755), .ZN(n13574) );
  OR2_X1 U7786 ( .A1(n11268), .A2(n12081), .ZN(n11310) );
  NAND2_X1 U7787 ( .A1(n9185), .A2(n9184), .ZN(n7152) );
  AND2_X1 U7788 ( .A1(n7541), .A2(n6580), .ZN(n7473) );
  INV_X1 U7789 ( .A(n9226), .ZN(n9239) );
  XNOR2_X1 U7790 ( .A(n10366), .B(n8150), .ZN(n10367) );
  AND2_X1 U7791 ( .A1(n7364), .A2(n13824), .ZN(n7363) );
  NAND2_X1 U7792 ( .A1(n13849), .A2(n11959), .ZN(n7364) );
  NAND2_X1 U7793 ( .A1(n6905), .A2(n11959), .ZN(n6903) );
  NAND2_X1 U7794 ( .A1(n6707), .A2(n6706), .ZN(n6884) );
  INV_X1 U7795 ( .A(n13912), .ZN(n6706) );
  INV_X1 U7796 ( .A(n13910), .ZN(n6707) );
  NAND2_X1 U7797 ( .A1(n7664), .A2(n14435), .ZN(n7723) );
  AOI21_X1 U7798 ( .B1(n14104), .B2(n6967), .A(n6966), .ZN(n6965) );
  INV_X1 U7799 ( .A(n8197), .ZN(n6967) );
  INV_X1 U7800 ( .A(n8479), .ZN(n6966) );
  NAND2_X1 U7801 ( .A1(n6965), .A2(n14100), .ZN(n6964) );
  AOI21_X1 U7802 ( .B1(n7524), .B2(n7522), .A(n7521), .ZN(n7520) );
  INV_X1 U7803 ( .A(n8325), .ZN(n7521) );
  AOI21_X1 U7804 ( .B1(n7228), .B2(n11753), .A(n6609), .ZN(n6937) );
  NAND2_X1 U7805 ( .A1(n11282), .A2(n11608), .ZN(n11355) );
  NAND2_X1 U7806 ( .A1(n8173), .A2(n7747), .ZN(n8437) );
  NAND2_X1 U7807 ( .A1(n7718), .A2(n8171), .ZN(n8168) );
  NOR2_X1 U7808 ( .A1(n6829), .A2(n14435), .ZN(n6831) );
  OR2_X1 U7809 ( .A1(n7664), .A2(n7691), .ZN(n6829) );
  NOR2_X1 U7810 ( .A1(n7703), .A2(n7690), .ZN(n6832) );
  NAND2_X1 U7811 ( .A1(n8107), .A2(n7519), .ZN(n7518) );
  AND2_X1 U7812 ( .A1(n8448), .A2(n8106), .ZN(n7519) );
  NAND2_X1 U7813 ( .A1(n14211), .A2(n14329), .ZN(n14196) );
  NAND2_X1 U7814 ( .A1(n7011), .A2(n7010), .ZN(n11755) );
  INV_X1 U7815 ( .A(n14373), .ZN(n7010) );
  OR2_X1 U7816 ( .A1(n8152), .A2(n14061), .ZN(n8243) );
  NAND2_X1 U7817 ( .A1(n7622), .A2(n7623), .ZN(n7624) );
  INV_X1 U7818 ( .A(n7652), .ZN(n8201) );
  NAND2_X1 U7819 ( .A1(n7619), .A2(n7618), .ZN(n7620) );
  NAND2_X1 U7820 ( .A1(n7415), .A2(n6567), .ZN(n7619) );
  NAND2_X1 U7821 ( .A1(n7606), .A2(n7605), .ZN(n7958) );
  CLKBUF_X1 U7822 ( .A(n7959), .Z(n7923) );
  NAND2_X1 U7823 ( .A1(n7594), .A2(n7593), .ZN(n7881) );
  XNOR2_X1 U7824 ( .A(n7592), .B(SI_12_), .ZN(n7864) );
  XNOR2_X1 U7825 ( .A(n7588), .B(SI_11_), .ZN(n7846) );
  NAND2_X1 U7826 ( .A1(n7582), .A2(SI_9_), .ZN(n7584) );
  NAND2_X1 U7827 ( .A1(n7573), .A2(SI_6_), .ZN(n7575) );
  NAND2_X1 U7828 ( .A1(n7383), .A2(n7389), .ZN(n7385) );
  OAI22_X1 U7829 ( .A1(n14507), .A2(n14454), .B1(P1_ADDR_REG_6__SCAN_IN), .B2(
        n14453), .ZN(n14455) );
  OR2_X1 U7830 ( .A1(n11046), .A2(n11047), .ZN(n11044) );
  AND2_X1 U7831 ( .A1(n12695), .A2(n7305), .ZN(n7304) );
  OR2_X1 U7832 ( .A1(n12660), .A2(n7306), .ZN(n7305) );
  INV_X1 U7833 ( .A(n9688), .ZN(n7306) );
  AND2_X1 U7834 ( .A1(n9740), .A2(n9627), .ZN(n6709) );
  AND2_X1 U7835 ( .A1(n10835), .A2(n7312), .ZN(n7311) );
  NAND2_X1 U7836 ( .A1(n10650), .A2(n9651), .ZN(n7312) );
  NAND2_X1 U7837 ( .A1(n10481), .A2(n9645), .ZN(n10478) );
  NOR2_X1 U7838 ( .A1(n11642), .A2(n7338), .ZN(n7337) );
  INV_X1 U7839 ( .A(n9676), .ZN(n7338) );
  NAND2_X1 U7840 ( .A1(n12374), .A2(n7264), .ZN(n12573) );
  NAND2_X1 U7841 ( .A1(n14614), .A2(n12376), .ZN(n7264) );
  NAND2_X1 U7842 ( .A1(n7199), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n7198) );
  NAND2_X1 U7843 ( .A1(n6717), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n7196) );
  INV_X1 U7844 ( .A(n15037), .ZN(n6717) );
  XNOR2_X1 U7845 ( .A(n10897), .B(n10896), .ZN(n15087) );
  INV_X1 U7846 ( .A(n6742), .ZN(n6741) );
  NAND2_X1 U7847 ( .A1(n6854), .A2(n6858), .ZN(n6853) );
  INV_X1 U7848 ( .A(n6855), .ZN(n6854) );
  AOI21_X1 U7849 ( .B1(n12344), .B2(n6859), .A(n6856), .ZN(n6855) );
  INV_X1 U7850 ( .A(n12330), .ZN(n6856) );
  NAND2_X1 U7851 ( .A1(n12318), .A2(n12319), .ZN(n12317) );
  XNOR2_X1 U7852 ( .A(n10904), .B(n10883), .ZN(n15108) );
  NAND2_X1 U7853 ( .A1(n10906), .A2(n10907), .ZN(n11248) );
  OR2_X1 U7854 ( .A1(n11254), .A2(n11253), .ZN(n6868) );
  XNOR2_X1 U7855 ( .A(n11490), .B(n11484), .ZN(n11250) );
  INV_X1 U7856 ( .A(n6866), .ZN(n11500) );
  XNOR2_X1 U7857 ( .A(n12822), .B(n12833), .ZN(n12808) );
  OR2_X1 U7858 ( .A1(n12835), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n7201) );
  NOR2_X1 U7859 ( .A1(n12808), .A2(n12809), .ZN(n12823) );
  NAND2_X1 U7860 ( .A1(n12802), .A2(n12804), .ZN(n12818) );
  OR2_X1 U7861 ( .A1(n14603), .A2(n14602), .ZN(n14601) );
  NAND2_X1 U7862 ( .A1(n6719), .A2(n12560), .ZN(n12875) );
  INV_X1 U7863 ( .A(n12873), .ZN(n6719) );
  AND2_X1 U7864 ( .A1(n12901), .A2(n12554), .ZN(n12888) );
  NAND2_X1 U7865 ( .A1(n6577), .A2(n12542), .ZN(n6986) );
  NAND2_X1 U7866 ( .A1(n6987), .A2(n6577), .ZN(n6985) );
  OAI21_X1 U7867 ( .B1(n9059), .B2(n12543), .A(n12923), .ZN(n6987) );
  OAI21_X1 U7868 ( .B1(n8960), .B2(n8961), .A(n6623), .ZN(n7434) );
  AND2_X1 U7869 ( .A1(n12958), .A2(n12953), .ZN(n9056) );
  NAND2_X1 U7870 ( .A1(n12937), .A2(n9059), .ZN(n12941) );
  NAND2_X1 U7871 ( .A1(n7438), .A2(n8914), .ZN(n12954) );
  AND2_X1 U7872 ( .A1(n8913), .A2(n8912), .ZN(n12985) );
  OR2_X1 U7873 ( .A1(n13015), .A2(n12523), .ZN(n7008) );
  AND2_X1 U7874 ( .A1(n8868), .A2(n12518), .ZN(n13013) );
  AND3_X1 U7875 ( .A1(n8880), .A2(n8879), .A3(n8878), .ZN(n13009) );
  NAND2_X1 U7876 ( .A1(n13039), .A2(n7452), .ZN(n13020) );
  NOR2_X1 U7877 ( .A1(n13023), .A2(n7453), .ZN(n7452) );
  INV_X1 U7878 ( .A(n8829), .ZN(n7453) );
  NAND2_X1 U7879 ( .A1(n9052), .A2(n13041), .ZN(n13045) );
  OAI21_X1 U7880 ( .B1(n13051), .B2(n8812), .A(n8811), .ZN(n13036) );
  OR2_X1 U7881 ( .A1(n13036), .A2(n13041), .ZN(n13039) );
  INV_X1 U7882 ( .A(n12734), .ZN(n13068) );
  AND2_X1 U7883 ( .A1(n12502), .A2(n12508), .ZN(n13071) );
  INV_X1 U7884 ( .A(n12735), .ZN(n13054) );
  NAND2_X1 U7885 ( .A1(n8756), .A2(n7432), .ZN(n11791) );
  INV_X1 U7886 ( .A(n11441), .ZN(n13066) );
  AOI21_X1 U7887 ( .B1(n7001), .B2(n7000), .A(n6999), .ZN(n6998) );
  NAND2_X1 U7888 ( .A1(n11449), .A2(n12469), .ZN(n7426) );
  NOR2_X1 U7889 ( .A1(n6558), .A2(n12463), .ZN(n7004) );
  NAND2_X1 U7890 ( .A1(n11342), .A2(n12471), .ZN(n11449) );
  AOI21_X1 U7891 ( .B1(n6991), .B2(n6994), .A(n6989), .ZN(n6988) );
  AOI21_X1 U7892 ( .B1(n11174), .B2(n6989), .A(n8656), .ZN(n11208) );
  AND2_X1 U7893 ( .A1(n6994), .A2(n8619), .ZN(n7443) );
  OR2_X1 U7894 ( .A1(n11070), .A2(n12437), .ZN(n11072) );
  NAND2_X1 U7895 ( .A1(n11054), .A2(n12384), .ZN(n11056) );
  NAND2_X1 U7896 ( .A1(n9045), .A2(n12446), .ZN(n11054) );
  INV_X1 U7897 ( .A(n14614), .ZN(n14620) );
  NAND2_X1 U7898 ( .A1(n8820), .A2(n8819), .ZN(n13126) );
  BUF_X1 U7899 ( .A(n12363), .Z(n12370) );
  NAND2_X1 U7900 ( .A1(n12549), .A2(n12581), .ZN(n13069) );
  AND2_X1 U7901 ( .A1(n9089), .A2(n9088), .ZN(n9805) );
  NAND2_X1 U7902 ( .A1(n8997), .A2(n8998), .ZN(n7250) );
  NAND2_X1 U7903 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n8900), .ZN(n8901) );
  AND2_X1 U7904 ( .A1(n12615), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n7267) );
  NAND2_X1 U7905 ( .A1(n8757), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n7273) );
  INV_X1 U7906 ( .A(n7260), .ZN(n7259) );
  AOI21_X1 U7907 ( .B1(n7260), .B2(n7258), .A(n6619), .ZN(n7257) );
  INV_X1 U7908 ( .A(n8680), .ZN(n7258) );
  CLKBUF_X1 U7909 ( .A(n8681), .Z(n6693) );
  NAND2_X1 U7910 ( .A1(n8628), .A2(n8627), .ZN(n8649) );
  AND2_X1 U7911 ( .A1(n8633), .A2(n8646), .ZN(n10899) );
  AND2_X1 U7912 ( .A1(n10028), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n8575) );
  INV_X1 U7913 ( .A(n11659), .ZN(n7114) );
  INV_X1 U7914 ( .A(n13271), .ZN(n7137) );
  NAND2_X1 U7915 ( .A1(n7128), .A2(n6573), .ZN(n7127) );
  NOR2_X1 U7916 ( .A1(n7124), .A2(n7123), .ZN(n7122) );
  NOR2_X1 U7917 ( .A1(n7128), .A2(n6573), .ZN(n7123) );
  NOR2_X1 U7918 ( .A1(n7130), .A2(n7127), .ZN(n7124) );
  INV_X1 U7919 ( .A(n10310), .ZN(n6685) );
  OR2_X1 U7920 ( .A1(n10784), .A2(n10783), .ZN(n10936) );
  AND2_X1 U7921 ( .A1(n10938), .A2(n7139), .ZN(n7138) );
  OR2_X1 U7922 ( .A1(n9476), .A2(n9164), .ZN(n9165) );
  NOR2_X1 U7923 ( .A1(n14892), .A2(n6914), .ZN(n14909) );
  AND2_X1 U7924 ( .A1(n14900), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n6914) );
  OR2_X1 U7925 ( .A1(n14909), .A2(n14910), .ZN(n6913) );
  XNOR2_X1 U7926 ( .A(n6911), .B(n14920), .ZN(n14919) );
  OR2_X1 U7927 ( .A1(n13426), .A2(n13442), .ZN(n13424) );
  AND2_X1 U7928 ( .A1(n13443), .A2(n13442), .ZN(n13649) );
  NAND2_X1 U7929 ( .A1(n9573), .A2(n7100), .ZN(n7099) );
  OR2_X1 U7930 ( .A1(n13531), .A2(n9462), .ZN(n7169) );
  AND2_X1 U7931 ( .A1(n9441), .A2(n9440), .ZN(n13550) );
  NAND2_X1 U7932 ( .A1(n9562), .A2(n7094), .ZN(n13623) );
  AND2_X1 U7933 ( .A1(n13616), .A2(n9561), .ZN(n7094) );
  NAND2_X1 U7934 ( .A1(n11803), .A2(n9559), .ZN(n11845) );
  NOR2_X1 U7935 ( .A1(n11810), .A2(n13726), .ZN(n11848) );
  NAND2_X1 U7936 ( .A1(n11263), .A2(n9550), .ZN(n7093) );
  NAND2_X1 U7937 ( .A1(n7093), .A2(n7092), .ZN(n11302) );
  AND2_X1 U7938 ( .A1(n12263), .A2(n9551), .ZN(n7092) );
  NAND2_X1 U7939 ( .A1(n7174), .A2(n6601), .ZN(n11264) );
  NAND2_X1 U7940 ( .A1(n11005), .A2(n12260), .ZN(n7174) );
  NAND2_X1 U7941 ( .A1(n11003), .A2(n9549), .ZN(n11263) );
  OAI21_X1 U7942 ( .B1(n10716), .B2(n12060), .A(n9269), .ZN(n10918) );
  NOR2_X1 U7943 ( .A1(n7193), .A2(n7191), .ZN(n7190) );
  NOR2_X1 U7944 ( .A1(n12257), .A2(n7090), .ZN(n7089) );
  INV_X1 U7945 ( .A(n9546), .ZN(n7090) );
  OAI21_X1 U7946 ( .B1(n10659), .B2(n9224), .A(n9225), .ZN(n10844) );
  OR2_X1 U7947 ( .A1(n10844), .A2(n9543), .ZN(n10845) );
  NAND2_X1 U7948 ( .A1(n10237), .A2(n10240), .ZN(n10236) );
  NAND2_X1 U7949 ( .A1(n9537), .A2(n9536), .ZN(n7071) );
  INV_X1 U7950 ( .A(n12248), .ZN(n10078) );
  NAND2_X1 U7951 ( .A1(n7145), .A2(n12613), .ZN(n13624) );
  XNOR2_X1 U7952 ( .A(n9578), .B(n12289), .ZN(n7145) );
  OR2_X1 U7953 ( .A1(n6975), .A2(n14999), .ZN(n7538) );
  NAND2_X1 U7955 ( .A1(n9190), .A2(n9189), .ZN(n12021) );
  AND2_X1 U7956 ( .A1(n9376), .A2(n9375), .ZN(n9389) );
  AND2_X1 U7957 ( .A1(n7365), .A2(n7358), .ZN(n7357) );
  INV_X1 U7958 ( .A(n7366), .ZN(n7365) );
  NAND2_X1 U7959 ( .A1(n7361), .A2(n7359), .ZN(n7358) );
  OAI21_X1 U7960 ( .B1(n13898), .B2(n7368), .A(n7367), .ZN(n7366) );
  NAND2_X1 U7961 ( .A1(n6561), .A2(n6599), .ZN(n6885) );
  NAND2_X1 U7962 ( .A1(n13855), .A2(n7369), .ZN(n13812) );
  NOR2_X1 U7963 ( .A1(n13815), .A2(n7370), .ZN(n7369) );
  INV_X1 U7964 ( .A(n11930), .ZN(n7370) );
  NAND2_X1 U7965 ( .A1(n10041), .A2(n10360), .ZN(n10362) );
  INV_X1 U7966 ( .A(n13898), .ZN(n6895) );
  AOI21_X1 U7967 ( .B1(n6898), .B2(n6903), .A(n6897), .ZN(n6896) );
  INV_X1 U7968 ( .A(n7368), .ZN(n6897) );
  NOR2_X1 U7969 ( .A1(n8468), .A2(n8467), .ZN(n7044) );
  NAND2_X1 U7970 ( .A1(n6798), .A2(n6797), .ZN(n8411) );
  OR2_X1 U7971 ( .A1(n8381), .A2(n8382), .ZN(n6797) );
  AND2_X1 U7972 ( .A1(n8466), .A2(n7037), .ZN(n7036) );
  AND2_X1 U7973 ( .A1(n8050), .A2(n8049), .ZN(n13817) );
  INV_X1 U7974 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n14442) );
  XNOR2_X1 U7975 ( .A(n8379), .B(n13917), .ZN(n8451) );
  INV_X1 U7976 ( .A(n8449), .ZN(n8499) );
  NAND2_X1 U7977 ( .A1(n14103), .A2(n14104), .ZN(n14102) );
  NAND2_X1 U7978 ( .A1(n7213), .A2(n8446), .ZN(n14119) );
  AND2_X1 U7979 ( .A1(n6960), .A2(n14158), .ZN(n6959) );
  NAND2_X1 U7980 ( .A1(n14174), .A2(n8192), .ZN(n6960) );
  NAND2_X1 U7981 ( .A1(n8191), .A2(n8190), .ZN(n14172) );
  NAND2_X1 U7982 ( .A1(n14175), .A2(n14174), .ZN(n14173) );
  NOR2_X1 U7983 ( .A1(n14205), .A2(n6943), .ZN(n6942) );
  INV_X1 U7984 ( .A(n8342), .ZN(n6943) );
  INV_X1 U7985 ( .A(n8010), .ZN(n14224) );
  NAND2_X1 U7986 ( .A1(n11749), .A2(n8184), .ZN(n14274) );
  NAND2_X1 U7988 ( .A1(n6938), .A2(n7526), .ZN(n11749) );
  INV_X1 U7989 ( .A(n11751), .ZN(n6938) );
  AOI21_X1 U7990 ( .B1(n7224), .B2(n7226), .A(n6611), .ZN(n7222) );
  NOR2_X1 U7991 ( .A1(n11633), .A2(n6711), .ZN(n7513) );
  INV_X1 U7992 ( .A(n7898), .ZN(n6711) );
  INV_X1 U7993 ( .A(n13932), .ZN(n11550) );
  NAND2_X1 U7994 ( .A1(n6941), .A2(n8177), .ZN(n11016) );
  NAND2_X1 U7995 ( .A1(n6935), .A2(n6933), .ZN(n10592) );
  AND2_X1 U7996 ( .A1(n6934), .A2(n10594), .ZN(n6933) );
  NAND2_X1 U7997 ( .A1(n7782), .A2(n10589), .ZN(n6934) );
  NAND2_X1 U7998 ( .A1(n10295), .A2(n8172), .ZN(n10286) );
  AND2_X1 U7999 ( .A1(n10048), .A2(n8158), .ZN(n14247) );
  AND2_X1 U8000 ( .A1(n10048), .A2(n13965), .ZN(n14757) );
  NAND2_X1 U8001 ( .A1(n8166), .A2(n8165), .ZN(n8167) );
  INV_X1 U8002 ( .A(n12593), .ZN(n8166) );
  NAND2_X1 U8003 ( .A1(n8002), .A2(n8001), .ZN(n14345) );
  NAND2_X1 U8004 ( .A1(n8243), .A2(n8244), .ZN(n14783) );
  NAND2_X1 U8005 ( .A1(n8153), .A2(n6549), .ZN(n14793) );
  AOI21_X1 U8006 ( .B1(n7400), .B2(n7398), .A(n6669), .ZN(n7397) );
  INV_X1 U8007 ( .A(n7400), .ZN(n7399) );
  XNOR2_X1 U8008 ( .A(n8093), .B(n8092), .ZN(n11816) );
  XNOR2_X1 U8009 ( .A(n8029), .B(n8028), .ZN(n11134) );
  OAI22_X1 U8010 ( .A1(n7917), .A2(n7916), .B1(n7915), .B2(SI_14_), .ZN(n7920)
         );
  OR2_X1 U8011 ( .A1(n7866), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n7867) );
  INV_X1 U8012 ( .A(n7572), .ZN(n7381) );
  INV_X1 U8013 ( .A(n7568), .ZN(n7382) );
  AND2_X1 U8014 ( .A1(n7387), .A2(n7386), .ZN(n7679) );
  AOI21_X1 U8015 ( .B1(n7388), .B2(n15478), .A(n7695), .ZN(n7387) );
  INV_X1 U8016 ( .A(n7384), .ZN(n6746) );
  NAND2_X1 U8017 ( .A1(n7385), .A2(n7558), .ZN(n7681) );
  NAND2_X1 U8018 ( .A1(n14557), .A2(n14556), .ZN(n7283) );
  NAND2_X1 U8019 ( .A1(n14561), .A2(P2_ADDR_REG_10__SCAN_IN), .ZN(n7289) );
  AOI21_X1 U8020 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(n14466), .A(n14465), .ZN(
        n14527) );
  NOR2_X1 U8021 ( .A1(n14523), .A2(n14522), .ZN(n14465) );
  NAND2_X1 U8022 ( .A1(n7299), .A2(n11103), .ZN(n7298) );
  INV_X1 U8023 ( .A(n14704), .ZN(n7299) );
  NAND2_X1 U8024 ( .A1(n8886), .A2(n8885), .ZN(n12644) );
  AND2_X1 U8025 ( .A1(n8894), .A2(n8893), .ZN(n12974) );
  INV_X1 U8026 ( .A(n12737), .ZN(n11720) );
  NAND4_X1 U8027 ( .A1(n8664), .A2(n8663), .A3(n8662), .A4(n8661), .ZN(n12740)
         );
  XNOR2_X1 U8028 ( .A(n12818), .B(n12824), .ZN(n12803) );
  NAND2_X1 U8029 ( .A1(n12803), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n12819) );
  OR2_X1 U8030 ( .A1(n14579), .A2(n6736), .ZN(n6735) );
  INV_X1 U8031 ( .A(n12855), .ZN(n6736) );
  NAND2_X1 U8032 ( .A1(n6735), .A2(n6727), .ZN(n6726) );
  AOI21_X1 U8033 ( .B1(n12855), .B2(n6734), .A(n6723), .ZN(n6727) );
  NAND2_X1 U8034 ( .A1(n6737), .A2(n14593), .ZN(n6723) );
  AND2_X1 U8035 ( .A1(n6731), .A2(n6729), .ZN(n6728) );
  NAND2_X1 U8036 ( .A1(n6737), .A2(n6730), .ZN(n6729) );
  OAI21_X1 U8037 ( .B1(n12855), .B2(n6733), .A(n6724), .ZN(n6731) );
  INV_X1 U8038 ( .A(n6738), .ZN(n6730) );
  NAND2_X1 U8039 ( .A1(n6871), .A2(n6870), .ZN(n6869) );
  INV_X1 U8040 ( .A(n12869), .ZN(n6870) );
  NAND2_X1 U8041 ( .A1(n6872), .A2(n15085), .ZN(n6871) );
  OR2_X1 U8042 ( .A1(n14611), .A2(n9004), .ZN(n12883) );
  AND2_X1 U8043 ( .A1(n12920), .A2(n12919), .ZN(n12922) );
  AND2_X1 U8044 ( .A1(n8920), .A2(n8919), .ZN(n12969) );
  NAND2_X1 U8045 ( .A1(n8594), .A2(SI_23_), .ZN(n8919) );
  OR2_X1 U8046 ( .A1(n15200), .A2(n9726), .ZN(n15118) );
  AND2_X1 U8047 ( .A1(n11996), .A2(n9072), .ZN(n9127) );
  AND2_X1 U8048 ( .A1(n9110), .A2(n9109), .ZN(n15206) );
  INV_X1 U8049 ( .A(n13542), .ZN(n13686) );
  NOR2_X1 U8050 ( .A1(n7119), .A2(n13348), .ZN(n7117) );
  NOR2_X1 U8051 ( .A1(n7125), .A2(n7120), .ZN(n7119) );
  NOR2_X1 U8052 ( .A1(n7126), .A2(n6573), .ZN(n7125) );
  INV_X1 U8053 ( .A(n7122), .ZN(n7120) );
  NAND2_X1 U8054 ( .A1(n7122), .A2(n7127), .ZN(n7121) );
  OR2_X1 U8055 ( .A1(n9403), .A2(n10030), .ZN(n9161) );
  INV_X1 U8056 ( .A(n6682), .ZN(n6681) );
  OAI22_X1 U8057 ( .A1(n9177), .A2(n9800), .B1(n9841), .B2(n9860), .ZN(n6682)
         );
  NAND2_X1 U8058 ( .A1(n9472), .A2(n9471), .ZN(n13503) );
  NAND2_X1 U8059 ( .A1(n9464), .A2(n9463), .ZN(n13681) );
  NAND2_X1 U8060 ( .A1(n9445), .A2(n9444), .ZN(n13690) );
  OAI211_X1 U8061 ( .C1(n12613), .C2(n12288), .A(n12295), .B(n12287), .ZN(
        n12303) );
  OR2_X1 U8062 ( .A1(n9496), .A2(n9859), .ZN(n9154) );
  NAND2_X1 U8063 ( .A1(n10108), .A2(n10107), .ZN(n10261) );
  AND2_X1 U8064 ( .A1(n6910), .A2(n6909), .ZN(n10108) );
  NAND2_X1 U8065 ( .A1(n10106), .A2(n10922), .ZN(n6909) );
  NAND2_X1 U8066 ( .A1(n13410), .A2(n14929), .ZN(n6919) );
  INV_X1 U8067 ( .A(n6917), .ZN(n6916) );
  OAI21_X1 U8068 ( .B1(n13411), .B2(n14922), .A(n6918), .ZN(n6917) );
  NOR2_X1 U8069 ( .A1(n14914), .A2(n12613), .ZN(n6918) );
  XNOR2_X1 U8070 ( .A(n13432), .B(n13434), .ZN(n13653) );
  NAND2_X1 U8071 ( .A1(n7078), .A2(n7080), .ZN(n13561) );
  NAND2_X1 U8072 ( .A1(n7086), .A2(n7082), .ZN(n7078) );
  OR2_X1 U8073 ( .A1(n9799), .A2(n6790), .ZN(n9242) );
  NAND2_X1 U8074 ( .A1(n10021), .A2(n14953), .ZN(n13535) );
  NAND2_X1 U8075 ( .A1(n6791), .A2(n12168), .ZN(n9229) );
  INV_X1 U8076 ( .A(n9802), .ZN(n6791) );
  NAND2_X1 U8077 ( .A1(n13450), .A2(n9582), .ZN(n13655) );
  INV_X1 U8078 ( .A(n9581), .ZN(n9582) );
  NAND2_X1 U8079 ( .A1(n8054), .A2(n8053), .ZN(n14160) );
  AOI21_X1 U8080 ( .B1(n7345), .B2(n7347), .A(n7343), .ZN(n7342) );
  INV_X1 U8081 ( .A(n13798), .ZN(n7343) );
  NAND2_X1 U8082 ( .A1(n7660), .A2(n7659), .ZN(n14085) );
  XNOR2_X1 U8083 ( .A(n6932), .B(n8200), .ZN(n12605) );
  INV_X1 U8084 ( .A(n8451), .ZN(n8200) );
  NAND2_X1 U8085 ( .A1(n8497), .A2(n8199), .ZN(n6932) );
  NOR2_X1 U8086 ( .A1(n6598), .A2(n8477), .ZN(n8484) );
  NAND2_X1 U8087 ( .A1(n7515), .A2(n8021), .ZN(n14188) );
  NAND2_X1 U8088 ( .A1(n7943), .A2(n7942), .ZN(n11898) );
  OR2_X1 U8089 ( .A1(n7711), .A2(n9800), .ZN(n7231) );
  NAND2_X1 U8090 ( .A1(n11872), .A2(n8418), .ZN(n8113) );
  NAND2_X1 U8091 ( .A1(n14438), .A2(n7716), .ZN(n14410) );
  XNOR2_X1 U8092 ( .A(n14491), .B(n6696), .ZN(n15531) );
  INV_X1 U8093 ( .A(n14561), .ZN(n7288) );
  INV_X1 U8094 ( .A(n6697), .ZN(n14693) );
  AND2_X1 U8095 ( .A1(n14547), .A2(n14548), .ZN(n14573) );
  INV_X1 U8096 ( .A(n8267), .ZN(n7065) );
  INV_X1 U8097 ( .A(n12030), .ZN(n6774) );
  NOR2_X1 U8098 ( .A1(n12033), .A2(n12030), .ZN(n6773) );
  INV_X1 U8099 ( .A(n12049), .ZN(n7467) );
  NAND2_X1 U8100 ( .A1(n6803), .A2(n7047), .ZN(n6802) );
  NAND2_X1 U8101 ( .A1(n8283), .A2(n7048), .ZN(n7047) );
  AND2_X1 U8102 ( .A1(n7486), .A2(n7484), .ZN(n6759) );
  NAND2_X1 U8103 ( .A1(n6556), .A2(n7488), .ZN(n6760) );
  NAND2_X1 U8104 ( .A1(n7485), .A2(n7481), .ZN(n12072) );
  INV_X1 U8105 ( .A(n7482), .ZN(n7481) );
  OAI21_X1 U8106 ( .B1(n7486), .B2(n7484), .A(n7483), .ZN(n7482) );
  INV_X1 U8107 ( .A(n7480), .ZN(n7478) );
  NAND2_X1 U8108 ( .A1(n12078), .A2(n6594), .ZN(n7480) );
  INV_X1 U8109 ( .A(n12083), .ZN(n6776) );
  OR2_X1 U8110 ( .A1(n8294), .A2(n6826), .ZN(n6823) );
  AOI21_X1 U8111 ( .B1(n6821), .B2(n6826), .A(n6819), .ZN(n6818) );
  MUX2_X1 U8112 ( .A(n8320), .B(n8319), .S(n8376), .Z(n8328) );
  NAND2_X1 U8113 ( .A1(n7457), .A2(n7454), .ZN(n12097) );
  INV_X1 U8114 ( .A(n12102), .ZN(n6771) );
  INV_X1 U8115 ( .A(n12113), .ZN(n6769) );
  NOR2_X1 U8116 ( .A1(n12115), .A2(n6559), .ZN(n7469) );
  INV_X1 U8117 ( .A(n12135), .ZN(n6750) );
  INV_X1 U8118 ( .A(n6641), .ZN(n6751) );
  NOR2_X1 U8119 ( .A1(n8359), .A2(n8358), .ZN(n7062) );
  NAND2_X1 U8120 ( .A1(n8360), .A2(n7063), .ZN(n7061) );
  NAND2_X1 U8121 ( .A1(n8362), .A2(n7064), .ZN(n7063) );
  AOI21_X1 U8122 ( .B1(n6811), .B2(n6810), .A(n6809), .ZN(n6808) );
  AOI21_X1 U8123 ( .B1(n12141), .B2(n7492), .A(n6621), .ZN(n7491) );
  NOR2_X1 U8124 ( .A1(n7496), .A2(n12138), .ZN(n7492) );
  INV_X1 U8125 ( .A(n8704), .ZN(n7256) );
  NOR2_X1 U8126 ( .A1(n11310), .A2(n12087), .ZN(n11311) );
  NOR2_X1 U8127 ( .A1(n11753), .A2(n8336), .ZN(n7522) );
  NOR2_X1 U8128 ( .A1(n8353), .A2(n14199), .ZN(n7026) );
  INV_X1 U8129 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n7506) );
  NAND2_X1 U8130 ( .A1(n7405), .A2(SI_26_), .ZN(n7404) );
  INV_X1 U8131 ( .A(n8091), .ZN(n7405) );
  AOI21_X1 U8132 ( .B1(n7624), .B2(n7377), .A(n8062), .ZN(n7376) );
  AND2_X1 U8133 ( .A1(n7417), .A2(n7615), .ZN(n7416) );
  NAND2_X1 U8134 ( .A1(n7418), .A2(n7607), .ZN(n7417) );
  NAND2_X1 U8135 ( .A1(n7958), .A2(n7418), .ZN(n7415) );
  OAI21_X1 U8136 ( .B1(n7880), .B2(n7414), .A(n7546), .ZN(n7413) );
  INV_X1 U8137 ( .A(n7601), .ZN(n7410) );
  NAND2_X1 U8138 ( .A1(n7602), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n6710) );
  INV_X1 U8139 ( .A(n6691), .ZN(n14447) );
  OAI21_X1 U8140 ( .B1(n14495), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n6612), .ZN(
        n6691) );
  INV_X1 U8141 ( .A(n7319), .ZN(n7318) );
  AOI21_X1 U8142 ( .B1(n7319), .B2(n7317), .A(n7316), .ZN(n7315) );
  INV_X1 U8143 ( .A(n9699), .ZN(n7316) );
  NAND2_X1 U8144 ( .A1(n10880), .A2(n10900), .ZN(n6858) );
  AND2_X1 U8145 ( .A1(n6877), .A2(n12824), .ZN(n6874) );
  INV_X1 U8146 ( .A(n12863), .ZN(n6877) );
  INV_X1 U8147 ( .A(n7436), .ZN(n7435) );
  NAND2_X1 U8148 ( .A1(n8748), .A2(n11439), .ZN(n8767) );
  NOR2_X1 U8149 ( .A1(n8730), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n8748) );
  OR2_X1 U8150 ( .A1(n8688), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8714) );
  AND2_X1 U8151 ( .A1(n8658), .A2(n8657), .ZN(n8671) );
  AOI21_X1 U8152 ( .B1(n6993), .B2(n12384), .A(n6992), .ZN(n6991) );
  INV_X1 U8153 ( .A(n12447), .ZN(n6992) );
  INV_X1 U8154 ( .A(n12446), .ZN(n6993) );
  INV_X1 U8155 ( .A(n10397), .ZN(n9041) );
  NOR2_X1 U8156 ( .A1(n7245), .A2(n8982), .ZN(n7243) );
  OAI21_X1 U8157 ( .B1(n7247), .B2(n7246), .A(n6677), .ZN(n7245) );
  INV_X1 U8158 ( .A(n12359), .ZN(n7246) );
  NAND2_X1 U8159 ( .A1(n12607), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n7249) );
  NAND2_X1 U8160 ( .A1(n6839), .A2(n6838), .ZN(n8537) );
  NAND2_X1 U8161 ( .A1(n8522), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n6838) );
  NAND2_X1 U8162 ( .A1(n6840), .A2(P3_IR_REG_27__SCAN_IN), .ZN(n6839) );
  INV_X1 U8163 ( .A(n8697), .ZN(n6720) );
  INV_X1 U8164 ( .A(n8930), .ZN(n7270) );
  INV_X1 U8165 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n8856) );
  INV_X1 U8166 ( .A(n7257), .ZN(n7254) );
  NAND2_X1 U8167 ( .A1(n7259), .A2(n7256), .ZN(n7253) );
  NAND2_X1 U8168 ( .A1(n13277), .A2(n7129), .ZN(n7128) );
  INV_X1 U8169 ( .A(n13278), .ZN(n7129) );
  NOR2_X1 U8170 ( .A1(n13279), .A2(n13254), .ZN(n7130) );
  NAND2_X1 U8171 ( .A1(n7144), .A2(n12289), .ZN(n10428) );
  OR2_X1 U8172 ( .A1(n12219), .A2(n12182), .ZN(n12231) );
  INV_X1 U8173 ( .A(n6923), .ZN(n6921) );
  NAND2_X1 U8174 ( .A1(n6913), .A2(n6912), .ZN(n6911) );
  NAND2_X1 U8175 ( .A1(n14913), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n6912) );
  AND2_X1 U8176 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(n9495), .ZN(n9506) );
  NOR2_X1 U8177 ( .A1(n7184), .A2(n7187), .ZN(n7183) );
  INV_X1 U8178 ( .A(n7187), .ZN(n7182) );
  NAND2_X1 U8179 ( .A1(n7183), .A2(n7179), .ZN(n7178) );
  INV_X1 U8180 ( .A(n12244), .ZN(n7179) );
  OR2_X1 U8181 ( .A1(n13287), .A2(n13463), .ZN(n9514) );
  INV_X1 U8182 ( .A(n9572), .ZN(n7102) );
  NOR2_X1 U8183 ( .A1(n6590), .A2(n6786), .ZN(n6785) );
  AOI21_X1 U8184 ( .B1(n7170), .B2(n7173), .A(n6564), .ZN(n7167) );
  INV_X1 U8185 ( .A(n7170), .ZN(n7168) );
  OR2_X1 U8186 ( .A1(n13686), .A2(n13354), .ZN(n12274) );
  INV_X1 U8187 ( .A(n9447), .ZN(n9448) );
  NAND2_X1 U8188 ( .A1(n9448), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n9456) );
  INV_X1 U8189 ( .A(n7161), .ZN(n7160) );
  NOR2_X1 U8190 ( .A1(n13711), .A2(n12125), .ZN(n6972) );
  NOR2_X1 U8191 ( .A1(n12105), .A2(n11418), .ZN(n6969) );
  NAND2_X1 U8192 ( .A1(n11311), .A2(n9580), .ZN(n11418) );
  NOR2_X1 U8193 ( .A1(n12052), .A2(n10785), .ZN(n7193) );
  NAND2_X1 U8194 ( .A1(n10845), .A2(n6592), .ZN(n7192) );
  NAND2_X1 U8195 ( .A1(n12052), .A2(n10785), .ZN(n7194) );
  AND2_X1 U8196 ( .A1(n10530), .A2(n10529), .ZN(n11997) );
  NAND2_X1 U8197 ( .A1(n13479), .A2(n6976), .ZN(n13441) );
  NAND2_X1 U8198 ( .A1(n13460), .A2(n13471), .ZN(n6796) );
  NAND2_X1 U8199 ( .A1(n6794), .A2(n9576), .ZN(n6793) );
  NAND2_X1 U8200 ( .A1(n6796), .A2(n6578), .ZN(n6794) );
  AND3_X1 U8201 ( .A1(n10984), .A2(n6979), .A3(n6555), .ZN(n11011) );
  NAND2_X1 U8202 ( .A1(n10984), .A2(n6555), .ZN(n10923) );
  OAI21_X1 U8203 ( .B1(n7067), .B2(n7068), .A(n9542), .ZN(n10855) );
  OAI21_X1 U8204 ( .B1(n10240), .B2(n7069), .A(n9541), .ZN(n7068) );
  NOR2_X1 U8205 ( .A1(n10237), .A2(n7069), .ZN(n7067) );
  XNOR2_X1 U8206 ( .A(n10946), .B(n9196), .ZN(n10144) );
  INV_X1 U8207 ( .A(n7148), .ZN(n7146) );
  INV_X1 U8208 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n9295) );
  OR2_X1 U8209 ( .A1(n9239), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n9251) );
  AND2_X1 U8210 ( .A1(n9310), .A2(n9214), .ZN(n9226) );
  OR2_X1 U8211 ( .A1(n11971), .A2(n11970), .ZN(n7367) );
  INV_X1 U8212 ( .A(n11959), .ZN(n7359) );
  NOR2_X1 U8213 ( .A1(n13898), .A2(n7362), .ZN(n7361) );
  INV_X1 U8214 ( .A(n7363), .ZN(n7362) );
  AND2_X1 U8215 ( .A1(n7927), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n7944) );
  INV_X1 U8216 ( .A(n11159), .ZN(n6888) );
  OR2_X1 U8217 ( .A1(n7055), .A2(n8378), .ZN(n7054) );
  NOR2_X1 U8218 ( .A1(n8374), .A2(n8373), .ZN(n7053) );
  OR2_X1 U8219 ( .A1(n8468), .A2(n6695), .ZN(n8453) );
  NAND2_X1 U8220 ( .A1(n7046), .A2(n6627), .ZN(n7040) );
  NAND2_X1 U8221 ( .A1(n7041), .A2(n8410), .ZN(n7039) );
  NOR2_X1 U8222 ( .A1(n8494), .A2(n14085), .ZN(n7019) );
  NOR2_X1 U8223 ( .A1(n6958), .A2(n6957), .ZN(n6956) );
  INV_X1 U8224 ( .A(n8192), .ZN(n6957) );
  INV_X1 U8225 ( .A(n8194), .ZN(n6958) );
  NAND2_X1 U8226 ( .A1(n6955), .A2(n8194), .ZN(n6954) );
  INV_X1 U8227 ( .A(n6959), .ZN(n6955) );
  NOR2_X1 U8228 ( .A1(n7025), .A2(n14160), .ZN(n7024) );
  INV_X1 U8229 ( .A(n7026), .ZN(n7025) );
  AOI21_X1 U8230 ( .B1(n11279), .B2(n7511), .A(n7510), .ZN(n7509) );
  INV_X1 U8231 ( .A(n7845), .ZN(n7511) );
  NAND2_X1 U8232 ( .A1(n7509), .A2(n7512), .ZN(n7507) );
  AOI21_X1 U8233 ( .B1(n10496), .B2(n7221), .A(n7215), .ZN(n7214) );
  INV_X1 U8234 ( .A(n8174), .ZN(n7215) );
  NAND3_X1 U8235 ( .A1(n10307), .A2(n7016), .A3(n7014), .ZN(n7017) );
  AND2_X1 U8236 ( .A1(n7015), .A2(n10642), .ZN(n7014) );
  NOR2_X1 U8237 ( .A1(n8248), .A2(n8170), .ZN(n10182) );
  NAND2_X1 U8238 ( .A1(n14211), .A2(n7026), .ZN(n14176) );
  NAND2_X1 U8239 ( .A1(n8130), .A2(n8129), .ZN(n8391) );
  NOR2_X1 U8240 ( .A1(n7401), .A2(n7632), .ZN(n7400) );
  INV_X1 U8241 ( .A(n7403), .ZN(n7401) );
  INV_X1 U8242 ( .A(n7404), .ZN(n7398) );
  NAND2_X1 U8243 ( .A1(n8093), .A2(n7404), .ZN(n7402) );
  NAND2_X1 U8244 ( .A1(n8091), .A2(n13216), .ZN(n7403) );
  NAND2_X1 U8245 ( .A1(n7415), .A2(n7416), .ZN(n8024) );
  INV_X1 U8246 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n7647) );
  INV_X1 U8247 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n7646) );
  INV_X1 U8248 ( .A(n7899), .ZN(n7916) );
  NAND2_X1 U8249 ( .A1(n7411), .A2(n7596), .ZN(n7914) );
  OR2_X1 U8250 ( .A1(n7853), .A2(n7852), .ZN(n7866) );
  AOI21_X1 U8251 ( .B1(n7583), .B2(n7395), .A(n6617), .ZN(n7393) );
  INV_X1 U8252 ( .A(n7395), .ZN(n7394) );
  OR2_X1 U8253 ( .A1(n7819), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n7820) );
  NAND2_X1 U8254 ( .A1(n7579), .A2(SI_8_), .ZN(n7581) );
  NAND2_X1 U8255 ( .A1(n7576), .A2(SI_7_), .ZN(n7578) );
  NAND2_X2 U8256 ( .A1(n6684), .A2(n6683), .ZN(n7658) );
  INV_X1 U8257 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n14444) );
  XNOR2_X1 U8258 ( .A(n14445), .B(n14446), .ZN(n14495) );
  XNOR2_X1 U8259 ( .A(n14448), .B(n14447), .ZN(n14485) );
  NOR2_X1 U8260 ( .A1(n14458), .A2(n14457), .ZN(n14484) );
  NOR2_X1 U8261 ( .A1(n14510), .A2(n14456), .ZN(n14457) );
  AOI21_X1 U8262 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(n14460), .A(n14459), .ZN(
        n14517) );
  NOR2_X1 U8263 ( .A1(n14484), .A2(n14483), .ZN(n14459) );
  NOR2_X1 U8264 ( .A1(n6560), .A2(n7287), .ZN(n7286) );
  AOI21_X1 U8265 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(n14464), .A(n14463), .ZN(
        n14523) );
  OR2_X1 U8266 ( .A1(n11437), .A2(n9674), .ZN(n7339) );
  NOR2_X1 U8267 ( .A1(n12640), .A2(n7320), .ZN(n7319) );
  INV_X1 U8268 ( .A(n9695), .ZN(n7320) );
  NAND2_X1 U8269 ( .A1(n12680), .A2(n12679), .ZN(n7321) );
  AOI21_X1 U8270 ( .B1(n7309), .B2(n7311), .A(n6579), .ZN(n7307) );
  INV_X1 U8271 ( .A(n9651), .ZN(n7309) );
  INV_X1 U8272 ( .A(n7311), .ZN(n7310) );
  AND2_X1 U8273 ( .A1(n9666), .A2(n7323), .ZN(n7322) );
  INV_X1 U8274 ( .A(n7327), .ZN(n7323) );
  INV_X1 U8275 ( .A(n7325), .ZN(n7324) );
  OAI21_X1 U8276 ( .B1(n7327), .B2(n9669), .A(n9670), .ZN(n7325) );
  NAND2_X1 U8277 ( .A1(n11119), .A2(n9669), .ZN(n11514) );
  OR2_X1 U8278 ( .A1(n8767), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8785) );
  NOR2_X1 U8279 ( .A1(n8785), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n8805) );
  AND2_X1 U8280 ( .A1(n14620), .A2(n14610), .ZN(n12574) );
  NAND2_X1 U8281 ( .A1(n7200), .A2(n10205), .ZN(n10327) );
  NAND2_X1 U8282 ( .A1(n10345), .A2(n10203), .ZN(n7200) );
  AND2_X1 U8283 ( .A1(n10223), .A2(n6862), .ZN(n10337) );
  NAND2_X1 U8284 ( .A1(n10220), .A2(n10345), .ZN(n6862) );
  AOI21_X1 U8285 ( .B1(n10336), .B2(n6862), .A(n10229), .ZN(n15042) );
  OR2_X1 U8286 ( .A1(n15067), .A2(n15066), .ZN(n15064) );
  NOR2_X1 U8287 ( .A1(n10895), .A2(n10860), .ZN(n7205) );
  OR2_X1 U8288 ( .A1(n15075), .A2(n8603), .ZN(n15073) );
  AND2_X1 U8289 ( .A1(n12345), .A2(n7212), .ZN(n10862) );
  NAND2_X1 U8290 ( .A1(n12351), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n7212) );
  NOR2_X1 U8291 ( .A1(n6860), .A2(n6852), .ZN(n6851) );
  INV_X1 U8292 ( .A(n6858), .ZN(n6852) );
  NAND2_X1 U8293 ( .A1(n12332), .A2(n10902), .ZN(n12318) );
  INV_X1 U8294 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n15461) );
  OR2_X1 U8295 ( .A1(n10867), .A2(n15444), .ZN(n7208) );
  OR2_X1 U8296 ( .A1(n15093), .A2(n15444), .ZN(n7209) );
  AOI21_X1 U8297 ( .B1(n6845), .B2(n6848), .A(n6843), .ZN(n6842) );
  INV_X1 U8298 ( .A(n15096), .ZN(n6843) );
  NAND2_X1 U8299 ( .A1(n15107), .A2(n10905), .ZN(n10906) );
  AND2_X1 U8300 ( .A1(n6866), .A2(n6865), .ZN(n12753) );
  NOR2_X1 U8301 ( .A1(n11502), .A2(n11499), .ZN(n6865) );
  NAND2_X1 U8302 ( .A1(n11491), .A2(n11492), .ZN(n11495) );
  NAND2_X1 U8303 ( .A1(n11495), .A2(n11494), .ZN(n12750) );
  NAND2_X1 U8304 ( .A1(n12750), .A2(n6743), .ZN(n12771) );
  OR2_X1 U8305 ( .A1(n12751), .A2(n11493), .ZN(n6743) );
  NOR2_X1 U8306 ( .A1(n12753), .A2(n6863), .ZN(n12757) );
  NOR2_X1 U8307 ( .A1(n6864), .A2(n12751), .ZN(n6863) );
  INV_X1 U8308 ( .A(n12755), .ZN(n6864) );
  INV_X1 U8309 ( .A(n12835), .ZN(n7203) );
  OR2_X1 U8310 ( .A1(n12800), .A2(n12801), .ZN(n7204) );
  OAI211_X1 U8311 ( .C1(n12808), .C2(n6876), .A(n6875), .B(n12862), .ZN(n14585) );
  NAND2_X1 U8312 ( .A1(n6878), .A2(n6877), .ZN(n6876) );
  NAND2_X1 U8313 ( .A1(n12825), .A2(n6874), .ZN(n6875) );
  INV_X1 U8314 ( .A(n12809), .ZN(n6878) );
  AND2_X1 U8315 ( .A1(n12845), .A2(n12844), .ZN(n12846) );
  INV_X1 U8316 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n6734) );
  NOR2_X1 U8317 ( .A1(n6732), .A2(n6725), .ZN(n6724) );
  NOR2_X1 U8318 ( .A1(n6733), .A2(n6734), .ZN(n6725) );
  NAND2_X1 U8319 ( .A1(n12856), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n6738) );
  XNOR2_X1 U8320 ( .A(n6873), .B(n12868), .ZN(n6872) );
  NOR2_X1 U8321 ( .A1(n14595), .A2(n6588), .ZN(n6873) );
  AND2_X1 U8322 ( .A1(n12365), .A2(n12364), .ZN(n12377) );
  OR2_X1 U8323 ( .A1(n9062), .A2(n12561), .ZN(n9063) );
  OR2_X1 U8324 ( .A1(n8970), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8985) );
  AND2_X1 U8325 ( .A1(n8875), .A2(n8874), .ZN(n8887) );
  OR2_X1 U8326 ( .A1(n8843), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8862) );
  NOR2_X1 U8327 ( .A1(n8862), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8875) );
  NAND2_X1 U8328 ( .A1(n8822), .A2(n8821), .ZN(n8843) );
  AND2_X1 U8329 ( .A1(n8805), .A2(n8804), .ZN(n8822) );
  NAND2_X1 U8330 ( .A1(n8793), .A2(n8792), .ZN(n13051) );
  OAI21_X1 U8331 ( .B1(n8756), .B2(n7431), .A(n7429), .ZN(n8793) );
  INV_X1 U8332 ( .A(n7430), .ZN(n7429) );
  NAND2_X1 U8333 ( .A1(n13057), .A2(n13056), .ZN(n13055) );
  AND2_X1 U8334 ( .A1(n12509), .A2(n13042), .ZN(n13056) );
  NAND2_X1 U8335 ( .A1(n13072), .A2(n13071), .ZN(n13070) );
  NAND2_X1 U8336 ( .A1(n12413), .A2(n12477), .ZN(n7003) );
  INV_X1 U8337 ( .A(n7424), .ZN(n7423) );
  OAI21_X1 U8338 ( .B1(n12469), .B2(n6576), .A(n8720), .ZN(n7424) );
  INV_X1 U8339 ( .A(n11518), .ZN(n11624) );
  NAND2_X1 U8340 ( .A1(n11208), .A2(n12457), .ZN(n11341) );
  INV_X1 U8341 ( .A(n12389), .ZN(n12457) );
  NAND2_X1 U8342 ( .A1(n7442), .A2(n7441), .ZN(n11174) );
  AOI21_X1 U8343 ( .B1(n7443), .B2(n12437), .A(n6589), .ZN(n7441) );
  OR2_X1 U8344 ( .A1(n8620), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8638) );
  INV_X1 U8345 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n10836) );
  NAND2_X1 U8346 ( .A1(n8599), .A2(n10836), .ZN(n8620) );
  NAND2_X1 U8347 ( .A1(n11200), .A2(n8580), .ZN(n10728) );
  INV_X1 U8348 ( .A(n12433), .ZN(n10727) );
  NAND2_X1 U8349 ( .A1(n15122), .A2(n8569), .ZN(n11198) );
  NAND2_X1 U8350 ( .A1(n15122), .A2(n7427), .ZN(n11200) );
  NOR2_X1 U8351 ( .A1(n12385), .A2(n7428), .ZN(n7427) );
  INV_X1 U8352 ( .A(n8569), .ZN(n7428) );
  NAND2_X1 U8353 ( .A1(n12422), .A2(n12418), .ZN(n15142) );
  NAND2_X1 U8354 ( .A1(n15142), .A2(n15141), .ZN(n15140) );
  NAND2_X1 U8355 ( .A1(n8594), .A2(SI_1_), .ZN(n8542) );
  NAND2_X1 U8356 ( .A1(n8905), .A2(n8904), .ZN(n12686) );
  NAND2_X1 U8357 ( .A1(n8594), .A2(SI_22_), .ZN(n8904) );
  NAND2_X1 U8358 ( .A1(n8594), .A2(n9764), .ZN(n8654) );
  AND3_X1 U8359 ( .A1(n8636), .A2(n8635), .A3(n8634), .ZN(n15178) );
  NAND2_X1 U8360 ( .A1(n8594), .A2(SI_6_), .ZN(n8636) );
  NAND2_X1 U8361 ( .A1(n7242), .A2(n6570), .ZN(n12367) );
  NAND2_X1 U8362 ( .A1(n7447), .A2(n8536), .ZN(n7446) );
  INV_X1 U8363 ( .A(n7448), .ZN(n7447) );
  INV_X1 U8364 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n8523) );
  NAND2_X1 U8365 ( .A1(n7248), .A2(n7249), .ZN(n7247) );
  AND2_X1 U8366 ( .A1(n9077), .A2(n9076), .ZN(n9089) );
  OAI21_X1 U8367 ( .B1(n9078), .B2(P3_IR_REG_25__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9075) );
  NAND2_X1 U8368 ( .A1(n9022), .A2(n9021), .ZN(n9025) );
  NAND2_X1 U8369 ( .A1(n15400), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n7266) );
  INV_X1 U8370 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n8835) );
  OR2_X1 U8371 ( .A1(n8838), .A2(P3_IR_REG_18__SCAN_IN), .ZN(n8855) );
  AND3_X1 U8372 ( .A1(n8511), .A2(n8512), .A3(n7330), .ZN(n8817) );
  NOR2_X1 U8373 ( .A1(n8514), .A2(P3_IR_REG_15__SCAN_IN), .ZN(n7330) );
  NAND2_X1 U8374 ( .A1(n6705), .A2(n6704), .ZN(n8667) );
  INV_X1 U8375 ( .A(n8651), .ZN(n6704) );
  OR2_X1 U8376 ( .A1(n8632), .A2(P3_IR_REG_6__SCAN_IN), .ZN(n8646) );
  OR2_X1 U8377 ( .A1(n8646), .A2(P3_IR_REG_7__SCAN_IN), .ZN(n8677) );
  XNOR2_X1 U8378 ( .A(n9801), .B(P2_DATAO_REG_6__SCAN_IN), .ZN(n8648) );
  AND2_X1 U8379 ( .A1(n8627), .A2(n8614), .ZN(n8615) );
  NAND2_X1 U8380 ( .A1(n10030), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n8561) );
  OAI22_X1 U8381 ( .A1(n10204), .A2(n6722), .B1(P3_IR_REG_31__SCAN_IN), .B2(
        P3_IR_REG_2__SCAN_IN), .ZN(n8558) );
  NAND2_X1 U8382 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_2__SCAN_IN), .ZN(
        n6722) );
  XNOR2_X1 U8383 ( .A(n12021), .B(n13236), .ZN(n10312) );
  AOI21_X1 U8384 ( .B1(n7135), .B2(n7134), .A(n6618), .ZN(n7133) );
  INV_X1 U8385 ( .A(n11864), .ZN(n7134) );
  INV_X1 U8386 ( .A(n7130), .ZN(n7126) );
  NAND2_X1 U8387 ( .A1(n9380), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n9415) );
  NAND2_X1 U8388 ( .A1(n13324), .A2(n13243), .ZN(n13244) );
  NOR2_X1 U8389 ( .A1(n11407), .A2(n7142), .ZN(n7141) );
  INV_X1 U8390 ( .A(n11404), .ZN(n7142) );
  NAND2_X1 U8391 ( .A1(n11863), .A2(n11864), .ZN(n11875) );
  NOR2_X1 U8392 ( .A1(n9473), .A2(n13298), .ZN(n9486) );
  AND2_X1 U8393 ( .A1(n9578), .A2(n10529), .ZN(n10015) );
  CLKBUF_X1 U8394 ( .A(n11830), .Z(n11698) );
  OR2_X1 U8395 ( .A1(n9345), .A2(n9344), .ZN(n9355) );
  AND2_X1 U8396 ( .A1(n12192), .A2(n6763), .ZN(n6762) );
  NAND2_X1 U8397 ( .A1(n6766), .A2(n6765), .ZN(n6763) );
  NOR2_X1 U8398 ( .A1(n7148), .A2(n7151), .ZN(n7147) );
  NAND2_X1 U8399 ( .A1(n9896), .A2(n6908), .ZN(n14818) );
  OR2_X1 U8400 ( .A1(n9861), .A2(n9862), .ZN(n6908) );
  NAND2_X1 U8401 ( .A1(n14818), .A2(n14819), .ZN(n14817) );
  NAND2_X1 U8402 ( .A1(n14817), .A2(n6907), .ZN(n14830) );
  OR2_X1 U8403 ( .A1(n14825), .A2(n9864), .ZN(n6907) );
  NAND2_X1 U8404 ( .A1(n14830), .A2(n14831), .ZN(n14829) );
  OR2_X1 U8405 ( .A1(n9984), .A2(n9985), .ZN(n6910) );
  OR2_X1 U8406 ( .A1(n14871), .A2(n14872), .ZN(n14869) );
  NAND2_X1 U8407 ( .A1(n6924), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n6923) );
  AND2_X1 U8408 ( .A1(n11099), .A2(n11100), .ZN(n13401) );
  AND2_X1 U8409 ( .A1(n6976), .A2(n6975), .ZN(n6974) );
  OAI21_X1 U8410 ( .B1(n9491), .B2(n7180), .A(n7177), .ZN(n13435) );
  INV_X1 U8411 ( .A(n7183), .ZN(n7180) );
  AND2_X1 U8412 ( .A1(n7178), .A2(n7181), .ZN(n7177) );
  NAND2_X1 U8413 ( .A1(n7186), .A2(n7182), .ZN(n7181) );
  NOR2_X1 U8414 ( .A1(n13471), .A2(n7098), .ZN(n7097) );
  INV_X1 U8415 ( .A(n9574), .ZN(n7098) );
  NAND2_X1 U8416 ( .A1(n13479), .A2(n13485), .ZN(n13480) );
  NAND2_X1 U8417 ( .A1(n7164), .A2(n7167), .ZN(n13492) );
  OR2_X1 U8418 ( .A1(n13531), .A2(n7168), .ZN(n7164) );
  NOR2_X1 U8419 ( .A1(n9456), .A2(n13263), .ZN(n9466) );
  OR2_X1 U8420 ( .A1(n13538), .A2(n13681), .ZN(n13518) );
  INV_X1 U8421 ( .A(n9567), .ZN(n7081) );
  NOR2_X1 U8422 ( .A1(n13569), .A2(n7088), .ZN(n7084) );
  AND2_X1 U8423 ( .A1(n11848), .A2(n6634), .ZN(n13588) );
  AND2_X1 U8424 ( .A1(n7533), .A2(n9387), .ZN(n7175) );
  NAND2_X1 U8425 ( .A1(n11848), .A2(n6972), .ZN(n7532) );
  NAND2_X1 U8426 ( .A1(n7176), .A2(n9387), .ZN(n13617) );
  NAND2_X1 U8427 ( .A1(n11848), .A2(n13765), .ZN(n13632) );
  NAND2_X1 U8428 ( .A1(n6969), .A2(n6968), .ZN(n11810) );
  INV_X1 U8429 ( .A(n7107), .ZN(n7106) );
  OAI21_X1 U8430 ( .B1(n12270), .B2(n7108), .A(n9558), .ZN(n7107) );
  NAND2_X1 U8431 ( .A1(n9556), .A2(n9557), .ZN(n7108) );
  NOR2_X1 U8432 ( .A1(n12270), .A2(n7110), .ZN(n7109) );
  INV_X1 U8433 ( .A(n9557), .ZN(n7110) );
  NAND2_X1 U8434 ( .A1(n7104), .A2(n7103), .ZN(n11803) );
  AND2_X1 U8435 ( .A1(n7106), .A2(n12266), .ZN(n7103) );
  NAND2_X1 U8436 ( .A1(n6782), .A2(n12105), .ZN(n6779) );
  NAND2_X1 U8437 ( .A1(n6781), .A2(n6605), .ZN(n6780) );
  INV_X1 U8438 ( .A(n6969), .ZN(n11692) );
  NOR2_X1 U8439 ( .A1(n9303), .A2(n9302), .ZN(n9317) );
  OR2_X1 U8440 ( .A1(n9287), .A2(n10115), .ZN(n9303) );
  NAND2_X1 U8441 ( .A1(n9272), .A2(n9271), .ZN(n12068) );
  OR2_X1 U8442 ( .A1(n9839), .A2(n6790), .ZN(n9272) );
  NOR2_X1 U8443 ( .A1(n9244), .A2(n9243), .ZN(n9262) );
  AND2_X1 U8444 ( .A1(n7192), .A2(n7189), .ZN(n10716) );
  INV_X1 U8445 ( .A(n7193), .ZN(n7189) );
  AND2_X1 U8446 ( .A1(n14974), .A2(n10851), .ZN(n10984) );
  NAND2_X1 U8447 ( .A1(n10984), .A2(n14981), .ZN(n10983) );
  AND2_X1 U8448 ( .A1(n9237), .A2(n9238), .ZN(n12254) );
  NAND2_X1 U8449 ( .A1(n7153), .A2(n9212), .ZN(n10659) );
  NOR2_X1 U8450 ( .A1(n10664), .A2(n6721), .ZN(n10851) );
  OR2_X1 U8451 ( .A1(n10239), .A2(n12025), .ZN(n10664) );
  NOR2_X1 U8452 ( .A1(n10074), .A2(n12016), .ZN(n10146) );
  NAND2_X1 U8453 ( .A1(n10146), .A2(n10946), .ZN(n10239) );
  NAND2_X1 U8454 ( .A1(n7406), .A2(n6663), .ZN(n12166) );
  NAND2_X1 U8455 ( .A1(n12195), .A2(n12194), .ZN(n13426) );
  NAND2_X1 U8456 ( .A1(n6792), .A2(n12168), .ZN(n12195) );
  INV_X1 U8457 ( .A(n14432), .ZN(n6792) );
  NAND2_X1 U8458 ( .A1(n6680), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9156) );
  OR2_X1 U8459 ( .A1(n9591), .A2(P2_IR_REG_25__SCAN_IN), .ZN(n9594) );
  AND2_X1 U8461 ( .A1(n9188), .A2(n9199), .ZN(n9863) );
  OR2_X1 U8462 ( .A1(n7348), .A2(n7346), .ZN(n7345) );
  AND2_X1 U8463 ( .A1(n13890), .A2(n7349), .ZN(n7348) );
  INV_X1 U8464 ( .A(n7351), .ZN(n7346) );
  OR2_X1 U8465 ( .A1(n13841), .A2(n7350), .ZN(n7349) );
  NAND2_X1 U8466 ( .A1(n7351), .A2(n11909), .ZN(n7347) );
  OAI21_X1 U8467 ( .B1(n7357), .B2(n7356), .A(n6620), .ZN(n7354) );
  INV_X1 U8468 ( .A(n7361), .ZN(n7360) );
  INV_X1 U8469 ( .A(n13783), .ZN(n7356) );
  INV_X1 U8470 ( .A(n10356), .ZN(n10357) );
  NAND2_X1 U8471 ( .A1(n6708), .A2(n6884), .ZN(n13830) );
  AND2_X1 U8472 ( .A1(n6584), .A2(n13831), .ZN(n6708) );
  NAND2_X1 U8473 ( .A1(n7944), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n8004) );
  NOR2_X1 U8474 ( .A1(n8055), .A2(n13792), .ZN(n8066) );
  NAND2_X1 U8475 ( .A1(n11156), .A2(n6575), .ZN(n11368) );
  NAND2_X1 U8476 ( .A1(n10038), .A2(n10037), .ZN(n10360) );
  OR2_X1 U8477 ( .A1(n8044), .A2(n13869), .ZN(n8055) );
  OR2_X1 U8478 ( .A1(n11936), .A2(n11935), .ZN(n11937) );
  OR2_X1 U8479 ( .A1(n7839), .A2(n7838), .ZN(n7857) );
  CLKBUF_X1 U8480 ( .A(n13876), .Z(n13877) );
  NAND2_X1 U8481 ( .A1(n6902), .A2(n6901), .ZN(n6900) );
  INV_X1 U8482 ( .A(n13790), .ZN(n6901) );
  INV_X1 U8483 ( .A(n6903), .ZN(n6902) );
  NOR2_X1 U8484 ( .A1(n7664), .A2(n7503), .ZN(n7505) );
  NAND2_X1 U8485 ( .A1(n6828), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n7503) );
  NAND2_X1 U8486 ( .A1(n7019), .A2(n7018), .ZN(n14073) );
  INV_X1 U8487 ( .A(n7019), .ZN(n8495) );
  AND2_X1 U8488 ( .A1(n6964), .A2(n8474), .ZN(n6963) );
  NOR2_X1 U8489 ( .A1(n8448), .A2(n14755), .ZN(n6716) );
  INV_X1 U8490 ( .A(n7021), .ZN(n14110) );
  INV_X1 U8491 ( .A(n8446), .ZN(n14123) );
  AOI21_X1 U8492 ( .B1(n7528), .B2(n6961), .A(n6583), .ZN(n7527) );
  OAI21_X1 U8493 ( .B1(n14172), .B2(n6952), .A(n6950), .ZN(n14141) );
  AOI21_X1 U8494 ( .B1(n6954), .B2(n6951), .A(n8075), .ZN(n6950) );
  INV_X1 U8495 ( .A(n6954), .ZN(n6952) );
  INV_X1 U8496 ( .A(n6956), .ZN(n6951) );
  NAND2_X1 U8497 ( .A1(n6949), .A2(n6954), .ZN(n7547) );
  NAND2_X1 U8498 ( .A1(n14172), .A2(n6956), .ZN(n6949) );
  INV_X1 U8499 ( .A(n7222), .ZN(n6931) );
  OR2_X1 U8500 ( .A1(n7857), .A2(n11549), .ZN(n7871) );
  NOR2_X1 U8501 ( .A1(n7871), .A2(n7870), .ZN(n7890) );
  NAND2_X1 U8502 ( .A1(n7013), .A2(n7012), .ZN(n11281) );
  NAND2_X1 U8503 ( .A1(n11183), .A2(n7845), .ZN(n11280) );
  NAND2_X1 U8504 ( .A1(n11280), .A2(n11279), .ZN(n11461) );
  NAND2_X1 U8505 ( .A1(n6554), .A2(n11018), .ZN(n6940) );
  AOI21_X1 U8506 ( .B1(n11021), .B2(n6554), .A(n6610), .ZN(n6939) );
  NOR2_X2 U8507 ( .A1(n10969), .A2(n7017), .ZN(n10815) );
  AND3_X1 U8508 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n7776) );
  NAND2_X1 U8509 ( .A1(n7214), .A2(n7216), .ZN(n10539) );
  NAND2_X1 U8510 ( .A1(n7218), .A2(n7217), .ZN(n10491) );
  NAND2_X1 U8511 ( .A1(n10285), .A2(n8173), .ZN(n10492) );
  NAND2_X1 U8512 ( .A1(n10286), .A2(n10287), .ZN(n10285) );
  NOR2_X1 U8513 ( .A1(n6832), .A2(n6831), .ZN(n6830) );
  NAND2_X1 U8514 ( .A1(n8421), .A2(n8420), .ZN(n8454) );
  NAND2_X1 U8515 ( .A1(n8417), .A2(n8418), .ZN(n8421) );
  NAND2_X1 U8516 ( .A1(n7518), .A2(n6585), .ZN(n8491) );
  NAND2_X1 U8517 ( .A1(n7963), .A2(n7962), .ZN(n14358) );
  NAND2_X1 U8518 ( .A1(n7731), .A2(n7732), .ZN(n10379) );
  NAND2_X1 U8519 ( .A1(n8413), .A2(n8412), .ZN(n8416) );
  XNOR2_X1 U8520 ( .A(n8391), .B(n8390), .ZN(n13774) );
  OAI21_X1 U8521 ( .B1(n8052), .B2(n7377), .A(n7624), .ZN(n8063) );
  XNOR2_X1 U8522 ( .A(n7992), .B(n7991), .ZN(n10991) );
  NAND2_X1 U8523 ( .A1(n7818), .A2(n7584), .ZN(n7830) );
  NAND2_X1 U8524 ( .A1(n7816), .A2(n7815), .ZN(n7818) );
  OR2_X1 U8525 ( .A1(n7751), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n7753) );
  INV_X1 U8526 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n7645) );
  CLKBUF_X1 U8527 ( .A(n7684), .Z(n7685) );
  INV_X1 U8528 ( .A(n7280), .ZN(n14487) );
  OAI21_X1 U8529 ( .B1(n14441), .B2(n14489), .A(n7281), .ZN(n7280) );
  NAND2_X1 U8530 ( .A1(n14442), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n7281) );
  NOR2_X1 U8531 ( .A1(n14504), .A2(n14505), .ZN(n14506) );
  NOR2_X1 U8532 ( .A1(n14452), .A2(n14451), .ZN(n14507) );
  NAND2_X1 U8533 ( .A1(n14512), .A2(n14513), .ZN(n14514) );
  OAI21_X1 U8534 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(n14468), .A(n14467), .ZN(
        n14529) );
  OAI21_X1 U8535 ( .B1(n7292), .B2(n7297), .A(n14891), .ZN(n7291) );
  NAND2_X1 U8536 ( .A1(n7339), .A2(n9676), .ZN(n11641) );
  INV_X1 U8537 ( .A(n12969), .ZN(n13101) );
  NAND2_X1 U8538 ( .A1(n11122), .A2(n9666), .ZN(n11119) );
  CLKBUF_X1 U8539 ( .A(n11044), .Z(n11122) );
  OR2_X1 U8540 ( .A1(n9643), .A2(n15137), .ZN(n10480) );
  AOI21_X1 U8541 ( .B1(n7304), .B2(n7306), .A(n6593), .ZN(n7302) );
  NAND2_X1 U8542 ( .A1(n7321), .A2(n9695), .ZN(n12639) );
  NAND2_X1 U8543 ( .A1(n7308), .A2(n7311), .ZN(n11107) );
  NAND2_X1 U8544 ( .A1(n10651), .A2(n9651), .ZN(n7308) );
  NAND2_X1 U8545 ( .A1(n10648), .A2(n9651), .ZN(n10834) );
  NAND2_X1 U8546 ( .A1(n7314), .A2(n7313), .ZN(n10648) );
  INV_X1 U8547 ( .A(n10650), .ZN(n7313) );
  INV_X1 U8548 ( .A(n10651), .ZN(n7314) );
  NAND2_X1 U8549 ( .A1(n7303), .A2(n9688), .ZN(n12696) );
  NAND2_X1 U8550 ( .A1(n12661), .A2(n12660), .ZN(n7303) );
  NAND2_X1 U8551 ( .A1(n7336), .A2(n7334), .ZN(n11710) );
  AOI21_X1 U8552 ( .B1(n7337), .B2(n9674), .A(n7335), .ZN(n7334) );
  INV_X1 U8553 ( .A(n9680), .ZN(n7335) );
  INV_X1 U8554 ( .A(n12926), .ZN(n12657) );
  NAND4_X1 U8555 ( .A1(n8676), .A2(n8675), .A3(n8674), .A4(n8673), .ZN(n12739)
         );
  AND2_X1 U8556 ( .A1(n7196), .A2(n7195), .ZN(n15055) );
  XNOR2_X1 U8557 ( .A(n10861), .B(n10896), .ZN(n15075) );
  AOI21_X1 U8558 ( .B1(n15087), .B2(P3_REG1_REG_5__SCAN_IN), .A(n6741), .ZN(
        n12349) );
  OAI21_X1 U8559 ( .B1(n12343), .B2(n12344), .A(n6859), .ZN(n12329) );
  NAND2_X1 U8560 ( .A1(n6850), .A2(n6853), .ZN(n12313) );
  NAND2_X1 U8561 ( .A1(n12343), .A2(n6851), .ZN(n6850) );
  NAND2_X1 U8562 ( .A1(n7207), .A2(n7206), .ZN(n11245) );
  INV_X1 U8563 ( .A(n6868), .ZN(n11256) );
  XNOR2_X1 U8564 ( .A(n12771), .B(n12783), .ZN(n12752) );
  NOR2_X1 U8565 ( .A1(n12749), .A2(n11722), .ZN(n12767) );
  OAI21_X1 U8566 ( .B1(n12749), .B2(n7211), .A(n7210), .ZN(n12798) );
  NAND2_X1 U8567 ( .A1(n12787), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n7211) );
  INV_X1 U8568 ( .A(n7204), .ZN(n12834) );
  NOR2_X1 U8569 ( .A1(n12823), .A2(n6879), .ZN(n12864) );
  NAND2_X1 U8570 ( .A1(n12819), .A2(n12820), .ZN(n12849) );
  XNOR2_X1 U8571 ( .A(n12846), .B(n14580), .ZN(n14577) );
  NAND2_X1 U8572 ( .A1(n12860), .A2(n6738), .ZN(n6732) );
  AND2_X1 U8573 ( .A1(n12372), .A2(n12371), .ZN(n14614) );
  INV_X1 U8574 ( .A(n12377), .ZN(n14623) );
  XNOR2_X1 U8575 ( .A(n12379), .B(n9065), .ZN(n11993) );
  AND2_X1 U8576 ( .A1(n9003), .A2(n9002), .ZN(n14611) );
  AND2_X1 U8577 ( .A1(n12878), .A2(n12877), .ZN(n13081) );
  AOI211_X1 U8578 ( .C1(n12945), .C2(n13085), .A(n12893), .B(n12892), .ZN(
        n13087) );
  OR2_X1 U8579 ( .A1(n12937), .A2(n6986), .ZN(n6982) );
  NAND2_X1 U8580 ( .A1(n8969), .A2(n8968), .ZN(n12913) );
  NAND2_X1 U8581 ( .A1(n12542), .A2(n12941), .ZN(n12924) );
  AND3_X1 U8582 ( .A1(n12965), .A2(n12964), .A3(n12963), .ZN(n13104) );
  NAND2_X1 U8583 ( .A1(n8897), .A2(n8896), .ZN(n12972) );
  NAND2_X1 U8584 ( .A1(n8873), .A2(n8872), .ZN(n13000) );
  NAND2_X1 U8585 ( .A1(n8594), .A2(SI_20_), .ZN(n8872) );
  NAND2_X1 U8586 ( .A1(n13020), .A2(n8849), .ZN(n13008) );
  NAND2_X1 U8587 ( .A1(n13039), .A2(n8829), .ZN(n13022) );
  NAND2_X1 U8588 ( .A1(n13045), .A2(n12516), .ZN(n13030) );
  NAND2_X1 U8589 ( .A1(n8842), .A2(n8841), .ZN(n13122) );
  NAND2_X1 U8590 ( .A1(n11791), .A2(n8773), .ZN(n13063) );
  AND2_X1 U8591 ( .A1(n15132), .A2(n11448), .ZN(n13077) );
  NAND2_X1 U8592 ( .A1(n8766), .A2(n8765), .ZN(n13140) );
  NAND2_X1 U8593 ( .A1(n8756), .A2(n8755), .ZN(n11788) );
  NAND2_X1 U8594 ( .A1(n7426), .A2(n8702), .ZN(n11526) );
  NAND2_X1 U8595 ( .A1(n7005), .A2(n12459), .ZN(n11339) );
  NAND2_X1 U8596 ( .A1(n11072), .A2(n7443), .ZN(n11061) );
  NAND2_X1 U8597 ( .A1(n8594), .A2(n9787), .ZN(n8578) );
  AND2_X1 U8598 ( .A1(n10804), .A2(n9071), .ZN(n15134) );
  INV_X1 U8599 ( .A(n15118), .ZN(n15150) );
  NAND2_X1 U8600 ( .A1(n8860), .A2(n8859), .ZN(n13175) );
  AND2_X1 U8601 ( .A1(n8803), .A2(n8802), .ZN(n13184) );
  XNOR2_X1 U8602 ( .A(n12360), .B(n9016), .ZN(n13201) );
  NAND2_X1 U8603 ( .A1(n7244), .A2(n7247), .ZN(n12360) );
  NAND2_X1 U8604 ( .A1(n7250), .A2(n6674), .ZN(n7244) );
  INV_X1 U8605 ( .A(n7271), .ZN(n8931) );
  OAI21_X1 U8606 ( .B1(n6693), .B2(n7259), .A(n7257), .ZN(n8705) );
  NAND2_X1 U8607 ( .A1(n7262), .A2(n8682), .ZN(n8695) );
  NAND2_X1 U8608 ( .A1(n6693), .A2(n8680), .ZN(n7262) );
  NAND2_X1 U8609 ( .A1(n7239), .A2(n7237), .ZN(n8613) );
  NAND2_X1 U8610 ( .A1(n7239), .A2(n8588), .ZN(n8592) );
  INV_X1 U8611 ( .A(n10893), .ZN(n15045) );
  XOR2_X1 U8612 ( .A(n13278), .B(n13277), .Z(n13279) );
  NAND2_X1 U8613 ( .A1(n7131), .A2(n7133), .ZN(n13272) );
  NAND2_X1 U8614 ( .A1(n7143), .A2(n11404), .ZN(n11406) );
  NAND2_X1 U8615 ( .A1(n9365), .A2(n9364), .ZN(n13726) );
  AOI21_X1 U8616 ( .B1(n10440), .B2(n10439), .A(n10438), .ZN(n10471) );
  NAND2_X1 U8617 ( .A1(n10936), .A2(n10935), .ZN(n10937) );
  NAND2_X1 U8618 ( .A1(n9327), .A2(n9326), .ZN(n12092) );
  AND2_X1 U8619 ( .A1(n10023), .A2(n12305), .ZN(n13342) );
  NAND2_X1 U8620 ( .A1(n11875), .A2(n11874), .ZN(n13223) );
  INV_X1 U8621 ( .A(n12300), .ZN(n12301) );
  NAND4_X1 U8622 ( .A1(n9195), .A2(n9194), .A3(n9193), .A4(n9192), .ZN(n13372)
         );
  OR2_X1 U8623 ( .A1(n6546), .A2(n9173), .ZN(n9174) );
  OR2_X1 U8624 ( .A1(n9496), .A2(n9163), .ZN(n9167) );
  INV_X1 U8625 ( .A(n6910), .ZN(n10105) );
  NAND2_X1 U8626 ( .A1(n10261), .A2(n6651), .ZN(n10263) );
  NOR2_X1 U8627 ( .A1(n6923), .A2(n13393), .ZN(n13392) );
  NAND2_X1 U8628 ( .A1(n6922), .A2(n6924), .ZN(n11086) );
  INV_X1 U8629 ( .A(n13393), .ZN(n6922) );
  INV_X1 U8630 ( .A(n6913), .ZN(n14908) );
  NAND2_X1 U8631 ( .A1(n7099), .A2(n9574), .ZN(n13472) );
  NAND2_X1 U8632 ( .A1(n7099), .A2(n7097), .ZN(n13660) );
  NAND2_X1 U8633 ( .A1(n11872), .A2(n12168), .ZN(n9493) );
  NAND2_X1 U8634 ( .A1(n9573), .A2(n9572), .ZN(n13487) );
  NAND2_X1 U8635 ( .A1(n7169), .A2(n7172), .ZN(n13510) );
  AND2_X1 U8636 ( .A1(n9455), .A2(n9454), .ZN(n13542) );
  NAND2_X1 U8637 ( .A1(n7158), .A2(n9431), .ZN(n13566) );
  NAND2_X1 U8638 ( .A1(n13585), .A2(n13582), .ZN(n7158) );
  NAND2_X1 U8639 ( .A1(n7085), .A2(n7087), .ZN(n13570) );
  NAND2_X1 U8640 ( .A1(n7086), .A2(n6574), .ZN(n7085) );
  NAND2_X1 U8641 ( .A1(n9562), .A2(n9561), .ZN(n13621) );
  NAND2_X1 U8642 ( .A1(n7105), .A2(n9557), .ZN(n11690) );
  OR2_X1 U8643 ( .A1(n11570), .A2(n9556), .ZN(n7105) );
  NAND2_X1 U8644 ( .A1(n7093), .A2(n9551), .ZN(n11304) );
  NAND2_X1 U8645 ( .A1(n7174), .A2(n9294), .ZN(n11266) );
  CLKBUF_X1 U8646 ( .A(n12068), .Z(n6703) );
  NAND2_X1 U8647 ( .A1(n7091), .A2(n9546), .ZN(n10713) );
  OR2_X1 U8648 ( .A1(n9835), .A2(n6790), .ZN(n9260) );
  NAND2_X1 U8649 ( .A1(n10845), .A2(n9238), .ZN(n10979) );
  NAND2_X1 U8650 ( .A1(n10236), .A2(n9540), .ZN(n10658) );
  NAND2_X1 U8651 ( .A1(n7070), .A2(n9537), .ZN(n10073) );
  OR2_X1 U8652 ( .A1(n12247), .A2(n9536), .ZN(n7070) );
  OR2_X1 U8653 ( .A1(n14947), .A2(n10615), .ZN(n13610) );
  OR2_X1 U8654 ( .A1(n14947), .A2(n7536), .ZN(n14939) );
  NAND2_X1 U8655 ( .A1(n9300), .A2(n9299), .ZN(n12081) );
  INV_X1 U8656 ( .A(n12166), .ZN(n12165) );
  OAI21_X1 U8657 ( .B1(n13653), .B2(n13730), .A(n7111), .ZN(n13740) );
  AND2_X1 U8658 ( .A1(n13652), .A2(n13654), .ZN(n7111) );
  AND2_X1 U8659 ( .A1(n13651), .A2(n7538), .ZN(n13652) );
  OR2_X1 U8660 ( .A1(n13695), .A2(n13694), .ZN(n13751) );
  AND2_X1 U8661 ( .A1(n9433), .A2(n9432), .ZN(n13755) );
  INV_X1 U8662 ( .A(n12092), .ZN(n9580) );
  AND2_X1 U8663 ( .A1(n11481), .A2(n9602), .ZN(n14953) );
  NAND2_X1 U8664 ( .A1(n13771), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9147) );
  NAND2_X1 U8665 ( .A1(n9597), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9158) );
  NAND2_X1 U8666 ( .A1(n9389), .A2(n9388), .ZN(n9404) );
  INV_X1 U8667 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n9834) );
  INV_X1 U8668 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n9798) );
  INV_X1 U8669 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n9801) );
  INV_X1 U8670 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n9795) );
  INV_X1 U8671 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n15480) );
  OAI211_X1 U8672 ( .C1(P2_IR_REG_31__SCAN_IN), .C2(P2_IR_REG_1__SCAN_IN), .A(
        n9179), .B(n6925), .ZN(n9860) );
  NAND2_X1 U8673 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n6607), .ZN(n6925) );
  NAND2_X1 U8674 ( .A1(n7903), .A2(n7902), .ZN(n14680) );
  INV_X1 U8675 ( .A(n11374), .ZN(n6887) );
  NAND2_X1 U8676 ( .A1(n6886), .A2(n6885), .ZN(n11375) );
  NAND2_X1 U8677 ( .A1(n13877), .A2(n10370), .ZN(n10373) );
  NAND2_X1 U8678 ( .A1(n7341), .A2(n7345), .ZN(n13799) );
  OR2_X1 U8679 ( .A1(n13840), .A2(n7347), .ZN(n7341) );
  INV_X1 U8680 ( .A(n7352), .ZN(n11985) );
  OAI21_X1 U8681 ( .B1(n13848), .B2(n7355), .A(n7353), .ZN(n7352) );
  OR2_X1 U8682 ( .A1(n7360), .A2(n7356), .ZN(n7355) );
  INV_X1 U8683 ( .A(n7354), .ZN(n7353) );
  NAND2_X1 U8684 ( .A1(n11156), .A2(n11155), .ZN(n11158) );
  INV_X1 U8685 ( .A(n14792), .ZN(n13807) );
  NAND2_X1 U8686 ( .A1(n13855), .A2(n11930), .ZN(n13814) );
  NAND2_X1 U8687 ( .A1(n13797), .A2(n11923), .ZN(n13857) );
  NAND2_X1 U8688 ( .A1(n11544), .A2(n11543), .ZN(n11547) );
  NAND2_X1 U8689 ( .A1(n7856), .A2(n7855), .ZN(n11555) );
  OAI22_X1 U8690 ( .A1(n9797), .A2(n7711), .B1(n7727), .B2(n9754), .ZN(n6948)
         );
  INV_X1 U8691 ( .A(n7733), .ZN(n13885) );
  AND2_X1 U8692 ( .A1(n13818), .A2(n14247), .ZN(n14665) );
  NAND2_X1 U8693 ( .A1(n13839), .A2(n11909), .ZN(n13889) );
  INV_X1 U8694 ( .A(n14674), .ZN(n13880) );
  NAND2_X1 U8695 ( .A1(n6896), .A2(n6895), .ZN(n6894) );
  OAI21_X1 U8696 ( .B1(n6896), .B2(n13898), .A(n6890), .ZN(n6889) );
  NAND2_X1 U8697 ( .A1(n6896), .A2(n6891), .ZN(n6890) );
  NAND2_X1 U8698 ( .A1(n6895), .A2(n6899), .ZN(n6891) );
  AND2_X1 U8699 ( .A1(n10378), .A2(n11477), .ZN(n14684) );
  NAND2_X1 U8700 ( .A1(n6687), .A2(n6565), .ZN(n6694) );
  AND2_X1 U8701 ( .A1(n7036), .A2(n7042), .ZN(n7034) );
  INV_X1 U8702 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n10032) );
  INV_X1 U8703 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n10028) );
  INV_X1 U8704 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n10030) );
  AND2_X1 U8705 ( .A1(n14108), .A2(n14107), .ZN(n14296) );
  OAI21_X1 U8706 ( .B1(n14172), .B2(n14174), .A(n8192), .ZN(n14159) );
  NAND2_X1 U8707 ( .A1(n6953), .A2(n6959), .ZN(n14157) );
  NAND2_X1 U8708 ( .A1(n14172), .A2(n8192), .ZN(n6953) );
  NAND2_X1 U8709 ( .A1(n14173), .A2(n7528), .ZN(n14156) );
  NAND2_X1 U8710 ( .A1(n14224), .A2(n8011), .ZN(n14204) );
  NAND2_X1 U8711 ( .A1(n6944), .A2(n8342), .ZN(n14206) );
  OR2_X1 U8712 ( .A1(n14252), .A2(n14251), .ZN(n14354) );
  NAND2_X1 U8713 ( .A1(n11749), .A2(n7228), .ZN(n14279) );
  OAI21_X1 U8714 ( .B1(n6690), .B2(n7526), .A(n7524), .ZN(n14263) );
  NAND2_X1 U8715 ( .A1(n11754), .A2(n11753), .ZN(n11752) );
  NAND2_X1 U8716 ( .A1(n6690), .A2(n7937), .ZN(n11754) );
  NAND2_X1 U8717 ( .A1(n7926), .A2(n7925), .ZN(n14373) );
  NAND2_X1 U8718 ( .A1(n11459), .A2(n7224), .ZN(n6928) );
  NAND2_X1 U8719 ( .A1(n11352), .A2(n7898), .ZN(n11629) );
  NAND2_X1 U8720 ( .A1(n11459), .A2(n11464), .ZN(n7223) );
  NAND2_X1 U8721 ( .A1(n11016), .A2(n8178), .ZN(n11185) );
  AND2_X1 U8722 ( .A1(n14256), .A2(n14803), .ZN(n14235) );
  NAND2_X1 U8723 ( .A1(n10592), .A2(n8175), .ZN(n10807) );
  INV_X1 U8724 ( .A(n14284), .ZN(n14261) );
  AND2_X1 U8725 ( .A1(n14256), .A2(n14061), .ZN(n14284) );
  INV_X1 U8726 ( .A(n8454), .ZN(n14390) );
  NOR2_X1 U8727 ( .A1(n12605), .A2(n14761), .ZN(n6700) );
  NAND2_X1 U8728 ( .A1(n11816), .A2(n8418), .ZN(n8095) );
  OR3_X1 U8729 ( .A1(n14333), .A2(n14332), .A3(n14331), .ZN(n14412) );
  NAND2_X1 U8730 ( .A1(n8014), .A2(n8013), .ZN(n14415) );
  NAND2_X1 U8731 ( .A1(n7869), .A2(n7868), .ZN(n11599) );
  AND2_X1 U8732 ( .A1(n9914), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9780) );
  NAND2_X1 U8733 ( .A1(n8130), .A2(n7640), .ZN(n13776) );
  XNOR2_X1 U8734 ( .A(n8043), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n14438) );
  INV_X1 U8735 ( .A(n8152), .ZN(n14439) );
  NAND2_X1 U8736 ( .A1(n8140), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8145) );
  INV_X1 U8737 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n10070) );
  INV_X1 U8738 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n15281) );
  INV_X1 U8739 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n9794) );
  INV_X1 U8740 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n9773) );
  OAI21_X1 U8741 ( .B1(n7569), .B2(n7571), .A(n7380), .ZN(n7770) );
  INV_X1 U8742 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n9772) );
  NAND2_X1 U8743 ( .A1(n7750), .A2(n7749), .ZN(n7748) );
  OR2_X1 U8744 ( .A1(n7750), .A2(n7749), .ZN(n6689) );
  NAND2_X1 U8745 ( .A1(n7569), .A2(n7568), .ZN(n7750) );
  INV_X1 U8746 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n9768) );
  NAND2_X1 U8747 ( .A1(n7682), .A2(n6745), .ZN(n9800) );
  NAND2_X1 U8748 ( .A1(n6746), .A2(n7558), .ZN(n6745) );
  NAND2_X1 U8749 ( .A1(n15531), .A2(n15532), .ZN(n14492) );
  NOR2_X1 U8750 ( .A1(n15527), .A2(n14498), .ZN(n15520) );
  XNOR2_X1 U8751 ( .A(n14506), .B(n7284), .ZN(n14557) );
  INV_X1 U8752 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n7284) );
  XNOR2_X1 U8753 ( .A(n14511), .B(n7282), .ZN(n15525) );
  OAI21_X1 U8754 ( .B1(n14526), .B2(n7279), .A(n6568), .ZN(n14701) );
  NAND2_X1 U8755 ( .A1(n6697), .A2(n6562), .ZN(n7279) );
  NAND2_X1 U8756 ( .A1(n14704), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n7297) );
  NOR2_X1 U8757 ( .A1(n14708), .A2(n7295), .ZN(n7294) );
  INV_X1 U8758 ( .A(n7297), .ZN(n7295) );
  AND2_X1 U8759 ( .A1(n14541), .A2(n14540), .ZN(n14710) );
  AND2_X1 U8760 ( .A1(n14545), .A2(n14544), .ZN(n14564) );
  OAI211_X1 U8761 ( .C1(n6735), .C2(n6732), .A(n6728), .B(n6726), .ZN(n12870)
         );
  OAI21_X1 U8762 ( .B1(n12375), .B2(n13188), .A(n9111), .ZN(n9112) );
  NAND2_X1 U8763 ( .A1(n7121), .A2(n13326), .ZN(n7118) );
  NAND2_X1 U8764 ( .A1(n6920), .A2(n6915), .ZN(n13414) );
  NAND2_X1 U8765 ( .A1(n13412), .A2(n12613), .ZN(n6920) );
  NAND2_X1 U8766 ( .A1(n6919), .A2(n6916), .ZN(n6915) );
  AOI21_X1 U8767 ( .B1(n13655), .B2(n15007), .A(n6664), .ZN(n9618) );
  AND2_X1 U8768 ( .A1(n6650), .A2(n9622), .ZN(n9623) );
  OAI21_X1 U8769 ( .B1(n8488), .B2(n14809), .A(n6714), .ZN(n8486) );
  OR2_X1 U8770 ( .A1(n14811), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n6714) );
  AND2_X1 U8771 ( .A1(n7539), .A2(n8505), .ZN(n8506) );
  OAI21_X1 U8772 ( .B1(n8488), .B2(n14804), .A(n6715), .ZN(n8489) );
  OR2_X1 U8773 ( .A1(n14806), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n6715) );
  NAND2_X1 U8774 ( .A1(n7290), .A2(n14521), .ZN(n14560) );
  NOR2_X1 U8775 ( .A1(n14697), .A2(n14696), .ZN(n14695) );
  NOR2_X1 U8776 ( .A1(n14526), .A2(n14693), .ZN(n14697) );
  OAI21_X1 U8777 ( .B1(n14573), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n7275), .ZN(
        n7274) );
  AND2_X1 U8778 ( .A1(n8179), .A2(n8178), .ZN(n6554) );
  AND2_X1 U8779 ( .A1(n14981), .A2(n7191), .ZN(n6555) );
  INV_X1 U8780 ( .A(n7002), .ZN(n7001) );
  NAND2_X1 U8781 ( .A1(n12476), .A2(n7003), .ZN(n7002) );
  INV_X2 U8782 ( .A(n10429), .ZN(n13603) );
  INV_X2 U8783 ( .A(n13603), .ZN(n10574) );
  INV_X1 U8784 ( .A(n13583), .ZN(n7086) );
  OR2_X1 U8785 ( .A1(n12056), .A2(n12055), .ZN(n6556) );
  NAND2_X1 U8786 ( .A1(n7689), .A2(n10178), .ZN(n8434) );
  INV_X1 U8787 ( .A(n14174), .ZN(n6961) );
  INV_X1 U8788 ( .A(n8448), .ZN(n8474) );
  INV_X1 U8789 ( .A(n7571), .ZN(n7749) );
  NAND2_X1 U8790 ( .A1(n9757), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n6557) );
  NOR2_X1 U8791 ( .A1(n12739), .A2(n15193), .ZN(n6558) );
  AOI21_X1 U8792 ( .B1(n7159), .B2(n7160), .A(n7157), .ZN(n7156) );
  OR2_X1 U8793 ( .A1(n12106), .A2(n12107), .ZN(n6559) );
  NOR2_X1 U8794 ( .A1(n14561), .A2(P2_ADDR_REG_10__SCAN_IN), .ZN(n6560) );
  INV_X1 U8795 ( .A(n12479), .ZN(n6999) );
  OR2_X1 U8796 ( .A1(n11367), .A2(n11366), .ZN(n6561) );
  OR2_X1 U8797 ( .A1(n14696), .A2(P2_ADDR_REG_12__SCAN_IN), .ZN(n6562) );
  AND2_X1 U8798 ( .A1(n12447), .A2(n12448), .ZN(n12384) );
  INV_X1 U8799 ( .A(n12384), .ZN(n6994) );
  AND2_X1 U8800 ( .A1(n11460), .A2(n7863), .ZN(n11279) );
  INV_X1 U8801 ( .A(n11279), .ZN(n7512) );
  AND2_X1 U8802 ( .A1(n13661), .A2(n13352), .ZN(n6563) );
  INV_X1 U8803 ( .A(n8301), .ZN(n7057) );
  AND2_X1 U8804 ( .A1(n13681), .A2(n13299), .ZN(n6564) );
  AND2_X1 U8805 ( .A1(n7036), .A2(n6646), .ZN(n6565) );
  AND2_X1 U8806 ( .A1(n8269), .A2(n7065), .ZN(n6566) );
  INV_X1 U8807 ( .A(n7496), .ZN(n7495) );
  OAI21_X1 U8808 ( .B1(n7500), .B2(n7498), .A(n7497), .ZN(n7496) );
  INV_X1 U8809 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n9405) );
  AND2_X1 U8810 ( .A1(n7416), .A2(n6657), .ZN(n6567) );
  INV_X1 U8811 ( .A(n11621), .ZN(n6996) );
  NAND2_X1 U8812 ( .A1(n14696), .A2(P2_ADDR_REG_12__SCAN_IN), .ZN(n6568) );
  AND2_X1 U8813 ( .A1(n7781), .A2(n10589), .ZN(n10543) );
  AND2_X1 U8814 ( .A1(n7506), .A2(n7372), .ZN(n6569) );
  INV_X1 U8815 ( .A(n14061), .ZN(n7373) );
  NAND2_X1 U8816 ( .A1(n7837), .A2(n7836), .ZN(n11373) );
  INV_X1 U8817 ( .A(n11373), .ZN(n7012) );
  INV_X1 U8818 ( .A(n12060), .ZN(n7191) );
  OR2_X1 U8819 ( .A1(n7245), .A2(n6676), .ZN(n6570) );
  NAND2_X4 U8820 ( .A1(n10036), .A2(n8149), .ZN(n11149) );
  OR2_X1 U8821 ( .A1(n10883), .A2(n10866), .ZN(n6571) );
  OR2_X1 U8822 ( .A1(n7444), .A2(n8697), .ZN(n6572) );
  XNOR2_X1 U8823 ( .A(n13287), .B(n13283), .ZN(n6573) );
  INV_X1 U8824 ( .A(n13029), .ZN(n13023) );
  OR2_X1 U8825 ( .A1(n13703), .A2(n13356), .ZN(n6574) );
  INV_X1 U8826 ( .A(n12275), .ZN(n7157) );
  AND2_X1 U8827 ( .A1(n12825), .A2(n12824), .ZN(n6879) );
  AND2_X1 U8828 ( .A1(n6888), .A2(n11155), .ZN(n6575) );
  OR2_X1 U8829 ( .A1(n7425), .A2(n8721), .ZN(n6576) );
  NAND2_X1 U8830 ( .A1(n12548), .A2(n12943), .ZN(n6577) );
  NAND2_X1 U8831 ( .A1(n13661), .A2(n9501), .ZN(n6578) );
  NAND4_X1 U8832 ( .A1(n11290), .A2(n9657), .A3(n11106), .A4(n9655), .ZN(n6579) );
  AND4_X1 U8833 ( .A1(n9600), .A2(n9589), .A3(n9145), .A4(n9595), .ZN(n6580)
         );
  OR2_X1 U8834 ( .A1(n9797), .A2(n9177), .ZN(n6581) );
  INV_X1 U8835 ( .A(n11753), .ZN(n7526) );
  AND2_X1 U8836 ( .A1(n13479), .A2(n6978), .ZN(n6582) );
  AND2_X1 U8837 ( .A1(n14160), .A2(n14140), .ZN(n6583) );
  NAND2_X1 U8838 ( .A1(n11897), .A2(n11896), .ZN(n6584) );
  OR2_X1 U8839 ( .A1(n14095), .A2(n14106), .ZN(n6585) );
  INV_X1 U8840 ( .A(n6848), .ZN(n6847) );
  NAND2_X1 U8841 ( .A1(n6853), .A2(n6849), .ZN(n6848) );
  INV_X1 U8842 ( .A(n13471), .ZN(n7184) );
  NAND2_X1 U8843 ( .A1(n9379), .A2(n9378), .ZN(n12125) );
  OR2_X1 U8844 ( .A1(n7470), .A2(n7471), .ZN(n6586) );
  INV_X1 U8845 ( .A(n12413), .ZN(n7000) );
  XNOR2_X1 U8846 ( .A(n13650), .B(n13351), .ZN(n13433) );
  INV_X1 U8847 ( .A(n13433), .ZN(n13434) );
  AND2_X1 U8848 ( .A1(n12568), .A2(n14620), .ZN(n6587) );
  AND2_X1 U8849 ( .A1(n12867), .A2(n14592), .ZN(n6588) );
  AND2_X1 U8850 ( .A1(n14173), .A2(n8051), .ZN(n14155) );
  NAND2_X1 U8851 ( .A1(n13430), .A2(n9514), .ZN(n12279) );
  NAND2_X1 U8852 ( .A1(n8132), .A2(n8131), .ZN(n8379) );
  INV_X1 U8853 ( .A(n8379), .ZN(n7018) );
  AND2_X1 U8854 ( .A1(n12742), .A2(n11065), .ZN(n6589) );
  AND2_X1 U8855 ( .A1(n6787), .A2(n6789), .ZN(n6590) );
  AND3_X1 U8856 ( .A1(n9166), .A2(n9165), .A3(n9168), .ZN(n6591) );
  NAND2_X1 U8857 ( .A1(n8065), .A2(n8064), .ZN(n14148) );
  INV_X1 U8858 ( .A(n8355), .ZN(n6815) );
  AND2_X1 U8859 ( .A1(n9238), .A2(n7194), .ZN(n6592) );
  NAND2_X1 U8860 ( .A1(n9485), .A2(n9484), .ZN(n13670) );
  INV_X1 U8861 ( .A(n12106), .ZN(n7470) );
  AND2_X1 U8862 ( .A1(n9689), .A2(n12733), .ZN(n6593) );
  AND2_X1 U8863 ( .A1(n12074), .A2(n12073), .ZN(n6594) );
  NAND2_X1 U8864 ( .A1(n8031), .A2(n8030), .ZN(n14199) );
  INV_X1 U8865 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n13195) );
  NAND2_X1 U8866 ( .A1(n9424), .A2(n9423), .ZN(n13703) );
  INV_X1 U8867 ( .A(n7173), .ZN(n7172) );
  NOR2_X1 U8868 ( .A1(n13542), .A2(n13354), .ZN(n7173) );
  NAND2_X1 U8869 ( .A1(n14211), .A2(n7024), .ZN(n7027) );
  AND2_X1 U8870 ( .A1(n13755), .A2(n13355), .ZN(n6595) );
  INV_X1 U8871 ( .A(n14100), .ZN(n14104) );
  NAND2_X1 U8872 ( .A1(n8479), .A2(n8105), .ZN(n14100) );
  AND2_X1 U8873 ( .A1(n8328), .A2(n8331), .ZN(n6596) );
  AND2_X1 U8874 ( .A1(n7493), .A2(n7491), .ZN(n6597) );
  AND2_X1 U8875 ( .A1(n8478), .A2(n6716), .ZN(n6598) );
  NAND2_X1 U8876 ( .A1(n11364), .A2(n11365), .ZN(n6599) );
  INV_X1 U8877 ( .A(n7083), .ZN(n7082) );
  NAND2_X1 U8878 ( .A1(n9567), .A2(n6574), .ZN(n7083) );
  AND2_X1 U8879 ( .A1(n11545), .A2(n11543), .ZN(n6600) );
  AND2_X1 U8880 ( .A1(n9308), .A2(n9294), .ZN(n6601) );
  AND2_X1 U8881 ( .A1(n6885), .A2(n6887), .ZN(n6602) );
  INV_X1 U8882 ( .A(n7101), .ZN(n7100) );
  OR2_X1 U8883 ( .A1(n9575), .A2(n7102), .ZN(n7101) );
  NAND2_X1 U8884 ( .A1(n7204), .A2(n7203), .ZN(n6603) );
  AND2_X1 U8885 ( .A1(n6561), .A2(n6575), .ZN(n6604) );
  NAND2_X1 U8886 ( .A1(n12105), .A2(n9334), .ZN(n6605) );
  INV_X1 U8887 ( .A(n6899), .ZN(n6898) );
  NAND2_X1 U8888 ( .A1(n7363), .A2(n6900), .ZN(n6899) );
  NOR2_X1 U8889 ( .A1(n7469), .A2(n6769), .ZN(n6606) );
  AND2_X1 U8890 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n6607) );
  NOR2_X1 U8891 ( .A1(n13690), .A2(n13264), .ZN(n6608) );
  NOR2_X1 U8892 ( .A1(n14358), .A2(n14250), .ZN(n6609) );
  NOR2_X1 U8893 ( .A1(n11373), .A2(n11550), .ZN(n6610) );
  NOR2_X1 U8894 ( .A1(n11736), .A2(n14669), .ZN(n6611) );
  INV_X1 U8895 ( .A(n12450), .ZN(n6989) );
  INV_X1 U8896 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n8210) );
  OR2_X1 U8897 ( .A1(n14445), .A2(n14446), .ZN(n6612) );
  INV_X1 U8898 ( .A(n7088), .ZN(n7087) );
  NOR2_X1 U8899 ( .A1(n13591), .A2(n12143), .ZN(n7088) );
  AND2_X1 U8900 ( .A1(n6820), .A2(n6818), .ZN(n6613) );
  AND2_X1 U8901 ( .A1(n9175), .A2(n9176), .ZN(n6614) );
  AND2_X1 U8902 ( .A1(n12047), .A2(n12046), .ZN(n6615) );
  AND2_X1 U8903 ( .A1(n6982), .A2(n6985), .ZN(n6616) );
  AND2_X1 U8904 ( .A1(n7585), .A2(n9785), .ZN(n6617) );
  NOR2_X1 U8905 ( .A1(n13221), .A2(n13220), .ZN(n6618) );
  INV_X1 U8906 ( .A(n12070), .ZN(n7484) );
  INV_X1 U8907 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n7074) );
  INV_X1 U8908 ( .A(n7529), .ZN(n7528) );
  NAND2_X1 U8909 ( .A1(n8061), .A2(n8051), .ZN(n7529) );
  AND2_X1 U8910 ( .A1(n9838), .A2(P2_DATAO_REG_9__SCAN_IN), .ZN(n6619) );
  NAND2_X1 U8911 ( .A1(n8210), .A2(n7657), .ZN(n7531) );
  NAND2_X1 U8912 ( .A1(n11978), .A2(n11977), .ZN(n6620) );
  INV_X1 U8913 ( .A(n6812), .ZN(n6811) );
  NAND2_X1 U8914 ( .A1(n8358), .A2(n6813), .ZN(n6812) );
  NAND2_X1 U8915 ( .A1(n9768), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n8612) );
  AND2_X1 U8916 ( .A1(n7495), .A2(n7499), .ZN(n6621) );
  AND2_X1 U8917 ( .A1(n7530), .A2(n7661), .ZN(n6622) );
  INV_X1 U8918 ( .A(n12899), .ZN(n12902) );
  NAND2_X1 U8919 ( .A1(n12554), .A2(n12553), .ZN(n12899) );
  NAND2_X1 U8920 ( .A1(n8962), .A2(n7435), .ZN(n6623) );
  AND2_X1 U8921 ( .A1(n8521), .A2(n7449), .ZN(n6624) );
  INV_X1 U8922 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n7372) );
  OR2_X1 U8923 ( .A1(n14203), .A2(n7516), .ZN(n6625) );
  OR2_X1 U8924 ( .A1(n12574), .A2(n6587), .ZN(n6626) );
  INV_X1 U8925 ( .A(n6905), .ZN(n6904) );
  NAND2_X1 U8926 ( .A1(n9057), .A2(n12925), .ZN(n12542) );
  NAND2_X1 U8927 ( .A1(n12065), .A2(n12064), .ZN(n7488) );
  INV_X1 U8928 ( .A(n7186), .ZN(n7185) );
  NAND2_X1 U8929 ( .A1(n6578), .A2(n12279), .ZN(n7186) );
  INV_X1 U8930 ( .A(n12266), .ZN(n11805) );
  AND2_X1 U8931 ( .A1(n8409), .A2(n8408), .ZN(n6627) );
  NAND2_X1 U8932 ( .A1(n12170), .A2(n12169), .ZN(n13650) );
  INV_X1 U8933 ( .A(n13650), .ZN(n6975) );
  AND2_X1 U8934 ( .A1(n7257), .A2(n7256), .ZN(n6628) );
  INV_X1 U8935 ( .A(n8439), .ZN(n10812) );
  OR2_X1 U8936 ( .A1(n12078), .A2(n6594), .ZN(n6629) );
  OR2_X1 U8937 ( .A1(n14447), .A2(n14448), .ZN(n6630) );
  AND2_X1 U8938 ( .A1(n7133), .A2(n7137), .ZN(n6631) );
  AND2_X1 U8939 ( .A1(n8730), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n6632) );
  AND2_X1 U8940 ( .A1(n14521), .A2(n7289), .ZN(n6633) );
  AND2_X1 U8941 ( .A1(n6970), .A2(n13591), .ZN(n6634) );
  AND2_X1 U8942 ( .A1(n8962), .A2(n7439), .ZN(n6635) );
  AND2_X1 U8943 ( .A1(n6629), .A2(n12083), .ZN(n6636) );
  AND2_X1 U8944 ( .A1(n7488), .A2(n12070), .ZN(n6637) );
  AND2_X1 U8945 ( .A1(n9053), .A2(n12518), .ZN(n6638) );
  AND2_X1 U8946 ( .A1(n6586), .A2(n12114), .ZN(n6639) );
  NOR2_X1 U8947 ( .A1(n13222), .A2(n7136), .ZN(n7135) );
  AND2_X1 U8948 ( .A1(n12570), .A2(n12569), .ZN(n6640) );
  AND2_X1 U8949 ( .A1(n12132), .A2(n12131), .ZN(n6641) );
  AND2_X1 U8950 ( .A1(n7524), .A2(n8185), .ZN(n6642) );
  INV_X1 U8951 ( .A(n7042), .ZN(n7041) );
  AND2_X1 U8952 ( .A1(n9146), .A2(n6580), .ZN(n6643) );
  NOR2_X1 U8953 ( .A1(n7531), .A2(P1_IR_REG_28__SCAN_IN), .ZN(n7530) );
  AND2_X1 U8954 ( .A1(n7534), .A2(n8324), .ZN(n6644) );
  AND2_X1 U8955 ( .A1(n7507), .A2(n7878), .ZN(n6645) );
  OR2_X1 U8956 ( .A1(n7045), .A2(n8410), .ZN(n6646) );
  AND2_X1 U8957 ( .A1(n14262), .A2(n8184), .ZN(n7228) );
  OR2_X1 U8958 ( .A1(n7084), .A2(n7081), .ZN(n7080) );
  INV_X1 U8959 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n9157) );
  OR2_X1 U8960 ( .A1(n12144), .A2(n12145), .ZN(n7501) );
  OR2_X1 U8961 ( .A1(n7467), .A2(n6615), .ZN(n6647) );
  NAND2_X1 U8962 ( .A1(n8378), .A2(n7055), .ZN(n6648) );
  INV_X4 U8963 ( .A(n11940), .ZN(n11980) );
  INV_X1 U8964 ( .A(n13463), .ZN(n7188) );
  NOR2_X2 U8965 ( .A1(n8558), .A2(n8557), .ZN(n10892) );
  INV_X1 U8966 ( .A(n12147), .ZN(n7498) );
  NAND2_X1 U8967 ( .A1(n6936), .A2(n6937), .ZN(n14240) );
  INV_X1 U8968 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6713) );
  XOR2_X1 U8969 ( .A(n13542), .B(n13282), .Z(n6649) );
  NAND2_X1 U8970 ( .A1(n7223), .A2(n8182), .ZN(n11350) );
  NAND2_X1 U8971 ( .A1(n6928), .A2(n7222), .ZN(n11632) );
  OR2_X1 U8972 ( .A1(n9620), .A2(n14327), .ZN(n6650) );
  OR2_X1 U8973 ( .A1(n10262), .A2(n11010), .ZN(n6651) );
  AND2_X1 U8974 ( .A1(n14521), .A2(n7288), .ZN(n6652) );
  NOR2_X1 U8975 ( .A1(n12767), .A2(n12768), .ZN(n6653) );
  AND2_X1 U8976 ( .A1(n7104), .A2(n7106), .ZN(n6654) );
  INV_X1 U8977 ( .A(n6860), .ZN(n6859) );
  INV_X1 U8978 ( .A(n7011), .ZN(n11679) );
  NOR2_X1 U8979 ( .A1(n11635), .A2(n14680), .ZN(n7011) );
  NAND2_X1 U8980 ( .A1(n11848), .A2(n6970), .ZN(n6973) );
  INV_X1 U8981 ( .A(n13287), .ZN(n13658) );
  NAND2_X1 U8982 ( .A1(n9504), .A2(n9503), .ZN(n13287) );
  NOR2_X1 U8983 ( .A1(n14703), .A2(n14704), .ZN(n6655) );
  AND2_X1 U8984 ( .A1(n7321), .A2(n7319), .ZN(n6656) );
  AND2_X1 U8985 ( .A1(n7551), .A2(n7535), .ZN(n6657) );
  OR2_X1 U8986 ( .A1(n11908), .A2(n11907), .ZN(n11909) );
  AND2_X1 U8987 ( .A1(n8341), .A2(n8342), .ZN(n14223) );
  INV_X1 U8988 ( .A(n14223), .ZN(n7229) );
  OR2_X1 U8989 ( .A1(n13147), .A2(n13188), .ZN(n6658) );
  OR2_X1 U8990 ( .A1(n13147), .A2(n13138), .ZN(n6659) );
  NOR2_X1 U8991 ( .A1(n10881), .A2(n12324), .ZN(n6857) );
  AND2_X1 U8992 ( .A1(n9335), .A2(n9334), .ZN(n6660) );
  INV_X1 U8993 ( .A(n7331), .ZN(n8763) );
  AND2_X1 U8994 ( .A1(n7290), .A2(n6652), .ZN(n6661) );
  AND2_X1 U8995 ( .A1(n6883), .A2(n6584), .ZN(n6662) );
  INV_X1 U8996 ( .A(n12110), .ZN(n6968) );
  OR2_X1 U8997 ( .A1(n9502), .A2(n13769), .ZN(n6663) );
  INV_X1 U8998 ( .A(n6703), .ZN(n6979) );
  INV_X1 U8999 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n7155) );
  NAND2_X1 U9000 ( .A1(n7541), .A2(n9144), .ZN(n9583) );
  NAND2_X1 U9001 ( .A1(n10539), .A2(n10543), .ZN(n10538) );
  AND2_X1 U9002 ( .A1(n9579), .A2(n7536), .ZN(n10530) );
  AND2_X1 U9003 ( .A1(n15005), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6664) );
  INV_X1 U9004 ( .A(n8871), .ZN(n7268) );
  INV_X1 U9005 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n7150) );
  NAND2_X1 U9006 ( .A1(n9092), .A2(n9091), .ZN(n9625) );
  INV_X1 U9007 ( .A(n11460), .ZN(n7510) );
  NAND2_X1 U9008 ( .A1(n7473), .A2(n9144), .ZN(n9597) );
  NAND4_X1 U9009 ( .A1(n7371), .A2(n6569), .A3(n7649), .A4(n7743), .ZN(n7993)
         );
  AND2_X1 U9010 ( .A1(n6663), .A2(n13421), .ZN(n6665) );
  AND2_X1 U9011 ( .A1(n11016), .A2(n6554), .ZN(n6666) );
  OR2_X1 U9012 ( .A1(n11249), .A2(n10885), .ZN(n6667) );
  AND2_X1 U9013 ( .A1(n7339), .A2(n7337), .ZN(n6668) );
  INV_X1 U9014 ( .A(n7154), .ZN(n9376) );
  AND2_X1 U9015 ( .A1(n8108), .A2(SI_27_), .ZN(n6669) );
  INV_X1 U9016 ( .A(n7013), .ZN(n11189) );
  NOR2_X1 U9017 ( .A1(n11023), .A2(n11232), .ZN(n7013) );
  AND2_X1 U9018 ( .A1(n7209), .A2(n6571), .ZN(n6670) );
  AND2_X1 U9019 ( .A1(n11072), .A2(n8619), .ZN(n6671) );
  NAND2_X1 U9020 ( .A1(n11246), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n6672) );
  NAND2_X1 U9021 ( .A1(n7775), .A2(n7774), .ZN(n10767) );
  INV_X1 U9022 ( .A(n10767), .ZN(n7015) );
  AND2_X1 U9023 ( .A1(n10307), .A2(n10642), .ZN(n6673) );
  AND2_X1 U9024 ( .A1(n7249), .A2(n8999), .ZN(n6674) );
  AND2_X1 U9025 ( .A1(n15252), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n6675) );
  INV_X1 U9026 ( .A(n9014), .ZN(n7248) );
  NAND4_X1 U9027 ( .A1(n8546), .A2(n8545), .A3(n8544), .A4(n8543), .ZN(n15138)
         );
  INV_X1 U9028 ( .A(n14593), .ZN(n6733) );
  INV_X1 U9029 ( .A(n8173), .ZN(n7221) );
  INV_X1 U9030 ( .A(n12860), .ZN(n6737) );
  AND2_X1 U9031 ( .A1(n6674), .A2(n12359), .ZN(n6676) );
  NAND2_X1 U9032 ( .A1(n15332), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n6677) );
  INV_X1 U9033 ( .A(SI_1_), .ZN(n7389) );
  INV_X1 U9034 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n6740) );
  NOR2_X1 U9035 ( .A1(n12838), .A2(n12843), .ZN(n6678) );
  INV_X1 U9036 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n7287) );
  INV_X1 U9037 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n6696) );
  INV_X1 U9038 ( .A(SI_23_), .ZN(n7377) );
  INV_X1 U9039 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n7282) );
  OAI21_X2 U9040 ( .B1(n14175), .B2(n7529), .A(n7527), .ZN(n14138) );
  NAND2_X2 U9041 ( .A1(n7523), .A2(n7520), .ZN(n14242) );
  NAND2_X1 U9042 ( .A1(n11020), .A2(n7829), .ZN(n11184) );
  NAND2_X1 U9043 ( .A1(n10596), .A2(n7798), .ZN(n10813) );
  NOR2_X1 U9044 ( .A1(n14222), .A2(n14223), .ZN(n8010) );
  NAND2_X1 U9045 ( .A1(n6701), .A2(n6699), .ZN(n8241) );
  NAND2_X1 U9046 ( .A1(n14122), .A2(n8090), .ZN(n14101) );
  NAND2_X1 U9047 ( .A1(n6698), .A2(n11675), .ZN(n7938) );
  NAND2_X1 U9048 ( .A1(n11631), .A2(n7912), .ZN(n11674) );
  NAND2_X1 U9049 ( .A1(n6679), .A2(n6688), .ZN(n8261) );
  OAI21_X1 U9050 ( .B1(n7053), .B2(n7052), .A(n7054), .ZN(n8381) );
  NAND2_X1 U9051 ( .A1(n7030), .A2(n7028), .ZN(n8374) );
  AOI21_X1 U9052 ( .B1(n8276), .B2(n8278), .A(n6801), .ZN(n6800) );
  INV_X1 U9053 ( .A(n8411), .ZN(n6687) );
  OAI21_X1 U9054 ( .B1(n8264), .B2(n8263), .A(n8262), .ZN(n8266) );
  NAND2_X2 U9055 ( .A1(n8389), .A2(n8246), .ZN(n8340) );
  NAND3_X1 U9056 ( .A1(n7473), .A2(n9144), .A3(n9157), .ZN(n6680) );
  NAND2_X2 U9057 ( .A1(n6681), .A2(n9161), .ZN(n14934) );
  NAND2_X1 U9058 ( .A1(n7555), .A2(n7554), .ZN(n6683) );
  NAND2_X1 U9059 ( .A1(P1_ADDR_REG_19__SCAN_IN), .A2(n7556), .ZN(n6684) );
  OAI21_X2 U9060 ( .B1(n10575), .B2(n10576), .A(n10581), .ZN(n10771) );
  OAI21_X2 U9061 ( .B1(n13290), .B2(n13289), .A(n13239), .ZN(n13242) );
  OAI21_X2 U9062 ( .B1(n11142), .B2(n11141), .A(n11140), .ZN(n11400) );
  NAND2_X1 U9063 ( .A1(n9144), .A2(n7474), .ZN(n13771) );
  NAND2_X4 U9064 ( .A1(n9148), .A2(n9149), .ZN(n9496) );
  INV_X1 U9065 ( .A(n9146), .ZN(n7475) );
  NAND2_X2 U9066 ( .A1(n9167), .A2(n6591), .ZN(n13375) );
  NAND2_X1 U9067 ( .A1(n7132), .A2(n7135), .ZN(n7131) );
  NAND2_X1 U9068 ( .A1(n7113), .A2(n10136), .ZN(n10311) );
  NAND2_X1 U9069 ( .A1(n6686), .A2(n6685), .ZN(n10440) );
  NAND2_X1 U9070 ( .A1(n7802), .A2(n7801), .ZN(n9835) );
  NAND2_X1 U9071 ( .A1(n10783), .A2(n10935), .ZN(n7139) );
  NAND2_X1 U9072 ( .A1(n7562), .A2(SI_3_), .ZN(n7564) );
  NAND2_X1 U9073 ( .A1(n10776), .A2(n10775), .ZN(n10784) );
  INV_X1 U9074 ( .A(n10311), .ZN(n6686) );
  NAND2_X1 U9075 ( .A1(n10095), .A2(n10096), .ZN(n7113) );
  NAND2_X1 U9076 ( .A1(n10013), .A2(n10012), .ZN(n10094) );
  NAND2_X1 U9077 ( .A1(n7143), .A2(n7141), .ZN(n11427) );
  NAND2_X1 U9078 ( .A1(n13313), .A2(n13314), .ZN(n13312) );
  NAND2_X1 U9079 ( .A1(n11836), .A2(n11835), .ZN(n11838) );
  NAND2_X1 U9080 ( .A1(n11400), .A2(n11399), .ZN(n7143) );
  NAND2_X2 U9081 ( .A1(n9852), .A2(n13418), .ZN(n9841) );
  NAND2_X1 U9082 ( .A1(n13312), .A2(n13235), .ZN(n13290) );
  NAND2_X1 U9083 ( .A1(n11427), .A2(n11426), .ZN(n11660) );
  XNOR2_X1 U9084 ( .A(n14934), .B(n10428), .ZN(n10090) );
  NAND2_X1 U9085 ( .A1(n10471), .A2(n10441), .ZN(n10575) );
  NAND2_X1 U9086 ( .A1(n10994), .A2(n10993), .ZN(n11142) );
  NAND3_X1 U9087 ( .A1(n8254), .A2(n8255), .A3(n8253), .ZN(n6688) );
  OAI22_X1 U9088 ( .A1(n8268), .A2(n6566), .B1(n8269), .B2(n7065), .ZN(n8272)
         );
  NAND2_X1 U9089 ( .A1(n6823), .A2(n6824), .ZN(n8296) );
  NAND2_X1 U9090 ( .A1(n8375), .A2(n6648), .ZN(n7052) );
  OAI22_X1 U9091 ( .A1(n6802), .A2(n6800), .B1(n8283), .B2(n7048), .ZN(n8286)
         );
  NAND2_X1 U9092 ( .A1(n10441), .A2(n10434), .ZN(n10469) );
  NAND2_X1 U9093 ( .A1(n7140), .A2(n7138), .ZN(n10994) );
  OAI22_X1 U9094 ( .A1(n7062), .A2(n7061), .B1(n7064), .B2(n8362), .ZN(n8364)
         );
  AOI21_X1 U9095 ( .B1(n7033), .B2(n8369), .A(n7032), .ZN(n7031) );
  INV_X1 U9096 ( .A(n7038), .ZN(n7037) );
  NAND2_X1 U9097 ( .A1(n6689), .A2(n7748), .ZN(n9796) );
  XNOR2_X2 U9098 ( .A(n6881), .B(n7656), .ZN(n8158) );
  NAND2_X1 U9099 ( .A1(n12603), .A2(n14803), .ZN(n6701) );
  NAND2_X1 U9100 ( .A1(n7797), .A2(n10590), .ZN(n10596) );
  NAND2_X1 U9101 ( .A1(n8041), .A2(n8040), .ZN(n14175) );
  INV_X1 U9102 ( .A(n11674), .ZN(n6698) );
  XNOR2_X1 U9103 ( .A(n14514), .B(n14515), .ZN(n14558) );
  NOR2_X1 U9104 ( .A1(n14706), .A2(n7300), .ZN(n14541) );
  OAI21_X1 U9105 ( .B1(n6633), .B2(n6560), .A(n7285), .ZN(n14525) );
  INV_X1 U9106 ( .A(n14574), .ZN(n7275) );
  XNOR2_X1 U9107 ( .A(n7274), .B(n14575), .ZN(SUB_1596_U4) );
  NOR2_X1 U9108 ( .A1(n14711), .A2(n14542), .ZN(n14544) );
  NOR2_X1 U9109 ( .A1(n14565), .A2(n14546), .ZN(n14547) );
  NAND2_X1 U9110 ( .A1(n13080), .A2(n13139), .ZN(n6692) );
  NAND2_X1 U9111 ( .A1(n8725), .A2(n8724), .ZN(n8739) );
  NAND2_X1 U9112 ( .A1(n13083), .A2(n6659), .ZN(P3_U3487) );
  NAND2_X1 U9113 ( .A1(n13146), .A2(n6658), .ZN(P3_U3455) );
  INV_X1 U9114 ( .A(n8652), .ZN(n6705) );
  INV_X1 U9115 ( .A(n8465), .ZN(n8466) );
  NAND3_X1 U9116 ( .A1(n7035), .A2(n8469), .A3(n6694), .ZN(n8473) );
  NAND3_X1 U9117 ( .A1(n8450), .A2(n8451), .A3(n8452), .ZN(n6695) );
  NAND2_X1 U9118 ( .A1(n13323), .A2(n13325), .ZN(n13324) );
  OAI21_X1 U9119 ( .B1(SI_2_), .B2(n7559), .A(n7561), .ZN(n7707) );
  NOR2_X1 U9120 ( .A1(n14558), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n7276) );
  NOR2_X1 U9121 ( .A1(n14701), .A2(n14700), .ZN(n14531) );
  OR2_X1 U9122 ( .A1(n7816), .A2(n7815), .ZN(n7817) );
  AOI21_X2 U9123 ( .B1(n13297), .B2(n13296), .A(n6702), .ZN(n13338) );
  OAI22_X2 U9124 ( .A1(n13306), .A2(n13305), .B1(n13248), .B2(n13247), .ZN(
        n13297) );
  NAND2_X1 U9125 ( .A1(n7518), .A2(n7517), .ZN(n8493) );
  MUX2_X1 U9126 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n8241), .S(n14811), .Z(
        P1_U3557) );
  OAI21_X1 U9127 ( .B1(n12572), .B2(n12571), .A(n6640), .ZN(n12576) );
  AOI21_X4 U9128 ( .B1(n7271), .B2(n7270), .A(n6675), .ZN(n8943) );
  XNOR2_X1 U9129 ( .A(n9015), .B(n7248), .ZN(n13204) );
  NAND2_X1 U9130 ( .A1(n8964), .A2(n8963), .ZN(n7232) );
  NAND2_X1 U9131 ( .A1(n8979), .A2(n8980), .ZN(n8981) );
  NAND2_X1 U9132 ( .A1(n13812), .A2(n11937), .ZN(n13865) );
  NAND2_X1 U9133 ( .A1(n7344), .A2(n7342), .ZN(n13797) );
  NAND2_X1 U9134 ( .A1(n10478), .A2(n9648), .ZN(n10651) );
  NAND2_X1 U9135 ( .A1(n12652), .A2(n9714), .ZN(n12720) );
  INV_X4 U9136 ( .A(n10251), .ZN(n9644) );
  NAND2_X4 U9137 ( .A1(n7328), .A2(n6709), .ZN(n10251) );
  NAND2_X1 U9138 ( .A1(n6720), .A2(n6545), .ZN(n9080) );
  NAND2_X1 U9139 ( .A1(n7326), .A2(n7324), .ZN(n9673) );
  NAND2_X2 U9140 ( .A1(n13338), .A2(n13337), .ZN(n13336) );
  INV_X2 U9141 ( .A(n12021), .ZN(n10946) );
  NAND2_X1 U9142 ( .A1(n7590), .A2(n7589), .ZN(n7865) );
  NAND2_X1 U9143 ( .A1(n7785), .A2(n7784), .ZN(n7787) );
  NAND3_X1 U9144 ( .A1(n15481), .A2(n7553), .A3(P2_ADDR_REG_19__SCAN_IN), .ZN(
        n7556) );
  NAND2_X1 U9145 ( .A1(n7375), .A2(n7376), .ZN(n7627) );
  NAND2_X1 U9146 ( .A1(n7637), .A2(n7636), .ZN(n8130) );
  NAND2_X1 U9147 ( .A1(n7787), .A2(n7578), .ZN(n7800) );
  NAND2_X1 U9148 ( .A1(n8391), .A2(n8390), .ZN(n8395) );
  OAI21_X1 U9149 ( .B1(n8093), .B2(n7399), .A(n7397), .ZN(n7639) );
  NAND2_X1 U9150 ( .A1(n7772), .A2(n7575), .ZN(n7785) );
  OAI21_X1 U9151 ( .B1(n7045), .B2(n7040), .A(n7039), .ZN(n7038) );
  NAND2_X1 U9152 ( .A1(n7392), .A2(n7390), .ZN(n7590) );
  NAND2_X1 U9153 ( .A1(n6627), .A2(n7046), .ZN(n7043) );
  NAND2_X1 U9154 ( .A1(n7044), .A2(n7043), .ZN(n7042) );
  NAND2_X1 U9155 ( .A1(n14124), .A2(n14123), .ZN(n14122) );
  INV_X2 U9156 ( .A(n7959), .ZN(n7654) );
  OAI21_X2 U9157 ( .B1(n8209), .B2(n7531), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n6881) );
  NAND2_X1 U9158 ( .A1(n7515), .A2(n7514), .ZN(n8041) );
  NOR2_X1 U9159 ( .A1(n12766), .A2(n12783), .ZN(n12768) );
  AND2_X2 U9160 ( .A1(n12748), .A2(n12747), .ZN(n12766) );
  NAND2_X1 U9161 ( .A1(n12799), .A2(n12805), .ZN(n12832) );
  NAND2_X1 U9162 ( .A1(n12346), .A2(n12347), .ZN(n12345) );
  NOR2_X1 U9163 ( .A1(n14576), .A2(n12847), .ZN(n14603) );
  NAND4_X1 U9164 ( .A1(n14605), .A2(n14607), .A3(n14606), .A4(n14608), .ZN(
        P3_U3200) );
  NOR2_X2 U9165 ( .A1(n10863), .A2(n10864), .ZN(n12316) );
  NOR2_X1 U9166 ( .A1(n15053), .A2(n7205), .ZN(n10861) );
  NAND2_X1 U9167 ( .A1(n6718), .A2(n12008), .ZN(n12013) );
  NAND2_X1 U9168 ( .A1(n12007), .A2(n12006), .ZN(n6718) );
  INV_X1 U9169 ( .A(n12139), .ZN(n12141) );
  NAND2_X1 U9170 ( .A1(n6777), .A2(n6597), .ZN(n12149) );
  NAND2_X1 U9171 ( .A1(n12101), .A2(n6639), .ZN(n6770) );
  NAND2_X1 U9172 ( .A1(n7490), .A2(n7501), .ZN(n7489) );
  NAND2_X1 U9173 ( .A1(n6772), .A2(n6768), .ZN(n12124) );
  OAI21_X1 U9174 ( .B1(n12024), .B2(n7462), .A(n7461), .ZN(n12031) );
  NAND2_X1 U9175 ( .A1(n6764), .A2(n6762), .ZN(n12237) );
  AOI21_X1 U9176 ( .B1(n7115), .B2(n7114), .A(n7537), .ZN(n11665) );
  NAND2_X1 U9177 ( .A1(n7131), .A2(n6631), .ZN(n13269) );
  INV_X1 U9178 ( .A(n7235), .ZN(n7234) );
  NAND2_X1 U9179 ( .A1(n8616), .A2(n8615), .ZN(n8628) );
  NAND2_X1 U9180 ( .A1(n8799), .A2(n8798), .ZN(n8814) );
  OAI21_X1 U9181 ( .B1(n8883), .B2(n8882), .A(n7266), .ZN(n7265) );
  INV_X1 U9182 ( .A(n8870), .ZN(n7269) );
  OAI21_X1 U9183 ( .B1(n12903), .B2(n8978), .A(n8977), .ZN(n12890) );
  NAND2_X1 U9184 ( .A1(n12720), .A2(n12721), .ZN(n12719) );
  NAND2_X2 U9185 ( .A1(n9686), .A2(n9685), .ZN(n12661) );
  XNOR2_X2 U9186 ( .A(n12450), .B(n10251), .ZN(n11290) );
  NAND2_X1 U9187 ( .A1(n14579), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n14578) );
  NAND2_X1 U9188 ( .A1(n14578), .A2(n12855), .ZN(n14594) );
  INV_X1 U9189 ( .A(n10898), .ZN(n12348) );
  XNOR2_X2 U9190 ( .A(n9158), .B(n9157), .ZN(n13418) );
  XNOR2_X2 U9191 ( .A(n9156), .B(n9155), .ZN(n9852) );
  NAND2_X1 U9192 ( .A1(n6747), .A2(n6748), .ZN(n12139) );
  OR2_X1 U9193 ( .A1(n12136), .A2(n6749), .ZN(n6747) );
  NAND2_X1 U9194 ( .A1(n6753), .A2(n6752), .ZN(n12024) );
  OR2_X1 U9195 ( .A1(n6756), .A2(n12018), .ZN(n6752) );
  NAND2_X1 U9196 ( .A1(n6755), .A2(n6754), .ZN(n6753) );
  INV_X1 U9197 ( .A(n12017), .ZN(n6754) );
  NAND2_X1 U9198 ( .A1(n6756), .A2(n12018), .ZN(n6755) );
  NAND2_X1 U9199 ( .A1(n6758), .A2(n6757), .ZN(n6756) );
  NAND2_X1 U9200 ( .A1(n12012), .A2(n12013), .ZN(n6757) );
  OAI21_X1 U9201 ( .B1(n12012), .B2(n12013), .A(n12011), .ZN(n6758) );
  OAI21_X1 U9202 ( .B1(n12054), .B2(n6760), .A(n6759), .ZN(n12071) );
  OAI21_X1 U9203 ( .B1(n12155), .B2(n6761), .A(n6765), .ZN(n6764) );
  INV_X1 U9204 ( .A(n12158), .ZN(n6767) );
  OAI21_X1 U9205 ( .B1(n6771), .B2(n6770), .A(n6606), .ZN(n6768) );
  NAND3_X1 U9206 ( .A1(n7468), .A2(n6559), .A3(n12115), .ZN(n6772) );
  NAND2_X1 U9207 ( .A1(n12040), .A2(n12041), .ZN(n12039) );
  OAI22_X1 U9208 ( .A1(n12031), .A2(n6773), .B1(n6774), .B2(n12032), .ZN(
        n12040) );
  NAND3_X1 U9209 ( .A1(n7476), .A2(n7480), .A3(n6776), .ZN(n6775) );
  NAND3_X1 U9210 ( .A1(n7494), .A2(n7500), .A3(n7498), .ZN(n6777) );
  NAND2_X1 U9211 ( .A1(n9335), .A2(n6780), .ZN(n6778) );
  NAND2_X1 U9212 ( .A1(n6778), .A2(n6779), .ZN(n11688) );
  NAND2_X1 U9213 ( .A1(n6784), .A2(n6785), .ZN(n7163) );
  NAND2_X1 U9214 ( .A1(n13585), .A2(n6787), .ZN(n6784) );
  INV_X1 U9215 ( .A(n7156), .ZN(n6789) );
  OAI211_X2 U9216 ( .C1(n9862), .C2(n9496), .A(n6614), .B(n9174), .ZN(n13373)
         );
  NAND2_X1 U9217 ( .A1(n6799), .A2(n8380), .ZN(n6798) );
  NAND2_X1 U9218 ( .A1(n8381), .A2(n8382), .ZN(n6799) );
  NAND3_X1 U9219 ( .A1(n8281), .A2(n8279), .A3(n8280), .ZN(n6803) );
  NAND3_X1 U9220 ( .A1(n6622), .A2(n7654), .A3(n7653), .ZN(n14427) );
  NAND2_X1 U9221 ( .A1(n7654), .A2(n7653), .ZN(n8209) );
  NAND2_X1 U9222 ( .A1(n6804), .A2(n8343), .ZN(n8346) );
  NAND2_X1 U9223 ( .A1(n6805), .A2(n7550), .ZN(n6804) );
  NAND3_X1 U9224 ( .A1(n6807), .A2(n6806), .A3(n6644), .ZN(n6805) );
  NAND2_X1 U9225 ( .A1(n8329), .A2(n8321), .ZN(n6806) );
  NAND2_X1 U9226 ( .A1(n8329), .A2(n6596), .ZN(n6807) );
  OAI21_X1 U9227 ( .B1(n8356), .B2(n6816), .A(n6814), .ZN(n8359) );
  OAI21_X1 U9228 ( .B1(n8356), .B2(n6812), .A(n6808), .ZN(n8360) );
  NAND2_X1 U9229 ( .A1(n8294), .A2(n6821), .ZN(n6820) );
  INV_X1 U9230 ( .A(n7664), .ZN(n7502) );
  NAND3_X1 U9231 ( .A1(n6835), .A2(n6834), .A3(n6833), .ZN(n7652) );
  OAI21_X1 U9232 ( .B1(n12343), .B2(n6848), .A(n6845), .ZN(n15095) );
  NAND2_X1 U9233 ( .A1(n6844), .A2(n6842), .ZN(n15094) );
  NAND2_X1 U9234 ( .A1(n12343), .A2(n6845), .ZN(n6844) );
  NOR2_X1 U9235 ( .A1(n10878), .A2(n12351), .ZN(n6860) );
  NAND2_X2 U9236 ( .A1(n8511), .A2(n8512), .ZN(n8697) );
  NAND2_X1 U9237 ( .A1(n10336), .A2(n6861), .ZN(n10230) );
  AND2_X1 U9238 ( .A1(n10229), .A2(n6862), .ZN(n6861) );
  AOI21_X1 U9239 ( .B1(n12870), .B2(n15109), .A(n6869), .ZN(n12871) );
  NAND3_X1 U9240 ( .A1(n7654), .A2(n7653), .A3(n8210), .ZN(n6880) );
  XNOR2_X2 U9241 ( .A(n6882), .B(n7657), .ZN(n13962) );
  XNOR2_X1 U9242 ( .A(n11894), .B(n11895), .ZN(n13910) );
  CLKBUF_X1 U9243 ( .A(n6884), .Z(n6883) );
  INV_X1 U9244 ( .A(n6883), .ZN(n13911) );
  OR2_X1 U9245 ( .A1(n13789), .A2(n6894), .ZN(n6893) );
  NAND3_X1 U9246 ( .A1(n6893), .A2(n6892), .A3(n6889), .ZN(n13905) );
  NAND3_X1 U9247 ( .A1(n13789), .A2(n13898), .A3(n6898), .ZN(n6892) );
  NAND2_X1 U9248 ( .A1(n11952), .A2(n11951), .ZN(n6905) );
  NOR2_X1 U9249 ( .A1(n6921), .A2(n13393), .ZN(n13394) );
  NAND2_X1 U9250 ( .A1(n11088), .A2(n11085), .ZN(n6924) );
  NAND2_X1 U9251 ( .A1(n10297), .A2(n10296), .ZN(n10295) );
  NAND2_X1 U9252 ( .A1(n10181), .A2(n8171), .ZN(n10297) );
  NAND2_X1 U9253 ( .A1(n8429), .A2(n10182), .ZN(n10181) );
  NAND3_X1 U9254 ( .A1(n6927), .A2(n8314), .A3(n6926), .ZN(n11676) );
  NAND3_X1 U9255 ( .A1(n6929), .A2(n11633), .A3(n6931), .ZN(n6926) );
  NAND3_X1 U9256 ( .A1(n11459), .A2(n6929), .A3(n11633), .ZN(n6927) );
  NAND3_X1 U9257 ( .A1(n7214), .A2(n10589), .A3(n7216), .ZN(n6935) );
  NAND2_X1 U9258 ( .A1(n11751), .A2(n7228), .ZN(n6936) );
  INV_X1 U9259 ( .A(n11018), .ZN(n6941) );
  NAND2_X1 U9260 ( .A1(n6940), .A2(n6939), .ZN(n11277) );
  NAND2_X1 U9261 ( .A1(n6944), .A2(n6942), .ZN(n14208) );
  NAND2_X1 U9262 ( .A1(n8187), .A2(n8186), .ZN(n14221) );
  INV_X1 U9263 ( .A(n6948), .ZN(n6947) );
  NAND2_X1 U9264 ( .A1(n14119), .A2(n6965), .ZN(n6962) );
  NAND2_X1 U9265 ( .A1(n6962), .A2(n6963), .ZN(n8476) );
  NAND2_X1 U9266 ( .A1(n14119), .A2(n8197), .ZN(n14103) );
  INV_X1 U9267 ( .A(n6973), .ZN(n13606) );
  NAND2_X1 U9268 ( .A1(n13479), .A2(n6974), .ZN(n13442) );
  NAND2_X1 U9269 ( .A1(n11011), .A2(n15000), .ZN(n11268) );
  CLKBUF_X1 U9270 ( .A(n8586), .Z(n6980) );
  INV_X2 U9271 ( .A(n8586), .ZN(n8511) );
  NAND2_X2 U9272 ( .A1(n6981), .A2(n8520), .ZN(n9078) );
  NAND2_X1 U9273 ( .A1(n12937), .A2(n6985), .ZN(n6984) );
  OAI21_X1 U9274 ( .B1(n9045), .B2(n6994), .A(n6991), .ZN(n11169) );
  NAND2_X1 U9275 ( .A1(n6990), .A2(n6988), .ZN(n9046) );
  NAND2_X1 U9276 ( .A1(n9045), .A2(n6991), .ZN(n6990) );
  OAI21_X1 U9277 ( .B1(n11446), .B2(n7002), .A(n6998), .ZN(n11620) );
  NAND2_X1 U9278 ( .A1(n6997), .A2(n6995), .ZN(n9049) );
  NAND2_X1 U9279 ( .A1(n11446), .A2(n6998), .ZN(n6997) );
  OAI21_X1 U9280 ( .B1(n11446), .B2(n12477), .A(n12413), .ZN(n11525) );
  NAND2_X1 U9281 ( .A1(n7005), .A2(n7004), .ZN(n9048) );
  NAND2_X1 U9282 ( .A1(n13045), .A2(n7006), .ZN(n13032) );
  AOI21_X2 U9283 ( .B1(n7007), .B2(n7263), .A(n6626), .ZN(n12380) );
  NAND2_X1 U9284 ( .A1(n7008), .A2(n12518), .ZN(n13003) );
  NAND2_X1 U9285 ( .A1(n7008), .A2(n6638), .ZN(n13001) );
  NAND2_X2 U9286 ( .A1(n9030), .A2(n13205), .ZN(n8565) );
  XNOR2_X2 U9287 ( .A(n7009), .B(n8536), .ZN(n13205) );
  NOR2_X2 U9288 ( .A1(n11898), .A2(n11755), .ZN(n14264) );
  NOR2_X2 U9289 ( .A1(n11281), .A2(n11555), .ZN(n11282) );
  NAND3_X1 U9290 ( .A1(n7016), .A2(n10307), .A3(n10642), .ZN(n10548) );
  INV_X1 U9291 ( .A(n10744), .ZN(n7016) );
  INV_X1 U9292 ( .A(n7017), .ZN(n10601) );
  NOR2_X2 U9293 ( .A1(n14109), .A2(n14396), .ZN(n7021) );
  INV_X1 U9294 ( .A(n7027), .ZN(n14163) );
  NOR2_X2 U9295 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n7684) );
  INV_X1 U9296 ( .A(n7033), .ZN(n7029) );
  INV_X1 U9297 ( .A(n7031), .ZN(n7030) );
  INV_X1 U9298 ( .A(n8368), .ZN(n7032) );
  NAND2_X1 U9299 ( .A1(n8411), .A2(n7034), .ZN(n7035) );
  INV_X1 U9300 ( .A(n8427), .ZN(n7045) );
  INV_X1 U9301 ( .A(n8410), .ZN(n7046) );
  INV_X1 U9302 ( .A(n8282), .ZN(n7048) );
  XNOR2_X1 U9303 ( .A(n7733), .B(n10379), .ZN(n10300) );
  AND2_X1 U9304 ( .A1(n7724), .A2(n7725), .ZN(n7049) );
  INV_X1 U9305 ( .A(n8377), .ZN(n7055) );
  NAND2_X1 U9306 ( .A1(n7058), .A2(n7056), .ZN(n8300) );
  NAND2_X1 U9307 ( .A1(n8296), .A2(n7059), .ZN(n7058) );
  INV_X1 U9308 ( .A(n8361), .ZN(n7064) );
  NAND2_X1 U9309 ( .A1(n8272), .A2(n8273), .ZN(n8271) );
  NAND3_X1 U9310 ( .A1(n7654), .A2(n7530), .A3(n7653), .ZN(n7066) );
  NAND2_X1 U9311 ( .A1(n9537), .A2(n12247), .ZN(n7072) );
  XNOR2_X1 U9312 ( .A(n13374), .B(n14934), .ZN(n12247) );
  INV_X1 U9313 ( .A(n9183), .ZN(n7073) );
  NAND3_X1 U9314 ( .A1(n7072), .A2(n10078), .A3(n7071), .ZN(n10072) );
  XNOR2_X2 U9315 ( .A(n7075), .B(n7074), .ZN(n9149) );
  NAND3_X1 U9316 ( .A1(n6643), .A2(n9144), .A3(n7541), .ZN(n7076) );
  NAND2_X1 U9317 ( .A1(n13583), .A2(n7080), .ZN(n7077) );
  NAND2_X1 U9318 ( .A1(n7091), .A2(n7089), .ZN(n10715) );
  NAND2_X1 U9319 ( .A1(n13623), .A2(n9563), .ZN(n13596) );
  NAND2_X1 U9320 ( .A1(n11570), .A2(n7109), .ZN(n7104) );
  NAND2_X1 U9321 ( .A1(n7113), .A2(n7112), .ZN(n10097) );
  OR2_X1 U9322 ( .A1(n10095), .A2(n10096), .ZN(n7112) );
  NAND2_X1 U9323 ( .A1(n11830), .A2(n11829), .ZN(n11836) );
  NAND2_X1 U9324 ( .A1(n11665), .A2(n11666), .ZN(n11830) );
  INV_X1 U9325 ( .A(n11660), .ZN(n7115) );
  NAND2_X1 U9326 ( .A1(n13336), .A2(n7117), .ZN(n7116) );
  OAI211_X1 U9327 ( .C1(n13336), .C2(n7118), .A(n7116), .B(n13288), .ZN(
        P2_U3192) );
  NAND2_X1 U9328 ( .A1(n13336), .A2(n13255), .ZN(n13280) );
  INV_X1 U9329 ( .A(n11863), .ZN(n7132) );
  NAND2_X1 U9330 ( .A1(n10784), .A2(n10935), .ZN(n7140) );
  NAND3_X1 U9331 ( .A1(n9578), .A2(n12289), .A3(n12613), .ZN(n7144) );
  AND2_X1 U9332 ( .A1(n9376), .A2(n7146), .ZN(n9516) );
  NAND2_X1 U9333 ( .A1(n9376), .A2(n7147), .ZN(n9518) );
  INV_X1 U9334 ( .A(n9515), .ZN(n7151) );
  NAND2_X1 U9335 ( .A1(n13560), .A2(n9568), .ZN(n13529) );
  NAND2_X1 U9336 ( .A1(n13514), .A2(n9570), .ZN(n13491) );
  NAND2_X1 U9337 ( .A1(n10143), .A2(n12249), .ZN(n10142) );
  AND2_X2 U9338 ( .A1(n10010), .A2(n10009), .ZN(n10131) );
  NAND2_X2 U9339 ( .A1(n10533), .A2(n9579), .ZN(n10429) );
  AND4_X2 U9340 ( .A1(n9143), .A2(n9515), .A3(n9142), .A4(n9141), .ZN(n7541)
         );
  AND3_X4 U9341 ( .A1(n7231), .A2(n7688), .A3(n7230), .ZN(n14792) );
  AND2_X2 U9342 ( .A1(n10305), .A2(n7734), .ZN(n10307) );
  NOR2_X2 U9343 ( .A1(n14226), .A2(n14415), .ZN(n14211) );
  NAND2_X1 U9344 ( .A1(n7152), .A2(n10144), .ZN(n9198) );
  XNOR2_X1 U9345 ( .A(n7152), .B(n10144), .ZN(n10145) );
  NAND2_X1 U9346 ( .A1(n10241), .A2(n12251), .ZN(n7153) );
  NAND4_X1 U9347 ( .A1(n9311), .A2(n9201), .A3(n9140), .A4(n7155), .ZN(n7154)
         );
  INV_X1 U9348 ( .A(n9144), .ZN(n9351) );
  OAI21_X1 U9349 ( .B1(n13585), .B2(n7160), .A(n7159), .ZN(n13546) );
  NAND2_X1 U9350 ( .A1(n7163), .A2(n7165), .ZN(n9483) );
  NAND2_X1 U9351 ( .A1(n7176), .A2(n7175), .ZN(n9402) );
  NAND2_X1 U9352 ( .A1(n9491), .A2(n12244), .ZN(n13460) );
  NAND2_X1 U9353 ( .A1(n7192), .A2(n7190), .ZN(n9268) );
  INV_X1 U9354 ( .A(n7196), .ZN(n15036) );
  NAND2_X1 U9355 ( .A1(n7197), .A2(n15045), .ZN(n7195) );
  XNOR2_X1 U9356 ( .A(n7197), .B(n15045), .ZN(n15037) );
  NAND2_X1 U9357 ( .A1(n10858), .A2(n7198), .ZN(n7197) );
  INV_X1 U9358 ( .A(n10892), .ZN(n7199) );
  OR2_X1 U9359 ( .A1(n10327), .A2(n10219), .ZN(n10329) );
  XNOR2_X2 U9360 ( .A(n8539), .B(P3_IR_REG_1__SCAN_IN), .ZN(n10345) );
  NAND2_X1 U9361 ( .A1(n7203), .A2(n12800), .ZN(n7202) );
  NAND3_X1 U9362 ( .A1(n7202), .A2(n7201), .A3(n6678), .ZN(n12845) );
  INV_X1 U9363 ( .A(n7209), .ZN(n15092) );
  NAND2_X1 U9364 ( .A1(n12768), .A2(n12787), .ZN(n7210) );
  INV_X1 U9365 ( .A(n14120), .ZN(n7213) );
  NAND3_X1 U9366 ( .A1(n10286), .A2(n10287), .A3(n10496), .ZN(n7216) );
  INV_X1 U9367 ( .A(n10286), .ZN(n7219) );
  OAI21_X1 U9368 ( .B1(n10287), .B2(n7221), .A(n10496), .ZN(n7220) );
  NAND2_X1 U9369 ( .A1(n7219), .A2(n8173), .ZN(n7217) );
  INV_X1 U9370 ( .A(n7220), .ZN(n7218) );
  NAND2_X1 U9371 ( .A1(n10592), .A2(n7227), .ZN(n10805) );
  NAND2_X1 U9372 ( .A1(n13883), .A2(n14792), .ZN(n8247) );
  NAND2_X1 U9373 ( .A1(n8559), .A2(n8560), .ZN(n7233) );
  NAND2_X1 U9374 ( .A1(n8589), .A2(n7237), .ZN(n7236) );
  NAND2_X1 U9375 ( .A1(n7236), .A2(n7234), .ZN(n8616) );
  INV_X1 U9376 ( .A(n7238), .ZN(n7237) );
  INV_X1 U9377 ( .A(n8589), .ZN(n7240) );
  INV_X1 U9378 ( .A(n8591), .ZN(n7241) );
  NAND2_X1 U9379 ( .A1(n8997), .A2(n7243), .ZN(n7242) );
  NAND2_X1 U9380 ( .A1(n7250), .A2(n8999), .ZN(n9015) );
  NAND2_X1 U9381 ( .A1(n8681), .A2(n6628), .ZN(n7255) );
  AOI21_X2 U9382 ( .B1(n7269), .B2(n7268), .A(n7267), .ZN(n8883) );
  XNOR2_X2 U9383 ( .A(n8943), .B(P2_DATAO_REG_24__SCAN_IN), .ZN(n8944) );
  OR2_X2 U9384 ( .A1(n8918), .A2(n7272), .ZN(n7271) );
  XNOR2_X2 U9385 ( .A(n14449), .B(n14450), .ZN(n14501) );
  AND2_X2 U9386 ( .A1(n7277), .A2(n6630), .ZN(n14449) );
  NAND2_X1 U9387 ( .A1(n14559), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n7290) );
  NAND2_X1 U9388 ( .A1(n14559), .A2(n7286), .ZN(n7285) );
  NAND2_X1 U9389 ( .A1(n14703), .A2(n7298), .ZN(n7296) );
  AOI21_X1 U9390 ( .B1(n14703), .B2(n7293), .A(n7291), .ZN(n7300) );
  INV_X1 U9391 ( .A(n14708), .ZN(n7292) );
  AND2_X1 U9392 ( .A1(n7298), .A2(n14708), .ZN(n7293) );
  NAND2_X1 U9393 ( .A1(n7296), .A2(n7297), .ZN(n14707) );
  NAND2_X1 U9394 ( .A1(n12661), .A2(n7304), .ZN(n7301) );
  NAND2_X1 U9395 ( .A1(n7301), .A2(n7302), .ZN(n12632) );
  OAI21_X1 U9396 ( .B1(n10651), .B2(n7310), .A(n7307), .ZN(n9664) );
  NAND2_X1 U9397 ( .A1(n11044), .A2(n7322), .ZN(n7326) );
  NAND2_X1 U9398 ( .A1(n12419), .A2(n9626), .ZN(n12407) );
  NAND3_X1 U9399 ( .A1(n7329), .A2(n12419), .A3(n9626), .ZN(n7328) );
  INV_X1 U9400 ( .A(n9625), .ZN(n7329) );
  XNOR2_X2 U9401 ( .A(n9027), .B(n9026), .ZN(n12419) );
  INV_X1 U9402 ( .A(n9740), .ZN(n12578) );
  NAND3_X1 U9403 ( .A1(n8511), .A2(n8512), .A3(n7445), .ZN(n7331) );
  NAND2_X1 U9404 ( .A1(n11437), .A2(n7337), .ZN(n7336) );
  NAND2_X1 U9405 ( .A1(n13804), .A2(n7340), .ZN(n13878) );
  NAND2_X1 U9406 ( .A1(n10355), .A2(n10356), .ZN(n7340) );
  NAND2_X1 U9407 ( .A1(n13840), .A2(n7345), .ZN(n7344) );
  INV_X1 U9408 ( .A(n11909), .ZN(n7350) );
  NAND2_X1 U9409 ( .A1(n13840), .A2(n13841), .ZN(n13839) );
  NAND2_X1 U9410 ( .A1(n11915), .A2(n11914), .ZN(n7351) );
  OAI21_X1 U9411 ( .B1(n13848), .B2(n7360), .A(n7357), .ZN(n13782) );
  OAI21_X1 U9412 ( .B1(n13848), .B2(n13849), .A(n11959), .ZN(n13823) );
  NAND2_X1 U9413 ( .A1(n11965), .A2(n11964), .ZN(n7368) );
  AND4_X1 U9414 ( .A1(n7649), .A2(n6569), .A3(n7743), .A4(n7648), .ZN(n7971)
         );
  AND2_X2 U9415 ( .A1(n7648), .A2(n7970), .ZN(n7371) );
  NOR2_X2 U9416 ( .A1(n7993), .A2(P1_IR_REG_18__SCAN_IN), .ZN(n7997) );
  NAND3_X1 U9417 ( .A1(n13876), .A2(n10370), .A3(n10371), .ZN(n10625) );
  NAND3_X1 U9418 ( .A1(n8153), .A2(n6549), .A3(n14061), .ZN(n10823) );
  NAND3_X1 U9419 ( .A1(n13415), .A2(P3_ADDR_REG_19__SCAN_IN), .A3(n7374), .ZN(
        n7555) );
  NAND2_X1 U9420 ( .A1(n8052), .A2(n7624), .ZN(n7375) );
  NAND2_X1 U9421 ( .A1(n7569), .A2(n7380), .ZN(n7378) );
  NAND2_X1 U9422 ( .A1(n7378), .A2(n7379), .ZN(n7772) );
  INV_X1 U9423 ( .A(n7557), .ZN(n7383) );
  NAND2_X1 U9424 ( .A1(n7384), .A2(n7558), .ZN(n7706) );
  NAND2_X1 U9425 ( .A1(n7658), .A2(n15479), .ZN(n7386) );
  NAND2_X1 U9426 ( .A1(n7816), .A2(n7393), .ZN(n7392) );
  OAI21_X1 U9427 ( .B1(n7816), .B2(n7394), .A(n7393), .ZN(n7847) );
  AOI21_X1 U9428 ( .B1(n7393), .B2(n7394), .A(n7391), .ZN(n7390) );
  INV_X1 U9429 ( .A(n7639), .ZN(n7637) );
  NAND2_X1 U9430 ( .A1(n12160), .A2(n12168), .ZN(n7406) );
  NAND2_X1 U9431 ( .A1(n7881), .A2(n7412), .ZN(n7408) );
  NAND2_X1 U9432 ( .A1(n7881), .A2(n7880), .ZN(n7411) );
  NAND2_X1 U9433 ( .A1(n11342), .A2(n7421), .ZN(n7420) );
  NAND2_X1 U9434 ( .A1(n7420), .A2(n7423), .ZN(n11622) );
  NAND2_X1 U9435 ( .A1(n8568), .A2(n15115), .ZN(n15122) );
  AOI21_X1 U9436 ( .B1(n8897), .B2(n6635), .A(n7434), .ZN(n12903) );
  NAND2_X1 U9437 ( .A1(n11070), .A2(n7443), .ZN(n7442) );
  NAND2_X1 U9438 ( .A1(n7445), .A2(n8519), .ZN(n7444) );
  OR2_X2 U9439 ( .A1(n9078), .A2(n7448), .ZN(n8535) );
  NOR2_X2 U9440 ( .A1(n9078), .A2(n7446), .ZN(n8526) );
  NAND2_X1 U9441 ( .A1(n13020), .A2(n7450), .ZN(n13011) );
  NAND2_X1 U9442 ( .A1(n12097), .A2(n12098), .ZN(n12096) );
  NAND2_X1 U9443 ( .A1(n7456), .A2(n7455), .ZN(n7454) );
  INV_X1 U9444 ( .A(n12089), .ZN(n7455) );
  INV_X1 U9445 ( .A(n7460), .ZN(n7456) );
  NAND2_X1 U9446 ( .A1(n7459), .A2(n7458), .ZN(n7457) );
  NAND2_X1 U9447 ( .A1(n7460), .A2(n12089), .ZN(n7459) );
  INV_X1 U9448 ( .A(n12022), .ZN(n7463) );
  INV_X1 U9449 ( .A(n12023), .ZN(n7464) );
  NAND3_X1 U9450 ( .A1(n12045), .A2(n6647), .A3(n12044), .ZN(n7465) );
  NAND2_X1 U9451 ( .A1(n7465), .A2(n7466), .ZN(n12056) );
  AOI21_X1 U9452 ( .B1(n12056), .B2(n12055), .A(n12053), .ZN(n12054) );
  NAND3_X1 U9453 ( .A1(n12102), .A2(n12101), .A3(n6586), .ZN(n7468) );
  INV_X1 U9454 ( .A(n12107), .ZN(n7471) );
  NAND3_X1 U9455 ( .A1(n12072), .A2(n12071), .A3(n6629), .ZN(n7476) );
  NAND3_X1 U9456 ( .A1(n12072), .A2(n12071), .A3(n6636), .ZN(n7479) );
  NAND3_X1 U9457 ( .A1(n12057), .A2(n6556), .A3(n6637), .ZN(n7485) );
  NAND2_X1 U9458 ( .A1(n12141), .A2(n12142), .ZN(n7490) );
  NAND2_X1 U9459 ( .A1(n12140), .A2(n7495), .ZN(n7493) );
  OR2_X1 U9460 ( .A1(n7489), .A2(n12140), .ZN(n7494) );
  INV_X1 U9461 ( .A(n7703), .ZN(n7760) );
  AOI21_X1 U9462 ( .B1(n7760), .B2(P1_REG3_REG_1__SCAN_IN), .A(n7505), .ZN(
        n7504) );
  NAND3_X1 U9463 ( .A1(n7649), .A2(n7743), .A3(n7648), .ZN(n7921) );
  NAND2_X1 U9464 ( .A1(n11183), .A2(n7509), .ZN(n7508) );
  NAND2_X1 U9465 ( .A1(n14766), .A2(n10178), .ZN(n7719) );
  NAND2_X2 U9466 ( .A1(n11354), .A2(n11353), .ZN(n11352) );
  OR2_X2 U9467 ( .A1(n8010), .A2(n6625), .ZN(n7515) );
  NAND2_X1 U9468 ( .A1(n8107), .A2(n8106), .ZN(n8478) );
  NAND2_X1 U9469 ( .A1(n7938), .A2(n6642), .ZN(n7523) );
  OAI21_X1 U9470 ( .B1(n12888), .B2(n12889), .A(n12887), .ZN(n13085) );
  NAND2_X1 U9471 ( .A1(n12888), .A2(n12889), .ZN(n12887) );
  NOR2_X1 U9472 ( .A1(n14759), .A2(n13884), .ZN(n10305) );
  INV_X1 U9473 ( .A(n8834), .ZN(n8836) );
  NAND2_X1 U9474 ( .A1(n12719), .A2(n9715), .ZN(n12617) );
  INV_X1 U9475 ( .A(n15138), .ZN(n9042) );
  NAND2_X1 U9476 ( .A1(n13431), .A2(n13430), .ZN(n13432) );
  OAI21_X1 U9477 ( .B1(n13459), .B2(n13730), .A(n13453), .ZN(n9581) );
  CLKBUF_X1 U9478 ( .A(n9080), .Z(n9081) );
  NAND2_X1 U9479 ( .A1(n8482), .A2(n8448), .ZN(n8483) );
  INV_X1 U9480 ( .A(n15137), .ZN(n8567) );
  OR2_X1 U9481 ( .A1(n10796), .A2(n11531), .ZN(n8716) );
  OR2_X1 U9482 ( .A1(n10796), .A2(n10859), .ZN(n8553) );
  BUF_X2 U9483 ( .A(n8565), .Z(n10198) );
  INV_X1 U9484 ( .A(n6828), .ZN(n14435) );
  NAND2_X1 U9485 ( .A1(n7502), .A2(n14435), .ZN(n7699) );
  OAI22_X1 U9486 ( .A1(n12409), .A2(n12408), .B1(n12407), .B2(n12406), .ZN(
        n12580) );
  INV_X1 U9487 ( .A(n8530), .ZN(n12591) );
  INV_X1 U9488 ( .A(n13764), .ZN(n9616) );
  INV_X1 U9489 ( .A(n14142), .ZN(n8075) );
  OR2_X1 U9490 ( .A1(n13711), .A2(n12134), .ZN(n7533) );
  AND2_X1 U9491 ( .A1(n8327), .A2(n8326), .ZN(n7534) );
  OR2_X1 U9492 ( .A1(n8027), .A2(SI_21_), .ZN(n7535) );
  AND2_X1 U9493 ( .A1(n9408), .A2(n9520), .ZN(n7536) );
  INV_X1 U9494 ( .A(n13372), .ZN(n9196) );
  AND2_X1 U9495 ( .A1(n11664), .A2(n11663), .ZN(n7537) );
  OR2_X1 U9496 ( .A1(n9620), .A2(n14411), .ZN(n7539) );
  AND2_X1 U9497 ( .A1(n9303), .A2(n9302), .ZN(n7540) );
  AND2_X1 U9498 ( .A1(n7701), .A2(n7700), .ZN(n7542) );
  OR2_X1 U9499 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(n15020), .ZN(n7543) );
  OR2_X1 U9500 ( .A1(n14763), .A2(n14760), .ZN(n7544) );
  XNOR2_X1 U9501 ( .A(n12876), .B(n12375), .ZN(n12381) );
  AND2_X1 U9502 ( .A1(n8317), .A2(n8316), .ZN(n7545) );
  AND2_X1 U9503 ( .A1(n7598), .A2(n7599), .ZN(n7546) );
  AND2_X1 U9504 ( .A1(n9748), .A2(n9747), .ZN(n7548) );
  AND3_X1 U9505 ( .A1(n9721), .A2(n12722), .A3(n9720), .ZN(n7549) );
  AND3_X1 U9506 ( .A1(n14223), .A2(n8339), .A3(n8338), .ZN(n7550) );
  OR2_X1 U9507 ( .A1(n8022), .A2(SI_20_), .ZN(n7551) );
  INV_X1 U9508 ( .A(n11633), .ZN(n7911) );
  INV_X1 U9509 ( .A(n12263), .ZN(n9323) );
  AND2_X1 U9510 ( .A1(n12188), .A2(n12187), .ZN(n7552) );
  AOI22_X1 U9511 ( .A1(n12293), .A2(n13374), .B1(n12153), .B2(n14934), .ZN(
        n12012) );
  NAND2_X1 U9512 ( .A1(n8275), .A2(n8274), .ZN(n8280) );
  OAI21_X1 U9513 ( .B1(n12037), .B2(n12293), .A(n12036), .ZN(n12038) );
  OAI21_X1 U9514 ( .B1(n12112), .B2(n12293), .A(n12111), .ZN(n12113) );
  NOR2_X1 U9515 ( .A1(n12899), .A2(n12400), .ZN(n12401) );
  NAND2_X1 U9516 ( .A1(n12889), .A2(n12401), .ZN(n12402) );
  INV_X1 U9517 ( .A(n12193), .ZN(n12190) );
  NOR2_X1 U9518 ( .A1(n12560), .A2(n12402), .ZN(n12403) );
  INV_X1 U9519 ( .A(n15117), .ZN(n8566) );
  INV_X1 U9520 ( .A(n7956), .ZN(n7608) );
  NAND2_X1 U9521 ( .A1(n9065), .A2(n12403), .ZN(n12404) );
  INV_X1 U9522 ( .A(n13004), .ZN(n9053) );
  OR2_X1 U9523 ( .A1(n8714), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8730) );
  OR2_X1 U9524 ( .A1(n14637), .A2(n11518), .ZN(n8720) );
  INV_X1 U9525 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n8965) );
  INV_X1 U9526 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n8900) );
  INV_X1 U9527 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n9243) );
  NOR2_X1 U9528 ( .A1(n7929), .A2(n7928), .ZN(n7927) );
  NOR2_X1 U9529 ( .A1(n8016), .A2(n13859), .ZN(n8015) );
  NAND2_X1 U9530 ( .A1(n7620), .A2(SI_22_), .ZN(n7621) );
  INV_X1 U9531 ( .A(n7831), .ZN(n7585) );
  NOR2_X1 U9532 ( .A1(n14482), .A2(n14481), .ZN(n14463) );
  NOR2_X1 U9533 ( .A1(n8934), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n8951) );
  OR2_X1 U9534 ( .A1(n8921), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8934) );
  NAND2_X1 U9535 ( .A1(n8671), .A2(n15461), .ZN(n8688) );
  NOR2_X1 U9536 ( .A1(n8640), .A2(n12331), .ZN(n10863) );
  NAND2_X1 U9537 ( .A1(n13084), .A2(n9745), .ZN(n12879) );
  INV_X1 U9538 ( .A(n9028), .ZN(n9022) );
  INV_X1 U9539 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n8709) );
  INV_X1 U9540 ( .A(n12239), .ZN(n12240) );
  OR2_X1 U9541 ( .A1(n9415), .A2(n9414), .ZN(n9425) );
  OR2_X1 U9542 ( .A1(n9994), .A2(n9995), .ZN(n10112) );
  AND2_X1 U9543 ( .A1(n9366), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n9380) );
  NAND2_X1 U9544 ( .A1(n9317), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n9345) );
  OR2_X1 U9545 ( .A1(n9275), .A2(n9274), .ZN(n9287) );
  OR2_X1 U9546 ( .A1(n9283), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n9284) );
  INV_X1 U9547 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n7554) );
  INV_X1 U9548 ( .A(n11943), .ZN(n11944) );
  INV_X1 U9549 ( .A(n11548), .ZN(n11545) );
  NAND2_X1 U9550 ( .A1(n11900), .A2(n11901), .ZN(n11902) );
  INV_X1 U9551 ( .A(n11921), .ZN(n11922) );
  INV_X1 U9552 ( .A(n8067), .ZN(n8082) );
  OR2_X1 U9553 ( .A1(n8004), .A2(n7666), .ZN(n8016) );
  NOR2_X1 U9554 ( .A1(n7807), .A2(n7665), .ZN(n7823) );
  NAND2_X1 U9555 ( .A1(n8152), .A2(n12608), .ZN(n8155) );
  AND2_X1 U9556 ( .A1(n14439), .A2(n8157), .ZN(n10048) );
  XNOR2_X1 U9557 ( .A(n8416), .B(n8415), .ZN(n12160) );
  INV_X1 U9558 ( .A(n8205), .ZN(n8203) );
  INV_X4 U9559 ( .A(n7388), .ZN(n7602) );
  NOR2_X1 U9560 ( .A1(n7585), .A2(n9785), .ZN(n7586) );
  OR2_X1 U9561 ( .A1(n14480), .A2(n14479), .ZN(n14567) );
  NAND2_X1 U9562 ( .A1(n8887), .A2(n12641), .ZN(n8906) );
  INV_X1 U9563 ( .A(n12957), .ZN(n12925) );
  NOR2_X1 U9564 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_REG3_REG_3__SCAN_IN), 
        .ZN(n8599) );
  OR2_X1 U9565 ( .A1(n8906), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8921) );
  INV_X1 U9566 ( .A(n8866), .ZN(n10793) );
  NOR2_X1 U9567 ( .A1(n8985), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n9003) );
  INV_X1 U9568 ( .A(n12733), .ZN(n13037) );
  AND2_X1 U9569 ( .A1(n12474), .A2(n12478), .ZN(n11621) );
  NOR2_X1 U9570 ( .A1(n8638), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8658) );
  INV_X1 U9571 ( .A(n13138), .ZN(n9128) );
  NAND2_X1 U9572 ( .A1(n13204), .A2(n12362), .ZN(n9001) );
  AND2_X1 U9573 ( .A1(n9070), .A2(n10384), .ZN(n15147) );
  OR2_X1 U9574 ( .A1(n9067), .A2(n9066), .ZN(n9730) );
  NAND2_X1 U9575 ( .A1(n9772), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n8627) );
  AND3_X1 U9576 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .A3(P2_REG3_REG_5__SCAN_IN), .ZN(n9230) );
  NOR2_X1 U9577 ( .A1(n9355), .A2(n11701), .ZN(n9366) );
  OAI21_X1 U9578 ( .B1(n12303), .B2(n12299), .A(n12298), .ZN(n12300) );
  NOR2_X1 U9579 ( .A1(n9425), .A2(n13317), .ZN(n9434) );
  OR2_X1 U9580 ( .A1(n14861), .A2(n14860), .ZN(n14863) );
  XNOR2_X1 U9581 ( .A(n13661), .B(n13352), .ZN(n13471) );
  INV_X1 U9582 ( .A(n13479), .ZN(n13499) );
  INV_X1 U9583 ( .A(n10144), .ZN(n12249) );
  INV_X1 U9584 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n13732) );
  INV_X1 U9585 ( .A(n13363), .ZN(n11428) );
  AND2_X1 U9586 ( .A1(n9523), .A2(n12288), .ZN(n13600) );
  NAND2_X1 U9587 ( .A1(n9520), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9522) );
  NAND2_X1 U9588 ( .A1(n11945), .A2(n11944), .ZN(n11946) );
  AND2_X1 U9589 ( .A1(n7722), .A2(n7721), .ZN(n7726) );
  OR2_X1 U9590 ( .A1(n14373), .A2(n14666), .ZN(n8319) );
  INV_X1 U9591 ( .A(n14757), .ZN(n14276) );
  AND2_X1 U9592 ( .A1(n8223), .A2(n8222), .ZN(n9774) );
  NAND2_X1 U9593 ( .A1(n7627), .A2(n7626), .ZN(n8079) );
  XNOR2_X1 U9594 ( .A(n7595), .B(SI_13_), .ZN(n7880) );
  NOR2_X1 U9595 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n14501), .ZN(n14451) );
  INV_X1 U9596 ( .A(n15135), .ZN(n10252) );
  AND2_X1 U9597 ( .A1(n9742), .A2(n9741), .ZN(n12728) );
  AND2_X1 U9598 ( .A1(n8994), .A2(n8993), .ZN(n9745) );
  NOR2_X1 U9599 ( .A1(n12891), .A2(n13064), .ZN(n12892) );
  AND2_X1 U9600 ( .A1(n12471), .A2(n8686), .ZN(n12465) );
  INV_X1 U9601 ( .A(n14613), .ZN(n14617) );
  AND2_X1 U9602 ( .A1(n15132), .A2(n15131), .ZN(n15151) );
  INV_X1 U9603 ( .A(n15222), .ZN(n9126) );
  AND2_X1 U9604 ( .A1(n9118), .A2(n9117), .ZN(n10386) );
  NAND2_X1 U9605 ( .A1(n12416), .A2(n12419), .ZN(n15200) );
  AND4_X1 U9606 ( .A1(n9461), .A2(n9460), .A3(n9459), .A4(n9458), .ZN(n13549)
         );
  OR2_X1 U9607 ( .A1(n10114), .A2(n10113), .ZN(n10271) );
  AND2_X1 U9608 ( .A1(n9866), .A2(n9845), .ZN(n14914) );
  INV_X1 U9609 ( .A(n12279), .ZN(n9576) );
  INV_X1 U9610 ( .A(n13610), .ZN(n14935) );
  INV_X1 U9611 ( .A(n14939), .ZN(n13613) );
  INV_X1 U9612 ( .A(n13600), .ZN(n13618) );
  NAND2_X1 U9613 ( .A1(n15005), .A2(n13732), .ZN(n13733) );
  AND2_X1 U9614 ( .A1(n9258), .A2(n9283), .ZN(n9991) );
  OR2_X1 U9615 ( .A1(n7905), .A2(n7904), .ZN(n7929) );
  INV_X1 U9616 ( .A(n10360), .ZN(n10044) );
  AND2_X1 U9617 ( .A1(n13818), .A2(n14757), .ZN(n13900) );
  INV_X1 U9618 ( .A(n14746), .ZN(n14059) );
  INV_X1 U9619 ( .A(n14271), .ZN(n14258) );
  INV_X1 U9620 ( .A(n14755), .ZN(n14803) );
  OR3_X1 U9621 ( .A1(n10051), .A2(n8233), .A3(n8239), .ZN(n10509) );
  AND2_X1 U9622 ( .A1(n7887), .A2(n7900), .ZN(n10672) );
  NAND2_X1 U9623 ( .A1(n7706), .A2(n7560), .ZN(n7709) );
  AND2_X1 U9624 ( .A1(n10215), .A2(n10214), .ZN(n15106) );
  INV_X1 U9625 ( .A(n12702), .ZN(n12731) );
  INV_X1 U9626 ( .A(n9745), .ZN(n12906) );
  NAND4_X2 U9627 ( .A1(n8573), .A2(n8572), .A3(n8571), .A4(n8570), .ZN(n15120)
         );
  INV_X1 U9628 ( .A(n15023), .ZN(n15113) );
  INV_X1 U9629 ( .A(n15151), .ZN(n12916) );
  AND2_X1 U9630 ( .A1(n9132), .A2(n9131), .ZN(n9133) );
  AND2_X1 U9631 ( .A1(n9096), .A2(n9095), .ZN(n13192) );
  INV_X1 U9632 ( .A(SI_10_), .ZN(n9785) );
  INV_X1 U9633 ( .A(n10903), .ZN(n12324) );
  INV_X1 U9634 ( .A(n10896), .ZN(n15083) );
  INV_X1 U9635 ( .A(n13703), .ZN(n13591) );
  INV_X1 U9636 ( .A(n13549), .ZN(n13354) );
  OR2_X1 U9637 ( .A1(n9866), .A2(P2_U3088), .ZN(n14932) );
  OR2_X1 U9638 ( .A1(n14947), .A2(n10610), .ZN(n14942) );
  INV_X1 U9639 ( .A(n15019), .ZN(n15017) );
  INV_X1 U9640 ( .A(n15007), .ZN(n15005) );
  INV_X1 U9641 ( .A(n14949), .ZN(n14950) );
  INV_X1 U9642 ( .A(n14953), .ZN(n14956) );
  INV_X1 U9643 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n10069) );
  AND2_X1 U9644 ( .A1(n9930), .A2(n9916), .ZN(n14719) );
  OR2_X1 U9645 ( .A1(n10054), .A2(n10050), .ZN(n14674) );
  OR3_X1 U9646 ( .A1(n7969), .A2(n7968), .A3(n7967), .ZN(n13925) );
  OR3_X1 U9647 ( .A1(n8240), .A2(n10051), .A3(n10045), .ZN(n14809) );
  OR2_X1 U9648 ( .A1(n14806), .A2(n8235), .ZN(n8236) );
  OR2_X1 U9649 ( .A1(n10509), .A2(n8240), .ZN(n14804) );
  INV_X1 U9650 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n15454) );
  INV_X1 U9651 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n9757) );
  NAND2_X1 U9652 ( .A1(n9114), .A2(n9113), .ZN(P3_U3456) );
  NAND2_X1 U9653 ( .A1(n8507), .A2(n8506), .ZN(P1_U3524) );
  NAND2_X1 U9654 ( .A1(n7557), .A2(SI_1_), .ZN(n7558) );
  INV_X1 U9655 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n15478) );
  INV_X1 U9656 ( .A(SI_0_), .ZN(n7695) );
  MUX2_X1 U9657 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(P1_DATAO_REG_2__SCAN_IN), 
        .S(n7658), .Z(n7559) );
  NAND2_X1 U9658 ( .A1(n7559), .A2(SI_2_), .ZN(n7561) );
  INV_X1 U9659 ( .A(n7707), .ZN(n7560) );
  NAND2_X1 U9660 ( .A1(n7709), .A2(n7561), .ZN(n7730) );
  INV_X1 U9661 ( .A(n7729), .ZN(n7563) );
  NAND2_X1 U9662 ( .A1(n7730), .A2(n7563), .ZN(n7565) );
  NAND2_X1 U9663 ( .A1(n7565), .A2(n7564), .ZN(n7741) );
  MUX2_X1 U9664 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(P1_DATAO_REG_4__SCAN_IN), 
        .S(n7602), .Z(n7566) );
  INV_X1 U9665 ( .A(n7740), .ZN(n7567) );
  MUX2_X1 U9666 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n7658), .Z(n7570) );
  OAI21_X1 U9667 ( .B1(n7570), .B2(SI_5_), .A(n7572), .ZN(n7571) );
  MUX2_X1 U9668 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n7602), .Z(n7573) );
  OAI21_X1 U9669 ( .B1(SI_6_), .B2(n7573), .A(n7575), .ZN(n7574) );
  INV_X1 U9670 ( .A(n7574), .ZN(n7769) );
  MUX2_X1 U9671 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n7602), .Z(n7576) );
  OAI21_X1 U9672 ( .B1(n7576), .B2(SI_7_), .A(n7578), .ZN(n7577) );
  INV_X1 U9673 ( .A(n7577), .ZN(n7784) );
  MUX2_X1 U9674 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n7602), .Z(n7579) );
  OAI21_X1 U9675 ( .B1(SI_8_), .B2(n7579), .A(n7581), .ZN(n7580) );
  INV_X1 U9676 ( .A(n7580), .ZN(n7799) );
  MUX2_X1 U9677 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n7602), .Z(n7582) );
  OAI21_X1 U9678 ( .B1(n7582), .B2(SI_9_), .A(n7584), .ZN(n7583) );
  INV_X1 U9679 ( .A(n7583), .ZN(n7815) );
  MUX2_X1 U9680 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n7602), .Z(n7831) );
  MUX2_X1 U9681 ( .A(n10070), .B(n10069), .S(n8538), .Z(n7588) );
  INV_X1 U9682 ( .A(SI_11_), .ZN(n7587) );
  NAND2_X1 U9683 ( .A1(n7588), .A2(n7587), .ZN(n7589) );
  INV_X1 U9684 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n8740) );
  INV_X1 U9685 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n10122) );
  MUX2_X1 U9686 ( .A(n8740), .B(n10122), .S(n7602), .Z(n7592) );
  NAND2_X1 U9687 ( .A1(n7865), .A2(n7864), .ZN(n7594) );
  INV_X1 U9688 ( .A(SI_12_), .ZN(n7591) );
  NAND2_X1 U9689 ( .A1(n7592), .A2(n7591), .ZN(n7593) );
  INV_X1 U9690 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n10190) );
  MUX2_X1 U9691 ( .A(n15454), .B(n10190), .S(n7602), .Z(n7595) );
  INV_X1 U9692 ( .A(SI_13_), .ZN(n9909) );
  NAND2_X1 U9693 ( .A1(n7595), .A2(n9909), .ZN(n7596) );
  INV_X1 U9694 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10453) );
  INV_X1 U9695 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n10455) );
  MUX2_X1 U9696 ( .A(n10453), .B(n10455), .S(n7602), .Z(n7899) );
  NAND2_X1 U9697 ( .A1(n7916), .A2(SI_14_), .ZN(n7598) );
  INV_X1 U9698 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10558) );
  INV_X1 U9699 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n10559) );
  MUX2_X1 U9700 ( .A(n10558), .B(n10559), .S(n7602), .Z(n7918) );
  INV_X1 U9701 ( .A(n7918), .ZN(n7597) );
  NAND2_X1 U9702 ( .A1(n7597), .A2(SI_15_), .ZN(n7599) );
  NOR2_X1 U9703 ( .A1(n7916), .A2(SI_14_), .ZN(n7600) );
  INV_X1 U9704 ( .A(SI_15_), .ZN(n10104) );
  AOI22_X1 U9705 ( .A1(n7600), .A2(n7599), .B1(n10104), .B2(n7918), .ZN(n7601)
         );
  INV_X1 U9706 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n10421) );
  INV_X1 U9707 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n10424) );
  MUX2_X1 U9708 ( .A(n10421), .B(n10424), .S(n8538), .Z(n7604) );
  XNOR2_X1 U9709 ( .A(n7604), .B(SI_16_), .ZN(n7939) );
  NAND2_X1 U9710 ( .A1(n7940), .A2(n7939), .ZN(n7606) );
  INV_X1 U9711 ( .A(SI_16_), .ZN(n7603) );
  NAND2_X1 U9712 ( .A1(n7604), .A2(n7603), .ZN(n7605) );
  INV_X1 U9713 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n10508) );
  INV_X1 U9714 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n8832) );
  INV_X4 U9715 ( .A(n9769), .ZN(n8538) );
  MUX2_X1 U9716 ( .A(n10508), .B(n8832), .S(n8538), .Z(n7956) );
  NOR2_X1 U9717 ( .A1(n7608), .A2(SI_17_), .ZN(n7607) );
  NAND2_X1 U9718 ( .A1(n7608), .A2(SI_17_), .ZN(n7609) );
  INV_X1 U9719 ( .A(SI_18_), .ZN(n10427) );
  MUX2_X1 U9720 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(P1_DATAO_REG_18__SCAN_IN), 
        .S(n8538), .Z(n7984) );
  INV_X1 U9721 ( .A(n7984), .ZN(n7610) );
  MUX2_X1 U9722 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(P1_DATAO_REG_19__SCAN_IN), 
        .S(n8538), .Z(n7611) );
  NAND2_X1 U9723 ( .A1(n7611), .A2(SI_19_), .ZN(n7990) );
  OAI21_X1 U9724 ( .B1(n10427), .B2(n7610), .A(n7990), .ZN(n7616) );
  NOR2_X1 U9725 ( .A1(n7984), .A2(SI_18_), .ZN(n7614) );
  INV_X1 U9726 ( .A(n7611), .ZN(n7612) );
  INV_X1 U9727 ( .A(SI_19_), .ZN(n10476) );
  NAND2_X1 U9728 ( .A1(n7612), .A2(n10476), .ZN(n7989) );
  INV_X1 U9729 ( .A(n7989), .ZN(n7613) );
  AOI21_X1 U9730 ( .B1(n7614), .B2(n7990), .A(n7613), .ZN(n7615) );
  INV_X1 U9731 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n15251) );
  INV_X1 U9732 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n15400) );
  MUX2_X1 U9733 ( .A(n15251), .B(n15400), .S(n8538), .Z(n8012) );
  INV_X1 U9734 ( .A(n8012), .ZN(n8022) );
  MUX2_X1 U9735 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n8538), .Z(n8027) );
  INV_X1 U9736 ( .A(SI_20_), .ZN(n10802) );
  NOR2_X1 U9737 ( .A1(n8012), .A2(n10802), .ZN(n7617) );
  AOI22_X1 U9738 ( .A1(n7617), .A2(n7535), .B1(n8027), .B2(SI_21_), .ZN(n7618)
         );
  MUX2_X1 U9739 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(P1_DATAO_REG_22__SCAN_IN), 
        .S(n8538), .Z(n9443) );
  MUX2_X1 U9740 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n8538), .Z(n7623) );
  MUX2_X1 U9741 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n8538), .Z(n7625) );
  XNOR2_X1 U9742 ( .A(n7625), .B(SI_24_), .ZN(n8062) );
  NAND2_X1 U9743 ( .A1(n7625), .A2(SI_24_), .ZN(n7626) );
  INV_X1 U9744 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n11651) );
  MUX2_X1 U9745 ( .A(n8965), .B(n11651), .S(n8538), .Z(n7628) );
  INV_X1 U9746 ( .A(SI_25_), .ZN(n11801) );
  NAND2_X1 U9747 ( .A1(n7628), .A2(n11801), .ZN(n7631) );
  INV_X1 U9748 ( .A(n7628), .ZN(n7629) );
  NAND2_X1 U9749 ( .A1(n7629), .A2(SI_25_), .ZN(n7630) );
  NAND2_X1 U9750 ( .A1(n7631), .A2(n7630), .ZN(n8078) );
  OAI21_X2 U9751 ( .B1(n8079), .B2(n8078), .A(n7631), .ZN(n8093) );
  INV_X1 U9752 ( .A(SI_26_), .ZN(n13216) );
  INV_X1 U9753 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n11821) );
  INV_X1 U9754 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n11817) );
  MUX2_X1 U9755 ( .A(n11821), .B(n11817), .S(n8538), .Z(n8091) );
  MUX2_X1 U9756 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(P1_DATAO_REG_27__SCAN_IN), 
        .S(n8538), .Z(n8108) );
  NOR2_X1 U9757 ( .A1(n8108), .A2(SI_27_), .ZN(n7632) );
  INV_X1 U9758 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n12607) );
  INV_X1 U9759 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n13779) );
  MUX2_X1 U9760 ( .A(n12607), .B(n13779), .S(n8538), .Z(n7633) );
  INV_X1 U9761 ( .A(SI_28_), .ZN(n13206) );
  NAND2_X1 U9762 ( .A1(n7633), .A2(n13206), .ZN(n8129) );
  INV_X1 U9763 ( .A(n7633), .ZN(n7634) );
  NAND2_X1 U9764 ( .A1(n7634), .A2(SI_28_), .ZN(n7635) );
  NAND2_X1 U9765 ( .A1(n8129), .A2(n7635), .ZN(n7638) );
  NAND2_X1 U9766 ( .A1(n7639), .A2(n7638), .ZN(n7640) );
  NOR2_X1 U9767 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n7644) );
  AND4_X2 U9768 ( .A1(n7644), .A2(n7643), .A3(n7642), .A4(n7641), .ZN(n7649)
         );
  AND2_X2 U9769 ( .A1(n7684), .A2(n7645), .ZN(n7743) );
  INV_X2 U9770 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n7850) );
  AND4_X2 U9771 ( .A1(n7850), .A2(n7647), .A3(n7849), .A4(n7646), .ZN(n7648)
         );
  INV_X1 U9772 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n7650) );
  INV_X1 U9773 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n8202) );
  NAND4_X1 U9774 ( .A1(n7372), .A2(n7650), .A3(n8216), .A4(n8202), .ZN(n7651)
         );
  NOR2_X1 U9775 ( .A1(n7652), .A2(n7651), .ZN(n7653) );
  INV_X1 U9776 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n7655) );
  INV_X1 U9777 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n7656) );
  INV_X1 U9778 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n7657) );
  NAND2_X1 U9779 ( .A1(n13776), .A2(n8418), .ZN(n7660) );
  OR2_X1 U9780 ( .A1(n8419), .A2(n12607), .ZN(n7659) );
  INV_X1 U9781 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n7661) );
  INV_X2 U9782 ( .A(n7723), .ZN(n7697) );
  NAND2_X1 U9783 ( .A1(n7697), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n7675) );
  INV_X1 U9784 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n8504) );
  OR2_X1 U9785 ( .A1(n8385), .A2(n8504), .ZN(n7674) );
  NAND2_X1 U9786 ( .A1(n7776), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n7807) );
  NAND2_X1 U9787 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_REG3_REG_7__SCAN_IN), 
        .ZN(n7665) );
  NAND2_X1 U9788 ( .A1(n7823), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7839) );
  INV_X1 U9789 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n7838) );
  INV_X1 U9790 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n11549) );
  INV_X1 U9791 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n7870) );
  NAND2_X1 U9792 ( .A1(n7890), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n7905) );
  INV_X1 U9793 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n7904) );
  INV_X1 U9794 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n7928) );
  NAND2_X1 U9795 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_REG3_REG_19__SCAN_IN), 
        .ZN(n7666) );
  INV_X1 U9796 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n13859) );
  NAND2_X1 U9797 ( .A1(n8015), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n8044) );
  INV_X1 U9798 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n13869) );
  INV_X1 U9799 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n13792) );
  NAND2_X1 U9800 ( .A1(n8066), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n8067) );
  NAND2_X1 U9801 ( .A1(P1_REG3_REG_25__SCAN_IN), .A2(n8082), .ZN(n8097) );
  INV_X1 U9802 ( .A(n8097), .ZN(n7667) );
  NAND2_X1 U9803 ( .A1(n7667), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n8117) );
  INV_X1 U9804 ( .A(n8117), .ZN(n7668) );
  NAND2_X1 U9805 ( .A1(n7668), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n8119) );
  INV_X1 U9806 ( .A(n8119), .ZN(n7669) );
  NAND2_X1 U9807 ( .A1(n7669), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n12594) );
  INV_X1 U9808 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n7670) );
  NAND2_X1 U9809 ( .A1(n8119), .A2(n7670), .ZN(n7671) );
  NAND2_X1 U9810 ( .A1(n12594), .A2(n7671), .ZN(n14082) );
  OR2_X1 U9811 ( .A1(n8134), .A2(n14082), .ZN(n7673) );
  INV_X1 U9812 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n9621) );
  OR2_X1 U9813 ( .A1(n8115), .A2(n9621), .ZN(n7672) );
  NAND4_X1 U9814 ( .A1(n7675), .A2(n7674), .A3(n7673), .A4(n7672), .ZN(n13918)
         );
  INV_X1 U9815 ( .A(n13918), .ZN(n8128) );
  NAND2_X1 U9816 ( .A1(n7697), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n7678) );
  INV_X1 U9817 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n7676) );
  OR2_X1 U9818 ( .A1(n7699), .A2(n7676), .ZN(n7677) );
  INV_X1 U9819 ( .A(n7679), .ZN(n7680) );
  NAND2_X1 U9820 ( .A1(n7681), .A2(n7680), .ZN(n7682) );
  NAND2_X1 U9821 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n7683) );
  MUX2_X1 U9822 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7683), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n7687) );
  INV_X1 U9823 ( .A(n7685), .ZN(n7686) );
  NAND2_X1 U9824 ( .A1(n7687), .A2(n7686), .ZN(n9934) );
  OR2_X1 U9825 ( .A1(n7716), .A2(n9934), .ZN(n7688) );
  NAND2_X1 U9826 ( .A1(n7697), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n7694) );
  INV_X1 U9827 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n7690) );
  INV_X1 U9828 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n7691) );
  INV_X1 U9829 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n7692) );
  OR2_X1 U9830 ( .A1(n7699), .A2(n7692), .ZN(n7693) );
  NOR2_X1 U9831 ( .A1(n8538), .A2(n7695), .ZN(n7696) );
  XNOR2_X1 U9832 ( .A(n7696), .B(n15478), .ZN(n14440) );
  NAND2_X1 U9833 ( .A1(n7697), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n7701) );
  INV_X1 U9834 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n7698) );
  OR2_X1 U9835 ( .A1(n7699), .A2(n7698), .ZN(n7700) );
  INV_X1 U9836 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n7702) );
  OR2_X1 U9837 ( .A1(n8134), .A2(n7702), .ZN(n7705) );
  INV_X1 U9838 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n9918) );
  OR2_X1 U9839 ( .A1(n8115), .A2(n9918), .ZN(n7704) );
  NAND3_X1 U9840 ( .A1(n7542), .A2(n7705), .A3(n7704), .ZN(n10363) );
  INV_X1 U9841 ( .A(n7706), .ZN(n7708) );
  NAND2_X1 U9842 ( .A1(n7708), .A2(n7707), .ZN(n7710) );
  NAND2_X1 U9843 ( .A1(n7710), .A2(n7709), .ZN(n9797) );
  INV_X1 U9844 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n9754) );
  NOR2_X1 U9845 ( .A1(n7685), .A2(n7655), .ZN(n7712) );
  MUX2_X1 U9846 ( .A(n7655), .B(n7712), .S(P1_IR_REG_2__SCAN_IN), .Z(n7713) );
  INV_X1 U9847 ( .A(n7713), .ZN(n7715) );
  INV_X1 U9848 ( .A(n7743), .ZN(n7714) );
  NAND2_X1 U9849 ( .A1(n7715), .A2(n7714), .ZN(n14727) );
  OR2_X1 U9850 ( .A1(n7716), .A2(n14727), .ZN(n7717) );
  NAND2_X1 U9851 ( .A1(n13808), .A2(n10519), .ZN(n7718) );
  INV_X1 U9852 ( .A(n10363), .ZN(n14771) );
  NAND2_X1 U9853 ( .A1(n14771), .A2(n13884), .ZN(n8171) );
  NAND2_X1 U9854 ( .A1(n7719), .A2(n8168), .ZN(n10180) );
  NAND2_X1 U9855 ( .A1(n14771), .A2(n10519), .ZN(n8257) );
  NAND2_X1 U9856 ( .A1(n10180), .A2(n8257), .ZN(n10299) );
  INV_X1 U9857 ( .A(n8115), .ZN(n8069) );
  NAND2_X1 U9858 ( .A1(n8069), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n7722) );
  INV_X1 U9859 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n7720) );
  OR2_X1 U9860 ( .A1(n8385), .A2(n7720), .ZN(n7721) );
  OR2_X1 U9861 ( .A1(n8134), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n7725) );
  INV_X1 U9862 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n10521) );
  OR2_X1 U9863 ( .A1(n8384), .A2(n10521), .ZN(n7724) );
  INV_X2 U9864 ( .A(n7727), .ZN(n8000) );
  INV_X2 U9865 ( .A(n7716), .ZN(n7999) );
  OR2_X1 U9866 ( .A1(n7743), .A2(n7655), .ZN(n7728) );
  XNOR2_X1 U9867 ( .A(n7728), .B(P1_IR_REG_3__SCAN_IN), .ZN(n13957) );
  AOI22_X1 U9868 ( .A1(n6553), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(n7999), .B2(
        n13957), .ZN(n7732) );
  XNOR2_X1 U9869 ( .A(n7730), .B(n7729), .ZN(n9755) );
  NAND2_X1 U9870 ( .A1(n9755), .A2(n8418), .ZN(n7731) );
  NAND2_X1 U9871 ( .A1(n10299), .A2(n10300), .ZN(n10298) );
  NAND2_X1 U9872 ( .A1(n7733), .A2(n7734), .ZN(n7735) );
  NAND2_X1 U9873 ( .A1(n8133), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n7739) );
  INV_X1 U9874 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n10640) );
  OR2_X1 U9875 ( .A1(n8384), .A2(n10640), .ZN(n7738) );
  XNOR2_X1 U9876 ( .A(P1_REG3_REG_3__SCAN_IN), .B(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n10641) );
  OR2_X1 U9877 ( .A1(n8134), .A2(n10641), .ZN(n7737) );
  INV_X1 U9878 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n9922) );
  OR2_X1 U9879 ( .A1(n8115), .A2(n9922), .ZN(n7736) );
  INV_X1 U9880 ( .A(n13938), .ZN(n10493) );
  XNOR2_X1 U9881 ( .A(n7741), .B(n7740), .ZN(n9767) );
  NAND2_X1 U9882 ( .A1(n9767), .A2(n8418), .ZN(n7746) );
  INV_X1 U9883 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n7742) );
  NAND2_X1 U9884 ( .A1(n7743), .A2(n7742), .ZN(n7751) );
  NAND2_X1 U9885 ( .A1(n7751), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7744) );
  XNOR2_X1 U9886 ( .A(n7744), .B(P1_IR_REG_4__SCAN_IN), .ZN(n13977) );
  AOI22_X1 U9887 ( .A1(n8000), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n7999), .B2(
        n13977), .ZN(n7745) );
  NAND2_X1 U9888 ( .A1(n7746), .A2(n7745), .ZN(n10631) );
  NAND2_X1 U9889 ( .A1(n10493), .A2(n10631), .ZN(n8173) );
  NAND2_X1 U9890 ( .A1(n10642), .A2(n13938), .ZN(n7747) );
  OR2_X1 U9891 ( .A1(n10631), .A2(n13938), .ZN(n10495) );
  NAND2_X1 U9892 ( .A1(n10497), .A2(n10495), .ZN(n7768) );
  OR2_X1 U9893 ( .A1(n9796), .A2(n7711), .ZN(n7759) );
  NAND2_X1 U9894 ( .A1(n7753), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7752) );
  MUX2_X1 U9895 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7752), .S(
        P1_IR_REG_5__SCAN_IN), .Z(n7756) );
  INV_X1 U9896 ( .A(n7753), .ZN(n7755) );
  INV_X1 U9897 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n7754) );
  NAND2_X1 U9898 ( .A1(n7755), .A2(n7754), .ZN(n7788) );
  NAND2_X1 U9899 ( .A1(n7756), .A2(n7788), .ZN(n9953) );
  INV_X1 U9900 ( .A(n9953), .ZN(n7757) );
  AOI22_X1 U9901 ( .A1(n8000), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n7999), .B2(
        n7757), .ZN(n7758) );
  NAND2_X1 U9902 ( .A1(n7759), .A2(n7758), .ZN(n10744) );
  AOI21_X1 U9903 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(P1_REG3_REG_5__SCAN_IN), .ZN(n7761) );
  NOR2_X1 U9904 ( .A1(n7761), .A2(n7776), .ZN(n10704) );
  NAND2_X1 U9905 ( .A1(n7760), .A2(n10704), .ZN(n7767) );
  INV_X1 U9906 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n7762) );
  OR2_X1 U9907 ( .A1(n8385), .A2(n7762), .ZN(n7766) );
  INV_X1 U9908 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n7763) );
  OR2_X1 U9909 ( .A1(n8384), .A2(n7763), .ZN(n7765) );
  INV_X1 U9910 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n9923) );
  OR2_X1 U9911 ( .A1(n8115), .A2(n9923), .ZN(n7764) );
  NAND4_X1 U9912 ( .A1(n7767), .A2(n7766), .A3(n7765), .A4(n7764), .ZN(n13937)
         );
  INV_X1 U9913 ( .A(n13937), .ZN(n10540) );
  NAND2_X1 U9914 ( .A1(n10744), .A2(n10540), .ZN(n8174) );
  OAI21_X1 U9915 ( .B1(n10744), .B2(n10540), .A(n8174), .ZN(n8435) );
  NAND2_X1 U9916 ( .A1(n7768), .A2(n8435), .ZN(n10494) );
  NAND2_X1 U9917 ( .A1(n7016), .A2(n10540), .ZN(n10542) );
  NAND2_X1 U9918 ( .A1(n10494), .A2(n10542), .ZN(n7783) );
  OR2_X1 U9919 ( .A1(n7770), .A2(n7769), .ZN(n7771) );
  NAND2_X1 U9920 ( .A1(n7772), .A2(n7771), .ZN(n9802) );
  OR2_X1 U9921 ( .A1(n9802), .A2(n7711), .ZN(n7775) );
  NAND2_X1 U9922 ( .A1(n7788), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7773) );
  XNOR2_X1 U9923 ( .A(n7773), .B(P1_IR_REG_6__SCAN_IN), .ZN(n13989) );
  AOI22_X1 U9924 ( .A1(n8000), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n7999), .B2(
        n13989), .ZN(n7774) );
  NAND2_X1 U9925 ( .A1(n8133), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n7780) );
  INV_X1 U9926 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n10748) );
  OR2_X1 U9927 ( .A1(n8384), .A2(n10748), .ZN(n7779) );
  OAI21_X1 U9928 ( .B1(n7776), .B2(P1_REG3_REG_6__SCAN_IN), .A(n7807), .ZN(
        n10762) );
  OR2_X1 U9929 ( .A1(n8134), .A2(n10762), .ZN(n7778) );
  INV_X1 U9930 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n9924) );
  OR2_X1 U9931 ( .A1(n8115), .A2(n9924), .ZN(n7777) );
  NAND4_X1 U9932 ( .A1(n7780), .A2(n7779), .A3(n7778), .A4(n7777), .ZN(n13936)
         );
  INV_X1 U9933 ( .A(n13936), .ZN(n10597) );
  OR2_X1 U9934 ( .A1(n10767), .A2(n10597), .ZN(n7781) );
  NAND2_X1 U9935 ( .A1(n10767), .A2(n10597), .ZN(n10589) );
  INV_X1 U9936 ( .A(n10543), .ZN(n7782) );
  NAND2_X1 U9937 ( .A1(n7783), .A2(n7782), .ZN(n10541) );
  OR2_X1 U9938 ( .A1(n10767), .A2(n13936), .ZN(n10593) );
  NAND2_X1 U9939 ( .A1(n10541), .A2(n10593), .ZN(n7797) );
  OR2_X1 U9940 ( .A1(n7785), .A2(n7784), .ZN(n7786) );
  NAND2_X1 U9941 ( .A1(n7787), .A2(n7786), .ZN(n9799) );
  OR2_X1 U9942 ( .A1(n9799), .A2(n7711), .ZN(n7790) );
  NAND2_X1 U9943 ( .A1(n7853), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7804) );
  XNOR2_X1 U9944 ( .A(n7804), .B(P1_IR_REG_7__SCAN_IN), .ZN(n9941) );
  AOI22_X1 U9945 ( .A1(n8000), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n7999), .B2(
        n9941), .ZN(n7789) );
  NAND2_X1 U9946 ( .A1(n7790), .A2(n7789), .ZN(n10969) );
  NAND2_X1 U9947 ( .A1(n8133), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n7796) );
  INV_X1 U9948 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n7791) );
  OR2_X1 U9949 ( .A1(n8384), .A2(n7791), .ZN(n7795) );
  INV_X1 U9950 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n7792) );
  XNOR2_X1 U9951 ( .A(n7807), .B(n7792), .ZN(n10972) );
  OR2_X1 U9952 ( .A1(n8134), .A2(n10972), .ZN(n7794) );
  INV_X1 U9953 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n9926) );
  OR2_X1 U9954 ( .A1(n8115), .A2(n9926), .ZN(n7793) );
  NAND4_X1 U9955 ( .A1(n7796), .A2(n7795), .A3(n7794), .A4(n7793), .ZN(n13935)
         );
  XNOR2_X1 U9956 ( .A(n10969), .B(n13935), .ZN(n10594) );
  INV_X1 U9957 ( .A(n10594), .ZN(n10590) );
  OR2_X1 U9958 ( .A1(n10969), .A2(n13935), .ZN(n7798) );
  OR2_X1 U9959 ( .A1(n7800), .A2(n7799), .ZN(n7801) );
  OR2_X1 U9960 ( .A1(n9835), .A2(n7711), .ZN(n7806) );
  NAND2_X1 U9961 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n7803) );
  NAND2_X1 U9962 ( .A1(n7804), .A2(n7803), .ZN(n7819) );
  XNOR2_X1 U9963 ( .A(n7819), .B(n7850), .ZN(n9971) );
  AOI22_X1 U9964 ( .A1(n8000), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n7999), .B2(
        n9971), .ZN(n7805) );
  NAND2_X1 U9965 ( .A1(n7806), .A2(n7805), .ZN(n11164) );
  NAND2_X1 U9966 ( .A1(n8133), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n7813) );
  INV_X1 U9967 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n9942) );
  OR2_X1 U9968 ( .A1(n8384), .A2(n9942), .ZN(n7812) );
  INV_X1 U9969 ( .A(n7807), .ZN(n7808) );
  AOI21_X1 U9970 ( .B1(n7808), .B2(P1_REG3_REG_7__SCAN_IN), .A(
        P1_REG3_REG_8__SCAN_IN), .ZN(n7809) );
  OR2_X1 U9971 ( .A1(n7809), .A2(n7823), .ZN(n11162) );
  OR2_X1 U9972 ( .A1(n8134), .A2(n11162), .ZN(n7811) );
  INV_X1 U9973 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9965) );
  OR2_X1 U9974 ( .A1(n8115), .A2(n9965), .ZN(n7810) );
  NAND4_X1 U9975 ( .A1(n7813), .A2(n7812), .A3(n7811), .A4(n7810), .ZN(n13934)
         );
  XNOR2_X1 U9976 ( .A(n11164), .B(n13934), .ZN(n8439) );
  NAND2_X1 U9977 ( .A1(n10813), .A2(n10812), .ZN(n10811) );
  OR2_X1 U9978 ( .A1(n11164), .A2(n13934), .ZN(n7814) );
  NAND2_X1 U9979 ( .A1(n10811), .A2(n7814), .ZN(n11022) );
  NAND2_X1 U9980 ( .A1(n7818), .A2(n7817), .ZN(n9839) );
  OR2_X1 U9981 ( .A1(n9839), .A2(n7711), .ZN(n7822) );
  NAND2_X1 U9982 ( .A1(n7820), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7833) );
  XNOR2_X1 U9983 ( .A(n7833), .B(P1_IR_REG_9__SCAN_IN), .ZN(n9972) );
  AOI22_X1 U9984 ( .A1(n8000), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n7999), .B2(
        n9972), .ZN(n7821) );
  NAND2_X1 U9985 ( .A1(n8133), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n7828) );
  INV_X1 U9986 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n11025) );
  OR2_X1 U9987 ( .A1(n8384), .A2(n11025), .ZN(n7827) );
  OR2_X1 U9988 ( .A1(n7823), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7824) );
  NAND2_X1 U9989 ( .A1(n7839), .A2(n7824), .ZN(n11238) );
  OR2_X1 U9990 ( .A1(n8134), .A2(n11238), .ZN(n7826) );
  INV_X1 U9991 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10160) );
  OR2_X1 U9992 ( .A1(n8115), .A2(n10160), .ZN(n7825) );
  NAND4_X1 U9993 ( .A1(n7828), .A2(n7827), .A3(n7826), .A4(n7825), .ZN(n13933)
         );
  INV_X1 U9994 ( .A(n13933), .ZN(n11230) );
  XNOR2_X1 U9995 ( .A(n11232), .B(n11230), .ZN(n11021) );
  NAND2_X1 U9996 ( .A1(n11022), .A2(n11021), .ZN(n11020) );
  OR2_X1 U9997 ( .A1(n11232), .A2(n13933), .ZN(n7829) );
  XNOR2_X1 U9998 ( .A(n7831), .B(SI_10_), .ZN(n7832) );
  XNOR2_X1 U9999 ( .A(n7830), .B(n7832), .ZN(n9911) );
  NAND2_X1 U10000 ( .A1(n9911), .A2(n8418), .ZN(n7837) );
  INV_X1 U10001 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n7851) );
  NAND2_X1 U10002 ( .A1(n7833), .A2(n7851), .ZN(n7834) );
  NAND2_X1 U10003 ( .A1(n7834), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7835) );
  XNOR2_X1 U10004 ( .A(n7835), .B(P1_IR_REG_10__SCAN_IN), .ZN(n10167) );
  AOI22_X1 U10005 ( .A1(n10167), .A2(n7999), .B1(n8000), .B2(
        P2_DATAO_REG_10__SCAN_IN), .ZN(n7836) );
  NAND2_X1 U10006 ( .A1(n8133), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n7844) );
  INV_X1 U10007 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n11188) );
  OR2_X1 U10008 ( .A1(n8384), .A2(n11188), .ZN(n7843) );
  NAND2_X1 U10009 ( .A1(n7839), .A2(n7838), .ZN(n7840) );
  NAND2_X1 U10010 ( .A1(n7857), .A2(n7840), .ZN(n11377) );
  OR2_X1 U10011 ( .A1(n8134), .A2(n11377), .ZN(n7842) );
  INV_X1 U10012 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n10161) );
  OR2_X1 U10013 ( .A1(n8115), .A2(n10161), .ZN(n7841) );
  NAND4_X1 U10014 ( .A1(n7844), .A2(n7843), .A3(n7842), .A4(n7841), .ZN(n13932) );
  XNOR2_X1 U10015 ( .A(n11373), .B(n11550), .ZN(n11186) );
  OR2_X1 U10016 ( .A1(n11373), .A2(n13932), .ZN(n7845) );
  XNOR2_X1 U10017 ( .A(n7847), .B(n7846), .ZN(n10068) );
  NAND2_X1 U10018 ( .A1(n10068), .A2(n8418), .ZN(n7856) );
  INV_X1 U10019 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n7848) );
  NAND4_X1 U10020 ( .A1(n7851), .A2(n7850), .A3(n7849), .A4(n7848), .ZN(n7852)
         );
  NAND2_X1 U10021 ( .A1(n7866), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7854) );
  XNOR2_X1 U10022 ( .A(n7854), .B(P1_IR_REG_11__SCAN_IN), .ZN(n10402) );
  AOI22_X1 U10023 ( .A1(n8000), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n7999), 
        .B2(n10402), .ZN(n7855) );
  NAND2_X1 U10024 ( .A1(n8133), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n7862) );
  INV_X1 U10025 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n11284) );
  OR2_X1 U10026 ( .A1(n8384), .A2(n11284), .ZN(n7861) );
  INV_X1 U10027 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n10399) );
  OR2_X1 U10028 ( .A1(n8115), .A2(n10399), .ZN(n7860) );
  NAND2_X1 U10029 ( .A1(n7857), .A2(n11549), .ZN(n7858) );
  NAND2_X1 U10030 ( .A1(n7871), .A2(n7858), .ZN(n11553) );
  OR2_X1 U10031 ( .A1(n8134), .A2(n11553), .ZN(n7859) );
  NAND4_X1 U10032 ( .A1(n7862), .A2(n7861), .A3(n7860), .A4(n7859), .ZN(n13931) );
  OR2_X1 U10033 ( .A1(n11555), .A2(n13931), .ZN(n11460) );
  NAND2_X1 U10034 ( .A1(n11555), .A2(n13931), .ZN(n7863) );
  XNOR2_X1 U10035 ( .A(n7865), .B(n7864), .ZN(n10082) );
  NAND2_X1 U10036 ( .A1(n10082), .A2(n8418), .ZN(n7869) );
  NAND2_X1 U10037 ( .A1(n7867), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7883) );
  XNOR2_X1 U10038 ( .A(n7883), .B(P1_IR_REG_12__SCAN_IN), .ZN(n10566) );
  AOI22_X1 U10039 ( .A1(n8000), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n7999), 
        .B2(n10566), .ZN(n7868) );
  NAND2_X1 U10040 ( .A1(n8133), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n7877) );
  INV_X1 U10041 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n11472) );
  OR2_X1 U10042 ( .A1(n8384), .A2(n11472), .ZN(n7876) );
  AND2_X1 U10043 ( .A1(n7871), .A2(n7870), .ZN(n7872) );
  OR2_X1 U10044 ( .A1(n7872), .A2(n7890), .ZN(n11602) );
  OR2_X1 U10045 ( .A1(n8134), .A2(n11602), .ZN(n7875) );
  INV_X1 U10046 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n7873) );
  OR2_X1 U10047 ( .A1(n8115), .A2(n7873), .ZN(n7874) );
  NAND4_X1 U10048 ( .A1(n7877), .A2(n7876), .A3(n7875), .A4(n7874), .ZN(n13930) );
  XNOR2_X1 U10049 ( .A(n11599), .B(n13930), .ZN(n11464) );
  INV_X1 U10050 ( .A(n11464), .ZN(n7878) );
  OR2_X1 U10051 ( .A1(n11599), .A2(n13930), .ZN(n7879) );
  XNOR2_X1 U10052 ( .A(n7881), .B(n7880), .ZN(n10189) );
  NAND2_X1 U10053 ( .A1(n10189), .A2(n8418), .ZN(n7889) );
  INV_X1 U10054 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n7882) );
  AOI21_X1 U10055 ( .B1(n7883), .B2(n7882), .A(n7655), .ZN(n7884) );
  NAND2_X1 U10056 ( .A1(n7884), .A2(P1_IR_REG_13__SCAN_IN), .ZN(n7887) );
  INV_X1 U10057 ( .A(n7884), .ZN(n7886) );
  INV_X1 U10058 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n7885) );
  NAND2_X1 U10059 ( .A1(n7886), .A2(n7885), .ZN(n7900) );
  AOI22_X1 U10060 ( .A1(n7999), .A2(n10672), .B1(n8000), .B2(
        P2_DATAO_REG_13__SCAN_IN), .ZN(n7888) );
  NAND2_X1 U10061 ( .A1(n7697), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n7897) );
  OR2_X1 U10062 ( .A1(n7890), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n7891) );
  NAND2_X1 U10063 ( .A1(n7905), .A2(n7891), .ZN(n11739) );
  OR2_X1 U10064 ( .A1(n8134), .A2(n11739), .ZN(n7896) );
  INV_X1 U10065 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n7892) );
  OR2_X1 U10066 ( .A1(n8115), .A2(n7892), .ZN(n7895) );
  INV_X1 U10067 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n7893) );
  OR2_X1 U10068 ( .A1(n8385), .A2(n7893), .ZN(n7894) );
  NAND4_X1 U10069 ( .A1(n7897), .A2(n7896), .A3(n7895), .A4(n7894), .ZN(n13929) );
  XNOR2_X1 U10070 ( .A(n11736), .B(n13929), .ZN(n11351) );
  INV_X1 U10071 ( .A(n11351), .ZN(n11353) );
  OR2_X1 U10072 ( .A1(n11736), .A2(n13929), .ZN(n7898) );
  XNOR2_X1 U10073 ( .A(n7913), .B(n7899), .ZN(n10452) );
  NAND2_X1 U10074 ( .A1(n10452), .A2(n8418), .ZN(n7903) );
  NAND2_X1 U10075 ( .A1(n7900), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7901) );
  XNOR2_X1 U10076 ( .A(n7901), .B(P1_IR_REG_14__SCAN_IN), .ZN(n11319) );
  AOI22_X1 U10077 ( .A1(n11319), .A2(n7999), .B1(n8000), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n7902) );
  NAND2_X1 U10078 ( .A1(n7697), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n7910) );
  NAND2_X1 U10079 ( .A1(n7905), .A2(n7904), .ZN(n7906) );
  NAND2_X1 U10080 ( .A1(n7929), .A2(n7906), .ZN(n14683) );
  OR2_X1 U10081 ( .A1(n8134), .A2(n14683), .ZN(n7909) );
  INV_X1 U10082 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n11773) );
  OR2_X1 U10083 ( .A1(n8115), .A2(n11773), .ZN(n7908) );
  INV_X1 U10084 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n11776) );
  OR2_X1 U10085 ( .A1(n8385), .A2(n11776), .ZN(n7907) );
  NAND4_X1 U10086 ( .A1(n7910), .A2(n7909), .A3(n7908), .A4(n7907), .ZN(n13928) );
  INV_X1 U10087 ( .A(n13928), .ZN(n13906) );
  NAND2_X1 U10088 ( .A1(n14680), .A2(n13906), .ZN(n8308) );
  NAND2_X1 U10089 ( .A1(n14680), .A2(n13928), .ZN(n7912) );
  INV_X1 U10090 ( .A(n7913), .ZN(n7917) );
  INV_X1 U10091 ( .A(n7914), .ZN(n7915) );
  XNOR2_X1 U10092 ( .A(n7918), .B(SI_15_), .ZN(n7919) );
  XNOR2_X1 U10093 ( .A(n7920), .B(n7919), .ZN(n10557) );
  NAND2_X1 U10094 ( .A1(n10557), .A2(n8418), .ZN(n7926) );
  NAND2_X1 U10095 ( .A1(n7921), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7922) );
  MUX2_X1 U10096 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7922), .S(
        P1_IR_REG_15__SCAN_IN), .Z(n7924) );
  AND2_X1 U10097 ( .A1(n7924), .A2(n7923), .ZN(n11327) );
  AOI22_X1 U10098 ( .A1(n8000), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n7999), 
        .B2(n11327), .ZN(n7925) );
  NAND2_X1 U10099 ( .A1(n7697), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n7935) );
  INV_X1 U10100 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n14740) );
  OR2_X1 U10101 ( .A1(n8115), .A2(n14740), .ZN(n7934) );
  INV_X1 U10102 ( .A(n7927), .ZN(n7946) );
  NAND2_X1 U10103 ( .A1(n7929), .A2(n7928), .ZN(n7930) );
  NAND2_X1 U10104 ( .A1(n7946), .A2(n7930), .ZN(n13909) );
  OR2_X1 U10105 ( .A1(n8134), .A2(n13909), .ZN(n7933) );
  INV_X1 U10106 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n7931) );
  OR2_X1 U10107 ( .A1(n8385), .A2(n7931), .ZN(n7932) );
  NAND4_X1 U10108 ( .A1(n7935), .A2(n7934), .A3(n7933), .A4(n7932), .ZN(n13927) );
  INV_X1 U10109 ( .A(n13927), .ZN(n14666) );
  NAND2_X1 U10110 ( .A1(n14373), .A2(n14666), .ZN(n8320) );
  NAND2_X1 U10111 ( .A1(n8319), .A2(n8320), .ZN(n11675) );
  INV_X1 U10112 ( .A(n11675), .ZN(n7936) );
  OR2_X1 U10113 ( .A1(n14373), .A2(n13927), .ZN(n7937) );
  XNOR2_X1 U10114 ( .A(n7940), .B(n7939), .ZN(n10420) );
  NAND2_X1 U10115 ( .A1(n10420), .A2(n8418), .ZN(n7943) );
  NAND2_X1 U10116 ( .A1(n7923), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7941) );
  XNOR2_X1 U10117 ( .A(n7941), .B(P1_IR_REG_16__SCAN_IN), .ZN(n11561) );
  AOI22_X1 U10118 ( .A1(n8000), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n7999), 
        .B2(n11561), .ZN(n7942) );
  INV_X1 U10119 ( .A(n7944), .ZN(n7965) );
  INV_X1 U10120 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n7945) );
  NAND2_X1 U10121 ( .A1(n7946), .A2(n7945), .ZN(n7947) );
  AND2_X1 U10122 ( .A1(n7965), .A2(n7947), .ZN(n13836) );
  NAND2_X1 U10123 ( .A1(n7760), .A2(n13836), .ZN(n7954) );
  INV_X1 U10124 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n7948) );
  OR2_X1 U10125 ( .A1(n8385), .A2(n7948), .ZN(n7953) );
  INV_X1 U10126 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n7949) );
  OR2_X1 U10127 ( .A1(n8384), .A2(n7949), .ZN(n7952) );
  INV_X1 U10128 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n7950) );
  OR2_X1 U10129 ( .A1(n8115), .A2(n7950), .ZN(n7951) );
  NAND4_X1 U10130 ( .A1(n7954), .A2(n7953), .A3(n7952), .A4(n7951), .ZN(n13926) );
  INV_X1 U10131 ( .A(n13926), .ZN(n14277) );
  XNOR2_X1 U10132 ( .A(n11898), .B(n14277), .ZN(n11753) );
  OR2_X1 U10133 ( .A1(n11898), .A2(n13926), .ZN(n7955) );
  XNOR2_X1 U10134 ( .A(n7956), .B(SI_17_), .ZN(n7957) );
  XNOR2_X1 U10135 ( .A(n7958), .B(n7957), .ZN(n10456) );
  NAND2_X1 U10136 ( .A1(n10456), .A2(n8418), .ZN(n7963) );
  INV_X1 U10137 ( .A(n7971), .ZN(n7960) );
  NAND2_X1 U10138 ( .A1(n7960), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7961) );
  XNOR2_X1 U10139 ( .A(n7961), .B(P1_IR_REG_17__SCAN_IN), .ZN(n14039) );
  AOI22_X1 U10140 ( .A1(n6553), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n7999), 
        .B2(n14039), .ZN(n7962) );
  INV_X1 U10141 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n7964) );
  NAND2_X1 U10142 ( .A1(n7965), .A2(n7964), .ZN(n7966) );
  NAND2_X1 U10143 ( .A1(n8004), .A2(n7966), .ZN(n14268) );
  NOR2_X1 U10144 ( .A1(n14268), .A2(n8134), .ZN(n7969) );
  INV_X1 U10145 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n15262) );
  INV_X1 U10146 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n15434) );
  OAI22_X1 U10147 ( .A1(n8385), .A2(n15262), .B1(n8384), .B2(n15434), .ZN(
        n7968) );
  INV_X1 U10148 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n15280) );
  NOR2_X1 U10149 ( .A1(n8115), .A2(n15280), .ZN(n7967) );
  NOR2_X1 U10150 ( .A1(n14358), .A2(n13925), .ZN(n8336) );
  NAND2_X1 U10151 ( .A1(n14358), .A2(n13925), .ZN(n8325) );
  XNOR2_X1 U10152 ( .A(n7986), .B(SI_18_), .ZN(n7983) );
  XNOR2_X1 U10153 ( .A(n7983), .B(n7984), .ZN(n10830) );
  NAND2_X1 U10154 ( .A1(n10830), .A2(n8418), .ZN(n7974) );
  INV_X1 U10155 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n7970) );
  NAND2_X1 U10156 ( .A1(n7993), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7972) );
  XNOR2_X1 U10157 ( .A(n7972), .B(P1_IR_REG_18__SCAN_IN), .ZN(n14052) );
  AOI22_X1 U10158 ( .A1(n6553), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n7999), 
        .B2(n14052), .ZN(n7973) );
  XNOR2_X1 U10159 ( .A(n8004), .B(P1_REG3_REG_18__SCAN_IN), .ZN(n14253) );
  NAND2_X1 U10160 ( .A1(n14253), .A2(n7760), .ZN(n7979) );
  INV_X1 U10161 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n15416) );
  NAND2_X1 U10162 ( .A1(n7697), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n7976) );
  INV_X1 U10163 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n14355) );
  OR2_X1 U10164 ( .A1(n8115), .A2(n14355), .ZN(n7975) );
  OAI211_X1 U10165 ( .C1(n8385), .C2(n15416), .A(n7976), .B(n7975), .ZN(n7977)
         );
  INV_X1 U10166 ( .A(n7977), .ZN(n7978) );
  NAND2_X1 U10167 ( .A1(n7979), .A2(n7978), .ZN(n13924) );
  OR2_X1 U10168 ( .A1(n14350), .A2(n13924), .ZN(n7980) );
  NAND2_X1 U10169 ( .A1(n14242), .A2(n7980), .ZN(n7982) );
  NAND2_X1 U10170 ( .A1(n14350), .A2(n13924), .ZN(n7981) );
  NAND2_X1 U10171 ( .A1(n7982), .A2(n7981), .ZN(n14222) );
  INV_X1 U10172 ( .A(n7983), .ZN(n7985) );
  NAND2_X1 U10173 ( .A1(n7985), .A2(n7984), .ZN(n7988) );
  NAND2_X1 U10174 ( .A1(n7986), .A2(SI_18_), .ZN(n7987) );
  NAND2_X1 U10175 ( .A1(n7988), .A2(n7987), .ZN(n7992) );
  NAND2_X1 U10176 ( .A1(n7990), .A2(n7989), .ZN(n7991) );
  NAND2_X1 U10177 ( .A1(n10991), .A2(n8418), .ZN(n8002) );
  INV_X1 U10178 ( .A(n7997), .ZN(n7994) );
  NAND2_X1 U10179 ( .A1(n7994), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7995) );
  MUX2_X1 U10180 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7995), .S(
        P1_IR_REG_19__SCAN_IN), .Z(n7998) );
  INV_X1 U10181 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n7996) );
  NAND2_X1 U10182 ( .A1(n7997), .A2(n7996), .ZN(n8140) );
  NAND2_X1 U10183 ( .A1(n7998), .A2(n8140), .ZN(n14061) );
  AOI22_X1 U10184 ( .A1(n8000), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n7373), 
        .B2(n7999), .ZN(n8001) );
  INV_X1 U10185 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n8008) );
  INV_X1 U10186 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n13892) );
  INV_X1 U10187 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n8003) );
  OAI21_X1 U10188 ( .B1(n8004), .B2(n13892), .A(n8003), .ZN(n8005) );
  NAND2_X1 U10189 ( .A1(n8005), .A2(n8016), .ZN(n14228) );
  OR2_X1 U10190 ( .A1(n14228), .A2(n8134), .ZN(n8007) );
  AOI22_X1 U10191 ( .A1(n8133), .A2(P1_REG0_REG_19__SCAN_IN), .B1(n7697), .B2(
        P1_REG2_REG_19__SCAN_IN), .ZN(n8006) );
  OAI211_X1 U10192 ( .C1(n8115), .C2(n8008), .A(n8007), .B(n8006), .ZN(n14248)
         );
  INV_X1 U10193 ( .A(n14248), .ZN(n8009) );
  OR2_X1 U10194 ( .A1(n14345), .A2(n8009), .ZN(n8341) );
  NAND2_X1 U10195 ( .A1(n14345), .A2(n8009), .ZN(n8342) );
  OR2_X1 U10196 ( .A1(n14345), .A2(n14248), .ZN(n8011) );
  XNOR2_X1 U10197 ( .A(n8024), .B(SI_20_), .ZN(n8023) );
  XNOR2_X1 U10198 ( .A(n8023), .B(n8012), .ZN(n11033) );
  NAND2_X1 U10199 ( .A1(n11033), .A2(n8418), .ZN(n8014) );
  OR2_X1 U10200 ( .A1(n8419), .A2(n15251), .ZN(n8013) );
  INV_X1 U10201 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n8020) );
  INV_X1 U10202 ( .A(n8015), .ZN(n8033) );
  NAND2_X1 U10203 ( .A1(n8016), .A2(n13859), .ZN(n8017) );
  NAND2_X1 U10204 ( .A1(n8033), .A2(n8017), .ZN(n14212) );
  OR2_X1 U10205 ( .A1(n14212), .A2(n8134), .ZN(n8019) );
  AOI22_X1 U10206 ( .A1(n8133), .A2(P1_REG0_REG_20__SCAN_IN), .B1(n7697), .B2(
        P1_REG2_REG_20__SCAN_IN), .ZN(n8018) );
  OAI211_X1 U10207 ( .C1(n8115), .C2(n8020), .A(n8019), .B(n8018), .ZN(n13923)
         );
  XNOR2_X1 U10208 ( .A(n14415), .B(n13923), .ZN(n14203) );
  NAND2_X1 U10209 ( .A1(n14415), .A2(n13923), .ZN(n8021) );
  NAND2_X1 U10210 ( .A1(n8023), .A2(n8022), .ZN(n8026) );
  OR2_X1 U10211 ( .A1(n8024), .A2(n10802), .ZN(n8025) );
  NAND2_X1 U10212 ( .A1(n8026), .A2(n8025), .ZN(n8029) );
  XNOR2_X1 U10213 ( .A(n8027), .B(SI_21_), .ZN(n8028) );
  NAND2_X1 U10214 ( .A1(n11134), .A2(n8418), .ZN(n8031) );
  OR2_X1 U10215 ( .A1(n8419), .A2(n8900), .ZN(n8030) );
  INV_X1 U10216 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n8032) );
  NAND2_X1 U10217 ( .A1(n8033), .A2(n8032), .ZN(n8034) );
  NAND2_X1 U10218 ( .A1(n8044), .A2(n8034), .ZN(n14197) );
  OR2_X1 U10219 ( .A1(n14197), .A2(n8134), .ZN(n8039) );
  INV_X1 U10220 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n15436) );
  NAND2_X1 U10221 ( .A1(n7697), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n8036) );
  NAND2_X1 U10222 ( .A1(n8133), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n8035) );
  OAI211_X1 U10223 ( .C1(n15436), .C2(n8115), .A(n8036), .B(n8035), .ZN(n8037)
         );
  INV_X1 U10224 ( .A(n8037), .ZN(n8038) );
  NAND2_X1 U10225 ( .A1(n8039), .A2(n8038), .ZN(n13922) );
  INV_X1 U10226 ( .A(n13922), .ZN(n8189) );
  XNOR2_X1 U10227 ( .A(n14199), .B(n8189), .ZN(n14190) );
  INV_X1 U10228 ( .A(n14190), .ZN(n14187) );
  OR2_X1 U10229 ( .A1(n14199), .A2(n13922), .ZN(n8040) );
  OR2_X1 U10230 ( .A1(n8042), .A2(n8538), .ZN(n8043) );
  NAND2_X1 U10231 ( .A1(n8044), .A2(n13869), .ZN(n8045) );
  NAND2_X1 U10232 ( .A1(n8055), .A2(n8045), .ZN(n14178) );
  OR2_X1 U10233 ( .A1(n14178), .A2(n8134), .ZN(n8050) );
  INV_X1 U10234 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n14408) );
  NAND2_X1 U10235 ( .A1(n7697), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n8047) );
  NAND2_X1 U10236 ( .A1(n8069), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n8046) );
  OAI211_X1 U10237 ( .C1(n14408), .C2(n8385), .A(n8047), .B(n8046), .ZN(n8048)
         );
  INV_X1 U10238 ( .A(n8048), .ZN(n8049) );
  INV_X1 U10239 ( .A(n13817), .ZN(n13921) );
  XNOR2_X1 U10240 ( .A(n14410), .B(n13921), .ZN(n14174) );
  NAND2_X1 U10241 ( .A1(n14410), .A2(n13817), .ZN(n8051) );
  XNOR2_X1 U10242 ( .A(n8052), .B(SI_23_), .ZN(n11480) );
  NAND2_X1 U10243 ( .A1(n11480), .A2(n8418), .ZN(n8054) );
  INV_X1 U10244 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n11479) );
  OR2_X1 U10245 ( .A1(n8419), .A2(n11479), .ZN(n8053) );
  AND2_X1 U10246 ( .A1(n8055), .A2(n13792), .ZN(n8056) );
  OR2_X1 U10247 ( .A1(n8066), .A2(n8056), .ZN(n14165) );
  INV_X1 U10248 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n14164) );
  NAND2_X1 U10249 ( .A1(n8069), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n8058) );
  NAND2_X1 U10250 ( .A1(n8133), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n8057) );
  OAI211_X1 U10251 ( .C1(n8384), .C2(n14164), .A(n8058), .B(n8057), .ZN(n8059)
         );
  INV_X1 U10252 ( .A(n8059), .ZN(n8060) );
  OAI21_X1 U10253 ( .B1(n14165), .B2(n8134), .A(n8060), .ZN(n14140) );
  XNOR2_X1 U10254 ( .A(n14160), .B(n14140), .ZN(n14158) );
  INV_X1 U10255 ( .A(n14158), .ZN(n8061) );
  INV_X1 U10256 ( .A(n14138), .ZN(n8076) );
  XNOR2_X1 U10257 ( .A(n8063), .B(n8062), .ZN(n11613) );
  NAND2_X1 U10258 ( .A1(n11613), .A2(n8418), .ZN(n8065) );
  INV_X1 U10259 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n11617) );
  OR2_X1 U10260 ( .A1(n8419), .A2(n11617), .ZN(n8064) );
  OR2_X1 U10261 ( .A1(n8066), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n8068) );
  NAND2_X1 U10262 ( .A1(n8068), .A2(n8067), .ZN(n14149) );
  OR2_X1 U10263 ( .A1(n14149), .A2(n8134), .ZN(n8074) );
  INV_X1 U10264 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n14403) );
  NAND2_X1 U10265 ( .A1(n8069), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n8071) );
  NAND2_X1 U10266 ( .A1(n7697), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n8070) );
  OAI211_X1 U10267 ( .C1(n8385), .C2(n14403), .A(n8071), .B(n8070), .ZN(n8072)
         );
  INV_X1 U10268 ( .A(n8072), .ZN(n8073) );
  NAND2_X1 U10269 ( .A1(n8074), .A2(n8073), .ZN(n13920) );
  XNOR2_X1 U10270 ( .A(n14148), .B(n13920), .ZN(n14142) );
  NAND2_X1 U10271 ( .A1(n8076), .A2(n8075), .ZN(n14136) );
  OR2_X1 U10272 ( .A1(n14148), .A2(n13920), .ZN(n8077) );
  AND2_X2 U10273 ( .A1(n14136), .A2(n8077), .ZN(n14124) );
  XNOR2_X1 U10274 ( .A(n8079), .B(n8078), .ZN(n11649) );
  NAND2_X1 U10275 ( .A1(n11649), .A2(n8418), .ZN(n8081) );
  OR2_X1 U10276 ( .A1(n8419), .A2(n8965), .ZN(n8080) );
  NAND2_X1 U10277 ( .A1(n7697), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n8087) );
  INV_X1 U10278 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n15473) );
  OR2_X1 U10279 ( .A1(n8385), .A2(n15473), .ZN(n8086) );
  OAI21_X1 U10280 ( .B1(P1_REG3_REG_25__SCAN_IN), .B2(n8082), .A(n8097), .ZN(
        n14126) );
  OR2_X1 U10281 ( .A1(n8134), .A2(n14126), .ZN(n8085) );
  INV_X1 U10282 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n8083) );
  OR2_X1 U10283 ( .A1(n8115), .A2(n8083), .ZN(n8084) );
  NAND4_X1 U10284 ( .A1(n8087), .A2(n8086), .A3(n8085), .A4(n8084), .ZN(n14139) );
  INV_X1 U10285 ( .A(n14139), .ZN(n8088) );
  NAND2_X1 U10286 ( .A1(n14400), .A2(n8088), .ZN(n8197) );
  OR2_X1 U10287 ( .A1(n14400), .A2(n8088), .ZN(n8089) );
  NAND2_X1 U10288 ( .A1(n14400), .A2(n14139), .ZN(n8090) );
  XNOR2_X1 U10289 ( .A(n8091), .B(SI_26_), .ZN(n8092) );
  OR2_X1 U10290 ( .A1(n8419), .A2(n11821), .ZN(n8094) );
  NAND2_X1 U10291 ( .A1(n8133), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n8103) );
  INV_X1 U10292 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n14113) );
  OR2_X1 U10293 ( .A1(n8384), .A2(n14113), .ZN(n8102) );
  INV_X1 U10294 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n8096) );
  NAND2_X1 U10295 ( .A1(n8097), .A2(n8096), .ZN(n8098) );
  NAND2_X1 U10296 ( .A1(n8117), .A2(n8098), .ZN(n14112) );
  OR2_X1 U10297 ( .A1(n8134), .A2(n14112), .ZN(n8101) );
  INV_X1 U10298 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n8099) );
  OR2_X1 U10299 ( .A1(n8115), .A2(n8099), .ZN(n8100) );
  NAND4_X1 U10300 ( .A1(n8103), .A2(n8102), .A3(n8101), .A4(n8100), .ZN(n13919) );
  INV_X1 U10301 ( .A(n13919), .ZN(n8104) );
  NAND2_X1 U10302 ( .A1(n14396), .A2(n8104), .ZN(n8479) );
  OR2_X1 U10303 ( .A1(n14396), .A2(n8104), .ZN(n8105) );
  NAND2_X1 U10304 ( .A1(n14101), .A2(n14100), .ZN(n8107) );
  NAND2_X1 U10305 ( .A1(n14396), .A2(n13919), .ZN(n8106) );
  INV_X1 U10306 ( .A(n8108), .ZN(n8109) );
  XNOR2_X1 U10307 ( .A(n8109), .B(SI_27_), .ZN(n8110) );
  INV_X1 U10308 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n11873) );
  OR2_X1 U10309 ( .A1(n8419), .A2(n11873), .ZN(n8112) );
  NAND2_X1 U10310 ( .A1(n7697), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n8124) );
  INV_X1 U10311 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n8114) );
  OR2_X1 U10312 ( .A1(n8115), .A2(n8114), .ZN(n8123) );
  INV_X1 U10313 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n8116) );
  NAND2_X1 U10314 ( .A1(n8117), .A2(n8116), .ZN(n8118) );
  NAND2_X1 U10315 ( .A1(n8119), .A2(n8118), .ZN(n14092) );
  OR2_X1 U10316 ( .A1(n8134), .A2(n14092), .ZN(n8122) );
  INV_X1 U10317 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n8120) );
  OR2_X1 U10318 ( .A1(n8385), .A2(n8120), .ZN(n8121) );
  NAND4_X1 U10319 ( .A1(n8124), .A2(n8123), .A3(n8122), .A4(n8121), .ZN(n14106) );
  INV_X1 U10320 ( .A(n14106), .ZN(n8125) );
  NAND2_X1 U10321 ( .A1(n14095), .A2(n8125), .ZN(n8198) );
  OR2_X1 U10322 ( .A1(n14095), .A2(n8125), .ZN(n8126) );
  NAND2_X1 U10323 ( .A1(n8198), .A2(n8126), .ZN(n8448) );
  NAND2_X1 U10324 ( .A1(n14085), .A2(n8128), .ZN(n8199) );
  OAI21_X1 U10325 ( .B1(n9620), .B2(n8128), .A(n8493), .ZN(n8139) );
  INV_X1 U10326 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n14434) );
  INV_X1 U10327 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n15332) );
  MUX2_X1 U10328 ( .A(n14434), .B(n15332), .S(n8538), .Z(n8393) );
  XNOR2_X1 U10329 ( .A(n8393), .B(SI_29_), .ZN(n8390) );
  NAND2_X1 U10330 ( .A1(n13774), .A2(n8418), .ZN(n8132) );
  OR2_X1 U10331 ( .A1(n8419), .A2(n14434), .ZN(n8131) );
  NAND2_X1 U10332 ( .A1(n8133), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n8138) );
  NAND2_X1 U10333 ( .A1(n7697), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n8137) );
  OR2_X1 U10334 ( .A1(n8134), .A2(n12594), .ZN(n8136) );
  INV_X1 U10335 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n15333) );
  OR2_X1 U10336 ( .A1(n8115), .A2(n15333), .ZN(n8135) );
  NAND4_X1 U10337 ( .A1(n8138), .A2(n8137), .A3(n8136), .A4(n8135), .ZN(n13917) );
  XNOR2_X1 U10338 ( .A(n8139), .B(n8451), .ZN(n12603) );
  INV_X1 U10339 ( .A(n8140), .ZN(n8142) );
  INV_X1 U10340 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n8141) );
  NAND2_X1 U10341 ( .A1(n8142), .A2(n8141), .ZN(n8146) );
  INV_X1 U10342 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n8143) );
  NAND2_X2 U10343 ( .A1(n8157), .A2(n6548), .ZN(n10036) );
  INV_X1 U10344 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n8147) );
  OR2_X1 U10345 ( .A1(n10036), .A2(n8152), .ZN(n8151) );
  NAND2_X1 U10346 ( .A1(n11149), .A2(n8151), .ZN(n14755) );
  INV_X1 U10347 ( .A(n14148), .ZN(n14405) );
  INV_X1 U10348 ( .A(n11599), .ZN(n11608) );
  NAND2_X1 U10349 ( .A1(n14760), .A2(n14792), .ZN(n14759) );
  INV_X1 U10350 ( .A(n10969), .ZN(n10973) );
  INV_X1 U10351 ( .A(n11164), .ZN(n10818) );
  NAND2_X1 U10352 ( .A1(n10815), .A2(n10818), .ZN(n11023) );
  OR2_X2 U10353 ( .A1(n11355), .A2(n11736), .ZN(n11635) );
  INV_X1 U10354 ( .A(n14358), .ZN(n14272) );
  OR2_X2 U10355 ( .A1(n14265), .A2(n14350), .ZN(n14238) );
  OR2_X2 U10356 ( .A1(n14238), .A2(n14345), .ZN(n14226) );
  INV_X1 U10357 ( .A(n14199), .ZN(n14329) );
  INV_X1 U10358 ( .A(n14410), .ZN(n8353) );
  INV_X1 U10359 ( .A(n8155), .ZN(n8153) );
  INV_X1 U10360 ( .A(n6549), .ZN(n8425) );
  AOI21_X1 U10361 ( .B1(n8379), .B2(n8495), .A(n14793), .ZN(n8154) );
  NAND2_X1 U10362 ( .A1(n6549), .A2(n14061), .ZN(n8213) );
  INV_X1 U10363 ( .A(n8213), .ZN(n8156) );
  OR2_X1 U10364 ( .A1(n8155), .A2(n8156), .ZN(n14798) );
  INV_X1 U10365 ( .A(n8158), .ZN(n13965) );
  NAND2_X1 U10366 ( .A1(n14757), .A2(n13918), .ZN(n12597) );
  INV_X1 U10367 ( .A(P1_B_REG_SCAN_IN), .ZN(n8159) );
  OR2_X1 U10368 ( .A1(n13962), .A2(n8159), .ZN(n8160) );
  AND2_X1 U10369 ( .A1(n14247), .A2(n8160), .ZN(n14069) );
  INV_X1 U10370 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n15242) );
  OR2_X1 U10371 ( .A1(n8115), .A2(n15242), .ZN(n8163) );
  INV_X1 U10372 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n14076) );
  OR2_X1 U10373 ( .A1(n8384), .A2(n14076), .ZN(n8162) );
  INV_X1 U10374 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n15488) );
  OR2_X1 U10375 ( .A1(n8385), .A2(n15488), .ZN(n8161) );
  AND3_X1 U10376 ( .A1(n8163), .A2(n8162), .A3(n8161), .ZN(n8404) );
  INV_X1 U10377 ( .A(n8404), .ZN(n13916) );
  NAND2_X1 U10378 ( .A1(n14069), .A2(n13916), .ZN(n12595) );
  OAI211_X1 U10379 ( .C1(n7018), .C2(n14798), .A(n12597), .B(n12595), .ZN(
        n8164) );
  INV_X1 U10380 ( .A(n8164), .ZN(n8165) );
  INV_X1 U10381 ( .A(n8168), .ZN(n8429) );
  NAND2_X1 U10382 ( .A1(n14763), .A2(n14780), .ZN(n8430) );
  NAND2_X1 U10383 ( .A1(n10352), .A2(n13807), .ZN(n8169) );
  AND2_X1 U10384 ( .A1(n8430), .A2(n8169), .ZN(n8248) );
  INV_X1 U10385 ( .A(n8247), .ZN(n8170) );
  INV_X1 U10386 ( .A(n10300), .ZN(n10296) );
  NAND2_X1 U10387 ( .A1(n7733), .A2(n10379), .ZN(n8172) );
  INV_X1 U10388 ( .A(n8437), .ZN(n10287) );
  INV_X1 U10389 ( .A(n8435), .ZN(n10496) );
  INV_X1 U10390 ( .A(n13935), .ZN(n10961) );
  NAND2_X1 U10391 ( .A1(n10969), .A2(n10961), .ZN(n8175) );
  INV_X1 U10392 ( .A(n13934), .ZN(n11240) );
  OR2_X1 U10393 ( .A1(n11164), .A2(n11240), .ZN(n8176) );
  NAND2_X1 U10394 ( .A1(n10805), .A2(n8176), .ZN(n11018) );
  INV_X1 U10395 ( .A(n11021), .ZN(n8177) );
  NAND2_X1 U10396 ( .A1(n11232), .A2(n11230), .ZN(n8178) );
  INV_X1 U10397 ( .A(n11186), .ZN(n8179) );
  NAND2_X1 U10398 ( .A1(n11277), .A2(n7512), .ZN(n8181) );
  INV_X1 U10399 ( .A(n13931), .ZN(n11603) );
  OR2_X1 U10400 ( .A1(n11555), .A2(n11603), .ZN(n8180) );
  NAND2_X1 U10401 ( .A1(n8181), .A2(n8180), .ZN(n11459) );
  INV_X1 U10402 ( .A(n13930), .ZN(n11597) );
  OR2_X1 U10403 ( .A1(n11599), .A2(n11597), .ZN(n8182) );
  INV_X1 U10404 ( .A(n13929), .ZN(n14669) );
  NAND2_X1 U10405 ( .A1(n11676), .A2(n7936), .ZN(n8183) );
  NAND2_X1 U10406 ( .A1(n8183), .A2(n8319), .ZN(n11751) );
  NAND2_X1 U10407 ( .A1(n11898), .A2(n14277), .ZN(n8184) );
  INV_X1 U10408 ( .A(n8336), .ZN(n8185) );
  NAND2_X1 U10409 ( .A1(n8185), .A2(n8325), .ZN(n14262) );
  INV_X1 U10410 ( .A(n14262), .ZN(n14273) );
  INV_X1 U10411 ( .A(n13925), .ZN(n14250) );
  XNOR2_X1 U10412 ( .A(n14350), .B(n13924), .ZN(n14244) );
  NAND2_X1 U10413 ( .A1(n14240), .A2(n14244), .ZN(n8187) );
  INV_X1 U10414 ( .A(n13924), .ZN(n14275) );
  OR2_X1 U10415 ( .A1(n14350), .A2(n14275), .ZN(n8186) );
  INV_X1 U10416 ( .A(n14203), .ZN(n14205) );
  INV_X1 U10417 ( .A(n13923), .ZN(n13816) );
  OR2_X1 U10418 ( .A1(n14415), .A2(n13816), .ZN(n8188) );
  NAND2_X1 U10419 ( .A1(n14208), .A2(n8188), .ZN(n14189) );
  NAND2_X1 U10420 ( .A1(n14189), .A2(n14187), .ZN(n8191) );
  OR2_X1 U10421 ( .A1(n14199), .A2(n8189), .ZN(n8190) );
  OR2_X1 U10422 ( .A1(n14410), .A2(n13921), .ZN(n8192) );
  INV_X1 U10423 ( .A(n14140), .ZN(n8193) );
  NAND2_X1 U10424 ( .A1(n14160), .A2(n8193), .ZN(n8194) );
  INV_X1 U10425 ( .A(n13920), .ZN(n8195) );
  OR2_X1 U10426 ( .A1(n14148), .A2(n8195), .ZN(n8196) );
  NAND2_X1 U10427 ( .A1(n14141), .A2(n8196), .ZN(n14120) );
  NAND2_X1 U10428 ( .A1(n8476), .A2(n8198), .ZN(n8498) );
  NAND2_X1 U10429 ( .A1(n8498), .A2(n8499), .ZN(n8497) );
  OR2_X1 U10430 ( .A1(n12608), .A2(n6549), .ZN(n8244) );
  AND2_X1 U10431 ( .A1(n7971), .A2(n8201), .ZN(n8214) );
  NAND2_X1 U10432 ( .A1(n8214), .A2(n8216), .ZN(n8205) );
  NAND2_X1 U10433 ( .A1(n8203), .A2(n8202), .ZN(n8207) );
  NAND2_X1 U10434 ( .A1(n8207), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8204) );
  XNOR2_X1 U10435 ( .A(n8204), .B(P1_IR_REG_25__SCAN_IN), .ZN(n8221) );
  NAND2_X1 U10436 ( .A1(n8205), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8206) );
  NAND2_X1 U10437 ( .A1(n8208), .A2(n8207), .ZN(n8218) );
  NAND2_X1 U10438 ( .A1(n8209), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8211) );
  XNOR2_X1 U10439 ( .A(n8211), .B(n8210), .ZN(n11820) );
  NOR2_X1 U10440 ( .A1(n8218), .A2(n11820), .ZN(n8212) );
  NAND2_X1 U10441 ( .A1(n8221), .A2(n8212), .ZN(n10035) );
  INV_X1 U10442 ( .A(n10035), .ZN(n10039) );
  AOI21_X1 U10443 ( .B1(n10048), .B2(n8213), .A(n10039), .ZN(n10375) );
  INV_X1 U10444 ( .A(n8214), .ZN(n8215) );
  NAND2_X1 U10445 ( .A1(n8215), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8217) );
  XNOR2_X1 U10446 ( .A(n8217), .B(n8216), .ZN(n9914) );
  NAND2_X1 U10447 ( .A1(n10375), .A2(n9780), .ZN(n10051) );
  INV_X1 U10448 ( .A(n11820), .ZN(n8219) );
  OAI21_X1 U10449 ( .B1(n8218), .B2(P1_B_REG_SCAN_IN), .A(n8219), .ZN(n8220)
         );
  INV_X1 U10450 ( .A(n8220), .ZN(n8223) );
  INV_X1 U10451 ( .A(n8221), .ZN(n11652) );
  NAND3_X1 U10452 ( .A1(n11652), .A2(P1_B_REG_SCAN_IN), .A3(n8218), .ZN(n8222)
         );
  NOR4_X1 U10453 ( .A1(P1_D_REG_8__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_7__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n8231) );
  NOR4_X1 U10454 ( .A1(P1_D_REG_28__SCAN_IN), .A2(P1_D_REG_2__SCAN_IN), .A3(
        P1_D_REG_3__SCAN_IN), .A4(P1_D_REG_4__SCAN_IN), .ZN(n8230) );
  INV_X1 U10455 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n15240) );
  INV_X1 U10456 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n15356) );
  INV_X1 U10457 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n15389) );
  INV_X1 U10458 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n15418) );
  NAND4_X1 U10459 ( .A1(n15240), .A2(n15356), .A3(n15389), .A4(n15418), .ZN(
        n15468) );
  NOR4_X1 U10460 ( .A1(P1_D_REG_14__SCAN_IN), .A2(P1_D_REG_15__SCAN_IN), .A3(
        P1_D_REG_17__SCAN_IN), .A4(P1_D_REG_18__SCAN_IN), .ZN(n8227) );
  NOR4_X1 U10461 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n8226) );
  NOR4_X1 U10462 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_25__SCAN_IN), .A4(P1_D_REG_26__SCAN_IN), .ZN(n8225) );
  NOR4_X1 U10463 ( .A1(P1_D_REG_19__SCAN_IN), .A2(P1_D_REG_20__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n8224) );
  NAND4_X1 U10464 ( .A1(n8227), .A2(n8226), .A3(n8225), .A4(n8224), .ZN(n8228)
         );
  NOR4_X1 U10465 ( .A1(P1_D_REG_30__SCAN_IN), .A2(P1_D_REG_29__SCAN_IN), .A3(
        n15468), .A4(n8228), .ZN(n8229) );
  NAND3_X1 U10466 ( .A1(n8231), .A2(n8230), .A3(n8229), .ZN(n8232) );
  NAND2_X1 U10467 ( .A1(n9774), .A2(n8232), .ZN(n8238) );
  INV_X1 U10468 ( .A(n8238), .ZN(n8233) );
  INV_X1 U10469 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n9777) );
  AND2_X1 U10470 ( .A1(n8218), .A2(n11820), .ZN(n9776) );
  AOI21_X1 U10471 ( .B1(n9774), .B2(n9777), .A(n9776), .ZN(n8239) );
  NAND2_X1 U10472 ( .A1(n6549), .A2(n7373), .ZN(n14778) );
  OR2_X1 U10473 ( .A1(n8155), .A2(n14778), .ZN(n10056) );
  INV_X1 U10474 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n9781) );
  NAND2_X1 U10475 ( .A1(n9774), .A2(n9781), .ZN(n8234) );
  NAND2_X1 U10476 ( .A1(n11652), .A2(n11820), .ZN(n9778) );
  NAND2_X1 U10477 ( .A1(n8234), .A2(n9778), .ZN(n10510) );
  NAND2_X1 U10478 ( .A1(n10056), .A2(n10510), .ZN(n8240) );
  INV_X2 U10479 ( .A(n14804), .ZN(n14806) );
  NAND2_X1 U10480 ( .A1(n8241), .A2(n14806), .ZN(n8237) );
  INV_X1 U10481 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n8235) );
  NAND2_X1 U10482 ( .A1(n8237), .A2(n8236), .ZN(P1_U3525) );
  NAND2_X1 U10483 ( .A1(n8239), .A2(n8238), .ZN(n10045) );
  INV_X2 U10484 ( .A(n14809), .ZN(n14811) );
  NAND2_X1 U10485 ( .A1(n8152), .A2(n14061), .ZN(n8242) );
  AND2_X1 U10486 ( .A1(n8243), .A2(n8242), .ZN(n8245) );
  NAND2_X1 U10487 ( .A1(n8245), .A2(n12608), .ZN(n8405) );
  NAND2_X1 U10488 ( .A1(n8405), .A2(n8244), .ZN(n8389) );
  NAND2_X1 U10489 ( .A1(n8245), .A2(n8425), .ZN(n8246) );
  MUX2_X1 U10490 ( .A(n8248), .B(n8247), .S(n8340), .Z(n8251) );
  OR2_X1 U10491 ( .A1(n14763), .A2(n14780), .ZN(n8431) );
  INV_X1 U10492 ( .A(n10036), .ZN(n10034) );
  NAND2_X1 U10493 ( .A1(n8431), .A2(n10034), .ZN(n8249) );
  NAND3_X1 U10494 ( .A1(n8249), .A2(n8340), .A3(n8430), .ZN(n8250) );
  NAND2_X1 U10495 ( .A1(n8251), .A2(n8250), .ZN(n8255) );
  MUX2_X1 U10496 ( .A(n13808), .B(n13884), .S(n8340), .Z(n8256) );
  OAI21_X1 U10497 ( .B1(n10519), .B2(n14771), .A(n8256), .ZN(n8254) );
  MUX2_X1 U10498 ( .A(n14792), .B(n10352), .S(n8340), .Z(n8252) );
  NAND2_X1 U10499 ( .A1(n8252), .A2(n10178), .ZN(n8253) );
  INV_X1 U10500 ( .A(n8256), .ZN(n8258) );
  MUX2_X1 U10501 ( .A(n13885), .B(n10379), .S(n8340), .Z(n8259) );
  OAI21_X1 U10502 ( .B1(n7734), .B2(n7733), .A(n8259), .ZN(n8260) );
  NAND2_X1 U10503 ( .A1(n8261), .A2(n8260), .ZN(n8264) );
  MUX2_X1 U10504 ( .A(n10642), .B(n10493), .S(n8340), .Z(n8263) );
  MUX2_X1 U10505 ( .A(n13938), .B(n10631), .S(n8340), .Z(n8262) );
  NAND2_X1 U10506 ( .A1(n8264), .A2(n8263), .ZN(n8265) );
  NAND2_X1 U10507 ( .A1(n8266), .A2(n8265), .ZN(n8268) );
  MUX2_X1 U10508 ( .A(n13937), .B(n10744), .S(n8340), .Z(n8269) );
  MUX2_X1 U10509 ( .A(n10744), .B(n13937), .S(n8340), .Z(n8267) );
  MUX2_X1 U10510 ( .A(n10767), .B(n13936), .S(n8403), .Z(n8273) );
  MUX2_X1 U10511 ( .A(n13936), .B(n10767), .S(n8403), .Z(n8270) );
  NAND2_X1 U10512 ( .A1(n8271), .A2(n8270), .ZN(n8281) );
  INV_X1 U10513 ( .A(n8272), .ZN(n8275) );
  INV_X1 U10514 ( .A(n8273), .ZN(n8274) );
  NAND2_X1 U10515 ( .A1(n8281), .A2(n8280), .ZN(n8276) );
  MUX2_X1 U10516 ( .A(n13935), .B(n10969), .S(n8403), .Z(n8278) );
  MUX2_X1 U10517 ( .A(n10969), .B(n13935), .S(n8403), .Z(n8277) );
  INV_X1 U10518 ( .A(n8278), .ZN(n8279) );
  INV_X1 U10519 ( .A(n8340), .ZN(n8367) );
  MUX2_X1 U10520 ( .A(n13934), .B(n11164), .S(n8367), .Z(n8283) );
  MUX2_X1 U10521 ( .A(n13934), .B(n11164), .S(n8403), .Z(n8282) );
  MUX2_X1 U10522 ( .A(n13933), .B(n11232), .S(n8340), .Z(n8287) );
  NAND2_X1 U10523 ( .A1(n8286), .A2(n8287), .ZN(n8285) );
  MUX2_X1 U10524 ( .A(n13933), .B(n11232), .S(n8367), .Z(n8284) );
  NAND2_X1 U10525 ( .A1(n8285), .A2(n8284), .ZN(n8291) );
  INV_X1 U10526 ( .A(n8286), .ZN(n8289) );
  INV_X1 U10527 ( .A(n8287), .ZN(n8288) );
  NAND2_X1 U10528 ( .A1(n8289), .A2(n8288), .ZN(n8290) );
  NAND2_X1 U10529 ( .A1(n8291), .A2(n8290), .ZN(n8294) );
  MUX2_X1 U10530 ( .A(n13932), .B(n11373), .S(n8367), .Z(n8293) );
  MUX2_X1 U10531 ( .A(n13932), .B(n11373), .S(n8403), .Z(n8292) );
  MUX2_X1 U10532 ( .A(n13931), .B(n11555), .S(n8403), .Z(n8297) );
  MUX2_X1 U10533 ( .A(n13931), .B(n11555), .S(n8376), .Z(n8295) );
  INV_X1 U10534 ( .A(n8297), .ZN(n8298) );
  MUX2_X1 U10535 ( .A(n13930), .B(n11599), .S(n8367), .Z(n8301) );
  MUX2_X1 U10536 ( .A(n13930), .B(n11599), .S(n8340), .Z(n8299) );
  NAND2_X1 U10537 ( .A1(n8300), .A2(n8299), .ZN(n8307) );
  NAND2_X1 U10538 ( .A1(n6613), .A2(n7057), .ZN(n8306) );
  MUX2_X1 U10539 ( .A(n13929), .B(n11736), .S(n8376), .Z(n8311) );
  NOR2_X1 U10540 ( .A1(n8403), .A2(n13929), .ZN(n8303) );
  NOR2_X1 U10541 ( .A1(n11736), .A2(n8367), .ZN(n8302) );
  OR3_X1 U10542 ( .A1(n8311), .A2(n8303), .A3(n8302), .ZN(n8304) );
  AND2_X1 U10543 ( .A1(n11633), .A2(n8304), .ZN(n8305) );
  NAND3_X1 U10544 ( .A1(n8307), .A2(n8306), .A3(n8305), .ZN(n8318) );
  NAND2_X1 U10545 ( .A1(n8320), .A2(n8308), .ZN(n8313) );
  NOR2_X1 U10546 ( .A1(n8340), .A2(n14669), .ZN(n8309) );
  AOI21_X1 U10547 ( .B1(n11736), .B2(n8340), .A(n8309), .ZN(n8310) );
  AND2_X1 U10548 ( .A1(n8311), .A2(n8310), .ZN(n8312) );
  AOI22_X1 U10549 ( .A1(n8313), .A2(n8376), .B1(n11633), .B2(n8312), .ZN(n8317) );
  NAND2_X1 U10550 ( .A1(n8319), .A2(n8314), .ZN(n8315) );
  NAND2_X1 U10551 ( .A1(n8315), .A2(n8403), .ZN(n8316) );
  NAND2_X1 U10552 ( .A1(n8318), .A2(n7545), .ZN(n8329) );
  MUX2_X1 U10553 ( .A(n13926), .B(n11898), .S(n8376), .Z(n8322) );
  AND2_X1 U10554 ( .A1(n8328), .A2(n8322), .ZN(n8321) );
  INV_X1 U10555 ( .A(n8322), .ZN(n8323) );
  MUX2_X1 U10556 ( .A(n13926), .B(n11898), .S(n8403), .Z(n8330) );
  OR2_X1 U10557 ( .A1(n8323), .A2(n8330), .ZN(n8324) );
  XNOR2_X1 U10558 ( .A(n14350), .B(n8376), .ZN(n8332) );
  XNOR2_X1 U10559 ( .A(n8340), .B(n13924), .ZN(n8335) );
  NAND2_X1 U10560 ( .A1(n8332), .A2(n8335), .ZN(n8327) );
  MUX2_X1 U10561 ( .A(n13925), .B(n14358), .S(n8376), .Z(n8337) );
  NAND2_X1 U10562 ( .A1(n8337), .A2(n8325), .ZN(n8326) );
  INV_X1 U10563 ( .A(n8330), .ZN(n8331) );
  INV_X1 U10564 ( .A(n8332), .ZN(n8334) );
  OAI21_X1 U10565 ( .B1(n8337), .B2(n8336), .A(n8335), .ZN(n8333) );
  NAND2_X1 U10566 ( .A1(n8334), .A2(n8333), .ZN(n8339) );
  OR3_X1 U10567 ( .A1(n8337), .A2(n8336), .A3(n8335), .ZN(n8338) );
  MUX2_X1 U10568 ( .A(n8342), .B(n8341), .S(n8340), .Z(n8343) );
  INV_X1 U10569 ( .A(n14415), .ZN(n14213) );
  MUX2_X1 U10570 ( .A(n13816), .B(n14213), .S(n8403), .Z(n8345) );
  MUX2_X1 U10571 ( .A(n13923), .B(n14415), .S(n8376), .Z(n8344) );
  NAND2_X1 U10572 ( .A1(n8346), .A2(n8345), .ZN(n8347) );
  NAND2_X1 U10573 ( .A1(n8348), .A2(n8347), .ZN(n8350) );
  MUX2_X1 U10574 ( .A(n13922), .B(n14199), .S(n8376), .Z(n8351) );
  MUX2_X1 U10575 ( .A(n13922), .B(n14199), .S(n8403), .Z(n8349) );
  INV_X1 U10576 ( .A(n8351), .ZN(n8352) );
  MUX2_X1 U10577 ( .A(n13921), .B(n8353), .S(n8403), .Z(n8355) );
  MUX2_X1 U10578 ( .A(n13817), .B(n14410), .S(n8376), .Z(n8354) );
  MUX2_X1 U10579 ( .A(n14140), .B(n14160), .S(n8376), .Z(n8358) );
  MUX2_X1 U10580 ( .A(n14140), .B(n14160), .S(n8403), .Z(n8357) );
  MUX2_X1 U10581 ( .A(n13920), .B(n14148), .S(n8340), .Z(n8362) );
  MUX2_X1 U10582 ( .A(n13920), .B(n14148), .S(n8376), .Z(n8361) );
  MUX2_X1 U10583 ( .A(n14139), .B(n14400), .S(n8376), .Z(n8365) );
  MUX2_X1 U10584 ( .A(n14139), .B(n14400), .S(n8403), .Z(n8363) );
  INV_X1 U10585 ( .A(n8365), .ZN(n8366) );
  MUX2_X1 U10586 ( .A(n13919), .B(n14396), .S(n8403), .Z(n8369) );
  MUX2_X1 U10587 ( .A(n13919), .B(n14396), .S(n8367), .Z(n8368) );
  INV_X1 U10588 ( .A(n8369), .ZN(n8370) );
  MUX2_X1 U10589 ( .A(n14106), .B(n14095), .S(n8376), .Z(n8373) );
  NAND2_X1 U10590 ( .A1(n8374), .A2(n8373), .ZN(n8372) );
  MUX2_X1 U10591 ( .A(n14106), .B(n14095), .S(n8403), .Z(n8371) );
  NAND2_X1 U10592 ( .A1(n8372), .A2(n8371), .ZN(n8375) );
  MUX2_X1 U10593 ( .A(n13918), .B(n14085), .S(n8403), .Z(n8378) );
  MUX2_X1 U10594 ( .A(n13918), .B(n14085), .S(n8376), .Z(n8377) );
  MUX2_X1 U10595 ( .A(n13917), .B(n8379), .S(n8376), .Z(n8382) );
  MUX2_X1 U10596 ( .A(n13917), .B(n8379), .S(n8340), .Z(n8380) );
  INV_X1 U10597 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n14289) );
  OR2_X1 U10598 ( .A1(n8115), .A2(n14289), .ZN(n8388) );
  INV_X1 U10599 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n8383) );
  OR2_X1 U10600 ( .A1(n8384), .A2(n8383), .ZN(n8387) );
  INV_X1 U10601 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n14388) );
  OR2_X1 U10602 ( .A1(n8385), .A2(n14388), .ZN(n8386) );
  AND3_X1 U10603 ( .A1(n8388), .A2(n8387), .A3(n8386), .ZN(n8428) );
  AOI21_X1 U10604 ( .B1(n8389), .B2(n8428), .A(n8404), .ZN(n8402) );
  INV_X1 U10605 ( .A(SI_29_), .ZN(n8392) );
  NAND2_X1 U10606 ( .A1(n8393), .A2(n8392), .ZN(n8394) );
  NAND2_X1 U10607 ( .A1(n8395), .A2(n8394), .ZN(n8398) );
  MUX2_X1 U10608 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n8538), .Z(n8396) );
  NAND2_X1 U10609 ( .A1(n8396), .A2(SI_30_), .ZN(n8412) );
  OAI21_X1 U10610 ( .B1(SI_30_), .B2(n8396), .A(n8412), .ZN(n8397) );
  NAND2_X1 U10611 ( .A1(n8398), .A2(n8397), .ZN(n8399) );
  INV_X1 U10612 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n14431) );
  OR2_X1 U10613 ( .A1(n8419), .A2(n14431), .ZN(n8400) );
  OR2_X1 U10614 ( .A1(n8403), .A2(n8428), .ZN(n8406) );
  AOI21_X1 U10615 ( .B1(n8406), .B2(n8405), .A(n8404), .ZN(n8407) );
  AOI21_X1 U10616 ( .B1(n14291), .B2(n8403), .A(n8407), .ZN(n8408) );
  NOR2_X1 U10617 ( .A1(n8409), .A2(n8408), .ZN(n8410) );
  MUX2_X1 U10618 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n8538), .Z(n8414) );
  XNOR2_X1 U10619 ( .A(n8414), .B(SI_31_), .ZN(n8415) );
  INV_X1 U10620 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n14430) );
  OR2_X1 U10621 ( .A1(n8419), .A2(n14430), .ZN(n8420) );
  NOR2_X1 U10622 ( .A1(n8454), .A2(n8376), .ZN(n8459) );
  INV_X1 U10623 ( .A(n8428), .ZN(n14068) );
  AND2_X1 U10624 ( .A1(n8152), .A2(n6549), .ZN(n8422) );
  OR2_X1 U10625 ( .A1(n10048), .A2(n8422), .ZN(n8424) );
  OR2_X1 U10626 ( .A1(n14778), .A2(n12608), .ZN(n8423) );
  NAND2_X1 U10627 ( .A1(n8424), .A2(n8423), .ZN(n8467) );
  NAND2_X1 U10628 ( .A1(n12608), .A2(n8425), .ZN(n8463) );
  NAND2_X1 U10629 ( .A1(n8467), .A2(n8463), .ZN(n8455) );
  NOR2_X1 U10630 ( .A1(n8457), .A2(n14068), .ZN(n8426) );
  INV_X1 U10631 ( .A(n8430), .ZN(n8433) );
  INV_X1 U10632 ( .A(n8431), .ZN(n8432) );
  NOR2_X1 U10633 ( .A1(n8433), .A2(n8432), .ZN(n14781) );
  NAND3_X1 U10634 ( .A1(n8429), .A2(n14781), .A3(n8434), .ZN(n8436) );
  NOR4_X1 U10635 ( .A1(n10300), .A2(n8437), .A3(n8436), .A4(n8435), .ZN(n8438)
         );
  NAND4_X1 U10636 ( .A1(n8439), .A2(n10543), .A3(n8438), .A4(n10594), .ZN(
        n8440) );
  NOR4_X1 U10637 ( .A1(n11279), .A2(n11186), .A3(n11021), .A4(n8440), .ZN(
        n8441) );
  NAND4_X1 U10638 ( .A1(n14262), .A2(n8441), .A3(n11351), .A4(n11464), .ZN(
        n8442) );
  NOR4_X1 U10639 ( .A1(n11753), .A2(n11675), .A3(n8442), .A4(n7911), .ZN(n8443) );
  NAND4_X1 U10640 ( .A1(n14223), .A2(n14203), .A3(n8443), .A4(n14244), .ZN(
        n8444) );
  NOR3_X1 U10641 ( .A1(n14174), .A2(n14190), .A3(n8444), .ZN(n8445) );
  NAND4_X1 U10642 ( .A1(n8446), .A2(n8445), .A3(n14142), .A4(n14158), .ZN(
        n8447) );
  NOR4_X1 U10643 ( .A1(n8449), .A2(n8448), .A3(n14100), .A4(n8447), .ZN(n8452)
         );
  XNOR2_X1 U10644 ( .A(n14291), .B(n13916), .ZN(n8450) );
  XNOR2_X1 U10645 ( .A(n8453), .B(n14061), .ZN(n8464) );
  NOR3_X1 U10646 ( .A1(n14390), .A2(n14068), .A3(n8455), .ZN(n8458) );
  NOR3_X1 U10647 ( .A1(n8457), .A2(n14068), .A3(n8467), .ZN(n8456) );
  AOI21_X1 U10648 ( .B1(n8458), .B2(n8457), .A(n8456), .ZN(n8462) );
  XOR2_X1 U10649 ( .A(n8467), .B(n8459), .Z(n8460) );
  NAND3_X1 U10650 ( .A1(n8460), .A2(n14390), .A3(n14068), .ZN(n8461) );
  OAI211_X1 U10651 ( .C1(n8464), .C2(n8463), .A(n8462), .B(n8461), .ZN(n8465)
         );
  OR2_X1 U10652 ( .A1(n9914), .A2(P1_U3086), .ZN(n11477) );
  INV_X1 U10653 ( .A(n11477), .ZN(n8469) );
  NOR3_X1 U10654 ( .A1(n10051), .A2(n14276), .A3(n13962), .ZN(n8471) );
  OAI21_X1 U10655 ( .B1(n14439), .B2(n11477), .A(P1_B_REG_SCAN_IN), .ZN(n8470)
         );
  OR2_X1 U10656 ( .A1(n8471), .A2(n8470), .ZN(n8472) );
  NAND2_X1 U10657 ( .A1(n8473), .A2(n8472), .ZN(P1_U3242) );
  INV_X1 U10658 ( .A(n14798), .ZN(n14372) );
  NAND2_X1 U10659 ( .A1(n14811), .A2(n14372), .ZN(n14327) );
  INV_X1 U10660 ( .A(n14327), .ZN(n14341) );
  NAND2_X1 U10661 ( .A1(n14095), .A2(n14341), .ZN(n8487) );
  AOI22_X1 U10662 ( .A1(n14247), .A2(n13918), .B1(n14757), .B2(n13919), .ZN(
        n8475) );
  OAI21_X1 U10663 ( .B1(n8476), .B2(n14761), .A(n8475), .ZN(n8477) );
  NAND3_X1 U10664 ( .A1(n14102), .A2(n8479), .A3(n14783), .ZN(n8480) );
  AOI21_X1 U10665 ( .B1(n14095), .B2(n14110), .A(n14793), .ZN(n8485) );
  NAND2_X1 U10666 ( .A1(n8485), .A2(n8494), .ZN(n14096) );
  NAND2_X1 U10667 ( .A1(n14099), .A2(n14096), .ZN(n8488) );
  NAND2_X1 U10668 ( .A1(n8487), .A2(n8486), .ZN(P1_U3555) );
  NAND2_X1 U10669 ( .A1(n14806), .A2(n14372), .ZN(n14411) );
  INV_X1 U10670 ( .A(n14411), .ZN(n14416) );
  NAND2_X1 U10671 ( .A1(n14095), .A2(n14416), .ZN(n8490) );
  NAND2_X1 U10672 ( .A1(n8490), .A2(n8489), .ZN(P1_U3523) );
  NAND2_X1 U10673 ( .A1(n8491), .A2(n8499), .ZN(n8492) );
  NAND2_X1 U10674 ( .A1(n8493), .A2(n8492), .ZN(n14081) );
  AOI21_X1 U10675 ( .B1(n14085), .B2(n8494), .A(n14793), .ZN(n8496) );
  NAND2_X1 U10676 ( .A1(n8496), .A2(n8495), .ZN(n14087) );
  OAI21_X1 U10677 ( .B1(n8499), .B2(n8498), .A(n8497), .ZN(n8500) );
  NAND2_X1 U10678 ( .A1(n8500), .A2(n14783), .ZN(n8502) );
  AOI22_X1 U10679 ( .A1(n14247), .A2(n13917), .B1(n14757), .B2(n14106), .ZN(
        n8501) );
  NAND2_X1 U10680 ( .A1(n8502), .A2(n8501), .ZN(n14080) );
  NOR2_X1 U10681 ( .A1(n8503), .A2(n14080), .ZN(n9619) );
  OR2_X1 U10682 ( .A1(n14806), .A2(n8504), .ZN(n8505) );
  NOR2_X1 U10683 ( .A1(P3_IR_REG_6__SCAN_IN), .A2(P3_IR_REG_5__SCAN_IN), .ZN(
        n8510) );
  AND4_X2 U10684 ( .A1(n8510), .A2(n8509), .A3(n8508), .A4(n15350), .ZN(n8512)
         );
  NOR2_X1 U10685 ( .A1(P3_IR_REG_20__SCAN_IN), .A2(P3_IR_REG_21__SCAN_IN), 
        .ZN(n8518) );
  NOR2_X1 U10686 ( .A1(P3_IR_REG_22__SCAN_IN), .A2(P3_IR_REG_19__SCAN_IN), 
        .ZN(n8517) );
  NOR2_X1 U10687 ( .A1(P3_IR_REG_18__SCAN_IN), .A2(P3_IR_REG_16__SCAN_IN), 
        .ZN(n8516) );
  NOR2_X1 U10688 ( .A1(P3_IR_REG_17__SCAN_IN), .A2(P3_IR_REG_15__SCAN_IN), 
        .ZN(n8515) );
  INV_X1 U10689 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n8521) );
  INV_X1 U10690 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n8522) );
  NAND2_X1 U10691 ( .A1(n8526), .A2(n8523), .ZN(n13196) );
  INV_X1 U10692 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n8524) );
  XNOR2_X2 U10693 ( .A(n8525), .B(P3_IR_REG_30__SCAN_IN), .ZN(n8530) );
  XNOR2_X2 U10694 ( .A(n8527), .B(n8523), .ZN(n8529) );
  AND2_X2 U10695 ( .A1(n12591), .A2(n8528), .ZN(n9032) );
  NAND2_X1 U10696 ( .A1(n9032), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n8534) );
  NAND2_X1 U10697 ( .A1(n8637), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n8533) );
  NAND2_X1 U10698 ( .A1(n8601), .A2(P3_REG0_REG_1__SCAN_IN), .ZN(n8532) );
  NAND2_X4 U10699 ( .A1(n8530), .A2(n8529), .ZN(n10796) );
  INV_X1 U10700 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n10219) );
  OR2_X1 U10701 ( .A1(n10796), .A2(n10219), .ZN(n8531) );
  INV_X1 U10702 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n8536) );
  NAND2_X1 U10703 ( .A1(n8537), .A2(n8535), .ZN(n9030) );
  AND2_X2 U10704 ( .A1(n8565), .A2(n8538), .ZN(n8594) );
  AND2_X2 U10705 ( .A1(n8565), .A2(n9769), .ZN(n9017) );
  XNOR2_X1 U10706 ( .A(n8559), .B(n8560), .ZN(n9765) );
  NAND2_X1 U10707 ( .A1(n9017), .A2(n9765), .ZN(n8541) );
  INV_X2 U10708 ( .A(n8565), .ZN(n8858) );
  NAND2_X1 U10709 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(n15507), .ZN(n8539) );
  NAND2_X1 U10710 ( .A1(n8858), .A2(n10345), .ZN(n8540) );
  NAND2_X1 U10711 ( .A1(n15121), .A2(n8551), .ZN(n12418) );
  NAND2_X1 U10712 ( .A1(n9032), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n8546) );
  NAND2_X1 U10713 ( .A1(n8637), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n8545) );
  NAND2_X1 U10714 ( .A1(n8601), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n8544) );
  OR2_X1 U10715 ( .A1(n10796), .A2(n15495), .ZN(n8543) );
  INV_X1 U10716 ( .A(n15507), .ZN(n8550) );
  NOR2_X1 U10717 ( .A1(n15479), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n8547) );
  NOR2_X1 U10718 ( .A1(n8560), .A2(n8547), .ZN(n8548) );
  NAND2_X1 U10719 ( .A1(n7602), .A2(SI_0_), .ZN(n9169) );
  OAI21_X1 U10720 ( .B1(n8538), .B2(n8548), .A(n9169), .ZN(n13219) );
  INV_X1 U10721 ( .A(n13219), .ZN(n8549) );
  MUX2_X1 U10722 ( .A(n8550), .B(n8549), .S(n10198), .Z(n10397) );
  INV_X1 U10723 ( .A(n10397), .ZN(n10155) );
  NAND2_X1 U10724 ( .A1(n15138), .A2(n10155), .ZN(n15141) );
  INV_X1 U10725 ( .A(n8551), .ZN(n8552) );
  OR2_X1 U10726 ( .A1(n15121), .A2(n8552), .ZN(n15123) );
  NAND2_X1 U10727 ( .A1(n15140), .A2(n15123), .ZN(n8568) );
  NAND2_X1 U10728 ( .A1(n9032), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n8556) );
  NAND2_X1 U10729 ( .A1(n8637), .A2(P3_REG3_REG_2__SCAN_IN), .ZN(n8555) );
  NAND2_X1 U10730 ( .A1(n8601), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n8554) );
  INV_X1 U10731 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n10859) );
  NAND4_X4 U10732 ( .A1(n8556), .A2(n8555), .A3(n8554), .A4(n8553), .ZN(n15137) );
  INV_X1 U10733 ( .A(n8586), .ZN(n8557) );
  XNOR2_X1 U10734 ( .A(n10028), .B(P2_DATAO_REG_2__SCAN_IN), .ZN(n8562) );
  XNOR2_X1 U10735 ( .A(n8576), .B(n8562), .ZN(n9793) );
  NAND2_X1 U10736 ( .A1(n9017), .A2(n9793), .ZN(n8564) );
  INV_X1 U10737 ( .A(SI_2_), .ZN(n15292) );
  NAND2_X1 U10738 ( .A1(n8594), .A2(n15292), .ZN(n8563) );
  OAI211_X1 U10739 ( .C1(n10892), .C2(n8565), .A(n8564), .B(n8563), .ZN(n15117) );
  NAND2_X1 U10740 ( .A1(n15137), .A2(n15117), .ZN(n12426) );
  NAND2_X1 U10741 ( .A1(n8567), .A2(n8566), .ZN(n12427) );
  AND2_X1 U10742 ( .A1(n12426), .A2(n12427), .ZN(n15124) );
  INV_X1 U10743 ( .A(n15124), .ZN(n15115) );
  OR2_X1 U10744 ( .A1(n15137), .A2(n8566), .ZN(n8569) );
  NAND2_X1 U10745 ( .A1(n9032), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n8573) );
  INV_X1 U10746 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n15459) );
  NAND2_X1 U10747 ( .A1(n8637), .A2(n15459), .ZN(n8572) );
  NAND2_X1 U10748 ( .A1(n8861), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n8571) );
  INV_X1 U10749 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n10869) );
  OR2_X1 U10750 ( .A1(n10796), .A2(n10869), .ZN(n8570) );
  NAND2_X1 U10751 ( .A1(n6980), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8574) );
  XNOR2_X1 U10752 ( .A(n8574), .B(P3_IR_REG_3__SCAN_IN), .ZN(n10893) );
  XNOR2_X1 U10753 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .ZN(n8577) );
  XNOR2_X1 U10754 ( .A(n8589), .B(n8577), .ZN(n9786) );
  NAND2_X1 U10755 ( .A1(n9017), .A2(n9786), .ZN(n8579) );
  INV_X1 U10756 ( .A(SI_3_), .ZN(n9787) );
  OAI211_X1 U10757 ( .C1(n10893), .C2(n10198), .A(n8579), .B(n8578), .ZN(
        n15161) );
  OR2_X1 U10758 ( .A1(n15120), .A2(n15161), .ZN(n12431) );
  NAND2_X1 U10759 ( .A1(n15120), .A2(n15161), .ZN(n12430) );
  AND2_X2 U10760 ( .A1(n12431), .A2(n12430), .ZN(n12385) );
  INV_X1 U10761 ( .A(n15161), .ZN(n10484) );
  NAND2_X1 U10762 ( .A1(n15120), .A2(n10484), .ZN(n8580) );
  NAND2_X1 U10763 ( .A1(n9032), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n8585) );
  AND2_X1 U10764 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n8581) );
  OR2_X1 U10765 ( .A1(n8581), .A2(n8599), .ZN(n10734) );
  NAND2_X1 U10766 ( .A1(n8988), .A2(n10734), .ZN(n8584) );
  NAND2_X1 U10767 ( .A1(n8861), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n8583) );
  INV_X1 U10768 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n10860) );
  OR2_X1 U10769 ( .A1(n10796), .A2(n10860), .ZN(n8582) );
  NAND4_X1 U10770 ( .A1(n8585), .A2(n8584), .A3(n8583), .A4(n8582), .ZN(n12744) );
  NOR2_X1 U10771 ( .A1(n6980), .A2(P3_IR_REG_3__SCAN_IN), .ZN(n8630) );
  INV_X1 U10772 ( .A(n8630), .ZN(n8587) );
  NAND2_X1 U10773 ( .A1(n8587), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8609) );
  XNOR2_X1 U10774 ( .A(n8609), .B(P3_IR_REG_4__SCAN_IN), .ZN(n10895) );
  NAND2_X1 U10775 ( .A1(n10032), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n8588) );
  NAND2_X1 U10776 ( .A1(n15480), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n8590) );
  NAND2_X1 U10777 ( .A1(n8612), .A2(n8590), .ZN(n8591) );
  NAND2_X1 U10778 ( .A1(n8592), .A2(n8591), .ZN(n8593) );
  NAND2_X1 U10779 ( .A1(n8613), .A2(n8593), .ZN(n9761) );
  NAND2_X1 U10780 ( .A1(n9017), .A2(n9761), .ZN(n8596) );
  INV_X1 U10782 ( .A(SI_4_), .ZN(n9762) );
  NAND2_X1 U10783 ( .A1(n12363), .A2(n9762), .ZN(n8595) );
  OAI211_X1 U10784 ( .C1(n10895), .C2(n10198), .A(n8596), .B(n8595), .ZN(
        n15168) );
  OR2_X1 U10785 ( .A1(n12744), .A2(n15168), .ZN(n12440) );
  NAND2_X1 U10786 ( .A1(n12744), .A2(n15168), .ZN(n12439) );
  NAND2_X1 U10787 ( .A1(n10728), .A2(n10727), .ZN(n8598) );
  INV_X1 U10788 ( .A(n15168), .ZN(n10735) );
  NAND2_X1 U10789 ( .A1(n12744), .A2(n10735), .ZN(n8597) );
  NAND2_X1 U10790 ( .A1(n8598), .A2(n8597), .ZN(n11070) );
  NAND2_X1 U10791 ( .A1(n9032), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n8607) );
  OR2_X1 U10792 ( .A1(n8599), .A2(n10836), .ZN(n8600) );
  NAND2_X1 U10793 ( .A1(n8620), .A2(n8600), .ZN(n11078) );
  NAND2_X1 U10794 ( .A1(n8988), .A2(n11078), .ZN(n8606) );
  NAND2_X1 U10795 ( .A1(n8861), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n8605) );
  INV_X1 U10796 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n8603) );
  OR2_X1 U10797 ( .A1(n10796), .A2(n8603), .ZN(n8604) );
  NAND4_X1 U10798 ( .A1(n8607), .A2(n8606), .A3(n8605), .A4(n8604), .ZN(n12743) );
  INV_X1 U10799 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n8608) );
  NAND2_X1 U10800 ( .A1(n8609), .A2(n8608), .ZN(n8610) );
  NAND2_X1 U10801 ( .A1(n8610), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8611) );
  XNOR2_X1 U10802 ( .A(n8611), .B(P3_IR_REG_5__SCAN_IN), .ZN(n10896) );
  NAND2_X1 U10803 ( .A1(n9795), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n8614) );
  OAI21_X1 U10804 ( .B1(n8616), .B2(n8615), .A(n8628), .ZN(n9788) );
  NAND2_X1 U10805 ( .A1(n12362), .A2(n9788), .ZN(n8618) );
  INV_X1 U10806 ( .A(SI_5_), .ZN(n9789) );
  NAND2_X1 U10807 ( .A1(n12363), .A2(n9789), .ZN(n8617) );
  OAI211_X1 U10808 ( .C1(n10896), .C2(n10198), .A(n8618), .B(n8617), .ZN(
        n15173) );
  OR2_X1 U10809 ( .A1(n12743), .A2(n15173), .ZN(n12446) );
  NAND2_X1 U10810 ( .A1(n12743), .A2(n15173), .ZN(n12436) );
  INV_X1 U10811 ( .A(n15173), .ZN(n11079) );
  OR2_X1 U10812 ( .A1(n12743), .A2(n11079), .ZN(n8619) );
  NAND2_X1 U10813 ( .A1(n9032), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n8626) );
  NAND2_X1 U10814 ( .A1(n8620), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8621) );
  NAND2_X1 U10815 ( .A1(n8638), .A2(n8621), .ZN(n12714) );
  NAND2_X1 U10816 ( .A1(n8988), .A2(n12714), .ZN(n8625) );
  NAND2_X1 U10817 ( .A1(n8861), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n8624) );
  INV_X1 U10818 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n8622) );
  OR2_X1 U10819 ( .A1(n10796), .A2(n8622), .ZN(n8623) );
  XNOR2_X1 U10820 ( .A(n8649), .B(n8648), .ZN(n9758) );
  NAND2_X1 U10821 ( .A1(n9017), .A2(n9758), .ZN(n8635) );
  NOR2_X1 U10822 ( .A1(P3_IR_REG_5__SCAN_IN), .A2(P3_IR_REG_4__SCAN_IN), .ZN(
        n8629) );
  NAND2_X1 U10823 ( .A1(n8630), .A2(n8629), .ZN(n8632) );
  NAND2_X1 U10824 ( .A1(n8632), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8631) );
  MUX2_X1 U10825 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8631), .S(
        P3_IR_REG_6__SCAN_IN), .Z(n8633) );
  NAND2_X1 U10826 ( .A1(n8858), .A2(n10899), .ZN(n8634) );
  NAND2_X1 U10827 ( .A1(n12742), .A2(n15178), .ZN(n12448) );
  INV_X1 U10828 ( .A(n15178), .ZN(n11065) );
  NAND2_X1 U10829 ( .A1(n9032), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n8644) );
  AND2_X1 U10830 ( .A1(n8638), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8639) );
  OR2_X1 U10831 ( .A1(n8639), .A2(n8658), .ZN(n11179) );
  NAND2_X1 U10832 ( .A1(n8988), .A2(n11179), .ZN(n8643) );
  NAND2_X1 U10833 ( .A1(n8601), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n8642) );
  INV_X1 U10834 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n8640) );
  OR2_X1 U10835 ( .A1(n10796), .A2(n8640), .ZN(n8641) );
  NAND4_X1 U10836 ( .A1(n8644), .A2(n8643), .A3(n8642), .A4(n8641), .ZN(n12741) );
  NAND2_X1 U10837 ( .A1(n8646), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8645) );
  MUX2_X1 U10838 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8645), .S(
        P3_IR_REG_7__SCAN_IN), .Z(n8647) );
  NAND2_X1 U10839 ( .A1(n8647), .A2(n8677), .ZN(n12338) );
  INV_X1 U10840 ( .A(n12338), .ZN(n10900) );
  NAND2_X1 U10841 ( .A1(n9798), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n8650) );
  NAND2_X1 U10842 ( .A1(n8666), .A2(n8650), .ZN(n8651) );
  NAND2_X1 U10843 ( .A1(n8652), .A2(n8651), .ZN(n8653) );
  NAND2_X1 U10844 ( .A1(n8667), .A2(n8653), .ZN(n9763) );
  NAND2_X1 U10845 ( .A1(n9017), .A2(n9763), .ZN(n8655) );
  INV_X1 U10846 ( .A(SI_7_), .ZN(n9764) );
  OAI211_X1 U10847 ( .C1(n10900), .C2(n10198), .A(n8655), .B(n8654), .ZN(
        n15183) );
  NAND2_X1 U10848 ( .A1(n12741), .A2(n15183), .ZN(n12453) );
  AND2_X2 U10849 ( .A1(n12454), .A2(n12453), .ZN(n12450) );
  INV_X1 U10850 ( .A(n15183), .ZN(n11180) );
  AND2_X1 U10851 ( .A1(n12741), .A2(n11180), .ZN(n8656) );
  NAND2_X1 U10852 ( .A1(n10792), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n8664) );
  INV_X1 U10853 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n8657) );
  NOR2_X1 U10854 ( .A1(n8658), .A2(n8657), .ZN(n8659) );
  OR2_X1 U10855 ( .A1(n8671), .A2(n8659), .ZN(n11294) );
  NAND2_X1 U10856 ( .A1(n8988), .A2(n11294), .ZN(n8663) );
  NAND2_X1 U10857 ( .A1(n8861), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n8662) );
  INV_X1 U10858 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n8660) );
  OR2_X1 U10859 ( .A1(n10796), .A2(n8660), .ZN(n8661) );
  NAND2_X1 U10860 ( .A1(n8677), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8665) );
  XNOR2_X1 U10861 ( .A(n8665), .B(P3_IR_REG_8__SCAN_IN), .ZN(n10903) );
  NAND2_X1 U10862 ( .A1(n12363), .A2(SI_8_), .ZN(n8670) );
  XNOR2_X1 U10863 ( .A(n9834), .B(P2_DATAO_REG_8__SCAN_IN), .ZN(n8668) );
  XNOR2_X1 U10864 ( .A(n6693), .B(n8668), .ZN(n9790) );
  NAND2_X1 U10865 ( .A1(n9017), .A2(n9790), .ZN(n8669) );
  OAI211_X1 U10866 ( .C1(n10198), .C2(n12324), .A(n8670), .B(n8669), .ZN(
        n12460) );
  XNOR2_X1 U10867 ( .A(n12740), .B(n12460), .ZN(n12389) );
  NAND2_X1 U10868 ( .A1(n9032), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n8676) );
  OR2_X1 U10869 ( .A1(n8671), .A2(n15461), .ZN(n8672) );
  NAND2_X1 U10870 ( .A1(n8688), .A2(n8672), .ZN(n11048) );
  NAND2_X1 U10871 ( .A1(n8988), .A2(n11048), .ZN(n8675) );
  NAND2_X1 U10872 ( .A1(n8861), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n8674) );
  INV_X1 U10873 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n15444) );
  OR2_X1 U10874 ( .A1(n10796), .A2(n15444), .ZN(n8673) );
  OAI21_X1 U10875 ( .B1(n8677), .B2(P3_IR_REG_8__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8679) );
  INV_X1 U10876 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n8678) );
  XNOR2_X1 U10877 ( .A(n8679), .B(n8678), .ZN(n15101) );
  INV_X1 U10878 ( .A(n15101), .ZN(n10883) );
  NAND2_X1 U10879 ( .A1(n9834), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n8680) );
  INV_X1 U10880 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n9833) );
  NAND2_X1 U10881 ( .A1(n9833), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n8682) );
  XNOR2_X1 U10882 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(P2_DATAO_REG_9__SCAN_IN), 
        .ZN(n8683) );
  XNOR2_X1 U10883 ( .A(n8695), .B(n8683), .ZN(n9782) );
  NAND2_X1 U10884 ( .A1(n9782), .A2(n12362), .ZN(n8685) );
  INV_X1 U10885 ( .A(SI_9_), .ZN(n9783) );
  NAND2_X1 U10886 ( .A1(n12363), .A2(n9783), .ZN(n8684) );
  OAI211_X1 U10887 ( .C1(n10883), .C2(n10198), .A(n8685), .B(n8684), .ZN(
        n15193) );
  INV_X1 U10888 ( .A(n15193), .ZN(n12414) );
  NAND2_X1 U10889 ( .A1(n12739), .A2(n12414), .ZN(n12471) );
  OR2_X1 U10890 ( .A1(n12739), .A2(n12414), .ZN(n8686) );
  OR2_X1 U10891 ( .A1(n12740), .A2(n12460), .ZN(n11340) );
  AND2_X1 U10892 ( .A1(n12465), .A2(n11340), .ZN(n8687) );
  NAND2_X1 U10893 ( .A1(n11341), .A2(n8687), .ZN(n11342) );
  NAND2_X1 U10894 ( .A1(n10792), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n8693) );
  NAND2_X1 U10895 ( .A1(n8688), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8689) );
  NAND2_X1 U10896 ( .A1(n8714), .A2(n8689), .ZN(n11452) );
  NAND2_X1 U10897 ( .A1(n8988), .A2(n11452), .ZN(n8692) );
  NAND2_X1 U10898 ( .A1(n8861), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n8691) );
  INV_X1 U10899 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n11454) );
  OR2_X1 U10900 ( .A1(n10796), .A2(n11454), .ZN(n8690) );
  NAND4_X1 U10901 ( .A1(n8693), .A2(n8692), .A3(n8691), .A4(n8690), .ZN(n12738) );
  INV_X1 U10902 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n9840) );
  INV_X1 U10903 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n9838) );
  NAND2_X1 U10904 ( .A1(n15281), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n8703) );
  INV_X1 U10905 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n9913) );
  NAND2_X1 U10906 ( .A1(n9913), .A2(P2_DATAO_REG_10__SCAN_IN), .ZN(n8696) );
  NAND2_X1 U10907 ( .A1(n8703), .A2(n8696), .ZN(n8704) );
  XNOR2_X1 U10908 ( .A(n8705), .B(n8704), .ZN(n9784) );
  NAND2_X1 U10909 ( .A1(n9784), .A2(n12362), .ZN(n8700) );
  NAND2_X1 U10910 ( .A1(n8697), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8698) );
  XNOR2_X1 U10911 ( .A(n8698), .B(n15498), .ZN(n11246) );
  AOI22_X1 U10912 ( .A1(n12370), .A2(n9785), .B1(n8858), .B2(n11246), .ZN(
        n8699) );
  NAND2_X1 U10913 ( .A1(n8700), .A2(n8699), .ZN(n15199) );
  OR2_X1 U10914 ( .A1(n12738), .A2(n15199), .ZN(n12413) );
  AND2_X1 U10915 ( .A1(n12738), .A2(n15199), .ZN(n12477) );
  INV_X1 U10916 ( .A(n12477), .ZN(n8701) );
  NAND2_X1 U10917 ( .A1(n12413), .A2(n8701), .ZN(n12469) );
  INV_X1 U10918 ( .A(n15199), .ZN(n11456) );
  NAND2_X1 U10919 ( .A1(n11456), .A2(n12738), .ZN(n8702) );
  XNOR2_X1 U10920 ( .A(n10069), .B(P2_DATAO_REG_11__SCAN_IN), .ZN(n8706) );
  XNOR2_X1 U10921 ( .A(n8723), .B(n8706), .ZN(n9803) );
  NAND2_X1 U10922 ( .A1(n9803), .A2(n12362), .ZN(n8713) );
  NOR2_X1 U10923 ( .A1(n8697), .A2(P3_IR_REG_10__SCAN_IN), .ZN(n8710) );
  NOR2_X1 U10924 ( .A1(n8710), .A2(n13195), .ZN(n8707) );
  MUX2_X1 U10925 ( .A(n13195), .B(n8707), .S(P3_IR_REG_11__SCAN_IN), .Z(n8708)
         );
  INV_X1 U10926 ( .A(n8708), .ZN(n8711) );
  NAND2_X1 U10927 ( .A1(n8710), .A2(n15342), .ZN(n8743) );
  AND2_X1 U10928 ( .A1(n8711), .A2(n8743), .ZN(n11484) );
  AOI22_X1 U10929 ( .A1(n12370), .A2(SI_11_), .B1(n8858), .B2(n11484), .ZN(
        n8712) );
  NAND2_X1 U10930 ( .A1(n8713), .A2(n8712), .ZN(n14637) );
  NAND2_X1 U10931 ( .A1(n9032), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n8719) );
  NAND2_X1 U10932 ( .A1(n8714), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8715) );
  NAND2_X1 U10933 ( .A1(n8730), .A2(n8715), .ZN(n11529) );
  NAND2_X1 U10934 ( .A1(n8988), .A2(n11529), .ZN(n8718) );
  NAND2_X1 U10935 ( .A1(n8861), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n8717) );
  INV_X1 U10936 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n11531) );
  NAND4_X1 U10937 ( .A1(n8719), .A2(n8718), .A3(n8717), .A4(n8716), .ZN(n11518) );
  AND2_X1 U10938 ( .A1(n14637), .A2(n11518), .ZN(n8721) );
  NAND2_X1 U10939 ( .A1(n10069), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n8722) );
  NAND2_X1 U10940 ( .A1(n8723), .A2(n8722), .ZN(n8725) );
  NAND2_X1 U10941 ( .A1(n10070), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n8724) );
  XNOR2_X1 U10942 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .ZN(n8738) );
  INV_X1 U10943 ( .A(n8738), .ZN(n8726) );
  XNOR2_X1 U10944 ( .A(n8739), .B(n8726), .ZN(n9836) );
  NAND2_X1 U10945 ( .A1(n9836), .A2(n12362), .ZN(n8729) );
  NAND2_X1 U10946 ( .A1(n8743), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8727) );
  XNOR2_X1 U10947 ( .A(n8727), .B(P3_IR_REG_12__SCAN_IN), .ZN(n12751) );
  AOI22_X1 U10948 ( .A1(n12370), .A2(SI_12_), .B1(n8858), .B2(n12751), .ZN(
        n8728) );
  NAND2_X1 U10949 ( .A1(n8729), .A2(n8728), .ZN(n14633) );
  NAND2_X1 U10950 ( .A1(n10792), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n8734) );
  NAND2_X1 U10951 ( .A1(n8861), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n8733) );
  OR2_X1 U10952 ( .A1(n6632), .A2(n8748), .ZN(n11583) );
  NAND2_X1 U10953 ( .A1(n8988), .A2(n11583), .ZN(n8732) );
  INV_X1 U10954 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n12746) );
  OR2_X1 U10955 ( .A1(n10796), .A2(n12746), .ZN(n8731) );
  NAND4_X1 U10956 ( .A1(n8734), .A2(n8733), .A3(n8732), .A4(n8731), .ZN(n12737) );
  NAND2_X1 U10957 ( .A1(n14633), .A2(n12737), .ZN(n8735) );
  NAND2_X1 U10958 ( .A1(n11622), .A2(n8735), .ZN(n8737) );
  OR2_X1 U10959 ( .A1(n14633), .A2(n12737), .ZN(n8736) );
  NAND2_X1 U10960 ( .A1(n8737), .A2(n8736), .ZN(n11718) );
  NAND2_X1 U10961 ( .A1(n8739), .A2(n8738), .ZN(n8742) );
  NAND2_X1 U10962 ( .A1(n8740), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n8741) );
  NAND2_X2 U10963 ( .A1(n8742), .A2(n8741), .ZN(n8758) );
  XNOR2_X2 U10964 ( .A(n8758), .B(P2_DATAO_REG_13__SCAN_IN), .ZN(n8757) );
  XNOR2_X1 U10965 ( .A(n8757), .B(P1_DATAO_REG_13__SCAN_IN), .ZN(n9908) );
  NAND2_X1 U10966 ( .A1(n9908), .A2(n12362), .ZN(n8747) );
  OR2_X1 U10967 ( .A1(n8743), .A2(P3_IR_REG_12__SCAN_IN), .ZN(n8761) );
  NAND2_X1 U10968 ( .A1(n8761), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8745) );
  XNOR2_X1 U10969 ( .A(n8745), .B(n8744), .ZN(n12772) );
  AOI22_X1 U10970 ( .A1(n12370), .A2(n9909), .B1(n8858), .B2(n12772), .ZN(
        n8746) );
  NAND2_X1 U10971 ( .A1(n8747), .A2(n8746), .ZN(n14625) );
  NAND2_X1 U10972 ( .A1(n9032), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n8753) );
  INV_X1 U10973 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n11439) );
  OR2_X1 U10974 ( .A1(n8748), .A2(n11439), .ZN(n8749) );
  NAND2_X1 U10975 ( .A1(n8767), .A2(n8749), .ZN(n11438) );
  NAND2_X1 U10976 ( .A1(n8988), .A2(n11438), .ZN(n8752) );
  NAND2_X1 U10977 ( .A1(n8861), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n8751) );
  INV_X1 U10978 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n11722) );
  OR2_X1 U10979 ( .A1(n10796), .A2(n11722), .ZN(n8750) );
  NAND4_X1 U10980 ( .A1(n8753), .A2(n8752), .A3(n8751), .A4(n8750), .ZN(n12736) );
  NOR2_X1 U10981 ( .A1(n14625), .A2(n12736), .ZN(n12490) );
  INV_X1 U10982 ( .A(n12490), .ZN(n8754) );
  NAND2_X1 U10983 ( .A1(n14625), .A2(n12736), .ZN(n12489) );
  NAND2_X1 U10984 ( .A1(n8754), .A2(n12489), .ZN(n12488) );
  NAND2_X1 U10985 ( .A1(n11718), .A2(n12488), .ZN(n8756) );
  INV_X1 U10986 ( .A(n12736), .ZN(n11789) );
  NAND2_X1 U10987 ( .A1(n14625), .A2(n11789), .ZN(n8755) );
  NAND2_X1 U10988 ( .A1(n8758), .A2(n15454), .ZN(n8759) );
  XNOR2_X1 U10989 ( .A(n10455), .B(P2_DATAO_REG_14__SCAN_IN), .ZN(n8760) );
  XNOR2_X1 U10990 ( .A(n8775), .B(n8760), .ZN(n10000) );
  NAND2_X1 U10991 ( .A1(n10000), .A2(n12362), .ZN(n8766) );
  OAI21_X1 U10992 ( .B1(n8761), .B2(P3_IR_REG_13__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8762) );
  MUX2_X1 U10993 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8762), .S(
        P3_IR_REG_14__SCAN_IN), .Z(n8764) );
  AND2_X1 U10994 ( .A1(n8764), .A2(n7331), .ZN(n12776) );
  AOI22_X1 U10995 ( .A1(n12370), .A2(SI_14_), .B1(n8858), .B2(n12776), .ZN(
        n8765) );
  NAND2_X1 U10996 ( .A1(n10792), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n8772) );
  NAND2_X1 U10997 ( .A1(n8767), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8768) );
  NAND2_X1 U10998 ( .A1(n8785), .A2(n8768), .ZN(n11643) );
  NAND2_X1 U10999 ( .A1(n8988), .A2(n11643), .ZN(n8771) );
  NAND2_X1 U11000 ( .A1(n8861), .A2(P3_REG0_REG_14__SCAN_IN), .ZN(n8770) );
  INV_X1 U11001 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n12769) );
  OR2_X1 U11002 ( .A1(n10796), .A2(n12769), .ZN(n8769) );
  NAND4_X1 U11003 ( .A1(n8772), .A2(n8771), .A3(n8770), .A4(n8769), .ZN(n11441) );
  OR2_X1 U11004 ( .A1(n13140), .A2(n13066), .ZN(n12497) );
  NAND2_X1 U11005 ( .A1(n13140), .A2(n13066), .ZN(n12496) );
  NAND2_X1 U11006 ( .A1(n12497), .A2(n12496), .ZN(n12492) );
  NAND2_X1 U11007 ( .A1(n13140), .A2(n11441), .ZN(n8773) );
  AND2_X1 U11008 ( .A1(n10453), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n8774) );
  NAND2_X1 U11009 ( .A1(n10455), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n8776) );
  NAND2_X1 U11010 ( .A1(n10558), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n8794) );
  NAND2_X1 U11011 ( .A1(n10559), .A2(P2_DATAO_REG_15__SCAN_IN), .ZN(n8777) );
  NAND2_X1 U11012 ( .A1(n8794), .A2(n8777), .ZN(n8795) );
  INV_X1 U11013 ( .A(n8795), .ZN(n8778) );
  XNOR2_X1 U11014 ( .A(n8796), .B(n8778), .ZN(n10102) );
  NAND2_X1 U11015 ( .A1(n10102), .A2(n12362), .ZN(n8784) );
  NOR2_X1 U11016 ( .A1(n8763), .A2(n13195), .ZN(n8779) );
  MUX2_X1 U11017 ( .A(n13195), .B(n8779), .S(P3_IR_REG_15__SCAN_IN), .Z(n8780)
         );
  INV_X1 U11018 ( .A(n8780), .ZN(n8782) );
  INV_X1 U11019 ( .A(n8817), .ZN(n8781) );
  NAND2_X1 U11020 ( .A1(n8782), .A2(n8781), .ZN(n12833) );
  INV_X1 U11021 ( .A(n12833), .ZN(n12824) );
  AOI22_X1 U11022 ( .A1(n12370), .A2(SI_15_), .B1(n8858), .B2(n12824), .ZN(
        n8783) );
  NAND2_X1 U11023 ( .A1(n8784), .A2(n8783), .ZN(n11712) );
  NAND2_X1 U11024 ( .A1(n10792), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n8790) );
  AND2_X1 U11025 ( .A1(n8785), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n8786) );
  OR2_X1 U11026 ( .A1(n8786), .A2(n8805), .ZN(n13073) );
  NAND2_X1 U11027 ( .A1(n8988), .A2(n13073), .ZN(n8789) );
  NAND2_X1 U11028 ( .A1(n10793), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n8788) );
  INV_X1 U11029 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n12801) );
  OR2_X1 U11030 ( .A1(n10796), .A2(n12801), .ZN(n8787) );
  NAND4_X1 U11031 ( .A1(n8790), .A2(n8789), .A3(n8788), .A4(n8787), .ZN(n12735) );
  OR2_X1 U11032 ( .A1(n11712), .A2(n12735), .ZN(n8791) );
  NAND2_X1 U11033 ( .A1(n11712), .A2(n12735), .ZN(n8792) );
  OAI21_X2 U11034 ( .B1(n8796), .B2(n8795), .A(n8794), .ZN(n8799) );
  NAND2_X1 U11035 ( .A1(n10421), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n8813) );
  NAND2_X1 U11036 ( .A1(n10424), .A2(P2_DATAO_REG_16__SCAN_IN), .ZN(n8797) );
  AND2_X1 U11037 ( .A1(n8813), .A2(n8797), .ZN(n8798) );
  OR2_X1 U11038 ( .A1(n8799), .A2(n8798), .ZN(n8800) );
  AND2_X1 U11039 ( .A1(n8814), .A2(n8800), .ZN(n10249) );
  NAND2_X1 U11040 ( .A1(n10249), .A2(n12362), .ZN(n8803) );
  OR2_X1 U11041 ( .A1(n8817), .A2(n13195), .ZN(n8801) );
  XNOR2_X1 U11042 ( .A(n8801), .B(P3_IR_REG_16__SCAN_IN), .ZN(n12837) );
  AOI22_X1 U11043 ( .A1(n12370), .A2(SI_16_), .B1(n8858), .B2(n12837), .ZN(
        n8802) );
  NAND2_X1 U11044 ( .A1(n10792), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n8810) );
  INV_X1 U11045 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n8804) );
  NOR2_X1 U11046 ( .A1(n8805), .A2(n8804), .ZN(n8806) );
  OR2_X1 U11047 ( .A1(n8822), .A2(n8806), .ZN(n13058) );
  NAND2_X1 U11048 ( .A1(n8988), .A2(n13058), .ZN(n8809) );
  NAND2_X1 U11049 ( .A1(n10793), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n8808) );
  INV_X1 U11050 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n12836) );
  OR2_X1 U11051 ( .A1(n10796), .A2(n12836), .ZN(n8807) );
  NAND4_X1 U11052 ( .A1(n8810), .A2(n8809), .A3(n8808), .A4(n8807), .ZN(n12734) );
  NOR2_X1 U11053 ( .A1(n13184), .A2(n13068), .ZN(n8812) );
  NAND2_X1 U11054 ( .A1(n13184), .A2(n13068), .ZN(n8811) );
  XNOR2_X1 U11055 ( .A(n10508), .B(P1_DATAO_REG_17__SCAN_IN), .ZN(n8815) );
  XNOR2_X1 U11056 ( .A(n8831), .B(n8815), .ZN(n10292) );
  NAND2_X1 U11057 ( .A1(n10292), .A2(n12362), .ZN(n8820) );
  INV_X1 U11058 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n8816) );
  NAND2_X1 U11059 ( .A1(n8817), .A2(n8816), .ZN(n8834) );
  NAND2_X1 U11060 ( .A1(n8834), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8818) );
  XNOR2_X1 U11061 ( .A(n8818), .B(P3_IR_REG_17__SCAN_IN), .ZN(n14580) );
  AOI22_X1 U11062 ( .A1(n12370), .A2(SI_17_), .B1(n8858), .B2(n14580), .ZN(
        n8819) );
  NAND2_X1 U11063 ( .A1(n10792), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n8828) );
  INV_X1 U11064 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n8821) );
  OR2_X1 U11065 ( .A1(n8822), .A2(n8821), .ZN(n8823) );
  NAND2_X1 U11066 ( .A1(n8843), .A2(n8823), .ZN(n13046) );
  NAND2_X1 U11067 ( .A1(n8988), .A2(n13046), .ZN(n8827) );
  NAND2_X1 U11068 ( .A1(n8861), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n8826) );
  INV_X1 U11069 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n8824) );
  OR2_X1 U11070 ( .A1(n10796), .A2(n8824), .ZN(n8825) );
  NAND4_X1 U11071 ( .A1(n8828), .A2(n8827), .A3(n8826), .A4(n8825), .ZN(n11782) );
  XNOR2_X1 U11072 ( .A(n13126), .B(n11782), .ZN(n13041) );
  NAND2_X1 U11073 ( .A1(n13126), .A2(n11782), .ZN(n8829) );
  AND2_X1 U11074 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n10508), .ZN(n8830) );
  NAND2_X1 U11075 ( .A1(n8832), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n8833) );
  INV_X1 U11076 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n10833) );
  INV_X1 U11077 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n10831) );
  AOI22_X1 U11078 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(n10833), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n10831), .ZN(n8850) );
  XNOR2_X1 U11079 ( .A(n8853), .B(n8850), .ZN(n10425) );
  NAND2_X1 U11080 ( .A1(n10425), .A2(n12362), .ZN(n8842) );
  NAND2_X1 U11081 ( .A1(n8836), .A2(n8835), .ZN(n8838) );
  NAND2_X1 U11082 ( .A1(n8838), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8837) );
  MUX2_X1 U11083 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8837), .S(
        P3_IR_REG_18__SCAN_IN), .Z(n8840) );
  INV_X1 U11084 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n8839) );
  NAND2_X1 U11085 ( .A1(n8840), .A2(n8855), .ZN(n12856) );
  INV_X1 U11086 ( .A(n12856), .ZN(n14592) );
  AOI22_X1 U11087 ( .A1(n12370), .A2(SI_18_), .B1(n8858), .B2(n14592), .ZN(
        n8841) );
  NAND2_X1 U11088 ( .A1(n8843), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8844) );
  NAND2_X1 U11089 ( .A1(n8862), .A2(n8844), .ZN(n12697) );
  NAND2_X1 U11090 ( .A1(n12697), .A2(n8988), .ZN(n8848) );
  NAND2_X1 U11091 ( .A1(n10792), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n8847) );
  NAND2_X1 U11092 ( .A1(n10793), .A2(P3_REG0_REG_18__SCAN_IN), .ZN(n8846) );
  INV_X1 U11093 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n13027) );
  OR2_X1 U11094 ( .A1(n10796), .A2(n13027), .ZN(n8845) );
  NAND4_X1 U11095 ( .A1(n8848), .A2(n8847), .A3(n8846), .A4(n8845), .ZN(n12733) );
  NAND2_X1 U11096 ( .A1(n13122), .A2(n13037), .ZN(n12517) );
  NAND2_X1 U11097 ( .A1(n12513), .A2(n12517), .ZN(n13029) );
  OR2_X1 U11098 ( .A1(n13122), .A2(n12733), .ZN(n8849) );
  INV_X1 U11099 ( .A(n8850), .ZN(n8852) );
  NAND2_X1 U11100 ( .A1(n10831), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n8851) );
  OAI21_X2 U11101 ( .B1(n8853), .B2(n8852), .A(n8851), .ZN(n8870) );
  INV_X1 U11102 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n12615) );
  INV_X1 U11103 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n10992) );
  AOI22_X1 U11104 ( .A1(P2_DATAO_REG_19__SCAN_IN), .A2(
        P1_DATAO_REG_19__SCAN_IN), .B1(n12615), .B2(n10992), .ZN(n8871) );
  XNOR2_X1 U11105 ( .A(n8870), .B(n7268), .ZN(n10477) );
  NAND2_X1 U11106 ( .A1(n10477), .A2(n12362), .ZN(n8860) );
  NAND2_X1 U11107 ( .A1(n8855), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8854) );
  MUX2_X1 U11108 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8854), .S(
        P3_IR_REG_19__SCAN_IN), .Z(n8857) );
  NAND2_X1 U11109 ( .A1(n8857), .A2(n9028), .ZN(n12859) );
  AOI22_X1 U11110 ( .A1(n12370), .A2(n10476), .B1(n8858), .B2(n12859), .ZN(
        n8859) );
  INV_X1 U11111 ( .A(n8861), .ZN(n8866) );
  INV_X1 U11112 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n13173) );
  AND2_X1 U11113 ( .A1(n8862), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8863) );
  OR2_X1 U11114 ( .A1(n8863), .A2(n8875), .ZN(n13016) );
  NAND2_X1 U11115 ( .A1(n13016), .A2(n8988), .ZN(n8865) );
  INV_X1 U11116 ( .A(n10796), .ZN(n8877) );
  AOI22_X1 U11117 ( .A1(n8877), .A2(P3_REG2_REG_19__SCAN_IN), .B1(n10792), 
        .B2(P3_REG1_REG_19__SCAN_IN), .ZN(n8864) );
  OAI211_X1 U11118 ( .C1(n8866), .C2(n13173), .A(n8865), .B(n8864), .ZN(n12995) );
  INV_X1 U11119 ( .A(n12523), .ZN(n8868) );
  INV_X1 U11120 ( .A(n13175), .ZN(n8867) );
  INV_X1 U11121 ( .A(n12995), .ZN(n13025) );
  NAND2_X1 U11122 ( .A1(n8867), .A2(n13025), .ZN(n12518) );
  OR2_X1 U11123 ( .A1(n13175), .A2(n13025), .ZN(n8869) );
  NAND2_X1 U11124 ( .A1(n13011), .A2(n8869), .ZN(n12994) );
  AOI22_X1 U11125 ( .A1(P2_DATAO_REG_20__SCAN_IN), .A2(
        P1_DATAO_REG_20__SCAN_IN), .B1(n15400), .B2(n15251), .ZN(n8882) );
  XNOR2_X1 U11126 ( .A(n8883), .B(n8882), .ZN(n10801) );
  NAND2_X1 U11127 ( .A1(n10801), .A2(n12362), .ZN(n8873) );
  INV_X1 U11128 ( .A(P3_REG3_REG_20__SCAN_IN), .ZN(n8874) );
  NOR2_X1 U11129 ( .A1(n8875), .A2(n8874), .ZN(n8876) );
  OR2_X1 U11130 ( .A1(n8887), .A2(n8876), .ZN(n12999) );
  NAND2_X1 U11131 ( .A1(n12999), .A2(n8988), .ZN(n8880) );
  AOI22_X1 U11132 ( .A1(n8877), .A2(P3_REG2_REG_20__SCAN_IN), .B1(n10792), 
        .B2(P3_REG1_REG_20__SCAN_IN), .ZN(n8879) );
  NAND2_X1 U11133 ( .A1(n10793), .A2(P3_REG0_REG_20__SCAN_IN), .ZN(n8878) );
  NAND2_X1 U11134 ( .A1(n12994), .A2(n13004), .ZN(n12993) );
  INV_X1 U11135 ( .A(n13009), .ZN(n12529) );
  NAND2_X1 U11136 ( .A1(n13000), .A2(n12529), .ZN(n8881) );
  NAND2_X1 U11137 ( .A1(n12993), .A2(n8881), .ZN(n12983) );
  INV_X1 U11138 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n11135) );
  AOI22_X1 U11139 ( .A1(P2_DATAO_REG_21__SCAN_IN), .A2(n11135), .B1(
        P1_DATAO_REG_21__SCAN_IN), .B2(n8900), .ZN(n8898) );
  INV_X1 U11140 ( .A(n8898), .ZN(n8884) );
  XNOR2_X1 U11141 ( .A(n8899), .B(n8884), .ZN(n11031) );
  NAND2_X1 U11142 ( .A1(n11031), .A2(n12362), .ZN(n8886) );
  NAND2_X1 U11143 ( .A1(n12363), .A2(SI_21_), .ZN(n8885) );
  INV_X1 U11144 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n12641) );
  OR2_X1 U11145 ( .A1(n8887), .A2(n12641), .ZN(n8888) );
  NAND2_X1 U11146 ( .A1(n8906), .A2(n8888), .ZN(n12988) );
  NAND2_X1 U11147 ( .A1(n12988), .A2(n8988), .ZN(n8894) );
  INV_X1 U11148 ( .A(P3_REG2_REG_21__SCAN_IN), .ZN(n8891) );
  NAND2_X1 U11149 ( .A1(n10792), .A2(P3_REG1_REG_21__SCAN_IN), .ZN(n8890) );
  NAND2_X1 U11150 ( .A1(n10793), .A2(P3_REG0_REG_21__SCAN_IN), .ZN(n8889) );
  OAI211_X1 U11151 ( .C1(n8891), .C2(n10796), .A(n8890), .B(n8889), .ZN(n8892)
         );
  INV_X1 U11152 ( .A(n8892), .ZN(n8893) );
  INV_X1 U11153 ( .A(n12974), .ZN(n12996) );
  OR2_X1 U11154 ( .A1(n12644), .A2(n12996), .ZN(n8895) );
  NAND2_X1 U11155 ( .A1(n12983), .A2(n8895), .ZN(n8897) );
  NAND2_X1 U11156 ( .A1(n12644), .A2(n12996), .ZN(n8896) );
  NAND2_X1 U11157 ( .A1(n8899), .A2(n8898), .ZN(n8902) );
  INV_X1 U11158 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8903) );
  INV_X1 U11159 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n15312) );
  AOI22_X1 U11160 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(
        P2_DATAO_REG_22__SCAN_IN), .B1(n8903), .B2(n15312), .ZN(n8916) );
  XNOR2_X1 U11161 ( .A(n8917), .B(n8916), .ZN(n11132) );
  NAND2_X1 U11162 ( .A1(n11132), .A2(n9017), .ZN(n8905) );
  NAND2_X1 U11163 ( .A1(n8906), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8907) );
  NAND2_X1 U11164 ( .A1(n8921), .A2(n8907), .ZN(n12978) );
  NAND2_X1 U11165 ( .A1(n12978), .A2(n8988), .ZN(n8913) );
  INV_X1 U11166 ( .A(P3_REG2_REG_22__SCAN_IN), .ZN(n8910) );
  NAND2_X1 U11167 ( .A1(n10793), .A2(P3_REG0_REG_22__SCAN_IN), .ZN(n8909) );
  NAND2_X1 U11168 ( .A1(n10792), .A2(P3_REG1_REG_22__SCAN_IN), .ZN(n8908) );
  OAI211_X1 U11169 ( .C1(n10796), .C2(n8910), .A(n8909), .B(n8908), .ZN(n8911)
         );
  INV_X1 U11170 ( .A(n8911), .ZN(n8912) );
  INV_X1 U11171 ( .A(n12985), .ZN(n12956) );
  AND2_X1 U11172 ( .A1(n12686), .A2(n12956), .ZN(n8915) );
  OR2_X1 U11173 ( .A1(n12686), .A2(n12956), .ZN(n8914) );
  NOR2_X1 U11174 ( .A1(n8917), .A2(n8916), .ZN(n8918) );
  INV_X1 U11175 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n15252) );
  AOI22_X1 U11176 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(
        P2_DATAO_REG_23__SCAN_IN), .B1(n11479), .B2(n15252), .ZN(n8930) );
  XNOR2_X1 U11177 ( .A(n8931), .B(n8930), .ZN(n11383) );
  NAND2_X1 U11178 ( .A1(n11383), .A2(n9017), .ZN(n8920) );
  NAND2_X1 U11179 ( .A1(n8921), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8922) );
  NAND2_X1 U11180 ( .A1(n8934), .A2(n8922), .ZN(n12967) );
  NAND2_X1 U11181 ( .A1(n12967), .A2(n8988), .ZN(n8928) );
  INV_X1 U11182 ( .A(P3_REG2_REG_23__SCAN_IN), .ZN(n8925) );
  NAND2_X1 U11183 ( .A1(n10793), .A2(P3_REG0_REG_23__SCAN_IN), .ZN(n8924) );
  NAND2_X1 U11184 ( .A1(n10792), .A2(P3_REG1_REG_23__SCAN_IN), .ZN(n8923) );
  OAI211_X1 U11185 ( .C1(n10796), .C2(n8925), .A(n8924), .B(n8923), .ZN(n8926)
         );
  INV_X1 U11186 ( .A(n8926), .ZN(n8927) );
  NAND2_X1 U11187 ( .A1(n8928), .A2(n8927), .ZN(n12732) );
  NAND2_X1 U11188 ( .A1(n12969), .A2(n12732), .ZN(n9058) );
  INV_X1 U11189 ( .A(n12732), .ZN(n12975) );
  NAND2_X1 U11190 ( .A1(n13101), .A2(n12975), .ZN(n8929) );
  NAND2_X1 U11191 ( .A1(n9058), .A2(n8929), .ZN(n12960) );
  NAND2_X1 U11192 ( .A1(n13101), .A2(n12732), .ZN(n12935) );
  INV_X1 U11193 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n11615) );
  XNOR2_X1 U11194 ( .A(n11615), .B(n8944), .ZN(n11745) );
  NAND2_X1 U11195 ( .A1(n11745), .A2(n12362), .ZN(n8933) );
  NAND2_X1 U11196 ( .A1(n12370), .A2(SI_24_), .ZN(n8932) );
  AND2_X1 U11197 ( .A1(n8934), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n8935) );
  OR2_X1 U11198 ( .A1(n8935), .A2(n8951), .ZN(n12948) );
  NAND2_X1 U11199 ( .A1(n12948), .A2(n8988), .ZN(n8941) );
  INV_X1 U11200 ( .A(P3_REG2_REG_24__SCAN_IN), .ZN(n8938) );
  NAND2_X1 U11201 ( .A1(n10793), .A2(P3_REG0_REG_24__SCAN_IN), .ZN(n8937) );
  NAND2_X1 U11202 ( .A1(n10792), .A2(P3_REG1_REG_24__SCAN_IN), .ZN(n8936) );
  OAI211_X1 U11203 ( .C1(n10796), .C2(n8938), .A(n8937), .B(n8936), .ZN(n8939)
         );
  INV_X1 U11204 ( .A(n8939), .ZN(n8940) );
  NAND2_X1 U11205 ( .A1(n8941), .A2(n8940), .ZN(n12957) );
  NAND2_X1 U11206 ( .A1(n9057), .A2(n12957), .ZN(n8942) );
  AND2_X1 U11207 ( .A1(n12935), .A2(n8942), .ZN(n12918) );
  NAND2_X1 U11208 ( .A1(n8943), .A2(n11617), .ZN(n8946) );
  NAND2_X1 U11209 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n8944), .ZN(n8945) );
  AOI22_X1 U11210 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n8965), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n11651), .ZN(n8963) );
  INV_X1 U11211 ( .A(n8963), .ZN(n8947) );
  XNOR2_X1 U11212 ( .A(n8964), .B(n8947), .ZN(n11799) );
  NAND2_X1 U11213 ( .A1(n11799), .A2(n12362), .ZN(n8949) );
  NAND2_X1 U11214 ( .A1(n12363), .A2(SI_25_), .ZN(n8948) );
  NAND2_X2 U11215 ( .A1(n8949), .A2(n8948), .ZN(n12548) );
  INV_X1 U11216 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n8950) );
  NAND2_X1 U11217 ( .A1(n8951), .A2(n8950), .ZN(n8970) );
  OR2_X1 U11218 ( .A1(n8951), .A2(n8950), .ZN(n8952) );
  NAND2_X1 U11219 ( .A1(n8970), .A2(n8952), .ZN(n12930) );
  NAND2_X1 U11220 ( .A1(n12930), .A2(n8988), .ZN(n8958) );
  INV_X1 U11221 ( .A(P3_REG2_REG_25__SCAN_IN), .ZN(n8955) );
  NAND2_X1 U11222 ( .A1(n10793), .A2(P3_REG0_REG_25__SCAN_IN), .ZN(n8954) );
  NAND2_X1 U11223 ( .A1(n10792), .A2(P3_REG1_REG_25__SCAN_IN), .ZN(n8953) );
  OAI211_X1 U11224 ( .C1(n10796), .C2(n8955), .A(n8954), .B(n8953), .ZN(n8956)
         );
  INV_X1 U11225 ( .A(n8956), .ZN(n8957) );
  NAND2_X1 U11226 ( .A1(n8958), .A2(n8957), .ZN(n12905) );
  NAND2_X1 U11227 ( .A1(n12548), .A2(n12905), .ZN(n8959) );
  AND2_X1 U11228 ( .A1(n12918), .A2(n8959), .ZN(n8962) );
  INV_X1 U11229 ( .A(n8959), .ZN(n8961) );
  INV_X1 U11230 ( .A(n12923), .ZN(n12921) );
  NAND2_X1 U11231 ( .A1(n13159), .A2(n12925), .ZN(n12919) );
  AND2_X1 U11232 ( .A1(n12921), .A2(n12919), .ZN(n8960) );
  AOI22_X1 U11233 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(n11817), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n11821), .ZN(n8980) );
  INV_X1 U11234 ( .A(n8980), .ZN(n8967) );
  XNOR2_X1 U11235 ( .A(n8979), .B(n8967), .ZN(n13214) );
  NAND2_X1 U11236 ( .A1(n13214), .A2(n12362), .ZN(n8969) );
  NAND2_X1 U11237 ( .A1(n12363), .A2(SI_26_), .ZN(n8968) );
  NAND2_X1 U11238 ( .A1(n8970), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8971) );
  NAND2_X1 U11239 ( .A1(n8985), .A2(n8971), .ZN(n12909) );
  NAND2_X1 U11240 ( .A1(n12909), .A2(n8988), .ZN(n8976) );
  INV_X1 U11241 ( .A(P3_REG2_REG_26__SCAN_IN), .ZN(n12910) );
  NAND2_X1 U11242 ( .A1(n10793), .A2(P3_REG0_REG_26__SCAN_IN), .ZN(n8973) );
  NAND2_X1 U11243 ( .A1(n10792), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n8972) );
  OAI211_X1 U11244 ( .C1(n10796), .C2(n12910), .A(n8973), .B(n8972), .ZN(n8974) );
  INV_X1 U11245 ( .A(n8974), .ZN(n8975) );
  AND2_X1 U11246 ( .A1(n12913), .A2(n12657), .ZN(n8978) );
  OAI21_X2 U11247 ( .B1(P2_DATAO_REG_26__SCAN_IN), .B2(n11817), .A(n8981), 
        .ZN(n8997) );
  INV_X1 U11248 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n12312) );
  AOI22_X1 U11249 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(n12312), .B1(
        P1_DATAO_REG_27__SCAN_IN), .B2(n11873), .ZN(n8998) );
  INV_X1 U11250 ( .A(n8998), .ZN(n8982) );
  XNOR2_X1 U11251 ( .A(n8997), .B(n8982), .ZN(n13208) );
  NAND2_X1 U11252 ( .A1(n13208), .A2(n12362), .ZN(n8984) );
  NAND2_X1 U11253 ( .A1(n12363), .A2(SI_27_), .ZN(n8983) );
  INV_X1 U11254 ( .A(n9003), .ZN(n8987) );
  NAND2_X1 U11255 ( .A1(n8985), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n8986) );
  NAND2_X1 U11256 ( .A1(n8987), .A2(n8986), .ZN(n12894) );
  NAND2_X1 U11257 ( .A1(n12894), .A2(n8988), .ZN(n8994) );
  INV_X1 U11258 ( .A(P3_REG2_REG_27__SCAN_IN), .ZN(n8991) );
  NAND2_X1 U11259 ( .A1(n10792), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n8990) );
  NAND2_X1 U11260 ( .A1(n10793), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n8989) );
  OAI211_X1 U11261 ( .C1(n8991), .C2(n10796), .A(n8990), .B(n8989), .ZN(n8992)
         );
  INV_X1 U11262 ( .A(n8992), .ZN(n8993) );
  OR2_X2 U11263 ( .A1(n13084), .A2(n9745), .ZN(n12559) );
  NAND2_X1 U11264 ( .A1(n12890), .A2(n12382), .ZN(n8996) );
  OR2_X1 U11265 ( .A1(n13084), .A2(n12906), .ZN(n8995) );
  NAND2_X1 U11266 ( .A1(n8996), .A2(n8995), .ZN(n12873) );
  NAND2_X1 U11267 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n11873), .ZN(n8999) );
  AOI22_X1 U11268 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(n13779), .B1(
        P1_DATAO_REG_28__SCAN_IN), .B2(n12607), .ZN(n9014) );
  NAND2_X1 U11269 ( .A1(n12363), .A2(SI_28_), .ZN(n9000) );
  NAND2_X2 U11270 ( .A1(n9001), .A2(n9000), .ZN(n12882) );
  INV_X1 U11271 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n9002) );
  NOR2_X1 U11272 ( .A1(n9003), .A2(n9002), .ZN(n9004) );
  INV_X1 U11273 ( .A(P3_REG2_REG_28__SCAN_IN), .ZN(n9007) );
  NAND2_X1 U11274 ( .A1(n10792), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n9006) );
  NAND2_X1 U11275 ( .A1(n10793), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n9005) );
  OAI211_X1 U11276 ( .C1(n9007), .C2(n10796), .A(n9006), .B(n9005), .ZN(n9008)
         );
  AOI21_X1 U11277 ( .B1(n12883), .B2(n8988), .A(n9008), .ZN(n15223) );
  OR2_X2 U11278 ( .A1(n12882), .A2(n15223), .ZN(n12562) );
  NAND2_X1 U11279 ( .A1(n12882), .A2(n15223), .ZN(n9061) );
  NAND2_X2 U11280 ( .A1(n12562), .A2(n9061), .ZN(n12560) );
  INV_X1 U11281 ( .A(n15223), .ZN(n12622) );
  NAND2_X1 U11282 ( .A1(n12882), .A2(n12622), .ZN(n9009) );
  NAND2_X1 U11283 ( .A1(n12875), .A2(n9009), .ZN(n9020) );
  NAND2_X1 U11284 ( .A1(n14611), .A2(n8988), .ZN(n10799) );
  INV_X1 U11285 ( .A(P3_REG2_REG_29__SCAN_IN), .ZN(n11991) );
  NAND2_X1 U11286 ( .A1(n10792), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n9011) );
  INV_X1 U11287 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n15437) );
  OR2_X1 U11288 ( .A1(n8866), .A2(n15437), .ZN(n9010) );
  OAI211_X1 U11289 ( .C1(n11991), .C2(n10796), .A(n9011), .B(n9010), .ZN(n9012) );
  INV_X1 U11290 ( .A(n9012), .ZN(n9013) );
  NAND2_X1 U11291 ( .A1(n10799), .A2(n9013), .ZN(n12876) );
  AOI22_X1 U11292 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n14434), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n15332), .ZN(n9016) );
  NAND2_X1 U11293 ( .A1(n9017), .A2(n13201), .ZN(n9019) );
  NAND2_X1 U11294 ( .A1(n12363), .A2(SI_29_), .ZN(n9018) );
  XNOR2_X1 U11295 ( .A(n9020), .B(n9065), .ZN(n9040) );
  INV_X1 U11296 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n9021) );
  OAI21_X1 U11297 ( .B1(n9025), .B2(P3_IR_REG_21__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9023) );
  MUX2_X1 U11298 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9023), .S(
        P3_IR_REG_22__SCAN_IN), .Z(n9024) );
  OR2_X1 U11299 ( .A1(n12416), .A2(n12859), .ZN(n9121) );
  NAND2_X1 U11300 ( .A1(n9025), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9027) );
  INV_X1 U11301 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n9026) );
  INV_X1 U11302 ( .A(n12419), .ZN(n10733) );
  NAND2_X1 U11303 ( .A1(n9028), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9029) );
  XNOR2_X1 U11304 ( .A(n9029), .B(P3_IR_REG_20__SCAN_IN), .ZN(n9626) );
  NAND2_X1 U11305 ( .A1(n10733), .A2(n9626), .ZN(n12408) );
  NAND2_X1 U11306 ( .A1(n9121), .A2(n12408), .ZN(n15143) );
  OR2_X2 U11307 ( .A1(n12416), .A2(n12419), .ZN(n9115) );
  INV_X1 U11308 ( .A(n13205), .ZN(n10201) );
  INV_X1 U11309 ( .A(n9030), .ZN(n10218) );
  NAND2_X1 U11310 ( .A1(n10201), .A2(n10218), .ZN(n10202) );
  NAND2_X1 U11311 ( .A1(n10198), .A2(n10202), .ZN(n12581) );
  INV_X1 U11312 ( .A(n12581), .ZN(n9031) );
  NAND2_X1 U11313 ( .A1(n12549), .A2(n9031), .ZN(n13067) );
  INV_X1 U11314 ( .A(P3_REG2_REG_30__SCAN_IN), .ZN(n9035) );
  NAND2_X1 U11315 ( .A1(n10793), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n9034) );
  NAND2_X1 U11316 ( .A1(n9032), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n9033) );
  OAI211_X1 U11317 ( .C1(n10796), .C2(n9035), .A(n9034), .B(n9033), .ZN(n9036)
         );
  INV_X1 U11318 ( .A(n9036), .ZN(n9037) );
  AND2_X1 U11319 ( .A1(n10799), .A2(n9037), .ZN(n12373) );
  INV_X1 U11320 ( .A(P3_B_REG_SCAN_IN), .ZN(n15484) );
  NOR2_X1 U11321 ( .A1(n13205), .A2(n15484), .ZN(n9038) );
  OR2_X1 U11322 ( .A1(n13069), .A2(n9038), .ZN(n14609) );
  OAI22_X1 U11323 ( .A1(n15223), .A2(n13067), .B1(n12373), .B2(n14609), .ZN(
        n9039) );
  AOI21_X1 U11324 ( .B1(n9040), .B2(n15143), .A(n9039), .ZN(n11996) );
  AND2_X2 U11325 ( .A1(n9042), .A2(n9041), .ZN(n15135) );
  NAND2_X1 U11326 ( .A1(n12418), .A2(n15135), .ZN(n9634) );
  NAND2_X1 U11327 ( .A1(n9634), .A2(n12422), .ZN(n15116) );
  NAND2_X1 U11328 ( .A1(n15116), .A2(n15124), .ZN(n9043) );
  NAND2_X1 U11329 ( .A1(n9043), .A2(n12427), .ZN(n11195) );
  NAND2_X1 U11330 ( .A1(n11195), .A2(n12385), .ZN(n11197) );
  NAND2_X1 U11331 ( .A1(n11197), .A2(n12431), .ZN(n10729) );
  NAND2_X1 U11332 ( .A1(n10729), .A2(n12433), .ZN(n9044) );
  NAND2_X1 U11333 ( .A1(n9044), .A2(n12440), .ZN(n11068) );
  NAND2_X1 U11334 ( .A1(n11068), .A2(n12437), .ZN(n9045) );
  NAND2_X1 U11335 ( .A1(n9046), .A2(n12454), .ZN(n11207) );
  INV_X1 U11336 ( .A(n12460), .ZN(n15188) );
  OR2_X1 U11337 ( .A1(n12740), .A2(n15188), .ZN(n12459) );
  NAND2_X1 U11338 ( .A1(n12739), .A2(n15193), .ZN(n9047) );
  NAND2_X1 U11339 ( .A1(n9048), .A2(n9047), .ZN(n11446) );
  OR2_X1 U11340 ( .A1(n14637), .A2(n11624), .ZN(n12473) );
  NAND2_X1 U11341 ( .A1(n14637), .A2(n11624), .ZN(n12479) );
  OR2_X1 U11342 ( .A1(n14633), .A2(n11720), .ZN(n12474) );
  NAND2_X1 U11343 ( .A1(n14633), .A2(n11720), .ZN(n12478) );
  INV_X1 U11344 ( .A(n12492), .ZN(n9050) );
  OR2_X1 U11345 ( .A1(n11712), .A2(n13054), .ZN(n12502) );
  NAND2_X1 U11346 ( .A1(n11712), .A2(n13054), .ZN(n12508) );
  NAND2_X1 U11347 ( .A1(n13070), .A2(n12508), .ZN(n13057) );
  NAND2_X1 U11348 ( .A1(n13184), .A2(n12734), .ZN(n12509) );
  INV_X1 U11349 ( .A(n13184), .ZN(n9051) );
  NAND2_X1 U11350 ( .A1(n9051), .A2(n13068), .ZN(n13042) );
  NAND2_X1 U11351 ( .A1(n13055), .A2(n13042), .ZN(n9052) );
  INV_X1 U11352 ( .A(n11782), .ZN(n13053) );
  NAND2_X1 U11353 ( .A1(n13126), .A2(n13053), .ZN(n12516) );
  NAND2_X1 U11354 ( .A1(n13032), .A2(n12513), .ZN(n13015) );
  OR2_X1 U11355 ( .A1(n13000), .A2(n13009), .ZN(n12528) );
  NAND2_X1 U11356 ( .A1(n13001), .A2(n12528), .ZN(n12987) );
  NAND2_X1 U11357 ( .A1(n12644), .A2(n12974), .ZN(n9055) );
  NOR2_X1 U11358 ( .A1(n12644), .A2(n12974), .ZN(n9054) );
  AOI21_X2 U11359 ( .B1(n12987), .B2(n9055), .A(n9054), .ZN(n12977) );
  NAND2_X1 U11360 ( .A1(n12977), .A2(n12410), .ZN(n12959) );
  NAND2_X1 U11361 ( .A1(n12686), .A2(n12985), .ZN(n12958) );
  NAND2_X1 U11362 ( .A1(n12959), .A2(n9056), .ZN(n12937) );
  NAND2_X1 U11363 ( .A1(n13159), .A2(n12957), .ZN(n12540) );
  NAND2_X1 U11364 ( .A1(n12540), .A2(n12542), .ZN(n12938) );
  INV_X1 U11365 ( .A(n9058), .ZN(n12939) );
  NOR2_X1 U11366 ( .A1(n12938), .A2(n12939), .ZN(n9059) );
  INV_X1 U11367 ( .A(n12905), .ZN(n12943) );
  NAND2_X1 U11368 ( .A1(n12913), .A2(n12926), .ZN(n12553) );
  INV_X2 U11369 ( .A(n12382), .ZN(n12889) );
  AND2_X1 U11370 ( .A1(n12889), .A2(n12562), .ZN(n9060) );
  NAND2_X1 U11371 ( .A1(n12888), .A2(n9060), .ZN(n9064) );
  INV_X1 U11372 ( .A(n12562), .ZN(n9062) );
  AND2_X1 U11373 ( .A1(n9061), .A2(n12879), .ZN(n12561) );
  INV_X1 U11374 ( .A(n9626), .ZN(n10804) );
  NAND2_X1 U11375 ( .A1(n12419), .A2(n10804), .ZN(n9119) );
  XNOR2_X1 U11376 ( .A(n9119), .B(n12416), .ZN(n9067) );
  AND2_X1 U11377 ( .A1(n12419), .A2(n12859), .ZN(n9066) );
  AND2_X1 U11378 ( .A1(n15200), .A2(n12578), .ZN(n9068) );
  NAND2_X1 U11379 ( .A1(n9730), .A2(n9068), .ZN(n9070) );
  NAND2_X1 U11380 ( .A1(n9626), .A2(n12859), .ZN(n9069) );
  OR2_X1 U11381 ( .A1(n12416), .A2(n9069), .ZN(n10384) );
  INV_X1 U11382 ( .A(n12859), .ZN(n9071) );
  NAND2_X1 U11383 ( .A1(n12416), .A2(n15134), .ZN(n15194) );
  NAND2_X1 U11384 ( .A1(n15147), .A2(n15194), .ZN(n13139) );
  NAND2_X1 U11385 ( .A1(n11993), .A2(n13139), .ZN(n9072) );
  INV_X1 U11386 ( .A(n9121), .ZN(n9074) );
  INV_X1 U11387 ( .A(n12407), .ZN(n9073) );
  NAND2_X1 U11388 ( .A1(n9074), .A2(n9073), .ZN(n9735) );
  MUX2_X1 U11389 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9075), .S(
        P3_IR_REG_26__SCAN_IN), .Z(n9077) );
  NAND2_X1 U11390 ( .A1(n9078), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9079) );
  XNOR2_X1 U11391 ( .A(n9079), .B(P3_IR_REG_25__SCAN_IN), .ZN(n9094) );
  NAND2_X1 U11392 ( .A1(n9081), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9082) );
  XNOR2_X1 U11393 ( .A(n9082), .B(P3_IR_REG_24__SCAN_IN), .ZN(n9090) );
  AND2_X1 U11394 ( .A1(n9094), .A2(n9090), .ZN(n9083) );
  NAND2_X1 U11395 ( .A1(n9089), .A2(n9083), .ZN(n9753) );
  NAND2_X1 U11396 ( .A1(n6572), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9085) );
  XNOR2_X1 U11397 ( .A(n9085), .B(n9084), .ZN(n10197) );
  AND2_X1 U11398 ( .A1(n10197), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13193) );
  NAND2_X1 U11399 ( .A1(n9753), .A2(n13193), .ZN(n10200) );
  NOR2_X1 U11400 ( .A1(n10200), .A2(n9740), .ZN(n9086) );
  NAND2_X1 U11401 ( .A1(n12549), .A2(n9086), .ZN(n12582) );
  OAI21_X1 U11402 ( .B1(n9735), .B2(n10200), .A(n12582), .ZN(n9107) );
  XNOR2_X1 U11403 ( .A(n9090), .B(P3_B_REG_SCAN_IN), .ZN(n9087) );
  OR2_X1 U11404 ( .A1(n9087), .A2(n9094), .ZN(n9088) );
  INV_X1 U11405 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n15450) );
  NAND2_X1 U11406 ( .A1(n9805), .A2(n15450), .ZN(n9092) );
  INV_X1 U11407 ( .A(n9089), .ZN(n13218) );
  INV_X1 U11408 ( .A(n9090), .ZN(n11748) );
  NAND2_X1 U11409 ( .A1(n13218), .A2(n11748), .ZN(n9091) );
  INV_X1 U11410 ( .A(P3_D_REG_1__SCAN_IN), .ZN(n9093) );
  NAND2_X1 U11411 ( .A1(n9805), .A2(n9093), .ZN(n9096) );
  INV_X1 U11412 ( .A(n9094), .ZN(n11802) );
  NAND2_X1 U11413 ( .A1(n13218), .A2(n11802), .ZN(n9095) );
  NOR4_X1 U11414 ( .A1(P3_D_REG_9__SCAN_IN), .A2(P3_D_REG_17__SCAN_IN), .A3(
        P3_D_REG_22__SCAN_IN), .A4(P3_D_REG_25__SCAN_IN), .ZN(n9105) );
  INV_X1 U11415 ( .A(P3_D_REG_7__SCAN_IN), .ZN(n15226) );
  INV_X1 U11416 ( .A(P3_D_REG_28__SCAN_IN), .ZN(n15254) );
  INV_X1 U11417 ( .A(P3_D_REG_14__SCAN_IN), .ZN(n15265) );
  INV_X1 U11418 ( .A(P3_D_REG_26__SCAN_IN), .ZN(n15365) );
  NAND4_X1 U11419 ( .A1(n15226), .A2(n15254), .A3(n15265), .A4(n15365), .ZN(
        n9102) );
  NOR4_X1 U11420 ( .A1(P3_D_REG_21__SCAN_IN), .A2(P3_D_REG_12__SCAN_IN), .A3(
        P3_D_REG_11__SCAN_IN), .A4(P3_D_REG_16__SCAN_IN), .ZN(n9100) );
  NOR4_X1 U11421 ( .A1(P3_D_REG_10__SCAN_IN), .A2(P3_D_REG_24__SCAN_IN), .A3(
        P3_D_REG_29__SCAN_IN), .A4(P3_D_REG_31__SCAN_IN), .ZN(n9099) );
  NOR4_X1 U11422 ( .A1(P3_D_REG_6__SCAN_IN), .A2(P3_D_REG_3__SCAN_IN), .A3(
        P3_D_REG_5__SCAN_IN), .A4(P3_D_REG_8__SCAN_IN), .ZN(n9098) );
  NOR4_X1 U11423 ( .A1(P3_D_REG_15__SCAN_IN), .A2(P3_D_REG_30__SCAN_IN), .A3(
        P3_D_REG_13__SCAN_IN), .A4(P3_D_REG_23__SCAN_IN), .ZN(n9097) );
  NAND4_X1 U11424 ( .A1(n9100), .A2(n9099), .A3(n9098), .A4(n9097), .ZN(n9101)
         );
  NOR4_X1 U11425 ( .A1(P3_D_REG_4__SCAN_IN), .A2(P3_D_REG_2__SCAN_IN), .A3(
        n9102), .A4(n9101), .ZN(n9104) );
  NOR4_X1 U11426 ( .A1(P3_D_REG_20__SCAN_IN), .A2(P3_D_REG_19__SCAN_IN), .A3(
        P3_D_REG_18__SCAN_IN), .A4(P3_D_REG_27__SCAN_IN), .ZN(n9103) );
  NAND3_X1 U11427 ( .A1(n9105), .A2(n9104), .A3(n9103), .ZN(n9106) );
  NAND2_X1 U11428 ( .A1(n9805), .A2(n9106), .ZN(n9116) );
  AND3_X1 U11429 ( .A1(n7329), .A2(n13192), .A3(n9116), .ZN(n9729) );
  NAND2_X1 U11430 ( .A1(n9107), .A2(n9729), .ZN(n9110) );
  NAND2_X1 U11431 ( .A1(n9625), .A2(n9116), .ZN(n9108) );
  NOR2_X1 U11432 ( .A1(n9108), .A2(n13192), .ZN(n9737) );
  INV_X1 U11433 ( .A(n10200), .ZN(n9725) );
  AND2_X1 U11434 ( .A1(n9737), .A2(n9725), .ZN(n9742) );
  NAND2_X1 U11435 ( .A1(n9742), .A2(n9730), .ZN(n9109) );
  OR2_X1 U11436 ( .A1(n15206), .A2(n15200), .ZN(n13188) );
  NAND2_X1 U11437 ( .A1(n15206), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n9111) );
  INV_X1 U11438 ( .A(n9112), .ZN(n9113) );
  MUX2_X1 U11439 ( .A(n9740), .B(n10384), .S(n9115), .Z(n10385) );
  NAND2_X1 U11440 ( .A1(n10385), .A2(n13192), .ZN(n9125) );
  XNOR2_X1 U11441 ( .A(n13192), .B(n9625), .ZN(n9118) );
  AND2_X1 U11442 ( .A1(n9725), .A2(n9116), .ZN(n9117) );
  NAND2_X1 U11443 ( .A1(n9119), .A2(n12416), .ZN(n9120) );
  NAND3_X1 U11444 ( .A1(n9121), .A2(n9740), .A3(n9120), .ZN(n9122) );
  NAND2_X1 U11445 ( .A1(n9122), .A2(n9115), .ZN(n9123) );
  INV_X1 U11446 ( .A(n13192), .ZN(n10388) );
  NAND2_X1 U11447 ( .A1(n9123), .A2(n10388), .ZN(n9124) );
  AND3_X2 U11448 ( .A1(n9125), .A2(n10386), .A3(n9124), .ZN(n15222) );
  INV_X1 U11449 ( .A(n12375), .ZN(n9129) );
  INV_X1 U11450 ( .A(n15200), .ZN(n14638) );
  NAND2_X1 U11451 ( .A1(n15222), .A2(n14638), .ZN(n13138) );
  NAND2_X1 U11452 ( .A1(n9129), .A2(n9128), .ZN(n9132) );
  INV_X1 U11453 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n9130) );
  OR2_X1 U11454 ( .A1(n15222), .A2(n9130), .ZN(n9131) );
  NAND2_X1 U11455 ( .A1(n9134), .A2(n9133), .ZN(P3_U3488) );
  NOR2_X1 U11456 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n9137) );
  AND4_X2 U11457 ( .A1(n9137), .A2(n9136), .A3(n9135), .A4(n9295), .ZN(n9311)
         );
  NOR3_X2 U11458 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), 
        .A3(P2_IR_REG_13__SCAN_IN), .ZN(n9140) );
  NOR2_X1 U11459 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), 
        .ZN(n9143) );
  NOR2_X1 U11460 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), 
        .ZN(n9142) );
  NOR2_X1 U11461 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), 
        .ZN(n9141) );
  INV_X1 U11462 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n9145) );
  INV_X1 U11463 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n9595) );
  INV_X1 U11464 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n9155) );
  AND2_X1 U11465 ( .A1(n9155), .A2(n9157), .ZN(n9146) );
  INV_X1 U11466 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n13767) );
  INV_X1 U11467 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n9859) );
  INV_X1 U11468 ( .A(n12612), .ZN(n9148) );
  INV_X1 U11469 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n10027) );
  OR2_X1 U11470 ( .A1(n9476), .A2(n10027), .ZN(n9153) );
  NAND2_X1 U11471 ( .A1(n12162), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n9152) );
  INV_X1 U11472 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n9150) );
  OR2_X1 U11473 ( .A1(n6546), .A2(n9150), .ZN(n9151) );
  NAND4_X2 U11474 ( .A1(n9154), .A2(n9153), .A3(n9152), .A4(n9151), .ZN(n13374) );
  INV_X1 U11475 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n9160) );
  INV_X1 U11476 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n9159) );
  NAND2_X1 U11477 ( .A1(n9160), .A2(n9159), .ZN(n9179) );
  INV_X1 U11478 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n9162) );
  OR2_X1 U11479 ( .A1(n9172), .A2(n9162), .ZN(n9168) );
  INV_X1 U11480 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n9163) );
  NAND2_X1 U11481 ( .A1(n12162), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n9166) );
  INV_X1 U11482 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n9164) );
  XNOR2_X1 U11483 ( .A(n9169), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n13781) );
  INV_X1 U11484 ( .A(n12002), .ZN(n12003) );
  OR2_X1 U11485 ( .A1(n13375), .A2(n12003), .ZN(n10009) );
  INV_X1 U11486 ( .A(n10009), .ZN(n10062) );
  NAND2_X1 U11487 ( .A1(n12247), .A2(n10062), .ZN(n9171) );
  INV_X1 U11488 ( .A(n14934), .ZN(n10193) );
  OR2_X1 U11489 ( .A1(n13374), .A2(n10193), .ZN(n9170) );
  NAND2_X1 U11490 ( .A1(n9171), .A2(n9170), .ZN(n10077) );
  NAND2_X1 U11491 ( .A1(n12162), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n9176) );
  INV_X1 U11492 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n10101) );
  OR2_X1 U11493 ( .A1(n9476), .A2(n10101), .ZN(n9175) );
  INV_X1 U11494 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n9862) );
  INV_X1 U11495 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n9173) );
  NAND2_X1 U11496 ( .A1(n9179), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9178) );
  MUX2_X1 U11497 ( .A(n9178), .B(P2_IR_REG_31__SCAN_IN), .S(n9180), .Z(n9182)
         );
  INV_X1 U11498 ( .A(n9179), .ZN(n9181) );
  NAND2_X1 U11499 ( .A1(n9181), .A2(n9180), .ZN(n9187) );
  NAND2_X1 U11500 ( .A1(n9182), .A2(n9187), .ZN(n9861) );
  OAI22_X1 U11501 ( .A1(n9403), .A2(n10028), .B1(n9841), .B2(n9861), .ZN(n9183) );
  NAND2_X1 U11502 ( .A1(n10077), .A2(n12248), .ZN(n9185) );
  INV_X1 U11503 ( .A(n12016), .ZN(n11039) );
  OR2_X1 U11504 ( .A1(n13373), .A2(n11039), .ZN(n9184) );
  NAND2_X1 U11505 ( .A1(n9755), .A2(n12168), .ZN(n9190) );
  INV_X2 U11506 ( .A(n9403), .ZN(n9392) );
  INV_X2 U11507 ( .A(n9841), .ZN(n9391) );
  NAND2_X1 U11508 ( .A1(n9187), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9186) );
  MUX2_X1 U11509 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9186), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n9188) );
  OR2_X1 U11510 ( .A1(n9187), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n9199) );
  AOI22_X1 U11511 ( .A1(n9392), .A2(P1_DATAO_REG_3__SCAN_IN), .B1(n9391), .B2(
        n9863), .ZN(n9189) );
  NAND2_X1 U11512 ( .A1(n12162), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n9195) );
  OR2_X1 U11513 ( .A1(n9476), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n9194) );
  INV_X1 U11514 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n9864) );
  OR2_X1 U11515 ( .A1(n9496), .A2(n9864), .ZN(n9193) );
  INV_X1 U11516 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n9191) );
  OR2_X1 U11517 ( .A1(n6546), .A2(n9191), .ZN(n9192) );
  OR2_X1 U11518 ( .A1(n13372), .A2(n10946), .ZN(n9197) );
  NAND2_X1 U11519 ( .A1(n9198), .A2(n9197), .ZN(n10241) );
  NAND2_X1 U11520 ( .A1(n9767), .A2(n12168), .ZN(n9205) );
  NAND2_X1 U11521 ( .A1(n9199), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9200) );
  MUX2_X1 U11522 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9200), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n9203) );
  INV_X1 U11523 ( .A(n9310), .ZN(n9202) );
  NAND2_X1 U11524 ( .A1(n9203), .A2(n9202), .ZN(n14837) );
  INV_X1 U11525 ( .A(n14837), .ZN(n9850) );
  AOI22_X1 U11526 ( .A1(n9392), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n9391), .B2(
        n9850), .ZN(n9204) );
  NAND2_X1 U11527 ( .A1(n9524), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n9210) );
  INV_X2 U11528 ( .A(n12162), .ZN(n12196) );
  INV_X1 U11529 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n9206) );
  OR2_X1 U11530 ( .A1(n12196), .A2(n9206), .ZN(n9209) );
  XNOR2_X1 U11531 ( .A(P2_REG3_REG_3__SCAN_IN), .B(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n10616) );
  OR2_X1 U11532 ( .A1(n9525), .A2(n10616), .ZN(n9208) );
  INV_X1 U11533 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n10613) );
  OR2_X1 U11534 ( .A1(n9496), .A2(n10613), .ZN(n9207) );
  NAND4_X1 U11535 ( .A1(n9210), .A2(n9209), .A3(n9208), .A4(n9207), .ZN(n13371) );
  XNOR2_X1 U11536 ( .A(n12025), .B(n13371), .ZN(n12251) );
  INV_X1 U11537 ( .A(n13371), .ZN(n9211) );
  NAND2_X1 U11538 ( .A1(n9211), .A2(n12025), .ZN(n9212) );
  NOR2_X1 U11539 ( .A1(n9310), .A2(n9405), .ZN(n9213) );
  MUX2_X1 U11540 ( .A(n9405), .B(n9213), .S(P2_IR_REG_5__SCAN_IN), .Z(n9215)
         );
  INV_X1 U11541 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n9214) );
  NOR2_X1 U11542 ( .A1(n9215), .A2(n9226), .ZN(n9871) );
  AOI22_X1 U11543 ( .A1(n9392), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n9391), .B2(
        n9871), .ZN(n9216) );
  INV_X1 U11544 ( .A(n9476), .ZN(n9436) );
  AOI21_X1 U11545 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(P2_REG3_REG_3__SCAN_IN), 
        .A(P2_REG3_REG_5__SCAN_IN), .ZN(n9217) );
  NOR2_X1 U11546 ( .A1(n9217), .A2(n9230), .ZN(n10665) );
  NAND2_X1 U11547 ( .A1(n9436), .A2(n10665), .ZN(n9223) );
  INV_X1 U11548 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n9218) );
  OR2_X1 U11549 ( .A1(n6546), .A2(n9218), .ZN(n9222) );
  INV_X1 U11550 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n9219) );
  OR2_X1 U11551 ( .A1(n12196), .A2(n9219), .ZN(n9221) );
  INV_X1 U11552 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n10663) );
  OR2_X1 U11553 ( .A1(n9496), .A2(n10663), .ZN(n9220) );
  NAND4_X1 U11554 ( .A1(n9223), .A2(n9222), .A3(n9221), .A4(n9220), .ZN(n13370) );
  INV_X1 U11555 ( .A(n13370), .ZN(n12037) );
  AND2_X1 U11556 ( .A1(n6721), .A2(n12037), .ZN(n9224) );
  INV_X1 U11557 ( .A(n6721), .ZN(n10667) );
  NAND2_X1 U11558 ( .A1(n10667), .A2(n13370), .ZN(n9225) );
  NAND2_X1 U11559 ( .A1(n9239), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9227) );
  XNOR2_X1 U11560 ( .A(n9227), .B(P2_IR_REG_6__SCAN_IN), .ZN(n9987) );
  AOI22_X1 U11561 ( .A1(n9392), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n9391), .B2(
        n9987), .ZN(n9228) );
  NAND2_X1 U11562 ( .A1(n9229), .A2(n9228), .ZN(n12048) );
  INV_X1 U11563 ( .A(n12048), .ZN(n14974) );
  NAND2_X1 U11564 ( .A1(n12162), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n9235) );
  INV_X1 U11565 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n10850) );
  OR2_X1 U11566 ( .A1(n9496), .A2(n10850), .ZN(n9234) );
  NAND2_X1 U11567 ( .A1(n9230), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n9244) );
  OAI21_X1 U11568 ( .B1(n9230), .B2(P2_REG3_REG_6__SCAN_IN), .A(n9244), .ZN(
        n10849) );
  OR2_X1 U11569 ( .A1(n9525), .A2(n10849), .ZN(n9233) );
  INV_X1 U11570 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n9231) );
  OR2_X1 U11571 ( .A1(n6546), .A2(n9231), .ZN(n9232) );
  NAND4_X1 U11572 ( .A1(n9235), .A2(n9234), .A3(n9233), .A4(n9232), .ZN(n13369) );
  NAND2_X1 U11573 ( .A1(n14974), .A2(n13369), .ZN(n9237) );
  INV_X1 U11574 ( .A(n13369), .ZN(n9236) );
  NAND2_X1 U11575 ( .A1(n12048), .A2(n9236), .ZN(n9238) );
  INV_X1 U11576 ( .A(n12254), .ZN(n9543) );
  NAND2_X1 U11577 ( .A1(n9251), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9240) );
  XNOR2_X1 U11578 ( .A(n9240), .B(P2_IR_REG_7__SCAN_IN), .ZN(n13376) );
  AOI22_X1 U11579 ( .A1(n9392), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n9391), .B2(
        n13376), .ZN(n9241) );
  NAND2_X1 U11580 ( .A1(n9242), .A2(n9241), .ZN(n12052) );
  NAND2_X1 U11581 ( .A1(n12162), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n9250) );
  INV_X1 U11582 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n10986) );
  OR2_X1 U11583 ( .A1(n9496), .A2(n10986), .ZN(n9249) );
  AND2_X1 U11584 ( .A1(n9244), .A2(n9243), .ZN(n9245) );
  OR2_X1 U11585 ( .A1(n9245), .A2(n9262), .ZN(n10985) );
  OR2_X1 U11586 ( .A1(n9525), .A2(n10985), .ZN(n9248) );
  INV_X1 U11587 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n9246) );
  OR2_X1 U11588 ( .A1(n6546), .A2(n9246), .ZN(n9247) );
  NAND4_X1 U11589 ( .A1(n9250), .A2(n9249), .A3(n9248), .A4(n9247), .ZN(n13368) );
  INV_X1 U11590 ( .A(n13368), .ZN(n10785) );
  INV_X1 U11591 ( .A(n9251), .ZN(n9253) );
  INV_X1 U11592 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n9252) );
  NAND2_X1 U11593 ( .A1(n9253), .A2(n9252), .ZN(n9255) );
  NAND2_X1 U11594 ( .A1(n9255), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9254) );
  MUX2_X1 U11595 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9254), .S(
        P2_IR_REG_8__SCAN_IN), .Z(n9258) );
  INV_X1 U11596 ( .A(n9255), .ZN(n9257) );
  INV_X1 U11597 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n9256) );
  NAND2_X1 U11598 ( .A1(n9257), .A2(n9256), .ZN(n9283) );
  AOI22_X1 U11599 ( .A1(n9392), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n9391), .B2(
        n9991), .ZN(n9259) );
  NAND2_X1 U11600 ( .A1(n9524), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n9267) );
  INV_X1 U11601 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n9261) );
  OR2_X1 U11602 ( .A1(n12196), .A2(n9261), .ZN(n9266) );
  NAND2_X1 U11603 ( .A1(n9262), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n9275) );
  OR2_X1 U11604 ( .A1(n9262), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n9263) );
  NAND2_X1 U11605 ( .A1(n9275), .A2(n9263), .ZN(n10786) );
  OR2_X1 U11606 ( .A1(n9525), .A2(n10786), .ZN(n9265) );
  INV_X1 U11607 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n10720) );
  OR2_X1 U11608 ( .A1(n9496), .A2(n10720), .ZN(n9264) );
  NAND4_X1 U11609 ( .A1(n9267), .A2(n9266), .A3(n9265), .A4(n9264), .ZN(n13367) );
  NAND2_X1 U11610 ( .A1(n9268), .A2(n13367), .ZN(n9269) );
  NAND2_X1 U11611 ( .A1(n9283), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9270) );
  XNOR2_X1 U11612 ( .A(n9270), .B(P2_IR_REG_9__SCAN_IN), .ZN(n10110) );
  AOI22_X1 U11613 ( .A1(n9392), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n9391), .B2(
        n10110), .ZN(n9271) );
  NAND2_X1 U11614 ( .A1(n9524), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n9280) );
  INV_X1 U11615 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n9273) );
  OR2_X1 U11616 ( .A1(n12196), .A2(n9273), .ZN(n9279) );
  INV_X1 U11617 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n9274) );
  NAND2_X1 U11618 ( .A1(n9275), .A2(n9274), .ZN(n9276) );
  NAND2_X1 U11619 ( .A1(n9287), .A2(n9276), .ZN(n10940) );
  OR2_X1 U11620 ( .A1(n9525), .A2(n10940), .ZN(n9278) );
  INV_X1 U11621 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n10922) );
  OR2_X1 U11622 ( .A1(n9496), .A2(n10922), .ZN(n9277) );
  NAND4_X1 U11623 ( .A1(n9280), .A2(n9279), .A3(n9278), .A4(n9277), .ZN(n13366) );
  XNOR2_X1 U11624 ( .A(n6703), .B(n13366), .ZN(n12258) );
  NAND2_X1 U11625 ( .A1(n10918), .A2(n12258), .ZN(n9282) );
  INV_X1 U11626 ( .A(n13366), .ZN(n10787) );
  OR2_X1 U11627 ( .A1(n6703), .A2(n10787), .ZN(n9281) );
  NAND2_X1 U11628 ( .A1(n9911), .A2(n12168), .ZN(n9286) );
  NAND2_X1 U11629 ( .A1(n9284), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9296) );
  XNOR2_X1 U11630 ( .A(n9296), .B(P2_IR_REG_10__SCAN_IN), .ZN(n10269) );
  AOI22_X1 U11631 ( .A1(n9392), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n9391), 
        .B2(n10269), .ZN(n9285) );
  NAND2_X1 U11632 ( .A1(n9524), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n9292) );
  INV_X1 U11633 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n10109) );
  OR2_X1 U11634 ( .A1(n12196), .A2(n10109), .ZN(n9291) );
  INV_X1 U11635 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n10115) );
  NAND2_X1 U11636 ( .A1(n9287), .A2(n10115), .ZN(n9288) );
  NAND2_X1 U11637 ( .A1(n9303), .A2(n9288), .ZN(n11009) );
  OR2_X1 U11638 ( .A1(n9525), .A2(n11009), .ZN(n9290) );
  INV_X1 U11639 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n11010) );
  OR2_X1 U11640 ( .A1(n9496), .A2(n11010), .ZN(n9289) );
  NAND4_X1 U11641 ( .A1(n9292), .A2(n9291), .A3(n9290), .A4(n9289), .ZN(n13365) );
  NAND2_X1 U11642 ( .A1(n12075), .A2(n13365), .ZN(n9549) );
  OR2_X1 U11643 ( .A1(n12075), .A2(n13365), .ZN(n9293) );
  NAND2_X1 U11644 ( .A1(n9549), .A2(n9293), .ZN(n12260) );
  INV_X1 U11645 ( .A(n13365), .ZN(n12077) );
  OR2_X1 U11646 ( .A1(n12075), .A2(n12077), .ZN(n9294) );
  NAND2_X1 U11647 ( .A1(n10068), .A2(n12168), .ZN(n9300) );
  NAND2_X1 U11648 ( .A1(n9296), .A2(n9295), .ZN(n9297) );
  NAND2_X1 U11649 ( .A1(n9297), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9298) );
  XNOR2_X1 U11650 ( .A(n9298), .B(P2_IR_REG_11__SCAN_IN), .ZN(n11089) );
  AOI22_X1 U11651 ( .A1(n9392), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n9391), 
        .B2(n11089), .ZN(n9299) );
  NAND2_X1 U11652 ( .A1(n12162), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n9307) );
  INV_X1 U11653 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n9301) );
  OR2_X1 U11654 ( .A1(n6546), .A2(n9301), .ZN(n9306) );
  INV_X1 U11655 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n9302) );
  OR2_X1 U11656 ( .A1(n7540), .A2(n9317), .ZN(n11270) );
  OR2_X1 U11657 ( .A1(n9525), .A2(n11270), .ZN(n9305) );
  INV_X1 U11658 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n11083) );
  OR2_X1 U11659 ( .A1(n9496), .A2(n11083), .ZN(n9304) );
  NAND4_X1 U11660 ( .A1(n9307), .A2(n9306), .A3(n9305), .A4(n9304), .ZN(n13364) );
  INV_X1 U11661 ( .A(n13364), .ZN(n10995) );
  XNOR2_X1 U11662 ( .A(n12081), .B(n10995), .ZN(n12262) );
  INV_X1 U11663 ( .A(n12262), .ZN(n9308) );
  NAND2_X1 U11664 ( .A1(n12081), .A2(n10995), .ZN(n9309) );
  NAND2_X1 U11665 ( .A1(n10082), .A2(n12168), .ZN(n9316) );
  NAND2_X1 U11666 ( .A1(n9311), .A2(n9310), .ZN(n9313) );
  NAND2_X1 U11667 ( .A1(n9313), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9312) );
  MUX2_X1 U11668 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9312), .S(
        P2_IR_REG_12__SCAN_IN), .Z(n9314) );
  OR2_X1 U11669 ( .A1(n9313), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n9336) );
  AND2_X1 U11670 ( .A1(n9314), .A2(n9336), .ZN(n14857) );
  AOI22_X1 U11671 ( .A1(n9392), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n9391), 
        .B2(n14857), .ZN(n9315) );
  NAND2_X1 U11672 ( .A1(n9524), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n9322) );
  INV_X1 U11673 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n11093) );
  OR2_X1 U11674 ( .A1(n12196), .A2(n11093), .ZN(n9321) );
  OR2_X1 U11675 ( .A1(n9317), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n9318) );
  NAND2_X1 U11676 ( .A1(n9345), .A2(n9318), .ZN(n11409) );
  OR2_X1 U11677 ( .A1(n9476), .A2(n11409), .ZN(n9320) );
  INV_X1 U11678 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n11309) );
  OR2_X1 U11679 ( .A1(n9496), .A2(n11309), .ZN(n9319) );
  NAND4_X1 U11680 ( .A1(n9322), .A2(n9321), .A3(n9320), .A4(n9319), .ZN(n13363) );
  XNOR2_X1 U11681 ( .A(n12087), .B(n11428), .ZN(n12263) );
  NAND2_X1 U11682 ( .A1(n11306), .A2(n9323), .ZN(n11305) );
  OR2_X1 U11683 ( .A1(n12087), .A2(n11428), .ZN(n9324) );
  NAND2_X1 U11684 ( .A1(n11305), .A2(n9324), .ZN(n11415) );
  NAND2_X1 U11685 ( .A1(n10189), .A2(n12168), .ZN(n9327) );
  NAND2_X1 U11686 ( .A1(n9336), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9325) );
  XNOR2_X1 U11687 ( .A(n9325), .B(P2_IR_REG_13__SCAN_IN), .ZN(n14878) );
  AOI22_X1 U11688 ( .A1(n9392), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n9391), 
        .B2(n14878), .ZN(n9326) );
  NAND2_X1 U11689 ( .A1(n12162), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n9333) );
  INV_X1 U11690 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n9343) );
  XNOR2_X1 U11691 ( .A(n9345), .B(n9343), .ZN(n11429) );
  OR2_X1 U11692 ( .A1(n9525), .A2(n11429), .ZN(n9332) );
  INV_X1 U11693 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n9328) );
  OR2_X1 U11694 ( .A1(n9496), .A2(n9328), .ZN(n9331) );
  INV_X1 U11695 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n9329) );
  OR2_X1 U11696 ( .A1(n6546), .A2(n9329), .ZN(n9330) );
  NAND4_X1 U11697 ( .A1(n9333), .A2(n9332), .A3(n9331), .A4(n9330), .ZN(n13362) );
  INV_X1 U11698 ( .A(n13362), .ZN(n12094) );
  XNOR2_X1 U11699 ( .A(n12092), .B(n12094), .ZN(n12264) );
  INV_X1 U11700 ( .A(n12264), .ZN(n11414) );
  NAND2_X1 U11701 ( .A1(n11415), .A2(n11414), .ZN(n9335) );
  OR2_X1 U11702 ( .A1(n12092), .A2(n12094), .ZN(n9334) );
  NAND2_X1 U11703 ( .A1(n10452), .A2(n12168), .ZN(n9340) );
  OAI21_X1 U11704 ( .B1(n9336), .B2(P2_IR_REG_13__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9337) );
  MUX2_X1 U11705 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9337), .S(
        P2_IR_REG_14__SCAN_IN), .Z(n9338) );
  NAND2_X1 U11706 ( .A1(n9338), .A2(n9351), .ZN(n11088) );
  INV_X1 U11707 ( .A(n11088), .ZN(n13402) );
  AOI22_X1 U11708 ( .A1(n9392), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n9391), 
        .B2(n13402), .ZN(n9339) );
  INV_X1 U11710 ( .A(n12105), .ZN(n14650) );
  NAND2_X1 U11711 ( .A1(n9524), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n9350) );
  INV_X1 U11712 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n9341) );
  OR2_X1 U11713 ( .A1(n12196), .A2(n9341), .ZN(n9349) );
  INV_X1 U11714 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n9342) );
  OAI21_X1 U11715 ( .B1(n9345), .B2(n9343), .A(n9342), .ZN(n9346) );
  NAND2_X1 U11716 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_REG3_REG_14__SCAN_IN), 
        .ZN(n9344) );
  NAND2_X1 U11717 ( .A1(n9346), .A2(n9355), .ZN(n11668) );
  OR2_X1 U11718 ( .A1(n9525), .A2(n11668), .ZN(n9348) );
  INV_X1 U11719 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n11572) );
  OR2_X1 U11720 ( .A1(n9496), .A2(n11572), .ZN(n9347) );
  NAND4_X1 U11721 ( .A1(n9350), .A2(n9349), .A3(n9348), .A4(n9347), .ZN(n13361) );
  INV_X1 U11722 ( .A(n13361), .ZN(n11430) );
  NAND2_X1 U11723 ( .A1(n10557), .A2(n12168), .ZN(n9354) );
  NAND2_X1 U11724 ( .A1(n9351), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9352) );
  XNOR2_X1 U11725 ( .A(n9352), .B(n7155), .ZN(n13404) );
  INV_X1 U11726 ( .A(n13404), .ZN(n14888) );
  AOI22_X1 U11727 ( .A1(n9392), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n9391), 
        .B2(n14888), .ZN(n9353) );
  INV_X1 U11728 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n11701) );
  AND2_X1 U11729 ( .A1(n9355), .A2(n11701), .ZN(n9356) );
  NOR2_X1 U11730 ( .A1(n9366), .A2(n9356), .ZN(n11705) );
  NAND2_X1 U11731 ( .A1(n9436), .A2(n11705), .ZN(n9361) );
  INV_X1 U11732 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n14884) );
  OR2_X1 U11733 ( .A1(n12196), .A2(n14884), .ZN(n9360) );
  INV_X1 U11734 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n11768) );
  OR2_X1 U11735 ( .A1(n6546), .A2(n11768), .ZN(n9359) );
  INV_X1 U11736 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n9357) );
  OR2_X1 U11737 ( .A1(n9496), .A2(n9357), .ZN(n9358) );
  NAND4_X1 U11738 ( .A1(n9361), .A2(n9360), .A3(n9359), .A4(n9358), .ZN(n13360) );
  XNOR2_X1 U11739 ( .A(n12110), .B(n13360), .ZN(n12270) );
  INV_X1 U11740 ( .A(n12270), .ZN(n11687) );
  INV_X1 U11741 ( .A(n13360), .ZN(n12112) );
  OR2_X1 U11742 ( .A1(n12110), .A2(n12112), .ZN(n9362) );
  OAI21_X1 U11743 ( .B1(n11688), .B2(n11687), .A(n9362), .ZN(n11806) );
  NAND2_X1 U11744 ( .A1(n10420), .A2(n12168), .ZN(n9365) );
  NAND2_X1 U11745 ( .A1(n7154), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9363) );
  XNOR2_X1 U11746 ( .A(n9363), .B(P2_IR_REG_16__SCAN_IN), .ZN(n14900) );
  AOI22_X1 U11747 ( .A1(n9392), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n9391), 
        .B2(n14900), .ZN(n9364) );
  NOR2_X1 U11748 ( .A1(n9366), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n9367) );
  OR2_X1 U11749 ( .A1(n9380), .A2(n9367), .ZN(n11840) );
  INV_X1 U11750 ( .A(n9496), .ZN(n12161) );
  NAND2_X1 U11751 ( .A1(n12161), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n9368) );
  OAI21_X1 U11752 ( .B1(n11840), .B2(n9525), .A(n9368), .ZN(n9372) );
  INV_X1 U11753 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n9370) );
  NAND2_X1 U11754 ( .A1(n12162), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n9369) );
  OAI21_X1 U11755 ( .B1(n6546), .B2(n9370), .A(n9369), .ZN(n9371) );
  OR2_X1 U11756 ( .A1(n9372), .A2(n9371), .ZN(n13359) );
  INV_X1 U11757 ( .A(n13359), .ZN(n9373) );
  XNOR2_X1 U11758 ( .A(n13726), .B(n9373), .ZN(n12266) );
  NAND2_X1 U11759 ( .A1(n11806), .A2(n11805), .ZN(n11804) );
  OR2_X1 U11760 ( .A1(n13726), .A2(n9373), .ZN(n9374) );
  NAND2_X1 U11761 ( .A1(n11804), .A2(n9374), .ZN(n11846) );
  NAND2_X1 U11762 ( .A1(n10456), .A2(n12168), .ZN(n9379) );
  INV_X1 U11763 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n9375) );
  OR2_X1 U11764 ( .A1(n9389), .A2(n9405), .ZN(n9377) );
  XNOR2_X1 U11765 ( .A(n9377), .B(P2_IR_REG_17__SCAN_IN), .ZN(n14913) );
  AOI22_X1 U11766 ( .A1(n9392), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n9391), 
        .B2(n14913), .ZN(n9378) );
  OR2_X1 U11767 ( .A1(n9380), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n9381) );
  NAND2_X1 U11768 ( .A1(n9415), .A2(n9381), .ZN(n11866) );
  NAND2_X1 U11769 ( .A1(n9524), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n9383) );
  NAND2_X1 U11770 ( .A1(n12162), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n9382) );
  AND2_X1 U11771 ( .A1(n9383), .A2(n9382), .ZN(n9385) );
  NAND2_X1 U11772 ( .A1(n12161), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n9384) );
  OAI211_X1 U11773 ( .C1(n11866), .C2(n9525), .A(n9385), .B(n9384), .ZN(n13358) );
  INV_X1 U11774 ( .A(n13358), .ZN(n13628) );
  NAND2_X1 U11775 ( .A1(n12125), .A2(n13628), .ZN(n9386) );
  OR2_X1 U11776 ( .A1(n12125), .A2(n13628), .ZN(n9387) );
  NAND2_X1 U11777 ( .A1(n10830), .A2(n12168), .ZN(n9394) );
  INV_X1 U11778 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n9388) );
  NAND2_X1 U11779 ( .A1(n9404), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9390) );
  XNOR2_X1 U11780 ( .A(n9390), .B(n7150), .ZN(n14920) );
  INV_X1 U11781 ( .A(n14920), .ZN(n13397) );
  AOI22_X1 U11782 ( .A1(n9392), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n9391), 
        .B2(n13397), .ZN(n9393) );
  XNOR2_X1 U11783 ( .A(n9415), .B(P2_REG3_REG_18__SCAN_IN), .ZN(n13634) );
  NAND2_X1 U11784 ( .A1(n13634), .A2(n9436), .ZN(n9400) );
  INV_X1 U11785 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n14924) );
  NAND2_X1 U11786 ( .A1(n9524), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n9397) );
  INV_X1 U11787 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n9395) );
  OR2_X1 U11788 ( .A1(n9496), .A2(n9395), .ZN(n9396) );
  OAI211_X1 U11789 ( .C1(n12196), .C2(n14924), .A(n9397), .B(n9396), .ZN(n9398) );
  INV_X1 U11790 ( .A(n9398), .ZN(n9399) );
  NAND2_X1 U11791 ( .A1(n9400), .A2(n9399), .ZN(n13357) );
  INV_X1 U11792 ( .A(n13357), .ZN(n12134) );
  NAND2_X1 U11793 ( .A1(n13711), .A2(n12134), .ZN(n9401) );
  NAND2_X1 U11794 ( .A1(n9402), .A2(n9401), .ZN(n13598) );
  NAND2_X1 U11795 ( .A1(n10991), .A2(n12168), .ZN(n9411) );
  OR2_X1 U11796 ( .A1(n9516), .A2(n9405), .ZN(n9406) );
  MUX2_X1 U11797 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9406), .S(
        P2_IR_REG_19__SCAN_IN), .Z(n9408) );
  INV_X1 U11798 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n9407) );
  NAND2_X1 U11799 ( .A1(n9516), .A2(n9407), .ZN(n9520) );
  INV_X2 U11800 ( .A(n7536), .ZN(n12613) );
  OAI22_X1 U11801 ( .A1(n9502), .A2(n12615), .B1(n12613), .B2(n9841), .ZN(
        n9409) );
  INV_X1 U11802 ( .A(n9409), .ZN(n9410) );
  INV_X1 U11803 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n9419) );
  INV_X1 U11804 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n9413) );
  INV_X1 U11805 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n9412) );
  OAI21_X1 U11806 ( .B1(n9415), .B2(n9413), .A(n9412), .ZN(n9416) );
  NAND2_X1 U11807 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(P2_REG3_REG_19__SCAN_IN), 
        .ZN(n9414) );
  NAND2_X1 U11808 ( .A1(n9416), .A2(n9425), .ZN(n13607) );
  OR2_X1 U11809 ( .A1(n13607), .A2(n9476), .ZN(n9418) );
  AOI22_X1 U11810 ( .A1(n12162), .A2(P2_REG1_REG_19__SCAN_IN), .B1(n12161), 
        .B2(P2_REG2_REG_19__SCAN_IN), .ZN(n9417) );
  OAI211_X1 U11811 ( .C1(n6546), .C2(n9419), .A(n9418), .B(n9417), .ZN(n13625)
         );
  INV_X1 U11812 ( .A(n13625), .ZN(n9420) );
  XNOR2_X1 U11813 ( .A(n13708), .B(n9420), .ZN(n13597) );
  INV_X1 U11814 ( .A(n13597), .ZN(n13595) );
  NAND2_X1 U11815 ( .A1(n13598), .A2(n13595), .ZN(n9422) );
  NAND2_X1 U11816 ( .A1(n13708), .A2(n9420), .ZN(n9421) );
  NAND2_X1 U11817 ( .A1(n9422), .A2(n9421), .ZN(n13585) );
  NAND2_X1 U11818 ( .A1(n11033), .A2(n12168), .ZN(n9424) );
  OR2_X1 U11819 ( .A1(n9502), .A2(n15400), .ZN(n9423) );
  INV_X1 U11820 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n13317) );
  AND2_X1 U11821 ( .A1(n9425), .A2(n13317), .ZN(n9426) );
  OR2_X1 U11822 ( .A1(n9426), .A2(n9434), .ZN(n13316) );
  INV_X1 U11823 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n15465) );
  NAND2_X1 U11824 ( .A1(n12161), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n9428) );
  NAND2_X1 U11825 ( .A1(n12162), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n9427) );
  OAI211_X1 U11826 ( .C1(n6546), .C2(n15465), .A(n9428), .B(n9427), .ZN(n9429)
         );
  INV_X1 U11827 ( .A(n9429), .ZN(n9430) );
  OAI21_X1 U11828 ( .B1(n13316), .B2(n9525), .A(n9430), .ZN(n13356) );
  INV_X1 U11829 ( .A(n13356), .ZN(n12143) );
  XNOR2_X1 U11830 ( .A(n13703), .B(n12143), .ZN(n13584) );
  INV_X1 U11831 ( .A(n13584), .ZN(n13582) );
  NAND2_X1 U11832 ( .A1(n13703), .A2(n12143), .ZN(n9431) );
  NAND2_X1 U11833 ( .A1(n11134), .A2(n12168), .ZN(n9433) );
  OR2_X1 U11834 ( .A1(n9502), .A2(n11135), .ZN(n9432) );
  OR2_X1 U11835 ( .A1(n9434), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n9435) );
  NAND2_X1 U11836 ( .A1(n9434), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n9447) );
  AND2_X1 U11837 ( .A1(n9435), .A2(n9447), .ZN(n13575) );
  NAND2_X1 U11838 ( .A1(n13575), .A2(n9436), .ZN(n9441) );
  INV_X1 U11839 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n13753) );
  NAND2_X1 U11840 ( .A1(n12162), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n9438) );
  NAND2_X1 U11841 ( .A1(n12161), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n9437) );
  OAI211_X1 U11842 ( .C1(n6546), .C2(n13753), .A(n9438), .B(n9437), .ZN(n9439)
         );
  INV_X1 U11843 ( .A(n9439), .ZN(n9440) );
  INV_X1 U11844 ( .A(n13550), .ZN(n13355) );
  NOR2_X1 U11845 ( .A1(n13755), .A2(n13355), .ZN(n9442) );
  XNOR2_X1 U11846 ( .A(n8042), .B(n9443), .ZN(n11167) );
  NAND2_X1 U11847 ( .A1(n11167), .A2(n12168), .ZN(n9445) );
  OR2_X1 U11848 ( .A1(n9502), .A2(n15312), .ZN(n9444) );
  NAND2_X1 U11849 ( .A1(n12162), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n9453) );
  INV_X1 U11850 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n9446) );
  OR2_X1 U11851 ( .A1(n9496), .A2(n9446), .ZN(n9452) );
  OAI21_X1 U11852 ( .B1(P2_REG3_REG_22__SCAN_IN), .B2(n9448), .A(n9456), .ZN(
        n13556) );
  OR2_X1 U11853 ( .A1(n9476), .A2(n13556), .ZN(n9451) );
  INV_X1 U11854 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n9449) );
  OR2_X1 U11855 ( .A1(n6546), .A2(n9449), .ZN(n9450) );
  NAND4_X1 U11856 ( .A1(n9453), .A2(n9452), .A3(n9451), .A4(n9450), .ZN(n13532) );
  XNOR2_X1 U11857 ( .A(n13690), .B(n13532), .ZN(n12275) );
  INV_X1 U11858 ( .A(n13532), .ZN(n13264) );
  NAND2_X1 U11859 ( .A1(n11480), .A2(n12168), .ZN(n9455) );
  OR2_X1 U11860 ( .A1(n9502), .A2(n15252), .ZN(n9454) );
  NAND2_X1 U11861 ( .A1(n9524), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n9461) );
  INV_X1 U11862 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n15327) );
  OR2_X1 U11863 ( .A1(n12196), .A2(n15327), .ZN(n9460) );
  INV_X1 U11864 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n13541) );
  OR2_X1 U11865 ( .A1(n9496), .A2(n13541), .ZN(n9459) );
  INV_X1 U11866 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n13263) );
  AOI21_X1 U11867 ( .B1(n9456), .B2(n13263), .A(n9466), .ZN(n9457) );
  INV_X1 U11868 ( .A(n9457), .ZN(n13536) );
  OR2_X1 U11869 ( .A1(n9525), .A2(n13536), .ZN(n9458) );
  AND2_X1 U11870 ( .A1(n13542), .A2(n13354), .ZN(n9462) );
  NAND2_X1 U11871 ( .A1(n11613), .A2(n12168), .ZN(n9464) );
  OR2_X1 U11872 ( .A1(n9502), .A2(n11615), .ZN(n9463) );
  NAND2_X1 U11873 ( .A1(n12162), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n9470) );
  INV_X1 U11874 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n9465) );
  OR2_X1 U11875 ( .A1(n6546), .A2(n9465), .ZN(n9469) );
  NAND2_X1 U11876 ( .A1(n9466), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n9473) );
  OAI21_X1 U11877 ( .B1(P2_REG3_REG_24__SCAN_IN), .B2(n9466), .A(n9473), .ZN(
        n13521) );
  OR2_X1 U11878 ( .A1(n9525), .A2(n13521), .ZN(n9468) );
  INV_X1 U11879 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n13522) );
  OR2_X1 U11880 ( .A1(n9496), .A2(n13522), .ZN(n9467) );
  NAND4_X1 U11881 ( .A1(n9470), .A2(n9469), .A3(n9468), .A4(n9467), .ZN(n13533) );
  XNOR2_X1 U11882 ( .A(n13681), .B(n13533), .ZN(n13509) );
  INV_X1 U11883 ( .A(n13533), .ZN(n13299) );
  NAND2_X1 U11884 ( .A1(n11649), .A2(n12168), .ZN(n9472) );
  OR2_X1 U11885 ( .A1(n9502), .A2(n11651), .ZN(n9471) );
  NAND2_X1 U11886 ( .A1(n9524), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n9480) );
  INV_X1 U11887 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n13678) );
  OR2_X1 U11888 ( .A1(n12196), .A2(n13678), .ZN(n9479) );
  INV_X1 U11889 ( .A(n9473), .ZN(n9475) );
  INV_X1 U11890 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n13298) );
  INV_X1 U11891 ( .A(n9486), .ZN(n9474) );
  OAI21_X1 U11892 ( .B1(P2_REG3_REG_25__SCAN_IN), .B2(n9475), .A(n9474), .ZN(
        n13501) );
  OR2_X1 U11893 ( .A1(n9476), .A2(n13501), .ZN(n9478) );
  INV_X1 U11894 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n13502) );
  OR2_X1 U11895 ( .A1(n9496), .A2(n13502), .ZN(n9477) );
  NAND4_X1 U11896 ( .A1(n9480), .A2(n9479), .A3(n9478), .A4(n9477), .ZN(n13353) );
  XNOR2_X1 U11897 ( .A(n13503), .B(n13353), .ZN(n13493) );
  INV_X1 U11898 ( .A(n13353), .ZN(n9481) );
  NAND2_X1 U11899 ( .A1(n13503), .A2(n9481), .ZN(n9482) );
  NAND2_X1 U11900 ( .A1(n9483), .A2(n9482), .ZN(n13476) );
  NAND2_X1 U11901 ( .A1(n11816), .A2(n12168), .ZN(n9485) );
  OR2_X1 U11902 ( .A1(n9502), .A2(n11817), .ZN(n9484) );
  NAND2_X1 U11903 ( .A1(n12161), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n9490) );
  INV_X1 U11904 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n15435) );
  OR2_X1 U11905 ( .A1(n6546), .A2(n15435), .ZN(n9489) );
  INV_X1 U11906 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n15486) );
  OR2_X1 U11907 ( .A1(n12196), .A2(n15486), .ZN(n9488) );
  NAND2_X1 U11908 ( .A1(n9486), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n9494) );
  OAI21_X1 U11909 ( .B1(P2_REG3_REG_26__SCAN_IN), .B2(n9486), .A(n9494), .ZN(
        n13482) );
  OR2_X1 U11910 ( .A1(n9525), .A2(n13482), .ZN(n9487) );
  NAND4_X1 U11911 ( .A1(n9490), .A2(n9489), .A3(n9488), .A4(n9487), .ZN(n13495) );
  INV_X1 U11912 ( .A(n13495), .ZN(n13300) );
  OR2_X1 U11913 ( .A1(n13670), .A2(n13300), .ZN(n12245) );
  NAND2_X1 U11914 ( .A1(n13476), .A2(n12245), .ZN(n9491) );
  NAND2_X1 U11915 ( .A1(n13670), .A2(n13300), .ZN(n12244) );
  OR2_X1 U11916 ( .A1(n9502), .A2(n12312), .ZN(n9492) );
  NAND2_X1 U11917 ( .A1(n9524), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n9500) );
  INV_X1 U11918 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n13667) );
  OR2_X1 U11919 ( .A1(n12196), .A2(n13667), .ZN(n9499) );
  INV_X1 U11920 ( .A(n9494), .ZN(n9495) );
  INV_X1 U11921 ( .A(n9506), .ZN(n9508) );
  OAI21_X1 U11922 ( .B1(P2_REG3_REG_27__SCAN_IN), .B2(n9495), .A(n9508), .ZN(
        n13466) );
  OR2_X1 U11923 ( .A1(n9525), .A2(n13466), .ZN(n9498) );
  INV_X1 U11924 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n13467) );
  OR2_X1 U11925 ( .A1(n9496), .A2(n13467), .ZN(n9497) );
  NAND4_X1 U11926 ( .A1(n9500), .A2(n9499), .A3(n9498), .A4(n9497), .ZN(n13352) );
  INV_X1 U11927 ( .A(n13352), .ZN(n9501) );
  NAND2_X1 U11928 ( .A1(n13776), .A2(n12168), .ZN(n9504) );
  OR2_X1 U11929 ( .A1(n9502), .A2(n13779), .ZN(n9503) );
  NAND2_X1 U11930 ( .A1(n9524), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n9513) );
  INV_X1 U11931 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n9505) );
  OR2_X1 U11932 ( .A1(n12196), .A2(n9505), .ZN(n9512) );
  NAND2_X1 U11933 ( .A1(n9506), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n13444) );
  INV_X1 U11934 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n9507) );
  NAND2_X1 U11935 ( .A1(n9508), .A2(n9507), .ZN(n9509) );
  NAND2_X1 U11936 ( .A1(n13444), .A2(n9509), .ZN(n13451) );
  OR2_X1 U11937 ( .A1(n9525), .A2(n13451), .ZN(n9511) );
  INV_X1 U11938 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n13454) );
  OR2_X1 U11939 ( .A1(n9496), .A2(n13454), .ZN(n9510) );
  NAND4_X1 U11940 ( .A1(n9513), .A2(n9512), .A3(n9511), .A4(n9510), .ZN(n13463) );
  NAND2_X1 U11941 ( .A1(n13287), .A2(n13463), .ZN(n13430) );
  NAND2_X1 U11942 ( .A1(n9578), .A2(n7536), .ZN(n9523) );
  NAND2_X1 U11943 ( .A1(n9518), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9519) );
  XNOR2_X1 U11944 ( .A(n9519), .B(P2_IR_REG_21__SCAN_IN), .ZN(n10529) );
  INV_X1 U11945 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n9521) );
  XNOR2_X2 U11946 ( .A(n9522), .B(n9521), .ZN(n9579) );
  INV_X1 U11947 ( .A(n9579), .ZN(n12246) );
  NAND2_X1 U11948 ( .A1(n10529), .A2(n12246), .ZN(n12288) );
  AND2_X2 U11949 ( .A1(n10015), .A2(n9852), .ZN(n13496) );
  NAND2_X1 U11950 ( .A1(n9524), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n9530) );
  NAND2_X1 U11951 ( .A1(n12162), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n9529) );
  OR2_X1 U11952 ( .A1(n9525), .A2(n13444), .ZN(n9528) );
  INV_X1 U11953 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n9526) );
  OR2_X1 U11954 ( .A1(n9496), .A2(n9526), .ZN(n9527) );
  NAND4_X1 U11955 ( .A1(n9530), .A2(n9529), .A3(n9528), .A4(n9527), .ZN(n13351) );
  NAND2_X1 U11956 ( .A1(n13496), .A2(n13351), .ZN(n9533) );
  INV_X1 U11957 ( .A(n9852), .ZN(n9531) );
  NAND2_X1 U11958 ( .A1(n10015), .A2(n9531), .ZN(n13627) );
  INV_X1 U11959 ( .A(n13627), .ZN(n13462) );
  NAND2_X1 U11960 ( .A1(n13462), .A2(n13352), .ZN(n9532) );
  NAND2_X1 U11961 ( .A1(n9533), .A2(n9532), .ZN(n13284) );
  INV_X1 U11962 ( .A(n13284), .ZN(n9534) );
  NAND2_X1 U11963 ( .A1(n13375), .A2(n12002), .ZN(n10532) );
  INV_X1 U11964 ( .A(n10532), .ZN(n9536) );
  OR2_X1 U11965 ( .A1(n13374), .A2(n14934), .ZN(n9537) );
  OR2_X1 U11966 ( .A1(n13373), .A2(n12016), .ZN(n9538) );
  NAND2_X1 U11967 ( .A1(n10072), .A2(n9538), .ZN(n10143) );
  OR2_X1 U11968 ( .A1(n13372), .A2(n12021), .ZN(n9539) );
  NAND2_X1 U11969 ( .A1(n10142), .A2(n9539), .ZN(n10237) );
  INV_X1 U11970 ( .A(n12251), .ZN(n10240) );
  OR2_X1 U11971 ( .A1(n12025), .A2(n13371), .ZN(n9540) );
  NAND2_X1 U11972 ( .A1(n6721), .A2(n13370), .ZN(n9541) );
  NAND2_X1 U11973 ( .A1(n10667), .A2(n12037), .ZN(n9542) );
  NAND2_X1 U11974 ( .A1(n10855), .A2(n9543), .ZN(n9545) );
  OR2_X1 U11975 ( .A1(n12048), .A2(n13369), .ZN(n9544) );
  NAND2_X1 U11976 ( .A1(n9545), .A2(n9544), .ZN(n10982) );
  XNOR2_X1 U11977 ( .A(n12052), .B(n10785), .ZN(n12256) );
  OR2_X1 U11978 ( .A1(n12052), .A2(n13368), .ZN(n9546) );
  XNOR2_X1 U11979 ( .A(n12060), .B(n13367), .ZN(n12257) );
  NAND2_X1 U11980 ( .A1(n12060), .A2(n13367), .ZN(n9547) );
  NAND2_X1 U11981 ( .A1(n10715), .A2(n9547), .ZN(n10914) );
  INV_X1 U11982 ( .A(n12258), .ZN(n10917) );
  NAND2_X1 U11983 ( .A1(n10914), .A2(n10917), .ZN(n10916) );
  NAND2_X1 U11984 ( .A1(n6703), .A2(n13366), .ZN(n9548) );
  NAND2_X1 U11985 ( .A1(n10916), .A2(n9548), .ZN(n11001) );
  INV_X1 U11986 ( .A(n12260), .ZN(n11004) );
  NAND2_X1 U11987 ( .A1(n11001), .A2(n11004), .ZN(n11003) );
  OR2_X1 U11988 ( .A1(n12081), .A2(n13364), .ZN(n9550) );
  NAND2_X1 U11989 ( .A1(n12081), .A2(n13364), .ZN(n9551) );
  OR2_X1 U11990 ( .A1(n12087), .A2(n13363), .ZN(n9552) );
  NAND2_X1 U11991 ( .A1(n11302), .A2(n9552), .ZN(n11417) );
  NAND2_X1 U11992 ( .A1(n12092), .A2(n13362), .ZN(n9553) );
  NAND2_X1 U11993 ( .A1(n11417), .A2(n9553), .ZN(n9555) );
  OR2_X1 U11994 ( .A1(n12092), .A2(n13362), .ZN(n9554) );
  NAND2_X1 U11995 ( .A1(n9555), .A2(n9554), .ZN(n11570) );
  NOR2_X1 U11996 ( .A1(n12105), .A2(n13361), .ZN(n9556) );
  NAND2_X1 U11997 ( .A1(n12105), .A2(n13361), .ZN(n9557) );
  OR2_X1 U11998 ( .A1(n12110), .A2(n13360), .ZN(n9558) );
  NAND2_X1 U11999 ( .A1(n13726), .A2(n13359), .ZN(n9559) );
  XNOR2_X1 U12000 ( .A(n12125), .B(n13358), .ZN(n12267) );
  INV_X1 U12001 ( .A(n12267), .ZN(n9560) );
  NAND2_X1 U12002 ( .A1(n11845), .A2(n9560), .ZN(n9562) );
  NAND2_X1 U12003 ( .A1(n12125), .A2(n13358), .ZN(n9561) );
  XNOR2_X1 U12004 ( .A(n13711), .B(n12134), .ZN(n13616) );
  INV_X1 U12005 ( .A(n13616), .ZN(n13620) );
  OR2_X1 U12006 ( .A1(n13711), .A2(n13357), .ZN(n9563) );
  NAND2_X1 U12007 ( .A1(n13708), .A2(n13625), .ZN(n9564) );
  NAND2_X1 U12008 ( .A1(n13596), .A2(n9564), .ZN(n9566) );
  OR2_X1 U12009 ( .A1(n13708), .A2(n13625), .ZN(n9565) );
  NAND2_X1 U12010 ( .A1(n9566), .A2(n9565), .ZN(n13583) );
  XNOR2_X1 U12011 ( .A(n13574), .B(n13550), .ZN(n13565) );
  INV_X1 U12012 ( .A(n13565), .ZN(n13569) );
  NAND2_X1 U12013 ( .A1(n13755), .A2(n13550), .ZN(n9567) );
  NAND2_X1 U12014 ( .A1(n13690), .A2(n13532), .ZN(n9568) );
  NAND2_X1 U12015 ( .A1(n13529), .A2(n12274), .ZN(n9569) );
  NAND2_X1 U12016 ( .A1(n13686), .A2(n13354), .ZN(n12273) );
  NAND2_X1 U12017 ( .A1(n9569), .A2(n12273), .ZN(n13512) );
  INV_X1 U12018 ( .A(n13509), .ZN(n13511) );
  NAND2_X1 U12019 ( .A1(n13512), .A2(n13511), .ZN(n13514) );
  NAND2_X1 U12020 ( .A1(n13681), .A2(n13533), .ZN(n9570) );
  OR2_X1 U12021 ( .A1(n13503), .A2(n13353), .ZN(n9571) );
  NAND2_X1 U12022 ( .A1(n13491), .A2(n9571), .ZN(n9573) );
  NAND2_X1 U12023 ( .A1(n13503), .A2(n13353), .ZN(n9572) );
  AND2_X1 U12024 ( .A1(n13670), .A2(n13495), .ZN(n9575) );
  OR2_X1 U12025 ( .A1(n13670), .A2(n13495), .ZN(n9574) );
  NAND2_X1 U12026 ( .A1(n9577), .A2(n9576), .ZN(n13431) );
  OAI21_X1 U12027 ( .B1(n9577), .B2(n9576), .A(n13431), .ZN(n13459) );
  INV_X1 U12028 ( .A(n9578), .ZN(n12000) );
  NAND2_X1 U12029 ( .A1(n12000), .A2(n10530), .ZN(n14970) );
  INV_X1 U12030 ( .A(n12075), .ZN(n15000) );
  INV_X1 U12031 ( .A(n12052), .ZN(n14981) );
  OR2_X1 U12032 ( .A1(n14934), .A2(n12002), .ZN(n10074) );
  INV_X1 U12033 ( .A(n12125), .ZN(n13765) );
  NAND2_X1 U12034 ( .A1(n13588), .A2(n13755), .ZN(n13571) );
  NAND2_X1 U12035 ( .A1(n13555), .A2(n13542), .ZN(n13538) );
  NOR2_X2 U12036 ( .A1(n13518), .A2(n13503), .ZN(n13479) );
  INV_X2 U12037 ( .A(n10019), .ZN(n10533) );
  OAI211_X1 U12038 ( .C1(n13658), .C2(n6582), .A(n13603), .B(n13441), .ZN(
        n13453) );
  INV_X1 U12039 ( .A(n9583), .ZN(n9584) );
  NAND2_X1 U12040 ( .A1(n9584), .A2(n9600), .ZN(n9588) );
  INV_X1 U12041 ( .A(n9588), .ZN(n9585) );
  NAND2_X1 U12042 ( .A1(n9585), .A2(n9589), .ZN(n9591) );
  NAND2_X1 U12043 ( .A1(n9591), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9586) );
  MUX2_X1 U12044 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9586), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n9587) );
  NAND2_X1 U12045 ( .A1(n9587), .A2(n9594), .ZN(n11650) );
  NAND2_X1 U12046 ( .A1(n9588), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9590) );
  MUX2_X1 U12047 ( .A(n9590), .B(P2_IR_REG_31__SCAN_IN), .S(n9589), .Z(n9592)
         );
  NAND2_X1 U12048 ( .A1(n9592), .A2(n9591), .ZN(n11614) );
  XNOR2_X1 U12049 ( .A(n11614), .B(P2_B_REG_SCAN_IN), .ZN(n9593) );
  AND2_X1 U12050 ( .A1(n11650), .A2(n9593), .ZN(n9599) );
  NAND2_X1 U12051 ( .A1(n9594), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9596) );
  MUX2_X1 U12052 ( .A(n9596), .B(P2_IR_REG_31__SCAN_IN), .S(n9595), .Z(n9598)
         );
  NAND2_X1 U12053 ( .A1(n9598), .A2(n9597), .ZN(n11818) );
  NOR2_X1 U12054 ( .A1(n9599), .A2(n11818), .ZN(n14948) );
  INV_X1 U12055 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n14957) );
  AOI22_X1 U12056 ( .A1(n14948), .A2(n14957), .B1(n11818), .B2(n11650), .ZN(
        n10004) );
  NAND2_X1 U12057 ( .A1(n9583), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9601) );
  XNOR2_X1 U12058 ( .A(n9601), .B(n9600), .ZN(n11481) );
  NOR3_X1 U12059 ( .A1(n11818), .A2(n11650), .A3(n11614), .ZN(n9751) );
  INV_X1 U12060 ( .A(n9751), .ZN(n10006) );
  AND2_X1 U12061 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10006), .ZN(n9602) );
  OR2_X1 U12062 ( .A1(n10004), .A2(n14956), .ZN(n14954) );
  NOR4_X1 U12063 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_17__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_19__SCAN_IN), .ZN(n9606) );
  NOR4_X1 U12064 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_12__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_15__SCAN_IN), .ZN(n9605) );
  NOR4_X1 U12065 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n9604) );
  NOR4_X1 U12066 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_23__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n9603) );
  NAND4_X1 U12067 ( .A1(n9606), .A2(n9605), .A3(n9604), .A4(n9603), .ZN(n9612)
         );
  NOR2_X1 U12068 ( .A1(P2_D_REG_20__SCAN_IN), .A2(P2_D_REG_8__SCAN_IN), .ZN(
        n9610) );
  NOR4_X1 U12069 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n9609) );
  NOR4_X1 U12070 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_10__SCAN_IN), .A4(P2_D_REG_11__SCAN_IN), .ZN(n9608) );
  NOR4_X1 U12071 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_2__SCAN_IN), .A3(
        P2_D_REG_3__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n9607) );
  NAND4_X1 U12072 ( .A1(n9610), .A2(n9609), .A3(n9608), .A4(n9607), .ZN(n9611)
         );
  OAI21_X1 U12073 ( .B1(n9612), .B2(n9611), .A(n14948), .ZN(n10003) );
  NAND2_X1 U12074 ( .A1(n10533), .A2(n10530), .ZN(n10020) );
  NAND2_X1 U12075 ( .A1(n9579), .A2(n12613), .ZN(n12204) );
  NAND2_X1 U12076 ( .A1(n10015), .A2(n12204), .ZN(n10527) );
  NAND3_X1 U12077 ( .A1(n10003), .A2(n10020), .A3(n10527), .ZN(n9613) );
  NOR2_X1 U12078 ( .A1(n14954), .A2(n9613), .ZN(n10061) );
  INV_X1 U12079 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n14951) );
  NAND2_X1 U12080 ( .A1(n14948), .A2(n14951), .ZN(n9615) );
  NAND2_X1 U12081 ( .A1(n11818), .A2(n11614), .ZN(n9614) );
  NAND2_X1 U12082 ( .A1(n9615), .A2(n9614), .ZN(n14952) );
  AND2_X2 U12083 ( .A1(n10061), .A2(n14952), .ZN(n15007) );
  NAND2_X1 U12084 ( .A1(n10533), .A2(n12204), .ZN(n14999) );
  INV_X1 U12085 ( .A(n14999), .ZN(n14965) );
  NAND2_X1 U12086 ( .A1(n15007), .A2(n14965), .ZN(n13764) );
  NAND2_X1 U12087 ( .A1(n13287), .A2(n9616), .ZN(n9617) );
  NAND2_X1 U12088 ( .A1(n9618), .A2(n9617), .ZN(P2_U3495) );
  OR2_X1 U12089 ( .A1(n14811), .A2(n9621), .ZN(n9622) );
  NAND2_X1 U12090 ( .A1(n9624), .A2(n9623), .ZN(P1_U3556) );
  OR2_X1 U12091 ( .A1(n12419), .A2(n9626), .ZN(n9627) );
  XNOR2_X1 U12092 ( .A(n13084), .B(n10251), .ZN(n9722) );
  NAND2_X1 U12093 ( .A1(n9722), .A2(n9745), .ZN(n9720) );
  INV_X1 U12094 ( .A(n9722), .ZN(n9628) );
  NAND2_X1 U12095 ( .A1(n9628), .A2(n12906), .ZN(n9629) );
  AND2_X1 U12096 ( .A1(n9720), .A2(n9629), .ZN(n12618) );
  XNOR2_X1 U12097 ( .A(n12913), .B(n10251), .ZN(n9630) );
  NAND2_X1 U12098 ( .A1(n9630), .A2(n12926), .ZN(n9715) );
  INV_X1 U12099 ( .A(n9630), .ZN(n9631) );
  NAND2_X1 U12100 ( .A1(n9631), .A2(n12657), .ZN(n9632) );
  AND2_X1 U12101 ( .A1(n9715), .A2(n9632), .ZN(n12721) );
  XNOR2_X1 U12102 ( .A(n14637), .B(n9644), .ZN(n11513) );
  INV_X1 U12103 ( .A(n15141), .ZN(n9633) );
  AOI21_X1 U12104 ( .B1(n9634), .B2(n10251), .A(n9633), .ZN(n9640) );
  OR2_X1 U12105 ( .A1(n15121), .A2(n10251), .ZN(n9635) );
  NAND2_X1 U12106 ( .A1(n12422), .A2(n9635), .ZN(n9636) );
  OR2_X1 U12107 ( .A1(n8551), .A2(n10251), .ZN(n9637) );
  NAND2_X1 U12108 ( .A1(n9636), .A2(n9637), .ZN(n9641) );
  INV_X1 U12109 ( .A(n9637), .ZN(n9638) );
  NAND2_X1 U12110 ( .A1(n9638), .A2(n15121), .ZN(n9639) );
  AND2_X1 U12111 ( .A1(n9641), .A2(n9639), .ZN(n10255) );
  NAND2_X1 U12112 ( .A1(n9640), .A2(n10255), .ZN(n10254) );
  NAND2_X1 U12113 ( .A1(n10254), .A2(n9641), .ZN(n10411) );
  XNOR2_X1 U12114 ( .A(n15117), .B(n9644), .ZN(n9642) );
  XNOR2_X1 U12115 ( .A(n9642), .B(n15137), .ZN(n10412) );
  NAND2_X1 U12116 ( .A1(n10411), .A2(n10412), .ZN(n10481) );
  INV_X1 U12117 ( .A(n9642), .ZN(n9643) );
  XNOR2_X1 U12118 ( .A(n15161), .B(n9644), .ZN(n9646) );
  XNOR2_X1 U12119 ( .A(n9646), .B(n15120), .ZN(n10479) );
  AND2_X1 U12120 ( .A1(n10480), .A2(n10479), .ZN(n9645) );
  INV_X1 U12121 ( .A(n9646), .ZN(n9647) );
  NAND2_X1 U12122 ( .A1(n9647), .A2(n15120), .ZN(n9648) );
  XNOR2_X1 U12123 ( .A(n15168), .B(n10251), .ZN(n9649) );
  OR2_X1 U12124 ( .A1(n9649), .A2(n12744), .ZN(n9651) );
  NAND2_X1 U12125 ( .A1(n9649), .A2(n12744), .ZN(n9650) );
  NAND2_X1 U12126 ( .A1(n9651), .A2(n9650), .ZN(n10650) );
  XNOR2_X1 U12127 ( .A(n15173), .B(n9644), .ZN(n9652) );
  XNOR2_X1 U12128 ( .A(n9652), .B(n12743), .ZN(n10835) );
  XNOR2_X1 U12129 ( .A(n12460), .B(n10251), .ZN(n9659) );
  XNOR2_X1 U12130 ( .A(n9659), .B(n12740), .ZN(n9657) );
  INV_X1 U12131 ( .A(n9652), .ZN(n9653) );
  OR2_X1 U12132 ( .A1(n9653), .A2(n12743), .ZN(n11106) );
  XNOR2_X1 U12133 ( .A(n15178), .B(n9644), .ZN(n11108) );
  INV_X1 U12134 ( .A(n12742), .ZN(n9654) );
  NAND2_X1 U12135 ( .A1(n11108), .A2(n9654), .ZN(n9655) );
  INV_X1 U12136 ( .A(n9657), .ZN(n11292) );
  INV_X1 U12137 ( .A(n11108), .ZN(n9656) );
  NAND2_X1 U12138 ( .A1(n9656), .A2(n12742), .ZN(n11109) );
  OAI21_X1 U12139 ( .B1(n11292), .B2(n11109), .A(n11290), .ZN(n9662) );
  INV_X1 U12140 ( .A(n11290), .ZN(n11110) );
  NAND2_X1 U12141 ( .A1(n9657), .A2(n12741), .ZN(n9658) );
  NAND2_X1 U12142 ( .A1(n11110), .A2(n9658), .ZN(n9661) );
  INV_X1 U12143 ( .A(n9659), .ZN(n9660) );
  AOI22_X1 U12144 ( .A1(n9662), .A2(n9661), .B1(n9660), .B2(n12740), .ZN(n9663) );
  NAND2_X1 U12145 ( .A1(n9664), .A2(n9663), .ZN(n11046) );
  XNOR2_X1 U12146 ( .A(n15193), .B(n10251), .ZN(n9665) );
  XNOR2_X1 U12147 ( .A(n9665), .B(n12739), .ZN(n11047) );
  XNOR2_X1 U12148 ( .A(n15199), .B(n9644), .ZN(n9667) );
  XNOR2_X1 U12149 ( .A(n9667), .B(n12738), .ZN(n11120) );
  OR2_X1 U12150 ( .A1(n9665), .A2(n12739), .ZN(n11121) );
  AND2_X1 U12151 ( .A1(n11120), .A2(n11121), .ZN(n9666) );
  INV_X1 U12152 ( .A(n9667), .ZN(n9668) );
  NAND2_X1 U12153 ( .A1(n9668), .A2(n12738), .ZN(n9669) );
  XNOR2_X1 U12154 ( .A(n14633), .B(n9644), .ZN(n11580) );
  AOI22_X1 U12155 ( .A1(n11580), .A2(n12737), .B1(n11513), .B2(n11518), .ZN(
        n9670) );
  INV_X1 U12156 ( .A(n11580), .ZN(n9671) );
  NAND2_X1 U12157 ( .A1(n9671), .A2(n11720), .ZN(n9672) );
  NAND2_X1 U12158 ( .A1(n9673), .A2(n9672), .ZN(n11437) );
  XNOR2_X1 U12159 ( .A(n14625), .B(n9644), .ZN(n11435) );
  AND2_X1 U12160 ( .A1(n11435), .A2(n11789), .ZN(n9674) );
  INV_X1 U12161 ( .A(n11435), .ZN(n9675) );
  NAND2_X1 U12162 ( .A1(n9675), .A2(n12736), .ZN(n9676) );
  XNOR2_X1 U12163 ( .A(n13140), .B(n10251), .ZN(n9677) );
  NAND2_X1 U12164 ( .A1(n9677), .A2(n13066), .ZN(n9680) );
  INV_X1 U12165 ( .A(n9677), .ZN(n9678) );
  NAND2_X1 U12166 ( .A1(n9678), .A2(n11441), .ZN(n9679) );
  NAND2_X1 U12167 ( .A1(n9680), .A2(n9679), .ZN(n11642) );
  XNOR2_X1 U12168 ( .A(n11712), .B(n10251), .ZN(n11708) );
  OAI21_X1 U12169 ( .B1(n11710), .B2(n13054), .A(n11708), .ZN(n9682) );
  NAND2_X1 U12170 ( .A1(n11710), .A2(n13054), .ZN(n9681) );
  NAND2_X1 U12171 ( .A1(n9682), .A2(n9681), .ZN(n11781) );
  XNOR2_X1 U12172 ( .A(n13184), .B(n9644), .ZN(n11779) );
  AND2_X1 U12173 ( .A1(n11779), .A2(n13068), .ZN(n9683) );
  INV_X1 U12174 ( .A(n11779), .ZN(n9684) );
  NAND2_X1 U12175 ( .A1(n9684), .A2(n12734), .ZN(n9685) );
  XNOR2_X1 U12176 ( .A(n13126), .B(n9644), .ZN(n9687) );
  XNOR2_X1 U12177 ( .A(n9687), .B(n13053), .ZN(n12660) );
  NAND2_X1 U12178 ( .A1(n9687), .A2(n11782), .ZN(n9688) );
  XNOR2_X1 U12179 ( .A(n13122), .B(n9644), .ZN(n9689) );
  XNOR2_X1 U12180 ( .A(n9689), .B(n13037), .ZN(n12695) );
  XNOR2_X1 U12181 ( .A(n13175), .B(n9644), .ZN(n9690) );
  XNOR2_X1 U12182 ( .A(n9690), .B(n12995), .ZN(n12633) );
  NAND2_X1 U12183 ( .A1(n12632), .A2(n12633), .ZN(n9693) );
  INV_X1 U12184 ( .A(n9690), .ZN(n9691) );
  NAND2_X1 U12185 ( .A1(n9691), .A2(n12995), .ZN(n9692) );
  NAND2_X1 U12186 ( .A1(n9693), .A2(n9692), .ZN(n12678) );
  XNOR2_X1 U12187 ( .A(n13000), .B(n9644), .ZN(n9694) );
  XNOR2_X1 U12188 ( .A(n9694), .B(n13009), .ZN(n12679) );
  NAND2_X1 U12189 ( .A1(n9694), .A2(n12529), .ZN(n9695) );
  XNOR2_X1 U12190 ( .A(n12644), .B(n10251), .ZN(n9696) );
  NAND2_X1 U12191 ( .A1(n9696), .A2(n12974), .ZN(n9699) );
  INV_X1 U12192 ( .A(n9696), .ZN(n9697) );
  NAND2_X1 U12193 ( .A1(n9697), .A2(n12996), .ZN(n9698) );
  NAND2_X1 U12194 ( .A1(n9699), .A2(n9698), .ZN(n12640) );
  XNOR2_X1 U12195 ( .A(n12686), .B(n10251), .ZN(n9700) );
  NAND2_X1 U12196 ( .A1(n9701), .A2(n9700), .ZN(n9703) );
  NAND2_X1 U12197 ( .A1(n12687), .A2(n9703), .ZN(n9705) );
  XNOR2_X1 U12198 ( .A(n12969), .B(n9644), .ZN(n9704) );
  NAND2_X2 U12199 ( .A1(n9705), .A2(n9704), .ZN(n12667) );
  OAI21_X1 U12200 ( .B1(n9705), .B2(n9704), .A(n12667), .ZN(n12626) );
  OR2_X2 U12201 ( .A1(n12626), .A2(n12732), .ZN(n12625) );
  NAND2_X1 U12202 ( .A1(n12625), .A2(n12667), .ZN(n9709) );
  XNOR2_X1 U12203 ( .A(n13159), .B(n9644), .ZN(n9706) );
  NAND2_X1 U12204 ( .A1(n9706), .A2(n12925), .ZN(n12649) );
  INV_X1 U12205 ( .A(n9706), .ZN(n9707) );
  NAND2_X1 U12206 ( .A1(n9707), .A2(n12957), .ZN(n9708) );
  AND2_X1 U12207 ( .A1(n12649), .A2(n9708), .ZN(n12668) );
  NAND2_X1 U12208 ( .A1(n9709), .A2(n12668), .ZN(n12648) );
  NAND2_X1 U12209 ( .A1(n12648), .A2(n12649), .ZN(n9713) );
  XNOR2_X1 U12210 ( .A(n12548), .B(n10251), .ZN(n9710) );
  NAND2_X1 U12211 ( .A1(n9710), .A2(n12943), .ZN(n9714) );
  INV_X1 U12212 ( .A(n9710), .ZN(n9711) );
  NAND2_X1 U12213 ( .A1(n9711), .A2(n12905), .ZN(n9712) );
  AND2_X1 U12214 ( .A1(n9714), .A2(n9712), .ZN(n12650) );
  NAND2_X1 U12215 ( .A1(n9713), .A2(n12650), .ZN(n12652) );
  NAND2_X1 U12216 ( .A1(n12618), .A2(n12617), .ZN(n12616) );
  XNOR2_X1 U12217 ( .A(n12560), .B(n10251), .ZN(n9721) );
  INV_X1 U12218 ( .A(n9721), .ZN(n9723) );
  AND2_X1 U12219 ( .A1(n9730), .A2(n15200), .ZN(n10153) );
  AND2_X1 U12220 ( .A1(n9729), .A2(n9725), .ZN(n9716) );
  NAND2_X1 U12221 ( .A1(n10153), .A2(n9716), .ZN(n9719) );
  INV_X1 U12222 ( .A(n9735), .ZN(n9717) );
  NAND2_X1 U12223 ( .A1(n9742), .A2(n9717), .ZN(n9718) );
  NAND2_X1 U12224 ( .A1(n9719), .A2(n9718), .ZN(n12722) );
  NAND2_X1 U12225 ( .A1(n9723), .A2(n12722), .ZN(n9750) );
  NAND2_X1 U12226 ( .A1(n12616), .A2(n7549), .ZN(n9749) );
  NAND4_X1 U12227 ( .A1(n9723), .A2(n9745), .A3(n9722), .A4(n12722), .ZN(n9748) );
  NOR2_X1 U12228 ( .A1(n15200), .A2(n10200), .ZN(n9724) );
  NAND2_X1 U12229 ( .A1(n9729), .A2(n9724), .ZN(n9727) );
  NAND2_X1 U12230 ( .A1(n9725), .A2(n15134), .ZN(n9726) );
  NAND2_X1 U12231 ( .A1(n9727), .A2(n15118), .ZN(n12702) );
  INV_X1 U12232 ( .A(n9737), .ZN(n9728) );
  OR3_X1 U12233 ( .A1(n12582), .A2(n9728), .A3(n12581), .ZN(n12726) );
  INV_X1 U12234 ( .A(n9729), .ZN(n9731) );
  NAND2_X1 U12235 ( .A1(n9731), .A2(n9730), .ZN(n9734) );
  OAI211_X1 U12236 ( .C1(n9115), .C2(n12578), .A(n10197), .B(n9753), .ZN(n9732) );
  INV_X1 U12237 ( .A(n9732), .ZN(n9733) );
  OAI211_X1 U12238 ( .C1(n9737), .C2(n9735), .A(n9734), .B(n9733), .ZN(n9736)
         );
  NAND2_X1 U12239 ( .A1(n9736), .A2(P3_STATE_REG_SCAN_IN), .ZN(n9739) );
  OR2_X1 U12240 ( .A1(n12582), .A2(n9737), .ZN(n9738) );
  NAND2_X1 U12241 ( .A1(n9739), .A2(n9738), .ZN(n12724) );
  AOI22_X1 U12242 ( .A1(n12883), .A2(n12724), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n9744) );
  NOR2_X1 U12243 ( .A1(n13069), .A2(n9740), .ZN(n9741) );
  NAND2_X1 U12244 ( .A1(n12876), .A2(n12728), .ZN(n9743) );
  OAI211_X1 U12245 ( .C1(n9745), .C2(n12726), .A(n9744), .B(n9743), .ZN(n9746)
         );
  AOI21_X1 U12246 ( .B1(n12882), .B2(n12702), .A(n9746), .ZN(n9747) );
  OAI211_X1 U12247 ( .C1(n12616), .C2(n9750), .A(n9749), .B(n7548), .ZN(
        P3_U3160) );
  NAND2_X1 U12248 ( .A1(n11481), .A2(n9751), .ZN(n9843) );
  NOR2_X1 U12249 ( .A1(P2_U3088), .A2(n9843), .ZN(P2_U3947) );
  INV_X1 U12250 ( .A(n9780), .ZN(n9752) );
  NOR2_X2 U12251 ( .A1(n10035), .A2(n9752), .ZN(P1_U4016) );
  INV_X1 U12252 ( .A(n13193), .ZN(n13191) );
  NOR2_X2 U12253 ( .A1(n9753), .A2(n13191), .ZN(P3_U3897) );
  AND2_X1 U12254 ( .A1(n8538), .A2(P1_U3086), .ZN(n10083) );
  INV_X2 U12255 ( .A(n10083), .ZN(n14433) );
  NOR2_X1 U12256 ( .A1(n8538), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14425) );
  OAI222_X1 U12257 ( .A1(n14433), .A2(n9754), .B1(n12610), .B2(n9797), .C1(
        n14727), .C2(P1_U3086), .ZN(P1_U3353) );
  INV_X1 U12258 ( .A(n9755), .ZN(n9770) );
  INV_X1 U12259 ( .A(n13957), .ZN(n9756) );
  OAI222_X1 U12260 ( .A1(n14433), .A2(n9757), .B1(n12610), .B2(n9770), .C1(
        P1_U3086), .C2(n9756), .ZN(P1_U3352) );
  INV_X1 U12261 ( .A(n9758), .ZN(n9760) );
  INV_X1 U12262 ( .A(SI_6_), .ZN(n9759) );
  INV_X1 U12263 ( .A(n10899), .ZN(n12351) );
  OAI222_X1 U12264 ( .A1(n13213), .A2(n9760), .B1(n13217), .B2(n9759), .C1(
        P3_U3151), .C2(n12351), .ZN(P3_U3289) );
  INV_X1 U12265 ( .A(n10895), .ZN(n15061) );
  OAI222_X1 U12266 ( .A1(P3_U3151), .A2(n15061), .B1(n13217), .B2(n9762), .C1(
        n13213), .C2(n9761), .ZN(P3_U3291) );
  OAI222_X1 U12267 ( .A1(P3_U3151), .A2(n12338), .B1(n13217), .B2(n9764), .C1(
        n13213), .C2(n9763), .ZN(P3_U3288) );
  INV_X1 U12268 ( .A(n10345), .ZN(n10221) );
  INV_X1 U12269 ( .A(n9765), .ZN(n9766) );
  OAI222_X1 U12270 ( .A1(P3_U3151), .A2(n10221), .B1(n13217), .B2(n7389), .C1(
        n9766), .C2(n13213), .ZN(P3_U3294) );
  INV_X1 U12271 ( .A(n9767), .ZN(n9771) );
  INV_X1 U12272 ( .A(n13977), .ZN(n13975) );
  OAI222_X1 U12273 ( .A1(n14433), .A2(n9768), .B1(n12610), .B2(n9771), .C1(
        P1_U3086), .C2(n13975), .ZN(P1_U3351) );
  NAND2_X1 U12274 ( .A1(n9769), .A2(P2_U3088), .ZN(n13768) );
  AND2_X1 U12275 ( .A1(n8538), .A2(P2_U3088), .ZN(n13775) );
  INV_X1 U12276 ( .A(n9863), .ZN(n14825) );
  OAI222_X1 U12277 ( .A1(n13768), .A2(n10032), .B1(n6551), .B2(n9770), .C1(
        P2_U3088), .C2(n14825), .ZN(P2_U3324) );
  OAI222_X1 U12278 ( .A1(n13768), .A2(n15480), .B1(n6551), .B2(n9771), .C1(
        P2_U3088), .C2(n14837), .ZN(P2_U3323) );
  OAI222_X1 U12279 ( .A1(n14433), .A2(n9772), .B1(n12610), .B2(n9796), .C1(
        n9953), .C2(P1_U3086), .ZN(P1_U3350) );
  OAI222_X1 U12280 ( .A1(n14433), .A2(n6713), .B1(n12610), .B2(n9800), .C1(
        n9934), .C2(P1_U3086), .ZN(P1_U3354) );
  INV_X1 U12281 ( .A(n13989), .ZN(n9925) );
  OAI222_X1 U12282 ( .A1(P1_U3086), .A2(n9925), .B1(n12610), .B2(n9802), .C1(
        n9773), .C2(n14433), .ZN(P1_U3349) );
  INV_X1 U12283 ( .A(n9774), .ZN(n9775) );
  NAND2_X1 U12284 ( .A1(n10035), .A2(n9780), .ZN(n10055) );
  INV_X1 U12285 ( .A(n10055), .ZN(n10046) );
  NAND2_X1 U12286 ( .A1(n9775), .A2(n10046), .ZN(n14789) );
  AOI22_X1 U12287 ( .A1(n14789), .A2(n9777), .B1(n9780), .B2(n9776), .ZN(
        P1_U3445) );
  INV_X1 U12288 ( .A(n9778), .ZN(n9779) );
  AOI22_X1 U12289 ( .A1(n14789), .A2(n9781), .B1(n9780), .B2(n9779), .ZN(
        P1_U3446) );
  OAI222_X1 U12290 ( .A1(P3_U3151), .A2(n15101), .B1(n13217), .B2(n9783), .C1(
        n13213), .C2(n9782), .ZN(P3_U3286) );
  OAI222_X1 U12291 ( .A1(P3_U3151), .A2(n11246), .B1(n13217), .B2(n9785), .C1(
        n13213), .C2(n9784), .ZN(P3_U3285) );
  OAI222_X1 U12292 ( .A1(P3_U3151), .A2(n15045), .B1(n13217), .B2(n9787), .C1(
        n13213), .C2(n9786), .ZN(P3_U3292) );
  OAI222_X1 U12293 ( .A1(P3_U3151), .A2(n15083), .B1(n13217), .B2(n9789), .C1(
        n13213), .C2(n9788), .ZN(P3_U3290) );
  INV_X1 U12294 ( .A(SI_8_), .ZN(n9792) );
  INV_X1 U12295 ( .A(n9790), .ZN(n9791) );
  OAI222_X1 U12296 ( .A1(P3_U3151), .A2(n12324), .B1(n13217), .B2(n9792), .C1(
        n13213), .C2(n9791), .ZN(P3_U3287) );
  OAI222_X1 U12297 ( .A1(n7199), .A2(P3_U3151), .B1(n13213), .B2(n9793), .C1(
        n15292), .C2(n13217), .ZN(P3_U3293) );
  INV_X1 U12298 ( .A(n9941), .ZN(n14001) );
  OAI222_X1 U12299 ( .A1(n14433), .A2(n9794), .B1(n12610), .B2(n9799), .C1(
        n14001), .C2(P1_U3086), .ZN(P1_U3348) );
  INV_X1 U12300 ( .A(n9871), .ZN(n9880) );
  INV_X1 U12301 ( .A(n13768), .ZN(n10457) );
  INV_X1 U12302 ( .A(n10457), .ZN(n13780) );
  OAI222_X1 U12303 ( .A1(P2_U3088), .A2(n9880), .B1(n6551), .B2(n9796), .C1(
        n9795), .C2(n13780), .ZN(P2_U3322) );
  OAI222_X1 U12304 ( .A1(P2_U3088), .A2(n9861), .B1(n6551), .B2(n9797), .C1(
        n10028), .C2(n13780), .ZN(P2_U3325) );
  INV_X1 U12305 ( .A(n13376), .ZN(n9983) );
  OAI222_X1 U12306 ( .A1(P2_U3088), .A2(n9983), .B1(n6551), .B2(n9799), .C1(
        n9798), .C2(n13780), .ZN(P2_U3320) );
  OAI222_X1 U12307 ( .A1(P2_U3088), .A2(n9860), .B1(n6551), .B2(n9800), .C1(
        n10030), .C2(n13780), .ZN(P2_U3326) );
  INV_X1 U12308 ( .A(n9987), .ZN(n9982) );
  OAI222_X1 U12309 ( .A1(P2_U3088), .A2(n9982), .B1(n6551), .B2(n9802), .C1(
        n9801), .C2(n13780), .ZN(P2_U3321) );
  INV_X1 U12310 ( .A(n13213), .ZN(n13202) );
  INV_X1 U12311 ( .A(n13217), .ZN(n13200) );
  AOI222_X1 U12312 ( .A1(n9803), .A2(n13202), .B1(n11484), .B2(
        P3_STATE_REG_SCAN_IN), .C1(SI_11_), .C2(n13200), .ZN(n9804) );
  INV_X1 U12313 ( .A(n9804), .ZN(P3_U3284) );
  NOR2_X1 U12314 ( .A1(n9805), .A2(n13191), .ZN(n9807) );
  INV_X1 U12315 ( .A(P3_D_REG_12__SCAN_IN), .ZN(n9806) );
  NOR2_X1 U12316 ( .A1(n9828), .A2(n9806), .ZN(P3_U3253) );
  NOR2_X1 U12317 ( .A1(n9807), .A2(n15265), .ZN(P3_U3251) );
  CLKBUF_X1 U12318 ( .A(n9807), .Z(n9828) );
  NOR2_X1 U12319 ( .A1(n9828), .A2(n15254), .ZN(P3_U3237) );
  INV_X1 U12320 ( .A(P3_D_REG_29__SCAN_IN), .ZN(n9808) );
  NOR2_X1 U12321 ( .A1(n9828), .A2(n9808), .ZN(P3_U3236) );
  INV_X1 U12322 ( .A(P3_D_REG_17__SCAN_IN), .ZN(n9809) );
  NOR2_X1 U12323 ( .A1(n9807), .A2(n9809), .ZN(P3_U3248) );
  INV_X1 U12324 ( .A(P3_D_REG_18__SCAN_IN), .ZN(n9810) );
  NOR2_X1 U12325 ( .A1(n9807), .A2(n9810), .ZN(P3_U3247) );
  INV_X1 U12326 ( .A(P3_D_REG_19__SCAN_IN), .ZN(n9811) );
  NOR2_X1 U12327 ( .A1(n9807), .A2(n9811), .ZN(P3_U3246) );
  INV_X1 U12328 ( .A(P3_D_REG_20__SCAN_IN), .ZN(n9812) );
  NOR2_X1 U12329 ( .A1(n9828), .A2(n9812), .ZN(P3_U3245) );
  INV_X1 U12330 ( .A(P3_D_REG_21__SCAN_IN), .ZN(n9813) );
  NOR2_X1 U12331 ( .A1(n9828), .A2(n9813), .ZN(P3_U3244) );
  INV_X1 U12332 ( .A(P3_D_REG_22__SCAN_IN), .ZN(n9814) );
  NOR2_X1 U12333 ( .A1(n9828), .A2(n9814), .ZN(P3_U3243) );
  INV_X1 U12334 ( .A(P3_D_REG_23__SCAN_IN), .ZN(n9815) );
  NOR2_X1 U12335 ( .A1(n9828), .A2(n9815), .ZN(P3_U3242) );
  INV_X1 U12336 ( .A(P3_D_REG_13__SCAN_IN), .ZN(n9816) );
  NOR2_X1 U12337 ( .A1(n9807), .A2(n9816), .ZN(P3_U3252) );
  INV_X1 U12338 ( .A(P3_D_REG_25__SCAN_IN), .ZN(n9817) );
  NOR2_X1 U12339 ( .A1(n9828), .A2(n9817), .ZN(P3_U3240) );
  NOR2_X1 U12340 ( .A1(n9828), .A2(n15365), .ZN(P3_U3239) );
  INV_X1 U12341 ( .A(P3_D_REG_27__SCAN_IN), .ZN(n9818) );
  NOR2_X1 U12342 ( .A1(n9828), .A2(n9818), .ZN(P3_U3238) );
  INV_X1 U12343 ( .A(P3_D_REG_10__SCAN_IN), .ZN(n9819) );
  NOR2_X1 U12344 ( .A1(n9807), .A2(n9819), .ZN(P3_U3255) );
  INV_X1 U12345 ( .A(P3_D_REG_30__SCAN_IN), .ZN(n9820) );
  NOR2_X1 U12346 ( .A1(n9828), .A2(n9820), .ZN(P3_U3235) );
  INV_X1 U12347 ( .A(P3_D_REG_31__SCAN_IN), .ZN(n9821) );
  NOR2_X1 U12348 ( .A1(n9828), .A2(n9821), .ZN(P3_U3234) );
  INV_X1 U12349 ( .A(P3_D_REG_9__SCAN_IN), .ZN(n15379) );
  NOR2_X1 U12350 ( .A1(n9807), .A2(n15379), .ZN(P3_U3256) );
  INV_X1 U12351 ( .A(P3_D_REG_8__SCAN_IN), .ZN(n9822) );
  NOR2_X1 U12352 ( .A1(n9807), .A2(n9822), .ZN(P3_U3257) );
  NOR2_X1 U12353 ( .A1(n9828), .A2(n15226), .ZN(P3_U3258) );
  INV_X1 U12354 ( .A(P3_D_REG_6__SCAN_IN), .ZN(n9823) );
  NOR2_X1 U12355 ( .A1(n9807), .A2(n9823), .ZN(P3_U3259) );
  INV_X1 U12356 ( .A(P3_D_REG_24__SCAN_IN), .ZN(n9824) );
  NOR2_X1 U12357 ( .A1(n9828), .A2(n9824), .ZN(P3_U3241) );
  INV_X1 U12358 ( .A(P3_D_REG_5__SCAN_IN), .ZN(n9825) );
  NOR2_X1 U12359 ( .A1(n9828), .A2(n9825), .ZN(P3_U3260) );
  INV_X1 U12360 ( .A(P3_D_REG_4__SCAN_IN), .ZN(n9826) );
  NOR2_X1 U12361 ( .A1(n9807), .A2(n9826), .ZN(P3_U3261) );
  INV_X1 U12362 ( .A(P3_D_REG_3__SCAN_IN), .ZN(n9827) );
  NOR2_X1 U12363 ( .A1(n9828), .A2(n9827), .ZN(P3_U3262) );
  INV_X1 U12364 ( .A(P3_D_REG_2__SCAN_IN), .ZN(n9829) );
  NOR2_X1 U12365 ( .A1(n9807), .A2(n9829), .ZN(P3_U3263) );
  INV_X1 U12366 ( .A(P3_D_REG_15__SCAN_IN), .ZN(n9830) );
  NOR2_X1 U12367 ( .A1(n9828), .A2(n9830), .ZN(P3_U3250) );
  INV_X1 U12368 ( .A(P3_D_REG_16__SCAN_IN), .ZN(n9831) );
  NOR2_X1 U12369 ( .A1(n9828), .A2(n9831), .ZN(P3_U3249) );
  INV_X1 U12370 ( .A(P3_D_REG_11__SCAN_IN), .ZN(n9832) );
  NOR2_X1 U12371 ( .A1(n9828), .A2(n9832), .ZN(P3_U3254) );
  INV_X1 U12372 ( .A(n9971), .ZN(n9966) );
  OAI222_X1 U12373 ( .A1(n14433), .A2(n9833), .B1(P1_U3086), .B2(n9966), .C1(
        n9835), .C2(n12610), .ZN(P1_U3347) );
  INV_X1 U12374 ( .A(n9991), .ZN(n14851) );
  OAI222_X1 U12375 ( .A1(P2_U3088), .A2(n14851), .B1(n6551), .B2(n9835), .C1(
        n9834), .C2(n13780), .ZN(P2_U3319) );
  AOI222_X1 U12376 ( .A1(n9836), .A2(n13202), .B1(n12751), .B2(
        P3_STATE_REG_SCAN_IN), .C1(SI_12_), .C2(n13200), .ZN(n9837) );
  INV_X1 U12377 ( .A(n9837), .ZN(P3_U3283) );
  INV_X1 U12378 ( .A(n10110), .ZN(n10106) );
  OAI222_X1 U12379 ( .A1(P2_U3088), .A2(n10106), .B1(n6551), .B2(n9839), .C1(
        n9838), .C2(n13780), .ZN(P2_U3318) );
  INV_X1 U12380 ( .A(n9972), .ZN(n10166) );
  OAI222_X1 U12381 ( .A1(n14433), .A2(n9840), .B1(n12610), .B2(n9839), .C1(
        n10166), .C2(P1_U3086), .ZN(P1_U3346) );
  NAND2_X1 U12382 ( .A1(n10015), .A2(n11481), .ZN(n9842) );
  NAND2_X1 U12383 ( .A1(n9842), .A2(n9841), .ZN(n9844) );
  NAND2_X1 U12384 ( .A1(n9844), .A2(n9843), .ZN(n9866) );
  AND2_X1 U12385 ( .A1(n9852), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9845) );
  INV_X1 U12386 ( .A(n14914), .ZN(n14921) );
  INV_X1 U12387 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n9857) );
  MUX2_X1 U12388 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n9219), .S(n9871), .Z(n9855)
         );
  INV_X1 U12389 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10065) );
  MUX2_X1 U12390 ( .A(n10065), .B(P2_REG1_REG_1__SCAN_IN), .S(n9860), .Z(n9893) );
  AND2_X1 U12391 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n9892) );
  NAND2_X1 U12392 ( .A1(n9893), .A2(n9892), .ZN(n9891) );
  INV_X1 U12393 ( .A(n9860), .ZN(n9890) );
  NAND2_X1 U12394 ( .A1(n9890), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n9846) );
  NAND2_X1 U12395 ( .A1(n9891), .A2(n9846), .ZN(n9903) );
  INV_X1 U12396 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n9847) );
  MUX2_X1 U12397 ( .A(n9847), .B(P2_REG1_REG_2__SCAN_IN), .S(n9861), .Z(n9904)
         );
  NAND2_X1 U12398 ( .A1(n9903), .A2(n9904), .ZN(n9902) );
  INV_X1 U12399 ( .A(n9861), .ZN(n9901) );
  NAND2_X1 U12400 ( .A1(n9901), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n9848) );
  NAND2_X1 U12401 ( .A1(n9902), .A2(n9848), .ZN(n14821) );
  INV_X1 U12402 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10148) );
  MUX2_X1 U12403 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n10148), .S(n9863), .Z(
        n14822) );
  NAND2_X1 U12404 ( .A1(n14821), .A2(n14822), .ZN(n14820) );
  NAND2_X1 U12405 ( .A1(n9863), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n9849) );
  NAND2_X1 U12406 ( .A1(n14820), .A2(n9849), .ZN(n14833) );
  MUX2_X1 U12407 ( .A(n9206), .B(P2_REG1_REG_4__SCAN_IN), .S(n14837), .Z(
        n14834) );
  NAND2_X1 U12408 ( .A1(n14833), .A2(n14834), .ZN(n14832) );
  NAND2_X1 U12409 ( .A1(n9850), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n9851) );
  NAND2_X1 U12410 ( .A1(n14832), .A2(n9851), .ZN(n9854) );
  OR2_X1 U12411 ( .A1(n9852), .A2(P2_U3088), .ZN(n13777) );
  INV_X1 U12412 ( .A(n13418), .ZN(n12306) );
  NOR2_X1 U12413 ( .A1(n13777), .A2(n12306), .ZN(n9853) );
  AND2_X1 U12414 ( .A1(n9866), .A2(n9853), .ZN(n14846) );
  NAND2_X1 U12415 ( .A1(n9854), .A2(n9855), .ZN(n9873) );
  OAI211_X1 U12416 ( .C1(n9855), .C2(n9854), .A(n14846), .B(n9873), .ZN(n9856)
         );
  NAND2_X1 U12417 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3088), .ZN(n10467) );
  OAI211_X1 U12418 ( .C1(n9857), .C2(n14932), .A(n9856), .B(n10467), .ZN(n9858) );
  INV_X1 U12419 ( .A(n9858), .ZN(n9870) );
  MUX2_X1 U12420 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n10663), .S(n9871), .Z(n9868) );
  MUX2_X1 U12421 ( .A(n9859), .B(P2_REG2_REG_1__SCAN_IN), .S(n9860), .Z(n9887)
         );
  NAND3_X1 U12422 ( .A1(n9887), .A2(P2_REG2_REG_0__SCAN_IN), .A3(
        P2_IR_REG_0__SCAN_IN), .ZN(n9885) );
  OAI21_X1 U12423 ( .B1(n9860), .B2(n9859), .A(n9885), .ZN(n9897) );
  MUX2_X1 U12424 ( .A(n9862), .B(P2_REG2_REG_2__SCAN_IN), .S(n9861), .Z(n9898)
         );
  NAND2_X1 U12425 ( .A1(n9897), .A2(n9898), .ZN(n9896) );
  MUX2_X1 U12426 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n9864), .S(n9863), .Z(n14819) );
  MUX2_X1 U12427 ( .A(n10613), .B(P2_REG2_REG_4__SCAN_IN), .S(n14837), .Z(
        n14831) );
  OAI21_X1 U12428 ( .B1(n10613), .B2(n14837), .A(n14829), .ZN(n9867) );
  NOR2_X1 U12429 ( .A1(n13777), .A2(n13418), .ZN(n9865) );
  AND2_X1 U12430 ( .A1(n9866), .A2(n9865), .ZN(n14929) );
  NAND2_X1 U12431 ( .A1(n9867), .A2(n9868), .ZN(n9879) );
  OAI211_X1 U12432 ( .C1(n9868), .C2(n9867), .A(n14929), .B(n9879), .ZN(n9869)
         );
  OAI211_X1 U12433 ( .C1(n14921), .C2(n9880), .A(n9870), .B(n9869), .ZN(
        P2_U3219) );
  INV_X1 U12434 ( .A(n14932), .ZN(n14813) );
  INV_X1 U12435 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n15011) );
  MUX2_X1 U12436 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n15011), .S(n9987), .Z(n9875) );
  NAND2_X1 U12437 ( .A1(n9871), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n9872) );
  NAND2_X1 U12438 ( .A1(n9873), .A2(n9872), .ZN(n9874) );
  NAND2_X1 U12439 ( .A1(n9874), .A2(n9875), .ZN(n9989) );
  OAI211_X1 U12440 ( .C1(n9875), .C2(n9874), .A(n14846), .B(n9989), .ZN(n9877)
         );
  NAND2_X1 U12441 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3088), .ZN(n9876) );
  NAND2_X1 U12442 ( .A1(n9877), .A2(n9876), .ZN(n9878) );
  AOI21_X1 U12443 ( .B1(n14813), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n9878), .ZN(
        n9884) );
  XOR2_X1 U12444 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n9987), .Z(n9882) );
  OAI21_X1 U12445 ( .B1(n10663), .B2(n9880), .A(n9879), .ZN(n9881) );
  NAND2_X1 U12446 ( .A1(n9881), .A2(n9882), .ZN(n9981) );
  OAI211_X1 U12447 ( .C1(n9882), .C2(n9881), .A(n14929), .B(n9981), .ZN(n9883)
         );
  OAI211_X1 U12448 ( .C1(n14921), .C2(n9982), .A(n9884), .B(n9883), .ZN(
        P2_U3220) );
  AND2_X1 U12449 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n9886) );
  OAI211_X1 U12450 ( .C1(n9887), .C2(n9886), .A(n14929), .B(n9885), .ZN(n9888)
         );
  OAI21_X1 U12451 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n10027), .A(n9888), .ZN(
        n9889) );
  AOI21_X1 U12452 ( .B1(n9890), .B2(n14914), .A(n9889), .ZN(n9895) );
  OAI211_X1 U12453 ( .C1(n9893), .C2(n9892), .A(n14846), .B(n9891), .ZN(n9894)
         );
  OAI211_X1 U12454 ( .C1(n6696), .C2(n14932), .A(n9895), .B(n9894), .ZN(
        P2_U3215) );
  INV_X1 U12455 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n9907) );
  OAI211_X1 U12456 ( .C1(n9898), .C2(n9897), .A(n14929), .B(n9896), .ZN(n9899)
         );
  OAI21_X1 U12457 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n10101), .A(n9899), .ZN(
        n9900) );
  AOI21_X1 U12458 ( .B1(n9901), .B2(n14914), .A(n9900), .ZN(n9906) );
  OAI211_X1 U12459 ( .C1(n9904), .C2(n9903), .A(n14846), .B(n9902), .ZN(n9905)
         );
  OAI211_X1 U12460 ( .C1(n9907), .C2(n14932), .A(n9906), .B(n9905), .ZN(
        P2_U3216) );
  OAI222_X1 U12461 ( .A1(P3_U3151), .A2(n12772), .B1(n13217), .B2(n9909), .C1(
        n13213), .C2(n9908), .ZN(P3_U3282) );
  INV_X1 U12462 ( .A(P3_DATAO_REG_14__SCAN_IN), .ZN(n15469) );
  NAND2_X1 U12463 ( .A1(n11441), .A2(P3_U3897), .ZN(n9910) );
  OAI21_X1 U12464 ( .B1(P3_U3897), .B2(n15469), .A(n9910), .ZN(P3_U3505) );
  INV_X1 U12465 ( .A(n9911), .ZN(n9912) );
  INV_X1 U12466 ( .A(n10167), .ZN(n14019) );
  OAI222_X1 U12467 ( .A1(n14433), .A2(n15281), .B1(n12610), .B2(n9912), .C1(
        P1_U3086), .C2(n14019), .ZN(P1_U3345) );
  INV_X1 U12468 ( .A(n10269), .ZN(n10262) );
  OAI222_X1 U12469 ( .A1(n13768), .A2(n9913), .B1(n6551), .B2(n9912), .C1(
        P2_U3088), .C2(n10262), .ZN(P2_U3317) );
  NAND2_X1 U12470 ( .A1(n10048), .A2(n9914), .ZN(n9915) );
  NAND2_X1 U12471 ( .A1(n9915), .A2(n7716), .ZN(n9930) );
  AND2_X1 U12472 ( .A1(n10055), .A2(n11477), .ZN(n9929) );
  INV_X1 U12473 ( .A(n9929), .ZN(n9916) );
  CLKBUF_X1 U12474 ( .A(P1_U4016), .Z(n13967) );
  NOR2_X1 U12475 ( .A1(n14719), .A2(n13967), .ZN(P1_U3085) );
  MUX2_X1 U12476 ( .A(n9965), .B(P1_REG1_REG_8__SCAN_IN), .S(n9971), .Z(n9928)
         );
  MUX2_X1 U12477 ( .A(n9918), .B(P1_REG1_REG_2__SCAN_IN), .S(n14727), .Z(
        n14720) );
  INV_X1 U12478 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n15442) );
  MUX2_X1 U12479 ( .A(n15442), .B(P1_REG1_REG_1__SCAN_IN), .S(n9934), .Z(
        n13943) );
  AND2_X1 U12480 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n13942) );
  NAND2_X1 U12481 ( .A1(n13943), .A2(n13942), .ZN(n14721) );
  INV_X1 U12482 ( .A(n9934), .ZN(n13941) );
  NAND2_X1 U12483 ( .A1(n13941), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n14722) );
  NAND2_X1 U12484 ( .A1(n14721), .A2(n14722), .ZN(n9917) );
  NAND2_X1 U12485 ( .A1(n14720), .A2(n9917), .ZN(n14725) );
  OR2_X1 U12486 ( .A1(n14727), .A2(n9918), .ZN(n9919) );
  NAND2_X1 U12487 ( .A1(n14725), .A2(n9919), .ZN(n13950) );
  INV_X1 U12488 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n9920) );
  XNOR2_X1 U12489 ( .A(n13957), .B(n9920), .ZN(n13951) );
  NAND2_X1 U12490 ( .A1(n13950), .A2(n13951), .ZN(n13949) );
  NAND2_X1 U12491 ( .A1(n13957), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n9921) );
  NAND2_X1 U12492 ( .A1(n13949), .A2(n9921), .ZN(n13972) );
  XNOR2_X1 U12493 ( .A(n13977), .B(n9922), .ZN(n13973) );
  NAND2_X1 U12494 ( .A1(n13972), .A2(n13973), .ZN(n13971) );
  OAI21_X1 U12495 ( .B1(n9922), .B2(n13975), .A(n13971), .ZN(n9951) );
  MUX2_X1 U12496 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n9923), .S(n9953), .Z(n9952)
         );
  NOR2_X1 U12497 ( .A1(n9951), .A2(n9952), .ZN(n9950) );
  AOI21_X1 U12498 ( .B1(n9953), .B2(n9923), .A(n9950), .ZN(n13991) );
  XOR2_X1 U12499 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n13989), .Z(n13992) );
  NAND2_X1 U12500 ( .A1(n13991), .A2(n13992), .ZN(n13990) );
  OAI21_X1 U12501 ( .B1(n9925), .B2(n9924), .A(n13990), .ZN(n14006) );
  MUX2_X1 U12502 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n9926), .S(n9941), .Z(n14005) );
  NAND2_X1 U12503 ( .A1(n14006), .A2(n14005), .ZN(n14004) );
  OAI21_X1 U12504 ( .B1(n14001), .B2(n9926), .A(n14004), .ZN(n9927) );
  NOR2_X1 U12505 ( .A1(n9927), .A2(n9928), .ZN(n9964) );
  AOI21_X1 U12506 ( .B1(n9928), .B2(n9927), .A(n9964), .ZN(n9948) );
  OR2_X1 U12507 ( .A1(n9930), .A2(n9929), .ZN(n14717) );
  INV_X1 U12508 ( .A(n13962), .ZN(n14714) );
  OR2_X1 U12509 ( .A1(n14717), .A2(n14714), .ZN(n14040) );
  AND2_X1 U12510 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n9932) );
  OR2_X1 U12511 ( .A1(n14717), .A2(n13965), .ZN(n14744) );
  NOR2_X1 U12512 ( .A1(n14744), .A2(n9966), .ZN(n9931) );
  AOI211_X1 U12513 ( .C1(n14719), .C2(P1_ADDR_REG_8__SCAN_IN), .A(n9932), .B(
        n9931), .ZN(n9947) );
  OR2_X1 U12514 ( .A1(n8158), .A2(n13962), .ZN(n9933) );
  OR2_X1 U12515 ( .A1(n14717), .A2(n9933), .ZN(n14746) );
  MUX2_X1 U12516 ( .A(n15433), .B(P1_REG2_REG_2__SCAN_IN), .S(n14727), .Z(
        n9936) );
  INV_X1 U12517 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n9935) );
  MUX2_X1 U12518 ( .A(n9935), .B(P1_REG2_REG_1__SCAN_IN), .S(n9934), .Z(n13945) );
  AND2_X1 U12519 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n13964) );
  NAND2_X1 U12520 ( .A1(n13945), .A2(n13964), .ZN(n13944) );
  OAI21_X1 U12521 ( .B1(n9935), .B2(n9934), .A(n13944), .ZN(n14726) );
  NAND2_X1 U12522 ( .A1(n9936), .A2(n14726), .ZN(n14728) );
  INV_X1 U12523 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n15433) );
  OR2_X1 U12524 ( .A1(n14727), .A2(n15433), .ZN(n13953) );
  NAND2_X1 U12525 ( .A1(n14728), .A2(n13953), .ZN(n9938) );
  MUX2_X1 U12526 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n10521), .S(n13957), .Z(
        n9937) );
  NAND2_X1 U12527 ( .A1(n9938), .A2(n9937), .ZN(n13980) );
  NAND2_X1 U12528 ( .A1(n13957), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n13979) );
  NAND2_X1 U12529 ( .A1(n13980), .A2(n13979), .ZN(n9940) );
  MUX2_X1 U12530 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n10640), .S(n13977), .Z(
        n9939) );
  NAND2_X1 U12531 ( .A1(n9940), .A2(n9939), .ZN(n13982) );
  NAND2_X1 U12532 ( .A1(n13977), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n9957) );
  MUX2_X1 U12533 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n7763), .S(n9953), .Z(n9956)
         );
  AOI21_X1 U12534 ( .B1(n13982), .B2(n9957), .A(n9956), .ZN(n13995) );
  NOR2_X1 U12535 ( .A1(n9953), .A2(n7763), .ZN(n13994) );
  MUX2_X1 U12536 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n10748), .S(n13989), .Z(
        n13993) );
  OAI21_X1 U12537 ( .B1(n13995), .B2(n13994), .A(n13993), .ZN(n14010) );
  NAND2_X1 U12538 ( .A1(n13989), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n14009) );
  MUX2_X1 U12539 ( .A(n7791), .B(P1_REG2_REG_7__SCAN_IN), .S(n9941), .Z(n14008) );
  AOI21_X1 U12540 ( .B1(n14010), .B2(n14009), .A(n14008), .ZN(n14007) );
  NOR2_X1 U12541 ( .A1(n14001), .A2(n7791), .ZN(n9944) );
  MUX2_X1 U12542 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n9942), .S(n9971), .Z(n9943)
         );
  OAI21_X1 U12543 ( .B1(n14007), .B2(n9944), .A(n9943), .ZN(n9975) );
  OR3_X1 U12544 ( .A1(n14007), .A2(n9944), .A3(n9943), .ZN(n9945) );
  NAND3_X1 U12545 ( .A1(n14059), .A2(n9975), .A3(n9945), .ZN(n9946) );
  OAI211_X1 U12546 ( .C1(n9948), .C2(n14040), .A(n9947), .B(n9946), .ZN(
        P1_U3251) );
  INV_X1 U12547 ( .A(P3_DATAO_REG_17__SCAN_IN), .ZN(n15228) );
  NAND2_X1 U12548 ( .A1(n11782), .A2(P3_U3897), .ZN(n9949) );
  OAI21_X1 U12549 ( .B1(P3_U3897), .B2(n15228), .A(n9949), .ZN(P3_U3508) );
  AOI21_X1 U12550 ( .B1(n9952), .B2(n9951), .A(n9950), .ZN(n9962) );
  AND2_X1 U12551 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n9955) );
  NOR2_X1 U12552 ( .A1(n14744), .A2(n9953), .ZN(n9954) );
  AOI211_X1 U12553 ( .C1(n14719), .C2(P1_ADDR_REG_5__SCAN_IN), .A(n9955), .B(
        n9954), .ZN(n9961) );
  INV_X1 U12554 ( .A(n13995), .ZN(n9959) );
  NAND3_X1 U12555 ( .A1(n13982), .A2(n9957), .A3(n9956), .ZN(n9958) );
  NAND3_X1 U12556 ( .A1(n14059), .A2(n9959), .A3(n9958), .ZN(n9960) );
  OAI211_X1 U12557 ( .C1(n9962), .C2(n14040), .A(n9961), .B(n9960), .ZN(
        P1_U3248) );
  INV_X1 U12558 ( .A(P3_DATAO_REG_11__SCAN_IN), .ZN(n15264) );
  NAND2_X1 U12559 ( .A1(n11518), .A2(P3_U3897), .ZN(n9963) );
  OAI21_X1 U12560 ( .B1(P3_U3897), .B2(n15264), .A(n9963), .ZN(P3_U3502) );
  MUX2_X1 U12561 ( .A(n10160), .B(P1_REG1_REG_9__SCAN_IN), .S(n9972), .Z(n9968) );
  AOI21_X1 U12562 ( .B1(n9966), .B2(n9965), .A(n9964), .ZN(n9967) );
  NOR2_X1 U12563 ( .A1(n9967), .A2(n9968), .ZN(n10159) );
  AOI21_X1 U12564 ( .B1(n9968), .B2(n9967), .A(n10159), .ZN(n9980) );
  INV_X1 U12565 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n11239) );
  NOR2_X1 U12566 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n11239), .ZN(n9970) );
  NOR2_X1 U12567 ( .A1(n14744), .A2(n10166), .ZN(n9969) );
  AOI211_X1 U12568 ( .C1(n14719), .C2(P1_ADDR_REG_9__SCAN_IN), .A(n9970), .B(
        n9969), .ZN(n9979) );
  NAND2_X1 U12569 ( .A1(n9971), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n9974) );
  MUX2_X1 U12570 ( .A(n11025), .B(P1_REG2_REG_9__SCAN_IN), .S(n9972), .Z(n9973) );
  AOI21_X1 U12571 ( .B1(n9975), .B2(n9974), .A(n9973), .ZN(n14024) );
  INV_X1 U12572 ( .A(n14024), .ZN(n9977) );
  NAND3_X1 U12573 ( .A1(n9975), .A2(n9974), .A3(n9973), .ZN(n9976) );
  NAND3_X1 U12574 ( .A1(n9977), .A2(n14059), .A3(n9976), .ZN(n9978) );
  OAI211_X1 U12575 ( .C1(n9980), .C2(n14040), .A(n9979), .B(n9978), .ZN(
        P1_U3252) );
  MUX2_X1 U12576 ( .A(n10922), .B(P2_REG2_REG_9__SCAN_IN), .S(n10110), .Z(
        n9985) );
  OAI21_X1 U12577 ( .B1(n10850), .B2(n9982), .A(n9981), .ZN(n13382) );
  XOR2_X1 U12578 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n13376), .Z(n13383) );
  NAND2_X1 U12579 ( .A1(n13382), .A2(n13383), .ZN(n13381) );
  OAI21_X1 U12580 ( .B1(n10986), .B2(n9983), .A(n13381), .ZN(n14844) );
  MUX2_X1 U12581 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n10720), .S(n9991), .Z(
        n14843) );
  NAND2_X1 U12582 ( .A1(n14844), .A2(n14843), .ZN(n14842) );
  OAI21_X1 U12583 ( .B1(n10720), .B2(n14851), .A(n14842), .ZN(n9984) );
  AOI21_X1 U12584 ( .B1(n9985), .B2(n9984), .A(n10105), .ZN(n9999) );
  INV_X1 U12585 ( .A(n14929), .ZN(n14907) );
  AND2_X1 U12586 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3088), .ZN(n10942) );
  NOR2_X1 U12587 ( .A1(n14932), .A2(n7287), .ZN(n9986) );
  AOI211_X1 U12588 ( .C1(n14914), .C2(n10110), .A(n10942), .B(n9986), .ZN(
        n9998) );
  MUX2_X1 U12589 ( .A(n9273), .B(P2_REG1_REG_9__SCAN_IN), .S(n10110), .Z(n9995) );
  NAND2_X1 U12590 ( .A1(n9987), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n9988) );
  NAND2_X1 U12591 ( .A1(n9989), .A2(n9988), .ZN(n13385) );
  INV_X1 U12592 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n15013) );
  MUX2_X1 U12593 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n15013), .S(n13376), .Z(
        n13386) );
  NAND2_X1 U12594 ( .A1(n13385), .A2(n13386), .ZN(n13384) );
  NAND2_X1 U12595 ( .A1(n13376), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n9990) );
  NAND2_X1 U12596 ( .A1(n13384), .A2(n9990), .ZN(n14847) );
  MUX2_X1 U12597 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n9261), .S(n9991), .Z(n14848) );
  NAND2_X1 U12598 ( .A1(n14847), .A2(n14848), .ZN(n14845) );
  NAND2_X1 U12599 ( .A1(n9991), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n9992) );
  NAND2_X1 U12600 ( .A1(n14845), .A2(n9992), .ZN(n9994) );
  INV_X1 U12601 ( .A(n10112), .ZN(n9993) );
  AOI21_X1 U12602 ( .B1(n9995), .B2(n9994), .A(n9993), .ZN(n9996) );
  INV_X1 U12603 ( .A(n14846), .ZN(n14922) );
  OR2_X1 U12604 ( .A1(n9996), .A2(n14922), .ZN(n9997) );
  OAI211_X1 U12605 ( .C1(n9999), .C2(n14907), .A(n9998), .B(n9997), .ZN(
        P2_U3223) );
  INV_X1 U12606 ( .A(n12776), .ZN(n12781) );
  INV_X1 U12607 ( .A(SI_14_), .ZN(n10002) );
  INV_X1 U12608 ( .A(n10000), .ZN(n10001) );
  OAI222_X1 U12609 ( .A1(P3_U3151), .A2(n12781), .B1(n13217), .B2(n10002), 
        .C1(n13213), .C2(n10001), .ZN(P3_U3281) );
  AND2_X1 U12610 ( .A1(n10004), .A2(n10003), .ZN(n10526) );
  INV_X1 U12611 ( .A(n10526), .ZN(n10005) );
  OAI21_X1 U12612 ( .B1(n10005), .B2(n14952), .A(n10020), .ZN(n10008) );
  AND3_X1 U12613 ( .A1(n10527), .A2(n11481), .A3(n10006), .ZN(n10007) );
  NAND2_X1 U12614 ( .A1(n10008), .A2(n10007), .ZN(n10137) );
  NOR2_X1 U12615 ( .A1(n10137), .A2(P2_U3088), .ZN(n10128) );
  NAND2_X1 U12616 ( .A1(n10429), .A2(n13374), .ZN(n10091) );
  XNOR2_X1 U12617 ( .A(n10090), .B(n10091), .ZN(n10013) );
  NAND2_X1 U12618 ( .A1(n13603), .A2(n12002), .ZN(n10010) );
  NAND2_X1 U12619 ( .A1(n13282), .A2(n12003), .ZN(n10011) );
  NAND2_X1 U12620 ( .A1(n10131), .A2(n10011), .ZN(n10012) );
  OAI21_X1 U12621 ( .B1(n10013), .B2(n10012), .A(n10094), .ZN(n10018) );
  NOR2_X1 U12622 ( .A1(n14952), .A2(n14956), .ZN(n10014) );
  AND2_X1 U12623 ( .A1(n10526), .A2(n10014), .ZN(n10023) );
  INV_X1 U12624 ( .A(n10015), .ZN(n10016) );
  AND2_X1 U12625 ( .A1(n14999), .A2(n10016), .ZN(n10017) );
  NAND2_X1 U12626 ( .A1(n10023), .A2(n10017), .ZN(n13348) );
  INV_X1 U12627 ( .A(n13348), .ZN(n13326) );
  NAND2_X1 U12628 ( .A1(n10018), .A2(n13326), .ZN(n10026) );
  NOR2_X1 U12629 ( .A1(n10019), .A2(n9579), .ZN(n10614) );
  NAND2_X1 U12630 ( .A1(n10023), .A2(n10614), .ZN(n10022) );
  INV_X1 U12631 ( .A(n10020), .ZN(n10021) );
  NAND2_X1 U12632 ( .A1(n10022), .A2(n13535), .ZN(n13346) );
  INV_X1 U12633 ( .A(n12204), .ZN(n12305) );
  INV_X1 U12634 ( .A(n13375), .ZN(n10130) );
  INV_X1 U12635 ( .A(n13496), .ZN(n13548) );
  INV_X1 U12636 ( .A(n13373), .ZN(n10024) );
  OAI22_X1 U12637 ( .A1(n10130), .A2(n13627), .B1(n13548), .B2(n10024), .ZN(
        n10063) );
  AOI22_X1 U12638 ( .A1(n14934), .A2(n13346), .B1(n13342), .B2(n10063), .ZN(
        n10025) );
  OAI211_X1 U12639 ( .C1(n10128), .C2(n10027), .A(n10026), .B(n10025), .ZN(
        P2_U3194) );
  MUX2_X1 U12640 ( .A(n10028), .B(n14771), .S(n13967), .Z(n10029) );
  INV_X1 U12641 ( .A(n10029), .ZN(P1_U3562) );
  MUX2_X1 U12642 ( .A(n10030), .B(n10352), .S(n13967), .Z(n10031) );
  INV_X1 U12643 ( .A(n10031), .ZN(P1_U3561) );
  MUX2_X1 U12644 ( .A(n10032), .B(n7733), .S(n13967), .Z(n10033) );
  INV_X1 U12645 ( .A(n10033), .ZN(P1_U3563) );
  INV_X1 U12646 ( .A(n14763), .ZN(n13939) );
  NAND2_X2 U12647 ( .A1(n10034), .A2(n10035), .ZN(n11939) );
  NAND2_X1 U12648 ( .A1(n13939), .A2(n10626), .ZN(n10038) );
  AOI22_X1 U12649 ( .A1(n11980), .A2(n14780), .B1(n10039), .B2(
        P1_REG1_REG_0__SCAN_IN), .ZN(n10037) );
  AOI22_X1 U12650 ( .A1(n10626), .A2(n14780), .B1(n10039), .B2(
        P1_IR_REG_0__SCAN_IN), .ZN(n10040) );
  OAI21_X1 U12651 ( .B1(n10354), .B2(n14763), .A(n10040), .ZN(n10043) );
  INV_X1 U12652 ( .A(n10043), .ZN(n10041) );
  INV_X1 U12653 ( .A(n10362), .ZN(n10042) );
  AOI21_X1 U12654 ( .B1(n10044), .B2(n10043), .A(n10042), .ZN(n13963) );
  OR2_X1 U12655 ( .A1(n10045), .A2(n10510), .ZN(n10052) );
  INV_X1 U12656 ( .A(n10052), .ZN(n10047) );
  NAND2_X1 U12657 ( .A1(n10047), .A2(n10046), .ZN(n10054) );
  INV_X1 U12658 ( .A(n10048), .ZN(n10049) );
  NAND2_X1 U12659 ( .A1(n14798), .A2(n10049), .ZN(n10050) );
  NOR2_X1 U12660 ( .A1(n10051), .A2(n10052), .ZN(n13818) );
  INV_X1 U12661 ( .A(n14247), .ZN(n14770) );
  NOR2_X1 U12662 ( .A1(n14770), .A2(n10352), .ZN(n14779) );
  INV_X1 U12663 ( .A(n10051), .ZN(n10053) );
  NAND2_X1 U12664 ( .A1(n10052), .A2(n10056), .ZN(n10376) );
  NAND2_X1 U12665 ( .A1(n10053), .A2(n10376), .ZN(n13882) );
  AOI22_X1 U12666 ( .A1(n13818), .A2(n14779), .B1(n13882), .B2(
        P1_REG3_REG_0__SCAN_IN), .ZN(n10059) );
  OR2_X1 U12667 ( .A1(n8155), .A2(n6549), .ZN(n14772) );
  OR2_X1 U12668 ( .A1(n10054), .A2(n14772), .ZN(n10057) );
  OR2_X2 U12669 ( .A1(n10056), .A2(n10055), .ZN(n14777) );
  NAND2_X1 U12670 ( .A1(n10057), .A2(n14777), .ZN(n14679) );
  NAND2_X1 U12671 ( .A1(n14679), .A2(n14780), .ZN(n10058) );
  OAI211_X1 U12672 ( .C1(n13963), .C2(n14674), .A(n10059), .B(n10058), .ZN(
        P1_U3232) );
  INV_X1 U12673 ( .A(n14952), .ZN(n10060) );
  AND2_X2 U12674 ( .A1(n10061), .A2(n10060), .ZN(n15019) );
  XNOR2_X1 U12675 ( .A(n12247), .B(n10532), .ZN(n14941) );
  XNOR2_X1 U12676 ( .A(n12247), .B(n10062), .ZN(n10064) );
  AOI21_X1 U12677 ( .B1(n10064), .B2(n13618), .A(n10063), .ZN(n14946) );
  OAI211_X1 U12678 ( .C1(n10193), .C2(n12003), .A(n13603), .B(n10074), .ZN(
        n14940) );
  OAI211_X1 U12679 ( .C1(n13730), .C2(n14941), .A(n14946), .B(n14940), .ZN(
        n10195) );
  NAND2_X1 U12680 ( .A1(n15019), .A2(n14965), .ZN(n13724) );
  OAI22_X1 U12681 ( .A1(n13724), .A2(n10193), .B1(n15019), .B2(n10065), .ZN(
        n10066) );
  AOI21_X1 U12682 ( .B1(n15019), .B2(n10195), .A(n10066), .ZN(n10067) );
  INV_X1 U12683 ( .A(n10067), .ZN(P2_U3500) );
  INV_X1 U12684 ( .A(n11089), .ZN(n11084) );
  INV_X1 U12685 ( .A(n10068), .ZN(n10071) );
  OAI222_X1 U12686 ( .A1(P2_U3088), .A2(n11084), .B1(n6551), .B2(n10071), .C1(
        n10069), .C2(n13780), .ZN(P2_U3316) );
  INV_X1 U12687 ( .A(n10402), .ZN(n10400) );
  OAI222_X1 U12688 ( .A1(P1_U3086), .A2(n10400), .B1(n12610), .B2(n10071), 
        .C1(n10070), .C2(n14433), .ZN(P1_U3344) );
  INV_X1 U12689 ( .A(n13730), .ZN(n14983) );
  OAI21_X1 U12690 ( .B1(n10073), .B2(n10078), .A(n10072), .ZN(n11035) );
  INV_X1 U12691 ( .A(n10146), .ZN(n10076) );
  NAND2_X1 U12692 ( .A1(n10074), .A2(n12016), .ZN(n10075) );
  AND3_X1 U12693 ( .A1(n13603), .A2(n10076), .A3(n10075), .ZN(n11036) );
  XNOR2_X1 U12694 ( .A(n10078), .B(n10077), .ZN(n10080) );
  INV_X1 U12695 ( .A(n13374), .ZN(n12010) );
  OAI22_X1 U12696 ( .A1(n12010), .A2(n13627), .B1(n13548), .B2(n9196), .ZN(
        n10098) );
  INV_X1 U12697 ( .A(n10098), .ZN(n10079) );
  OAI21_X1 U12698 ( .B1(n10080), .B2(n13600), .A(n10079), .ZN(n11042) );
  AOI211_X1 U12699 ( .C1(n14983), .C2(n11035), .A(n11036), .B(n11042), .ZN(
        n10152) );
  INV_X1 U12700 ( .A(n13724), .ZN(n11388) );
  AOI22_X1 U12701 ( .A1(n11388), .A2(n12016), .B1(n15017), .B2(
        P2_REG1_REG_2__SCAN_IN), .ZN(n10081) );
  OAI21_X1 U12702 ( .B1(n10152), .B2(n15017), .A(n10081), .ZN(P2_U3501) );
  INV_X1 U12703 ( .A(n10082), .ZN(n10123) );
  AOI22_X1 U12704 ( .A1(n10566), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n10083), .ZN(n10084) );
  OAI21_X1 U12705 ( .B1(n10123), .B2(n12610), .A(n10084), .ZN(P1_U3343) );
  XNOR2_X1 U12706 ( .A(n10428), .B(n11039), .ZN(n10085) );
  NAND2_X1 U12707 ( .A1(n10429), .A2(n13373), .ZN(n10086) );
  NAND2_X1 U12708 ( .A1(n10085), .A2(n10086), .ZN(n10136) );
  INV_X1 U12709 ( .A(n10085), .ZN(n10088) );
  INV_X1 U12710 ( .A(n10086), .ZN(n10087) );
  NAND2_X1 U12711 ( .A1(n10088), .A2(n10087), .ZN(n10089) );
  AND2_X1 U12712 ( .A1(n10089), .A2(n10136), .ZN(n10096) );
  INV_X1 U12713 ( .A(n10090), .ZN(n10092) );
  NAND2_X1 U12714 ( .A1(n10092), .A2(n10091), .ZN(n10093) );
  NAND2_X1 U12715 ( .A1(n10094), .A2(n10093), .ZN(n10095) );
  NAND2_X1 U12716 ( .A1(n10097), .A2(n13326), .ZN(n10100) );
  AOI22_X1 U12717 ( .A1(n12016), .A2(n13346), .B1(n13342), .B2(n10098), .ZN(
        n10099) );
  OAI211_X1 U12718 ( .C1(n10128), .C2(n10101), .A(n10100), .B(n10099), .ZN(
        P2_U3209) );
  INV_X1 U12719 ( .A(n10102), .ZN(n10103) );
  OAI222_X1 U12720 ( .A1(P3_U3151), .A2(n12833), .B1(n13217), .B2(n10104), 
        .C1(n13213), .C2(n10103), .ZN(P3_U3280) );
  XNOR2_X1 U12721 ( .A(n10269), .B(n11010), .ZN(n10107) );
  OAI211_X1 U12722 ( .C1(n10108), .C2(n10107), .A(n10261), .B(n14929), .ZN(
        n10121) );
  MUX2_X1 U12723 ( .A(n10109), .B(P2_REG1_REG_10__SCAN_IN), .S(n10269), .Z(
        n10113) );
  OR2_X1 U12724 ( .A1(n10110), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n10111) );
  NAND2_X1 U12725 ( .A1(n10112), .A2(n10111), .ZN(n10114) );
  AOI21_X1 U12726 ( .B1(n10113), .B2(n10114), .A(n14922), .ZN(n10119) );
  INV_X1 U12727 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n14562) );
  NAND2_X1 U12728 ( .A1(n14914), .A2(n10269), .ZN(n10117) );
  NOR2_X1 U12729 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10115), .ZN(n10997) );
  INV_X1 U12730 ( .A(n10997), .ZN(n10116) );
  OAI211_X1 U12731 ( .C1(n14562), .C2(n14932), .A(n10117), .B(n10116), .ZN(
        n10118) );
  AOI21_X1 U12732 ( .B1(n10119), .B2(n10271), .A(n10118), .ZN(n10120) );
  NAND2_X1 U12733 ( .A1(n10121), .A2(n10120), .ZN(P2_U3224) );
  INV_X1 U12734 ( .A(n14857), .ZN(n11094) );
  OAI222_X1 U12735 ( .A1(P2_U3088), .A2(n11094), .B1(n6551), .B2(n10123), .C1(
        n10122), .C2(n13780), .ZN(P2_U3315) );
  INV_X1 U12736 ( .A(n12722), .ZN(n12704) );
  AND2_X1 U12737 ( .A1(n15138), .A2(n10397), .ZN(n12415) );
  INV_X1 U12738 ( .A(n12415), .ZN(n12417) );
  AND2_X1 U12739 ( .A1(n12417), .A2(n10252), .ZN(n12386) );
  NOR2_X1 U12740 ( .A1(n12724), .A2(P3_U3151), .ZN(n10419) );
  INV_X1 U12741 ( .A(n10419), .ZN(n10124) );
  NAND2_X1 U12742 ( .A1(n10124), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n10126) );
  AOI22_X1 U12743 ( .A1(n12728), .A2(n15121), .B1(n10155), .B2(n12702), .ZN(
        n10125) );
  OAI211_X1 U12744 ( .C1(n12704), .C2(n12386), .A(n10126), .B(n10125), .ZN(
        P3_U3172) );
  INV_X1 U12745 ( .A(P3_DATAO_REG_20__SCAN_IN), .ZN(n15470) );
  NAND2_X1 U12746 ( .A1(n12529), .A2(P3_U3897), .ZN(n10127) );
  OAI21_X1 U12747 ( .B1(P3_U3897), .B2(n15470), .A(n10127), .ZN(P3_U3511) );
  INV_X1 U12748 ( .A(n13346), .ZN(n13334) );
  INV_X1 U12749 ( .A(n10128), .ZN(n10129) );
  NAND2_X1 U12750 ( .A1(n13342), .A2(n13496), .ZN(n13329) );
  INV_X1 U12751 ( .A(n13329), .ZN(n11876) );
  AOI22_X1 U12752 ( .A1(n10129), .A2(P2_REG3_REG_0__SCAN_IN), .B1(n11876), 
        .B2(n13374), .ZN(n10135) );
  NOR3_X1 U12753 ( .A1(n13603), .A2(n12002), .A3(n10130), .ZN(n10133) );
  INV_X1 U12754 ( .A(n10131), .ZN(n10132) );
  OAI21_X1 U12755 ( .B1(n10133), .B2(n10132), .A(n13326), .ZN(n10134) );
  OAI211_X1 U12756 ( .C1(n13334), .C2(n12003), .A(n10135), .B(n10134), .ZN(
        P2_U3204) );
  NAND2_X1 U12757 ( .A1(n10429), .A2(n13372), .ZN(n10313) );
  XNOR2_X1 U12758 ( .A(n10312), .B(n10313), .ZN(n10310) );
  XNOR2_X1 U12759 ( .A(n10311), .B(n10310), .ZN(n10141) );
  NAND2_X1 U12760 ( .A1(n13342), .A2(n13462), .ZN(n13328) );
  INV_X1 U12761 ( .A(n13328), .ZN(n11671) );
  AOI22_X1 U12762 ( .A1(n11671), .A2(n13373), .B1(n11876), .B2(n13371), .ZN(
        n10140) );
  NAND2_X1 U12763 ( .A1(n10137), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13344) );
  INV_X1 U12764 ( .A(n13344), .ZN(n13320) );
  INV_X1 U12765 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n15293) );
  OAI22_X1 U12766 ( .A1(n13334), .A2(n10946), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n15293), .ZN(n10138) );
  AOI21_X1 U12767 ( .B1(n13320), .B2(n15293), .A(n10138), .ZN(n10139) );
  OAI211_X1 U12768 ( .C1(n10141), .C2(n13348), .A(n10140), .B(n10139), .ZN(
        P2_U3190) );
  OAI21_X1 U12769 ( .B1(n10143), .B2(n12249), .A(n10142), .ZN(n10951) );
  INV_X1 U12770 ( .A(n10951), .ZN(n10147) );
  AOI222_X1 U12771 ( .A1(n13618), .A2(n10145), .B1(n13371), .B2(n13496), .C1(
        n13373), .C2(n13462), .ZN(n10947) );
  OAI211_X1 U12772 ( .C1(n10146), .C2(n10946), .A(n13603), .B(n10239), .ZN(
        n10945) );
  OAI211_X1 U12773 ( .C1(n13730), .C2(n10147), .A(n10947), .B(n10945), .ZN(
        n10176) );
  OAI22_X1 U12774 ( .A1(n13724), .A2(n10946), .B1(n15019), .B2(n10148), .ZN(
        n10149) );
  AOI21_X1 U12775 ( .B1(n10176), .B2(n15019), .A(n10149), .ZN(n10150) );
  INV_X1 U12776 ( .A(n10150), .ZN(P2_U3502) );
  AOI22_X1 U12777 ( .A1(n9616), .A2(n12016), .B1(n15005), .B2(
        P2_REG0_REG_2__SCAN_IN), .ZN(n10151) );
  OAI21_X1 U12778 ( .B1(n10152), .B2(n15005), .A(n10151), .ZN(P2_U3436) );
  NOR2_X1 U12779 ( .A1(n10153), .A2(n15143), .ZN(n10154) );
  INV_X1 U12780 ( .A(n15121), .ZN(n10414) );
  OAI22_X1 U12781 ( .A1(n12386), .A2(n10154), .B1(n10414), .B2(n13069), .ZN(
        n10394) );
  INV_X1 U12782 ( .A(n10394), .ZN(n10158) );
  INV_X1 U12783 ( .A(n13188), .ZN(n10156) );
  AOI22_X1 U12784 ( .A1(n10156), .A2(n10155), .B1(n15206), .B2(
        P3_REG0_REG_0__SCAN_IN), .ZN(n10157) );
  OAI21_X1 U12785 ( .B1(n10158), .B2(n15206), .A(n10157), .ZN(P3_U3390) );
  MUX2_X1 U12786 ( .A(n10399), .B(P1_REG1_REG_11__SCAN_IN), .S(n10402), .Z(
        n10163) );
  AOI21_X1 U12787 ( .B1(n10166), .B2(n10160), .A(n10159), .ZN(n14018) );
  MUX2_X1 U12788 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n10161), .S(n10167), .Z(
        n14017) );
  NAND2_X1 U12789 ( .A1(n14018), .A2(n14017), .ZN(n14016) );
  OAI21_X1 U12790 ( .B1(n14019), .B2(n10161), .A(n14016), .ZN(n10162) );
  NOR2_X1 U12791 ( .A1(n10162), .A2(n10163), .ZN(n10398) );
  AOI21_X1 U12792 ( .B1(n10163), .B2(n10162), .A(n10398), .ZN(n10174) );
  NOR2_X1 U12793 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n11549), .ZN(n10165) );
  NOR2_X1 U12794 ( .A1(n14744), .A2(n10400), .ZN(n10164) );
  AOI211_X1 U12795 ( .C1(n14719), .C2(P1_ADDR_REG_11__SCAN_IN), .A(n10165), 
        .B(n10164), .ZN(n10173) );
  NOR2_X1 U12796 ( .A1(n10166), .A2(n11025), .ZN(n14023) );
  MUX2_X1 U12797 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n11188), .S(n10167), .Z(
        n14022) );
  OAI21_X1 U12798 ( .B1(n14024), .B2(n14023), .A(n14022), .ZN(n14026) );
  NAND2_X1 U12799 ( .A1(n10167), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n10169) );
  MUX2_X1 U12800 ( .A(n11284), .B(P1_REG2_REG_11__SCAN_IN), .S(n10402), .Z(
        n10168) );
  AOI21_X1 U12801 ( .B1(n14026), .B2(n10169), .A(n10168), .ZN(n10401) );
  INV_X1 U12802 ( .A(n10401), .ZN(n10171) );
  NAND3_X1 U12803 ( .A1(n14026), .A2(n10169), .A3(n10168), .ZN(n10170) );
  NAND3_X1 U12804 ( .A1(n10171), .A2(n14059), .A3(n10170), .ZN(n10172) );
  OAI211_X1 U12805 ( .C1(n10174), .C2(n14040), .A(n10173), .B(n10172), .ZN(
        P1_U3254) );
  OAI22_X1 U12806 ( .A1(n13764), .A2(n10946), .B1(n15007), .B2(n9191), .ZN(
        n10175) );
  AOI21_X1 U12807 ( .B1(n10176), .B2(n15007), .A(n10175), .ZN(n10177) );
  INV_X1 U12808 ( .A(n10177), .ZN(P2_U3439) );
  NAND3_X1 U12809 ( .A1(n14766), .A2(n8429), .A3(n10178), .ZN(n10179) );
  AND2_X1 U12810 ( .A1(n10180), .A2(n10179), .ZN(n10186) );
  OAI21_X1 U12811 ( .B1(n8429), .B2(n10182), .A(n10181), .ZN(n10183) );
  NAND2_X1 U12812 ( .A1(n10183), .A2(n14783), .ZN(n10185) );
  INV_X1 U12813 ( .A(n10352), .ZN(n13883) );
  AOI22_X1 U12814 ( .A1(n14757), .A2(n13883), .B1(n13885), .B2(n14247), .ZN(
        n10184) );
  OAI211_X1 U12815 ( .C1(n10186), .C2(n14755), .A(n10185), .B(n10184), .ZN(
        n10514) );
  AOI211_X1 U12816 ( .C1(n13884), .C2(n14759), .A(n14793), .B(n10305), .ZN(
        n10516) );
  NOR2_X1 U12817 ( .A1(n10514), .A2(n10516), .ZN(n10451) );
  OAI22_X1 U12818 ( .A1(n14327), .A2(n10519), .B1(n14811), .B2(n9918), .ZN(
        n10187) );
  INV_X1 U12819 ( .A(n10187), .ZN(n10188) );
  OAI21_X1 U12820 ( .B1(n10451), .B2(n14809), .A(n10188), .ZN(P1_U3530) );
  INV_X1 U12821 ( .A(n14878), .ZN(n10191) );
  INV_X1 U12822 ( .A(n10189), .ZN(n10192) );
  OAI222_X1 U12823 ( .A1(P2_U3088), .A2(n10191), .B1(n6551), .B2(n10192), .C1(
        n10190), .C2(n13780), .ZN(P2_U3314) );
  INV_X1 U12824 ( .A(n10672), .ZN(n10676) );
  OAI222_X1 U12825 ( .A1(n14433), .A2(n15454), .B1(n12610), .B2(n10192), .C1(
        n10676), .C2(P1_U3086), .ZN(P1_U3342) );
  OAI22_X1 U12826 ( .A1(n13764), .A2(n10193), .B1(n15007), .B2(n9150), .ZN(
        n10194) );
  AOI21_X1 U12827 ( .B1(n15007), .B2(n10195), .A(n10194), .ZN(n10196) );
  INV_X1 U12828 ( .A(n10196), .ZN(P2_U3433) );
  INV_X1 U12829 ( .A(n10197), .ZN(n10199) );
  OAI21_X1 U12830 ( .B1(n9115), .B2(n10199), .A(n10198), .ZN(n10215) );
  NAND2_X1 U12831 ( .A1(n10199), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12586) );
  AND2_X1 U12832 ( .A1(n10200), .A2(n12586), .ZN(n10213) );
  OR2_X1 U12833 ( .A1(n10215), .A2(n10213), .ZN(n10208) );
  INV_X2 U12834 ( .A(P3_U3897), .ZN(n12745) );
  MUX2_X1 U12835 ( .A(n10208), .B(n12745), .S(n10201), .Z(n15100) );
  NOR2_X1 U12836 ( .A1(n10208), .A2(n10202), .ZN(n15023) );
  MUX2_X1 U12837 ( .A(n10859), .B(P3_REG2_REG_2__SCAN_IN), .S(n10892), .Z(
        n10207) );
  INV_X1 U12838 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n15495) );
  NOR2_X1 U12839 ( .A1(n15507), .A2(n15495), .ZN(n15022) );
  INV_X1 U12840 ( .A(n15022), .ZN(n10203) );
  NAND2_X1 U12841 ( .A1(n10204), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n10205) );
  NAND2_X1 U12842 ( .A1(n10329), .A2(n10205), .ZN(n10206) );
  NAND2_X1 U12843 ( .A1(n10207), .A2(n10206), .ZN(n10858) );
  OAI21_X1 U12844 ( .B1(n10207), .B2(n10206), .A(n10858), .ZN(n10234) );
  NOR2_X2 U12845 ( .A1(n10208), .A2(n10218), .ZN(n15109) );
  INV_X1 U12846 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n10225) );
  MUX2_X1 U12847 ( .A(n10225), .B(P3_REG1_REG_2__SCAN_IN), .S(n10892), .Z(
        n10211) );
  NAND2_X1 U12848 ( .A1(P3_REG1_REG_0__SCAN_IN), .A2(n8550), .ZN(n15020) );
  NAND2_X1 U12849 ( .A1(n10345), .A2(n15020), .ZN(n10209) );
  NAND2_X1 U12850 ( .A1(n10209), .A2(n7543), .ZN(n10332) );
  INV_X1 U12851 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n10331) );
  OR2_X1 U12852 ( .A1(n10332), .A2(n10331), .ZN(n10334) );
  NAND2_X1 U12853 ( .A1(n10334), .A2(n7543), .ZN(n10210) );
  NAND2_X1 U12854 ( .A1(n10211), .A2(n10210), .ZN(n10891) );
  OAI21_X1 U12855 ( .B1(n10211), .B2(n10210), .A(n10891), .ZN(n10212) );
  NAND2_X1 U12856 ( .A1(n15109), .A2(n10212), .ZN(n10217) );
  INV_X1 U12857 ( .A(n10213), .ZN(n10214) );
  AOI22_X1 U12858 ( .A1(n15106), .A2(P3_ADDR_REG_2__SCAN_IN), .B1(
        P3_REG3_REG_2__SCAN_IN), .B2(P3_U3151), .ZN(n10216) );
  NAND2_X1 U12859 ( .A1(n10217), .A2(n10216), .ZN(n10233) );
  MUX2_X1 U12860 ( .A(n10219), .B(n10331), .S(n13209), .Z(n10220) );
  INV_X1 U12861 ( .A(n10220), .ZN(n10222) );
  NAND2_X1 U12862 ( .A1(n10222), .A2(n10221), .ZN(n10223) );
  INV_X1 U12863 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n10224) );
  MUX2_X1 U12864 ( .A(n15495), .B(n10224), .S(n13209), .Z(n15025) );
  NAND2_X1 U12865 ( .A1(n15025), .A2(n15507), .ZN(n15034) );
  INV_X1 U12866 ( .A(n15034), .ZN(n10338) );
  NAND2_X1 U12867 ( .A1(n10337), .A2(n10338), .ZN(n10336) );
  MUX2_X1 U12868 ( .A(n10859), .B(n10225), .S(n13209), .Z(n10226) );
  NAND2_X1 U12869 ( .A1(n10226), .A2(n10892), .ZN(n15038) );
  INV_X1 U12870 ( .A(n10226), .ZN(n10227) );
  NAND2_X1 U12871 ( .A1(n10227), .A2(n7199), .ZN(n10228) );
  NAND2_X1 U12872 ( .A1(n15038), .A2(n10228), .ZN(n10229) );
  INV_X1 U12873 ( .A(n15042), .ZN(n10231) );
  NAND2_X1 U12874 ( .A1(P3_U3897), .A2(n13205), .ZN(n15102) );
  AOI21_X1 U12875 ( .B1(n10231), .B2(n10230), .A(n15102), .ZN(n10232) );
  AOI211_X1 U12876 ( .C1(n15023), .C2(n10234), .A(n10233), .B(n10232), .ZN(
        n10235) );
  OAI21_X1 U12877 ( .B1(n7199), .B2(n15100), .A(n10235), .ZN(P3_U3184) );
  OAI21_X1 U12878 ( .B1(n10237), .B2(n10240), .A(n10236), .ZN(n10608) );
  INV_X1 U12879 ( .A(n10664), .ZN(n10238) );
  AOI211_X1 U12880 ( .C1(n12025), .C2(n10239), .A(n10574), .B(n10238), .ZN(
        n10618) );
  XNOR2_X1 U12881 ( .A(n10241), .B(n10240), .ZN(n10242) );
  AOI22_X1 U12882 ( .A1(n13462), .A2(n13372), .B1(n13496), .B2(n13370), .ZN(
        n10323) );
  OAI21_X1 U12883 ( .B1(n10242), .B2(n13600), .A(n10323), .ZN(n10611) );
  AOI211_X1 U12884 ( .C1(n14983), .C2(n10608), .A(n10618), .B(n10611), .ZN(
        n10248) );
  INV_X1 U12885 ( .A(n12025), .ZN(n12029) );
  OAI22_X1 U12886 ( .A1(n13724), .A2(n12029), .B1(n15019), .B2(n9206), .ZN(
        n10243) );
  INV_X1 U12887 ( .A(n10243), .ZN(n10244) );
  OAI21_X1 U12888 ( .B1(n10248), .B2(n15017), .A(n10244), .ZN(P2_U3503) );
  INV_X1 U12889 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10245) );
  OAI22_X1 U12890 ( .A1(n13764), .A2(n12029), .B1(n15007), .B2(n10245), .ZN(
        n10246) );
  INV_X1 U12891 ( .A(n10246), .ZN(n10247) );
  OAI21_X1 U12892 ( .B1(n10248), .B2(n15005), .A(n10247), .ZN(P2_U3442) );
  AOI222_X1 U12893 ( .A1(n10249), .A2(n13202), .B1(n12837), .B2(
        P3_STATE_REG_SCAN_IN), .C1(SI_16_), .C2(n13200), .ZN(n10250) );
  INV_X1 U12894 ( .A(n10250), .ZN(P3_U3279) );
  INV_X1 U12895 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n10260) );
  NAND3_X1 U12896 ( .A1(n15142), .A2(n10252), .A3(n10251), .ZN(n10253) );
  OAI211_X1 U12897 ( .C1(n10255), .C2(n15141), .A(n10254), .B(n10253), .ZN(
        n10256) );
  NAND2_X1 U12898 ( .A1(n10256), .A2(n12722), .ZN(n10259) );
  OAI22_X1 U12899 ( .A1(n9042), .A2(n12726), .B1(n12731), .B2(n8551), .ZN(
        n10257) );
  AOI21_X1 U12900 ( .B1(n12728), .B2(n15137), .A(n10257), .ZN(n10258) );
  OAI211_X1 U12901 ( .C1(n10419), .C2(n10260), .A(n10259), .B(n10258), .ZN(
        P3_U3162) );
  XNOR2_X1 U12902 ( .A(n11089), .B(P2_REG2_REG_11__SCAN_IN), .ZN(n10264) );
  NOR2_X1 U12903 ( .A1(n10263), .A2(n10264), .ZN(n11082) );
  AOI21_X1 U12904 ( .B1(n10264), .B2(n10263), .A(n11082), .ZN(n10277) );
  INV_X1 U12905 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n10267) );
  NAND2_X1 U12906 ( .A1(n14914), .A2(n11089), .ZN(n10266) );
  NAND2_X1 U12907 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(P2_U3088), .ZN(n10265)
         );
  OAI211_X1 U12908 ( .C1(n10267), .C2(n14932), .A(n10266), .B(n10265), .ZN(
        n10268) );
  INV_X1 U12909 ( .A(n10268), .ZN(n10276) );
  NAND2_X1 U12910 ( .A1(n10269), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n10270) );
  NAND2_X1 U12911 ( .A1(n10271), .A2(n10270), .ZN(n10274) );
  INV_X1 U12912 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n10272) );
  MUX2_X1 U12913 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n10272), .S(n11089), .Z(
        n10273) );
  NAND2_X1 U12914 ( .A1(n10274), .A2(n10273), .ZN(n11091) );
  OAI211_X1 U12915 ( .C1(n10274), .C2(n10273), .A(n11091), .B(n14846), .ZN(
        n10275) );
  OAI211_X1 U12916 ( .C1(n10277), .C2(n14907), .A(n10276), .B(n10275), .ZN(
        P2_U3225) );
  INV_X1 U12917 ( .A(n10278), .ZN(n10280) );
  INV_X1 U12918 ( .A(n10497), .ZN(n10279) );
  AOI21_X1 U12919 ( .B1(n10280), .B2(n10287), .A(n10279), .ZN(n10647) );
  INV_X1 U12920 ( .A(n10307), .ZN(n10281) );
  AOI211_X1 U12921 ( .C1(n10631), .C2(n10281), .A(n14793), .B(n6673), .ZN(
        n10644) );
  OR2_X1 U12922 ( .A1(n14276), .A2(n7733), .ZN(n10283) );
  NAND2_X1 U12923 ( .A1(n14247), .A2(n13937), .ZN(n10282) );
  AND2_X1 U12924 ( .A1(n10283), .A2(n10282), .ZN(n10637) );
  INV_X1 U12925 ( .A(n10637), .ZN(n10284) );
  NOR2_X1 U12926 ( .A1(n10644), .A2(n10284), .ZN(n10289) );
  OAI21_X1 U12927 ( .B1(n10287), .B2(n10286), .A(n10285), .ZN(n10288) );
  NAND2_X1 U12928 ( .A1(n10288), .A2(n14783), .ZN(n10638) );
  OAI211_X1 U12929 ( .C1(n10647), .C2(n14755), .A(n10289), .B(n10638), .ZN(
        n10461) );
  OAI22_X1 U12930 ( .A1(n14327), .A2(n10642), .B1(n14811), .B2(n9922), .ZN(
        n10290) );
  AOI21_X1 U12931 ( .B1(n10461), .B2(n14811), .A(n10290), .ZN(n10291) );
  INV_X1 U12932 ( .A(n10291), .ZN(P1_U3532) );
  INV_X1 U12933 ( .A(n14580), .ZN(n12865) );
  INV_X1 U12934 ( .A(SI_17_), .ZN(n10294) );
  INV_X1 U12935 ( .A(n10292), .ZN(n10293) );
  OAI222_X1 U12936 ( .A1(P3_U3151), .A2(n12865), .B1(n13217), .B2(n10294), 
        .C1(n13213), .C2(n10293), .ZN(P3_U3278) );
  OAI21_X1 U12937 ( .B1(n10297), .B2(n10296), .A(n10295), .ZN(n10304) );
  OAI22_X1 U12938 ( .A1(n10493), .A2(n14770), .B1(n14276), .B2(n14771), .ZN(
        n10303) );
  OAI21_X1 U12939 ( .B1(n10300), .B2(n10299), .A(n10298), .ZN(n10301) );
  AND2_X1 U12940 ( .A1(n10301), .A2(n14803), .ZN(n10302) );
  AOI211_X1 U12941 ( .C1(n14783), .C2(n10304), .A(n10303), .B(n10302), .ZN(
        n10520) );
  NOR2_X1 U12942 ( .A1(n10305), .A2(n7734), .ZN(n10306) );
  OR3_X1 U12943 ( .A1(n10307), .A2(n10306), .A3(n14793), .ZN(n10522) );
  NAND2_X1 U12944 ( .A1(n10520), .A2(n10522), .ZN(n10464) );
  OAI22_X1 U12945 ( .A1(n14327), .A2(n7734), .B1(n14811), .B2(n9920), .ZN(
        n10308) );
  AOI21_X1 U12946 ( .B1(n10464), .B2(n14811), .A(n10308), .ZN(n10309) );
  INV_X1 U12947 ( .A(n10309), .ZN(P1_U3531) );
  INV_X1 U12948 ( .A(n10312), .ZN(n10315) );
  INV_X1 U12949 ( .A(n10313), .ZN(n10314) );
  NAND2_X1 U12950 ( .A1(n10315), .A2(n10314), .ZN(n10436) );
  AND2_X1 U12951 ( .A1(n10440), .A2(n10436), .ZN(n10321) );
  XNOR2_X1 U12952 ( .A(n13282), .B(n12025), .ZN(n10319) );
  INV_X1 U12953 ( .A(n10319), .ZN(n10317) );
  AND2_X1 U12954 ( .A1(n10429), .A2(n13371), .ZN(n10318) );
  INV_X1 U12955 ( .A(n10318), .ZN(n10316) );
  NAND2_X1 U12956 ( .A1(n10317), .A2(n10316), .ZN(n10468) );
  NAND2_X1 U12957 ( .A1(n10319), .A2(n10318), .ZN(n10435) );
  AND2_X1 U12958 ( .A1(n10468), .A2(n10435), .ZN(n10320) );
  NAND2_X1 U12959 ( .A1(n10321), .A2(n10320), .ZN(n10470) );
  OAI21_X1 U12960 ( .B1(n10321), .B2(n10320), .A(n10470), .ZN(n10322) );
  NAND2_X1 U12961 ( .A1(n10322), .A2(n13326), .ZN(n10326) );
  INV_X1 U12962 ( .A(n13342), .ZN(n13318) );
  NAND2_X1 U12963 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3088), .ZN(n14839) );
  OAI21_X1 U12964 ( .B1(n13318), .B2(n10323), .A(n14839), .ZN(n10324) );
  AOI21_X1 U12965 ( .B1(n12025), .B2(n13346), .A(n10324), .ZN(n10325) );
  OAI211_X1 U12966 ( .C1(n13344), .C2(n10616), .A(n10326), .B(n10325), .ZN(
        P2_U3202) );
  INV_X1 U12967 ( .A(n15100), .ZN(n15031) );
  NAND2_X1 U12968 ( .A1(n10327), .A2(n10219), .ZN(n10328) );
  NAND2_X1 U12969 ( .A1(n10329), .A2(n10328), .ZN(n10330) );
  NAND2_X1 U12970 ( .A1(n15023), .A2(n10330), .ZN(n10343) );
  AOI22_X1 U12971 ( .A1(n15106), .A2(P3_ADDR_REG_1__SCAN_IN), .B1(
        P3_REG3_REG_1__SCAN_IN), .B2(P3_U3151), .ZN(n10342) );
  NAND2_X1 U12972 ( .A1(n10332), .A2(n10331), .ZN(n10333) );
  NAND2_X1 U12973 ( .A1(n10334), .A2(n10333), .ZN(n10335) );
  NAND2_X1 U12974 ( .A1(n15109), .A2(n10335), .ZN(n10341) );
  OAI21_X1 U12975 ( .B1(n10338), .B2(n10337), .A(n10336), .ZN(n10339) );
  INV_X1 U12976 ( .A(n15102), .ZN(n15085) );
  NAND2_X1 U12977 ( .A1(n10339), .A2(n15085), .ZN(n10340) );
  NAND4_X1 U12978 ( .A1(n10343), .A2(n10342), .A3(n10341), .A4(n10340), .ZN(
        n10344) );
  AOI21_X1 U12979 ( .B1(n10345), .B2(n15031), .A(n10344), .ZN(n10346) );
  INV_X1 U12980 ( .A(n10346), .ZN(P3_U3183) );
  NOR2_X1 U12981 ( .A1(n15222), .A2(n10224), .ZN(n10347) );
  AOI21_X1 U12982 ( .B1(n10394), .B2(n15222), .A(n10347), .ZN(n10348) );
  OAI21_X1 U12983 ( .B1(n10397), .B2(n13138), .A(n10348), .ZN(P3_U3459) );
  OAI22_X1 U12984 ( .A1(n11938), .A2(n7733), .B1(n7734), .B2(n11939), .ZN(
        n10623) );
  NAND2_X1 U12985 ( .A1(n13885), .A2(n10626), .ZN(n10350) );
  NAND2_X1 U12986 ( .A1(n11980), .A2(n10379), .ZN(n10349) );
  NAND2_X1 U12987 ( .A1(n10350), .A2(n10349), .ZN(n10351) );
  XNOR2_X1 U12988 ( .A(n10351), .B(n11149), .ZN(n10622) );
  XNOR2_X1 U12989 ( .A(n10623), .B(n10622), .ZN(n10374) );
  NAND2_X1 U12990 ( .A1(n13883), .A2(n10626), .ZN(n10353) );
  OAI22_X1 U12991 ( .A1(n10354), .A2(n10352), .B1(n14792), .B2(n11939), .ZN(
        n10358) );
  INV_X1 U12992 ( .A(n10358), .ZN(n10355) );
  NAND2_X1 U12993 ( .A1(n10358), .A2(n10357), .ZN(n10359) );
  NAND2_X1 U12994 ( .A1(n10362), .A2(n10361), .ZN(n13805) );
  NAND2_X1 U12995 ( .A1(n13803), .A2(n13805), .ZN(n13804) );
  NAND2_X1 U12996 ( .A1(n10626), .A2(n13808), .ZN(n10365) );
  NAND2_X1 U12997 ( .A1(n11980), .A2(n13884), .ZN(n10364) );
  NAND2_X1 U12998 ( .A1(n10365), .A2(n10364), .ZN(n10366) );
  OAI22_X1 U12999 ( .A1(n11938), .A2(n14771), .B1(n10519), .B2(n11939), .ZN(
        n10369) );
  XNOR2_X1 U13000 ( .A(n10367), .B(n10369), .ZN(n13879) );
  NAND2_X1 U13001 ( .A1(n13878), .A2(n13879), .ZN(n13876) );
  INV_X1 U13002 ( .A(n10367), .ZN(n10368) );
  OR2_X1 U13003 ( .A1(n10369), .A2(n10368), .ZN(n10370) );
  INV_X1 U13004 ( .A(n10374), .ZN(n10371) );
  INV_X1 U13005 ( .A(n10625), .ZN(n10372) );
  AOI211_X1 U13006 ( .C1(n10374), .C2(n10373), .A(n14674), .B(n10372), .ZN(
        n10383) );
  NAND2_X1 U13007 ( .A1(n10376), .A2(n10375), .ZN(n10377) );
  NAND2_X1 U13008 ( .A1(n10377), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10378) );
  INV_X1 U13009 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n13955) );
  AOI22_X1 U13010 ( .A1(n14665), .A2(n13938), .B1(n14679), .B2(n10379), .ZN(
        n10381) );
  AOI22_X1 U13011 ( .A1(n13900), .A2(n13808), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(P1_U3086), .ZN(n10380) );
  OAI211_X1 U13012 ( .C1(n14684), .C2(P1_REG3_REG_3__SCAN_IN), .A(n10381), .B(
        n10380), .ZN(n10382) );
  OR2_X1 U13013 ( .A1(n10383), .A2(n10382), .ZN(P1_U3218) );
  AND2_X1 U13014 ( .A1(n9115), .A2(n10384), .ZN(n10389) );
  NAND2_X1 U13015 ( .A1(n10385), .A2(n10388), .ZN(n10387) );
  OAI211_X1 U13016 ( .C1(n10389), .C2(n10388), .A(n10387), .B(n10386), .ZN(
        n10392) );
  INV_X1 U13017 ( .A(n10392), .ZN(n10391) );
  NOR2_X1 U13018 ( .A1(n15200), .A2(n15134), .ZN(n10390) );
  NAND2_X1 U13019 ( .A1(n10391), .A2(n10390), .ZN(n14613) );
  NOR2_X1 U13020 ( .A1(n15132), .A2(n15495), .ZN(n10393) );
  AOI21_X1 U13021 ( .B1(n10394), .B2(n15132), .A(n10393), .ZN(n10396) );
  NAND2_X1 U13022 ( .A1(n15150), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n10395) );
  OAI211_X1 U13023 ( .C1(n14613), .C2(n10397), .A(n10396), .B(n10395), .ZN(
        P3_U3233) );
  XNOR2_X1 U13024 ( .A(n10566), .B(P1_REG1_REG_12__SCAN_IN), .ZN(n10561) );
  AOI21_X1 U13025 ( .B1(n10400), .B2(n10399), .A(n10398), .ZN(n10562) );
  XOR2_X1 U13026 ( .A(n10561), .B(n10562), .Z(n10410) );
  MUX2_X1 U13027 ( .A(P1_REG2_REG_12__SCAN_IN), .B(n11472), .S(n10566), .Z(
        n10404) );
  AOI21_X1 U13028 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n10402), .A(n10401), 
        .ZN(n10403) );
  NAND2_X1 U13029 ( .A1(n10403), .A2(n10404), .ZN(n10565) );
  OAI21_X1 U13030 ( .B1(n10404), .B2(n10403), .A(n10565), .ZN(n10408) );
  INV_X1 U13031 ( .A(n10566), .ZN(n10406) );
  AOI22_X1 U13032 ( .A1(n14719), .A2(P1_ADDR_REG_12__SCAN_IN), .B1(
        P1_REG3_REG_12__SCAN_IN), .B2(P1_U3086), .ZN(n10405) );
  OAI21_X1 U13033 ( .B1(n10406), .B2(n14744), .A(n10405), .ZN(n10407) );
  AOI21_X1 U13034 ( .B1(n10408), .B2(n14059), .A(n10407), .ZN(n10409) );
  OAI21_X1 U13035 ( .B1(n10410), .B2(n14040), .A(n10409), .ZN(P1_U3255) );
  INV_X1 U13036 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n10418) );
  OAI21_X1 U13037 ( .B1(n10412), .B2(n10411), .A(n10481), .ZN(n10413) );
  NAND2_X1 U13038 ( .A1(n10413), .A2(n12722), .ZN(n10417) );
  OAI22_X1 U13039 ( .A1(n10414), .A2(n12726), .B1(n12731), .B2(n15117), .ZN(
        n10415) );
  AOI21_X1 U13040 ( .B1(n12728), .B2(n15120), .A(n10415), .ZN(n10416) );
  OAI211_X1 U13041 ( .C1(n10419), .C2(n10418), .A(n10417), .B(n10416), .ZN(
        P3_U3177) );
  INV_X1 U13042 ( .A(n10420), .ZN(n10423) );
  INV_X1 U13043 ( .A(n11561), .ZN(n11336) );
  OAI222_X1 U13044 ( .A1(n14433), .A2(n10421), .B1(n12610), .B2(n10423), .C1(
        n11336), .C2(P1_U3086), .ZN(P1_U3339) );
  INV_X1 U13045 ( .A(n14900), .ZN(n10422) );
  OAI222_X1 U13046 ( .A1(n13768), .A2(n10424), .B1(n6551), .B2(n10423), .C1(
        n10422), .C2(P2_U3088), .ZN(P2_U3311) );
  INV_X1 U13047 ( .A(n10425), .ZN(n10426) );
  OAI222_X1 U13048 ( .A1(P3_U3151), .A2(n12856), .B1(n13217), .B2(n10427), 
        .C1(n13213), .C2(n10426), .ZN(P3_U3277) );
  INV_X2 U13049 ( .A(n10428), .ZN(n13236) );
  XNOR2_X1 U13050 ( .A(n12048), .B(n13236), .ZN(n10577) );
  NAND2_X1 U13051 ( .A1(n10574), .A2(n13369), .ZN(n10578) );
  NAND2_X1 U13052 ( .A1(n10429), .A2(n13370), .ZN(n10431) );
  NAND2_X1 U13053 ( .A1(n10430), .A2(n10431), .ZN(n10441) );
  INV_X1 U13054 ( .A(n10430), .ZN(n10433) );
  INV_X1 U13055 ( .A(n10431), .ZN(n10432) );
  NAND2_X1 U13056 ( .A1(n10433), .A2(n10432), .ZN(n10434) );
  NAND2_X1 U13057 ( .A1(n10436), .A2(n10435), .ZN(n10437) );
  NOR2_X1 U13058 ( .A1(n10469), .A2(n10437), .ZN(n10439) );
  NOR2_X1 U13059 ( .A1(n10469), .A2(n10468), .ZN(n10438) );
  XOR2_X1 U13060 ( .A(n10575), .B(n10576), .Z(n10447) );
  NAND2_X1 U13061 ( .A1(n13496), .A2(n13368), .ZN(n10443) );
  NAND2_X1 U13062 ( .A1(n13462), .A2(n13370), .ZN(n10442) );
  NAND2_X1 U13063 ( .A1(n10443), .A2(n10442), .ZN(n10847) );
  AOI22_X1 U13064 ( .A1(n13342), .A2(n10847), .B1(P2_REG3_REG_6__SCAN_IN), 
        .B2(P2_U3088), .ZN(n10445) );
  NAND2_X1 U13065 ( .A1(n13346), .A2(n12048), .ZN(n10444) );
  OAI211_X1 U13066 ( .C1(n13344), .C2(n10849), .A(n10445), .B(n10444), .ZN(
        n10446) );
  AOI21_X1 U13067 ( .B1(n10447), .B2(n13326), .A(n10446), .ZN(n10448) );
  INV_X1 U13068 ( .A(n10448), .ZN(P2_U3211) );
  OAI22_X1 U13069 ( .A1(n14411), .A2(n10519), .B1(n14806), .B2(n7698), .ZN(
        n10449) );
  INV_X1 U13070 ( .A(n10449), .ZN(n10450) );
  OAI21_X1 U13071 ( .B1(n10451), .B2(n14804), .A(n10450), .ZN(P1_U3465) );
  INV_X1 U13072 ( .A(n10452), .ZN(n10454) );
  INV_X1 U13073 ( .A(n11319), .ZN(n11325) );
  OAI222_X1 U13074 ( .A1(n14433), .A2(n10453), .B1(n12610), .B2(n10454), .C1(
        n11325), .C2(P1_U3086), .ZN(P1_U3341) );
  OAI222_X1 U13075 ( .A1(n13768), .A2(n10455), .B1(n6551), .B2(n10454), .C1(
        n11088), .C2(P2_U3088), .ZN(P2_U3313) );
  INV_X1 U13076 ( .A(n10456), .ZN(n10507) );
  AOI22_X1 U13077 ( .A1(n14913), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n10457), .ZN(n10458) );
  OAI21_X1 U13078 ( .B1(n10507), .B2(n6551), .A(n10458), .ZN(P2_U3310) );
  INV_X1 U13079 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10459) );
  OAI22_X1 U13080 ( .A1(n14411), .A2(n10642), .B1(n14806), .B2(n10459), .ZN(
        n10460) );
  AOI21_X1 U13081 ( .B1(n10461), .B2(n14806), .A(n10460), .ZN(n10462) );
  INV_X1 U13082 ( .A(n10462), .ZN(P1_U3471) );
  OAI22_X1 U13083 ( .A1(n14411), .A2(n7734), .B1(n14806), .B2(n7720), .ZN(
        n10463) );
  AOI21_X1 U13084 ( .B1(n10464), .B2(n14806), .A(n10463), .ZN(n10465) );
  INV_X1 U13085 ( .A(n10465), .ZN(P1_U3468) );
  AOI22_X1 U13086 ( .A1(n13462), .A2(n13371), .B1(n13496), .B2(n13369), .ZN(
        n10660) );
  NAND2_X1 U13087 ( .A1(n13346), .A2(n6721), .ZN(n10466) );
  OAI211_X1 U13088 ( .C1(n13318), .C2(n10660), .A(n10467), .B(n10466), .ZN(
        n10474) );
  NAND3_X1 U13089 ( .A1(n10470), .A2(n10469), .A3(n10468), .ZN(n10472) );
  AOI21_X1 U13090 ( .B1(n10472), .B2(n10471), .A(n13348), .ZN(n10473) );
  AOI211_X1 U13091 ( .C1(n13320), .C2(n10665), .A(n10474), .B(n10473), .ZN(
        n10475) );
  INV_X1 U13092 ( .A(n10475), .ZN(P2_U3199) );
  OAI222_X1 U13093 ( .A1(n13213), .A2(n10477), .B1(n13217), .B2(n10476), .C1(
        P3_U3151), .C2(n12859), .ZN(P3_U3276) );
  INV_X1 U13094 ( .A(n10478), .ZN(n10483) );
  AOI21_X1 U13095 ( .B1(n10481), .B2(n10480), .A(n10479), .ZN(n10482) );
  NOR3_X1 U13096 ( .A1(n10483), .A2(n10482), .A3(n12704), .ZN(n10490) );
  NAND2_X1 U13097 ( .A1(n12724), .A2(n15459), .ZN(n10488) );
  INV_X1 U13098 ( .A(n12726), .ZN(n12709) );
  NOR2_X1 U13099 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15459), .ZN(n15043) );
  AOI21_X1 U13100 ( .B1(n12709), .B2(n15137), .A(n15043), .ZN(n10487) );
  NAND2_X1 U13101 ( .A1(n12728), .A2(n12744), .ZN(n10486) );
  NAND2_X1 U13102 ( .A1(n12702), .A2(n10484), .ZN(n10485) );
  NAND4_X1 U13103 ( .A1(n10488), .A2(n10487), .A3(n10486), .A4(n10485), .ZN(
        n10489) );
  OR2_X1 U13104 ( .A1(n10490), .A2(n10489), .ZN(P3_U3158) );
  OAI21_X1 U13105 ( .B1(n10496), .B2(n10492), .A(n10491), .ZN(n10501) );
  OAI22_X1 U13106 ( .A1(n10493), .A2(n14276), .B1(n14770), .B2(n10597), .ZN(
        n10500) );
  NAND3_X1 U13107 ( .A1(n10497), .A2(n10496), .A3(n10495), .ZN(n10498) );
  AOI21_X1 U13108 ( .B1(n10494), .B2(n10498), .A(n14755), .ZN(n10499) );
  AOI211_X1 U13109 ( .C1(n14783), .C2(n10501), .A(n10500), .B(n10499), .ZN(
        n10746) );
  INV_X1 U13110 ( .A(n14793), .ZN(n14365) );
  OAI211_X1 U13111 ( .C1(n6673), .C2(n7016), .A(n14365), .B(n10548), .ZN(
        n10741) );
  NAND2_X1 U13112 ( .A1(n10746), .A2(n10741), .ZN(n10505) );
  OAI22_X1 U13113 ( .A1(n14327), .A2(n7016), .B1(n14811), .B2(n9923), .ZN(
        n10502) );
  AOI21_X1 U13114 ( .B1(n10505), .B2(n14811), .A(n10502), .ZN(n10503) );
  INV_X1 U13115 ( .A(n10503), .ZN(P1_U3533) );
  OAI22_X1 U13116 ( .A1(n14411), .A2(n7016), .B1(n14806), .B2(n7762), .ZN(
        n10504) );
  AOI21_X1 U13117 ( .B1(n10505), .B2(n14806), .A(n10504), .ZN(n10506) );
  INV_X1 U13118 ( .A(n10506), .ZN(P1_U3474) );
  INV_X1 U13119 ( .A(n14039), .ZN(n14031) );
  OAI222_X1 U13120 ( .A1(n14433), .A2(n10508), .B1(n12610), .B2(n10507), .C1(
        n14031), .C2(P1_U3086), .ZN(P1_U3338) );
  INV_X1 U13121 ( .A(n10509), .ZN(n10512) );
  INV_X1 U13122 ( .A(n10510), .ZN(n10511) );
  NAND2_X1 U13123 ( .A1(n10512), .A2(n10511), .ZN(n12596) );
  INV_X2 U13124 ( .A(n14281), .ZN(n14256) );
  INV_X1 U13125 ( .A(n14772), .ZN(n10513) );
  NAND2_X1 U13126 ( .A1(n14256), .A2(n10513), .ZN(n14271) );
  MUX2_X1 U13127 ( .A(n10514), .B(P1_REG2_REG_2__SCAN_IN), .S(n14281), .Z(
        n10515) );
  INV_X1 U13128 ( .A(n10515), .ZN(n10518) );
  INV_X1 U13129 ( .A(n14777), .ZN(n14786) );
  AOI22_X1 U13130 ( .A1(n14284), .A2(n10516), .B1(P1_REG3_REG_2__SCAN_IN), 
        .B2(n14786), .ZN(n10517) );
  OAI211_X1 U13131 ( .C1(n10519), .C2(n14271), .A(n10518), .B(n10517), .ZN(
        P1_U3291) );
  MUX2_X1 U13132 ( .A(n10521), .B(n10520), .S(n14256), .Z(n10525) );
  INV_X1 U13133 ( .A(n10522), .ZN(n10523) );
  AOI22_X1 U13134 ( .A1(n14284), .A2(n10523), .B1(n14786), .B2(n13955), .ZN(
        n10524) );
  OAI211_X1 U13135 ( .C1(n7734), .C2(n14271), .A(n10525), .B(n10524), .ZN(
        P1_U3290) );
  NAND4_X1 U13136 ( .A1(n10527), .A2(n14953), .A3(n14952), .A4(n10526), .ZN(
        n10528) );
  AND2_X2 U13137 ( .A1(n13535), .A2(n10528), .ZN(n14947) );
  INV_X1 U13138 ( .A(n11997), .ZN(n10609) );
  NOR2_X1 U13139 ( .A1(n14947), .A2(n10609), .ZN(n13638) );
  INV_X1 U13140 ( .A(n13638), .ZN(n11317) );
  OR2_X1 U13141 ( .A1(n13375), .A2(n12002), .ZN(n10531) );
  NAND2_X1 U13142 ( .A1(n10532), .A2(n10531), .ZN(n14960) );
  NAND2_X1 U13143 ( .A1(n10533), .A2(n12002), .ZN(n14958) );
  AOI21_X1 U13144 ( .B1(n13600), .B2(n13624), .A(n14960), .ZN(n10534) );
  AOI21_X1 U13145 ( .B1(n13496), .B2(n13374), .A(n10534), .ZN(n14959) );
  OAI21_X1 U13146 ( .B1(n10530), .B2(n14958), .A(n14959), .ZN(n10535) );
  NAND2_X1 U13147 ( .A1(n10535), .A2(n13602), .ZN(n10537) );
  INV_X1 U13148 ( .A(n13535), .ZN(n14936) );
  AOI22_X1 U13149 ( .A1(n14947), .A2(P2_REG2_REG_0__SCAN_IN), .B1(n14936), 
        .B2(P2_REG3_REG_0__SCAN_IN), .ZN(n10536) );
  OAI211_X1 U13150 ( .C1(n11317), .C2(n14960), .A(n10537), .B(n10536), .ZN(
        P2_U3265) );
  OAI21_X1 U13151 ( .B1(n10543), .B2(n10539), .A(n10538), .ZN(n10547) );
  OAI22_X1 U13152 ( .A1(n10540), .A2(n14276), .B1(n14770), .B2(n10961), .ZN(
        n10546) );
  NAND3_X1 U13153 ( .A1(n10494), .A2(n10543), .A3(n10542), .ZN(n10544) );
  AOI21_X1 U13154 ( .B1(n10541), .B2(n10544), .A(n14755), .ZN(n10545) );
  AOI211_X1 U13155 ( .C1(n14783), .C2(n10547), .A(n10546), .B(n10545), .ZN(
        n10747) );
  NAND2_X1 U13156 ( .A1(n10548), .A2(n10767), .ZN(n10549) );
  NAND2_X1 U13157 ( .A1(n10549), .A2(n14365), .ZN(n10550) );
  OR2_X1 U13158 ( .A1(n10601), .A2(n10550), .ZN(n10752) );
  NAND2_X1 U13159 ( .A1(n10747), .A2(n10752), .ZN(n10555) );
  OAI22_X1 U13160 ( .A1(n14327), .A2(n7015), .B1(n14811), .B2(n9924), .ZN(
        n10551) );
  AOI21_X1 U13161 ( .B1(n10555), .B2(n14811), .A(n10551), .ZN(n10552) );
  INV_X1 U13162 ( .A(n10552), .ZN(P1_U3534) );
  INV_X1 U13163 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10553) );
  OAI22_X1 U13164 ( .A1(n14411), .A2(n7015), .B1(n14806), .B2(n10553), .ZN(
        n10554) );
  AOI21_X1 U13165 ( .B1(n10555), .B2(n14806), .A(n10554), .ZN(n10556) );
  INV_X1 U13166 ( .A(n10556), .ZN(P1_U3477) );
  INV_X1 U13167 ( .A(n11327), .ZN(n14745) );
  INV_X1 U13168 ( .A(n10557), .ZN(n10560) );
  OAI222_X1 U13169 ( .A1(P1_U3086), .A2(n14745), .B1(n12610), .B2(n10560), 
        .C1(n10558), .C2(n14433), .ZN(P1_U3340) );
  OAI222_X1 U13170 ( .A1(P2_U3088), .A2(n13404), .B1(n6551), .B2(n10560), .C1(
        n10559), .C2(n13780), .ZN(P2_U3312) );
  XNOR2_X1 U13171 ( .A(n10672), .B(P1_REG1_REG_13__SCAN_IN), .ZN(n10564) );
  OAI22_X1 U13172 ( .A1(n10562), .A2(n10561), .B1(P1_REG1_REG_12__SCAN_IN), 
        .B2(n10566), .ZN(n10563) );
  NOR2_X1 U13173 ( .A1(n10563), .A2(n10564), .ZN(n10671) );
  AOI211_X1 U13174 ( .C1(n10564), .C2(n10563), .A(n14040), .B(n10671), .ZN(
        n10573) );
  OAI21_X1 U13175 ( .B1(n10566), .B2(P1_REG2_REG_12__SCAN_IN), .A(n10565), 
        .ZN(n10568) );
  INV_X1 U13176 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n10675) );
  MUX2_X1 U13177 ( .A(n10675), .B(P1_REG2_REG_13__SCAN_IN), .S(n10672), .Z(
        n10567) );
  NOR2_X1 U13178 ( .A1(n10568), .A2(n10567), .ZN(n10682) );
  AOI211_X1 U13179 ( .C1(n10568), .C2(n10567), .A(n14746), .B(n10682), .ZN(
        n10572) );
  NAND2_X1 U13180 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n11740)
         );
  INV_X1 U13181 ( .A(n11740), .ZN(n10569) );
  AOI21_X1 U13182 ( .B1(n14719), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n10569), 
        .ZN(n10570) );
  OAI21_X1 U13183 ( .B1(n14744), .B2(n10676), .A(n10570), .ZN(n10571) );
  OR3_X1 U13184 ( .A1(n10573), .A2(n10572), .A3(n10571), .ZN(P1_U3256) );
  XNOR2_X1 U13185 ( .A(n12052), .B(n13282), .ZN(n10774) );
  NAND2_X1 U13186 ( .A1(n10574), .A2(n13368), .ZN(n10772) );
  XNOR2_X1 U13187 ( .A(n10774), .B(n10772), .ZN(n10770) );
  INV_X1 U13188 ( .A(n10577), .ZN(n10580) );
  INV_X1 U13189 ( .A(n10578), .ZN(n10579) );
  NAND2_X1 U13190 ( .A1(n10580), .A2(n10579), .ZN(n10581) );
  XOR2_X1 U13191 ( .A(n10771), .B(n10770), .Z(n10587) );
  NAND2_X1 U13192 ( .A1(n13496), .A2(n13367), .ZN(n10583) );
  NAND2_X1 U13193 ( .A1(n13462), .A2(n13369), .ZN(n10582) );
  NAND2_X1 U13194 ( .A1(n10583), .A2(n10582), .ZN(n10980) );
  NOR2_X1 U13195 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9243), .ZN(n13377) );
  AOI21_X1 U13196 ( .B1(n13342), .B2(n10980), .A(n13377), .ZN(n10585) );
  NAND2_X1 U13197 ( .A1(n13346), .A2(n12052), .ZN(n10584) );
  OAI211_X1 U13198 ( .C1(n13344), .C2(n10985), .A(n10585), .B(n10584), .ZN(
        n10586) );
  AOI21_X1 U13199 ( .B1(n10587), .B2(n13326), .A(n10586), .ZN(n10588) );
  INV_X1 U13200 ( .A(n10588), .ZN(P2_U3185) );
  NAND3_X1 U13201 ( .A1(n10538), .A2(n10590), .A3(n10589), .ZN(n10591) );
  AOI21_X1 U13202 ( .B1(n10592), .B2(n10591), .A(n14761), .ZN(n10600) );
  NAND3_X1 U13203 ( .A1(n10541), .A2(n10594), .A3(n10593), .ZN(n10595) );
  AOI21_X1 U13204 ( .B1(n10596), .B2(n10595), .A(n14755), .ZN(n10599) );
  OAI22_X1 U13205 ( .A1(n10597), .A2(n14276), .B1(n14770), .B2(n11240), .ZN(
        n10598) );
  OR3_X1 U13206 ( .A1(n10600), .A2(n10599), .A3(n10598), .ZN(n10974) );
  OAI21_X1 U13207 ( .B1(n10601), .B2(n10973), .A(n14365), .ZN(n10602) );
  NOR2_X1 U13208 ( .A1(n10602), .A2(n10815), .ZN(n10977) );
  NOR2_X1 U13209 ( .A1(n10974), .A2(n10977), .ZN(n10607) );
  INV_X1 U13210 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n10603) );
  OAI22_X1 U13211 ( .A1(n10973), .A2(n14411), .B1(n14806), .B2(n10603), .ZN(
        n10604) );
  INV_X1 U13212 ( .A(n10604), .ZN(n10605) );
  OAI21_X1 U13213 ( .B1(n10607), .B2(n14804), .A(n10605), .ZN(P1_U3480) );
  AOI22_X1 U13214 ( .A1(n14341), .A2(n10969), .B1(n14809), .B2(
        P1_REG1_REG_7__SCAN_IN), .ZN(n10606) );
  OAI21_X1 U13215 ( .B1(n10607), .B2(n14809), .A(n10606), .ZN(P1_U3535) );
  INV_X1 U13216 ( .A(n10608), .ZN(n10621) );
  AND2_X1 U13217 ( .A1(n13624), .A2(n10609), .ZN(n10610) );
  INV_X1 U13218 ( .A(n10611), .ZN(n10612) );
  MUX2_X1 U13219 ( .A(n10613), .B(n10612), .S(n13602), .Z(n10620) );
  INV_X1 U13220 ( .A(n10614), .ZN(n10615) );
  OAI22_X1 U13221 ( .A1(n13610), .A2(n12029), .B1(n13535), .B2(n10616), .ZN(
        n10617) );
  AOI21_X1 U13222 ( .B1(n10618), .B2(n13613), .A(n10617), .ZN(n10619) );
  OAI211_X1 U13223 ( .C1(n10621), .C2(n14942), .A(n10620), .B(n10619), .ZN(
        P2_U3261) );
  NAND2_X1 U13224 ( .A1(n10623), .A2(n10622), .ZN(n10624) );
  AND2_X1 U13225 ( .A1(n10631), .A2(n11975), .ZN(n10627) );
  AOI21_X1 U13226 ( .B1(n11979), .B2(n13938), .A(n10627), .ZN(n10692) );
  NAND2_X1 U13227 ( .A1(n10631), .A2(n11980), .ZN(n10629) );
  NAND2_X1 U13228 ( .A1(n13938), .A2(n11975), .ZN(n10628) );
  NAND2_X1 U13229 ( .A1(n10629), .A2(n10628), .ZN(n10630) );
  XNOR2_X1 U13230 ( .A(n10630), .B(n11149), .ZN(n10689) );
  XOR2_X1 U13231 ( .A(n10690), .B(n10689), .Z(n10635) );
  NOR2_X1 U13232 ( .A1(n14684), .A2(n10641), .ZN(n10634) );
  INV_X1 U13233 ( .A(n13818), .ZN(n13870) );
  NAND2_X1 U13234 ( .A1(n14679), .A2(n10631), .ZN(n10632) );
  NAND2_X1 U13235 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3086), .ZN(n13969) );
  OAI211_X1 U13236 ( .C1(n13870), .C2(n10637), .A(n10632), .B(n13969), .ZN(
        n10633) );
  AOI211_X1 U13237 ( .C1(n10635), .C2(n13880), .A(n10634), .B(n10633), .ZN(
        n10636) );
  INV_X1 U13238 ( .A(n10636), .ZN(P1_U3230) );
  INV_X1 U13239 ( .A(n14235), .ZN(n14286) );
  AND2_X1 U13240 ( .A1(n10638), .A2(n10637), .ZN(n10639) );
  MUX2_X1 U13241 ( .A(n10640), .B(n10639), .S(n14256), .Z(n10646) );
  OAI22_X1 U13242 ( .A1(n14271), .A2(n10642), .B1(n14777), .B2(n10641), .ZN(
        n10643) );
  AOI21_X1 U13243 ( .B1(n10644), .B2(n14284), .A(n10643), .ZN(n10645) );
  OAI211_X1 U13244 ( .C1(n10647), .C2(n14286), .A(n10646), .B(n10645), .ZN(
        P1_U3289) );
  INV_X1 U13245 ( .A(n10648), .ZN(n10649) );
  AOI21_X1 U13246 ( .B1(n10651), .B2(n10650), .A(n10649), .ZN(n10657) );
  INV_X1 U13247 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n10652) );
  NOR2_X1 U13248 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10652), .ZN(n15059) );
  AOI21_X1 U13249 ( .B1(n12709), .B2(n15120), .A(n15059), .ZN(n10654) );
  NAND2_X1 U13250 ( .A1(n12728), .A2(n12743), .ZN(n10653) );
  OAI211_X1 U13251 ( .C1(n12731), .C2(n15168), .A(n10654), .B(n10653), .ZN(
        n10655) );
  AOI21_X1 U13252 ( .B1(n10734), .B2(n12724), .A(n10655), .ZN(n10656) );
  OAI21_X1 U13253 ( .B1(n10657), .B2(n12704), .A(n10656), .ZN(P3_U3170) );
  XNOR2_X1 U13254 ( .A(n6721), .B(n13370), .ZN(n12252) );
  XNOR2_X1 U13255 ( .A(n10658), .B(n12252), .ZN(n14967) );
  XOR2_X1 U13256 ( .A(n12252), .B(n10659), .Z(n10661) );
  OAI21_X1 U13257 ( .B1(n10661), .B2(n13600), .A(n10660), .ZN(n14962) );
  INV_X1 U13258 ( .A(n14962), .ZN(n10662) );
  MUX2_X1 U13259 ( .A(n10663), .B(n10662), .S(n13602), .Z(n10670) );
  AOI211_X1 U13260 ( .C1(n6721), .C2(n10664), .A(n10574), .B(n10851), .ZN(
        n14963) );
  INV_X1 U13261 ( .A(n10665), .ZN(n10666) );
  OAI22_X1 U13262 ( .A1(n13610), .A2(n10667), .B1(n13535), .B2(n10666), .ZN(
        n10668) );
  AOI21_X1 U13263 ( .B1(n14963), .B2(n13613), .A(n10668), .ZN(n10669) );
  OAI211_X1 U13264 ( .C1(n14942), .C2(n14967), .A(n10670), .B(n10669), .ZN(
        P2_U3260) );
  XNOR2_X1 U13265 ( .A(n11319), .B(n11773), .ZN(n10674) );
  AOI21_X1 U13266 ( .B1(n10672), .B2(P1_REG1_REG_13__SCAN_IN), .A(n10671), 
        .ZN(n10673) );
  NAND2_X1 U13267 ( .A1(n10673), .A2(n10674), .ZN(n11318) );
  OAI21_X1 U13268 ( .B1(n10674), .B2(n10673), .A(n11318), .ZN(n10687) );
  INV_X1 U13269 ( .A(n14040), .ZN(n14749) );
  INV_X1 U13270 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n11326) );
  MUX2_X1 U13271 ( .A(n11326), .B(P1_REG2_REG_14__SCAN_IN), .S(n11319), .Z(
        n10678) );
  NOR2_X1 U13272 ( .A1(n10676), .A2(n10675), .ZN(n10680) );
  INV_X1 U13273 ( .A(n10680), .ZN(n10677) );
  NAND2_X1 U13274 ( .A1(n10678), .A2(n10677), .ZN(n10681) );
  MUX2_X1 U13275 ( .A(P1_REG2_REG_14__SCAN_IN), .B(n11326), .S(n11319), .Z(
        n10679) );
  OAI21_X1 U13276 ( .B1(n10682), .B2(n10680), .A(n10679), .ZN(n11324) );
  OAI211_X1 U13277 ( .C1(n10682), .C2(n10681), .A(n11324), .B(n14059), .ZN(
        n10685) );
  NAND2_X1 U13278 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n14681)
         );
  INV_X1 U13279 ( .A(n14681), .ZN(n10683) );
  AOI21_X1 U13280 ( .B1(n14719), .B2(P1_ADDR_REG_14__SCAN_IN), .A(n10683), 
        .ZN(n10684) );
  OAI211_X1 U13281 ( .C1(n14744), .C2(n11325), .A(n10685), .B(n10684), .ZN(
        n10686) );
  AOI21_X1 U13282 ( .B1(n10687), .B2(n14749), .A(n10686), .ZN(n10688) );
  INV_X1 U13283 ( .A(n10688), .ZN(P1_U3257) );
  NAND2_X1 U13284 ( .A1(n10690), .A2(n10689), .ZN(n10695) );
  INV_X1 U13285 ( .A(n10692), .ZN(n10693) );
  NAND2_X1 U13286 ( .A1(n10691), .A2(n10693), .ZN(n10694) );
  NAND2_X1 U13287 ( .A1(n10695), .A2(n10694), .ZN(n10754) );
  NAND2_X1 U13288 ( .A1(n10744), .A2(n11980), .ZN(n10697) );
  NAND2_X1 U13289 ( .A1(n13937), .A2(n11975), .ZN(n10696) );
  NAND2_X1 U13290 ( .A1(n10697), .A2(n10696), .ZN(n10698) );
  XNOR2_X1 U13291 ( .A(n10698), .B(n8150), .ZN(n10699) );
  AOI22_X1 U13292 ( .A1(n11979), .A2(n13937), .B1(n11975), .B2(n10744), .ZN(
        n10700) );
  NAND2_X1 U13293 ( .A1(n10699), .A2(n10700), .ZN(n10753) );
  INV_X1 U13294 ( .A(n10699), .ZN(n10702) );
  INV_X1 U13295 ( .A(n10700), .ZN(n10701) );
  NAND2_X1 U13296 ( .A1(n10702), .A2(n10701), .ZN(n10755) );
  NAND2_X1 U13297 ( .A1(n10753), .A2(n10755), .ZN(n10703) );
  XNOR2_X1 U13298 ( .A(n10754), .B(n10703), .ZN(n10710) );
  AOI22_X1 U13299 ( .A1(n13900), .A2(n13938), .B1(P1_REG3_REG_5__SCAN_IN), 
        .B2(P1_U3086), .ZN(n10708) );
  INV_X1 U13300 ( .A(n10704), .ZN(n10740) );
  OR2_X1 U13301 ( .A1(n14684), .A2(n10740), .ZN(n10707) );
  NAND2_X1 U13302 ( .A1(n14679), .A2(n10744), .ZN(n10706) );
  NAND2_X1 U13303 ( .A1(n14665), .A2(n13936), .ZN(n10705) );
  NAND4_X1 U13304 ( .A1(n10708), .A2(n10707), .A3(n10706), .A4(n10705), .ZN(
        n10709) );
  AOI21_X1 U13305 ( .B1(n10710), .B2(n13880), .A(n10709), .ZN(n10711) );
  INV_X1 U13306 ( .A(n10711), .ZN(P1_U3227) );
  INV_X1 U13307 ( .A(P3_DATAO_REG_26__SCAN_IN), .ZN(n15363) );
  NAND2_X1 U13308 ( .A1(n12657), .A2(P3_U3897), .ZN(n10712) );
  OAI21_X1 U13309 ( .B1(P3_U3897), .B2(n15363), .A(n10712), .ZN(P3_U3517) );
  NAND2_X1 U13310 ( .A1(n10713), .A2(n12257), .ZN(n10714) );
  NAND2_X1 U13311 ( .A1(n10715), .A2(n10714), .ZN(n14985) );
  XNOR2_X1 U13312 ( .A(n10716), .B(n12257), .ZN(n10717) );
  NAND2_X1 U13313 ( .A1(n10717), .A2(n13618), .ZN(n10719) );
  AOI22_X1 U13314 ( .A1(n13462), .A2(n13368), .B1(n13496), .B2(n13366), .ZN(
        n10718) );
  OAI211_X1 U13315 ( .C1(n14985), .C2(n13624), .A(n10719), .B(n10718), .ZN(
        n14987) );
  NAND2_X1 U13316 ( .A1(n14987), .A2(n13602), .ZN(n10725) );
  OAI22_X1 U13317 ( .A1(n13602), .A2(n10720), .B1(n10786), .B2(n13535), .ZN(
        n10723) );
  INV_X1 U13318 ( .A(n10983), .ZN(n10721) );
  OAI211_X1 U13319 ( .C1(n7191), .C2(n10721), .A(n13603), .B(n10923), .ZN(
        n14986) );
  NOR2_X1 U13320 ( .A1(n14986), .A2(n14939), .ZN(n10722) );
  AOI211_X1 U13321 ( .C1(n14935), .C2(n12060), .A(n10723), .B(n10722), .ZN(
        n10724) );
  OAI211_X1 U13322 ( .C1(n14985), .C2(n11317), .A(n10725), .B(n10724), .ZN(
        P2_U3257) );
  NAND2_X1 U13323 ( .A1(n12745), .A2(P3_DATAO_REG_30__SCAN_IN), .ZN(n10726) );
  OAI21_X1 U13324 ( .B1(n12373), .B2(n12745), .A(n10726), .ZN(P3_U3521) );
  XNOR2_X1 U13325 ( .A(n10728), .B(n10727), .ZN(n10732) );
  INV_X1 U13326 ( .A(n13067), .ZN(n15139) );
  INV_X1 U13327 ( .A(n13069), .ZN(n15136) );
  AOI22_X1 U13328 ( .A1(n15139), .A2(n15120), .B1(n12743), .B2(n15136), .ZN(
        n10731) );
  XNOR2_X1 U13329 ( .A(n10729), .B(n12433), .ZN(n15167) );
  INV_X1 U13330 ( .A(n15147), .ZN(n12945) );
  NAND2_X1 U13331 ( .A1(n15167), .A2(n12945), .ZN(n10730) );
  OAI211_X1 U13332 ( .C1(n10732), .C2(n13064), .A(n10731), .B(n10730), .ZN(
        n15171) );
  INV_X1 U13333 ( .A(n15171), .ZN(n10739) );
  INV_X2 U13334 ( .A(n15132), .ZN(n13074) );
  NAND2_X1 U13335 ( .A1(n10733), .A2(n15134), .ZN(n11447) );
  INV_X1 U13336 ( .A(n11447), .ZN(n15131) );
  AOI22_X1 U13337 ( .A1(n14617), .A2(n10735), .B1(n15150), .B2(n10734), .ZN(
        n10736) );
  OAI21_X1 U13338 ( .B1(n10860), .B2(n15132), .A(n10736), .ZN(n10737) );
  AOI21_X1 U13339 ( .B1(n15167), .B2(n15151), .A(n10737), .ZN(n10738) );
  OAI21_X1 U13340 ( .B1(n10739), .B2(n13074), .A(n10738), .ZN(P3_U3229) );
  OAI22_X1 U13341 ( .A1(n14256), .A2(n7763), .B1(n10740), .B2(n14777), .ZN(
        n10743) );
  NOR2_X1 U13342 ( .A1(n14261), .A2(n10741), .ZN(n10742) );
  AOI211_X1 U13343 ( .C1(n14258), .C2(n10744), .A(n10743), .B(n10742), .ZN(
        n10745) );
  OAI21_X1 U13344 ( .B1(n10746), .B2(n14281), .A(n10745), .ZN(P1_U3288) );
  MUX2_X1 U13345 ( .A(n10748), .B(n10747), .S(n14256), .Z(n10751) );
  INV_X1 U13346 ( .A(n10762), .ZN(n10749) );
  AOI22_X1 U13347 ( .A1(n14258), .A2(n10767), .B1(n10749), .B2(n14786), .ZN(
        n10750) );
  OAI211_X1 U13348 ( .C1(n14261), .C2(n10752), .A(n10751), .B(n10750), .ZN(
        P1_U3287) );
  NAND2_X1 U13349 ( .A1(n10754), .A2(n10753), .ZN(n10756) );
  NAND2_X1 U13350 ( .A1(n10756), .A2(n10755), .ZN(n10761) );
  NAND2_X1 U13351 ( .A1(n10767), .A2(n11980), .ZN(n10758) );
  NAND2_X1 U13352 ( .A1(n13936), .A2(n11975), .ZN(n10757) );
  NAND2_X1 U13353 ( .A1(n10758), .A2(n10757), .ZN(n10759) );
  XNOR2_X1 U13354 ( .A(n10759), .B(n11149), .ZN(n10953) );
  AOI22_X1 U13355 ( .A1(n10767), .A2(n11975), .B1(n11979), .B2(n13936), .ZN(
        n10954) );
  XNOR2_X1 U13356 ( .A(n10953), .B(n10954), .ZN(n10760) );
  NAND2_X1 U13357 ( .A1(n10761), .A2(n10760), .ZN(n10957) );
  OAI211_X1 U13358 ( .C1(n10761), .C2(n10760), .A(n10957), .B(n13880), .ZN(
        n10769) );
  NOR2_X1 U13359 ( .A1(n14684), .A2(n10762), .ZN(n10766) );
  NAND2_X1 U13360 ( .A1(n14665), .A2(n13935), .ZN(n10764) );
  NAND2_X1 U13361 ( .A1(n13900), .A2(n13937), .ZN(n10763) );
  NAND2_X1 U13362 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n13986) );
  NAND3_X1 U13363 ( .A1(n10764), .A2(n10763), .A3(n13986), .ZN(n10765) );
  AOI211_X1 U13364 ( .C1(n10767), .C2(n14679), .A(n10766), .B(n10765), .ZN(
        n10768) );
  NAND2_X1 U13365 ( .A1(n10769), .A2(n10768), .ZN(P1_U3239) );
  NAND2_X1 U13366 ( .A1(n10771), .A2(n10770), .ZN(n10776) );
  INV_X1 U13367 ( .A(n10772), .ZN(n10773) );
  NAND2_X1 U13368 ( .A1(n10774), .A2(n10773), .ZN(n10775) );
  NAND2_X1 U13369 ( .A1(n10574), .A2(n13367), .ZN(n10778) );
  INV_X1 U13370 ( .A(n10777), .ZN(n10780) );
  INV_X1 U13371 ( .A(n10778), .ZN(n10779) );
  NAND2_X1 U13372 ( .A1(n10780), .A2(n10779), .ZN(n10781) );
  NAND2_X1 U13373 ( .A1(n10935), .A2(n10781), .ZN(n10783) );
  INV_X1 U13374 ( .A(n10936), .ZN(n10782) );
  AOI21_X1 U13375 ( .B1(n10784), .B2(n10783), .A(n10782), .ZN(n10791) );
  NAND2_X1 U13376 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3088), .ZN(n14853) );
  OAI21_X1 U13377 ( .B1(n13328), .B2(n10785), .A(n14853), .ZN(n10789) );
  OAI22_X1 U13378 ( .A1(n13329), .A2(n10787), .B1(n13344), .B2(n10786), .ZN(
        n10788) );
  AOI211_X1 U13379 ( .C1(n12060), .C2(n13346), .A(n10789), .B(n10788), .ZN(
        n10790) );
  OAI21_X1 U13380 ( .B1(n10791), .B2(n13348), .A(n10790), .ZN(P2_U3193) );
  INV_X1 U13381 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n15294) );
  INV_X1 U13382 ( .A(P3_REG2_REG_31__SCAN_IN), .ZN(n14612) );
  NAND2_X1 U13383 ( .A1(n10792), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n10795) );
  NAND2_X1 U13384 ( .A1(n10793), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n10794) );
  OAI211_X1 U13385 ( .C1(n14612), .C2(n10796), .A(n10795), .B(n10794), .ZN(
        n10797) );
  INV_X1 U13386 ( .A(n10797), .ZN(n10798) );
  NAND2_X1 U13387 ( .A1(n10799), .A2(n10798), .ZN(n12376) );
  NAND2_X1 U13388 ( .A1(n12376), .A2(P3_U3897), .ZN(n10800) );
  OAI21_X1 U13389 ( .B1(P3_U3897), .B2(n15294), .A(n10800), .ZN(P3_U3522) );
  INV_X1 U13390 ( .A(n10801), .ZN(n10803) );
  OAI222_X1 U13391 ( .A1(P3_U3151), .A2(n10804), .B1(n13213), .B2(n10803), 
        .C1(n10802), .C2(n13217), .ZN(P3_U3275) );
  INV_X1 U13392 ( .A(n10805), .ZN(n10806) );
  AOI211_X1 U13393 ( .C1(n10812), .C2(n10807), .A(n14761), .B(n10806), .ZN(
        n10810) );
  NAND2_X1 U13394 ( .A1(n14757), .A2(n13935), .ZN(n10809) );
  NAND2_X1 U13395 ( .A1(n14247), .A2(n13933), .ZN(n10808) );
  NAND2_X1 U13396 ( .A1(n10809), .A2(n10808), .ZN(n11160) );
  OR2_X1 U13397 ( .A1(n10810), .A2(n11160), .ZN(n10826) );
  OAI21_X1 U13398 ( .B1(n10813), .B2(n10812), .A(n10811), .ZN(n10814) );
  INV_X1 U13399 ( .A(n10814), .ZN(n10829) );
  XNOR2_X1 U13400 ( .A(n10815), .B(n10818), .ZN(n10824) );
  OAI22_X1 U13401 ( .A1(n10829), .A2(n14755), .B1(n14793), .B2(n10824), .ZN(
        n10816) );
  NOR2_X1 U13402 ( .A1(n10826), .A2(n10816), .ZN(n10822) );
  INV_X1 U13403 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n10817) );
  OAI22_X1 U13404 ( .A1(n10818), .A2(n14411), .B1(n14806), .B2(n10817), .ZN(
        n10819) );
  INV_X1 U13405 ( .A(n10819), .ZN(n10820) );
  OAI21_X1 U13406 ( .B1(n10822), .B2(n14804), .A(n10820), .ZN(P1_U3483) );
  AOI22_X1 U13407 ( .A1(n11164), .A2(n14341), .B1(n14809), .B2(
        P1_REG1_REG_8__SCAN_IN), .ZN(n10821) );
  OAI21_X1 U13408 ( .B1(n10822), .B2(n14809), .A(n10821), .ZN(P1_U3536) );
  OAI22_X1 U13409 ( .A1(n10824), .A2(n10823), .B1(n11162), .B2(n14777), .ZN(
        n10825) );
  OAI21_X1 U13410 ( .B1(n10826), .B2(n10825), .A(n14256), .ZN(n10828) );
  AOI22_X1 U13411 ( .A1(n14258), .A2(n11164), .B1(n14281), .B2(
        P1_REG2_REG_8__SCAN_IN), .ZN(n10827) );
  OAI211_X1 U13412 ( .C1(n10829), .C2(n14286), .A(n10828), .B(n10827), .ZN(
        P1_U3285) );
  INV_X1 U13413 ( .A(n10830), .ZN(n10832) );
  INV_X1 U13414 ( .A(n14052), .ZN(n14046) );
  OAI222_X1 U13415 ( .A1(n14433), .A2(n10831), .B1(n12610), .B2(n10832), .C1(
        P1_U3086), .C2(n14046), .ZN(P1_U3337) );
  OAI222_X1 U13416 ( .A1(n13768), .A2(n10833), .B1(n6551), .B2(n10832), .C1(
        P2_U3088), .C2(n14920), .ZN(P2_U3309) );
  OAI21_X1 U13417 ( .B1(n10835), .B2(n10834), .A(n11107), .ZN(n10842) );
  NAND2_X1 U13418 ( .A1(n12724), .A2(n11078), .ZN(n10840) );
  NOR2_X1 U13419 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10836), .ZN(n15081) );
  AOI21_X1 U13420 ( .B1(n12709), .B2(n12744), .A(n15081), .ZN(n10839) );
  NAND2_X1 U13421 ( .A1(n12728), .A2(n12742), .ZN(n10838) );
  NAND2_X1 U13422 ( .A1(n12702), .A2(n11079), .ZN(n10837) );
  NAND4_X1 U13423 ( .A1(n10840), .A2(n10839), .A3(n10838), .A4(n10837), .ZN(
        n10841) );
  AOI21_X1 U13424 ( .B1(n10842), .B2(n12722), .A(n10841), .ZN(n10843) );
  INV_X1 U13425 ( .A(n10843), .ZN(P3_U3167) );
  INV_X1 U13426 ( .A(n10844), .ZN(n10846) );
  OAI21_X1 U13427 ( .B1(n10846), .B2(n12254), .A(n10845), .ZN(n10848) );
  AOI21_X1 U13428 ( .B1(n10848), .B2(n13618), .A(n10847), .ZN(n14973) );
  INV_X2 U13429 ( .A(n14947), .ZN(n13602) );
  OAI22_X1 U13430 ( .A1(n13602), .A2(n10850), .B1(n10849), .B2(n13535), .ZN(
        n10854) );
  OAI21_X1 U13431 ( .B1(n10851), .B2(n14974), .A(n13603), .ZN(n10852) );
  OR2_X1 U13432 ( .A1(n10852), .A2(n10984), .ZN(n14972) );
  NOR2_X1 U13433 ( .A1(n14972), .A2(n14939), .ZN(n10853) );
  AOI211_X1 U13434 ( .C1(n14935), .C2(n12048), .A(n10854), .B(n10853), .ZN(
        n10857) );
  XNOR2_X1 U13435 ( .A(n10855), .B(n12254), .ZN(n14971) );
  INV_X1 U13436 ( .A(n14971), .ZN(n14977) );
  INV_X1 U13437 ( .A(n14942), .ZN(n13579) );
  NAND2_X1 U13438 ( .A1(n14977), .A2(n13579), .ZN(n10856) );
  OAI211_X1 U13439 ( .C1(n14973), .C2(n14947), .A(n10857), .B(n10856), .ZN(
        P2_U3259) );
  MUX2_X1 U13440 ( .A(P3_REG2_REG_4__SCAN_IN), .B(n10860), .S(n10895), .Z(
        n15054) );
  NOR2_X1 U13441 ( .A1(n15055), .A2(n15054), .ZN(n15053) );
  OAI21_X1 U13442 ( .B1(n10861), .B2(n10896), .A(n15073), .ZN(n12346) );
  MUX2_X1 U13443 ( .A(n8622), .B(P3_REG2_REG_6__SCAN_IN), .S(n10899), .Z(
        n12347) );
  NOR2_X1 U13444 ( .A1(n10900), .A2(n10862), .ZN(n10864) );
  AOI22_X1 U13445 ( .A1(P3_REG2_REG_8__SCAN_IN), .A2(n10903), .B1(n12324), 
        .B2(n8660), .ZN(n12315) );
  NOR2_X1 U13446 ( .A1(n12316), .A2(n12315), .ZN(n10865) );
  AOI21_X1 U13447 ( .B1(P3_REG2_REG_8__SCAN_IN), .B2(n12324), .A(n10865), .ZN(
        n10866) );
  XNOR2_X1 U13448 ( .A(n10883), .B(n10866), .ZN(n15093) );
  INV_X1 U13449 ( .A(n11246), .ZN(n11249) );
  AOI22_X1 U13450 ( .A1(P3_REG2_REG_10__SCAN_IN), .A2(n11249), .B1(n11246), 
        .B2(n11454), .ZN(n10867) );
  AOI21_X1 U13451 ( .B1(n6670), .B2(n10867), .A(n11245), .ZN(n10913) );
  MUX2_X1 U13452 ( .A(P3_REG2_REG_4__SCAN_IN), .B(P3_REG1_REG_4__SCAN_IN), .S(
        n13209), .Z(n10876) );
  INV_X1 U13453 ( .A(n15038), .ZN(n10874) );
  INV_X1 U13454 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n10868) );
  MUX2_X1 U13455 ( .A(n10869), .B(n10868), .S(n13209), .Z(n10870) );
  NAND2_X1 U13456 ( .A1(n10870), .A2(n10893), .ZN(n10875) );
  INV_X1 U13457 ( .A(n10870), .ZN(n10871) );
  NAND2_X1 U13458 ( .A1(n10871), .A2(n15045), .ZN(n10872) );
  NAND2_X1 U13459 ( .A1(n10875), .A2(n10872), .ZN(n15039) );
  INV_X1 U13460 ( .A(n15039), .ZN(n10873) );
  OAI21_X1 U13461 ( .B1(n15042), .B2(n10874), .A(n10873), .ZN(n15040) );
  NAND2_X1 U13462 ( .A1(n15040), .A2(n10875), .ZN(n15058) );
  XNOR2_X1 U13463 ( .A(n10876), .B(n10895), .ZN(n15057) );
  NAND2_X1 U13464 ( .A1(n15058), .A2(n15057), .ZN(n15056) );
  OAI21_X1 U13465 ( .B1(n10876), .B2(n15061), .A(n15056), .ZN(n15080) );
  MUX2_X1 U13466 ( .A(P3_REG2_REG_5__SCAN_IN), .B(P3_REG1_REG_5__SCAN_IN), .S(
        n13209), .Z(n10877) );
  NAND2_X1 U13467 ( .A1(n10877), .A2(n15083), .ZN(n15076) );
  NOR2_X1 U13468 ( .A1(n10877), .A2(n15083), .ZN(n15078) );
  AOI21_X1 U13469 ( .B1(n15080), .B2(n15076), .A(n15078), .ZN(n12343) );
  MUX2_X1 U13470 ( .A(P3_REG2_REG_6__SCAN_IN), .B(P3_REG1_REG_6__SCAN_IN), .S(
        n13209), .Z(n10878) );
  XOR2_X1 U13471 ( .A(n10899), .B(n10878), .Z(n12344) );
  MUX2_X1 U13472 ( .A(P3_REG2_REG_7__SCAN_IN), .B(P3_REG1_REG_7__SCAN_IN), .S(
        n13209), .Z(n10879) );
  XNOR2_X1 U13473 ( .A(n10879), .B(n10900), .ZN(n12330) );
  INV_X1 U13474 ( .A(n10879), .ZN(n10880) );
  MUX2_X1 U13475 ( .A(P3_REG2_REG_8__SCAN_IN), .B(P3_REG1_REG_8__SCAN_IN), .S(
        n13209), .Z(n10881) );
  XNOR2_X1 U13476 ( .A(n10881), .B(n12324), .ZN(n12314) );
  MUX2_X1 U13477 ( .A(P3_REG2_REG_9__SCAN_IN), .B(P3_REG1_REG_9__SCAN_IN), .S(
        n13209), .Z(n10882) );
  NAND2_X1 U13478 ( .A1(n10882), .A2(n15101), .ZN(n15096) );
  INV_X1 U13479 ( .A(n10882), .ZN(n10884) );
  NAND2_X1 U13480 ( .A1(n10884), .A2(n10883), .ZN(n15098) );
  INV_X1 U13481 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n10885) );
  MUX2_X1 U13482 ( .A(n11454), .B(n10885), .S(n13209), .Z(n10886) );
  NAND2_X1 U13483 ( .A1(n10886), .A2(n11249), .ZN(n11252) );
  INV_X1 U13484 ( .A(n10886), .ZN(n10887) );
  NAND2_X1 U13485 ( .A1(n10887), .A2(n11246), .ZN(n10888) );
  NAND2_X1 U13486 ( .A1(n11252), .A2(n10888), .ZN(n10889) );
  AOI21_X1 U13487 ( .B1(n15094), .B2(n15098), .A(n10889), .ZN(n11254) );
  AND3_X1 U13488 ( .A1(n15094), .A2(n15098), .A3(n10889), .ZN(n10890) );
  OAI21_X1 U13489 ( .B1(n11254), .B2(n10890), .A(n15085), .ZN(n10912) );
  AOI22_X1 U13490 ( .A1(P3_REG1_REG_10__SCAN_IN), .A2(n11246), .B1(n11249), 
        .B2(n10885), .ZN(n10907) );
  INV_X1 U13491 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n15217) );
  AOI22_X1 U13492 ( .A1(P3_REG1_REG_8__SCAN_IN), .A2(n12324), .B1(n10903), 
        .B2(n15217), .ZN(n12319) );
  INV_X1 U13493 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n15213) );
  INV_X1 U13494 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n15210) );
  OAI21_X1 U13495 ( .B1(n10892), .B2(n10225), .A(n10891), .ZN(n10894) );
  XNOR2_X1 U13496 ( .A(n10894), .B(n10893), .ZN(n15048) );
  AOI22_X1 U13497 ( .A1(n15048), .A2(P3_REG1_REG_3__SCAN_IN), .B1(n15045), 
        .B2(n10894), .ZN(n15067) );
  MUX2_X1 U13498 ( .A(P3_REG1_REG_4__SCAN_IN), .B(n15210), .S(n10895), .Z(
        n15066) );
  OAI21_X1 U13499 ( .B1(n10895), .B2(n15210), .A(n15064), .ZN(n10897) );
  MUX2_X1 U13500 ( .A(P3_REG1_REG_6__SCAN_IN), .B(n15213), .S(n10899), .Z(
        n12350) );
  OAI21_X1 U13501 ( .B1(n10899), .B2(n15213), .A(n10898), .ZN(n10901) );
  NAND2_X1 U13502 ( .A1(n12338), .A2(n10901), .ZN(n10902) );
  XNOR2_X1 U13503 ( .A(n10901), .B(n10900), .ZN(n12333) );
  NAND2_X1 U13504 ( .A1(P3_REG1_REG_7__SCAN_IN), .A2(n12333), .ZN(n12332) );
  NAND2_X1 U13505 ( .A1(n15101), .A2(n10904), .ZN(n10905) );
  NAND2_X1 U13506 ( .A1(P3_REG1_REG_9__SCAN_IN), .A2(n15108), .ZN(n15107) );
  OAI21_X1 U13507 ( .B1(n10907), .B2(n10906), .A(n11248), .ZN(n10910) );
  INV_X1 U13508 ( .A(P3_REG3_REG_10__SCAN_IN), .ZN(n15462) );
  NOR2_X1 U13509 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15462), .ZN(n11123) );
  AOI21_X1 U13510 ( .B1(n15106), .B2(P3_ADDR_REG_10__SCAN_IN), .A(n11123), 
        .ZN(n10908) );
  OAI21_X1 U13511 ( .B1(n15100), .B2(n11246), .A(n10908), .ZN(n10909) );
  AOI21_X1 U13512 ( .B1(n10910), .B2(n15109), .A(n10909), .ZN(n10911) );
  OAI211_X1 U13513 ( .C1(n10913), .C2(n15113), .A(n10912), .B(n10911), .ZN(
        P3_U3192) );
  OR2_X1 U13514 ( .A1(n10914), .A2(n10917), .ZN(n10915) );
  NAND2_X1 U13515 ( .A1(n10916), .A2(n10915), .ZN(n14991) );
  XNOR2_X1 U13516 ( .A(n10918), .B(n10917), .ZN(n10919) );
  NAND2_X1 U13517 ( .A1(n10919), .A2(n13618), .ZN(n10921) );
  AOI22_X1 U13518 ( .A1(n13462), .A2(n13367), .B1(n13496), .B2(n13365), .ZN(
        n10920) );
  OAI211_X1 U13519 ( .C1(n13624), .C2(n14991), .A(n10921), .B(n10920), .ZN(
        n14993) );
  NAND2_X1 U13520 ( .A1(n14993), .A2(n13602), .ZN(n10929) );
  OAI22_X1 U13521 ( .A1(n13602), .A2(n10922), .B1(n10940), .B2(n13535), .ZN(
        n10927) );
  INV_X1 U13522 ( .A(n10923), .ZN(n10925) );
  INV_X1 U13523 ( .A(n11011), .ZN(n10924) );
  OAI211_X1 U13524 ( .C1(n6979), .C2(n10925), .A(n10924), .B(n13603), .ZN(
        n14992) );
  NOR2_X1 U13525 ( .A1(n14992), .A2(n14939), .ZN(n10926) );
  AOI211_X1 U13526 ( .C1(n14935), .C2(n6703), .A(n10927), .B(n10926), .ZN(
        n10928) );
  OAI211_X1 U13527 ( .C1(n14991), .C2(n11317), .A(n10929), .B(n10928), .ZN(
        P2_U3256) );
  NAND2_X1 U13528 ( .A1(n10574), .A2(n13366), .ZN(n10931) );
  INV_X1 U13529 ( .A(n10930), .ZN(n10933) );
  INV_X1 U13530 ( .A(n10931), .ZN(n10932) );
  NAND2_X1 U13531 ( .A1(n10933), .A2(n10932), .ZN(n10934) );
  AND2_X1 U13532 ( .A1(n10993), .A2(n10934), .ZN(n10938) );
  OAI21_X1 U13533 ( .B1(n10938), .B2(n10937), .A(n10994), .ZN(n10939) );
  NAND2_X1 U13534 ( .A1(n10939), .A2(n13326), .ZN(n10944) );
  OAI22_X1 U13535 ( .A1(n13329), .A2(n12077), .B1(n13344), .B2(n10940), .ZN(
        n10941) );
  AOI211_X1 U13536 ( .C1(n11671), .C2(n13367), .A(n10942), .B(n10941), .ZN(
        n10943) );
  OAI211_X1 U13537 ( .C1(n6979), .C2(n13334), .A(n10944), .B(n10943), .ZN(
        P2_U3203) );
  OAI22_X1 U13538 ( .A1(n10946), .A2(n13610), .B1(n14939), .B2(n10945), .ZN(
        n10950) );
  OAI21_X1 U13539 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(n13535), .A(n10947), .ZN(
        n10948) );
  MUX2_X1 U13540 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n10948), .S(n13602), .Z(
        n10949) );
  AOI211_X1 U13541 ( .C1(n13579), .C2(n10951), .A(n10950), .B(n10949), .ZN(
        n10952) );
  INV_X1 U13542 ( .A(n10952), .ZN(P2_U3262) );
  INV_X1 U13543 ( .A(n10953), .ZN(n10955) );
  OR2_X1 U13544 ( .A1(n10955), .A2(n10954), .ZN(n10956) );
  NAND2_X1 U13545 ( .A1(n10969), .A2(n11980), .ZN(n10959) );
  NAND2_X1 U13546 ( .A1(n13935), .A2(n11975), .ZN(n10958) );
  NAND2_X1 U13547 ( .A1(n10959), .A2(n10958), .ZN(n10960) );
  XNOR2_X1 U13548 ( .A(n10960), .B(n11149), .ZN(n11154) );
  NOR2_X1 U13549 ( .A1(n11938), .A2(n10961), .ZN(n10962) );
  AOI21_X1 U13550 ( .B1(n10969), .B2(n11975), .A(n10962), .ZN(n11152) );
  XNOR2_X1 U13551 ( .A(n11154), .B(n11152), .ZN(n10963) );
  OAI211_X1 U13552 ( .C1(n10964), .C2(n10963), .A(n11156), .B(n13880), .ZN(
        n10971) );
  NOR2_X1 U13553 ( .A1(n14684), .A2(n10972), .ZN(n10968) );
  NAND2_X1 U13554 ( .A1(n14665), .A2(n13934), .ZN(n10966) );
  NAND2_X1 U13555 ( .A1(n13900), .A2(n13936), .ZN(n10965) );
  NAND2_X1 U13556 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n14000) );
  NAND3_X1 U13557 ( .A1(n10966), .A2(n10965), .A3(n14000), .ZN(n10967) );
  AOI211_X1 U13558 ( .C1(n10969), .C2(n14679), .A(n10968), .B(n10967), .ZN(
        n10970) );
  NAND2_X1 U13559 ( .A1(n10971), .A2(n10970), .ZN(P1_U3213) );
  OAI22_X1 U13560 ( .A1(n14271), .A2(n10973), .B1(n10972), .B2(n14777), .ZN(
        n10976) );
  MUX2_X1 U13561 ( .A(n10974), .B(P1_REG2_REG_7__SCAN_IN), .S(n14281), .Z(
        n10975) );
  AOI211_X1 U13562 ( .C1(n14284), .C2(n10977), .A(n10976), .B(n10975), .ZN(
        n10978) );
  INV_X1 U13563 ( .A(n10978), .ZN(P1_U3286) );
  XOR2_X1 U13564 ( .A(n12256), .B(n10979), .Z(n10981) );
  AOI21_X1 U13565 ( .B1(n10981), .B2(n13618), .A(n10980), .ZN(n14980) );
  XNOR2_X1 U13566 ( .A(n10982), .B(n12256), .ZN(n14984) );
  OAI211_X1 U13567 ( .C1(n14981), .C2(n10984), .A(n13603), .B(n10983), .ZN(
        n14979) );
  OAI22_X1 U13568 ( .A1(n13602), .A2(n10986), .B1(n10985), .B2(n13535), .ZN(
        n10987) );
  AOI21_X1 U13569 ( .B1(n14935), .B2(n12052), .A(n10987), .ZN(n10988) );
  OAI21_X1 U13570 ( .B1(n14979), .B2(n14939), .A(n10988), .ZN(n10989) );
  AOI21_X1 U13571 ( .B1(n14984), .B2(n13579), .A(n10989), .ZN(n10990) );
  OAI21_X1 U13572 ( .B1(n14980), .B2(n14947), .A(n10990), .ZN(P2_U3258) );
  INV_X1 U13573 ( .A(n10991), .ZN(n12614) );
  OAI222_X1 U13574 ( .A1(n14433), .A2(n10992), .B1(n12610), .B2(n12614), .C1(
        n14061), .C2(P1_U3086), .ZN(P1_U3336) );
  XNOR2_X1 U13575 ( .A(n12075), .B(n13236), .ZN(n11136) );
  NAND2_X1 U13576 ( .A1(n10574), .A2(n13365), .ZN(n11137) );
  XNOR2_X1 U13577 ( .A(n11136), .B(n11137), .ZN(n11141) );
  XNOR2_X1 U13578 ( .A(n11142), .B(n11141), .ZN(n11000) );
  OAI22_X1 U13579 ( .A1(n13329), .A2(n10995), .B1(n13344), .B2(n11009), .ZN(
        n10996) );
  AOI211_X1 U13580 ( .C1(n11671), .C2(n13366), .A(n10997), .B(n10996), .ZN(
        n10999) );
  NAND2_X1 U13581 ( .A1(n12075), .A2(n13346), .ZN(n10998) );
  OAI211_X1 U13582 ( .C1(n11000), .C2(n13348), .A(n10999), .B(n10998), .ZN(
        P2_U3189) );
  OR2_X1 U13583 ( .A1(n11001), .A2(n11004), .ZN(n11002) );
  NAND2_X1 U13584 ( .A1(n11003), .A2(n11002), .ZN(n14997) );
  XNOR2_X1 U13585 ( .A(n11005), .B(n11004), .ZN(n11006) );
  NAND2_X1 U13586 ( .A1(n11006), .A2(n13618), .ZN(n11008) );
  AOI22_X1 U13587 ( .A1(n13462), .A2(n13366), .B1(n13496), .B2(n13364), .ZN(
        n11007) );
  OAI211_X1 U13588 ( .C1(n14997), .C2(n13624), .A(n11008), .B(n11007), .ZN(
        n15001) );
  NAND2_X1 U13589 ( .A1(n15001), .A2(n13602), .ZN(n11015) );
  OAI22_X1 U13590 ( .A1(n13602), .A2(n11010), .B1(n11009), .B2(n13535), .ZN(
        n11013) );
  OAI211_X1 U13591 ( .C1(n15000), .C2(n11011), .A(n13603), .B(n11268), .ZN(
        n14998) );
  NOR2_X1 U13592 ( .A1(n14998), .A2(n14939), .ZN(n11012) );
  AOI211_X1 U13593 ( .C1(n14935), .C2(n12075), .A(n11013), .B(n11012), .ZN(
        n11014) );
  OAI211_X1 U13594 ( .C1(n14997), .C2(n11317), .A(n11015), .B(n11014), .ZN(
        P2_U3255) );
  INV_X1 U13595 ( .A(n11016), .ZN(n11017) );
  AOI21_X1 U13596 ( .B1(n11021), .B2(n11018), .A(n11017), .ZN(n11019) );
  OAI222_X1 U13597 ( .A1(n14770), .A2(n11550), .B1(n14276), .B2(n11240), .C1(
        n14761), .C2(n11019), .ZN(n14800) );
  INV_X1 U13598 ( .A(n14800), .ZN(n11030) );
  OAI21_X1 U13599 ( .B1(n11022), .B2(n11021), .A(n11020), .ZN(n14802) );
  INV_X1 U13600 ( .A(n11023), .ZN(n11024) );
  INV_X1 U13601 ( .A(n11232), .ZN(n14799) );
  OAI211_X1 U13602 ( .C1(n11024), .C2(n14799), .A(n14365), .B(n11189), .ZN(
        n14797) );
  OAI22_X1 U13603 ( .A1(n14256), .A2(n11025), .B1(n11238), .B2(n14777), .ZN(
        n11026) );
  AOI21_X1 U13604 ( .B1(n11232), .B2(n14258), .A(n11026), .ZN(n11027) );
  OAI21_X1 U13605 ( .B1(n14797), .B2(n14261), .A(n11027), .ZN(n11028) );
  AOI21_X1 U13606 ( .B1(n14802), .B2(n14235), .A(n11028), .ZN(n11029) );
  OAI21_X1 U13607 ( .B1(n11030), .B2(n14281), .A(n11029), .ZN(P1_U3284) );
  INV_X1 U13608 ( .A(n11031), .ZN(n11032) );
  INV_X1 U13609 ( .A(SI_21_), .ZN(n15415) );
  OAI222_X1 U13610 ( .A1(n13213), .A2(n11032), .B1(n13217), .B2(n15415), .C1(
        P3_U3151), .C2(n12419), .ZN(P3_U3274) );
  INV_X1 U13611 ( .A(n11033), .ZN(n12592) );
  OAI222_X1 U13612 ( .A1(n14433), .A2(n15251), .B1(P1_U3086), .B2(n6549), .C1(
        n12610), .C2(n12592), .ZN(P1_U3335) );
  AND2_X1 U13613 ( .A1(n11035), .A2(n13579), .ZN(n11041) );
  NAND2_X1 U13614 ( .A1(n13613), .A2(n11036), .ZN(n11038) );
  AOI22_X1 U13615 ( .A1(n14947), .A2(P2_REG2_REG_2__SCAN_IN), .B1(n14936), 
        .B2(P2_REG3_REG_2__SCAN_IN), .ZN(n11037) );
  OAI211_X1 U13616 ( .C1(n11039), .C2(n13610), .A(n11038), .B(n11037), .ZN(
        n11040) );
  AOI211_X1 U13617 ( .C1(n13602), .C2(n11042), .A(n11041), .B(n11040), .ZN(
        n11043) );
  INV_X1 U13618 ( .A(n11043), .ZN(P2_U3263) );
  INV_X1 U13619 ( .A(n11122), .ZN(n11045) );
  AOI21_X1 U13620 ( .B1(n11047), .B2(n11046), .A(n11045), .ZN(n11053) );
  INV_X1 U13621 ( .A(n11048), .ZN(n11346) );
  INV_X1 U13622 ( .A(n12724), .ZN(n12700) );
  NOR2_X1 U13623 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15461), .ZN(n15105) );
  INV_X1 U13624 ( .A(n12740), .ZN(n12461) );
  NOR2_X1 U13625 ( .A1(n12461), .A2(n12726), .ZN(n11049) );
  AOI211_X1 U13626 ( .C1(n12728), .C2(n12738), .A(n15105), .B(n11049), .ZN(
        n11050) );
  OAI21_X1 U13627 ( .B1(n11346), .B2(n12700), .A(n11050), .ZN(n11051) );
  AOI21_X1 U13628 ( .B1(n12414), .B2(n12702), .A(n11051), .ZN(n11052) );
  OAI21_X1 U13629 ( .B1(n11053), .B2(n12704), .A(n11052), .ZN(P3_U3171) );
  OR2_X1 U13630 ( .A1(n11054), .A2(n12384), .ZN(n11055) );
  NAND2_X1 U13631 ( .A1(n11056), .A2(n11055), .ZN(n11060) );
  INV_X1 U13632 ( .A(n11060), .ZN(n15179) );
  NAND2_X1 U13633 ( .A1(n12743), .A2(n15139), .ZN(n11058) );
  NAND2_X1 U13634 ( .A1(n12741), .A2(n15136), .ZN(n11057) );
  NAND2_X1 U13635 ( .A1(n11058), .A2(n11057), .ZN(n11059) );
  AOI21_X1 U13636 ( .B1(n11060), .B2(n12945), .A(n11059), .ZN(n11063) );
  OAI211_X1 U13637 ( .C1(n6671), .C2(n6994), .A(n11061), .B(n15143), .ZN(
        n11062) );
  NAND2_X1 U13638 ( .A1(n11063), .A2(n11062), .ZN(n15180) );
  MUX2_X1 U13639 ( .A(n15180), .B(P3_REG2_REG_6__SCAN_IN), .S(n13074), .Z(
        n11064) );
  INV_X1 U13640 ( .A(n11064), .ZN(n11067) );
  AOI22_X1 U13641 ( .A1(n14617), .A2(n11065), .B1(n15150), .B2(n12714), .ZN(
        n11066) );
  OAI211_X1 U13642 ( .C1(n15179), .C2(n12916), .A(n11067), .B(n11066), .ZN(
        P3_U3227) );
  XNOR2_X1 U13643 ( .A(n11068), .B(n12437), .ZN(n11069) );
  INV_X1 U13644 ( .A(n11069), .ZN(n15174) );
  NAND2_X1 U13645 ( .A1(n11069), .A2(n12945), .ZN(n11076) );
  NAND2_X1 U13646 ( .A1(n11070), .A2(n12437), .ZN(n11071) );
  NAND2_X1 U13647 ( .A1(n11072), .A2(n11071), .ZN(n11073) );
  NAND2_X1 U13648 ( .A1(n11073), .A2(n15143), .ZN(n11075) );
  AOI22_X1 U13649 ( .A1(n15139), .A2(n12744), .B1(n12742), .B2(n15136), .ZN(
        n11074) );
  NAND3_X1 U13650 ( .A1(n11076), .A2(n11075), .A3(n11074), .ZN(n15175) );
  MUX2_X1 U13651 ( .A(n15175), .B(P3_REG2_REG_5__SCAN_IN), .S(n13074), .Z(
        n11077) );
  INV_X1 U13652 ( .A(n11077), .ZN(n11081) );
  AOI22_X1 U13653 ( .A1(n14617), .A2(n11079), .B1(n15150), .B2(n11078), .ZN(
        n11080) );
  OAI211_X1 U13654 ( .C1(n15174), .C2(n12916), .A(n11081), .B(n11080), .ZN(
        P3_U3228) );
  AOI21_X1 U13655 ( .B1(n11084), .B2(n11083), .A(n11082), .ZN(n14859) );
  XNOR2_X1 U13656 ( .A(n14857), .B(P2_REG2_REG_12__SCAN_IN), .ZN(n14858) );
  OAI22_X1 U13657 ( .A1(n14859), .A2(n14858), .B1(n14857), .B2(
        P2_REG2_REG_12__SCAN_IN), .ZN(n14874) );
  XNOR2_X1 U13658 ( .A(n14878), .B(P2_REG2_REG_13__SCAN_IN), .ZN(n14875) );
  NOR2_X1 U13659 ( .A1(n14874), .A2(n14875), .ZN(n14873) );
  AOI21_X1 U13660 ( .B1(P2_REG2_REG_13__SCAN_IN), .B2(n14878), .A(n14873), 
        .ZN(n11085) );
  NOR2_X1 U13661 ( .A1(n11085), .A2(n11088), .ZN(n13393) );
  AOI211_X1 U13662 ( .C1(n11572), .C2(n11086), .A(n14907), .B(n13392), .ZN(
        n11105) );
  INV_X1 U13663 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n11103) );
  NAND2_X1 U13664 ( .A1(n11088), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n11087) );
  OAI21_X1 U13665 ( .B1(n11088), .B2(P2_REG1_REG_14__SCAN_IN), .A(n11087), 
        .ZN(n11100) );
  NAND2_X1 U13666 ( .A1(n11089), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n11090) );
  NAND2_X1 U13667 ( .A1(n11091), .A2(n11090), .ZN(n14861) );
  NAND2_X1 U13668 ( .A1(n14857), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n11092) );
  OAI21_X1 U13669 ( .B1(n14857), .B2(P2_REG1_REG_12__SCAN_IN), .A(n11092), 
        .ZN(n14860) );
  NAND2_X1 U13670 ( .A1(n11094), .A2(n11093), .ZN(n11095) );
  NAND2_X1 U13671 ( .A1(n14863), .A2(n11095), .ZN(n14871) );
  INV_X1 U13672 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n11096) );
  MUX2_X1 U13673 ( .A(n11096), .B(P2_REG1_REG_13__SCAN_IN), .S(n14878), .Z(
        n14872) );
  NAND2_X1 U13674 ( .A1(n14878), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n11097) );
  NAND2_X1 U13675 ( .A1(n14869), .A2(n11097), .ZN(n11099) );
  INV_X1 U13676 ( .A(n13401), .ZN(n11098) );
  OAI211_X1 U13677 ( .C1(n11100), .C2(n11099), .A(n11098), .B(n14846), .ZN(
        n11102) );
  AND2_X1 U13678 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3088), .ZN(n11670) );
  AOI21_X1 U13679 ( .B1(n14914), .B2(n13402), .A(n11670), .ZN(n11101) );
  OAI211_X1 U13680 ( .C1(n14932), .C2(n11103), .A(n11102), .B(n11101), .ZN(
        n11104) );
  OR2_X1 U13681 ( .A1(n11105), .A2(n11104), .ZN(P2_U3228) );
  AND2_X1 U13682 ( .A1(n11107), .A2(n11106), .ZN(n12708) );
  XNOR2_X1 U13683 ( .A(n11108), .B(n12742), .ZN(n12707) );
  NAND2_X1 U13684 ( .A1(n12708), .A2(n12707), .ZN(n12706) );
  NAND2_X1 U13685 ( .A1(n12706), .A2(n11109), .ZN(n11291) );
  XNOR2_X1 U13686 ( .A(n11291), .B(n11110), .ZN(n11117) );
  NAND2_X1 U13687 ( .A1(n12724), .A2(n11179), .ZN(n11115) );
  INV_X1 U13688 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n11111) );
  NOR2_X1 U13689 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11111), .ZN(n12335) );
  AOI21_X1 U13690 ( .B1(n12709), .B2(n12742), .A(n12335), .ZN(n11114) );
  NAND2_X1 U13691 ( .A1(n12728), .A2(n12740), .ZN(n11113) );
  NAND2_X1 U13692 ( .A1(n12702), .A2(n11180), .ZN(n11112) );
  NAND4_X1 U13693 ( .A1(n11115), .A2(n11114), .A3(n11113), .A4(n11112), .ZN(
        n11116) );
  AOI21_X1 U13694 ( .B1(n11117), .B2(n12722), .A(n11116), .ZN(n11118) );
  INV_X1 U13695 ( .A(n11118), .ZN(P3_U3153) );
  NAND2_X1 U13696 ( .A1(n11119), .A2(n12722), .ZN(n11129) );
  AOI21_X1 U13697 ( .B1(n11122), .B2(n11121), .A(n11120), .ZN(n11128) );
  INV_X1 U13698 ( .A(n12728), .ZN(n12691) );
  NAND2_X1 U13699 ( .A1(n12724), .A2(n11452), .ZN(n11125) );
  AOI21_X1 U13700 ( .B1(n12709), .B2(n12739), .A(n11123), .ZN(n11124) );
  OAI211_X1 U13701 ( .C1(n11624), .C2(n12691), .A(n11125), .B(n11124), .ZN(
        n11126) );
  AOI21_X1 U13702 ( .B1(n11456), .B2(n12702), .A(n11126), .ZN(n11127) );
  OAI21_X1 U13703 ( .B1(n11129), .B2(n11128), .A(n11127), .ZN(P3_U3157) );
  INV_X1 U13704 ( .A(SI_22_), .ZN(n11130) );
  AOI22_X1 U13705 ( .A1(n12416), .A2(P3_STATE_REG_SCAN_IN), .B1(n11130), .B2(
        n13200), .ZN(n11131) );
  OAI21_X1 U13706 ( .B1(n11132), .B2(n13213), .A(n11131), .ZN(n11133) );
  INV_X1 U13707 ( .A(n11133), .ZN(P3_U3273) );
  INV_X1 U13708 ( .A(n11134), .ZN(n12609) );
  INV_X1 U13709 ( .A(n10529), .ZN(n12285) );
  OAI222_X1 U13710 ( .A1(n13768), .A2(n11135), .B1(n6551), .B2(n12609), .C1(
        P2_U3088), .C2(n12285), .ZN(P2_U3306) );
  INV_X1 U13711 ( .A(n11136), .ZN(n11139) );
  INV_X1 U13712 ( .A(n11137), .ZN(n11138) );
  NAND2_X1 U13713 ( .A1(n11139), .A2(n11138), .ZN(n11140) );
  XNOR2_X1 U13714 ( .A(n12081), .B(n13282), .ZN(n11403) );
  NAND2_X1 U13715 ( .A1(n10574), .A2(n13364), .ZN(n11401) );
  XNOR2_X1 U13716 ( .A(n11403), .B(n11401), .ZN(n11399) );
  XNOR2_X1 U13717 ( .A(n11400), .B(n11399), .ZN(n11146) );
  OAI22_X1 U13718 ( .A1(n13328), .A2(n12077), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9302), .ZN(n11144) );
  OAI22_X1 U13719 ( .A1(n13329), .A2(n11428), .B1(n13344), .B2(n11270), .ZN(
        n11143) );
  AOI211_X1 U13720 ( .C1(n12081), .C2(n13346), .A(n11144), .B(n11143), .ZN(
        n11145) );
  OAI21_X1 U13721 ( .B1(n11146), .B2(n13348), .A(n11145), .ZN(P2_U3208) );
  NAND2_X1 U13722 ( .A1(n11164), .A2(n11980), .ZN(n11148) );
  NAND2_X1 U13723 ( .A1(n13934), .A2(n11975), .ZN(n11147) );
  NAND2_X1 U13724 ( .A1(n11148), .A2(n11147), .ZN(n11150) );
  XNOR2_X1 U13725 ( .A(n11150), .B(n8150), .ZN(n11234) );
  NOR2_X1 U13726 ( .A1(n11938), .A2(n11240), .ZN(n11151) );
  AOI21_X1 U13727 ( .B1(n11164), .B2(n11975), .A(n11151), .ZN(n11233) );
  XNOR2_X1 U13728 ( .A(n11234), .B(n11233), .ZN(n11159) );
  INV_X1 U13729 ( .A(n11152), .ZN(n11153) );
  NAND2_X1 U13730 ( .A1(n11154), .A2(n11153), .ZN(n11155) );
  INV_X1 U13731 ( .A(n11368), .ZN(n11157) );
  AOI21_X1 U13732 ( .B1(n11159), .B2(n11158), .A(n11157), .ZN(n11166) );
  AOI22_X1 U13733 ( .A1(n13818), .A2(n11160), .B1(P1_REG3_REG_8__SCAN_IN), 
        .B2(P1_U3086), .ZN(n11161) );
  OAI21_X1 U13734 ( .B1(n14684), .B2(n11162), .A(n11161), .ZN(n11163) );
  AOI21_X1 U13735 ( .B1(n11164), .B2(n14679), .A(n11163), .ZN(n11165) );
  OAI21_X1 U13736 ( .B1(n11166), .B2(n14674), .A(n11165), .ZN(P1_U3221) );
  INV_X1 U13737 ( .A(n11167), .ZN(n11168) );
  OAI222_X1 U13738 ( .A1(n13768), .A2(n15312), .B1(n6551), .B2(n11168), .C1(
        n12000), .C2(P2_U3088), .ZN(P2_U3305) );
  XNOR2_X1 U13739 ( .A(n11169), .B(n12450), .ZN(n11173) );
  INV_X1 U13740 ( .A(n11173), .ZN(n15184) );
  NAND2_X1 U13741 ( .A1(n12742), .A2(n15139), .ZN(n11171) );
  NAND2_X1 U13742 ( .A1(n12740), .A2(n15136), .ZN(n11170) );
  NAND2_X1 U13743 ( .A1(n11171), .A2(n11170), .ZN(n11172) );
  AOI21_X1 U13744 ( .B1(n11173), .B2(n12945), .A(n11172), .ZN(n11177) );
  XNOR2_X1 U13745 ( .A(n11174), .B(n12450), .ZN(n11175) );
  NAND2_X1 U13746 ( .A1(n11175), .A2(n15143), .ZN(n11176) );
  NAND2_X1 U13747 ( .A1(n11177), .A2(n11176), .ZN(n15185) );
  MUX2_X1 U13748 ( .A(n15185), .B(P3_REG2_REG_7__SCAN_IN), .S(n13074), .Z(
        n11178) );
  INV_X1 U13749 ( .A(n11178), .ZN(n11182) );
  AOI22_X1 U13750 ( .A1(n14617), .A2(n11180), .B1(n15150), .B2(n11179), .ZN(
        n11181) );
  OAI211_X1 U13751 ( .C1(n15184), .C2(n12916), .A(n11182), .B(n11181), .ZN(
        P3_U3226) );
  OAI21_X1 U13752 ( .B1(n11184), .B2(n11186), .A(n11183), .ZN(n11221) );
  INV_X1 U13753 ( .A(n11221), .ZN(n11194) );
  AOI211_X1 U13754 ( .C1(n11186), .C2(n11185), .A(n14761), .B(n6666), .ZN(
        n11219) );
  NAND2_X1 U13755 ( .A1(n14757), .A2(n13933), .ZN(n11217) );
  INV_X1 U13756 ( .A(n11217), .ZN(n11187) );
  OAI21_X1 U13757 ( .B1(n11219), .B2(n11187), .A(n14256), .ZN(n11193) );
  OAI22_X1 U13758 ( .A1(n14256), .A2(n11188), .B1(n11377), .B2(n14777), .ZN(
        n11191) );
  OAI211_X1 U13759 ( .C1(n7012), .C2(n7013), .A(n14365), .B(n11281), .ZN(
        n11218) );
  NAND2_X1 U13760 ( .A1(n14247), .A2(n13931), .ZN(n11216) );
  AOI21_X1 U13761 ( .B1(n11218), .B2(n11216), .A(n14261), .ZN(n11190) );
  AOI211_X1 U13762 ( .C1(n14258), .C2(n11373), .A(n11191), .B(n11190), .ZN(
        n11192) );
  OAI211_X1 U13763 ( .C1(n11194), .C2(n14286), .A(n11193), .B(n11192), .ZN(
        P1_U3283) );
  OR2_X1 U13764 ( .A1(n11195), .A2(n12385), .ZN(n11196) );
  NAND2_X1 U13765 ( .A1(n11197), .A2(n11196), .ZN(n15164) );
  OAI22_X1 U13766 ( .A1(n14613), .A2(n15161), .B1(P3_REG3_REG_3__SCAN_IN), 
        .B2(n15118), .ZN(n11205) );
  NAND2_X1 U13767 ( .A1(n15164), .A2(n12945), .ZN(n11203) );
  AOI22_X1 U13768 ( .A1(n15139), .A2(n15137), .B1(n12744), .B2(n15136), .ZN(
        n11202) );
  NAND2_X1 U13769 ( .A1(n11198), .A2(n12385), .ZN(n11199) );
  NAND3_X1 U13770 ( .A1(n11200), .A2(n15143), .A3(n11199), .ZN(n11201) );
  NAND3_X1 U13771 ( .A1(n11203), .A2(n11202), .A3(n11201), .ZN(n15162) );
  MUX2_X1 U13772 ( .A(n15162), .B(P3_REG2_REG_3__SCAN_IN), .S(n13074), .Z(
        n11204) );
  AOI211_X1 U13773 ( .C1(n15151), .C2(n15164), .A(n11205), .B(n11204), .ZN(
        n11206) );
  INV_X1 U13774 ( .A(n11206), .ZN(P3_U3230) );
  XNOR2_X1 U13775 ( .A(n11207), .B(n12457), .ZN(n15189) );
  OAI21_X1 U13776 ( .B1(n12457), .B2(n11208), .A(n11341), .ZN(n11209) );
  NAND2_X1 U13777 ( .A1(n11209), .A2(n15143), .ZN(n11211) );
  AOI22_X1 U13778 ( .A1(n15139), .A2(n12741), .B1(n12739), .B2(n15136), .ZN(
        n11210) );
  OAI211_X1 U13779 ( .C1(n15147), .C2(n15189), .A(n11211), .B(n11210), .ZN(
        n15191) );
  NAND2_X1 U13780 ( .A1(n15191), .A2(n15132), .ZN(n11215) );
  INV_X1 U13781 ( .A(n11294), .ZN(n11212) );
  OAI22_X1 U13782 ( .A1(n14613), .A2(n15188), .B1(n11212), .B2(n15118), .ZN(
        n11213) );
  AOI21_X1 U13783 ( .B1(P3_REG2_REG_8__SCAN_IN), .B2(n13074), .A(n11213), .ZN(
        n11214) );
  OAI211_X1 U13784 ( .C1(n15189), .C2(n12916), .A(n11215), .B(n11214), .ZN(
        P3_U3225) );
  AND2_X1 U13785 ( .A1(n11217), .A2(n11216), .ZN(n11378) );
  NAND2_X1 U13786 ( .A1(n11218), .A2(n11378), .ZN(n11220) );
  AOI211_X1 U13787 ( .C1(n14803), .C2(n11221), .A(n11220), .B(n11219), .ZN(
        n11226) );
  INV_X1 U13788 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n11222) );
  OAI22_X1 U13789 ( .A1(n7012), .A2(n14411), .B1(n14806), .B2(n11222), .ZN(
        n11223) );
  INV_X1 U13790 ( .A(n11223), .ZN(n11224) );
  OAI21_X1 U13791 ( .B1(n11226), .B2(n14804), .A(n11224), .ZN(P1_U3489) );
  AOI22_X1 U13792 ( .A1(n11373), .A2(n14341), .B1(n14809), .B2(
        P1_REG1_REG_10__SCAN_IN), .ZN(n11225) );
  OAI21_X1 U13793 ( .B1(n11226), .B2(n14809), .A(n11225), .ZN(P1_U3538) );
  INV_X1 U13794 ( .A(n14679), .ZN(n13875) );
  NAND2_X1 U13795 ( .A1(n11232), .A2(n11980), .ZN(n11228) );
  NAND2_X1 U13796 ( .A1(n13933), .A2(n11975), .ZN(n11227) );
  NAND2_X1 U13797 ( .A1(n11228), .A2(n11227), .ZN(n11229) );
  XNOR2_X1 U13798 ( .A(n11229), .B(n11149), .ZN(n11361) );
  NOR2_X1 U13799 ( .A1(n11938), .A2(n11230), .ZN(n11231) );
  AOI21_X1 U13800 ( .B1(n11232), .B2(n11975), .A(n11231), .ZN(n11362) );
  XNOR2_X1 U13801 ( .A(n11361), .B(n11362), .ZN(n11366) );
  NAND2_X1 U13802 ( .A1(n11234), .A2(n11233), .ZN(n11364) );
  NAND2_X1 U13803 ( .A1(n11368), .A2(n11364), .ZN(n11236) );
  NAND2_X1 U13804 ( .A1(n11236), .A2(n11366), .ZN(n11235) );
  OAI21_X1 U13805 ( .B1(n11366), .B2(n11236), .A(n11235), .ZN(n11237) );
  NAND2_X1 U13806 ( .A1(n11237), .A2(n13880), .ZN(n11244) );
  NOR2_X1 U13807 ( .A1(n14684), .A2(n11238), .ZN(n11242) );
  INV_X1 U13808 ( .A(n13900), .ZN(n14668) );
  OAI22_X1 U13809 ( .A1(n14668), .A2(n11240), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n11239), .ZN(n11241) );
  AOI211_X1 U13810 ( .C1(n14665), .C2(n13932), .A(n11242), .B(n11241), .ZN(
        n11243) );
  OAI211_X1 U13811 ( .C1(n14799), .C2(n13875), .A(n11244), .B(n11243), .ZN(
        P1_U3231) );
  XNOR2_X1 U13812 ( .A(n11484), .B(n11483), .ZN(n11247) );
  NOR2_X1 U13813 ( .A1(n11531), .A2(n11247), .ZN(n11485) );
  AOI21_X1 U13814 ( .B1(n11531), .B2(n11247), .A(n11485), .ZN(n11262) );
  INV_X1 U13815 ( .A(n11484), .ZN(n11497) );
  NAND2_X1 U13816 ( .A1(P3_REG1_REG_11__SCAN_IN), .A2(n11250), .ZN(n11491) );
  OAI21_X1 U13817 ( .B1(P3_REG1_REG_11__SCAN_IN), .B2(n11250), .A(n11491), 
        .ZN(n11260) );
  INV_X1 U13818 ( .A(P3_REG3_REG_11__SCAN_IN), .ZN(n15413) );
  NOR2_X1 U13819 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15413), .ZN(n11519) );
  AOI21_X1 U13820 ( .B1(n15106), .B2(P3_ADDR_REG_11__SCAN_IN), .A(n11519), 
        .ZN(n11251) );
  OAI21_X1 U13821 ( .B1(n15100), .B2(n11497), .A(n11251), .ZN(n11259) );
  INV_X1 U13822 ( .A(n11252), .ZN(n11253) );
  MUX2_X1 U13823 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n13209), .Z(n11498) );
  XNOR2_X1 U13824 ( .A(n11498), .B(n11497), .ZN(n11255) );
  AOI21_X1 U13825 ( .B1(n11256), .B2(n11255), .A(n11500), .ZN(n11257) );
  NOR2_X1 U13826 ( .A1(n11257), .A2(n15102), .ZN(n11258) );
  AOI211_X1 U13827 ( .C1(n15109), .C2(n11260), .A(n11259), .B(n11258), .ZN(
        n11261) );
  OAI21_X1 U13828 ( .B1(n11262), .B2(n15113), .A(n11261), .ZN(P3_U3193) );
  XOR2_X1 U13829 ( .A(n12262), .B(n11263), .Z(n11387) );
  INV_X1 U13830 ( .A(n11387), .ZN(n11276) );
  INV_X1 U13831 ( .A(n11264), .ZN(n11265) );
  AOI21_X1 U13832 ( .B1(n12262), .B2(n11266), .A(n11265), .ZN(n11267) );
  OAI222_X1 U13833 ( .A1(n13548), .A2(n11428), .B1(n13627), .B2(n12077), .C1(
        n13600), .C2(n11267), .ZN(n11385) );
  INV_X1 U13834 ( .A(n12081), .ZN(n11390) );
  AOI21_X1 U13835 ( .B1(n11268), .B2(n12081), .A(n10574), .ZN(n11269) );
  AND2_X1 U13836 ( .A1(n11269), .A2(n11310), .ZN(n11386) );
  NAND2_X1 U13837 ( .A1(n11386), .A2(n13613), .ZN(n11273) );
  INV_X1 U13838 ( .A(n11270), .ZN(n11271) );
  AOI22_X1 U13839 ( .A1(n14947), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n14936), 
        .B2(n11271), .ZN(n11272) );
  OAI211_X1 U13840 ( .C1(n11390), .C2(n13610), .A(n11273), .B(n11272), .ZN(
        n11274) );
  AOI21_X1 U13841 ( .B1(n11385), .B2(n13602), .A(n11274), .ZN(n11275) );
  OAI21_X1 U13842 ( .B1(n11276), .B2(n14942), .A(n11275), .ZN(P2_U3254) );
  XNOR2_X1 U13843 ( .A(n11277), .B(n7512), .ZN(n11278) );
  OAI222_X1 U13844 ( .A1(n14770), .A2(n11597), .B1(n14276), .B2(n11550), .C1(
        n11278), .C2(n14761), .ZN(n14687) );
  INV_X1 U13845 ( .A(n14687), .ZN(n11289) );
  OAI21_X1 U13846 ( .B1(n11280), .B2(n11279), .A(n11461), .ZN(n14689) );
  INV_X1 U13847 ( .A(n11555), .ZN(n14686) );
  INV_X1 U13848 ( .A(n11281), .ZN(n11283) );
  INV_X1 U13849 ( .A(n11282), .ZN(n11471) );
  OAI211_X1 U13850 ( .C1(n14686), .C2(n11283), .A(n11471), .B(n14365), .ZN(
        n14685) );
  OAI22_X1 U13851 ( .A1(n14256), .A2(n11284), .B1(n11553), .B2(n14777), .ZN(
        n11285) );
  AOI21_X1 U13852 ( .B1(n11555), .B2(n14258), .A(n11285), .ZN(n11286) );
  OAI21_X1 U13853 ( .B1(n14685), .B2(n14261), .A(n11286), .ZN(n11287) );
  AOI21_X1 U13854 ( .B1(n14689), .B2(n14235), .A(n11287), .ZN(n11288) );
  OAI21_X1 U13855 ( .B1(n11289), .B2(n14281), .A(n11288), .ZN(P1_U3282) );
  MUX2_X1 U13856 ( .A(n12741), .B(n11291), .S(n11290), .Z(n11293) );
  XNOR2_X1 U13857 ( .A(n11293), .B(n11292), .ZN(n11300) );
  NAND2_X1 U13858 ( .A1(n12724), .A2(n11294), .ZN(n11298) );
  AND2_X1 U13859 ( .A1(P3_U3151), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n12321) );
  AOI21_X1 U13860 ( .B1(n12709), .B2(n12741), .A(n12321), .ZN(n11297) );
  NAND2_X1 U13861 ( .A1(n12702), .A2(n12460), .ZN(n11296) );
  NAND2_X1 U13862 ( .A1(n12728), .A2(n12739), .ZN(n11295) );
  NAND4_X1 U13863 ( .A1(n11298), .A2(n11297), .A3(n11296), .A4(n11295), .ZN(
        n11299) );
  AOI21_X1 U13864 ( .B1(n11300), .B2(n12722), .A(n11299), .ZN(n11301) );
  INV_X1 U13865 ( .A(n11301), .ZN(P3_U3161) );
  INV_X1 U13866 ( .A(n11302), .ZN(n11303) );
  AOI21_X1 U13867 ( .B1(n9323), .B2(n11304), .A(n11303), .ZN(n14655) );
  AOI22_X1 U13868 ( .A1(n13462), .A2(n13364), .B1(n13496), .B2(n13362), .ZN(
        n11308) );
  OAI211_X1 U13869 ( .C1(n11306), .C2(n9323), .A(n13618), .B(n11305), .ZN(
        n11307) );
  OAI211_X1 U13870 ( .C1(n14655), .C2(n13624), .A(n11308), .B(n11307), .ZN(
        n14658) );
  NAND2_X1 U13871 ( .A1(n14658), .A2(n13602), .ZN(n11316) );
  OAI22_X1 U13872 ( .A1(n13602), .A2(n11309), .B1(n11409), .B2(n13535), .ZN(
        n11314) );
  INV_X1 U13873 ( .A(n12087), .ZN(n14657) );
  INV_X1 U13874 ( .A(n11310), .ZN(n11312) );
  INV_X1 U13875 ( .A(n11311), .ZN(n11419) );
  OAI211_X1 U13876 ( .C1(n14657), .C2(n11312), .A(n13603), .B(n11419), .ZN(
        n14656) );
  NOR2_X1 U13877 ( .A1(n14656), .A2(n14939), .ZN(n11313) );
  AOI211_X1 U13878 ( .C1(n14935), .C2(n12087), .A(n11314), .B(n11313), .ZN(
        n11315) );
  OAI211_X1 U13879 ( .C1(n14655), .C2(n11317), .A(n11316), .B(n11315), .ZN(
        P2_U3253) );
  OAI21_X1 U13880 ( .B1(P1_REG1_REG_14__SCAN_IN), .B2(n11319), .A(n11318), 
        .ZN(n11320) );
  INV_X1 U13881 ( .A(n11320), .ZN(n11321) );
  XNOR2_X1 U13882 ( .A(n11320), .B(n11327), .ZN(n14741) );
  NAND2_X1 U13883 ( .A1(n14741), .A2(n14740), .ZN(n14739) );
  OAI21_X1 U13884 ( .B1(n11321), .B2(n11327), .A(n14739), .ZN(n11323) );
  XNOR2_X1 U13885 ( .A(n11561), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n11322) );
  NOR2_X1 U13886 ( .A1(n11322), .A2(n11323), .ZN(n11560) );
  AOI211_X1 U13887 ( .C1(n11323), .C2(n11322), .A(n11560), .B(n14040), .ZN(
        n11338) );
  OAI21_X1 U13888 ( .B1(n11326), .B2(n11325), .A(n11324), .ZN(n11328) );
  INV_X1 U13889 ( .A(n11328), .ZN(n11329) );
  XNOR2_X1 U13890 ( .A(n11328), .B(n11327), .ZN(n14743) );
  NOR2_X1 U13891 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n14743), .ZN(n14742) );
  AOI21_X1 U13892 ( .B1(n11329), .B2(n14745), .A(n14742), .ZN(n11332) );
  OR2_X1 U13893 ( .A1(n11561), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n11330) );
  NAND2_X1 U13894 ( .A1(n11561), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n11559) );
  AND2_X1 U13895 ( .A1(n11330), .A2(n11559), .ZN(n11331) );
  NAND2_X1 U13896 ( .A1(n11331), .A2(n11332), .ZN(n11558) );
  OAI211_X1 U13897 ( .C1(n11332), .C2(n11331), .A(n14059), .B(n11558), .ZN(
        n11335) );
  NAND2_X1 U13898 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n13834)
         );
  INV_X1 U13899 ( .A(n13834), .ZN(n11333) );
  AOI21_X1 U13900 ( .B1(n14719), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n11333), 
        .ZN(n11334) );
  OAI211_X1 U13901 ( .C1(n14744), .C2(n11336), .A(n11335), .B(n11334), .ZN(
        n11337) );
  OR2_X1 U13902 ( .A1(n11338), .A2(n11337), .ZN(P1_U3259) );
  XNOR2_X1 U13903 ( .A(n11339), .B(n12465), .ZN(n15195) );
  AND2_X1 U13904 ( .A1(n11341), .A2(n11340), .ZN(n11343) );
  OAI211_X1 U13905 ( .C1(n11343), .C2(n12465), .A(n15143), .B(n11342), .ZN(
        n11345) );
  AOI22_X1 U13906 ( .A1(n15139), .A2(n12740), .B1(n12738), .B2(n15136), .ZN(
        n11344) );
  OAI211_X1 U13907 ( .C1(n15147), .C2(n15195), .A(n11345), .B(n11344), .ZN(
        n15197) );
  NAND2_X1 U13908 ( .A1(n15197), .A2(n15132), .ZN(n11349) );
  OAI22_X1 U13909 ( .A1(n14613), .A2(n15193), .B1(n11346), .B2(n15118), .ZN(
        n11347) );
  AOI21_X1 U13910 ( .B1(P3_REG2_REG_9__SCAN_IN), .B2(n13074), .A(n11347), .ZN(
        n11348) );
  OAI211_X1 U13911 ( .C1(n15195), .C2(n12916), .A(n11349), .B(n11348), .ZN(
        P3_U3224) );
  XNOR2_X1 U13912 ( .A(n11350), .B(n11351), .ZN(n14386) );
  NAND2_X1 U13913 ( .A1(n14256), .A2(n14783), .ZN(n14237) );
  OAI21_X1 U13914 ( .B1(n11354), .B2(n11353), .A(n11352), .ZN(n14384) );
  INV_X1 U13915 ( .A(n11355), .ZN(n11470) );
  INV_X1 U13916 ( .A(n11736), .ZN(n14382) );
  OAI211_X1 U13917 ( .C1(n11470), .C2(n14382), .A(n14365), .B(n11635), .ZN(
        n14381) );
  AOI22_X1 U13918 ( .A1(n14757), .A2(n13930), .B1(n14247), .B2(n13928), .ZN(
        n14380) );
  OAI22_X1 U13919 ( .A1(n14281), .A2(n14380), .B1(n11739), .B2(n14777), .ZN(
        n11357) );
  NOR2_X1 U13920 ( .A1(n14382), .A2(n14271), .ZN(n11356) );
  AOI211_X1 U13921 ( .C1(n14281), .C2(P1_REG2_REG_13__SCAN_IN), .A(n11357), 
        .B(n11356), .ZN(n11358) );
  OAI21_X1 U13922 ( .B1(n14261), .B2(n14381), .A(n11358), .ZN(n11359) );
  AOI21_X1 U13923 ( .B1(n14384), .B2(n14235), .A(n11359), .ZN(n11360) );
  OAI21_X1 U13924 ( .B1(n14386), .B2(n14237), .A(n11360), .ZN(P1_U3280) );
  INV_X1 U13925 ( .A(n11361), .ZN(n11363) );
  NAND2_X1 U13926 ( .A1(n11363), .A2(n11362), .ZN(n11365) );
  INV_X1 U13927 ( .A(n11365), .ZN(n11367) );
  NAND2_X1 U13928 ( .A1(n11373), .A2(n11980), .ZN(n11370) );
  NAND2_X1 U13929 ( .A1(n13932), .A2(n11975), .ZN(n11369) );
  NAND2_X1 U13930 ( .A1(n11370), .A2(n11369), .ZN(n11371) );
  XNOR2_X1 U13931 ( .A(n11371), .B(n8150), .ZN(n11539) );
  NOR2_X1 U13932 ( .A1(n11938), .A2(n11550), .ZN(n11372) );
  AOI21_X1 U13933 ( .B1(n11373), .B2(n11975), .A(n11372), .ZN(n11540) );
  XNOR2_X1 U13934 ( .A(n11539), .B(n11540), .ZN(n11374) );
  AOI21_X1 U13935 ( .B1(n11375), .B2(n11374), .A(n14674), .ZN(n11376) );
  NAND2_X1 U13936 ( .A1(n11376), .A2(n11544), .ZN(n11382) );
  INV_X1 U13937 ( .A(n11377), .ZN(n11380) );
  INV_X1 U13938 ( .A(n14684), .ZN(n13891) );
  OAI22_X1 U13939 ( .A1(n13870), .A2(n11378), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7838), .ZN(n11379) );
  AOI21_X1 U13940 ( .B1(n11380), .B2(n13891), .A(n11379), .ZN(n11381) );
  OAI211_X1 U13941 ( .C1(n7012), .C2(n13875), .A(n11382), .B(n11381), .ZN(
        P1_U3217) );
  NAND2_X1 U13942 ( .A1(n11383), .A2(n13202), .ZN(n11384) );
  OAI211_X1 U13943 ( .C1(n7377), .C2(n13217), .A(n11384), .B(n12586), .ZN(
        P3_U3272) );
  AOI211_X1 U13944 ( .C1(n14983), .C2(n11387), .A(n11386), .B(n11385), .ZN(
        n11393) );
  AOI22_X1 U13945 ( .A1(n12081), .A2(n11388), .B1(n15017), .B2(
        P2_REG1_REG_11__SCAN_IN), .ZN(n11389) );
  OAI21_X1 U13946 ( .B1(n11393), .B2(n15017), .A(n11389), .ZN(P2_U3510) );
  OAI22_X1 U13947 ( .A1(n11390), .A2(n13764), .B1(n15007), .B2(n9301), .ZN(
        n11391) );
  INV_X1 U13948 ( .A(n11391), .ZN(n11392) );
  OAI21_X1 U13949 ( .B1(n11393), .B2(n15005), .A(n11392), .ZN(P2_U3463) );
  XNOR2_X1 U13950 ( .A(n12087), .B(n13236), .ZN(n11394) );
  NAND2_X1 U13951 ( .A1(n10574), .A2(n13363), .ZN(n11395) );
  NAND2_X1 U13952 ( .A1(n11394), .A2(n11395), .ZN(n11426) );
  INV_X1 U13953 ( .A(n11394), .ZN(n11397) );
  INV_X1 U13954 ( .A(n11395), .ZN(n11396) );
  NAND2_X1 U13955 ( .A1(n11397), .A2(n11396), .ZN(n11398) );
  NAND2_X1 U13956 ( .A1(n11426), .A2(n11398), .ZN(n11407) );
  INV_X1 U13957 ( .A(n11401), .ZN(n11402) );
  NAND2_X1 U13958 ( .A1(n11403), .A2(n11402), .ZN(n11404) );
  INV_X1 U13959 ( .A(n11427), .ZN(n11405) );
  AOI21_X1 U13960 ( .B1(n11407), .B2(n11406), .A(n11405), .ZN(n11413) );
  INV_X1 U13961 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n11408) );
  NOR2_X1 U13962 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n11408), .ZN(n14856) );
  OAI22_X1 U13963 ( .A1(n13329), .A2(n12094), .B1(n13344), .B2(n11409), .ZN(
        n11410) );
  AOI211_X1 U13964 ( .C1(n11671), .C2(n13364), .A(n14856), .B(n11410), .ZN(
        n11412) );
  NAND2_X1 U13965 ( .A1(n12087), .A2(n13346), .ZN(n11411) );
  OAI211_X1 U13966 ( .C1(n11413), .C2(n13348), .A(n11412), .B(n11411), .ZN(
        P2_U3196) );
  XNOR2_X1 U13967 ( .A(n11415), .B(n11414), .ZN(n11416) );
  OAI222_X1 U13968 ( .A1(n13548), .A2(n11430), .B1(n13627), .B2(n11428), .C1(
        n11416), .C2(n13600), .ZN(n11609) );
  INV_X1 U13969 ( .A(n11609), .ZN(n11425) );
  XNOR2_X1 U13970 ( .A(n11417), .B(n12264), .ZN(n11611) );
  INV_X1 U13971 ( .A(n11418), .ZN(n11571) );
  AOI211_X1 U13972 ( .C1(n12092), .C2(n11419), .A(n10574), .B(n11571), .ZN(
        n11610) );
  NAND2_X1 U13973 ( .A1(n11610), .A2(n13613), .ZN(n11422) );
  INV_X1 U13974 ( .A(n11429), .ZN(n11420) );
  AOI22_X1 U13975 ( .A1(n14947), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n14936), 
        .B2(n11420), .ZN(n11421) );
  OAI211_X1 U13976 ( .C1(n9580), .C2(n13610), .A(n11422), .B(n11421), .ZN(
        n11423) );
  AOI21_X1 U13977 ( .B1(n13579), .B2(n11611), .A(n11423), .ZN(n11424) );
  OAI21_X1 U13978 ( .B1(n11425), .B2(n14947), .A(n11424), .ZN(P2_U3252) );
  XNOR2_X1 U13979 ( .A(n12092), .B(n13236), .ZN(n11661) );
  NAND2_X1 U13980 ( .A1(n10574), .A2(n13362), .ZN(n11662) );
  XNOR2_X1 U13981 ( .A(n11661), .B(n11662), .ZN(n11659) );
  XNOR2_X1 U13982 ( .A(n11660), .B(n11659), .ZN(n11434) );
  OAI22_X1 U13983 ( .A1(n13328), .A2(n11428), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9343), .ZN(n11432) );
  OAI22_X1 U13984 ( .A1(n13329), .A2(n11430), .B1(n13344), .B2(n11429), .ZN(
        n11431) );
  AOI211_X1 U13985 ( .C1(n12092), .C2(n13346), .A(n11432), .B(n11431), .ZN(
        n11433) );
  OAI21_X1 U13986 ( .B1(n11434), .B2(n13348), .A(n11433), .ZN(P2_U3206) );
  XNOR2_X1 U13987 ( .A(n11435), .B(n11789), .ZN(n11436) );
  XNOR2_X1 U13988 ( .A(n11437), .B(n11436), .ZN(n11445) );
  INV_X1 U13989 ( .A(n14625), .ZN(n11724) );
  INV_X1 U13990 ( .A(n11438), .ZN(n11721) );
  NOR2_X1 U13991 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11439), .ZN(n12759) );
  NOR2_X1 U13992 ( .A1(n11720), .A2(n12726), .ZN(n11440) );
  AOI211_X1 U13993 ( .C1(n12728), .C2(n11441), .A(n12759), .B(n11440), .ZN(
        n11442) );
  OAI21_X1 U13994 ( .B1(n11721), .B2(n12700), .A(n11442), .ZN(n11443) );
  AOI21_X1 U13995 ( .B1(n11724), .B2(n12702), .A(n11443), .ZN(n11444) );
  OAI21_X1 U13996 ( .B1(n11445), .B2(n12704), .A(n11444), .ZN(P3_U3174) );
  INV_X1 U13997 ( .A(n12469), .ZN(n12390) );
  XNOR2_X1 U13998 ( .A(n11446), .B(n12390), .ZN(n15202) );
  NAND2_X1 U13999 ( .A1(n15147), .A2(n11447), .ZN(n11448) );
  INV_X1 U14000 ( .A(n13077), .ZN(n11795) );
  INV_X1 U14001 ( .A(n12739), .ZN(n11451) );
  XNOR2_X1 U14002 ( .A(n11449), .B(n12469), .ZN(n11450) );
  OAI222_X1 U14003 ( .A1(n13069), .A2(n11624), .B1(n13067), .B2(n11451), .C1(
        n11450), .C2(n13064), .ZN(n15204) );
  NAND2_X1 U14004 ( .A1(n15204), .A2(n15132), .ZN(n11458) );
  INV_X1 U14005 ( .A(n11452), .ZN(n11453) );
  OAI22_X1 U14006 ( .A1(n15132), .A2(n11454), .B1(n11453), .B2(n15118), .ZN(
        n11455) );
  AOI21_X1 U14007 ( .B1(n11456), .B2(n14617), .A(n11455), .ZN(n11457) );
  OAI211_X1 U14008 ( .C1(n15202), .C2(n11795), .A(n11458), .B(n11457), .ZN(
        P3_U3223) );
  NAND2_X1 U14009 ( .A1(n11459), .A2(n14783), .ZN(n11466) );
  INV_X1 U14010 ( .A(n11459), .ZN(n11463) );
  NOR2_X1 U14011 ( .A1(n7510), .A2(n14755), .ZN(n11462) );
  AOI22_X1 U14012 ( .A1(n11463), .A2(n14783), .B1(n11462), .B2(n11461), .ZN(
        n11465) );
  MUX2_X1 U14013 ( .A(n11466), .B(n11465), .S(n11464), .Z(n11468) );
  AOI22_X1 U14014 ( .A1(n14757), .A2(n13931), .B1(n14247), .B2(n13929), .ZN(
        n11467) );
  OAI211_X1 U14015 ( .C1(n11469), .C2(n14755), .A(n11468), .B(n11467), .ZN(
        n11509) );
  INV_X1 U14016 ( .A(n11509), .ZN(n11476) );
  AOI211_X1 U14017 ( .C1(n11599), .C2(n11471), .A(n14793), .B(n11470), .ZN(
        n11508) );
  NOR2_X1 U14018 ( .A1(n11608), .A2(n14271), .ZN(n11474) );
  OAI22_X1 U14019 ( .A1(n14256), .A2(n11472), .B1(n11602), .B2(n14777), .ZN(
        n11473) );
  AOI211_X1 U14020 ( .C1(n11508), .C2(n14284), .A(n11474), .B(n11473), .ZN(
        n11475) );
  OAI21_X1 U14021 ( .B1(n11476), .B2(n14281), .A(n11475), .ZN(P1_U3281) );
  NAND2_X1 U14022 ( .A1(n11480), .A2(n14425), .ZN(n11478) );
  OAI211_X1 U14023 ( .C1(n11479), .C2(n14433), .A(n11478), .B(n11477), .ZN(
        P1_U3332) );
  NAND2_X1 U14024 ( .A1(n11480), .A2(n13775), .ZN(n11482) );
  NOR2_X1 U14025 ( .A1(n11481), .A2(P2_U3088), .ZN(n12298) );
  INV_X1 U14026 ( .A(n12298), .ZN(n12308) );
  OAI211_X1 U14027 ( .C1(n15252), .C2(n13768), .A(n11482), .B(n12308), .ZN(
        P2_U3304) );
  NOR2_X1 U14028 ( .A1(n11484), .A2(n11483), .ZN(n11486) );
  NOR2_X1 U14029 ( .A1(n11486), .A2(n11485), .ZN(n11489) );
  MUX2_X1 U14030 ( .A(P3_REG2_REG_12__SCAN_IN), .B(n12746), .S(n12751), .Z(
        n11488) );
  OR2_X2 U14031 ( .A1(n11489), .A2(n11488), .ZN(n12748) );
  INV_X1 U14032 ( .A(n12748), .ZN(n11487) );
  AOI21_X1 U14033 ( .B1(n11489), .B2(n11488), .A(n11487), .ZN(n11507) );
  NAND2_X1 U14034 ( .A1(n11497), .A2(n11490), .ZN(n11492) );
  INV_X1 U14035 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n11493) );
  MUX2_X1 U14036 ( .A(n11493), .B(P3_REG1_REG_12__SCAN_IN), .S(n12751), .Z(
        n11494) );
  OAI21_X1 U14037 ( .B1(n11495), .B2(n11494), .A(n12750), .ZN(n11505) );
  INV_X1 U14038 ( .A(n12751), .ZN(n12754) );
  AND2_X1 U14039 ( .A1(P3_U3151), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n11585) );
  AOI21_X1 U14040 ( .B1(n15106), .B2(P3_ADDR_REG_12__SCAN_IN), .A(n11585), 
        .ZN(n11496) );
  OAI21_X1 U14041 ( .B1(n15100), .B2(n12754), .A(n11496), .ZN(n11504) );
  MUX2_X1 U14042 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n13209), .Z(n12755) );
  XOR2_X1 U14043 ( .A(n12751), .B(n12755), .Z(n11502) );
  NOR2_X1 U14044 ( .A1(n11498), .A2(n11497), .ZN(n11499) );
  OR2_X1 U14045 ( .A1(n11500), .A2(n11499), .ZN(n11501) );
  AOI211_X1 U14046 ( .C1(n11502), .C2(n11501), .A(n15102), .B(n12753), .ZN(
        n11503) );
  AOI211_X1 U14047 ( .C1(n15109), .C2(n11505), .A(n11504), .B(n11503), .ZN(
        n11506) );
  OAI21_X1 U14048 ( .B1(n11507), .B2(n15113), .A(n11506), .ZN(P3_U3194) );
  NOR2_X1 U14049 ( .A1(n11509), .A2(n11508), .ZN(n11512) );
  AOI22_X1 U14050 ( .A1(n11599), .A2(n14416), .B1(P1_REG0_REG_12__SCAN_IN), 
        .B2(n14804), .ZN(n11510) );
  OAI21_X1 U14051 ( .B1(n11512), .B2(n14804), .A(n11510), .ZN(P1_U3495) );
  AOI22_X1 U14052 ( .A1(n11599), .A2(n14341), .B1(P1_REG1_REG_12__SCAN_IN), 
        .B2(n14809), .ZN(n11511) );
  OAI21_X1 U14053 ( .B1(n11512), .B2(n14809), .A(n11511), .ZN(P1_U3540) );
  INV_X1 U14054 ( .A(n11514), .ZN(n11516) );
  INV_X1 U14055 ( .A(n11513), .ZN(n11515) );
  OR2_X1 U14056 ( .A1(n11514), .A2(n11513), .ZN(n11577) );
  OAI21_X1 U14057 ( .B1(n11516), .B2(n11515), .A(n11577), .ZN(n11517) );
  NOR2_X1 U14058 ( .A1(n11517), .A2(n11518), .ZN(n11579) );
  AOI21_X1 U14059 ( .B1(n11518), .B2(n11517), .A(n11579), .ZN(n11524) );
  NAND2_X1 U14060 ( .A1(n12724), .A2(n11529), .ZN(n11521) );
  AOI21_X1 U14061 ( .B1(n12709), .B2(n12738), .A(n11519), .ZN(n11520) );
  OAI211_X1 U14062 ( .C1(n11720), .C2(n12691), .A(n11521), .B(n11520), .ZN(
        n11522) );
  AOI21_X1 U14063 ( .B1(n14637), .B2(n12702), .A(n11522), .ZN(n11523) );
  OAI21_X1 U14064 ( .B1(n11524), .B2(n12704), .A(n11523), .ZN(P3_U3176) );
  INV_X1 U14065 ( .A(n12476), .ZN(n12483) );
  XNOR2_X1 U14066 ( .A(n11525), .B(n12483), .ZN(n14634) );
  INV_X1 U14067 ( .A(n12738), .ZN(n11528) );
  XNOR2_X1 U14068 ( .A(n11526), .B(n12483), .ZN(n11527) );
  OAI222_X1 U14069 ( .A1(n13069), .A2(n11720), .B1(n13067), .B2(n11528), .C1(
        n11527), .C2(n13064), .ZN(n14635) );
  NAND2_X1 U14070 ( .A1(n14635), .A2(n15132), .ZN(n11534) );
  INV_X1 U14071 ( .A(n11529), .ZN(n11530) );
  OAI22_X1 U14072 ( .A1(n15132), .A2(n11531), .B1(n11530), .B2(n15118), .ZN(
        n11532) );
  AOI21_X1 U14073 ( .B1(n14617), .B2(n14637), .A(n11532), .ZN(n11533) );
  OAI211_X1 U14074 ( .C1(n11795), .C2(n14634), .A(n11534), .B(n11533), .ZN(
        P3_U3222) );
  NAND2_X1 U14075 ( .A1(n11555), .A2(n11980), .ZN(n11536) );
  NAND2_X1 U14076 ( .A1(n13931), .A2(n11975), .ZN(n11535) );
  NAND2_X1 U14077 ( .A1(n11536), .A2(n11535), .ZN(n11537) );
  XNOR2_X1 U14078 ( .A(n11537), .B(n8150), .ZN(n11591) );
  NOR2_X1 U14079 ( .A1(n11938), .A2(n11603), .ZN(n11538) );
  AOI21_X1 U14080 ( .B1(n11555), .B2(n11975), .A(n11538), .ZN(n11590) );
  XNOR2_X1 U14081 ( .A(n11591), .B(n11590), .ZN(n11548) );
  INV_X1 U14082 ( .A(n11539), .ZN(n11542) );
  INV_X1 U14083 ( .A(n11540), .ZN(n11541) );
  NAND2_X1 U14084 ( .A1(n11542), .A2(n11541), .ZN(n11543) );
  INV_X1 U14085 ( .A(n11593), .ZN(n11546) );
  AOI21_X1 U14086 ( .B1(n11548), .B2(n11547), .A(n11546), .ZN(n11557) );
  OAI22_X1 U14087 ( .A1(n14668), .A2(n11550), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n11549), .ZN(n11551) );
  AOI21_X1 U14088 ( .B1(n14665), .B2(n13930), .A(n11551), .ZN(n11552) );
  OAI21_X1 U14089 ( .B1(n14684), .B2(n11553), .A(n11552), .ZN(n11554) );
  AOI21_X1 U14090 ( .B1(n11555), .B2(n14679), .A(n11554), .ZN(n11556) );
  OAI21_X1 U14091 ( .B1(n11557), .B2(n14674), .A(n11556), .ZN(P1_U3236) );
  NAND2_X1 U14092 ( .A1(n11559), .A2(n11558), .ZN(n14030) );
  XNOR2_X1 U14093 ( .A(n14039), .B(P1_REG2_REG_17__SCAN_IN), .ZN(n14032) );
  XNOR2_X1 U14094 ( .A(n14030), .B(n14032), .ZN(n11567) );
  AOI21_X1 U14095 ( .B1(n11561), .B2(P1_REG1_REG_16__SCAN_IN), .A(n11560), 
        .ZN(n11563) );
  XNOR2_X1 U14096 ( .A(n14039), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n11562) );
  NOR2_X1 U14097 ( .A1(n11562), .A2(n11563), .ZN(n14038) );
  AOI211_X1 U14098 ( .C1(n11563), .C2(n11562), .A(n14038), .B(n14040), .ZN(
        n11566) );
  NAND2_X1 U14099 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n13843)
         );
  NAND2_X1 U14100 ( .A1(n14719), .A2(P1_ADDR_REG_17__SCAN_IN), .ZN(n11564) );
  OAI211_X1 U14101 ( .C1(n14744), .C2(n14031), .A(n13843), .B(n11564), .ZN(
        n11565) );
  AOI211_X1 U14102 ( .C1(n11567), .C2(n14059), .A(n11566), .B(n11565), .ZN(
        n11568) );
  INV_X1 U14103 ( .A(n11568), .ZN(P1_U3260) );
  XNOR2_X1 U14104 ( .A(n12105), .B(n13361), .ZN(n12268) );
  XNOR2_X1 U14105 ( .A(n6660), .B(n12268), .ZN(n11569) );
  AOI222_X1 U14106 ( .A1(n13618), .A2(n11569), .B1(n13360), .B2(n13496), .C1(
        n13362), .C2(n13462), .ZN(n14651) );
  XOR2_X1 U14107 ( .A(n12268), .B(n11570), .Z(n14654) );
  OAI211_X1 U14108 ( .C1(n14650), .C2(n11571), .A(n13603), .B(n11692), .ZN(
        n14649) );
  OAI22_X1 U14109 ( .A1(n13602), .A2(n11572), .B1(n11668), .B2(n13535), .ZN(
        n11573) );
  AOI21_X1 U14110 ( .B1(n12105), .B2(n14935), .A(n11573), .ZN(n11574) );
  OAI21_X1 U14111 ( .B1(n14649), .B2(n14939), .A(n11574), .ZN(n11575) );
  AOI21_X1 U14112 ( .B1(n14654), .B2(n13579), .A(n11575), .ZN(n11576) );
  OAI21_X1 U14113 ( .B1(n14651), .B2(n14947), .A(n11576), .ZN(P2_U3251) );
  INV_X1 U14114 ( .A(n11577), .ZN(n11578) );
  NOR2_X1 U14115 ( .A1(n11579), .A2(n11578), .ZN(n11582) );
  XNOR2_X1 U14116 ( .A(n11580), .B(n11720), .ZN(n11581) );
  XNOR2_X1 U14117 ( .A(n11582), .B(n11581), .ZN(n11589) );
  INV_X1 U14118 ( .A(n11583), .ZN(n11625) );
  NOR2_X1 U14119 ( .A1(n11624), .A2(n12726), .ZN(n11584) );
  AOI211_X1 U14120 ( .C1(n12728), .C2(n12736), .A(n11585), .B(n11584), .ZN(
        n11586) );
  OAI21_X1 U14121 ( .B1(n11625), .B2(n12700), .A(n11586), .ZN(n11587) );
  AOI21_X1 U14122 ( .B1(n14633), .B2(n12702), .A(n11587), .ZN(n11588) );
  OAI21_X1 U14123 ( .B1(n11589), .B2(n12704), .A(n11588), .ZN(P3_U3164) );
  NAND2_X1 U14124 ( .A1(n11591), .A2(n11590), .ZN(n11592) );
  AND2_X2 U14125 ( .A1(n11593), .A2(n11592), .ZN(n11601) );
  NAND2_X1 U14126 ( .A1(n11599), .A2(n11980), .ZN(n11595) );
  NAND2_X1 U14127 ( .A1(n13930), .A2(n11975), .ZN(n11594) );
  NAND2_X1 U14128 ( .A1(n11595), .A2(n11594), .ZN(n11596) );
  XNOR2_X1 U14129 ( .A(n11596), .B(n11149), .ZN(n11729) );
  NOR2_X1 U14130 ( .A1(n11938), .A2(n11597), .ZN(n11598) );
  AOI21_X1 U14131 ( .B1(n11599), .B2(n11975), .A(n11598), .ZN(n11727) );
  XNOR2_X1 U14132 ( .A(n11729), .B(n11727), .ZN(n11600) );
  NAND2_X1 U14133 ( .A1(n11601), .A2(n11600), .ZN(n11731) );
  OAI211_X1 U14134 ( .C1(n11601), .C2(n11600), .A(n11731), .B(n13880), .ZN(
        n11607) );
  NOR2_X1 U14135 ( .A1(n14684), .A2(n11602), .ZN(n11605) );
  OAI22_X1 U14136 ( .A1(n14668), .A2(n11603), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7870), .ZN(n11604) );
  AOI211_X1 U14137 ( .C1(n14665), .C2(n13929), .A(n11605), .B(n11604), .ZN(
        n11606) );
  OAI211_X1 U14138 ( .C1(n11608), .C2(n13875), .A(n11607), .B(n11606), .ZN(
        P1_U3224) );
  AOI211_X1 U14139 ( .C1(n11611), .C2(n14983), .A(n11610), .B(n11609), .ZN(
        n11618) );
  MUX2_X1 U14140 ( .A(n11096), .B(n11618), .S(n15019), .Z(n11612) );
  OAI21_X1 U14141 ( .B1(n9580), .B2(n13724), .A(n11612), .ZN(P2_U3512) );
  INV_X1 U14142 ( .A(n11613), .ZN(n11616) );
  OAI222_X1 U14143 ( .A1(n13780), .A2(n11615), .B1(n6551), .B2(n11616), .C1(
        n11614), .C2(P2_U3088), .ZN(P2_U3303) );
  OAI222_X1 U14144 ( .A1(n14433), .A2(n11617), .B1(n12610), .B2(n11616), .C1(
        n8218), .C2(P1_U3086), .ZN(P1_U3331) );
  MUX2_X1 U14145 ( .A(n9329), .B(n11618), .S(n15007), .Z(n11619) );
  OAI21_X1 U14146 ( .B1(n9580), .B2(n13764), .A(n11619), .ZN(P2_U3469) );
  XNOR2_X1 U14147 ( .A(n11620), .B(n6996), .ZN(n14630) );
  XNOR2_X1 U14148 ( .A(n11622), .B(n11621), .ZN(n11623) );
  OAI222_X1 U14149 ( .A1(n13069), .A2(n11789), .B1(n13067), .B2(n11624), .C1(
        n13064), .C2(n11623), .ZN(n14631) );
  NAND2_X1 U14150 ( .A1(n14631), .A2(n15132), .ZN(n11628) );
  OAI22_X1 U14151 ( .A1(n15132), .A2(n12746), .B1(n11625), .B2(n15118), .ZN(
        n11626) );
  AOI21_X1 U14152 ( .B1(n14617), .B2(n14633), .A(n11626), .ZN(n11627) );
  OAI211_X1 U14153 ( .C1(n11795), .C2(n14630), .A(n11628), .B(n11627), .ZN(
        P3_U3221) );
  NAND2_X1 U14154 ( .A1(n11629), .A2(n11633), .ZN(n11630) );
  AND2_X1 U14155 ( .A1(n11631), .A2(n11630), .ZN(n11772) );
  INV_X1 U14156 ( .A(n11772), .ZN(n11640) );
  XNOR2_X1 U14157 ( .A(n11632), .B(n11633), .ZN(n11634) );
  OAI222_X1 U14158 ( .A1(n14770), .A2(n14666), .B1(n14276), .B2(n14669), .C1(
        n14761), .C2(n11634), .ZN(n11770) );
  NAND2_X1 U14159 ( .A1(n11770), .A2(n14256), .ZN(n11639) );
  AOI211_X1 U14160 ( .C1(n14680), .C2(n11635), .A(n14793), .B(n7011), .ZN(
        n11771) );
  INV_X1 U14161 ( .A(n14680), .ZN(n11778) );
  NOR2_X1 U14162 ( .A1(n11778), .A2(n14271), .ZN(n11637) );
  OAI22_X1 U14163 ( .A1(n14256), .A2(n11326), .B1(n14683), .B2(n14777), .ZN(
        n11636) );
  AOI211_X1 U14164 ( .C1(n11771), .C2(n14284), .A(n11637), .B(n11636), .ZN(
        n11638) );
  OAI211_X1 U14165 ( .C1(n11640), .C2(n14286), .A(n11639), .B(n11638), .ZN(
        P1_U3279) );
  AOI21_X1 U14166 ( .B1(n11642), .B2(n11641), .A(n6668), .ZN(n11648) );
  INV_X1 U14167 ( .A(n11643), .ZN(n11793) );
  INV_X1 U14168 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n15388) );
  NOR2_X1 U14169 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15388), .ZN(n12779) );
  NOR2_X1 U14170 ( .A1(n11789), .A2(n12726), .ZN(n11644) );
  AOI211_X1 U14171 ( .C1(n12728), .C2(n12735), .A(n12779), .B(n11644), .ZN(
        n11645) );
  OAI21_X1 U14172 ( .B1(n11793), .B2(n12700), .A(n11645), .ZN(n11646) );
  AOI21_X1 U14173 ( .B1(n13140), .B2(n12702), .A(n11646), .ZN(n11647) );
  OAI21_X1 U14174 ( .B1(n11648), .B2(n12704), .A(n11647), .ZN(P3_U3155) );
  INV_X1 U14175 ( .A(n11649), .ZN(n11653) );
  OAI222_X1 U14176 ( .A1(n13768), .A2(n11651), .B1(n6551), .B2(n11653), .C1(
        n11650), .C2(P2_U3088), .ZN(P2_U3302) );
  OAI222_X1 U14177 ( .A1(n14433), .A2(n8965), .B1(n12610), .B2(n11653), .C1(
        n11652), .C2(P1_U3086), .ZN(P1_U3330) );
  XNOR2_X1 U14178 ( .A(n12105), .B(n13236), .ZN(n11654) );
  NAND2_X1 U14179 ( .A1(n10574), .A2(n13361), .ZN(n11655) );
  NAND2_X1 U14180 ( .A1(n11654), .A2(n11655), .ZN(n11827) );
  INV_X1 U14181 ( .A(n11654), .ZN(n11657) );
  INV_X1 U14182 ( .A(n11655), .ZN(n11656) );
  NAND2_X1 U14183 ( .A1(n11657), .A2(n11656), .ZN(n11658) );
  AND2_X1 U14184 ( .A1(n11827), .A2(n11658), .ZN(n11666) );
  INV_X1 U14185 ( .A(n11661), .ZN(n11664) );
  INV_X1 U14186 ( .A(n11662), .ZN(n11663) );
  OAI21_X1 U14187 ( .B1(n11666), .B2(n11665), .A(n11698), .ZN(n11667) );
  NAND2_X1 U14188 ( .A1(n11667), .A2(n13326), .ZN(n11673) );
  OAI22_X1 U14189 ( .A1(n13329), .A2(n12112), .B1(n13344), .B2(n11668), .ZN(
        n11669) );
  AOI211_X1 U14190 ( .C1(n11671), .C2(n13362), .A(n11670), .B(n11669), .ZN(
        n11672) );
  OAI211_X1 U14191 ( .C1(n14650), .C2(n13334), .A(n11673), .B(n11672), .ZN(
        P2_U3187) );
  XNOR2_X1 U14192 ( .A(n11674), .B(n11675), .ZN(n14379) );
  INV_X1 U14193 ( .A(n14237), .ZN(n14218) );
  XNOR2_X1 U14194 ( .A(n11676), .B(n11675), .ZN(n14377) );
  INV_X1 U14195 ( .A(n13909), .ZN(n11682) );
  NAND2_X1 U14196 ( .A1(n14247), .A2(n13926), .ZN(n11678) );
  NAND2_X1 U14197 ( .A1(n14757), .A2(n13928), .ZN(n11677) );
  NAND2_X1 U14198 ( .A1(n11678), .A2(n11677), .ZN(n14371) );
  NAND2_X1 U14199 ( .A1(n14373), .A2(n11679), .ZN(n11680) );
  NAND2_X1 U14200 ( .A1(n11755), .A2(n11680), .ZN(n14375) );
  NOR2_X1 U14201 ( .A1(n14375), .A2(n10823), .ZN(n11681) );
  AOI211_X1 U14202 ( .C1(n14786), .C2(n11682), .A(n14371), .B(n11681), .ZN(
        n11684) );
  AOI22_X1 U14203 ( .A1(n14373), .A2(n14258), .B1(n14281), .B2(
        P1_REG2_REG_15__SCAN_IN), .ZN(n11683) );
  OAI21_X1 U14204 ( .B1(n11684), .B2(n14281), .A(n11683), .ZN(n11685) );
  AOI21_X1 U14205 ( .B1(n14218), .B2(n14377), .A(n11685), .ZN(n11686) );
  OAI21_X1 U14206 ( .B1(n14286), .B2(n14379), .A(n11686), .ZN(P1_U3278) );
  XNOR2_X1 U14207 ( .A(n11688), .B(n11687), .ZN(n11689) );
  AOI22_X1 U14208 ( .A1(n13462), .A2(n13361), .B1(n13496), .B2(n13359), .ZN(
        n11702) );
  OAI21_X1 U14209 ( .B1(n11689), .B2(n13600), .A(n11702), .ZN(n11763) );
  INV_X1 U14210 ( .A(n11763), .ZN(n11697) );
  XNOR2_X1 U14211 ( .A(n11690), .B(n12270), .ZN(n11765) );
  INV_X1 U14212 ( .A(n11810), .ZN(n11691) );
  AOI211_X1 U14213 ( .C1(n12110), .C2(n11692), .A(n10574), .B(n11691), .ZN(
        n11764) );
  NAND2_X1 U14214 ( .A1(n11764), .A2(n13613), .ZN(n11694) );
  AOI22_X1 U14215 ( .A1(n14947), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n14936), 
        .B2(n11705), .ZN(n11693) );
  OAI211_X1 U14216 ( .C1(n6968), .C2(n13610), .A(n11694), .B(n11693), .ZN(
        n11695) );
  AOI21_X1 U14217 ( .B1(n13579), .B2(n11765), .A(n11695), .ZN(n11696) );
  OAI21_X1 U14218 ( .B1(n11697), .B2(n14947), .A(n11696), .ZN(P2_U3250) );
  NAND2_X1 U14219 ( .A1(n11698), .A2(n11827), .ZN(n11700) );
  XNOR2_X1 U14220 ( .A(n12110), .B(n13236), .ZN(n11831) );
  NAND2_X1 U14221 ( .A1(n10574), .A2(n13360), .ZN(n11832) );
  XNOR2_X1 U14222 ( .A(n11831), .B(n11832), .ZN(n11699) );
  XNOR2_X1 U14223 ( .A(n11700), .B(n11699), .ZN(n11707) );
  OAI22_X1 U14224 ( .A1(n13318), .A2(n11702), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11701), .ZN(n11704) );
  NOR2_X1 U14225 ( .A1(n6968), .A2(n13334), .ZN(n11703) );
  AOI211_X1 U14226 ( .C1(n13320), .C2(n11705), .A(n11704), .B(n11703), .ZN(
        n11706) );
  OAI21_X1 U14227 ( .B1(n11707), .B2(n13348), .A(n11706), .ZN(P2_U3213) );
  XNOR2_X1 U14228 ( .A(n11708), .B(n13054), .ZN(n11709) );
  XNOR2_X1 U14229 ( .A(n11710), .B(n11709), .ZN(n11716) );
  NAND2_X1 U14230 ( .A1(n12728), .A2(n12734), .ZN(n11711) );
  NAND2_X1 U14231 ( .A1(P3_U3151), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n12810)
         );
  OAI211_X1 U14232 ( .C1(n13066), .C2(n12726), .A(n11711), .B(n12810), .ZN(
        n11714) );
  INV_X1 U14233 ( .A(n11712), .ZN(n13189) );
  NOR2_X1 U14234 ( .A1(n13189), .A2(n12731), .ZN(n11713) );
  AOI211_X1 U14235 ( .C1(n13073), .C2(n12724), .A(n11714), .B(n11713), .ZN(
        n11715) );
  OAI21_X1 U14236 ( .B1(n11716), .B2(n12704), .A(n11715), .ZN(P3_U3181) );
  XNOR2_X1 U14237 ( .A(n11717), .B(n12488), .ZN(n14626) );
  XOR2_X1 U14238 ( .A(n12488), .B(n11718), .Z(n11719) );
  OAI222_X1 U14239 ( .A1(n13069), .A2(n13066), .B1(n13067), .B2(n11720), .C1(
        n13064), .C2(n11719), .ZN(n14628) );
  NAND2_X1 U14240 ( .A1(n14628), .A2(n15132), .ZN(n11726) );
  OAI22_X1 U14241 ( .A1(n15132), .A2(n11722), .B1(n11721), .B2(n15118), .ZN(
        n11723) );
  AOI21_X1 U14242 ( .B1(n11724), .B2(n14617), .A(n11723), .ZN(n11725) );
  OAI211_X1 U14243 ( .C1(n11795), .C2(n14626), .A(n11726), .B(n11725), .ZN(
        P3_U3220) );
  INV_X1 U14244 ( .A(n11727), .ZN(n11728) );
  NAND2_X1 U14245 ( .A1(n11729), .A2(n11728), .ZN(n11730) );
  NAND2_X1 U14246 ( .A1(n11731), .A2(n11730), .ZN(n11738) );
  NAND2_X1 U14247 ( .A1(n11736), .A2(n11980), .ZN(n11733) );
  NAND2_X1 U14248 ( .A1(n13929), .A2(n11975), .ZN(n11732) );
  NAND2_X1 U14249 ( .A1(n11733), .A2(n11732), .ZN(n11734) );
  XNOR2_X1 U14250 ( .A(n11734), .B(n11149), .ZN(n11887) );
  NOR2_X1 U14251 ( .A1(n11938), .A2(n14669), .ZN(n11735) );
  AOI21_X1 U14252 ( .B1(n11736), .B2(n11975), .A(n11735), .ZN(n11885) );
  XNOR2_X1 U14253 ( .A(n11887), .B(n11885), .ZN(n11737) );
  NAND2_X1 U14254 ( .A1(n11738), .A2(n11737), .ZN(n14671) );
  OAI211_X1 U14255 ( .C1(n11738), .C2(n11737), .A(n14671), .B(n13880), .ZN(
        n11744) );
  INV_X1 U14256 ( .A(n11739), .ZN(n11742) );
  OAI21_X1 U14257 ( .B1(n13870), .B2(n14380), .A(n11740), .ZN(n11741) );
  AOI21_X1 U14258 ( .B1(n11742), .B2(n13891), .A(n11741), .ZN(n11743) );
  OAI211_X1 U14259 ( .C1(n14382), .C2(n13875), .A(n11744), .B(n11743), .ZN(
        P1_U3234) );
  INV_X1 U14260 ( .A(SI_24_), .ZN(n11747) );
  INV_X1 U14261 ( .A(n11745), .ZN(n11746) );
  OAI222_X1 U14262 ( .A1(P3_U3151), .A2(n11748), .B1(n13217), .B2(n11747), 
        .C1(n13213), .C2(n11746), .ZN(P3_U3271) );
  INV_X1 U14263 ( .A(n11749), .ZN(n11750) );
  AOI21_X1 U14264 ( .B1(n11753), .B2(n11751), .A(n11750), .ZN(n14370) );
  AOI22_X1 U14265 ( .A1(n11898), .A2(n14258), .B1(P1_REG2_REG_16__SCAN_IN), 
        .B2(n14281), .ZN(n11762) );
  OAI21_X1 U14266 ( .B1(n11754), .B2(n11753), .A(n11752), .ZN(n14367) );
  INV_X1 U14267 ( .A(n11898), .ZN(n14362) );
  XNOR2_X1 U14268 ( .A(n11755), .B(n14362), .ZN(n14366) );
  INV_X1 U14269 ( .A(n14366), .ZN(n11759) );
  NAND2_X1 U14270 ( .A1(n13925), .A2(n14247), .ZN(n11757) );
  NAND2_X1 U14271 ( .A1(n14757), .A2(n13927), .ZN(n11756) );
  NAND2_X1 U14272 ( .A1(n11757), .A2(n11756), .ZN(n14363) );
  AOI21_X1 U14273 ( .B1(n13836), .B2(n14786), .A(n14363), .ZN(n11758) );
  OAI21_X1 U14274 ( .B1(n11759), .B2(n10823), .A(n11758), .ZN(n11760) );
  AOI22_X1 U14275 ( .A1(n14367), .A2(n14235), .B1(n14256), .B2(n11760), .ZN(
        n11761) );
  OAI211_X1 U14276 ( .C1(n14370), .C2(n14237), .A(n11762), .B(n11761), .ZN(
        P1_U3277) );
  AOI211_X1 U14277 ( .C1(n14983), .C2(n11765), .A(n11764), .B(n11763), .ZN(
        n11767) );
  MUX2_X1 U14278 ( .A(n14884), .B(n11767), .S(n15019), .Z(n11766) );
  OAI21_X1 U14279 ( .B1(n6968), .B2(n13724), .A(n11766), .ZN(P2_U3514) );
  MUX2_X1 U14280 ( .A(n11768), .B(n11767), .S(n15007), .Z(n11769) );
  OAI21_X1 U14281 ( .B1(n6968), .B2(n13764), .A(n11769), .ZN(P2_U3475) );
  AOI211_X1 U14282 ( .C1(n14803), .C2(n11772), .A(n11771), .B(n11770), .ZN(
        n11775) );
  MUX2_X1 U14283 ( .A(n11773), .B(n11775), .S(n14811), .Z(n11774) );
  OAI21_X1 U14284 ( .B1(n11778), .B2(n14327), .A(n11774), .ZN(P1_U3542) );
  MUX2_X1 U14285 ( .A(n11776), .B(n11775), .S(n14806), .Z(n11777) );
  OAI21_X1 U14286 ( .B1(n11778), .B2(n14411), .A(n11777), .ZN(P1_U3501) );
  XNOR2_X1 U14287 ( .A(n11779), .B(n13068), .ZN(n11780) );
  XNOR2_X1 U14288 ( .A(n11781), .B(n11780), .ZN(n11787) );
  NAND2_X1 U14289 ( .A1(n12728), .A2(n11782), .ZN(n11783) );
  NAND2_X1 U14290 ( .A1(P3_U3151), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n12821)
         );
  OAI211_X1 U14291 ( .C1(n13054), .C2(n12726), .A(n11783), .B(n12821), .ZN(
        n11785) );
  NOR2_X1 U14292 ( .A1(n13184), .A2(n12731), .ZN(n11784) );
  AOI211_X1 U14293 ( .C1(n13058), .C2(n12724), .A(n11785), .B(n11784), .ZN(
        n11786) );
  OAI21_X1 U14294 ( .B1(n11787), .B2(n12704), .A(n11786), .ZN(P3_U3166) );
  AOI21_X1 U14295 ( .B1(n11788), .B2(n9050), .A(n13064), .ZN(n11792) );
  OAI22_X1 U14296 ( .A1(n11789), .A2(n13067), .B1(n13054), .B2(n13069), .ZN(
        n11790) );
  AOI21_X1 U14297 ( .B1(n11792), .B2(n11791), .A(n11790), .ZN(n13142) );
  OAI22_X1 U14298 ( .A1(n15132), .A2(n12769), .B1(n11793), .B2(n15118), .ZN(
        n11797) );
  XNOR2_X1 U14299 ( .A(n11794), .B(n9050), .ZN(n13143) );
  NOR2_X1 U14300 ( .A1(n13143), .A2(n11795), .ZN(n11796) );
  AOI211_X1 U14301 ( .C1(n14617), .C2(n13140), .A(n11797), .B(n11796), .ZN(
        n11798) );
  OAI21_X1 U14302 ( .B1(n13074), .B2(n13142), .A(n11798), .ZN(P3_U3219) );
  INV_X1 U14303 ( .A(n11799), .ZN(n11800) );
  OAI222_X1 U14304 ( .A1(P3_U3151), .A2(n11802), .B1(n13217), .B2(n11801), 
        .C1(n13213), .C2(n11800), .ZN(P3_U3270) );
  OAI21_X1 U14305 ( .B1(n6654), .B2(n12266), .A(n11803), .ZN(n13729) );
  OAI211_X1 U14306 ( .C1(n11806), .C2(n11805), .A(n11804), .B(n13618), .ZN(
        n11808) );
  AOI22_X1 U14307 ( .A1(n13496), .A2(n13358), .B1(n13462), .B2(n13360), .ZN(
        n11807) );
  AND2_X1 U14308 ( .A1(n11808), .A2(n11807), .ZN(n13728) );
  OAI21_X1 U14309 ( .B1(n11840), .B2(n13535), .A(n13728), .ZN(n11809) );
  NAND2_X1 U14310 ( .A1(n11809), .A2(n13602), .ZN(n11815) );
  AOI211_X1 U14311 ( .C1(n13726), .C2(n11810), .A(n10574), .B(n11848), .ZN(
        n13725) );
  INV_X1 U14312 ( .A(n13726), .ZN(n11812) );
  INV_X1 U14313 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n11811) );
  OAI22_X1 U14314 ( .A1(n11812), .A2(n13610), .B1(n13602), .B2(n11811), .ZN(
        n11813) );
  AOI21_X1 U14315 ( .B1(n13725), .B2(n13613), .A(n11813), .ZN(n11814) );
  OAI211_X1 U14316 ( .C1(n13729), .C2(n14942), .A(n11815), .B(n11814), .ZN(
        P2_U3249) );
  INV_X1 U14317 ( .A(n11816), .ZN(n11819) );
  OAI222_X1 U14318 ( .A1(n11818), .A2(P2_U3088), .B1(n6551), .B2(n11819), .C1(
        n11817), .C2(n13780), .ZN(P2_U3301) );
  OAI222_X1 U14319 ( .A1(n14433), .A2(n11821), .B1(P1_U3086), .B2(n11820), 
        .C1(n12610), .C2(n11819), .ZN(P1_U3329) );
  XNOR2_X1 U14320 ( .A(n13726), .B(n13236), .ZN(n11822) );
  NAND2_X1 U14321 ( .A1(n10574), .A2(n13359), .ZN(n11823) );
  NAND2_X1 U14322 ( .A1(n11822), .A2(n11823), .ZN(n11861) );
  INV_X1 U14323 ( .A(n11822), .ZN(n11825) );
  INV_X1 U14324 ( .A(n11823), .ZN(n11824) );
  NAND2_X1 U14325 ( .A1(n11825), .A2(n11824), .ZN(n11826) );
  NAND2_X1 U14326 ( .A1(n11861), .A2(n11826), .ZN(n11839) );
  INV_X1 U14327 ( .A(n11827), .ZN(n11828) );
  AOI21_X1 U14328 ( .B1(n11831), .B2(n11832), .A(n11828), .ZN(n11829) );
  INV_X1 U14329 ( .A(n11831), .ZN(n11834) );
  INV_X1 U14330 ( .A(n11832), .ZN(n11833) );
  NAND2_X1 U14331 ( .A1(n11834), .A2(n11833), .ZN(n11835) );
  OR2_X2 U14332 ( .A1(n11838), .A2(n11839), .ZN(n11862) );
  INV_X1 U14333 ( .A(n11862), .ZN(n11837) );
  AOI21_X1 U14334 ( .B1(n11839), .B2(n11838), .A(n11837), .ZN(n11844) );
  NAND2_X1 U14335 ( .A1(P2_U3088), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n14901)
         );
  OAI21_X1 U14336 ( .B1(n13328), .B2(n12112), .A(n14901), .ZN(n11842) );
  OAI22_X1 U14337 ( .A1(n13329), .A2(n13628), .B1(n13344), .B2(n11840), .ZN(
        n11841) );
  AOI211_X1 U14338 ( .C1(n13726), .C2(n13346), .A(n11842), .B(n11841), .ZN(
        n11843) );
  OAI21_X1 U14339 ( .B1(n11844), .B2(n13348), .A(n11843), .ZN(P2_U3198) );
  XNOR2_X1 U14340 ( .A(n11845), .B(n12267), .ZN(n13721) );
  INV_X1 U14341 ( .A(n13721), .ZN(n11855) );
  XNOR2_X1 U14342 ( .A(n11846), .B(n12267), .ZN(n11847) );
  AOI22_X1 U14343 ( .A1(n13357), .A2(n13496), .B1(n13462), .B2(n13359), .ZN(
        n11867) );
  OAI21_X1 U14344 ( .B1(n11847), .B2(n13600), .A(n11867), .ZN(n13719) );
  NAND2_X1 U14345 ( .A1(n13719), .A2(n13602), .ZN(n11854) );
  INV_X1 U14346 ( .A(n11848), .ZN(n11850) );
  INV_X1 U14347 ( .A(n13632), .ZN(n11849) );
  AOI211_X1 U14348 ( .C1(n12125), .C2(n11850), .A(n10574), .B(n11849), .ZN(
        n13720) );
  NOR2_X1 U14349 ( .A1(n13765), .A2(n13610), .ZN(n11852) );
  INV_X1 U14350 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n13390) );
  OAI22_X1 U14351 ( .A1(n13602), .A2(n13390), .B1(n11866), .B2(n13535), .ZN(
        n11851) );
  AOI211_X1 U14352 ( .C1(n13720), .C2(n13613), .A(n11852), .B(n11851), .ZN(
        n11853) );
  OAI211_X1 U14353 ( .C1(n11855), .C2(n14942), .A(n11854), .B(n11853), .ZN(
        P2_U3248) );
  XNOR2_X1 U14354 ( .A(n12125), .B(n13236), .ZN(n11856) );
  NAND2_X1 U14355 ( .A1(n13358), .A2(n10574), .ZN(n11857) );
  NAND2_X1 U14356 ( .A1(n11856), .A2(n11857), .ZN(n11874) );
  INV_X1 U14357 ( .A(n11856), .ZN(n11859) );
  INV_X1 U14358 ( .A(n11857), .ZN(n11858) );
  NAND2_X1 U14359 ( .A1(n11859), .A2(n11858), .ZN(n11860) );
  AND2_X1 U14360 ( .A1(n11874), .A2(n11860), .ZN(n11864) );
  OAI21_X1 U14361 ( .B1(n11864), .B2(n11863), .A(n11875), .ZN(n11865) );
  NAND2_X1 U14362 ( .A1(n11865), .A2(n13326), .ZN(n11871) );
  INV_X1 U14363 ( .A(n11866), .ZN(n11869) );
  NAND2_X1 U14364 ( .A1(P2_U3088), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n14915)
         );
  OAI21_X1 U14365 ( .B1(n13318), .B2(n11867), .A(n14915), .ZN(n11868) );
  AOI21_X1 U14366 ( .B1(n11869), .B2(n13320), .A(n11868), .ZN(n11870) );
  OAI211_X1 U14367 ( .C1(n13765), .C2(n13334), .A(n11871), .B(n11870), .ZN(
        P2_U3200) );
  INV_X1 U14368 ( .A(n11872), .ZN(n12311) );
  OAI222_X1 U14369 ( .A1(n14433), .A2(n11873), .B1(P1_U3086), .B2(n13962), 
        .C1(n12610), .C2(n12311), .ZN(P1_U3328) );
  XNOR2_X1 U14370 ( .A(n13711), .B(n13236), .ZN(n13221) );
  NAND2_X1 U14371 ( .A1(n13357), .A2(n10574), .ZN(n13220) );
  XNOR2_X1 U14372 ( .A(n13221), .B(n13220), .ZN(n13222) );
  XNOR2_X1 U14373 ( .A(n13223), .B(n13222), .ZN(n11880) );
  AOI22_X1 U14374 ( .A1(n11876), .A2(n13625), .B1(n13320), .B2(n13634), .ZN(
        n11877) );
  NAND2_X1 U14375 ( .A1(P2_U3088), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n14930)
         );
  OAI211_X1 U14376 ( .C1(n13628), .C2(n13328), .A(n11877), .B(n14930), .ZN(
        n11878) );
  AOI21_X1 U14377 ( .B1(n13711), .B2(n13346), .A(n11878), .ZN(n11879) );
  OAI21_X1 U14378 ( .B1(n11880), .B2(n13348), .A(n11879), .ZN(P2_U3210) );
  NAND2_X1 U14379 ( .A1(n14680), .A2(n11980), .ZN(n11882) );
  NAND2_X1 U14380 ( .A1(n13928), .A2(n11975), .ZN(n11881) );
  NAND2_X1 U14381 ( .A1(n11882), .A2(n11881), .ZN(n11883) );
  XNOR2_X1 U14382 ( .A(n11883), .B(n8150), .ZN(n11891) );
  NOR2_X1 U14383 ( .A1(n11938), .A2(n13906), .ZN(n11884) );
  AOI21_X1 U14384 ( .B1(n14680), .B2(n11975), .A(n11884), .ZN(n11890) );
  XNOR2_X1 U14385 ( .A(n11891), .B(n11890), .ZN(n14672) );
  INV_X1 U14386 ( .A(n14672), .ZN(n11888) );
  INV_X1 U14387 ( .A(n11885), .ZN(n11886) );
  NAND2_X1 U14388 ( .A1(n11887), .A2(n11886), .ZN(n14670) );
  AND2_X1 U14389 ( .A1(n11888), .A2(n14670), .ZN(n11889) );
  NAND2_X1 U14390 ( .A1(n14671), .A2(n11889), .ZN(n14676) );
  NAND2_X1 U14391 ( .A1(n11891), .A2(n11890), .ZN(n11892) );
  NAND2_X1 U14392 ( .A1(n14676), .A2(n11892), .ZN(n11894) );
  AOI22_X1 U14393 ( .A1(n14373), .A2(n11980), .B1(n11975), .B2(n13927), .ZN(
        n11893) );
  XNOR2_X1 U14394 ( .A(n11893), .B(n11149), .ZN(n11895) );
  AOI22_X1 U14395 ( .A1(n14373), .A2(n11975), .B1(n11979), .B2(n13927), .ZN(
        n13912) );
  INV_X1 U14396 ( .A(n11894), .ZN(n11897) );
  INV_X1 U14397 ( .A(n11895), .ZN(n11896) );
  AOI22_X1 U14398 ( .A1(n11898), .A2(n11975), .B1(n11979), .B2(n13926), .ZN(
        n11901) );
  AOI22_X1 U14399 ( .A1(n11898), .A2(n11980), .B1(n11975), .B2(n13926), .ZN(
        n11899) );
  XNOR2_X1 U14400 ( .A(n11899), .B(n11149), .ZN(n11900) );
  XOR2_X1 U14401 ( .A(n11901), .B(n11900), .Z(n13831) );
  NAND2_X1 U14402 ( .A1(n13830), .A2(n11902), .ZN(n13840) );
  NAND2_X1 U14403 ( .A1(n14358), .A2(n11980), .ZN(n11904) );
  NAND2_X1 U14404 ( .A1(n13925), .A2(n11975), .ZN(n11903) );
  NAND2_X1 U14405 ( .A1(n11904), .A2(n11903), .ZN(n11905) );
  XNOR2_X1 U14406 ( .A(n11905), .B(n11149), .ZN(n11908) );
  AOI22_X1 U14407 ( .A1(n14358), .A2(n11975), .B1(n11979), .B2(n13925), .ZN(
        n11906) );
  XNOR2_X1 U14408 ( .A(n11908), .B(n11906), .ZN(n13841) );
  INV_X1 U14409 ( .A(n11906), .ZN(n11907) );
  NAND2_X1 U14410 ( .A1(n14350), .A2(n11980), .ZN(n11911) );
  NAND2_X1 U14411 ( .A1(n13924), .A2(n11975), .ZN(n11910) );
  NAND2_X1 U14412 ( .A1(n11911), .A2(n11910), .ZN(n11912) );
  XNOR2_X1 U14413 ( .A(n11912), .B(n11149), .ZN(n11913) );
  AOI22_X1 U14414 ( .A1(n14350), .A2(n10626), .B1(n11979), .B2(n13924), .ZN(
        n11914) );
  XNOR2_X1 U14415 ( .A(n11913), .B(n11914), .ZN(n13890) );
  INV_X1 U14416 ( .A(n11913), .ZN(n11915) );
  NAND2_X1 U14417 ( .A1(n14345), .A2(n6547), .ZN(n11917) );
  NAND2_X1 U14418 ( .A1(n14248), .A2(n11975), .ZN(n11916) );
  NAND2_X1 U14419 ( .A1(n11917), .A2(n11916), .ZN(n11918) );
  XNOR2_X1 U14420 ( .A(n11918), .B(n11149), .ZN(n11920) );
  AND2_X1 U14421 ( .A1(n11979), .A2(n14248), .ZN(n11919) );
  AOI21_X1 U14422 ( .B1(n14345), .B2(n11975), .A(n11919), .ZN(n11921) );
  XNOR2_X1 U14423 ( .A(n11920), .B(n11921), .ZN(n13798) );
  NAND2_X1 U14424 ( .A1(n11920), .A2(n11922), .ZN(n11923) );
  AND2_X1 U14425 ( .A1(n13923), .A2(n11979), .ZN(n11924) );
  AOI21_X1 U14426 ( .B1(n14415), .B2(n11975), .A(n11924), .ZN(n11927) );
  AOI22_X1 U14427 ( .A1(n14415), .A2(n11980), .B1(n11975), .B2(n13923), .ZN(
        n11925) );
  XNOR2_X1 U14428 ( .A(n11925), .B(n11149), .ZN(n11926) );
  XOR2_X1 U14429 ( .A(n11927), .B(n11926), .Z(n13856) );
  INV_X1 U14430 ( .A(n11926), .ZN(n11929) );
  INV_X1 U14431 ( .A(n11927), .ZN(n11928) );
  NAND2_X1 U14432 ( .A1(n11929), .A2(n11928), .ZN(n11930) );
  AOI22_X1 U14433 ( .A1(n14199), .A2(n10626), .B1(n11979), .B2(n13922), .ZN(
        n11934) );
  NAND2_X1 U14434 ( .A1(n14199), .A2(n6547), .ZN(n11932) );
  NAND2_X1 U14435 ( .A1(n13922), .A2(n11975), .ZN(n11931) );
  NAND2_X1 U14436 ( .A1(n11932), .A2(n11931), .ZN(n11933) );
  XNOR2_X1 U14437 ( .A(n11933), .B(n11149), .ZN(n11936) );
  XOR2_X1 U14438 ( .A(n11934), .B(n11936), .Z(n13815) );
  INV_X1 U14439 ( .A(n11934), .ZN(n11935) );
  OAI22_X1 U14440 ( .A1(n14410), .A2(n11939), .B1(n13817), .B2(n11938), .ZN(
        n11943) );
  OAI22_X1 U14441 ( .A1(n14410), .A2(n11940), .B1(n13817), .B2(n11939), .ZN(
        n11941) );
  XNOR2_X1 U14442 ( .A(n11941), .B(n11149), .ZN(n11942) );
  XOR2_X1 U14443 ( .A(n11943), .B(n11942), .Z(n13866) );
  NAND2_X1 U14444 ( .A1(n13865), .A2(n13866), .ZN(n13864) );
  INV_X1 U14445 ( .A(n11942), .ZN(n11945) );
  NAND2_X1 U14446 ( .A1(n14160), .A2(n11980), .ZN(n11948) );
  NAND2_X1 U14447 ( .A1(n14140), .A2(n11975), .ZN(n11947) );
  NAND2_X1 U14448 ( .A1(n11948), .A2(n11947), .ZN(n11949) );
  XNOR2_X1 U14449 ( .A(n11949), .B(n11149), .ZN(n11950) );
  AOI22_X1 U14450 ( .A1(n14160), .A2(n11975), .B1(n11979), .B2(n14140), .ZN(
        n11951) );
  XNOR2_X1 U14451 ( .A(n11950), .B(n11951), .ZN(n13790) );
  INV_X1 U14452 ( .A(n11950), .ZN(n11952) );
  AOI22_X1 U14453 ( .A1(n14148), .A2(n11975), .B1(n11979), .B2(n13920), .ZN(
        n11956) );
  NAND2_X1 U14454 ( .A1(n14148), .A2(n11980), .ZN(n11954) );
  NAND2_X1 U14455 ( .A1(n13920), .A2(n11975), .ZN(n11953) );
  NAND2_X1 U14456 ( .A1(n11954), .A2(n11953), .ZN(n11955) );
  XNOR2_X1 U14457 ( .A(n11955), .B(n11149), .ZN(n11958) );
  XOR2_X1 U14458 ( .A(n11956), .B(n11958), .Z(n13849) );
  INV_X1 U14459 ( .A(n11956), .ZN(n11957) );
  OR2_X1 U14460 ( .A1(n11958), .A2(n11957), .ZN(n11959) );
  NAND2_X1 U14461 ( .A1(n14400), .A2(n11980), .ZN(n11961) );
  NAND2_X1 U14462 ( .A1(n14139), .A2(n11975), .ZN(n11960) );
  NAND2_X1 U14463 ( .A1(n11961), .A2(n11960), .ZN(n11962) );
  XNOR2_X1 U14464 ( .A(n11962), .B(n11149), .ZN(n11963) );
  AOI22_X1 U14465 ( .A1(n14400), .A2(n11975), .B1(n11979), .B2(n14139), .ZN(
        n11964) );
  XNOR2_X1 U14466 ( .A(n11963), .B(n11964), .ZN(n13824) );
  INV_X1 U14467 ( .A(n11963), .ZN(n11965) );
  AOI22_X1 U14468 ( .A1(n14396), .A2(n11975), .B1(n11979), .B2(n13919), .ZN(
        n11969) );
  NAND2_X1 U14469 ( .A1(n14396), .A2(n11980), .ZN(n11967) );
  NAND2_X1 U14470 ( .A1(n13919), .A2(n10626), .ZN(n11966) );
  NAND2_X1 U14471 ( .A1(n11967), .A2(n11966), .ZN(n11968) );
  XNOR2_X1 U14472 ( .A(n11968), .B(n11149), .ZN(n11971) );
  XOR2_X1 U14473 ( .A(n11969), .B(n11971), .Z(n13898) );
  INV_X1 U14474 ( .A(n11969), .ZN(n11970) );
  NAND2_X1 U14475 ( .A1(n14095), .A2(n6547), .ZN(n11973) );
  NAND2_X1 U14476 ( .A1(n14106), .A2(n11975), .ZN(n11972) );
  NAND2_X1 U14477 ( .A1(n11973), .A2(n11972), .ZN(n11974) );
  XNOR2_X1 U14478 ( .A(n11974), .B(n11149), .ZN(n11976) );
  AOI22_X1 U14479 ( .A1(n14095), .A2(n11975), .B1(n11979), .B2(n14106), .ZN(
        n11977) );
  XNOR2_X1 U14480 ( .A(n11976), .B(n11977), .ZN(n13783) );
  INV_X1 U14481 ( .A(n11976), .ZN(n11978) );
  AOI22_X1 U14482 ( .A1(n14085), .A2(n11975), .B1(n11979), .B2(n13918), .ZN(
        n11983) );
  AOI22_X1 U14483 ( .A1(n14085), .A2(n11980), .B1(n10626), .B2(n13918), .ZN(
        n11981) );
  XNOR2_X1 U14484 ( .A(n11981), .B(n11149), .ZN(n11982) );
  XOR2_X1 U14485 ( .A(n11983), .B(n11982), .Z(n11984) );
  XNOR2_X1 U14486 ( .A(n11985), .B(n11984), .ZN(n11990) );
  AOI22_X1 U14487 ( .A1(n14665), .A2(n13917), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n11987) );
  NAND2_X1 U14488 ( .A1(n13900), .A2(n14106), .ZN(n11986) );
  OAI211_X1 U14489 ( .C1(n14684), .C2(n14082), .A(n11987), .B(n11986), .ZN(
        n11988) );
  AOI21_X1 U14490 ( .B1(n14085), .B2(n14679), .A(n11988), .ZN(n11989) );
  OAI21_X1 U14491 ( .B1(n11990), .B2(n14674), .A(n11989), .ZN(P1_U3220) );
  OAI22_X1 U14492 ( .A1(n14613), .A2(n12375), .B1(n15132), .B2(n11991), .ZN(
        n11992) );
  AOI21_X1 U14493 ( .B1(n14611), .B2(n15150), .A(n11992), .ZN(n11995) );
  NAND2_X1 U14494 ( .A1(n11993), .A2(n13077), .ZN(n11994) );
  OAI211_X1 U14495 ( .C1(n11996), .C2(n13074), .A(n11995), .B(n11994), .ZN(
        P3_U3204) );
  AOI22_X1 U14496 ( .A1(n13703), .A2(n12215), .B1(n12214), .B2(n13356), .ZN(
        n12145) );
  NAND2_X1 U14497 ( .A1(n13708), .A2(n12214), .ZN(n11999) );
  NAND2_X1 U14498 ( .A1(n13625), .A2(n12215), .ZN(n11998) );
  NAND2_X1 U14499 ( .A1(n11999), .A2(n11998), .ZN(n12138) );
  INV_X1 U14500 ( .A(n12138), .ZN(n12142) );
  NAND2_X1 U14501 ( .A1(n12293), .A2(n13375), .ZN(n12006) );
  AOI21_X1 U14502 ( .B1(n7536), .B2(n12000), .A(n12289), .ZN(n12001) );
  OAI21_X1 U14503 ( .B1(n12006), .B2(n12002), .A(n12001), .ZN(n12008) );
  NAND2_X1 U14504 ( .A1(n12002), .A2(n12293), .ZN(n12005) );
  NAND2_X1 U14505 ( .A1(n13375), .A2(n12003), .ZN(n12004) );
  NAND2_X1 U14506 ( .A1(n12005), .A2(n12004), .ZN(n12007) );
  NAND2_X1 U14507 ( .A1(n12293), .A2(n14934), .ZN(n12009) );
  OAI21_X1 U14508 ( .B1(n12010), .B2(n12293), .A(n12009), .ZN(n12011) );
  INV_X1 U14509 ( .A(n12153), .ZN(n12202) );
  NAND2_X1 U14510 ( .A1(n12202), .A2(n12016), .ZN(n12015) );
  NAND2_X1 U14511 ( .A1(n12153), .A2(n13373), .ZN(n12014) );
  NAND2_X1 U14512 ( .A1(n12015), .A2(n12014), .ZN(n12018) );
  AOI22_X1 U14513 ( .A1(n12202), .A2(n13373), .B1(n12153), .B2(n12016), .ZN(
        n12017) );
  NAND2_X1 U14514 ( .A1(n12202), .A2(n13372), .ZN(n12020) );
  NAND2_X1 U14515 ( .A1(n12153), .A2(n12021), .ZN(n12019) );
  NAND2_X1 U14516 ( .A1(n12020), .A2(n12019), .ZN(n12023) );
  AOI22_X1 U14517 ( .A1(n12202), .A2(n12021), .B1(n12153), .B2(n13372), .ZN(
        n12022) );
  NAND2_X1 U14518 ( .A1(n12215), .A2(n12025), .ZN(n12027) );
  NAND2_X1 U14520 ( .A1(n12203), .A2(n13371), .ZN(n12026) );
  NAND2_X1 U14521 ( .A1(n12027), .A2(n12026), .ZN(n12032) );
  NAND2_X1 U14522 ( .A1(n12215), .A2(n13371), .ZN(n12028) );
  OAI21_X1 U14523 ( .B1(n12029), .B2(n12293), .A(n12028), .ZN(n12030) );
  INV_X1 U14524 ( .A(n12032), .ZN(n12033) );
  NAND2_X1 U14525 ( .A1(n6721), .A2(n12203), .ZN(n12035) );
  NAND2_X1 U14526 ( .A1(n12215), .A2(n13370), .ZN(n12034) );
  NAND2_X1 U14527 ( .A1(n12035), .A2(n12034), .ZN(n12041) );
  NAND2_X1 U14528 ( .A1(n6721), .A2(n12215), .ZN(n12036) );
  NAND2_X1 U14529 ( .A1(n12039), .A2(n12038), .ZN(n12045) );
  INV_X1 U14530 ( .A(n12040), .ZN(n12043) );
  INV_X1 U14531 ( .A(n12041), .ZN(n12042) );
  NAND2_X1 U14532 ( .A1(n12043), .A2(n12042), .ZN(n12044) );
  NAND2_X1 U14533 ( .A1(n12048), .A2(n12215), .ZN(n12047) );
  NAND2_X1 U14534 ( .A1(n12214), .A2(n13369), .ZN(n12046) );
  AOI22_X1 U14535 ( .A1(n12048), .A2(n12203), .B1(n13369), .B2(n12215), .ZN(
        n12049) );
  NAND2_X1 U14536 ( .A1(n12052), .A2(n12214), .ZN(n12051) );
  NAND2_X1 U14537 ( .A1(n12215), .A2(n13368), .ZN(n12050) );
  NAND2_X1 U14538 ( .A1(n12051), .A2(n12050), .ZN(n12055) );
  AOI22_X1 U14539 ( .A1(n12052), .A2(n12215), .B1(n12214), .B2(n13368), .ZN(
        n12053) );
  INV_X1 U14540 ( .A(n12054), .ZN(n12057) );
  NAND2_X1 U14541 ( .A1(n12060), .A2(n12215), .ZN(n12059) );
  NAND2_X1 U14542 ( .A1(n12214), .A2(n13367), .ZN(n12058) );
  NAND2_X1 U14543 ( .A1(n12059), .A2(n12058), .ZN(n12064) );
  INV_X1 U14544 ( .A(n13367), .ZN(n12062) );
  NAND2_X1 U14545 ( .A1(n12060), .A2(n12214), .ZN(n12061) );
  OAI21_X1 U14546 ( .B1(n12062), .B2(n12214), .A(n12061), .ZN(n12063) );
  INV_X1 U14547 ( .A(n12063), .ZN(n12065) );
  NAND2_X1 U14548 ( .A1(n6703), .A2(n12214), .ZN(n12067) );
  NAND2_X1 U14549 ( .A1(n12215), .A2(n13366), .ZN(n12066) );
  NAND2_X1 U14550 ( .A1(n12067), .A2(n12066), .ZN(n12070) );
  AOI22_X1 U14551 ( .A1(n6703), .A2(n12215), .B1(n12214), .B2(n13366), .ZN(
        n12069) );
  NAND2_X1 U14552 ( .A1(n12075), .A2(n12215), .ZN(n12074) );
  NAND2_X1 U14553 ( .A1(n12214), .A2(n13365), .ZN(n12073) );
  NAND2_X1 U14554 ( .A1(n12075), .A2(n12214), .ZN(n12076) );
  OAI21_X1 U14555 ( .B1(n12077), .B2(n12214), .A(n12076), .ZN(n12078) );
  NAND2_X1 U14556 ( .A1(n12081), .A2(n12214), .ZN(n12080) );
  NAND2_X1 U14557 ( .A1(n12215), .A2(n13364), .ZN(n12079) );
  NAND2_X1 U14558 ( .A1(n12080), .A2(n12079), .ZN(n12083) );
  AOI22_X1 U14559 ( .A1(n12081), .A2(n12215), .B1(n12214), .B2(n13364), .ZN(
        n12082) );
  NAND2_X1 U14560 ( .A1(n12087), .A2(n12215), .ZN(n12086) );
  NAND2_X1 U14561 ( .A1(n12214), .A2(n13363), .ZN(n12085) );
  NAND2_X1 U14562 ( .A1(n12086), .A2(n12085), .ZN(n12089) );
  AOI22_X1 U14563 ( .A1(n12087), .A2(n12203), .B1(n13363), .B2(n12215), .ZN(
        n12088) );
  NAND2_X1 U14564 ( .A1(n12092), .A2(n12214), .ZN(n12091) );
  NAND2_X1 U14565 ( .A1(n12215), .A2(n13362), .ZN(n12090) );
  NAND2_X1 U14566 ( .A1(n12091), .A2(n12090), .ZN(n12098) );
  NAND2_X1 U14567 ( .A1(n12092), .A2(n12215), .ZN(n12093) );
  OAI21_X1 U14568 ( .B1(n12094), .B2(n12293), .A(n12093), .ZN(n12095) );
  NAND2_X1 U14569 ( .A1(n12096), .A2(n12095), .ZN(n12102) );
  INV_X1 U14570 ( .A(n12097), .ZN(n12100) );
  INV_X1 U14571 ( .A(n12098), .ZN(n12099) );
  NAND2_X1 U14572 ( .A1(n12100), .A2(n12099), .ZN(n12101) );
  NAND2_X1 U14573 ( .A1(n12105), .A2(n12215), .ZN(n12104) );
  NAND2_X1 U14574 ( .A1(n12214), .A2(n13361), .ZN(n12103) );
  NAND2_X1 U14575 ( .A1(n12104), .A2(n12103), .ZN(n12107) );
  AOI22_X1 U14576 ( .A1(n12105), .A2(n12203), .B1(n13361), .B2(n12215), .ZN(
        n12106) );
  NAND2_X1 U14577 ( .A1(n12110), .A2(n12214), .ZN(n12109) );
  NAND2_X1 U14578 ( .A1(n12215), .A2(n13360), .ZN(n12108) );
  NAND2_X1 U14579 ( .A1(n12109), .A2(n12108), .ZN(n12114) );
  NAND2_X1 U14580 ( .A1(n12110), .A2(n12215), .ZN(n12111) );
  INV_X1 U14581 ( .A(n12114), .ZN(n12115) );
  NAND2_X1 U14582 ( .A1(n13726), .A2(n12215), .ZN(n12117) );
  NAND2_X1 U14583 ( .A1(n12214), .A2(n13359), .ZN(n12116) );
  NAND2_X1 U14584 ( .A1(n12117), .A2(n12116), .ZN(n12123) );
  AOI22_X1 U14585 ( .A1(n13726), .A2(n12203), .B1(n13359), .B2(n12215), .ZN(
        n12118) );
  AOI21_X1 U14586 ( .B1(n12124), .B2(n12123), .A(n12118), .ZN(n12130) );
  AOI22_X1 U14587 ( .A1(n12125), .A2(n12215), .B1(n12214), .B2(n13358), .ZN(
        n12121) );
  NAND2_X1 U14588 ( .A1(n12125), .A2(n12214), .ZN(n12120) );
  NAND2_X1 U14589 ( .A1(n13358), .A2(n12215), .ZN(n12119) );
  NAND2_X1 U14590 ( .A1(n12120), .A2(n12119), .ZN(n12127) );
  NAND2_X1 U14591 ( .A1(n12121), .A2(n12127), .ZN(n12122) );
  OAI21_X1 U14592 ( .B1(n12124), .B2(n12123), .A(n12122), .ZN(n12129) );
  NOR2_X1 U14593 ( .A1(n12125), .A2(n13358), .ZN(n12126) );
  OR2_X1 U14594 ( .A1(n12127), .A2(n12126), .ZN(n12128) );
  OAI21_X1 U14595 ( .B1(n12130), .B2(n12129), .A(n12128), .ZN(n12136) );
  NAND2_X1 U14596 ( .A1(n13711), .A2(n12215), .ZN(n12132) );
  NAND2_X1 U14597 ( .A1(n13357), .A2(n12214), .ZN(n12131) );
  NAND2_X1 U14598 ( .A1(n13711), .A2(n12214), .ZN(n12133) );
  OAI21_X1 U14599 ( .B1(n12134), .B2(n12214), .A(n12133), .ZN(n12135) );
  AOI22_X1 U14600 ( .A1(n13708), .A2(n12215), .B1(n12214), .B2(n13625), .ZN(
        n12137) );
  AOI21_X1 U14601 ( .B1(n12139), .B2(n12138), .A(n12137), .ZN(n12140) );
  OAI22_X1 U14602 ( .A1(n13591), .A2(n12293), .B1(n12143), .B2(n12214), .ZN(
        n12144) );
  OAI22_X1 U14603 ( .A1(n13755), .A2(n12293), .B1(n13550), .B2(n12214), .ZN(
        n12147) );
  AOI22_X1 U14604 ( .A1(n13574), .A2(n12215), .B1(n12214), .B2(n13355), .ZN(
        n12146) );
  AOI22_X1 U14605 ( .A1(n13690), .A2(n12202), .B1(n12214), .B2(n13532), .ZN(
        n12148) );
  AOI22_X1 U14606 ( .A1(n13690), .A2(n12203), .B1(n13532), .B2(n12202), .ZN(
        n12151) );
  INV_X1 U14607 ( .A(n12148), .ZN(n12150) );
  OAI22_X1 U14608 ( .A1(n12152), .A2(n12151), .B1(n12150), .B2(n12149), .ZN(
        n12156) );
  OAI22_X1 U14609 ( .A1(n13542), .A2(n12293), .B1(n13549), .B2(n12153), .ZN(
        n12157) );
  AOI22_X1 U14610 ( .A1(n13686), .A2(n12202), .B1(n12214), .B2(n13354), .ZN(
        n12154) );
  AOI21_X1 U14611 ( .B1(n12156), .B2(n12157), .A(n12154), .ZN(n12155) );
  AOI22_X1 U14612 ( .A1(n13681), .A2(n12202), .B1(n12214), .B2(n13533), .ZN(
        n12159) );
  AOI22_X1 U14613 ( .A1(n13681), .A2(n12203), .B1(n13533), .B2(n12215), .ZN(
        n12158) );
  INV_X1 U14614 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n13769) );
  NAND2_X1 U14615 ( .A1(n12161), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n12164) );
  NAND2_X1 U14616 ( .A1(n12162), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n12163) );
  OAI211_X1 U14617 ( .C1(n6546), .C2(n13732), .A(n12164), .B(n12163), .ZN(
        n13420) );
  NAND2_X1 U14618 ( .A1(n12166), .A2(n13420), .ZN(n12167) );
  NAND2_X1 U14619 ( .A1(n12291), .A2(n12167), .ZN(n12283) );
  NAND2_X1 U14620 ( .A1(n13774), .A2(n12168), .ZN(n12170) );
  OR2_X1 U14621 ( .A1(n9502), .A2(n15332), .ZN(n12169) );
  AND2_X1 U14622 ( .A1(n12215), .A2(n13351), .ZN(n12171) );
  AOI21_X1 U14623 ( .B1(n13650), .B2(n12203), .A(n12171), .ZN(n12211) );
  NAND2_X1 U14624 ( .A1(n13650), .A2(n12215), .ZN(n12173) );
  NAND2_X1 U14625 ( .A1(n12214), .A2(n13351), .ZN(n12172) );
  NAND2_X1 U14626 ( .A1(n12173), .A2(n12172), .ZN(n12210) );
  NAND2_X1 U14627 ( .A1(n12211), .A2(n12210), .ZN(n12222) );
  AND2_X1 U14628 ( .A1(n12215), .A2(n13463), .ZN(n12174) );
  AOI21_X1 U14629 ( .B1(n13287), .B2(n12203), .A(n12174), .ZN(n12221) );
  NAND2_X1 U14630 ( .A1(n13287), .A2(n12215), .ZN(n12176) );
  NAND2_X1 U14631 ( .A1(n12214), .A2(n13463), .ZN(n12175) );
  NAND2_X1 U14632 ( .A1(n12176), .A2(n12175), .ZN(n12220) );
  NAND2_X1 U14633 ( .A1(n12221), .A2(n12220), .ZN(n12177) );
  AND2_X1 U14634 ( .A1(n12222), .A2(n12177), .ZN(n12178) );
  NAND2_X1 U14635 ( .A1(n12283), .A2(n12178), .ZN(n12219) );
  AND2_X1 U14636 ( .A1(n12215), .A2(n13352), .ZN(n12179) );
  AOI21_X1 U14637 ( .B1(n13661), .B2(n12203), .A(n12179), .ZN(n12218) );
  NAND2_X1 U14638 ( .A1(n13661), .A2(n12215), .ZN(n12181) );
  NAND2_X1 U14639 ( .A1(n12214), .A2(n13352), .ZN(n12180) );
  NAND2_X1 U14640 ( .A1(n12181), .A2(n12180), .ZN(n12217) );
  AND2_X1 U14641 ( .A1(n12218), .A2(n12217), .ZN(n12182) );
  AND2_X1 U14642 ( .A1(n12215), .A2(n13495), .ZN(n12183) );
  AOI21_X1 U14643 ( .B1(n13670), .B2(n12203), .A(n12183), .ZN(n12230) );
  NAND2_X1 U14644 ( .A1(n13670), .A2(n12215), .ZN(n12185) );
  NAND2_X1 U14645 ( .A1(n12214), .A2(n13495), .ZN(n12184) );
  NAND2_X1 U14646 ( .A1(n12185), .A2(n12184), .ZN(n12229) );
  AND2_X1 U14647 ( .A1(n12230), .A2(n12229), .ZN(n12186) );
  NAND2_X1 U14648 ( .A1(n13503), .A2(n12203), .ZN(n12188) );
  NAND2_X1 U14649 ( .A1(n12215), .A2(n13353), .ZN(n12187) );
  AND2_X1 U14650 ( .A1(n12214), .A2(n13353), .ZN(n12189) );
  AOI21_X1 U14651 ( .B1(n13503), .B2(n12202), .A(n12189), .ZN(n12193) );
  NAND2_X1 U14652 ( .A1(n7552), .A2(n12190), .ZN(n12191) );
  NOR2_X1 U14653 ( .A1(n7552), .A2(n12190), .ZN(n12235) );
  INV_X1 U14654 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n12611) );
  OR2_X1 U14655 ( .A1(n9502), .A2(n12611), .ZN(n12194) );
  INV_X1 U14656 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n15329) );
  OR2_X1 U14657 ( .A1(n12196), .A2(n15329), .ZN(n12200) );
  INV_X1 U14658 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n12197) );
  OR2_X1 U14659 ( .A1(n9496), .A2(n12197), .ZN(n12199) );
  INV_X1 U14660 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n13737) );
  OR2_X1 U14661 ( .A1(n6546), .A2(n13737), .ZN(n12198) );
  AND3_X1 U14662 ( .A1(n12200), .A2(n12199), .A3(n12198), .ZN(n13436) );
  NOR2_X1 U14663 ( .A1(n13436), .A2(n12293), .ZN(n12201) );
  AOI21_X1 U14664 ( .B1(n13426), .B2(n12202), .A(n12201), .ZN(n12239) );
  NAND2_X1 U14665 ( .A1(n13426), .A2(n12203), .ZN(n12209) );
  NAND2_X1 U14666 ( .A1(n12215), .A2(n13420), .ZN(n12292) );
  NAND2_X1 U14667 ( .A1(n9578), .A2(n10530), .ZN(n12287) );
  AND2_X1 U14668 ( .A1(n12204), .A2(n10529), .ZN(n12205) );
  AND2_X1 U14669 ( .A1(n12287), .A2(n12205), .ZN(n12206) );
  NAND2_X1 U14670 ( .A1(n12292), .A2(n12206), .ZN(n12207) );
  INV_X1 U14671 ( .A(n13436), .ZN(n13350) );
  NAND2_X1 U14672 ( .A1(n12207), .A2(n13350), .ZN(n12208) );
  NAND2_X1 U14673 ( .A1(n12209), .A2(n12208), .ZN(n12238) );
  INV_X1 U14674 ( .A(n12210), .ZN(n12213) );
  INV_X1 U14675 ( .A(n12211), .ZN(n12212) );
  AOI22_X1 U14676 ( .A1(n12239), .A2(n12238), .B1(n12213), .B2(n12212), .ZN(
        n12228) );
  AOI22_X1 U14677 ( .A1(n12166), .A2(n12215), .B1(n12214), .B2(n13420), .ZN(
        n12216) );
  AND2_X1 U14678 ( .A1(n12216), .A2(n12291), .ZN(n12227) );
  OR3_X1 U14679 ( .A1(n12219), .A2(n12218), .A3(n12217), .ZN(n12226) );
  INV_X1 U14680 ( .A(n12220), .ZN(n12224) );
  INV_X1 U14681 ( .A(n12221), .ZN(n12223) );
  NAND4_X1 U14682 ( .A1(n12283), .A2(n12224), .A3(n12223), .A4(n12222), .ZN(
        n12225) );
  OAI211_X1 U14683 ( .C1(n12228), .C2(n12227), .A(n12226), .B(n12225), .ZN(
        n12233) );
  NOR3_X1 U14684 ( .A1(n12231), .A2(n12230), .A3(n12229), .ZN(n12232) );
  AOI211_X1 U14685 ( .C1(n12235), .C2(n12234), .A(n12233), .B(n12232), .ZN(
        n12236) );
  NAND2_X1 U14686 ( .A1(n12237), .A2(n12236), .ZN(n12243) );
  INV_X1 U14687 ( .A(n12238), .ZN(n12241) );
  NAND2_X1 U14688 ( .A1(n12241), .A2(n12240), .ZN(n12242) );
  NAND2_X1 U14689 ( .A1(n12243), .A2(n12242), .ZN(n12304) );
  XNOR2_X1 U14690 ( .A(n13426), .B(n13436), .ZN(n12281) );
  NAND2_X1 U14691 ( .A1(n12245), .A2(n12244), .ZN(n13486) );
  NAND4_X1 U14692 ( .A1(n12248), .A2(n12247), .A3(n12246), .A4(n14960), .ZN(
        n12250) );
  NOR2_X1 U14693 ( .A1(n12250), .A2(n12249), .ZN(n12253) );
  NAND4_X1 U14694 ( .A1(n12254), .A2(n12253), .A3(n12252), .A4(n12251), .ZN(
        n12255) );
  NOR2_X1 U14695 ( .A1(n12256), .A2(n12255), .ZN(n12259) );
  NAND4_X1 U14696 ( .A1(n12260), .A2(n12259), .A3(n12258), .A4(n12257), .ZN(
        n12261) );
  OR4_X1 U14697 ( .A1(n12264), .A2(n12263), .A3(n12262), .A4(n12261), .ZN(
        n12265) );
  NOR2_X1 U14698 ( .A1(n12266), .A2(n12265), .ZN(n12269) );
  NAND4_X1 U14699 ( .A1(n12270), .A2(n12269), .A3(n12268), .A4(n12267), .ZN(
        n12271) );
  OR4_X1 U14700 ( .A1(n13584), .A2(n13597), .A3(n13616), .A4(n12271), .ZN(
        n12272) );
  NOR2_X1 U14701 ( .A1(n13565), .A2(n12272), .ZN(n12276) );
  NAND2_X1 U14702 ( .A1(n12274), .A2(n12273), .ZN(n13530) );
  NAND4_X1 U14703 ( .A1(n13509), .A2(n12276), .A3(n13530), .A4(n12275), .ZN(
        n12277) );
  NOR2_X1 U14704 ( .A1(n13486), .A2(n12277), .ZN(n12278) );
  NAND4_X1 U14705 ( .A1(n12279), .A2(n12278), .A3(n13471), .A4(n13493), .ZN(
        n12280) );
  NOR2_X1 U14706 ( .A1(n12281), .A2(n12280), .ZN(n12282) );
  NAND3_X1 U14707 ( .A1(n12283), .A2(n12282), .A3(n13433), .ZN(n12284) );
  XNOR2_X1 U14708 ( .A(n12284), .B(n7536), .ZN(n12286) );
  NAND2_X1 U14709 ( .A1(n12286), .A2(n12285), .ZN(n12295) );
  NOR2_X1 U14710 ( .A1(n9578), .A2(n12289), .ZN(n12290) );
  AOI211_X1 U14711 ( .C1(n10529), .C2(n12613), .A(n12305), .B(n12290), .ZN(
        n12294) );
  OAI211_X1 U14712 ( .C1(n12165), .C2(n12293), .A(n12292), .B(n12291), .ZN(
        n12299) );
  OAI211_X1 U14713 ( .C1(n12295), .C2(n10530), .A(n12294), .B(n12299), .ZN(
        n12296) );
  INV_X1 U14714 ( .A(n12296), .ZN(n12297) );
  NAND2_X1 U14715 ( .A1(n12304), .A2(n12297), .ZN(n12302) );
  OAI211_X1 U14716 ( .C1(n12304), .C2(n12303), .A(n12302), .B(n12301), .ZN(
        n12310) );
  NAND4_X1 U14717 ( .A1(n13462), .A2(n12306), .A3(n14953), .A4(n12305), .ZN(
        n12307) );
  OAI211_X1 U14718 ( .C1(n9578), .C2(n12308), .A(n12307), .B(P2_B_REG_SCAN_IN), 
        .ZN(n12309) );
  NAND2_X1 U14719 ( .A1(n12310), .A2(n12309), .ZN(P2_U3328) );
  OAI222_X1 U14720 ( .A1(n13768), .A2(n12312), .B1(n6551), .B2(n12311), .C1(
        n13418), .C2(P2_U3088), .ZN(P2_U3300) );
  XOR2_X1 U14721 ( .A(n12314), .B(n12313), .Z(n12328) );
  XNOR2_X1 U14722 ( .A(n12316), .B(n12315), .ZN(n12326) );
  OAI21_X1 U14723 ( .B1(n12319), .B2(n12318), .A(n12317), .ZN(n12320) );
  NAND2_X1 U14724 ( .A1(n12320), .A2(n15109), .ZN(n12323) );
  AOI21_X1 U14725 ( .B1(n15106), .B2(P3_ADDR_REG_8__SCAN_IN), .A(n12321), .ZN(
        n12322) );
  OAI211_X1 U14726 ( .C1(n15100), .C2(n12324), .A(n12323), .B(n12322), .ZN(
        n12325) );
  AOI21_X1 U14727 ( .B1(n15023), .B2(n12326), .A(n12325), .ZN(n12327) );
  OAI21_X1 U14728 ( .B1(n12328), .B2(n15102), .A(n12327), .ZN(P3_U3190) );
  XOR2_X1 U14729 ( .A(n12330), .B(n12329), .Z(n12342) );
  XNOR2_X1 U14730 ( .A(n8640), .B(n12331), .ZN(n12340) );
  OAI21_X1 U14731 ( .B1(P3_REG1_REG_7__SCAN_IN), .B2(n12333), .A(n12332), .ZN(
        n12334) );
  NAND2_X1 U14732 ( .A1(n12334), .A2(n15109), .ZN(n12337) );
  AOI21_X1 U14733 ( .B1(n15106), .B2(P3_ADDR_REG_7__SCAN_IN), .A(n12335), .ZN(
        n12336) );
  OAI211_X1 U14734 ( .C1(n15100), .C2(n12338), .A(n12337), .B(n12336), .ZN(
        n12339) );
  AOI21_X1 U14735 ( .B1(n15023), .B2(n12340), .A(n12339), .ZN(n12341) );
  OAI21_X1 U14736 ( .B1(n12342), .B2(n15102), .A(n12341), .ZN(P3_U3189) );
  XOR2_X1 U14737 ( .A(n12344), .B(n12343), .Z(n12358) );
  OAI21_X1 U14738 ( .B1(n12347), .B2(n12346), .A(n12345), .ZN(n12356) );
  AOI21_X1 U14739 ( .B1(n12350), .B2(n12349), .A(n12348), .ZN(n12354) );
  INV_X1 U14740 ( .A(n15109), .ZN(n15069) );
  INV_X1 U14741 ( .A(P3_REG3_REG_6__SCAN_IN), .ZN(n15460) );
  NOR2_X1 U14742 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15460), .ZN(n12710) );
  NOR2_X1 U14743 ( .A1(n15100), .A2(n12351), .ZN(n12352) );
  AOI211_X1 U14744 ( .C1(n15106), .C2(P3_ADDR_REG_6__SCAN_IN), .A(n12710), .B(
        n12352), .ZN(n12353) );
  OAI21_X1 U14745 ( .B1(n12354), .B2(n15069), .A(n12353), .ZN(n12355) );
  AOI21_X1 U14746 ( .B1(n15023), .B2(n12356), .A(n12355), .ZN(n12357) );
  OAI21_X1 U14747 ( .B1(n12358), .B2(n15102), .A(n12357), .ZN(P3_U3188) );
  NAND2_X1 U14748 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n14434), .ZN(n12359) );
  AOI22_X1 U14749 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(
        P1_DATAO_REG_30__SCAN_IN), .B1(n12611), .B2(n14431), .ZN(n12361) );
  XNOR2_X1 U14750 ( .A(n12367), .B(n12361), .ZN(n12588) );
  NAND2_X1 U14751 ( .A1(n12588), .A2(n12362), .ZN(n12365) );
  NAND2_X1 U14752 ( .A1(n12363), .A2(SI_30_), .ZN(n12364) );
  NOR2_X1 U14753 ( .A1(n14623), .A2(n12373), .ZN(n12568) );
  NAND2_X1 U14754 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(n12611), .ZN(n12366) );
  AOI22_X1 U14755 ( .A1(n12367), .A2(n12366), .B1(P1_DATAO_REG_30__SCAN_IN), 
        .B2(n14431), .ZN(n12369) );
  AOI22_X1 U14756 ( .A1(P2_DATAO_REG_31__SCAN_IN), .A2(n13769), .B1(
        P1_DATAO_REG_31__SCAN_IN), .B2(n14430), .ZN(n12368) );
  XNOR2_X1 U14757 ( .A(n12369), .B(n12368), .ZN(n13194) );
  NAND2_X1 U14758 ( .A1(n13194), .A2(n9017), .ZN(n12372) );
  NAND2_X1 U14759 ( .A1(n12370), .A2(SI_31_), .ZN(n12371) );
  INV_X1 U14760 ( .A(n12376), .ZN(n14610) );
  NAND2_X1 U14761 ( .A1(n12876), .A2(n12375), .ZN(n12569) );
  NAND2_X1 U14762 ( .A1(n14623), .A2(n12373), .ZN(n12374) );
  OR2_X1 U14763 ( .A1(n12876), .A2(n12375), .ZN(n12567) );
  OAI21_X1 U14764 ( .B1(n12377), .B2(n12376), .A(n12567), .ZN(n12378) );
  XOR2_X1 U14765 ( .A(n12859), .B(n12380), .Z(n12409) );
  INV_X1 U14766 ( .A(n12938), .ZN(n12546) );
  XNOR2_X1 U14767 ( .A(n12644), .B(n12974), .ZN(n12986) );
  NAND2_X1 U14768 ( .A1(n12410), .A2(n12958), .ZN(n12976) );
  INV_X1 U14769 ( .A(n12976), .ZN(n12397) );
  INV_X1 U14770 ( .A(n13071), .ZN(n12395) );
  INV_X1 U14771 ( .A(n13056), .ZN(n12394) );
  INV_X1 U14772 ( .A(n15142), .ZN(n12383) );
  NAND4_X1 U14773 ( .A1(n12386), .A2(n12385), .A3(n12384), .A4(n12383), .ZN(
        n12388) );
  NAND4_X1 U14774 ( .A1(n12450), .A2(n15124), .A3(n12433), .A4(n12437), .ZN(
        n12387) );
  NOR3_X1 U14775 ( .A1(n12388), .A2(n12387), .A3(n12465), .ZN(n12391) );
  NAND4_X1 U14776 ( .A1(n12391), .A2(n12476), .A3(n12390), .A4(n12389), .ZN(
        n12392) );
  OR4_X1 U14777 ( .A1(n12492), .A2(n12488), .A3(n12392), .A4(n6996), .ZN(
        n12393) );
  NOR4_X1 U14778 ( .A1(n13029), .A2(n12395), .A3(n12394), .A4(n12393), .ZN(
        n12396) );
  NAND4_X1 U14779 ( .A1(n13013), .A2(n12397), .A3(n12396), .A4(n13041), .ZN(
        n12398) );
  NOR4_X1 U14780 ( .A1(n12986), .A2(n13004), .A3(n12960), .A4(n12398), .ZN(
        n12399) );
  NAND3_X1 U14781 ( .A1(n12546), .A2(n12399), .A3(n12923), .ZN(n12400) );
  XOR2_X1 U14782 ( .A(n12859), .B(n12405), .Z(n12406) );
  INV_X1 U14783 ( .A(n12410), .ZN(n12412) );
  INV_X1 U14784 ( .A(n12958), .ZN(n12411) );
  MUX2_X1 U14785 ( .A(n12412), .B(n12411), .S(n9115), .Z(n12539) );
  MUX2_X1 U14786 ( .A(n12414), .B(n12739), .S(n9115), .Z(n12470) );
  INV_X1 U14787 ( .A(n12418), .ZN(n12425) );
  OAI21_X1 U14788 ( .B1(n12415), .B2(n12419), .A(n9115), .ZN(n12421) );
  INV_X1 U14789 ( .A(n12416), .ZN(n12583) );
  NAND3_X1 U14790 ( .A1(n12418), .A2(n12417), .A3(n12583), .ZN(n12420) );
  AOI22_X1 U14791 ( .A1(n12421), .A2(n12420), .B1(n15135), .B2(n12419), .ZN(
        n12423) );
  MUX2_X1 U14792 ( .A(n12549), .B(n12423), .S(n12422), .Z(n12424) );
  AOI211_X1 U14793 ( .C1(n12425), .C2(n9115), .A(n15115), .B(n12424), .ZN(
        n12435) );
  NAND2_X1 U14794 ( .A1(n12430), .A2(n12426), .ZN(n12429) );
  NAND2_X1 U14795 ( .A1(n12431), .A2(n12427), .ZN(n12428) );
  MUX2_X1 U14796 ( .A(n12429), .B(n12428), .S(n9115), .Z(n12434) );
  MUX2_X1 U14797 ( .A(n12431), .B(n12430), .S(n9115), .Z(n12432) );
  OAI211_X1 U14798 ( .C1(n12435), .C2(n12434), .A(n12433), .B(n12432), .ZN(
        n12438) );
  NAND2_X1 U14799 ( .A1(n12448), .A2(n12436), .ZN(n12441) );
  AOI22_X1 U14800 ( .A1(n12438), .A2(n12437), .B1(n9115), .B2(n12441), .ZN(
        n12445) );
  INV_X1 U14801 ( .A(n12439), .ZN(n12443) );
  NOR2_X1 U14802 ( .A1(n12441), .A2(n12440), .ZN(n12442) );
  MUX2_X1 U14803 ( .A(n12443), .B(n12442), .S(n9115), .Z(n12444) );
  NOR2_X1 U14804 ( .A1(n12445), .A2(n12444), .ZN(n12452) );
  AOI21_X1 U14805 ( .B1(n12447), .B2(n12446), .A(n9115), .ZN(n12451) );
  MUX2_X1 U14806 ( .A(n12448), .B(n12447), .S(n9115), .Z(n12449) );
  OAI211_X1 U14807 ( .C1(n12452), .C2(n12451), .A(n12450), .B(n12449), .ZN(
        n12467) );
  INV_X1 U14808 ( .A(n12453), .ZN(n12456) );
  INV_X1 U14809 ( .A(n12454), .ZN(n12455) );
  MUX2_X1 U14810 ( .A(n12456), .B(n12455), .S(n12549), .Z(n12458) );
  NOR2_X1 U14811 ( .A1(n12458), .A2(n12457), .ZN(n12466) );
  INV_X1 U14812 ( .A(n12459), .ZN(n12463) );
  NOR2_X1 U14813 ( .A1(n12461), .A2(n12460), .ZN(n12462) );
  MUX2_X1 U14814 ( .A(n12463), .B(n12462), .S(n12549), .Z(n12464) );
  AOI211_X1 U14815 ( .C1(n12467), .C2(n12466), .A(n12465), .B(n12464), .ZN(
        n12468) );
  AOI211_X1 U14816 ( .C1(n12471), .C2(n12470), .A(n12469), .B(n12468), .ZN(
        n12472) );
  AOI21_X1 U14817 ( .B1(n7000), .B2(n9115), .A(n12472), .ZN(n12484) );
  INV_X1 U14818 ( .A(n12473), .ZN(n12475) );
  INV_X1 U14819 ( .A(n12474), .ZN(n12485) );
  AOI211_X1 U14820 ( .C1(n12477), .C2(n12476), .A(n12475), .B(n12485), .ZN(
        n12481) );
  INV_X1 U14821 ( .A(n12478), .ZN(n12486) );
  NOR2_X1 U14822 ( .A1(n12486), .A2(n6999), .ZN(n12480) );
  MUX2_X1 U14823 ( .A(n12481), .B(n12480), .S(n9115), .Z(n12482) );
  OAI21_X1 U14824 ( .B1(n12484), .B2(n12483), .A(n12482), .ZN(n12495) );
  MUX2_X1 U14825 ( .A(n12486), .B(n12485), .S(n9115), .Z(n12487) );
  NOR2_X1 U14826 ( .A1(n12488), .A2(n12487), .ZN(n12494) );
  INV_X1 U14827 ( .A(n12489), .ZN(n12491) );
  MUX2_X1 U14828 ( .A(n12491), .B(n12490), .S(n9115), .Z(n12493) );
  AOI211_X1 U14829 ( .C1(n12495), .C2(n12494), .A(n12493), .B(n12492), .ZN(
        n12501) );
  INV_X1 U14830 ( .A(n12496), .ZN(n12499) );
  INV_X1 U14831 ( .A(n12497), .ZN(n12498) );
  MUX2_X1 U14832 ( .A(n12499), .B(n12498), .S(n9115), .Z(n12500) );
  OAI21_X1 U14833 ( .B1(n12501), .B2(n12500), .A(n13071), .ZN(n12507) );
  INV_X1 U14834 ( .A(n12509), .ZN(n12504) );
  INV_X1 U14835 ( .A(n12502), .ZN(n12503) );
  OAI21_X1 U14836 ( .B1(n12504), .B2(n12503), .A(n9115), .ZN(n12506) );
  INV_X1 U14837 ( .A(n13042), .ZN(n12505) );
  AOI21_X1 U14838 ( .B1(n12507), .B2(n12506), .A(n12505), .ZN(n12511) );
  AOI21_X1 U14839 ( .B1(n13042), .B2(n12508), .A(n9115), .ZN(n12510) );
  OAI22_X1 U14840 ( .A1(n12511), .A2(n12510), .B1(n12509), .B2(n9115), .ZN(
        n12512) );
  NAND3_X1 U14841 ( .A1(n12512), .A2(n13023), .A3(n13041), .ZN(n12527) );
  NOR2_X1 U14842 ( .A1(n13126), .A2(n13053), .ZN(n12515) );
  INV_X1 U14843 ( .A(n12513), .ZN(n12514) );
  AOI211_X1 U14844 ( .C1(n12515), .C2(n12517), .A(n12514), .B(n12523), .ZN(
        n12522) );
  INV_X1 U14845 ( .A(n12516), .ZN(n12520) );
  INV_X1 U14846 ( .A(n12517), .ZN(n12519) );
  INV_X1 U14847 ( .A(n12518), .ZN(n12524) );
  AOI211_X1 U14848 ( .C1(n13023), .C2(n12520), .A(n12519), .B(n12524), .ZN(
        n12521) );
  MUX2_X1 U14849 ( .A(n12522), .B(n12521), .S(n9115), .Z(n12526) );
  MUX2_X1 U14850 ( .A(n12524), .B(n12523), .S(n9115), .Z(n12525) );
  AOI211_X1 U14851 ( .C1(n12527), .C2(n12526), .A(n13004), .B(n12525), .ZN(
        n12533) );
  INV_X1 U14852 ( .A(n12528), .ZN(n12531) );
  INV_X1 U14853 ( .A(n13000), .ZN(n13171) );
  NOR2_X1 U14854 ( .A1(n13171), .A2(n12529), .ZN(n12530) );
  MUX2_X1 U14855 ( .A(n12531), .B(n12530), .S(n9115), .Z(n12532) );
  NOR3_X1 U14856 ( .A1(n12533), .A2(n12986), .A3(n12532), .ZN(n12537) );
  NOR2_X1 U14857 ( .A1(n12644), .A2(n12549), .ZN(n12535) );
  INV_X1 U14858 ( .A(n12644), .ZN(n13167) );
  NOR2_X1 U14859 ( .A1(n13167), .A2(n9115), .ZN(n12534) );
  MUX2_X1 U14860 ( .A(n12535), .B(n12534), .S(n12974), .Z(n12536) );
  NOR3_X1 U14861 ( .A1(n12537), .A2(n12536), .A3(n12976), .ZN(n12538) );
  OAI33_X1 U14862 ( .A1(n9115), .A2(n12969), .A3(n12732), .B1(n12960), .B2(
        n12539), .B3(n12538), .ZN(n12547) );
  NAND2_X1 U14863 ( .A1(n12542), .A2(n12939), .ZN(n12541) );
  NAND2_X1 U14864 ( .A1(n12541), .A2(n12540), .ZN(n12544) );
  INV_X1 U14865 ( .A(n12542), .ZN(n12543) );
  MUX2_X1 U14866 ( .A(n12544), .B(n12543), .S(n12549), .Z(n12545) );
  AOI21_X1 U14867 ( .B1(n12547), .B2(n12546), .A(n12545), .ZN(n12552) );
  INV_X1 U14868 ( .A(n12548), .ZN(n13155) );
  MUX2_X1 U14869 ( .A(n12549), .B(n12548), .S(n12905), .Z(n12550) );
  AOI21_X1 U14870 ( .B1(n13155), .B2(n9115), .A(n12550), .ZN(n12551) );
  AOI211_X1 U14871 ( .C1(n12552), .C2(n12923), .A(n12551), .B(n12899), .ZN(
        n12558) );
  INV_X1 U14872 ( .A(n12553), .ZN(n12556) );
  INV_X1 U14873 ( .A(n12554), .ZN(n12555) );
  MUX2_X1 U14874 ( .A(n12556), .B(n12555), .S(n9115), .Z(n12557) );
  OAI211_X1 U14875 ( .C1(n12558), .C2(n12557), .A(n12881), .B(n12889), .ZN(
        n12565) );
  OAI21_X1 U14876 ( .B1(n12560), .B2(n12559), .A(n12565), .ZN(n12566) );
  INV_X1 U14877 ( .A(n12561), .ZN(n12563) );
  OAI21_X1 U14878 ( .B1(n12563), .B2(n9115), .A(n12562), .ZN(n12564) );
  AOI22_X1 U14879 ( .A1(n12566), .A2(n9115), .B1(n12565), .B2(n12564), .ZN(
        n12572) );
  INV_X1 U14880 ( .A(n12567), .ZN(n12571) );
  INV_X1 U14881 ( .A(n12568), .ZN(n12570) );
  INV_X1 U14882 ( .A(n12573), .ZN(n12575) );
  AOI21_X1 U14883 ( .B1(n12576), .B2(n12575), .A(n12574), .ZN(n12577) );
  MUX2_X1 U14884 ( .A(n15134), .B(n12578), .S(n12577), .Z(n12579) );
  NOR3_X1 U14885 ( .A1(n12582), .A2(n13205), .A3(n12581), .ZN(n12585) );
  OAI21_X1 U14886 ( .B1(n12583), .B2(n12586), .A(P3_B_REG_SCAN_IN), .ZN(n12584) );
  OAI22_X1 U14887 ( .A1(n12587), .A2(n12586), .B1(n12585), .B2(n12584), .ZN(
        P3_U3296) );
  INV_X1 U14888 ( .A(n12588), .ZN(n12590) );
  INV_X1 U14889 ( .A(SI_30_), .ZN(n12589) );
  OAI222_X1 U14890 ( .A1(P3_U3151), .A2(n12591), .B1(n13213), .B2(n12590), 
        .C1(n12589), .C2(n13217), .ZN(P3_U3265) );
  OAI222_X1 U14891 ( .A1(n13768), .A2(n15400), .B1(n6551), .B2(n12592), .C1(
        n9579), .C2(P2_U3088), .ZN(P2_U3307) );
  NAND2_X1 U14892 ( .A1(n12593), .A2(n14284), .ZN(n12601) );
  OAI22_X1 U14893 ( .A1(n12596), .A2(n12595), .B1(n12594), .B2(n14777), .ZN(
        n12599) );
  NOR2_X1 U14894 ( .A1(n14281), .A2(n12597), .ZN(n12598) );
  AOI211_X1 U14895 ( .C1(n14281), .C2(P1_REG2_REG_29__SCAN_IN), .A(n12599), 
        .B(n12598), .ZN(n12600) );
  OAI211_X1 U14896 ( .C1(n7018), .C2(n14271), .A(n12601), .B(n12600), .ZN(
        n12602) );
  AOI21_X1 U14897 ( .B1(n12603), .B2(n14235), .A(n12602), .ZN(n12604) );
  OAI21_X1 U14898 ( .B1(n12605), .B2(n14237), .A(n12604), .ZN(P1_U3356) );
  INV_X1 U14899 ( .A(n13776), .ZN(n12606) );
  OAI222_X1 U14900 ( .A1(n14433), .A2(n12607), .B1(n12610), .B2(n12606), .C1(
        n8158), .C2(P1_U3086), .ZN(P1_U3327) );
  OAI222_X1 U14901 ( .A1(n14433), .A2(n8900), .B1(n12610), .B2(n12609), .C1(
        n12608), .C2(P1_U3086), .ZN(P1_U3334) );
  OAI222_X1 U14902 ( .A1(n13768), .A2(n12615), .B1(n6551), .B2(n12614), .C1(
        P2_U3088), .C2(n12613), .ZN(P2_U3308) );
  INV_X1 U14903 ( .A(n13084), .ZN(n12896) );
  OAI21_X1 U14904 ( .B1(n12618), .B2(n12617), .A(n12616), .ZN(n12619) );
  NAND2_X1 U14905 ( .A1(n12619), .A2(n12722), .ZN(n12624) );
  AOI22_X1 U14906 ( .A1(n12894), .A2(n12724), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12620) );
  OAI21_X1 U14907 ( .B1(n12926), .B2(n12726), .A(n12620), .ZN(n12621) );
  AOI21_X1 U14908 ( .B1(n12622), .B2(n12728), .A(n12621), .ZN(n12623) );
  OAI211_X1 U14909 ( .C1(n12896), .C2(n12731), .A(n12624), .B(n12623), .ZN(
        P3_U3154) );
  INV_X1 U14910 ( .A(n12625), .ZN(n12670) );
  AOI21_X1 U14911 ( .B1(n12732), .B2(n12626), .A(n12670), .ZN(n12631) );
  AOI22_X1 U14912 ( .A1(n12956), .A2(n12709), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12628) );
  NAND2_X1 U14913 ( .A1(n12967), .A2(n12724), .ZN(n12627) );
  OAI211_X1 U14914 ( .C1(n12925), .C2(n12691), .A(n12628), .B(n12627), .ZN(
        n12629) );
  AOI21_X1 U14915 ( .B1(n13101), .B2(n12702), .A(n12629), .ZN(n12630) );
  OAI21_X1 U14916 ( .B1(n12631), .B2(n12704), .A(n12630), .ZN(P3_U3156) );
  XNOR2_X1 U14917 ( .A(n12632), .B(n12633), .ZN(n12638) );
  NAND2_X1 U14918 ( .A1(n12709), .A2(n12733), .ZN(n12634) );
  NAND2_X1 U14919 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n12858)
         );
  OAI211_X1 U14920 ( .C1(n13009), .C2(n12691), .A(n12634), .B(n12858), .ZN(
        n12636) );
  NOR2_X1 U14921 ( .A1(n13175), .A2(n12731), .ZN(n12635) );
  AOI211_X1 U14922 ( .C1(n13016), .C2(n12724), .A(n12636), .B(n12635), .ZN(
        n12637) );
  OAI21_X1 U14923 ( .B1(n12638), .B2(n12704), .A(n12637), .ZN(P3_U3159) );
  AOI21_X1 U14924 ( .B1(n12640), .B2(n12639), .A(n6656), .ZN(n12647) );
  OAI22_X1 U14925 ( .A1(n13009), .A2(n12726), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12641), .ZN(n12643) );
  NOR2_X1 U14926 ( .A1(n12985), .A2(n12691), .ZN(n12642) );
  AOI211_X1 U14927 ( .C1(n12988), .C2(n12724), .A(n12643), .B(n12642), .ZN(
        n12646) );
  NAND2_X1 U14928 ( .A1(n12644), .A2(n12702), .ZN(n12645) );
  OAI211_X1 U14929 ( .C1(n12647), .C2(n12704), .A(n12646), .B(n12645), .ZN(
        P3_U3163) );
  INV_X1 U14930 ( .A(n12648), .ZN(n12671) );
  INV_X1 U14931 ( .A(n12649), .ZN(n12651) );
  NOR3_X1 U14932 ( .A1(n12671), .A2(n12651), .A3(n12650), .ZN(n12654) );
  INV_X1 U14933 ( .A(n12652), .ZN(n12653) );
  OAI21_X1 U14934 ( .B1(n12654), .B2(n12653), .A(n12722), .ZN(n12659) );
  AOI22_X1 U14935 ( .A1(n12930), .A2(n12724), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12655) );
  OAI21_X1 U14936 ( .B1(n12925), .B2(n12726), .A(n12655), .ZN(n12656) );
  AOI21_X1 U14937 ( .B1(n12657), .B2(n12728), .A(n12656), .ZN(n12658) );
  OAI211_X1 U14938 ( .C1(n13155), .C2(n12731), .A(n12659), .B(n12658), .ZN(
        P3_U3165) );
  XNOR2_X1 U14939 ( .A(n12661), .B(n12660), .ZN(n12666) );
  NAND2_X1 U14940 ( .A1(n12728), .A2(n12733), .ZN(n12662) );
  NAND2_X1 U14941 ( .A1(P3_U3151), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n14581)
         );
  OAI211_X1 U14942 ( .C1(n13068), .C2(n12726), .A(n12662), .B(n14581), .ZN(
        n12664) );
  INV_X1 U14943 ( .A(n13126), .ZN(n13048) );
  NOR2_X1 U14944 ( .A1(n13048), .A2(n12731), .ZN(n12663) );
  AOI211_X1 U14945 ( .C1(n13046), .C2(n12724), .A(n12664), .B(n12663), .ZN(
        n12665) );
  OAI21_X1 U14946 ( .B1(n12666), .B2(n12704), .A(n12665), .ZN(P3_U3168) );
  INV_X1 U14947 ( .A(n12667), .ZN(n12669) );
  NOR3_X1 U14948 ( .A1(n12670), .A2(n12669), .A3(n12668), .ZN(n12672) );
  OAI21_X1 U14949 ( .B1(n12672), .B2(n12671), .A(n12722), .ZN(n12677) );
  INV_X1 U14950 ( .A(n12948), .ZN(n12674) );
  AOI22_X1 U14951 ( .A1(n12732), .A2(n12709), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12673) );
  OAI21_X1 U14952 ( .B1(n12674), .B2(n12700), .A(n12673), .ZN(n12675) );
  AOI21_X1 U14953 ( .B1(n12728), .B2(n12905), .A(n12675), .ZN(n12676) );
  OAI211_X1 U14954 ( .C1(n13159), .C2(n12731), .A(n12677), .B(n12676), .ZN(
        P3_U3169) );
  CLKBUF_X1 U14955 ( .A(n12678), .Z(n12680) );
  XNOR2_X1 U14956 ( .A(n12680), .B(n12679), .ZN(n12685) );
  AOI22_X1 U14957 ( .A1(n12995), .A2(n12709), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12682) );
  NAND2_X1 U14958 ( .A1(n12724), .A2(n12999), .ZN(n12681) );
  OAI211_X1 U14959 ( .C1(n12974), .C2(n12691), .A(n12682), .B(n12681), .ZN(
        n12683) );
  AOI21_X1 U14960 ( .B1(n13000), .B2(n12702), .A(n12683), .ZN(n12684) );
  OAI21_X1 U14961 ( .B1(n12685), .B2(n12704), .A(n12684), .ZN(P3_U3173) );
  INV_X1 U14962 ( .A(n12686), .ZN(n13164) );
  OAI21_X1 U14963 ( .B1(n12985), .B2(n12688), .A(n12687), .ZN(n12689) );
  NAND2_X1 U14964 ( .A1(n12689), .A2(n12722), .ZN(n12694) );
  AOI22_X1 U14965 ( .A1(n12996), .A2(n12709), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12690) );
  OAI21_X1 U14966 ( .B1(n12975), .B2(n12691), .A(n12690), .ZN(n12692) );
  AOI21_X1 U14967 ( .B1(n12978), .B2(n12724), .A(n12692), .ZN(n12693) );
  OAI211_X1 U14968 ( .C1(n13164), .C2(n12731), .A(n12694), .B(n12693), .ZN(
        P3_U3175) );
  XNOR2_X1 U14969 ( .A(n12696), .B(n12695), .ZN(n12705) );
  INV_X1 U14970 ( .A(n12697), .ZN(n13026) );
  NAND2_X1 U14971 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n14606)
         );
  OAI21_X1 U14972 ( .B1(n13053), .B2(n12726), .A(n14606), .ZN(n12698) );
  AOI21_X1 U14973 ( .B1(n12728), .B2(n12995), .A(n12698), .ZN(n12699) );
  OAI21_X1 U14974 ( .B1(n13026), .B2(n12700), .A(n12699), .ZN(n12701) );
  AOI21_X1 U14975 ( .B1(n13122), .B2(n12702), .A(n12701), .ZN(n12703) );
  OAI21_X1 U14976 ( .B1(n12705), .B2(n12704), .A(n12703), .ZN(P3_U3178) );
  OAI211_X1 U14977 ( .C1(n12708), .C2(n12707), .A(n12706), .B(n12722), .ZN(
        n12718) );
  NAND2_X1 U14978 ( .A1(n12709), .A2(n12743), .ZN(n12712) );
  INV_X1 U14979 ( .A(n12710), .ZN(n12711) );
  OAI211_X1 U14980 ( .C1(n12731), .C2(n15178), .A(n12712), .B(n12711), .ZN(
        n12713) );
  INV_X1 U14981 ( .A(n12713), .ZN(n12717) );
  NAND2_X1 U14982 ( .A1(n12724), .A2(n12714), .ZN(n12716) );
  NAND2_X1 U14983 ( .A1(n12728), .A2(n12741), .ZN(n12715) );
  NAND4_X1 U14984 ( .A1(n12718), .A2(n12717), .A3(n12716), .A4(n12715), .ZN(
        P3_U3179) );
  INV_X1 U14985 ( .A(n12913), .ZN(n13151) );
  OAI21_X1 U14986 ( .B1(n12721), .B2(n12720), .A(n12719), .ZN(n12723) );
  NAND2_X1 U14987 ( .A1(n12723), .A2(n12722), .ZN(n12730) );
  AOI22_X1 U14988 ( .A1(n12909), .A2(n12724), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12725) );
  OAI21_X1 U14989 ( .B1(n12943), .B2(n12726), .A(n12725), .ZN(n12727) );
  AOI21_X1 U14990 ( .B1(n12906), .B2(n12728), .A(n12727), .ZN(n12729) );
  OAI211_X1 U14991 ( .C1(n13151), .C2(n12731), .A(n12730), .B(n12729), .ZN(
        P3_U3180) );
  MUX2_X1 U14992 ( .A(n12876), .B(P3_DATAO_REG_29__SCAN_IN), .S(n12745), .Z(
        P3_U3520) );
  MUX2_X1 U14993 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(n12906), .S(P3_U3897), .Z(
        P3_U3518) );
  MUX2_X1 U14994 ( .A(n12905), .B(P3_DATAO_REG_25__SCAN_IN), .S(n12745), .Z(
        P3_U3516) );
  MUX2_X1 U14995 ( .A(n12957), .B(P3_DATAO_REG_24__SCAN_IN), .S(n12745), .Z(
        P3_U3515) );
  MUX2_X1 U14996 ( .A(n12732), .B(P3_DATAO_REG_23__SCAN_IN), .S(n12745), .Z(
        P3_U3514) );
  MUX2_X1 U14997 ( .A(n12956), .B(P3_DATAO_REG_22__SCAN_IN), .S(n12745), .Z(
        P3_U3513) );
  MUX2_X1 U14998 ( .A(n12996), .B(P3_DATAO_REG_21__SCAN_IN), .S(n12745), .Z(
        P3_U3512) );
  MUX2_X1 U14999 ( .A(n12995), .B(P3_DATAO_REG_19__SCAN_IN), .S(n12745), .Z(
        P3_U3510) );
  MUX2_X1 U15000 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(n12733), .S(P3_U3897), .Z(
        P3_U3509) );
  MUX2_X1 U15001 ( .A(n12734), .B(P3_DATAO_REG_16__SCAN_IN), .S(n12745), .Z(
        P3_U3507) );
  MUX2_X1 U15002 ( .A(n12735), .B(P3_DATAO_REG_15__SCAN_IN), .S(n12745), .Z(
        P3_U3506) );
  MUX2_X1 U15003 ( .A(n12736), .B(P3_DATAO_REG_13__SCAN_IN), .S(n12745), .Z(
        P3_U3504) );
  MUX2_X1 U15004 ( .A(n12737), .B(P3_DATAO_REG_12__SCAN_IN), .S(n12745), .Z(
        P3_U3503) );
  MUX2_X1 U15005 ( .A(n12738), .B(P3_DATAO_REG_10__SCAN_IN), .S(n12745), .Z(
        P3_U3501) );
  MUX2_X1 U15006 ( .A(n12739), .B(P3_DATAO_REG_9__SCAN_IN), .S(n12745), .Z(
        P3_U3500) );
  MUX2_X1 U15007 ( .A(n12740), .B(P3_DATAO_REG_8__SCAN_IN), .S(n12745), .Z(
        P3_U3499) );
  MUX2_X1 U15008 ( .A(n12741), .B(P3_DATAO_REG_7__SCAN_IN), .S(n12745), .Z(
        P3_U3498) );
  MUX2_X1 U15009 ( .A(n12742), .B(P3_DATAO_REG_6__SCAN_IN), .S(n12745), .Z(
        P3_U3497) );
  MUX2_X1 U15010 ( .A(n12743), .B(P3_DATAO_REG_5__SCAN_IN), .S(n12745), .Z(
        P3_U3496) );
  MUX2_X1 U15011 ( .A(n12744), .B(P3_DATAO_REG_4__SCAN_IN), .S(n12745), .Z(
        P3_U3495) );
  MUX2_X1 U15012 ( .A(n15120), .B(P3_DATAO_REG_3__SCAN_IN), .S(n12745), .Z(
        P3_U3494) );
  MUX2_X1 U15013 ( .A(n15137), .B(P3_DATAO_REG_2__SCAN_IN), .S(n12745), .Z(
        P3_U3493) );
  MUX2_X1 U15014 ( .A(n15121), .B(P3_DATAO_REG_1__SCAN_IN), .S(n12745), .Z(
        P3_U3492) );
  MUX2_X1 U15015 ( .A(n15138), .B(P3_DATAO_REG_0__SCAN_IN), .S(n12745), .Z(
        P3_U3491) );
  INV_X1 U15016 ( .A(n12772), .ZN(n12783) );
  OR2_X1 U15017 ( .A1(n12751), .A2(n12746), .ZN(n12747) );
  AOI21_X1 U15018 ( .B1(n11722), .B2(n12749), .A(n12767), .ZN(n12765) );
  NAND2_X1 U15019 ( .A1(P3_REG1_REG_13__SCAN_IN), .A2(n12752), .ZN(n12773) );
  OAI21_X1 U15020 ( .B1(P3_REG1_REG_13__SCAN_IN), .B2(n12752), .A(n12773), 
        .ZN(n12763) );
  MUX2_X1 U15021 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n13209), .Z(n12782) );
  XNOR2_X1 U15022 ( .A(n12782), .B(n12783), .ZN(n12756) );
  NAND2_X1 U15023 ( .A1(n12757), .A2(n12756), .ZN(n12790) );
  OAI21_X1 U15024 ( .B1(n12757), .B2(n12756), .A(n12790), .ZN(n12758) );
  NAND2_X1 U15025 ( .A1(n12758), .A2(n15085), .ZN(n12761) );
  AOI21_X1 U15026 ( .B1(n15106), .B2(P3_ADDR_REG_13__SCAN_IN), .A(n12759), 
        .ZN(n12760) );
  OAI211_X1 U15027 ( .C1(n15100), .C2(n12772), .A(n12761), .B(n12760), .ZN(
        n12762) );
  AOI21_X1 U15028 ( .B1(n15109), .B2(n12763), .A(n12762), .ZN(n12764) );
  OAI21_X1 U15029 ( .B1(n12765), .B2(n15113), .A(n12764), .ZN(P3_U3195) );
  NAND2_X1 U15030 ( .A1(n12781), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n12805) );
  NAND2_X1 U15031 ( .A1(n12776), .A2(n12769), .ZN(n12770) );
  NAND2_X1 U15032 ( .A1(n12805), .A2(n12770), .ZN(n12785) );
  AOI21_X1 U15033 ( .B1(n6653), .B2(n12785), .A(n12798), .ZN(n12797) );
  NAND2_X1 U15034 ( .A1(n12772), .A2(n12771), .ZN(n12774) );
  NAND2_X1 U15035 ( .A1(n12774), .A2(n12773), .ZN(n12778) );
  NAND2_X1 U15036 ( .A1(n12781), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n12804) );
  INV_X1 U15037 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n12775) );
  NAND2_X1 U15038 ( .A1(n12776), .A2(n12775), .ZN(n12777) );
  AND2_X1 U15039 ( .A1(n12804), .A2(n12777), .ZN(n12786) );
  NAND2_X1 U15040 ( .A1(n12786), .A2(n12778), .ZN(n12802) );
  OAI21_X1 U15041 ( .B1(n12778), .B2(n12786), .A(n12802), .ZN(n12795) );
  AOI21_X1 U15042 ( .B1(n15106), .B2(P3_ADDR_REG_14__SCAN_IN), .A(n12779), 
        .ZN(n12780) );
  OAI21_X1 U15043 ( .B1(n15100), .B2(n12781), .A(n12780), .ZN(n12794) );
  INV_X1 U15044 ( .A(n12782), .ZN(n12784) );
  NAND2_X1 U15045 ( .A1(n12784), .A2(n12783), .ZN(n12789) );
  INV_X1 U15046 ( .A(n12785), .ZN(n12787) );
  MUX2_X1 U15047 ( .A(n12787), .B(n12786), .S(n13209), .Z(n12788) );
  NAND3_X1 U15048 ( .A1(n12790), .A2(n12789), .A3(n12788), .ZN(n12807) );
  INV_X1 U15049 ( .A(n12807), .ZN(n12792) );
  AOI21_X1 U15050 ( .B1(n12790), .B2(n12789), .A(n12788), .ZN(n12791) );
  NOR3_X1 U15051 ( .A1(n12792), .A2(n12791), .A3(n15102), .ZN(n12793) );
  AOI211_X1 U15052 ( .C1(n15109), .C2(n12795), .A(n12794), .B(n12793), .ZN(
        n12796) );
  OAI21_X1 U15053 ( .B1(n12797), .B2(n15113), .A(n12796), .ZN(P3_U3196) );
  INV_X1 U15054 ( .A(n12798), .ZN(n12799) );
  XNOR2_X1 U15055 ( .A(n12833), .B(n12832), .ZN(n12800) );
  AOI21_X1 U15056 ( .B1(n12801), .B2(n12800), .A(n12834), .ZN(n12817) );
  OAI21_X1 U15057 ( .B1(P3_REG1_REG_15__SCAN_IN), .B2(n12803), .A(n12819), 
        .ZN(n12815) );
  MUX2_X1 U15058 ( .A(P3_REG2_REG_15__SCAN_IN), .B(P3_REG1_REG_15__SCAN_IN), 
        .S(n13209), .Z(n12809) );
  MUX2_X1 U15059 ( .A(n12805), .B(n12804), .S(n13209), .Z(n12806) );
  NAND2_X1 U15060 ( .A1(n12807), .A2(n12806), .ZN(n12822) );
  AOI21_X1 U15061 ( .B1(n12809), .B2(n12808), .A(n12823), .ZN(n12813) );
  INV_X1 U15062 ( .A(n15106), .ZN(n15028) );
  INV_X1 U15063 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n14475) );
  OAI21_X1 U15064 ( .B1(n15028), .B2(n14475), .A(n12810), .ZN(n12811) );
  AOI21_X1 U15065 ( .B1(n12824), .B2(n15031), .A(n12811), .ZN(n12812) );
  OAI21_X1 U15066 ( .B1(n12813), .B2(n15102), .A(n12812), .ZN(n12814) );
  AOI21_X1 U15067 ( .B1(n15109), .B2(n12815), .A(n12814), .ZN(n12816) );
  OAI21_X1 U15068 ( .B1(n12817), .B2(n15113), .A(n12816), .ZN(P3_U3197) );
  NAND2_X1 U15069 ( .A1(n12833), .A2(n12818), .ZN(n12820) );
  INV_X1 U15070 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n13132) );
  XNOR2_X1 U15071 ( .A(n12837), .B(n13132), .ZN(n12852) );
  XNOR2_X1 U15072 ( .A(n12849), .B(n12852), .ZN(n12842) );
  INV_X1 U15073 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n14537) );
  OAI21_X1 U15074 ( .B1(n15028), .B2(n14537), .A(n12821), .ZN(n12831) );
  INV_X1 U15075 ( .A(n12822), .ZN(n12825) );
  MUX2_X1 U15076 ( .A(n12836), .B(n13132), .S(n13209), .Z(n12826) );
  NAND2_X1 U15077 ( .A1(n12826), .A2(n12837), .ZN(n12862) );
  INV_X1 U15078 ( .A(n12862), .ZN(n12827) );
  NOR2_X1 U15079 ( .A1(n12837), .A2(n12836), .ZN(n12843) );
  NOR2_X1 U15080 ( .A1(n12837), .A2(n13132), .ZN(n12850) );
  MUX2_X1 U15081 ( .A(n12843), .B(n12850), .S(n13209), .Z(n12863) );
  NOR2_X1 U15082 ( .A1(n12827), .A2(n12863), .ZN(n12828) );
  XNOR2_X1 U15083 ( .A(n12864), .B(n12828), .ZN(n12829) );
  NOR2_X1 U15084 ( .A1(n12829), .A2(n15102), .ZN(n12830) );
  AOI211_X1 U15085 ( .C1(n15031), .C2(n12837), .A(n12831), .B(n12830), .ZN(
        n12841) );
  AND2_X1 U15086 ( .A1(n12833), .A2(n12832), .ZN(n12835) );
  AND2_X1 U15087 ( .A1(n12837), .A2(n12836), .ZN(n12838) );
  OAI21_X1 U15088 ( .B1(n6603), .B2(n6678), .A(n12845), .ZN(n12839) );
  NAND2_X1 U15089 ( .A1(n12839), .A2(n15023), .ZN(n12840) );
  OAI211_X1 U15090 ( .C1(n15069), .C2(n12842), .A(n12841), .B(n12840), .ZN(
        P3_U3198) );
  INV_X1 U15091 ( .A(n12843), .ZN(n12844) );
  NOR2_X1 U15092 ( .A1(n14580), .A2(n12846), .ZN(n12847) );
  NOR2_X1 U15093 ( .A1(n8824), .A2(n14577), .ZN(n14576) );
  XNOR2_X1 U15094 ( .A(n12856), .B(P3_REG2_REG_18__SCAN_IN), .ZN(n14602) );
  OAI21_X1 U15095 ( .B1(n14592), .B2(n13027), .A(n14601), .ZN(n12848) );
  XNOR2_X1 U15096 ( .A(n12859), .B(P3_REG2_REG_19__SCAN_IN), .ZN(n12861) );
  XNOR2_X1 U15097 ( .A(n12848), .B(n12861), .ZN(n12872) );
  INV_X1 U15098 ( .A(n12849), .ZN(n12853) );
  INV_X1 U15099 ( .A(n12850), .ZN(n12851) );
  OAI21_X1 U15100 ( .B1(n12853), .B2(n12852), .A(n12851), .ZN(n12854) );
  NAND2_X1 U15101 ( .A1(n12865), .A2(n12854), .ZN(n12855) );
  XNOR2_X1 U15102 ( .A(n12854), .B(n14580), .ZN(n14579) );
  XNOR2_X1 U15103 ( .A(n14592), .B(P3_REG1_REG_18__SCAN_IN), .ZN(n14593) );
  XNOR2_X1 U15104 ( .A(n12859), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n12860) );
  NAND2_X1 U15105 ( .A1(n15106), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n12857) );
  OAI211_X1 U15106 ( .C1(n15100), .C2(n12859), .A(n12858), .B(n12857), .ZN(
        n12869) );
  MUX2_X1 U15107 ( .A(n12861), .B(n12860), .S(n13209), .Z(n12868) );
  MUX2_X1 U15108 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n13209), .Z(n12866) );
  XNOR2_X1 U15109 ( .A(n12866), .B(n12865), .ZN(n14586) );
  NOR2_X1 U15110 ( .A1(n14585), .A2(n14586), .ZN(n14584) );
  AOI21_X1 U15111 ( .B1(n12866), .B2(n12865), .A(n14584), .ZN(n12867) );
  XNOR2_X1 U15112 ( .A(n12867), .B(n14592), .ZN(n14596) );
  MUX2_X1 U15113 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n13209), .Z(n14597) );
  NOR2_X1 U15114 ( .A1(n14596), .A2(n14597), .ZN(n14595) );
  OAI21_X1 U15115 ( .B1(n12872), .B2(n15113), .A(n12871), .ZN(P3_U3201) );
  NAND2_X1 U15116 ( .A1(n12873), .A2(n12881), .ZN(n12874) );
  NAND3_X1 U15117 ( .A1(n12875), .A2(n15143), .A3(n12874), .ZN(n12878) );
  AOI22_X1 U15118 ( .A1(n12906), .A2(n15139), .B1(n15136), .B2(n12876), .ZN(
        n12877) );
  NAND2_X1 U15119 ( .A1(n12887), .A2(n12879), .ZN(n12880) );
  XNOR2_X1 U15120 ( .A(n12881), .B(n12880), .ZN(n13080) );
  INV_X1 U15121 ( .A(n12882), .ZN(n13147) );
  AOI22_X1 U15122 ( .A1(n12883), .A2(n15150), .B1(n13074), .B2(
        P3_REG2_REG_28__SCAN_IN), .ZN(n12884) );
  OAI21_X1 U15123 ( .B1(n13147), .B2(n14613), .A(n12884), .ZN(n12885) );
  AOI21_X1 U15124 ( .B1(n13080), .B2(n13077), .A(n12885), .ZN(n12886) );
  OAI21_X1 U15125 ( .B1(n13081), .B2(n13074), .A(n12886), .ZN(P3_U3205) );
  OAI22_X1 U15126 ( .A1(n15223), .A2(n13069), .B1(n12926), .B2(n13067), .ZN(
        n12893) );
  XNOR2_X1 U15127 ( .A(n12890), .B(n12889), .ZN(n12891) );
  AOI22_X1 U15128 ( .A1(n12894), .A2(n15150), .B1(n13074), .B2(
        P3_REG2_REG_27__SCAN_IN), .ZN(n12895) );
  OAI21_X1 U15129 ( .B1(n12896), .B2(n14613), .A(n12895), .ZN(n12897) );
  AOI21_X1 U15130 ( .B1(n13085), .B2(n15151), .A(n12897), .ZN(n12898) );
  OAI21_X1 U15131 ( .B1(n13087), .B2(n13074), .A(n12898), .ZN(P3_U3206) );
  NAND2_X1 U15132 ( .A1(n6616), .A2(n12899), .ZN(n12900) );
  NAND2_X1 U15133 ( .A1(n12901), .A2(n12900), .ZN(n13088) );
  XNOR2_X1 U15134 ( .A(n12903), .B(n12902), .ZN(n12904) );
  NAND2_X1 U15135 ( .A1(n12904), .A2(n15143), .ZN(n12908) );
  AOI22_X1 U15136 ( .A1(n12906), .A2(n15136), .B1(n15139), .B2(n12905), .ZN(
        n12907) );
  OAI211_X1 U15137 ( .C1(n15147), .C2(n13088), .A(n12908), .B(n12907), .ZN(
        n13089) );
  NAND2_X1 U15138 ( .A1(n13089), .A2(n15132), .ZN(n12915) );
  INV_X1 U15139 ( .A(n12909), .ZN(n12911) );
  OAI22_X1 U15140 ( .A1(n12911), .A2(n15118), .B1(n15132), .B2(n12910), .ZN(
        n12912) );
  AOI21_X1 U15141 ( .B1(n12913), .B2(n14617), .A(n12912), .ZN(n12914) );
  OAI211_X1 U15142 ( .C1(n12916), .C2(n13088), .A(n12915), .B(n12914), .ZN(
        P3_U3207) );
  NAND2_X1 U15143 ( .A1(n12917), .A2(n12918), .ZN(n12920) );
  XNOR2_X1 U15144 ( .A(n12922), .B(n12921), .ZN(n12929) );
  XNOR2_X1 U15145 ( .A(n12924), .B(n12923), .ZN(n13094) );
  OAI22_X1 U15146 ( .A1(n12926), .A2(n13069), .B1(n12925), .B2(n13067), .ZN(
        n12927) );
  AOI21_X1 U15147 ( .B1(n13094), .B2(n12945), .A(n12927), .ZN(n12928) );
  OAI21_X1 U15148 ( .B1(n12929), .B2(n13064), .A(n12928), .ZN(n13093) );
  INV_X1 U15149 ( .A(n13093), .ZN(n12934) );
  AOI22_X1 U15150 ( .A1(n12930), .A2(n15150), .B1(n13074), .B2(
        P3_REG2_REG_25__SCAN_IN), .ZN(n12931) );
  OAI21_X1 U15151 ( .B1(n13155), .B2(n14613), .A(n12931), .ZN(n12932) );
  AOI21_X1 U15152 ( .B1(n13094), .B2(n15151), .A(n12932), .ZN(n12933) );
  OAI21_X1 U15153 ( .B1(n12934), .B2(n13074), .A(n12933), .ZN(P3_U3208) );
  NAND2_X1 U15154 ( .A1(n12917), .A2(n12935), .ZN(n12936) );
  XNOR2_X1 U15155 ( .A(n12936), .B(n12938), .ZN(n12947) );
  INV_X1 U15156 ( .A(n12937), .ZN(n12940) );
  OAI21_X1 U15157 ( .B1(n12940), .B2(n12939), .A(n12938), .ZN(n12942) );
  NAND2_X1 U15158 ( .A1(n12942), .A2(n12941), .ZN(n13098) );
  OAI22_X1 U15159 ( .A1(n12943), .A2(n13069), .B1(n12975), .B2(n13067), .ZN(
        n12944) );
  AOI21_X1 U15160 ( .B1(n13098), .B2(n12945), .A(n12944), .ZN(n12946) );
  OAI21_X1 U15161 ( .B1(n12947), .B2(n13064), .A(n12946), .ZN(n13097) );
  INV_X1 U15162 ( .A(n13097), .ZN(n12952) );
  AOI22_X1 U15163 ( .A1(n12948), .A2(n15150), .B1(n13074), .B2(
        P3_REG2_REG_24__SCAN_IN), .ZN(n12949) );
  OAI21_X1 U15164 ( .B1(n13159), .B2(n14613), .A(n12949), .ZN(n12950) );
  AOI21_X1 U15165 ( .B1(n13098), .B2(n15151), .A(n12950), .ZN(n12951) );
  OAI21_X1 U15166 ( .B1(n12952), .B2(n13074), .A(n12951), .ZN(P3_U3209) );
  NAND2_X1 U15167 ( .A1(n12954), .A2(n12953), .ZN(n12955) );
  NAND3_X1 U15168 ( .A1(n12917), .A2(n15143), .A3(n12955), .ZN(n12965) );
  AOI22_X1 U15169 ( .A1(n12957), .A2(n15136), .B1(n15139), .B2(n12956), .ZN(
        n12964) );
  NAND2_X1 U15170 ( .A1(n12959), .A2(n12958), .ZN(n12961) );
  NAND2_X1 U15171 ( .A1(n12961), .A2(n12960), .ZN(n12962) );
  NAND2_X1 U15172 ( .A1(n12937), .A2(n12962), .ZN(n12966) );
  OR2_X1 U15173 ( .A1(n12966), .A2(n15147), .ZN(n12963) );
  INV_X1 U15174 ( .A(n12966), .ZN(n13102) );
  AOI22_X1 U15175 ( .A1(n12967), .A2(n15150), .B1(n13074), .B2(
        P3_REG2_REG_23__SCAN_IN), .ZN(n12968) );
  OAI21_X1 U15176 ( .B1(n12969), .B2(n14613), .A(n12968), .ZN(n12970) );
  AOI21_X1 U15177 ( .B1(n13102), .B2(n15151), .A(n12970), .ZN(n12971) );
  OAI21_X1 U15178 ( .B1(n13104), .B2(n13074), .A(n12971), .ZN(P3_U3210) );
  XNOR2_X1 U15179 ( .A(n12972), .B(n12976), .ZN(n12973) );
  OAI222_X1 U15180 ( .A1(n13069), .A2(n12975), .B1(n13067), .B2(n12974), .C1(
        n12973), .C2(n13064), .ZN(n13105) );
  INV_X1 U15181 ( .A(n13105), .ZN(n12982) );
  XOR2_X1 U15182 ( .A(n12977), .B(n12976), .Z(n13106) );
  AOI22_X1 U15183 ( .A1(n12978), .A2(n15150), .B1(n13074), .B2(
        P3_REG2_REG_22__SCAN_IN), .ZN(n12979) );
  OAI21_X1 U15184 ( .B1(n13164), .B2(n14613), .A(n12979), .ZN(n12980) );
  AOI21_X1 U15185 ( .B1(n13106), .B2(n13077), .A(n12980), .ZN(n12981) );
  OAI21_X1 U15186 ( .B1(n12982), .B2(n13074), .A(n12981), .ZN(P3_U3211) );
  XNOR2_X1 U15187 ( .A(n12983), .B(n12986), .ZN(n12984) );
  OAI222_X1 U15188 ( .A1(n13069), .A2(n12985), .B1(n13067), .B2(n13009), .C1(
        n13064), .C2(n12984), .ZN(n13109) );
  INV_X1 U15189 ( .A(n13109), .ZN(n12992) );
  XNOR2_X1 U15190 ( .A(n12987), .B(n12986), .ZN(n13110) );
  AOI22_X1 U15191 ( .A1(n13074), .A2(P3_REG2_REG_21__SCAN_IN), .B1(n12988), 
        .B2(n15150), .ZN(n12989) );
  OAI21_X1 U15192 ( .B1(n13167), .B2(n14613), .A(n12989), .ZN(n12990) );
  AOI21_X1 U15193 ( .B1(n13110), .B2(n13077), .A(n12990), .ZN(n12991) );
  OAI21_X1 U15194 ( .B1(n12992), .B2(n13074), .A(n12991), .ZN(P3_U3212) );
  OAI211_X1 U15195 ( .C1(n12994), .C2(n13004), .A(n12993), .B(n15143), .ZN(
        n12998) );
  AOI22_X1 U15196 ( .A1(n12996), .A2(n15136), .B1(n15139), .B2(n12995), .ZN(
        n12997) );
  NAND2_X1 U15197 ( .A1(n12998), .A2(n12997), .ZN(n13113) );
  AOI21_X1 U15198 ( .B1(n15150), .B2(n12999), .A(n13113), .ZN(n13007) );
  AOI22_X1 U15199 ( .A1(n13000), .A2(n14617), .B1(P3_REG2_REG_20__SCAN_IN), 
        .B2(n13074), .ZN(n13006) );
  INV_X1 U15200 ( .A(n13001), .ZN(n13002) );
  AOI21_X1 U15201 ( .B1(n13004), .B2(n13003), .A(n13002), .ZN(n13114) );
  NAND2_X1 U15202 ( .A1(n13114), .A2(n13077), .ZN(n13005) );
  OAI211_X1 U15203 ( .C1(n13007), .C2(n13074), .A(n13006), .B(n13005), .ZN(
        P3_U3213) );
  AOI21_X1 U15204 ( .B1(n13008), .B2(n13013), .A(n13064), .ZN(n13012) );
  OAI22_X1 U15205 ( .A1(n13009), .A2(n13069), .B1(n13037), .B2(n13067), .ZN(
        n13010) );
  AOI21_X1 U15206 ( .B1(n13012), .B2(n13011), .A(n13010), .ZN(n13119) );
  INV_X1 U15207 ( .A(n13013), .ZN(n13014) );
  XNOR2_X1 U15208 ( .A(n13015), .B(n13014), .ZN(n13117) );
  AOI22_X1 U15209 ( .A1(n13074), .A2(P3_REG2_REG_19__SCAN_IN), .B1(n15150), 
        .B2(n13016), .ZN(n13017) );
  OAI21_X1 U15210 ( .B1(n13175), .B2(n14613), .A(n13017), .ZN(n13018) );
  AOI21_X1 U15211 ( .B1(n13117), .B2(n13077), .A(n13018), .ZN(n13019) );
  OAI21_X1 U15212 ( .B1(n13119), .B2(n13074), .A(n13019), .ZN(P3_U3214) );
  INV_X1 U15213 ( .A(n13020), .ZN(n13021) );
  AOI21_X1 U15214 ( .B1(n13023), .B2(n13022), .A(n13021), .ZN(n13024) );
  OAI222_X1 U15215 ( .A1(n13069), .A2(n13025), .B1(n13067), .B2(n13053), .C1(
        n13064), .C2(n13024), .ZN(n13123) );
  INV_X1 U15216 ( .A(n13123), .ZN(n13035) );
  OAI22_X1 U15217 ( .A1(n15132), .A2(n13027), .B1(n13026), .B2(n15118), .ZN(
        n13028) );
  AOI21_X1 U15218 ( .B1(n13122), .B2(n14617), .A(n13028), .ZN(n13034) );
  NAND2_X1 U15219 ( .A1(n13030), .A2(n13029), .ZN(n13031) );
  AND2_X1 U15220 ( .A1(n13032), .A2(n13031), .ZN(n13124) );
  NAND2_X1 U15221 ( .A1(n13124), .A2(n13077), .ZN(n13033) );
  OAI211_X1 U15222 ( .C1(n13035), .C2(n13074), .A(n13034), .B(n13033), .ZN(
        P3_U3215) );
  AOI21_X1 U15223 ( .B1(n13036), .B2(n13041), .A(n13064), .ZN(n13040) );
  OAI22_X1 U15224 ( .A1(n13068), .A2(n13067), .B1(n13037), .B2(n13069), .ZN(
        n13038) );
  AOI21_X1 U15225 ( .B1(n13040), .B2(n13039), .A(n13038), .ZN(n13129) );
  INV_X1 U15226 ( .A(n13041), .ZN(n13043) );
  NAND3_X1 U15227 ( .A1(n13055), .A2(n13043), .A3(n13042), .ZN(n13044) );
  NAND2_X1 U15228 ( .A1(n13045), .A2(n13044), .ZN(n13127) );
  AOI22_X1 U15229 ( .A1(n13074), .A2(P3_REG2_REG_17__SCAN_IN), .B1(n15150), 
        .B2(n13046), .ZN(n13047) );
  OAI21_X1 U15230 ( .B1(n13048), .B2(n14613), .A(n13047), .ZN(n13049) );
  AOI21_X1 U15231 ( .B1(n13127), .B2(n13077), .A(n13049), .ZN(n13050) );
  OAI21_X1 U15232 ( .B1(n13129), .B2(n13074), .A(n13050), .ZN(P3_U3216) );
  XOR2_X1 U15233 ( .A(n13051), .B(n13056), .Z(n13052) );
  OAI222_X1 U15234 ( .A1(n13067), .A2(n13054), .B1(n13069), .B2(n13053), .C1(
        n13052), .C2(n13064), .ZN(n13130) );
  INV_X1 U15235 ( .A(n13130), .ZN(n13062) );
  OAI21_X1 U15236 ( .B1(n13057), .B2(n13056), .A(n13055), .ZN(n13131) );
  AOI22_X1 U15237 ( .A1(n13074), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n15150), 
        .B2(n13058), .ZN(n13059) );
  OAI21_X1 U15238 ( .B1(n13184), .B2(n14613), .A(n13059), .ZN(n13060) );
  AOI21_X1 U15239 ( .B1(n13131), .B2(n13077), .A(n13060), .ZN(n13061) );
  OAI21_X1 U15240 ( .B1(n13062), .B2(n13074), .A(n13061), .ZN(P3_U3217) );
  XOR2_X1 U15241 ( .A(n13063), .B(n13071), .Z(n13065) );
  OAI222_X1 U15242 ( .A1(n13069), .A2(n13068), .B1(n13067), .B2(n13066), .C1(
        n13065), .C2(n13064), .ZN(n13134) );
  INV_X1 U15243 ( .A(n13134), .ZN(n13079) );
  OAI21_X1 U15244 ( .B1(n13072), .B2(n13071), .A(n13070), .ZN(n13135) );
  AOI22_X1 U15245 ( .A1(n13074), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n15150), 
        .B2(n13073), .ZN(n13075) );
  OAI21_X1 U15246 ( .B1(n13189), .B2(n14613), .A(n13075), .ZN(n13076) );
  AOI21_X1 U15247 ( .B1(n13135), .B2(n13077), .A(n13076), .ZN(n13078) );
  OAI21_X1 U15248 ( .B1(n13079), .B2(n13074), .A(n13078), .ZN(P3_U3218) );
  INV_X1 U15249 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n13082) );
  MUX2_X1 U15250 ( .A(n13082), .B(n13145), .S(n15222), .Z(n13083) );
  INV_X1 U15251 ( .A(n15194), .ZN(n15165) );
  AOI22_X1 U15252 ( .A1(n13085), .A2(n15165), .B1(n14638), .B2(n13084), .ZN(
        n13086) );
  NAND2_X1 U15253 ( .A1(n13087), .A2(n13086), .ZN(n13148) );
  MUX2_X1 U15254 ( .A(P3_REG1_REG_27__SCAN_IN), .B(n13148), .S(n15222), .Z(
        P3_U3486) );
  INV_X1 U15255 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n13091) );
  INV_X1 U15256 ( .A(n13088), .ZN(n13090) );
  AOI21_X1 U15257 ( .B1(n15165), .B2(n13090), .A(n13089), .ZN(n13149) );
  MUX2_X1 U15258 ( .A(n13091), .B(n13149), .S(n15222), .Z(n13092) );
  OAI21_X1 U15259 ( .B1(n13151), .B2(n13138), .A(n13092), .ZN(P3_U3485) );
  INV_X1 U15260 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n13095) );
  AOI21_X1 U15261 ( .B1(n15165), .B2(n13094), .A(n13093), .ZN(n13152) );
  MUX2_X1 U15262 ( .A(n13095), .B(n13152), .S(n15222), .Z(n13096) );
  OAI21_X1 U15263 ( .B1(n13155), .B2(n13138), .A(n13096), .ZN(P3_U3484) );
  INV_X1 U15264 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n13099) );
  AOI21_X1 U15265 ( .B1(n15165), .B2(n13098), .A(n13097), .ZN(n13156) );
  MUX2_X1 U15266 ( .A(n13099), .B(n13156), .S(n15222), .Z(n13100) );
  OAI21_X1 U15267 ( .B1(n13159), .B2(n13138), .A(n13100), .ZN(P3_U3483) );
  AOI22_X1 U15268 ( .A1(n13102), .A2(n15165), .B1(n14638), .B2(n13101), .ZN(
        n13103) );
  NAND2_X1 U15269 ( .A1(n13104), .A2(n13103), .ZN(n13160) );
  MUX2_X1 U15270 ( .A(P3_REG1_REG_23__SCAN_IN), .B(n13160), .S(n15222), .Z(
        P3_U3482) );
  INV_X1 U15271 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n13107) );
  AOI21_X1 U15272 ( .B1(n13139), .B2(n13106), .A(n13105), .ZN(n13161) );
  MUX2_X1 U15273 ( .A(n13107), .B(n13161), .S(n15222), .Z(n13108) );
  OAI21_X1 U15274 ( .B1(n13164), .B2(n13138), .A(n13108), .ZN(P3_U3481) );
  INV_X1 U15275 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n13111) );
  AOI21_X1 U15276 ( .B1(n13110), .B2(n13139), .A(n13109), .ZN(n13165) );
  MUX2_X1 U15277 ( .A(n13111), .B(n13165), .S(n15222), .Z(n13112) );
  OAI21_X1 U15278 ( .B1(n13167), .B2(n13138), .A(n13112), .ZN(P3_U3480) );
  INV_X1 U15279 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n13115) );
  AOI21_X1 U15280 ( .B1(n13114), .B2(n13139), .A(n13113), .ZN(n13168) );
  MUX2_X1 U15281 ( .A(n13115), .B(n13168), .S(n15222), .Z(n13116) );
  OAI21_X1 U15282 ( .B1(n13171), .B2(n13138), .A(n13116), .ZN(P3_U3479) );
  INV_X1 U15283 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n13120) );
  NAND2_X1 U15284 ( .A1(n13117), .A2(n13139), .ZN(n13118) );
  AND2_X1 U15285 ( .A1(n13119), .A2(n13118), .ZN(n13172) );
  MUX2_X1 U15286 ( .A(n13120), .B(n13172), .S(n15222), .Z(n13121) );
  OAI21_X1 U15287 ( .B1(n13138), .B2(n13175), .A(n13121), .ZN(P3_U3478) );
  INV_X1 U15288 ( .A(n13122), .ZN(n13179) );
  INV_X1 U15289 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n15492) );
  AOI21_X1 U15290 ( .B1(n13124), .B2(n13139), .A(n13123), .ZN(n13176) );
  MUX2_X1 U15291 ( .A(n15492), .B(n13176), .S(n15222), .Z(n13125) );
  OAI21_X1 U15292 ( .B1(n13179), .B2(n13138), .A(n13125), .ZN(P3_U3477) );
  AOI22_X1 U15293 ( .A1(n13127), .A2(n13139), .B1(n14638), .B2(n13126), .ZN(
        n13128) );
  NAND2_X1 U15294 ( .A1(n13129), .A2(n13128), .ZN(n13180) );
  MUX2_X1 U15295 ( .A(P3_REG1_REG_17__SCAN_IN), .B(n13180), .S(n15222), .Z(
        P3_U3476) );
  AOI21_X1 U15296 ( .B1(n13139), .B2(n13131), .A(n13130), .ZN(n13181) );
  MUX2_X1 U15297 ( .A(n13132), .B(n13181), .S(n15222), .Z(n13133) );
  OAI21_X1 U15298 ( .B1(n13184), .B2(n13138), .A(n13133), .ZN(P3_U3475) );
  INV_X1 U15299 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n13136) );
  AOI21_X1 U15300 ( .B1(n13139), .B2(n13135), .A(n13134), .ZN(n13185) );
  MUX2_X1 U15301 ( .A(n13136), .B(n13185), .S(n15222), .Z(n13137) );
  OAI21_X1 U15302 ( .B1(n13189), .B2(n13138), .A(n13137), .ZN(P3_U3474) );
  INV_X1 U15303 ( .A(n13139), .ZN(n15201) );
  NAND2_X1 U15304 ( .A1(n13140), .A2(n14638), .ZN(n13141) );
  OAI211_X1 U15305 ( .C1(n15201), .C2(n13143), .A(n13142), .B(n13141), .ZN(
        n13190) );
  MUX2_X1 U15306 ( .A(P3_REG1_REG_14__SCAN_IN), .B(n13190), .S(n15222), .Z(
        P3_U3473) );
  INV_X1 U15307 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n13144) );
  MUX2_X1 U15308 ( .A(n13145), .B(n13144), .S(n15206), .Z(n13146) );
  INV_X2 U15309 ( .A(n15206), .ZN(n15205) );
  MUX2_X1 U15310 ( .A(P3_REG0_REG_27__SCAN_IN), .B(n13148), .S(n15205), .Z(
        P3_U3454) );
  INV_X1 U15311 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n15452) );
  MUX2_X1 U15312 ( .A(n15452), .B(n13149), .S(n15205), .Z(n13150) );
  OAI21_X1 U15313 ( .B1(n13151), .B2(n13188), .A(n13150), .ZN(P3_U3453) );
  INV_X1 U15314 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n13153) );
  MUX2_X1 U15315 ( .A(n13153), .B(n13152), .S(n15205), .Z(n13154) );
  OAI21_X1 U15316 ( .B1(n13155), .B2(n13188), .A(n13154), .ZN(P3_U3452) );
  INV_X1 U15317 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n13157) );
  MUX2_X1 U15318 ( .A(n13157), .B(n13156), .S(n15205), .Z(n13158) );
  OAI21_X1 U15319 ( .B1(n13159), .B2(n13188), .A(n13158), .ZN(P3_U3451) );
  MUX2_X1 U15320 ( .A(n13160), .B(P3_REG0_REG_23__SCAN_IN), .S(n15206), .Z(
        P3_U3450) );
  INV_X1 U15321 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n13162) );
  MUX2_X1 U15322 ( .A(n13162), .B(n13161), .S(n15205), .Z(n13163) );
  OAI21_X1 U15323 ( .B1(n13164), .B2(n13188), .A(n13163), .ZN(P3_U3449) );
  INV_X1 U15324 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n15284) );
  MUX2_X1 U15325 ( .A(n15284), .B(n13165), .S(n15205), .Z(n13166) );
  OAI21_X1 U15326 ( .B1(n13167), .B2(n13188), .A(n13166), .ZN(P3_U3448) );
  INV_X1 U15327 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n13169) );
  MUX2_X1 U15328 ( .A(n13169), .B(n13168), .S(n15205), .Z(n13170) );
  OAI21_X1 U15329 ( .B1(n13171), .B2(n13188), .A(n13170), .ZN(P3_U3447) );
  MUX2_X1 U15330 ( .A(n13173), .B(n13172), .S(n15205), .Z(n13174) );
  OAI21_X1 U15331 ( .B1(n13188), .B2(n13175), .A(n13174), .ZN(P3_U3446) );
  INV_X1 U15332 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n13177) );
  MUX2_X1 U15333 ( .A(n13177), .B(n13176), .S(n15205), .Z(n13178) );
  OAI21_X1 U15334 ( .B1(n13179), .B2(n13188), .A(n13178), .ZN(P3_U3444) );
  MUX2_X1 U15335 ( .A(P3_REG0_REG_17__SCAN_IN), .B(n13180), .S(n15205), .Z(
        P3_U3441) );
  INV_X1 U15336 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n13182) );
  MUX2_X1 U15337 ( .A(n13182), .B(n13181), .S(n15205), .Z(n13183) );
  OAI21_X1 U15338 ( .B1(n13184), .B2(n13188), .A(n13183), .ZN(P3_U3438) );
  INV_X1 U15339 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n13186) );
  MUX2_X1 U15340 ( .A(n13186), .B(n13185), .S(n15205), .Z(n13187) );
  OAI21_X1 U15341 ( .B1(n13189), .B2(n13188), .A(n13187), .ZN(P3_U3435) );
  MUX2_X1 U15342 ( .A(P3_REG0_REG_14__SCAN_IN), .B(n13190), .S(n15205), .Z(
        P3_U3432) );
  MUX2_X1 U15343 ( .A(n13192), .B(P3_D_REG_1__SCAN_IN), .S(n13191), .Z(
        P3_U3377) );
  MUX2_X1 U15344 ( .A(P3_D_REG_0__SCAN_IN), .B(n7329), .S(n13193), .Z(P3_U3376) );
  INV_X1 U15345 ( .A(n13194), .ZN(n13199) );
  NOR4_X1 U15346 ( .A1(n13196), .A2(P3_IR_REG_30__SCAN_IN), .A3(n13195), .A4(
        P3_U3151), .ZN(n13197) );
  AOI21_X1 U15347 ( .B1(n13200), .B2(SI_31_), .A(n13197), .ZN(n13198) );
  OAI21_X1 U15348 ( .B1(n13199), .B2(n13213), .A(n13198), .ZN(P3_U3264) );
  AOI22_X1 U15349 ( .A1(n13202), .A2(n13201), .B1(n13200), .B2(SI_29_), .ZN(
        n13203) );
  OAI21_X1 U15350 ( .B1(n8529), .B2(P3_U3151), .A(n13203), .ZN(P3_U3266) );
  INV_X1 U15351 ( .A(n13204), .ZN(n13207) );
  OAI222_X1 U15352 ( .A1(n13213), .A2(n13207), .B1(n13217), .B2(n13206), .C1(
        P3_U3151), .C2(n13205), .ZN(P3_U3267) );
  INV_X1 U15353 ( .A(n13208), .ZN(n13212) );
  INV_X1 U15354 ( .A(SI_27_), .ZN(n13211) );
  OAI222_X1 U15355 ( .A1(n13213), .A2(n13212), .B1(n13217), .B2(n13211), .C1(
        P3_U3151), .C2(n13209), .ZN(P3_U3268) );
  INV_X1 U15356 ( .A(n13214), .ZN(n13215) );
  OAI222_X1 U15357 ( .A1(P3_U3151), .A2(n13218), .B1(n13217), .B2(n13216), 
        .C1(n13213), .C2(n13215), .ZN(P3_U3269) );
  MUX2_X1 U15358 ( .A(n13219), .B(n15507), .S(P3_STATE_REG_SCAN_IN), .Z(
        P3_U3295) );
  XNOR2_X1 U15359 ( .A(n13708), .B(n13236), .ZN(n13224) );
  NAND2_X1 U15360 ( .A1(n13625), .A2(n10574), .ZN(n13225) );
  NAND2_X1 U15361 ( .A1(n13224), .A2(n13225), .ZN(n13229) );
  INV_X1 U15362 ( .A(n13224), .ZN(n13227) );
  INV_X1 U15363 ( .A(n13225), .ZN(n13226) );
  NAND2_X1 U15364 ( .A1(n13227), .A2(n13226), .ZN(n13228) );
  NAND2_X1 U15365 ( .A1(n13229), .A2(n13228), .ZN(n13271) );
  NAND2_X1 U15366 ( .A1(n13269), .A2(n13229), .ZN(n13313) );
  XNOR2_X1 U15367 ( .A(n13703), .B(n13236), .ZN(n13230) );
  NAND2_X1 U15368 ( .A1(n13356), .A2(n10574), .ZN(n13231) );
  NAND2_X1 U15369 ( .A1(n13230), .A2(n13231), .ZN(n13235) );
  INV_X1 U15370 ( .A(n13230), .ZN(n13233) );
  INV_X1 U15371 ( .A(n13231), .ZN(n13232) );
  NAND2_X1 U15372 ( .A1(n13233), .A2(n13232), .ZN(n13234) );
  AND2_X1 U15373 ( .A1(n13235), .A2(n13234), .ZN(n13314) );
  XNOR2_X1 U15374 ( .A(n13755), .B(n13236), .ZN(n13238) );
  NOR2_X1 U15375 ( .A1(n13550), .A2(n13603), .ZN(n13237) );
  XNOR2_X1 U15376 ( .A(n13238), .B(n13237), .ZN(n13289) );
  NAND2_X1 U15377 ( .A1(n13238), .A2(n13237), .ZN(n13239) );
  XOR2_X1 U15378 ( .A(n13282), .B(n13690), .Z(n13240) );
  XNOR2_X1 U15379 ( .A(n13242), .B(n13240), .ZN(n13323) );
  NAND2_X1 U15380 ( .A1(n10574), .A2(n13532), .ZN(n13325) );
  INV_X1 U15381 ( .A(n13240), .ZN(n13241) );
  OR2_X1 U15382 ( .A1(n13242), .A2(n13241), .ZN(n13243) );
  NOR2_X1 U15383 ( .A1(n13603), .A2(n13549), .ZN(n13261) );
  INV_X1 U15384 ( .A(n13244), .ZN(n13245) );
  AOI22_X2 U15385 ( .A1(n13262), .A2(n13261), .B1(n13245), .B2(n6649), .ZN(
        n13306) );
  NAND2_X1 U15386 ( .A1(n10574), .A2(n13533), .ZN(n13247) );
  XNOR2_X1 U15387 ( .A(n13681), .B(n13282), .ZN(n13246) );
  XOR2_X1 U15388 ( .A(n13247), .B(n13246), .Z(n13305) );
  INV_X1 U15389 ( .A(n13246), .ZN(n13248) );
  XNOR2_X1 U15390 ( .A(n13503), .B(n13282), .ZN(n13250) );
  NAND2_X1 U15391 ( .A1(n10574), .A2(n13353), .ZN(n13249) );
  XNOR2_X1 U15392 ( .A(n13250), .B(n13249), .ZN(n13296) );
  INV_X1 U15393 ( .A(n13249), .ZN(n13251) );
  AND2_X1 U15394 ( .A1(n10574), .A2(n13495), .ZN(n13253) );
  XNOR2_X1 U15395 ( .A(n13670), .B(n13282), .ZN(n13252) );
  NOR2_X1 U15396 ( .A1(n13252), .A2(n13253), .ZN(n13254) );
  AOI21_X1 U15397 ( .B1(n13253), .B2(n13252), .A(n13254), .ZN(n13337) );
  INV_X1 U15398 ( .A(n13254), .ZN(n13255) );
  NAND2_X1 U15399 ( .A1(n10574), .A2(n13352), .ZN(n13278) );
  XNOR2_X1 U15400 ( .A(n13661), .B(n13282), .ZN(n13277) );
  XNOR2_X1 U15401 ( .A(n13280), .B(n13279), .ZN(n13260) );
  INV_X1 U15402 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n13256) );
  OAI22_X1 U15403 ( .A1(n13328), .A2(n13300), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13256), .ZN(n13258) );
  OAI22_X1 U15404 ( .A1(n13329), .A2(n7188), .B1(n13344), .B2(n13466), .ZN(
        n13257) );
  AOI211_X1 U15405 ( .C1(n13661), .C2(n13346), .A(n13258), .B(n13257), .ZN(
        n13259) );
  OAI21_X1 U15406 ( .B1(n13260), .B2(n13348), .A(n13259), .ZN(P2_U3186) );
  XNOR2_X1 U15407 ( .A(n13262), .B(n13261), .ZN(n13268) );
  OAI22_X1 U15408 ( .A1(n13328), .A2(n13264), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13263), .ZN(n13266) );
  OAI22_X1 U15409 ( .A1(n13329), .A2(n13299), .B1(n13344), .B2(n13536), .ZN(
        n13265) );
  AOI211_X1 U15410 ( .C1(n13686), .C2(n13346), .A(n13266), .B(n13265), .ZN(
        n13267) );
  OAI21_X1 U15411 ( .B1(n13268), .B2(n13348), .A(n13267), .ZN(P2_U3188) );
  INV_X1 U15412 ( .A(n13269), .ZN(n13270) );
  AOI21_X1 U15413 ( .B1(n13272), .B2(n13271), .A(n13270), .ZN(n13276) );
  NOR2_X1 U15414 ( .A1(n13344), .A2(n13607), .ZN(n13274) );
  AOI22_X1 U15415 ( .A1(n13356), .A2(n13496), .B1(n13462), .B2(n13357), .ZN(
        n13599) );
  NAND2_X1 U15416 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n13413)
         );
  OAI21_X1 U15417 ( .B1(n13318), .B2(n13599), .A(n13413), .ZN(n13273) );
  AOI211_X1 U15418 ( .C1(n13708), .C2(n13346), .A(n13274), .B(n13273), .ZN(
        n13275) );
  OAI21_X1 U15419 ( .B1(n13276), .B2(n13348), .A(n13275), .ZN(P2_U3191) );
  NAND2_X1 U15420 ( .A1(n10574), .A2(n13463), .ZN(n13281) );
  XNOR2_X1 U15421 ( .A(n13282), .B(n13281), .ZN(n13283) );
  AOI22_X1 U15422 ( .A1(n13342), .A2(n13284), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13285) );
  OAI21_X1 U15423 ( .B1(n13451), .B2(n13344), .A(n13285), .ZN(n13286) );
  AOI21_X1 U15424 ( .B1(n13287), .B2(n13346), .A(n13286), .ZN(n13288) );
  XNOR2_X1 U15425 ( .A(n13290), .B(n13289), .ZN(n13295) );
  AOI22_X1 U15426 ( .A1(n13356), .A2(n13462), .B1(n13496), .B2(n13532), .ZN(
        n13567) );
  INV_X1 U15427 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n13291) );
  OAI22_X1 U15428 ( .A1(n13318), .A2(n13567), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13291), .ZN(n13293) );
  NOR2_X1 U15429 ( .A1(n13755), .A2(n13334), .ZN(n13292) );
  AOI211_X1 U15430 ( .C1(n13320), .C2(n13575), .A(n13293), .B(n13292), .ZN(
        n13294) );
  OAI21_X1 U15431 ( .B1(n13295), .B2(n13348), .A(n13294), .ZN(P2_U3195) );
  XNOR2_X1 U15432 ( .A(n13297), .B(n13296), .ZN(n13304) );
  OAI22_X1 U15433 ( .A1(n13328), .A2(n13299), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13298), .ZN(n13302) );
  OAI22_X1 U15434 ( .A1(n13329), .A2(n13300), .B1(n13344), .B2(n13501), .ZN(
        n13301) );
  AOI211_X1 U15435 ( .C1(n13503), .C2(n13346), .A(n13302), .B(n13301), .ZN(
        n13303) );
  OAI21_X1 U15436 ( .B1(n13304), .B2(n13348), .A(n13303), .ZN(P2_U3197) );
  XNOR2_X1 U15437 ( .A(n13306), .B(n13305), .ZN(n13311) );
  NOR2_X1 U15438 ( .A1(n13344), .A2(n13521), .ZN(n13309) );
  AOI22_X1 U15439 ( .A1(n13354), .A2(n13462), .B1(n13496), .B2(n13353), .ZN(
        n13515) );
  INV_X1 U15440 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n13307) );
  OAI22_X1 U15441 ( .A1(n13318), .A2(n13515), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13307), .ZN(n13308) );
  AOI211_X1 U15442 ( .C1(n13681), .C2(n13346), .A(n13309), .B(n13308), .ZN(
        n13310) );
  OAI21_X1 U15443 ( .B1(n13311), .B2(n13348), .A(n13310), .ZN(P2_U3201) );
  OAI21_X1 U15444 ( .B1(n13314), .B2(n13313), .A(n13312), .ZN(n13315) );
  NAND2_X1 U15445 ( .A1(n13315), .A2(n13326), .ZN(n13322) );
  INV_X1 U15446 ( .A(n13316), .ZN(n13589) );
  AOI22_X1 U15447 ( .A1(n13355), .A2(n13496), .B1(n13462), .B2(n13625), .ZN(
        n13586) );
  OAI22_X1 U15448 ( .A1(n13586), .A2(n13318), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13317), .ZN(n13319) );
  AOI21_X1 U15449 ( .B1(n13589), .B2(n13320), .A(n13319), .ZN(n13321) );
  OAI211_X1 U15450 ( .C1(n13591), .C2(n13334), .A(n13322), .B(n13321), .ZN(
        P2_U3205) );
  INV_X1 U15451 ( .A(n13690), .ZN(n13335) );
  OAI21_X1 U15452 ( .B1(n13323), .B2(n13325), .A(n13324), .ZN(n13327) );
  NAND2_X1 U15453 ( .A1(n13327), .A2(n13326), .ZN(n13333) );
  NOR2_X1 U15454 ( .A1(n13328), .A2(n13550), .ZN(n13331) );
  OAI22_X1 U15455 ( .A1(n13329), .A2(n13549), .B1(n13344), .B2(n13556), .ZN(
        n13330) );
  AOI211_X1 U15456 ( .C1(P2_REG3_REG_22__SCAN_IN), .C2(P2_U3088), .A(n13331), 
        .B(n13330), .ZN(n13332) );
  OAI211_X1 U15457 ( .C1(n13335), .C2(n13334), .A(n13333), .B(n13332), .ZN(
        P2_U3207) );
  OAI21_X1 U15458 ( .B1(n13338), .B2(n13337), .A(n13336), .ZN(n13339) );
  INV_X1 U15459 ( .A(n13339), .ZN(n13349) );
  NAND2_X1 U15460 ( .A1(n13462), .A2(n13353), .ZN(n13341) );
  NAND2_X1 U15461 ( .A1(n13496), .A2(n13352), .ZN(n13340) );
  NAND2_X1 U15462 ( .A1(n13341), .A2(n13340), .ZN(n13477) );
  AOI22_X1 U15463 ( .A1(n13342), .A2(n13477), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13343) );
  OAI21_X1 U15464 ( .B1(n13482), .B2(n13344), .A(n13343), .ZN(n13345) );
  AOI21_X1 U15465 ( .B1(n13670), .B2(n13346), .A(n13345), .ZN(n13347) );
  OAI21_X1 U15466 ( .B1(n13349), .B2(n13348), .A(n13347), .ZN(P2_U3212) );
  MUX2_X1 U15467 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n13420), .S(n6550), .Z(
        P2_U3562) );
  MUX2_X1 U15468 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n13350), .S(n6550), .Z(
        P2_U3561) );
  MUX2_X1 U15469 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n13351), .S(n6550), .Z(
        P2_U3560) );
  MUX2_X1 U15470 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n13463), .S(n6550), .Z(
        P2_U3559) );
  MUX2_X1 U15471 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n13352), .S(n6550), .Z(
        P2_U3558) );
  MUX2_X1 U15472 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n13495), .S(n6550), .Z(
        P2_U3557) );
  MUX2_X1 U15473 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n13353), .S(n6550), .Z(
        P2_U3556) );
  MUX2_X1 U15474 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n13533), .S(n6550), .Z(
        P2_U3555) );
  MUX2_X1 U15475 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n13354), .S(n6550), .Z(
        P2_U3554) );
  MUX2_X1 U15476 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n13532), .S(n6550), .Z(
        P2_U3553) );
  MUX2_X1 U15477 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n13355), .S(n6550), .Z(
        P2_U3552) );
  MUX2_X1 U15478 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n13356), .S(n6550), .Z(
        P2_U3551) );
  MUX2_X1 U15479 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n13625), .S(n6550), .Z(
        P2_U3550) );
  MUX2_X1 U15480 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n13357), .S(n6550), .Z(
        P2_U3549) );
  MUX2_X1 U15481 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n13358), .S(n6550), .Z(
        P2_U3548) );
  MUX2_X1 U15482 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n13359), .S(n6550), .Z(
        P2_U3547) );
  MUX2_X1 U15483 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n13360), .S(n6550), .Z(
        P2_U3546) );
  MUX2_X1 U15484 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n13361), .S(n6550), .Z(
        P2_U3545) );
  MUX2_X1 U15485 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n13362), .S(n6550), .Z(
        P2_U3544) );
  MUX2_X1 U15486 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n13363), .S(n6550), .Z(
        P2_U3543) );
  MUX2_X1 U15487 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n13364), .S(n6550), .Z(
        P2_U3542) );
  MUX2_X1 U15488 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n13365), .S(n6550), .Z(
        P2_U3541) );
  MUX2_X1 U15489 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n13366), .S(n6550), .Z(
        P2_U3540) );
  MUX2_X1 U15490 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n13367), .S(n6550), .Z(
        P2_U3539) );
  MUX2_X1 U15491 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n13368), .S(n6550), .Z(
        P2_U3538) );
  MUX2_X1 U15492 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n13369), .S(n6550), .Z(
        P2_U3537) );
  MUX2_X1 U15493 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n13370), .S(n6550), .Z(
        P2_U3536) );
  MUX2_X1 U15494 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n13371), .S(n6550), .Z(
        P2_U3535) );
  MUX2_X1 U15495 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n13372), .S(n6550), .Z(
        P2_U3534) );
  MUX2_X1 U15496 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n13373), .S(n6550), .Z(
        P2_U3533) );
  MUX2_X1 U15497 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n13374), .S(n6550), .Z(
        P2_U3532) );
  MUX2_X1 U15498 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n13375), .S(n6550), .Z(
        P2_U3531) );
  NAND2_X1 U15499 ( .A1(n14914), .A2(n13376), .ZN(n13379) );
  INV_X1 U15500 ( .A(n13377), .ZN(n13378) );
  OAI211_X1 U15501 ( .C1(n7282), .C2(n14932), .A(n13379), .B(n13378), .ZN(
        n13380) );
  INV_X1 U15502 ( .A(n13380), .ZN(n13389) );
  OAI211_X1 U15503 ( .C1(n13383), .C2(n13382), .A(n14929), .B(n13381), .ZN(
        n13388) );
  OAI211_X1 U15504 ( .C1(n13386), .C2(n13385), .A(n14846), .B(n13384), .ZN(
        n13387) );
  NAND3_X1 U15505 ( .A1(n13389), .A2(n13388), .A3(n13387), .ZN(P2_U3221) );
  NOR2_X1 U15506 ( .A1(n14913), .A2(n13390), .ZN(n13391) );
  AOI21_X1 U15507 ( .B1(n14913), .B2(n13390), .A(n13391), .ZN(n14910) );
  NOR2_X1 U15508 ( .A1(n13394), .A2(n13404), .ZN(n13395) );
  XNOR2_X1 U15509 ( .A(n13404), .B(n13394), .ZN(n14882) );
  NOR2_X1 U15510 ( .A1(n9357), .A2(n14882), .ZN(n14881) );
  NOR2_X1 U15511 ( .A1(n13395), .A2(n14881), .ZN(n14894) );
  NAND2_X1 U15512 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n14900), .ZN(n13396) );
  OAI21_X1 U15513 ( .B1(n14900), .B2(P2_REG2_REG_16__SCAN_IN), .A(n13396), 
        .ZN(n14893) );
  NOR2_X1 U15514 ( .A1(n14894), .A2(n14893), .ZN(n14892) );
  NAND2_X1 U15515 ( .A1(n14919), .A2(n9395), .ZN(n14918) );
  NAND2_X1 U15516 ( .A1(n13398), .A2(n14920), .ZN(n13399) );
  NAND2_X1 U15517 ( .A1(n14918), .A2(n13399), .ZN(n13400) );
  XNOR2_X1 U15518 ( .A(n13400), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n13409) );
  XNOR2_X1 U15519 ( .A(n14913), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n14905) );
  AOI21_X1 U15520 ( .B1(n13402), .B2(P2_REG1_REG_14__SCAN_IN), .A(n13401), 
        .ZN(n13403) );
  NOR2_X1 U15521 ( .A1(n13403), .A2(n13404), .ZN(n13405) );
  XNOR2_X1 U15522 ( .A(n13404), .B(n13403), .ZN(n14885) );
  NOR2_X1 U15523 ( .A1(n14884), .A2(n14885), .ZN(n14883) );
  NOR2_X1 U15524 ( .A1(n13405), .A2(n14883), .ZN(n14897) );
  XNOR2_X1 U15525 ( .A(n14900), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n14896) );
  NOR2_X1 U15526 ( .A1(n14897), .A2(n14896), .ZN(n14895) );
  AOI21_X1 U15527 ( .B1(n14900), .B2(P2_REG1_REG_16__SCAN_IN), .A(n14895), 
        .ZN(n14906) );
  NOR2_X1 U15528 ( .A1(n14905), .A2(n14906), .ZN(n14904) );
  AOI21_X1 U15529 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(n14913), .A(n14904), 
        .ZN(n13406) );
  NOR2_X1 U15530 ( .A1(n13406), .A2(n14920), .ZN(n13407) );
  XNOR2_X1 U15531 ( .A(n13406), .B(n14920), .ZN(n14925) );
  NOR2_X1 U15532 ( .A1(n14924), .A2(n14925), .ZN(n14923) );
  NOR2_X1 U15533 ( .A1(n13407), .A2(n14923), .ZN(n13408) );
  XNOR2_X1 U15534 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n13408), .ZN(n13411) );
  AOI22_X1 U15535 ( .A1(n13409), .A2(n14929), .B1(n14846), .B2(n13411), .ZN(
        n13412) );
  INV_X1 U15536 ( .A(n13409), .ZN(n13410) );
  OAI211_X1 U15537 ( .C1(n13415), .C2(n14932), .A(n13414), .B(n13413), .ZN(
        P2_U3233) );
  XNOR2_X1 U15538 ( .A(n12166), .B(n13424), .ZN(n13416) );
  OR2_X1 U15539 ( .A1(n13416), .A2(n10574), .ZN(n13641) );
  INV_X1 U15540 ( .A(P2_B_REG_SCAN_IN), .ZN(n13417) );
  OR2_X1 U15541 ( .A1(n13418), .A2(n13417), .ZN(n13419) );
  NAND2_X1 U15542 ( .A1(n13496), .A2(n13419), .ZN(n13437) );
  INV_X1 U15543 ( .A(n13420), .ZN(n13421) );
  OR2_X1 U15544 ( .A1(n13437), .A2(n13421), .ZN(n13644) );
  NOR2_X1 U15545 ( .A1(n14947), .A2(n13644), .ZN(n13427) );
  NOR2_X1 U15546 ( .A1(n12165), .A2(n13610), .ZN(n13422) );
  AOI211_X1 U15547 ( .C1(n14947), .C2(P2_REG2_REG_31__SCAN_IN), .A(n13427), 
        .B(n13422), .ZN(n13423) );
  OAI21_X1 U15548 ( .B1(n13641), .B2(n14939), .A(n13423), .ZN(P2_U3234) );
  INV_X1 U15549 ( .A(n13426), .ZN(n13739) );
  INV_X1 U15550 ( .A(n13424), .ZN(n13425) );
  AOI211_X1 U15551 ( .C1(n13426), .C2(n13442), .A(n10574), .B(n13425), .ZN(
        n13646) );
  NAND2_X1 U15552 ( .A1(n13646), .A2(n13613), .ZN(n13429) );
  AOI21_X1 U15553 ( .B1(n14947), .B2(P2_REG2_REG_30__SCAN_IN), .A(n13427), 
        .ZN(n13428) );
  OAI211_X1 U15554 ( .C1(n13739), .C2(n13610), .A(n13429), .B(n13428), .ZN(
        P2_U3235) );
  XNOR2_X1 U15555 ( .A(n13435), .B(n13434), .ZN(n13440) );
  OAI22_X1 U15556 ( .A1(n7188), .A2(n13627), .B1(n13437), .B2(n13436), .ZN(
        n13438) );
  INV_X1 U15557 ( .A(n13438), .ZN(n13439) );
  OAI21_X1 U15558 ( .B1(n13440), .B2(n13600), .A(n13439), .ZN(n13648) );
  AOI21_X1 U15559 ( .B1(n13650), .B2(n13441), .A(n10574), .ZN(n13443) );
  NAND2_X1 U15560 ( .A1(n13649), .A2(n13613), .ZN(n13447) );
  INV_X1 U15561 ( .A(n13444), .ZN(n13445) );
  AOI22_X1 U15562 ( .A1(n14947), .A2(P2_REG2_REG_29__SCAN_IN), .B1(n14936), 
        .B2(n13445), .ZN(n13446) );
  OAI211_X1 U15563 ( .C1(n6975), .C2(n13610), .A(n13447), .B(n13446), .ZN(
        n13448) );
  AOI21_X1 U15564 ( .B1(n13648), .B2(n13602), .A(n13448), .ZN(n13449) );
  OAI21_X1 U15565 ( .B1(n13653), .B2(n14942), .A(n13449), .ZN(P2_U3236) );
  OAI21_X1 U15566 ( .B1(n13451), .B2(n13535), .A(n13450), .ZN(n13452) );
  NAND2_X1 U15567 ( .A1(n13452), .A2(n13602), .ZN(n13458) );
  INV_X1 U15568 ( .A(n13453), .ZN(n13456) );
  OAI22_X1 U15569 ( .A1(n13658), .A2(n13610), .B1(n13602), .B2(n13454), .ZN(
        n13455) );
  AOI21_X1 U15570 ( .B1(n13456), .B2(n13613), .A(n13455), .ZN(n13457) );
  OAI211_X1 U15571 ( .C1(n14942), .C2(n13459), .A(n13458), .B(n13457), .ZN(
        P2_U3237) );
  XNOR2_X1 U15572 ( .A(n13460), .B(n13471), .ZN(n13461) );
  NAND2_X1 U15573 ( .A1(n13461), .A2(n13618), .ZN(n13465) );
  AOI22_X1 U15574 ( .A1(n13496), .A2(n13463), .B1(n13462), .B2(n13495), .ZN(
        n13464) );
  NAND2_X1 U15575 ( .A1(n13465), .A2(n13464), .ZN(n13666) );
  INV_X1 U15576 ( .A(n13666), .ZN(n13475) );
  OAI22_X1 U15577 ( .A1(n13602), .A2(n13467), .B1(n13466), .B2(n13535), .ZN(
        n13470) );
  AND2_X1 U15578 ( .A1(n13661), .A2(n13480), .ZN(n13468) );
  OR3_X1 U15579 ( .A1(n13468), .A2(n6582), .A3(n10574), .ZN(n13662) );
  NOR2_X1 U15580 ( .A1(n13662), .A2(n14939), .ZN(n13469) );
  AOI211_X1 U15581 ( .C1(n14935), .C2(n13661), .A(n13470), .B(n13469), .ZN(
        n13474) );
  NAND2_X1 U15582 ( .A1(n13472), .A2(n13471), .ZN(n13659) );
  NAND3_X1 U15583 ( .A1(n13660), .A2(n13659), .A3(n13579), .ZN(n13473) );
  OAI211_X1 U15584 ( .C1(n13475), .C2(n14947), .A(n13474), .B(n13473), .ZN(
        P2_U3238) );
  XOR2_X1 U15585 ( .A(n13476), .B(n13486), .Z(n13478) );
  AOI21_X1 U15586 ( .B1(n13478), .B2(n13618), .A(n13477), .ZN(n13672) );
  INV_X1 U15587 ( .A(n13480), .ZN(n13481) );
  AOI211_X1 U15588 ( .C1(n13670), .C2(n13499), .A(n10574), .B(n13481), .ZN(
        n13669) );
  INV_X1 U15589 ( .A(n13670), .ZN(n13485) );
  INV_X1 U15590 ( .A(n13482), .ZN(n13483) );
  AOI22_X1 U15591 ( .A1(n14947), .A2(P2_REG2_REG_26__SCAN_IN), .B1(n14936), 
        .B2(n13483), .ZN(n13484) );
  OAI21_X1 U15592 ( .B1(n13485), .B2(n13610), .A(n13484), .ZN(n13489) );
  XNOR2_X1 U15593 ( .A(n13487), .B(n13486), .ZN(n13673) );
  NOR2_X1 U15594 ( .A1(n13673), .A2(n14942), .ZN(n13488) );
  AOI211_X1 U15595 ( .C1(n13669), .C2(n13613), .A(n13489), .B(n13488), .ZN(
        n13490) );
  OAI21_X1 U15596 ( .B1(n14947), .B2(n13672), .A(n13490), .ZN(P2_U3239) );
  XNOR2_X1 U15597 ( .A(n13491), .B(n13493), .ZN(n13674) );
  INV_X1 U15598 ( .A(n13674), .ZN(n13508) );
  XNOR2_X1 U15599 ( .A(n13492), .B(n13493), .ZN(n13494) );
  NAND2_X1 U15600 ( .A1(n13494), .A2(n13618), .ZN(n13498) );
  AOI22_X1 U15601 ( .A1(n13462), .A2(n13533), .B1(n13496), .B2(n13495), .ZN(
        n13497) );
  NAND2_X1 U15602 ( .A1(n13498), .A2(n13497), .ZN(n13676) );
  NAND2_X1 U15603 ( .A1(n13676), .A2(n13602), .ZN(n13507) );
  AOI21_X1 U15604 ( .B1(n13503), .B2(n13518), .A(n10574), .ZN(n13500) );
  AND2_X1 U15605 ( .A1(n13500), .A2(n13499), .ZN(n13675) );
  OAI22_X1 U15606 ( .A1(n13602), .A2(n13502), .B1(n13501), .B2(n13535), .ZN(
        n13505) );
  INV_X1 U15607 ( .A(n13503), .ZN(n13748) );
  NOR2_X1 U15608 ( .A1(n13748), .A2(n13610), .ZN(n13504) );
  AOI211_X1 U15609 ( .C1(n13675), .C2(n13613), .A(n13505), .B(n13504), .ZN(
        n13506) );
  OAI211_X1 U15610 ( .C1(n13508), .C2(n14942), .A(n13507), .B(n13506), .ZN(
        P2_U3240) );
  XNOR2_X1 U15611 ( .A(n13510), .B(n13509), .ZN(n13517) );
  OR2_X1 U15612 ( .A1(n13512), .A2(n13511), .ZN(n13513) );
  NAND2_X1 U15613 ( .A1(n13514), .A2(n13513), .ZN(n13684) );
  OAI21_X1 U15614 ( .B1(n13684), .B2(n13624), .A(n13515), .ZN(n13516) );
  AOI21_X1 U15615 ( .B1(n13618), .B2(n13517), .A(n13516), .ZN(n13683) );
  INV_X1 U15616 ( .A(n13518), .ZN(n13519) );
  AOI211_X1 U15617 ( .C1(n13681), .C2(n13538), .A(n10574), .B(n13519), .ZN(
        n13680) );
  INV_X1 U15618 ( .A(n13681), .ZN(n13520) );
  NOR2_X1 U15619 ( .A1(n13520), .A2(n13610), .ZN(n13524) );
  OAI22_X1 U15620 ( .A1(n13602), .A2(n13522), .B1(n13521), .B2(n13535), .ZN(
        n13523) );
  AOI211_X1 U15621 ( .C1(n13680), .C2(n13613), .A(n13524), .B(n13523), .ZN(
        n13527) );
  INV_X1 U15622 ( .A(n13684), .ZN(n13525) );
  NAND2_X1 U15623 ( .A1(n13525), .A2(n13638), .ZN(n13526) );
  OAI211_X1 U15624 ( .C1(n13683), .C2(n14947), .A(n13527), .B(n13526), .ZN(
        P2_U3241) );
  INV_X1 U15625 ( .A(n13530), .ZN(n13528) );
  XNOR2_X1 U15626 ( .A(n13529), .B(n13528), .ZN(n13689) );
  XOR2_X1 U15627 ( .A(n13531), .B(n13530), .Z(n13534) );
  AOI222_X1 U15628 ( .A1(n13618), .A2(n13534), .B1(n13533), .B2(n13496), .C1(
        n13532), .C2(n13462), .ZN(n13688) );
  OAI21_X1 U15629 ( .B1(n13536), .B2(n13535), .A(n13688), .ZN(n13537) );
  NAND2_X1 U15630 ( .A1(n13537), .A2(n13602), .ZN(n13545) );
  INV_X1 U15631 ( .A(n13555), .ZN(n13540) );
  INV_X1 U15632 ( .A(n13538), .ZN(n13539) );
  AOI211_X1 U15633 ( .C1(n13686), .C2(n13540), .A(n10574), .B(n13539), .ZN(
        n13685) );
  OAI22_X1 U15634 ( .A1(n13542), .A2(n13610), .B1(n13602), .B2(n13541), .ZN(
        n13543) );
  AOI21_X1 U15635 ( .B1(n13685), .B2(n13613), .A(n13543), .ZN(n13544) );
  OAI211_X1 U15636 ( .C1(n13689), .C2(n14942), .A(n13545), .B(n13544), .ZN(
        P2_U3242) );
  XNOR2_X1 U15637 ( .A(n13546), .B(n7157), .ZN(n13547) );
  NAND2_X1 U15638 ( .A1(n13547), .A2(n13618), .ZN(n13553) );
  OAI22_X1 U15639 ( .A1(n13550), .A2(n13627), .B1(n13549), .B2(n13548), .ZN(
        n13551) );
  INV_X1 U15640 ( .A(n13551), .ZN(n13552) );
  NAND2_X1 U15641 ( .A1(n13553), .A2(n13552), .ZN(n13695) );
  AND2_X1 U15642 ( .A1(n13571), .A2(n13690), .ZN(n13554) );
  OR3_X1 U15643 ( .A1(n13555), .A2(n13554), .A3(n10574), .ZN(n13692) );
  INV_X1 U15644 ( .A(n13556), .ZN(n13557) );
  AOI22_X1 U15645 ( .A1(n14947), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n14936), 
        .B2(n13557), .ZN(n13559) );
  NAND2_X1 U15646 ( .A1(n13690), .A2(n14935), .ZN(n13558) );
  OAI211_X1 U15647 ( .C1(n13692), .C2(n14939), .A(n13559), .B(n13558), .ZN(
        n13563) );
  OAI21_X1 U15648 ( .B1(n13561), .B2(n7157), .A(n13560), .ZN(n13693) );
  NOR2_X1 U15649 ( .A1(n13693), .A2(n14942), .ZN(n13562) );
  AOI211_X1 U15650 ( .C1(n13602), .C2(n13695), .A(n13563), .B(n13562), .ZN(
        n13564) );
  INV_X1 U15651 ( .A(n13564), .ZN(P2_U3243) );
  XNOR2_X1 U15652 ( .A(n13566), .B(n13565), .ZN(n13568) );
  OAI21_X1 U15653 ( .B1(n13568), .B2(n13600), .A(n13567), .ZN(n13696) );
  INV_X1 U15654 ( .A(n13696), .ZN(n13581) );
  XNOR2_X1 U15655 ( .A(n13570), .B(n13569), .ZN(n13698) );
  INV_X1 U15656 ( .A(n13588), .ZN(n13573) );
  INV_X1 U15657 ( .A(n13571), .ZN(n13572) );
  AOI211_X1 U15658 ( .C1(n13574), .C2(n13573), .A(n10574), .B(n13572), .ZN(
        n13697) );
  NAND2_X1 U15659 ( .A1(n13697), .A2(n13613), .ZN(n13577) );
  AOI22_X1 U15660 ( .A1(n14947), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n13575), 
        .B2(n14936), .ZN(n13576) );
  OAI211_X1 U15661 ( .C1(n13755), .C2(n13610), .A(n13577), .B(n13576), .ZN(
        n13578) );
  AOI21_X1 U15662 ( .B1(n13698), .B2(n13579), .A(n13578), .ZN(n13580) );
  OAI21_X1 U15663 ( .B1(n13581), .B2(n14947), .A(n13580), .ZN(P2_U3244) );
  XNOR2_X1 U15664 ( .A(n13583), .B(n13582), .ZN(n13705) );
  XNOR2_X1 U15665 ( .A(n13585), .B(n13584), .ZN(n13587) );
  OAI21_X1 U15666 ( .B1(n13587), .B2(n13600), .A(n13586), .ZN(n13701) );
  NAND2_X1 U15667 ( .A1(n13701), .A2(n13602), .ZN(n13594) );
  AOI211_X1 U15668 ( .C1(n13703), .C2(n6973), .A(n10574), .B(n13588), .ZN(
        n13702) );
  AOI22_X1 U15669 ( .A1(n14947), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n14936), 
        .B2(n13589), .ZN(n13590) );
  OAI21_X1 U15670 ( .B1(n13591), .B2(n13610), .A(n13590), .ZN(n13592) );
  AOI21_X1 U15671 ( .B1(n13702), .B2(n13613), .A(n13592), .ZN(n13593) );
  OAI211_X1 U15672 ( .C1(n13705), .C2(n14942), .A(n13594), .B(n13593), .ZN(
        P2_U3245) );
  XNOR2_X1 U15673 ( .A(n13596), .B(n13595), .ZN(n13710) );
  XNOR2_X1 U15674 ( .A(n13598), .B(n13597), .ZN(n13601) );
  OAI21_X1 U15675 ( .B1(n13601), .B2(n13600), .A(n13599), .ZN(n13706) );
  NAND2_X1 U15676 ( .A1(n13706), .A2(n13602), .ZN(n13615) );
  NAND2_X1 U15677 ( .A1(n7532), .A2(n13708), .ZN(n13604) );
  NAND2_X1 U15678 ( .A1(n13604), .A2(n13603), .ZN(n13605) );
  NOR2_X1 U15679 ( .A1(n13606), .A2(n13605), .ZN(n13707) );
  INV_X1 U15680 ( .A(n13708), .ZN(n13611) );
  INV_X1 U15681 ( .A(n13607), .ZN(n13608) );
  AOI22_X1 U15682 ( .A1(n14947), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n14936), 
        .B2(n13608), .ZN(n13609) );
  OAI21_X1 U15683 ( .B1(n13611), .B2(n13610), .A(n13609), .ZN(n13612) );
  AOI21_X1 U15684 ( .B1(n13707), .B2(n13613), .A(n13612), .ZN(n13614) );
  OAI211_X1 U15685 ( .C1(n13710), .C2(n14942), .A(n13615), .B(n13614), .ZN(
        P2_U3246) );
  XNOR2_X1 U15686 ( .A(n13617), .B(n13616), .ZN(n13619) );
  NAND2_X1 U15687 ( .A1(n13619), .A2(n13618), .ZN(n13631) );
  NAND2_X1 U15688 ( .A1(n13621), .A2(n13620), .ZN(n13622) );
  NAND2_X1 U15689 ( .A1(n13623), .A2(n13622), .ZN(n13712) );
  INV_X1 U15690 ( .A(n13624), .ZN(n14978) );
  NAND2_X1 U15691 ( .A1(n13625), .A2(n13496), .ZN(n13626) );
  OAI21_X1 U15692 ( .B1(n13628), .B2(n13627), .A(n13626), .ZN(n13629) );
  AOI21_X1 U15693 ( .B1(n13712), .B2(n14978), .A(n13629), .ZN(n13630) );
  NAND2_X1 U15694 ( .A1(n13631), .A2(n13630), .ZN(n13717) );
  INV_X1 U15695 ( .A(n13717), .ZN(n13640) );
  AOI21_X1 U15696 ( .B1(n13632), .B2(n13711), .A(n10574), .ZN(n13633) );
  NAND2_X1 U15697 ( .A1(n13633), .A2(n7532), .ZN(n13713) );
  AOI22_X1 U15698 ( .A1(n14947), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n14936), 
        .B2(n13634), .ZN(n13636) );
  NAND2_X1 U15699 ( .A1(n13711), .A2(n14935), .ZN(n13635) );
  OAI211_X1 U15700 ( .C1(n13713), .C2(n14939), .A(n13636), .B(n13635), .ZN(
        n13637) );
  AOI21_X1 U15701 ( .B1(n13712), .B2(n13638), .A(n13637), .ZN(n13639) );
  OAI21_X1 U15702 ( .B1(n13640), .B2(n14947), .A(n13639), .ZN(P2_U3247) );
  NAND2_X1 U15703 ( .A1(n13641), .A2(n13644), .ZN(n13731) );
  MUX2_X1 U15704 ( .A(n13731), .B(P2_REG1_REG_31__SCAN_IN), .S(n15017), .Z(
        n13642) );
  INV_X1 U15705 ( .A(n13642), .ZN(n13643) );
  OAI21_X1 U15706 ( .B1(n12165), .B2(n13724), .A(n13643), .ZN(P2_U3530) );
  INV_X1 U15707 ( .A(n13644), .ZN(n13645) );
  NOR2_X1 U15708 ( .A1(n13646), .A2(n13645), .ZN(n13736) );
  MUX2_X1 U15709 ( .A(n15329), .B(n13736), .S(n15019), .Z(n13647) );
  OAI21_X1 U15710 ( .B1(n13739), .B2(n13724), .A(n13647), .ZN(P2_U3529) );
  INV_X1 U15711 ( .A(n13648), .ZN(n13654) );
  INV_X1 U15712 ( .A(n13649), .ZN(n13651) );
  MUX2_X1 U15713 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n13740), .S(n15019), .Z(
        P2_U3528) );
  MUX2_X1 U15714 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n13655), .S(n15019), .Z(
        n13656) );
  INV_X1 U15715 ( .A(n13656), .ZN(n13657) );
  OAI21_X1 U15716 ( .B1(n13658), .B2(n13724), .A(n13657), .ZN(P2_U3527) );
  NAND3_X1 U15717 ( .A1(n13660), .A2(n13659), .A3(n14983), .ZN(n13664) );
  NAND2_X1 U15718 ( .A1(n13661), .A2(n14965), .ZN(n13663) );
  NAND3_X1 U15719 ( .A1(n13664), .A2(n13663), .A3(n13662), .ZN(n13665) );
  NOR2_X1 U15720 ( .A1(n13666), .A2(n13665), .ZN(n13741) );
  MUX2_X1 U15721 ( .A(n13667), .B(n13741), .S(n15019), .Z(n13668) );
  INV_X1 U15722 ( .A(n13668), .ZN(P2_U3526) );
  AOI21_X1 U15723 ( .B1(n14965), .B2(n13670), .A(n13669), .ZN(n13671) );
  OAI211_X1 U15724 ( .C1(n13730), .C2(n13673), .A(n13672), .B(n13671), .ZN(
        n13744) );
  MUX2_X1 U15725 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n13744), .S(n15019), .Z(
        P2_U3525) );
  AND2_X1 U15726 ( .A1(n13674), .A2(n14983), .ZN(n13677) );
  NOR3_X1 U15727 ( .A1(n13677), .A2(n13676), .A3(n13675), .ZN(n13746) );
  MUX2_X1 U15728 ( .A(n13746), .B(n13678), .S(n15017), .Z(n13679) );
  OAI21_X1 U15729 ( .B1(n13748), .B2(n13724), .A(n13679), .ZN(P2_U3524) );
  AOI21_X1 U15730 ( .B1(n14965), .B2(n13681), .A(n13680), .ZN(n13682) );
  OAI211_X1 U15731 ( .C1(n14970), .C2(n13684), .A(n13683), .B(n13682), .ZN(
        n13749) );
  MUX2_X1 U15732 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n13749), .S(n15019), .Z(
        P2_U3523) );
  AOI21_X1 U15733 ( .B1(n14965), .B2(n13686), .A(n13685), .ZN(n13687) );
  OAI211_X1 U15734 ( .C1(n13730), .C2(n13689), .A(n13688), .B(n13687), .ZN(
        n13750) );
  MUX2_X1 U15735 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n13750), .S(n15019), .Z(
        P2_U3522) );
  NAND2_X1 U15736 ( .A1(n13690), .A2(n14965), .ZN(n13691) );
  OAI211_X1 U15737 ( .C1(n13693), .C2(n13730), .A(n13692), .B(n13691), .ZN(
        n13694) );
  MUX2_X1 U15738 ( .A(n13751), .B(P2_REG1_REG_22__SCAN_IN), .S(n15017), .Z(
        P2_U3521) );
  INV_X1 U15739 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n13699) );
  AOI211_X1 U15740 ( .C1(n14983), .C2(n13698), .A(n13697), .B(n13696), .ZN(
        n13752) );
  MUX2_X1 U15741 ( .A(n13699), .B(n13752), .S(n15019), .Z(n13700) );
  OAI21_X1 U15742 ( .B1(n13755), .B2(n13724), .A(n13700), .ZN(P2_U3520) );
  AOI211_X1 U15743 ( .C1(n14965), .C2(n13703), .A(n13702), .B(n13701), .ZN(
        n13704) );
  OAI21_X1 U15744 ( .B1(n13730), .B2(n13705), .A(n13704), .ZN(n13756) );
  MUX2_X1 U15745 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n13756), .S(n15019), .Z(
        P2_U3519) );
  AOI211_X1 U15746 ( .C1(n14965), .C2(n13708), .A(n13707), .B(n13706), .ZN(
        n13709) );
  OAI21_X1 U15747 ( .B1(n13730), .B2(n13710), .A(n13709), .ZN(n13757) );
  MUX2_X1 U15748 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n13757), .S(n15019), .Z(
        P2_U3518) );
  INV_X1 U15749 ( .A(n13711), .ZN(n13715) );
  INV_X1 U15750 ( .A(n14970), .ZN(n15004) );
  NAND2_X1 U15751 ( .A1(n13712), .A2(n15004), .ZN(n13714) );
  OAI211_X1 U15752 ( .C1(n13715), .C2(n14999), .A(n13714), .B(n13713), .ZN(
        n13716) );
  NOR2_X1 U15753 ( .A1(n13717), .A2(n13716), .ZN(n13758) );
  MUX2_X1 U15754 ( .A(n14924), .B(n13758), .S(n15019), .Z(n13718) );
  INV_X1 U15755 ( .A(n13718), .ZN(P2_U3517) );
  INV_X1 U15756 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n13722) );
  AOI211_X1 U15757 ( .C1(n14983), .C2(n13721), .A(n13720), .B(n13719), .ZN(
        n13761) );
  MUX2_X1 U15758 ( .A(n13722), .B(n13761), .S(n15019), .Z(n13723) );
  OAI21_X1 U15759 ( .B1(n13765), .B2(n13724), .A(n13723), .ZN(P2_U3516) );
  AOI21_X1 U15760 ( .B1(n14965), .B2(n13726), .A(n13725), .ZN(n13727) );
  OAI211_X1 U15761 ( .C1(n13730), .C2(n13729), .A(n13728), .B(n13727), .ZN(
        n13766) );
  MUX2_X1 U15762 ( .A(n13766), .B(P2_REG1_REG_16__SCAN_IN), .S(n15017), .Z(
        P2_U3515) );
  OR2_X1 U15763 ( .A1(n13731), .A2(n15005), .ZN(n13734) );
  NAND2_X1 U15764 ( .A1(n13734), .A2(n13733), .ZN(n13735) );
  OAI21_X1 U15765 ( .B1(n12165), .B2(n13764), .A(n13735), .ZN(P2_U3498) );
  MUX2_X1 U15766 ( .A(n13737), .B(n13736), .S(n15007), .Z(n13738) );
  OAI21_X1 U15767 ( .B1(n13739), .B2(n13764), .A(n13738), .ZN(P2_U3497) );
  MUX2_X1 U15768 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n13740), .S(n15007), .Z(
        P2_U3496) );
  INV_X1 U15769 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n13742) );
  MUX2_X1 U15770 ( .A(n13742), .B(n13741), .S(n15007), .Z(n13743) );
  INV_X1 U15771 ( .A(n13743), .ZN(P2_U3494) );
  MUX2_X1 U15772 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n13744), .S(n15007), .Z(
        P2_U3493) );
  INV_X1 U15773 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n13745) );
  MUX2_X1 U15774 ( .A(n13746), .B(n13745), .S(n15005), .Z(n13747) );
  OAI21_X1 U15775 ( .B1(n13748), .B2(n13764), .A(n13747), .ZN(P2_U3492) );
  MUX2_X1 U15776 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n13749), .S(n15007), .Z(
        P2_U3491) );
  MUX2_X1 U15777 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n13750), .S(n15007), .Z(
        P2_U3490) );
  MUX2_X1 U15778 ( .A(n13751), .B(P2_REG0_REG_22__SCAN_IN), .S(n15005), .Z(
        P2_U3489) );
  MUX2_X1 U15779 ( .A(n13753), .B(n13752), .S(n15007), .Z(n13754) );
  OAI21_X1 U15780 ( .B1(n13755), .B2(n13764), .A(n13754), .ZN(P2_U3488) );
  MUX2_X1 U15781 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n13756), .S(n15007), .Z(
        P2_U3487) );
  MUX2_X1 U15782 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n13757), .S(n15007), .Z(
        P2_U3486) );
  INV_X1 U15783 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n13759) );
  MUX2_X1 U15784 ( .A(n13759), .B(n13758), .S(n15007), .Z(n13760) );
  INV_X1 U15785 ( .A(n13760), .ZN(P2_U3484) );
  INV_X1 U15786 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n13762) );
  MUX2_X1 U15787 ( .A(n13762), .B(n13761), .S(n15007), .Z(n13763) );
  OAI21_X1 U15788 ( .B1(n13765), .B2(n13764), .A(n13763), .ZN(P2_U3481) );
  MUX2_X1 U15789 ( .A(n13766), .B(P2_REG0_REG_16__SCAN_IN), .S(n15005), .Z(
        P2_U3478) );
  NAND3_X1 U15790 ( .A1(n13767), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .ZN(n13770) );
  OAI22_X1 U15791 ( .A1(n13771), .A2(n13770), .B1(n13769), .B2(n13768), .ZN(
        n13772) );
  AOI21_X1 U15792 ( .B1(n8417), .B2(n13775), .A(n13772), .ZN(n13773) );
  INV_X1 U15793 ( .A(n13773), .ZN(P2_U3296) );
  INV_X1 U15794 ( .A(n13774), .ZN(n14437) );
  NAND2_X1 U15795 ( .A1(n13776), .A2(n13775), .ZN(n13778) );
  OAI211_X1 U15796 ( .C1(n13780), .C2(n13779), .A(n13778), .B(n13777), .ZN(
        P2_U3299) );
  MUX2_X1 U15797 ( .A(n13781), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  XOR2_X1 U15798 ( .A(n13783), .B(n13782), .Z(n13788) );
  AOI22_X1 U15799 ( .A1(n14665), .A2(n13918), .B1(P1_REG3_REG_27__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13785) );
  NAND2_X1 U15800 ( .A1(n13900), .A2(n13919), .ZN(n13784) );
  OAI211_X1 U15801 ( .C1(n14684), .C2(n14092), .A(n13785), .B(n13784), .ZN(
        n13786) );
  AOI21_X1 U15802 ( .B1(n14095), .B2(n14679), .A(n13786), .ZN(n13787) );
  OAI21_X1 U15803 ( .B1(n13788), .B2(n14674), .A(n13787), .ZN(P1_U3214) );
  XOR2_X1 U15804 ( .A(n13790), .B(n13789), .Z(n13796) );
  NOR2_X1 U15805 ( .A1(n13817), .A2(n14276), .ZN(n13791) );
  AOI21_X1 U15806 ( .B1(n13920), .B2(n14247), .A(n13791), .ZN(n14312) );
  NOR2_X1 U15807 ( .A1(n14312), .A2(n13870), .ZN(n13794) );
  OAI22_X1 U15808 ( .A1(n14165), .A2(n14684), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13792), .ZN(n13793) );
  AOI211_X1 U15809 ( .C1(n14160), .C2(n14679), .A(n13794), .B(n13793), .ZN(
        n13795) );
  OAI21_X1 U15810 ( .B1(n13796), .B2(n14674), .A(n13795), .ZN(P1_U3216) );
  INV_X1 U15811 ( .A(n14345), .ZN(n14233) );
  OAI211_X1 U15812 ( .C1(n13799), .C2(n13798), .A(n13797), .B(n13880), .ZN(
        n13802) );
  OAI22_X1 U15813 ( .A1(n13816), .A2(n14770), .B1(n14275), .B2(n14276), .ZN(
        n14344) );
  AND2_X1 U15814 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n14064) );
  NOR2_X1 U15815 ( .A1(n14684), .A2(n14228), .ZN(n13800) );
  AOI211_X1 U15816 ( .C1(n13818), .C2(n14344), .A(n14064), .B(n13800), .ZN(
        n13801) );
  OAI211_X1 U15817 ( .C1(n14233), .C2(n13875), .A(n13802), .B(n13801), .ZN(
        P1_U3219) );
  OAI21_X1 U15818 ( .B1(n13803), .B2(n13805), .A(n13804), .ZN(n13806) );
  NAND2_X1 U15819 ( .A1(n13806), .A2(n13880), .ZN(n13811) );
  AOI22_X1 U15820 ( .A1(n13900), .A2(n13939), .B1(P1_REG3_REG_1__SCAN_IN), 
        .B2(n13882), .ZN(n13810) );
  AOI22_X1 U15821 ( .A1(n14665), .A2(n13808), .B1(n14679), .B2(n13807), .ZN(
        n13809) );
  NAND3_X1 U15822 ( .A1(n13811), .A2(n13810), .A3(n13809), .ZN(P1_U3222) );
  INV_X1 U15823 ( .A(n13812), .ZN(n13813) );
  AOI21_X1 U15824 ( .B1(n13815), .B2(n13814), .A(n13813), .ZN(n13822) );
  OAI22_X1 U15825 ( .A1(n13817), .A2(n14770), .B1(n13816), .B2(n14276), .ZN(
        n14192) );
  AOI22_X1 U15826 ( .A1(n14192), .A2(n13818), .B1(P1_REG3_REG_21__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13819) );
  OAI21_X1 U15827 ( .B1(n14684), .B2(n14197), .A(n13819), .ZN(n13820) );
  AOI21_X1 U15828 ( .B1(n14199), .B2(n14679), .A(n13820), .ZN(n13821) );
  OAI21_X1 U15829 ( .B1(n13822), .B2(n14674), .A(n13821), .ZN(P1_U3223) );
  XOR2_X1 U15830 ( .A(n13824), .B(n13823), .Z(n13829) );
  AND2_X1 U15831 ( .A1(n14247), .A2(n13919), .ZN(n13825) );
  AOI21_X1 U15832 ( .B1(n13920), .B2(n14757), .A(n13825), .ZN(n14300) );
  NOR2_X1 U15833 ( .A1(n14300), .A2(n13870), .ZN(n13827) );
  INV_X1 U15834 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n15391) );
  OAI22_X1 U15835 ( .A1(n14684), .A2(n14126), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15391), .ZN(n13826) );
  AOI211_X1 U15836 ( .C1(n14400), .C2(n14679), .A(n13827), .B(n13826), .ZN(
        n13828) );
  OAI21_X1 U15837 ( .B1(n13829), .B2(n14674), .A(n13828), .ZN(P1_U3225) );
  OAI21_X1 U15838 ( .B1(n13831), .B2(n6662), .A(n13830), .ZN(n13832) );
  NAND2_X1 U15839 ( .A1(n13832), .A2(n13880), .ZN(n13838) );
  NAND2_X1 U15840 ( .A1(n14665), .A2(n13925), .ZN(n13833) );
  OAI211_X1 U15841 ( .C1(n14668), .C2(n14666), .A(n13834), .B(n13833), .ZN(
        n13835) );
  AOI21_X1 U15842 ( .B1(n13836), .B2(n13891), .A(n13835), .ZN(n13837) );
  OAI211_X1 U15843 ( .C1(n14362), .C2(n13875), .A(n13838), .B(n13837), .ZN(
        P1_U3226) );
  OAI21_X1 U15844 ( .B1(n13841), .B2(n13840), .A(n13839), .ZN(n13842) );
  NAND2_X1 U15845 ( .A1(n13842), .A2(n13880), .ZN(n13847) );
  NOR2_X1 U15846 ( .A1(n14684), .A2(n14268), .ZN(n13845) );
  OAI21_X1 U15847 ( .B1(n14668), .B2(n14277), .A(n13843), .ZN(n13844) );
  AOI211_X1 U15848 ( .C1(n14665), .C2(n13924), .A(n13845), .B(n13844), .ZN(
        n13846) );
  OAI211_X1 U15849 ( .C1(n14272), .C2(n13875), .A(n13847), .B(n13846), .ZN(
        P1_U3228) );
  XOR2_X1 U15850 ( .A(n13849), .B(n13848), .Z(n13854) );
  NAND2_X1 U15851 ( .A1(n14140), .A2(n13900), .ZN(n13851) );
  AOI22_X1 U15852 ( .A1(n14665), .A2(n14139), .B1(P1_REG3_REG_24__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13850) );
  OAI211_X1 U15853 ( .C1(n14684), .C2(n14149), .A(n13851), .B(n13850), .ZN(
        n13852) );
  AOI21_X1 U15854 ( .B1(n14148), .B2(n14679), .A(n13852), .ZN(n13853) );
  OAI21_X1 U15855 ( .B1(n13854), .B2(n14674), .A(n13853), .ZN(P1_U3229) );
  OAI211_X1 U15856 ( .C1(n13857), .C2(n13856), .A(n13855), .B(n13880), .ZN(
        n13863) );
  INV_X1 U15857 ( .A(n14212), .ZN(n13861) );
  AND2_X1 U15858 ( .A1(n14248), .A2(n14757), .ZN(n13858) );
  AOI21_X1 U15859 ( .B1(n13922), .B2(n14247), .A(n13858), .ZN(n14335) );
  OAI22_X1 U15860 ( .A1(n14335), .A2(n13870), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13859), .ZN(n13860) );
  AOI21_X1 U15861 ( .B1(n13861), .B2(n13891), .A(n13860), .ZN(n13862) );
  OAI211_X1 U15862 ( .C1(n14213), .C2(n13875), .A(n13863), .B(n13862), .ZN(
        P1_U3233) );
  OAI21_X1 U15863 ( .B1(n13866), .B2(n13865), .A(n13864), .ZN(n13867) );
  NAND2_X1 U15864 ( .A1(n13867), .A2(n13880), .ZN(n13874) );
  INV_X1 U15865 ( .A(n14178), .ZN(n13872) );
  AND2_X1 U15866 ( .A1(n13922), .A2(n14757), .ZN(n13868) );
  AOI21_X1 U15867 ( .B1(n14140), .B2(n14247), .A(n13868), .ZN(n14321) );
  OAI22_X1 U15868 ( .A1(n14321), .A2(n13870), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13869), .ZN(n13871) );
  AOI21_X1 U15869 ( .B1(n13872), .B2(n13891), .A(n13871), .ZN(n13873) );
  OAI211_X1 U15870 ( .C1(n13875), .C2(n14410), .A(n13874), .B(n13873), .ZN(
        P1_U3235) );
  OAI21_X1 U15871 ( .B1(n13879), .B2(n13878), .A(n13877), .ZN(n13881) );
  NAND2_X1 U15872 ( .A1(n13881), .A2(n13880), .ZN(n13888) );
  AOI22_X1 U15873 ( .A1(n13900), .A2(n13883), .B1(P1_REG3_REG_2__SCAN_IN), 
        .B2(n13882), .ZN(n13887) );
  AOI22_X1 U15874 ( .A1(n14665), .A2(n13885), .B1(n14679), .B2(n13884), .ZN(
        n13886) );
  NAND3_X1 U15875 ( .A1(n13888), .A2(n13887), .A3(n13886), .ZN(P1_U3237) );
  XOR2_X1 U15876 ( .A(n13890), .B(n13889), .Z(n13897) );
  NAND2_X1 U15877 ( .A1(n13891), .A2(n14253), .ZN(n13894) );
  NOR2_X1 U15878 ( .A1(n13892), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14035) );
  AOI21_X1 U15879 ( .B1(n14665), .B2(n14248), .A(n14035), .ZN(n13893) );
  OAI211_X1 U15880 ( .C1(n14668), .C2(n14250), .A(n13894), .B(n13893), .ZN(
        n13895) );
  AOI21_X1 U15881 ( .B1(n14350), .B2(n14679), .A(n13895), .ZN(n13896) );
  OAI21_X1 U15882 ( .B1(n13897), .B2(n14674), .A(n13896), .ZN(P1_U3238) );
  AOI22_X1 U15883 ( .A1(n14665), .A2(n14106), .B1(P1_REG3_REG_26__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13902) );
  NAND2_X1 U15884 ( .A1(n13900), .A2(n14139), .ZN(n13901) );
  OAI211_X1 U15885 ( .C1(n14684), .C2(n14112), .A(n13902), .B(n13901), .ZN(
        n13903) );
  AOI21_X1 U15886 ( .B1(n14396), .B2(n14679), .A(n13903), .ZN(n13904) );
  OAI21_X1 U15887 ( .B1(n13905), .B2(n14674), .A(n13904), .ZN(P1_U3240) );
  NAND2_X1 U15888 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n14751)
         );
  OAI21_X1 U15889 ( .B1(n14668), .B2(n13906), .A(n14751), .ZN(n13907) );
  AOI21_X1 U15890 ( .B1(n14665), .B2(n13926), .A(n13907), .ZN(n13908) );
  OAI21_X1 U15891 ( .B1(n14684), .B2(n13909), .A(n13908), .ZN(n13914) );
  AOI211_X1 U15892 ( .C1(n13910), .C2(n13912), .A(n14674), .B(n13911), .ZN(
        n13913) );
  AOI211_X1 U15893 ( .C1(n14373), .C2(n14679), .A(n13914), .B(n13913), .ZN(
        n13915) );
  INV_X1 U15894 ( .A(n13915), .ZN(P1_U3241) );
  MUX2_X1 U15895 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n14068), .S(n13967), .Z(
        P1_U3591) );
  MUX2_X1 U15896 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n13916), .S(P1_U4016), .Z(
        P1_U3590) );
  MUX2_X1 U15897 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n13917), .S(n13967), .Z(
        P1_U3589) );
  MUX2_X1 U15898 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n13918), .S(P1_U4016), .Z(
        P1_U3588) );
  MUX2_X1 U15899 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n14106), .S(P1_U4016), .Z(
        P1_U3587) );
  MUX2_X1 U15900 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n13919), .S(P1_U4016), .Z(
        P1_U3586) );
  MUX2_X1 U15901 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n14139), .S(P1_U4016), .Z(
        P1_U3585) );
  MUX2_X1 U15902 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n13920), .S(P1_U4016), .Z(
        P1_U3584) );
  MUX2_X1 U15903 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n14140), .S(P1_U4016), .Z(
        P1_U3583) );
  MUX2_X1 U15904 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n13921), .S(P1_U4016), .Z(
        P1_U3582) );
  MUX2_X1 U15905 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n13922), .S(n13967), .Z(
        P1_U3581) );
  MUX2_X1 U15906 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n13923), .S(n13967), .Z(
        P1_U3580) );
  MUX2_X1 U15907 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n14248), .S(n13967), .Z(
        P1_U3579) );
  MUX2_X1 U15908 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n13924), .S(P1_U4016), .Z(
        P1_U3578) );
  MUX2_X1 U15909 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n13925), .S(P1_U4016), .Z(
        P1_U3577) );
  MUX2_X1 U15910 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n13926), .S(P1_U4016), .Z(
        P1_U3576) );
  MUX2_X1 U15911 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n13927), .S(P1_U4016), .Z(
        P1_U3575) );
  MUX2_X1 U15912 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n13928), .S(P1_U4016), .Z(
        P1_U3574) );
  MUX2_X1 U15913 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n13929), .S(P1_U4016), .Z(
        P1_U3573) );
  MUX2_X1 U15914 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n13930), .S(P1_U4016), .Z(
        P1_U3572) );
  MUX2_X1 U15915 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n13931), .S(P1_U4016), .Z(
        P1_U3571) );
  MUX2_X1 U15916 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n13932), .S(n13967), .Z(
        P1_U3570) );
  MUX2_X1 U15917 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n13933), .S(n13967), .Z(
        P1_U3569) );
  MUX2_X1 U15918 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n13934), .S(n13967), .Z(
        P1_U3568) );
  MUX2_X1 U15919 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n13935), .S(P1_U4016), .Z(
        P1_U3567) );
  MUX2_X1 U15920 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n13936), .S(n13967), .Z(
        P1_U3566) );
  MUX2_X1 U15921 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n13937), .S(n13967), .Z(
        P1_U3565) );
  MUX2_X1 U15922 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n13938), .S(n13967), .Z(
        P1_U3564) );
  MUX2_X1 U15923 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n13939), .S(n13967), .Z(
        P1_U3560) );
  INV_X1 U15924 ( .A(n14744), .ZN(n14735) );
  INV_X1 U15925 ( .A(n14719), .ZN(n14753) );
  INV_X1 U15926 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n14776) );
  OAI22_X1 U15927 ( .A1(n14753), .A2(n14442), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14776), .ZN(n13940) );
  AOI21_X1 U15928 ( .B1(n13941), .B2(n14735), .A(n13940), .ZN(n13948) );
  OAI211_X1 U15929 ( .C1(n13943), .C2(n13942), .A(n14749), .B(n14721), .ZN(
        n13947) );
  OAI211_X1 U15930 ( .C1(n13964), .C2(n13945), .A(n14059), .B(n13944), .ZN(
        n13946) );
  NAND3_X1 U15931 ( .A1(n13948), .A2(n13947), .A3(n13946), .ZN(P1_U3244) );
  OAI211_X1 U15932 ( .C1(n13951), .C2(n13950), .A(n14749), .B(n13949), .ZN(
        n13961) );
  MUX2_X1 U15933 ( .A(n10521), .B(P1_REG2_REG_3__SCAN_IN), .S(n13957), .Z(
        n13952) );
  NAND3_X1 U15934 ( .A1(n14728), .A2(n13953), .A3(n13952), .ZN(n13954) );
  NAND3_X1 U15935 ( .A1(n14059), .A2(n13980), .A3(n13954), .ZN(n13960) );
  NOR2_X1 U15936 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n13955), .ZN(n13956) );
  AOI21_X1 U15937 ( .B1(n14719), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n13956), .ZN(
        n13959) );
  NAND2_X1 U15938 ( .A1(n14735), .A2(n13957), .ZN(n13958) );
  NAND4_X1 U15939 ( .A1(n13961), .A2(n13960), .A3(n13959), .A4(n13958), .ZN(
        P1_U3246) );
  INV_X1 U15940 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n15326) );
  AOI21_X1 U15941 ( .B1(n14714), .B2(n15326), .A(n8158), .ZN(n14713) );
  MUX2_X1 U15942 ( .A(n13964), .B(n13963), .S(n13962), .Z(n13966) );
  NAND2_X1 U15943 ( .A1(n13966), .A2(n13965), .ZN(n13968) );
  OAI211_X1 U15944 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n14713), .A(n13968), .B(
        n13967), .ZN(n14736) );
  INV_X1 U15945 ( .A(n13969), .ZN(n13970) );
  AOI21_X1 U15946 ( .B1(n14719), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n13970), .ZN(
        n13985) );
  OAI21_X1 U15947 ( .B1(n13973), .B2(n13972), .A(n13971), .ZN(n13974) );
  OAI22_X1 U15948 ( .A1(n13975), .A2(n14744), .B1(n14040), .B2(n13974), .ZN(
        n13976) );
  INV_X1 U15949 ( .A(n13976), .ZN(n13984) );
  MUX2_X1 U15950 ( .A(n10640), .B(P1_REG2_REG_4__SCAN_IN), .S(n13977), .Z(
        n13978) );
  NAND3_X1 U15951 ( .A1(n13980), .A2(n13979), .A3(n13978), .ZN(n13981) );
  NAND3_X1 U15952 ( .A1(n14059), .A2(n13982), .A3(n13981), .ZN(n13983) );
  NAND4_X1 U15953 ( .A1(n14736), .A2(n13985), .A3(n13984), .A4(n13983), .ZN(
        P1_U3247) );
  INV_X1 U15954 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n13987) );
  OAI21_X1 U15955 ( .B1(n14753), .B2(n13987), .A(n13986), .ZN(n13988) );
  AOI21_X1 U15956 ( .B1(n13989), .B2(n14735), .A(n13988), .ZN(n13999) );
  OAI211_X1 U15957 ( .C1(n13992), .C2(n13991), .A(n14749), .B(n13990), .ZN(
        n13998) );
  OR3_X1 U15958 ( .A1(n13995), .A2(n13994), .A3(n13993), .ZN(n13996) );
  NAND3_X1 U15959 ( .A1(n14059), .A2(n14010), .A3(n13996), .ZN(n13997) );
  NAND3_X1 U15960 ( .A1(n13999), .A2(n13998), .A3(n13997), .ZN(P1_U3249) );
  INV_X1 U15961 ( .A(n14000), .ZN(n14003) );
  NOR2_X1 U15962 ( .A1(n14744), .A2(n14001), .ZN(n14002) );
  AOI211_X1 U15963 ( .C1(n14719), .C2(P1_ADDR_REG_7__SCAN_IN), .A(n14003), .B(
        n14002), .ZN(n14015) );
  OAI211_X1 U15964 ( .C1(n14006), .C2(n14005), .A(n14004), .B(n14749), .ZN(
        n14014) );
  INV_X1 U15965 ( .A(n14007), .ZN(n14012) );
  NAND3_X1 U15966 ( .A1(n14010), .A2(n14009), .A3(n14008), .ZN(n14011) );
  NAND3_X1 U15967 ( .A1(n14059), .A2(n14012), .A3(n14011), .ZN(n14013) );
  NAND3_X1 U15968 ( .A1(n14015), .A2(n14014), .A3(n14013), .ZN(P1_U3250) );
  OAI211_X1 U15969 ( .C1(n14018), .C2(n14017), .A(n14016), .B(n14749), .ZN(
        n14029) );
  NOR2_X1 U15970 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7838), .ZN(n14021) );
  NOR2_X1 U15971 ( .A1(n14744), .A2(n14019), .ZN(n14020) );
  AOI211_X1 U15972 ( .C1(n14719), .C2(P1_ADDR_REG_10__SCAN_IN), .A(n14021), 
        .B(n14020), .ZN(n14028) );
  OR3_X1 U15973 ( .A1(n14024), .A2(n14023), .A3(n14022), .ZN(n14025) );
  NAND3_X1 U15974 ( .A1(n14026), .A2(n14059), .A3(n14025), .ZN(n14027) );
  NAND3_X1 U15975 ( .A1(n14029), .A2(n14028), .A3(n14027), .ZN(P1_U3253) );
  INV_X1 U15976 ( .A(n14030), .ZN(n14033) );
  OAI22_X1 U15977 ( .A1(n14033), .A2(n14032), .B1(n14031), .B2(n15434), .ZN(
        n14051) );
  XNOR2_X1 U15978 ( .A(n14051), .B(n14046), .ZN(n14034) );
  NAND2_X1 U15979 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n14034), .ZN(n14054) );
  OAI211_X1 U15980 ( .C1(n14034), .C2(P1_REG2_REG_18__SCAN_IN), .A(n14059), 
        .B(n14054), .ZN(n14045) );
  INV_X1 U15981 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n14037) );
  INV_X1 U15982 ( .A(n14035), .ZN(n14036) );
  OAI21_X1 U15983 ( .B1(n14753), .B2(n14037), .A(n14036), .ZN(n14043) );
  AOI21_X1 U15984 ( .B1(P1_REG1_REG_17__SCAN_IN), .B2(n14039), .A(n14038), 
        .ZN(n14047) );
  XNOR2_X1 U15985 ( .A(n14047), .B(n14046), .ZN(n14041) );
  NOR2_X1 U15986 ( .A1(n14355), .A2(n14041), .ZN(n14049) );
  AOI211_X1 U15987 ( .C1(n14041), .C2(n14355), .A(n14049), .B(n14040), .ZN(
        n14042) );
  AOI211_X1 U15988 ( .C1(n14735), .C2(n14052), .A(n14043), .B(n14042), .ZN(
        n14044) );
  NAND2_X1 U15989 ( .A1(n14045), .A2(n14044), .ZN(P1_U3261) );
  NOR2_X1 U15990 ( .A1(n14047), .A2(n14046), .ZN(n14048) );
  NOR2_X1 U15991 ( .A1(n14049), .A2(n14048), .ZN(n14050) );
  XNOR2_X1 U15992 ( .A(n14050), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n14060) );
  INV_X1 U15993 ( .A(n14060), .ZN(n14057) );
  NAND2_X1 U15994 ( .A1(n14052), .A2(n14051), .ZN(n14053) );
  NAND2_X1 U15995 ( .A1(n14054), .A2(n14053), .ZN(n14055) );
  XOR2_X1 U15996 ( .A(n14055), .B(P1_REG2_REG_19__SCAN_IN), .Z(n14058) );
  OAI21_X1 U15997 ( .B1(n14058), .B2(n14746), .A(n14744), .ZN(n14056) );
  AOI21_X1 U15998 ( .B1(n14057), .B2(n14749), .A(n14056), .ZN(n14063) );
  AOI22_X1 U15999 ( .A1(n14060), .A2(n14749), .B1(n14059), .B2(n14058), .ZN(
        n14062) );
  MUX2_X1 U16000 ( .A(n14063), .B(n14062), .S(n14061), .Z(n14066) );
  INV_X1 U16001 ( .A(n14064), .ZN(n14065) );
  OAI211_X1 U16002 ( .C1(n7554), .C2(n14753), .A(n14066), .B(n14065), .ZN(
        P1_U3262) );
  NOR2_X2 U16003 ( .A1(n14291), .A2(n14073), .ZN(n14072) );
  XNOR2_X1 U16004 ( .A(n14390), .B(n14072), .ZN(n14067) );
  NAND2_X1 U16005 ( .A1(n14288), .A2(n14284), .ZN(n14071) );
  AND2_X1 U16006 ( .A1(n14069), .A2(n14068), .ZN(n14287) );
  INV_X1 U16007 ( .A(n14287), .ZN(n14292) );
  NOR2_X1 U16008 ( .A1(n14281), .A2(n14292), .ZN(n14077) );
  AOI21_X1 U16009 ( .B1(n14281), .B2(P1_REG2_REG_31__SCAN_IN), .A(n14077), 
        .ZN(n14070) );
  OAI211_X1 U16010 ( .C1(n14390), .C2(n14271), .A(n14071), .B(n14070), .ZN(
        P1_U3263) );
  INV_X1 U16011 ( .A(n14072), .ZN(n14075) );
  AOI21_X1 U16012 ( .B1(n14291), .B2(n14073), .A(n14793), .ZN(n14074) );
  NAND2_X1 U16013 ( .A1(n14075), .A2(n14074), .ZN(n14293) );
  NOR2_X1 U16014 ( .A1(n14256), .A2(n14076), .ZN(n14078) );
  AOI211_X1 U16015 ( .C1(n14291), .C2(n14258), .A(n14078), .B(n14077), .ZN(
        n14079) );
  OAI21_X1 U16016 ( .B1(n14293), .B2(n14261), .A(n14079), .ZN(P1_U3264) );
  INV_X1 U16017 ( .A(n14080), .ZN(n14091) );
  INV_X1 U16018 ( .A(n14081), .ZN(n14089) );
  INV_X1 U16019 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n14083) );
  OAI22_X1 U16020 ( .A1(n14256), .A2(n14083), .B1(n14082), .B2(n14777), .ZN(
        n14084) );
  AOI21_X1 U16021 ( .B1(n14085), .B2(n14258), .A(n14084), .ZN(n14086) );
  OAI21_X1 U16022 ( .B1(n14087), .B2(n14261), .A(n14086), .ZN(n14088) );
  AOI21_X1 U16023 ( .B1(n14089), .B2(n14235), .A(n14088), .ZN(n14090) );
  OAI21_X1 U16024 ( .B1(n14091), .B2(n14281), .A(n14090), .ZN(P1_U3265) );
  INV_X1 U16025 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n14093) );
  OAI22_X1 U16026 ( .A1(n14256), .A2(n14093), .B1(n14092), .B2(n14777), .ZN(
        n14094) );
  AOI21_X1 U16027 ( .B1(n14095), .B2(n14258), .A(n14094), .ZN(n14098) );
  OR2_X1 U16028 ( .A1(n14096), .A2(n14261), .ZN(n14097) );
  OAI211_X1 U16029 ( .C1(n14099), .C2(n14281), .A(n14098), .B(n14097), .ZN(
        P1_U3266) );
  XNOR2_X1 U16030 ( .A(n14101), .B(n14100), .ZN(n14297) );
  OAI21_X1 U16031 ( .B1(n14104), .B2(n14103), .A(n14102), .ZN(n14105) );
  NAND2_X1 U16032 ( .A1(n14105), .A2(n14783), .ZN(n14108) );
  AOI22_X1 U16033 ( .A1(n14247), .A2(n14106), .B1(n14757), .B2(n14139), .ZN(
        n14107) );
  INV_X1 U16034 ( .A(n14296), .ZN(n14117) );
  AOI21_X1 U16035 ( .B1(n14396), .B2(n14109), .A(n14793), .ZN(n14111) );
  NAND2_X1 U16036 ( .A1(n14111), .A2(n14110), .ZN(n14295) );
  OAI22_X1 U16037 ( .A1(n14256), .A2(n14113), .B1(n14112), .B2(n14777), .ZN(
        n14114) );
  AOI21_X1 U16038 ( .B1(n14396), .B2(n14258), .A(n14114), .ZN(n14115) );
  OAI21_X1 U16039 ( .B1(n14295), .B2(n14261), .A(n14115), .ZN(n14116) );
  AOI21_X1 U16040 ( .B1(n14117), .B2(n14256), .A(n14116), .ZN(n14118) );
  OAI21_X1 U16041 ( .B1(n14286), .B2(n14297), .A(n14118), .ZN(P1_U3267) );
  NAND2_X1 U16042 ( .A1(n14120), .A2(n14123), .ZN(n14121) );
  NAND2_X1 U16043 ( .A1(n14119), .A2(n14121), .ZN(n14302) );
  INV_X1 U16044 ( .A(n14302), .ZN(n14135) );
  OAI21_X1 U16045 ( .B1(n14124), .B2(n14123), .A(n14122), .ZN(n14305) );
  INV_X1 U16046 ( .A(n14305), .ZN(n14133) );
  XNOR2_X1 U16047 ( .A(n14146), .B(n14400), .ZN(n14125) );
  OR2_X1 U16048 ( .A1(n14125), .A2(n14793), .ZN(n14301) );
  INV_X1 U16049 ( .A(n14300), .ZN(n14129) );
  INV_X1 U16050 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n14127) );
  OAI22_X1 U16051 ( .A1(n14256), .A2(n14127), .B1(n14126), .B2(n14777), .ZN(
        n14128) );
  AOI21_X1 U16052 ( .B1(n14129), .B2(n14256), .A(n14128), .ZN(n14131) );
  NAND2_X1 U16053 ( .A1(n14400), .A2(n14258), .ZN(n14130) );
  OAI211_X1 U16054 ( .C1(n14301), .C2(n14261), .A(n14131), .B(n14130), .ZN(
        n14132) );
  AOI21_X1 U16055 ( .B1(n14133), .B2(n14235), .A(n14132), .ZN(n14134) );
  OAI21_X1 U16056 ( .B1(n14135), .B2(n14237), .A(n14134), .ZN(P1_U3268) );
  INV_X1 U16057 ( .A(n14136), .ZN(n14137) );
  AOI21_X1 U16058 ( .B1(n14142), .B2(n14138), .A(n14137), .ZN(n14145) );
  AOI22_X1 U16059 ( .A1(n14140), .A2(n14757), .B1(n14247), .B2(n14139), .ZN(
        n14144) );
  OAI211_X1 U16060 ( .C1(n7547), .C2(n14142), .A(n14783), .B(n14141), .ZN(
        n14143) );
  OAI211_X1 U16061 ( .C1(n14145), .C2(n14755), .A(n14144), .B(n14143), .ZN(
        n14309) );
  INV_X1 U16062 ( .A(n14309), .ZN(n14154) );
  INV_X1 U16063 ( .A(n14146), .ZN(n14147) );
  AOI211_X1 U16064 ( .C1(n14148), .C2(n7027), .A(n14793), .B(n14147), .ZN(
        n14308) );
  INV_X1 U16065 ( .A(n14149), .ZN(n14150) );
  AOI22_X1 U16066 ( .A1(n14150), .A2(n14786), .B1(n14281), .B2(
        P1_REG2_REG_24__SCAN_IN), .ZN(n14151) );
  OAI21_X1 U16067 ( .B1(n14405), .B2(n14271), .A(n14151), .ZN(n14152) );
  AOI21_X1 U16068 ( .B1(n14308), .B2(n14284), .A(n14152), .ZN(n14153) );
  OAI21_X1 U16069 ( .B1(n14154), .B2(n14281), .A(n14153), .ZN(P1_U3269) );
  OAI21_X1 U16070 ( .B1(n14155), .B2(n8061), .A(n14156), .ZN(n14318) );
  OAI21_X1 U16071 ( .B1(n14159), .B2(n14158), .A(n14157), .ZN(n14316) );
  INV_X1 U16072 ( .A(n14160), .ZN(n14313) );
  NAND2_X1 U16073 ( .A1(n14160), .A2(n14176), .ZN(n14161) );
  NAND2_X1 U16074 ( .A1(n14161), .A2(n14365), .ZN(n14162) );
  NOR2_X1 U16075 ( .A1(n14163), .A2(n14162), .ZN(n14315) );
  NAND2_X1 U16076 ( .A1(n14315), .A2(n14284), .ZN(n14169) );
  INV_X1 U16077 ( .A(n14312), .ZN(n14167) );
  OAI22_X1 U16078 ( .A1(n14165), .A2(n14777), .B1(n14256), .B2(n14164), .ZN(
        n14166) );
  AOI21_X1 U16079 ( .B1(n14167), .B2(n14256), .A(n14166), .ZN(n14168) );
  OAI211_X1 U16080 ( .C1(n14313), .C2(n14271), .A(n14169), .B(n14168), .ZN(
        n14170) );
  AOI21_X1 U16081 ( .B1(n14316), .B2(n14218), .A(n14170), .ZN(n14171) );
  OAI21_X1 U16082 ( .B1(n14286), .B2(n14318), .A(n14171), .ZN(P1_U3270) );
  XNOR2_X1 U16083 ( .A(n14172), .B(n14174), .ZN(n14324) );
  INV_X1 U16084 ( .A(n14324), .ZN(n14186) );
  OAI21_X1 U16085 ( .B1(n14175), .B2(n14174), .A(n14173), .ZN(n14319) );
  INV_X1 U16086 ( .A(n14196), .ZN(n14177) );
  OAI211_X1 U16087 ( .C1(n14177), .C2(n14410), .A(n14365), .B(n14176), .ZN(
        n14320) );
  NOR2_X1 U16088 ( .A1(n14320), .A2(n14261), .ZN(n14184) );
  INV_X1 U16089 ( .A(n14321), .ZN(n14181) );
  INV_X1 U16090 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n14179) );
  OAI22_X1 U16091 ( .A1(n14256), .A2(n14179), .B1(n14178), .B2(n14777), .ZN(
        n14180) );
  AOI21_X1 U16092 ( .B1(n14181), .B2(n14256), .A(n14180), .ZN(n14182) );
  OAI21_X1 U16093 ( .B1(n14410), .B2(n14271), .A(n14182), .ZN(n14183) );
  AOI211_X1 U16094 ( .C1(n14319), .C2(n14235), .A(n14184), .B(n14183), .ZN(
        n14185) );
  OAI21_X1 U16095 ( .B1(n14186), .B2(n14237), .A(n14185), .ZN(P1_U3271) );
  XNOR2_X1 U16096 ( .A(n14188), .B(n14187), .ZN(n14328) );
  INV_X1 U16097 ( .A(n14328), .ZN(n14202) );
  XNOR2_X1 U16098 ( .A(n14189), .B(n14190), .ZN(n14191) );
  NAND2_X1 U16099 ( .A1(n14191), .A2(n14783), .ZN(n14194) );
  INV_X1 U16100 ( .A(n14192), .ZN(n14193) );
  NAND2_X1 U16101 ( .A1(n14194), .A2(n14193), .ZN(n14333) );
  OR2_X1 U16102 ( .A1(n14211), .A2(n14329), .ZN(n14195) );
  NAND2_X1 U16103 ( .A1(n14196), .A2(n14195), .ZN(n14330) );
  OAI22_X1 U16104 ( .A1(n14330), .A2(n10823), .B1(n14197), .B2(n14777), .ZN(
        n14198) );
  OAI21_X1 U16105 ( .B1(n14333), .B2(n14198), .A(n14256), .ZN(n14201) );
  AOI22_X1 U16106 ( .A1(n14199), .A2(n14258), .B1(P1_REG2_REG_21__SCAN_IN), 
        .B2(n14281), .ZN(n14200) );
  OAI211_X1 U16107 ( .C1(n14202), .C2(n14286), .A(n14201), .B(n14200), .ZN(
        P1_U3272) );
  XNOR2_X1 U16108 ( .A(n14204), .B(n14203), .ZN(n14339) );
  NAND2_X1 U16109 ( .A1(n14206), .A2(n14205), .ZN(n14207) );
  NAND2_X1 U16110 ( .A1(n14208), .A2(n14207), .ZN(n14334) );
  INV_X1 U16111 ( .A(n14334), .ZN(n14219) );
  NAND2_X1 U16112 ( .A1(n14226), .A2(n14415), .ZN(n14209) );
  NAND2_X1 U16113 ( .A1(n14209), .A2(n14365), .ZN(n14210) );
  OR2_X1 U16114 ( .A1(n14211), .A2(n14210), .ZN(n14336) );
  OAI22_X1 U16115 ( .A1(n14281), .A2(n14335), .B1(n14212), .B2(n14777), .ZN(
        n14215) );
  NOR2_X1 U16116 ( .A1(n14213), .A2(n14271), .ZN(n14214) );
  AOI211_X1 U16117 ( .C1(n14281), .C2(P1_REG2_REG_20__SCAN_IN), .A(n14215), 
        .B(n14214), .ZN(n14216) );
  OAI21_X1 U16118 ( .B1(n14261), .B2(n14336), .A(n14216), .ZN(n14217) );
  AOI21_X1 U16119 ( .B1(n14219), .B2(n14218), .A(n14217), .ZN(n14220) );
  OAI21_X1 U16120 ( .B1(n14286), .B2(n14339), .A(n14220), .ZN(P1_U3273) );
  XNOR2_X1 U16121 ( .A(n14221), .B(n14223), .ZN(n14349) );
  INV_X1 U16122 ( .A(n14222), .ZN(n14225) );
  OAI21_X1 U16123 ( .B1(n14225), .B2(n7229), .A(n14224), .ZN(n14346) );
  INV_X1 U16124 ( .A(n14226), .ZN(n14227) );
  AOI211_X1 U16125 ( .C1(n14345), .C2(n14238), .A(n14793), .B(n14227), .ZN(
        n14343) );
  NAND2_X1 U16126 ( .A1(n14343), .A2(n14284), .ZN(n14232) );
  INV_X1 U16127 ( .A(n14344), .ZN(n14229) );
  OAI22_X1 U16128 ( .A1(n14229), .A2(n14281), .B1(n14228), .B2(n14777), .ZN(
        n14230) );
  AOI21_X1 U16129 ( .B1(P1_REG2_REG_19__SCAN_IN), .B2(n14281), .A(n14230), 
        .ZN(n14231) );
  OAI211_X1 U16130 ( .C1(n14233), .C2(n14271), .A(n14232), .B(n14231), .ZN(
        n14234) );
  AOI21_X1 U16131 ( .B1(n14346), .B2(n14235), .A(n14234), .ZN(n14236) );
  OAI21_X1 U16132 ( .B1(n14349), .B2(n14237), .A(n14236), .ZN(P1_U3274) );
  AOI21_X1 U16133 ( .B1(n14265), .B2(n14350), .A(n14793), .ZN(n14239) );
  NAND2_X1 U16134 ( .A1(n14239), .A2(n14238), .ZN(n14352) );
  NAND2_X1 U16135 ( .A1(n14240), .A2(n14783), .ZN(n14241) );
  OAI21_X1 U16136 ( .B1(n14242), .B2(n14755), .A(n14241), .ZN(n14246) );
  NAND2_X1 U16137 ( .A1(n14242), .A2(n14803), .ZN(n14243) );
  OAI21_X1 U16138 ( .B1(n14240), .B2(n14761), .A(n14243), .ZN(n14245) );
  MUX2_X1 U16139 ( .A(n14246), .B(n14245), .S(n14244), .Z(n14252) );
  NAND2_X1 U16140 ( .A1(n14248), .A2(n14247), .ZN(n14249) );
  OAI21_X1 U16141 ( .B1(n14250), .B2(n14276), .A(n14249), .ZN(n14251) );
  NAND2_X1 U16142 ( .A1(n14354), .A2(n14256), .ZN(n14260) );
  INV_X1 U16143 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n14255) );
  INV_X1 U16144 ( .A(n14253), .ZN(n14254) );
  OAI22_X1 U16145 ( .A1(n14256), .A2(n14255), .B1(n14254), .B2(n14777), .ZN(
        n14257) );
  AOI21_X1 U16146 ( .B1(n14350), .B2(n14258), .A(n14257), .ZN(n14259) );
  OAI211_X1 U16147 ( .C1(n14352), .C2(n14261), .A(n14260), .B(n14259), .ZN(
        P1_U3275) );
  XNOR2_X1 U16148 ( .A(n14263), .B(n14262), .ZN(n14361) );
  INV_X1 U16149 ( .A(n14264), .ZN(n14267) );
  INV_X1 U16150 ( .A(n14265), .ZN(n14266) );
  AOI211_X1 U16151 ( .C1(n14358), .C2(n14267), .A(n14793), .B(n14266), .ZN(
        n14357) );
  INV_X1 U16152 ( .A(n14268), .ZN(n14269) );
  AOI22_X1 U16153 ( .A1(n14281), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n14269), 
        .B2(n14786), .ZN(n14270) );
  OAI21_X1 U16154 ( .B1(n14272), .B2(n14271), .A(n14270), .ZN(n14283) );
  AOI21_X1 U16155 ( .B1(n14274), .B2(n14273), .A(n14761), .ZN(n14280) );
  OAI22_X1 U16156 ( .A1(n14277), .A2(n14276), .B1(n14275), .B2(n14770), .ZN(
        n14278) );
  AOI21_X1 U16157 ( .B1(n14280), .B2(n14279), .A(n14278), .ZN(n14360) );
  NOR2_X1 U16158 ( .A1(n14360), .A2(n14281), .ZN(n14282) );
  AOI211_X1 U16159 ( .C1(n14357), .C2(n14284), .A(n14283), .B(n14282), .ZN(
        n14285) );
  OAI21_X1 U16160 ( .B1(n14286), .B2(n14361), .A(n14285), .ZN(P1_U3276) );
  NOR2_X1 U16161 ( .A1(n14288), .A2(n14287), .ZN(n14387) );
  MUX2_X1 U16162 ( .A(n14289), .B(n14387), .S(n14811), .Z(n14290) );
  OAI21_X1 U16163 ( .B1(n14390), .B2(n14327), .A(n14290), .ZN(P1_U3559) );
  INV_X1 U16164 ( .A(n14291), .ZN(n14393) );
  AND2_X1 U16165 ( .A1(n14293), .A2(n14292), .ZN(n14391) );
  MUX2_X1 U16166 ( .A(n15242), .B(n14391), .S(n14811), .Z(n14294) );
  OAI21_X1 U16167 ( .B1(n14393), .B2(n14327), .A(n14294), .ZN(P1_U3558) );
  OAI211_X1 U16168 ( .C1(n14297), .C2(n14755), .A(n14296), .B(n14295), .ZN(
        n14394) );
  MUX2_X1 U16169 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n14394), .S(n14811), .Z(
        n14298) );
  AOI21_X1 U16170 ( .B1(n14341), .B2(n14396), .A(n14298), .ZN(n14299) );
  INV_X1 U16171 ( .A(n14299), .ZN(P1_U3554) );
  AND2_X1 U16172 ( .A1(n14301), .A2(n14300), .ZN(n14304) );
  NAND2_X1 U16173 ( .A1(n14302), .A2(n14783), .ZN(n14303) );
  OAI211_X1 U16174 ( .C1(n14305), .C2(n14755), .A(n14304), .B(n14303), .ZN(
        n14398) );
  MUX2_X1 U16175 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n14398), .S(n14811), .Z(
        n14306) );
  AOI21_X1 U16176 ( .B1(n14341), .B2(n14400), .A(n14306), .ZN(n14307) );
  INV_X1 U16177 ( .A(n14307), .ZN(P1_U3553) );
  INV_X1 U16178 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n14310) );
  NOR2_X1 U16179 ( .A1(n14309), .A2(n14308), .ZN(n14402) );
  MUX2_X1 U16180 ( .A(n14310), .B(n14402), .S(n14811), .Z(n14311) );
  OAI21_X1 U16181 ( .B1(n14405), .B2(n14327), .A(n14311), .ZN(P1_U3552) );
  OAI21_X1 U16182 ( .B1(n14313), .B2(n14798), .A(n14312), .ZN(n14314) );
  AOI211_X1 U16183 ( .C1(n14316), .C2(n14783), .A(n14315), .B(n14314), .ZN(
        n14317) );
  OAI21_X1 U16184 ( .B1(n14755), .B2(n14318), .A(n14317), .ZN(n14406) );
  MUX2_X1 U16185 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n14406), .S(n14811), .Z(
        P1_U3551) );
  INV_X1 U16186 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n14325) );
  INV_X1 U16187 ( .A(n14319), .ZN(n14322) );
  OAI211_X1 U16188 ( .C1(n14322), .C2(n14755), .A(n14321), .B(n14320), .ZN(
        n14323) );
  AOI21_X1 U16189 ( .B1(n14783), .B2(n14324), .A(n14323), .ZN(n14407) );
  MUX2_X1 U16190 ( .A(n14325), .B(n14407), .S(n14811), .Z(n14326) );
  OAI21_X1 U16191 ( .B1(n14327), .B2(n14410), .A(n14326), .ZN(P1_U3550) );
  AND2_X1 U16192 ( .A1(n14328), .A2(n14803), .ZN(n14332) );
  OAI22_X1 U16193 ( .A1(n14330), .A2(n14793), .B1(n14329), .B2(n14798), .ZN(
        n14331) );
  MUX2_X1 U16194 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n14412), .S(n14811), .Z(
        P1_U3549) );
  OR2_X1 U16195 ( .A1(n14334), .A2(n14761), .ZN(n14338) );
  AND2_X1 U16196 ( .A1(n14336), .A2(n14335), .ZN(n14337) );
  OAI211_X1 U16197 ( .C1(n14339), .C2(n14755), .A(n14338), .B(n14337), .ZN(
        n14413) );
  MUX2_X1 U16198 ( .A(n14413), .B(P1_REG1_REG_20__SCAN_IN), .S(n14809), .Z(
        n14340) );
  AOI21_X1 U16199 ( .B1(n14341), .B2(n14415), .A(n14340), .ZN(n14342) );
  INV_X1 U16200 ( .A(n14342), .ZN(P1_U3548) );
  AOI211_X1 U16201 ( .C1(n14372), .C2(n14345), .A(n14344), .B(n14343), .ZN(
        n14348) );
  NAND2_X1 U16202 ( .A1(n14346), .A2(n14803), .ZN(n14347) );
  OAI211_X1 U16203 ( .C1(n14349), .C2(n14761), .A(n14348), .B(n14347), .ZN(
        n14418) );
  MUX2_X1 U16204 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n14418), .S(n14811), .Z(
        P1_U3547) );
  NAND2_X1 U16205 ( .A1(n14350), .A2(n14372), .ZN(n14351) );
  NAND2_X1 U16206 ( .A1(n14352), .A2(n14351), .ZN(n14353) );
  NOR2_X1 U16207 ( .A1(n14354), .A2(n14353), .ZN(n14419) );
  MUX2_X1 U16208 ( .A(n14355), .B(n14419), .S(n14811), .Z(n14356) );
  INV_X1 U16209 ( .A(n14356), .ZN(P1_U3546) );
  AOI21_X1 U16210 ( .B1(n14372), .B2(n14358), .A(n14357), .ZN(n14359) );
  OAI211_X1 U16211 ( .C1(n14755), .C2(n14361), .A(n14360), .B(n14359), .ZN(
        n14421) );
  MUX2_X1 U16212 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n14421), .S(n14811), .Z(
        P1_U3545) );
  NOR2_X1 U16213 ( .A1(n14362), .A2(n14798), .ZN(n14364) );
  AOI211_X1 U16214 ( .C1(n14366), .C2(n14365), .A(n14364), .B(n14363), .ZN(
        n14369) );
  NAND2_X1 U16215 ( .A1(n14367), .A2(n14803), .ZN(n14368) );
  OAI211_X1 U16216 ( .C1(n14370), .C2(n14761), .A(n14369), .B(n14368), .ZN(
        n14422) );
  MUX2_X1 U16217 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n14422), .S(n14811), .Z(
        P1_U3544) );
  AOI21_X1 U16218 ( .B1(n14373), .B2(n14372), .A(n14371), .ZN(n14374) );
  OAI21_X1 U16219 ( .B1(n14375), .B2(n14793), .A(n14374), .ZN(n14376) );
  AOI21_X1 U16220 ( .B1(n14377), .B2(n14783), .A(n14376), .ZN(n14378) );
  OAI21_X1 U16221 ( .B1(n14755), .B2(n14379), .A(n14378), .ZN(n14423) );
  MUX2_X1 U16222 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n14423), .S(n14811), .Z(
        P1_U3543) );
  OAI211_X1 U16223 ( .C1(n14382), .C2(n14798), .A(n14381), .B(n14380), .ZN(
        n14383) );
  AOI21_X1 U16224 ( .B1(n14384), .B2(n14803), .A(n14383), .ZN(n14385) );
  OAI21_X1 U16225 ( .B1(n14386), .B2(n14761), .A(n14385), .ZN(n14424) );
  MUX2_X1 U16226 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n14424), .S(n14811), .Z(
        P1_U3541) );
  MUX2_X1 U16227 ( .A(n14388), .B(n14387), .S(n14806), .Z(n14389) );
  OAI21_X1 U16228 ( .B1(n14390), .B2(n14411), .A(n14389), .ZN(P1_U3527) );
  MUX2_X1 U16229 ( .A(n15488), .B(n14391), .S(n14806), .Z(n14392) );
  OAI21_X1 U16230 ( .B1(n14393), .B2(n14411), .A(n14392), .ZN(P1_U3526) );
  MUX2_X1 U16231 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n14394), .S(n14806), .Z(
        n14395) );
  AOI21_X1 U16232 ( .B1(n14416), .B2(n14396), .A(n14395), .ZN(n14397) );
  INV_X1 U16233 ( .A(n14397), .ZN(P1_U3522) );
  MUX2_X1 U16234 ( .A(n14398), .B(P1_REG0_REG_25__SCAN_IN), .S(n14804), .Z(
        n14399) );
  AOI21_X1 U16235 ( .B1(n14416), .B2(n14400), .A(n14399), .ZN(n14401) );
  INV_X1 U16236 ( .A(n14401), .ZN(P1_U3521) );
  MUX2_X1 U16237 ( .A(n14403), .B(n14402), .S(n14806), .Z(n14404) );
  OAI21_X1 U16238 ( .B1(n14405), .B2(n14411), .A(n14404), .ZN(P1_U3520) );
  MUX2_X1 U16239 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n14406), .S(n14806), .Z(
        P1_U3519) );
  MUX2_X1 U16240 ( .A(n14408), .B(n14407), .S(n14806), .Z(n14409) );
  OAI21_X1 U16241 ( .B1(n14411), .B2(n14410), .A(n14409), .ZN(P1_U3518) );
  MUX2_X1 U16242 ( .A(n14412), .B(P1_REG0_REG_21__SCAN_IN), .S(n14804), .Z(
        P1_U3517) );
  MUX2_X1 U16243 ( .A(n14413), .B(P1_REG0_REG_20__SCAN_IN), .S(n14804), .Z(
        n14414) );
  AOI21_X1 U16244 ( .B1(n14416), .B2(n14415), .A(n14414), .ZN(n14417) );
  INV_X1 U16245 ( .A(n14417), .ZN(P1_U3516) );
  MUX2_X1 U16246 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n14418), .S(n14806), .Z(
        P1_U3515) );
  MUX2_X1 U16247 ( .A(n15416), .B(n14419), .S(n14806), .Z(n14420) );
  INV_X1 U16248 ( .A(n14420), .ZN(P1_U3513) );
  MUX2_X1 U16249 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n14421), .S(n14806), .Z(
        P1_U3510) );
  MUX2_X1 U16250 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n14422), .S(n14806), .Z(
        P1_U3507) );
  MUX2_X1 U16251 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n14423), .S(n14806), .Z(
        P1_U3504) );
  MUX2_X1 U16252 ( .A(P1_REG0_REG_13__SCAN_IN), .B(n14424), .S(n14806), .Z(
        P1_U3498) );
  NAND2_X1 U16253 ( .A1(n8417), .A2(n14425), .ZN(n14429) );
  NAND2_X1 U16254 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_STATE_REG_SCAN_IN), 
        .ZN(n14426) );
  OR3_X1 U16255 ( .A1(n14427), .A2(P1_IR_REG_30__SCAN_IN), .A3(n14426), .ZN(
        n14428) );
  OAI211_X1 U16256 ( .C1(n14430), .C2(n14433), .A(n14429), .B(n14428), .ZN(
        P1_U3324) );
  OAI222_X1 U16257 ( .A1(n12610), .A2(n14432), .B1(P1_U3086), .B2(n7502), .C1(
        n14431), .C2(n14433), .ZN(P1_U3325) );
  OAI222_X1 U16258 ( .A1(n12610), .A2(n14437), .B1(P1_U3086), .B2(n14435), 
        .C1(n14434), .C2(n14433), .ZN(P1_U3326) );
  MUX2_X1 U16259 ( .A(n14439), .B(n14438), .S(P1_U3086), .Z(P1_U3333) );
  MUX2_X1 U16260 ( .A(n14440), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  NOR2_X1 U16261 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(n14537), .ZN(n14477) );
  INV_X1 U16262 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n14474) );
  INV_X1 U16263 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n14471) );
  INV_X1 U16264 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n14468) );
  XNOR2_X1 U16265 ( .A(P3_ADDR_REG_12__SCAN_IN), .B(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n14528) );
  INV_X1 U16266 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n14466) );
  INV_X1 U16267 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n14464) );
  INV_X1 U16268 ( .A(P3_ADDR_REG_9__SCAN_IN), .ZN(n14462) );
  XNOR2_X1 U16269 ( .A(P3_ADDR_REG_9__SCAN_IN), .B(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n14518) );
  INV_X1 U16270 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n14460) );
  INV_X1 U16271 ( .A(n14490), .ZN(n14441) );
  XNOR2_X1 U16272 ( .A(n14444), .B(P3_ADDR_REG_2__SCAN_IN), .ZN(n14488) );
  INV_X1 U16273 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n14448) );
  INV_X1 U16274 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n14450) );
  NOR2_X1 U16275 ( .A1(n14449), .A2(n14450), .ZN(n14452) );
  INV_X1 U16276 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n14453) );
  AND2_X1 U16277 ( .A1(n14453), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n14454) );
  NOR2_X1 U16278 ( .A1(P3_ADDR_REG_7__SCAN_IN), .A2(n14455), .ZN(n14458) );
  XNOR2_X1 U16279 ( .A(P3_ADDR_REG_7__SCAN_IN), .B(n14455), .ZN(n14510) );
  INV_X1 U16280 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n14456) );
  XNOR2_X1 U16281 ( .A(n14460), .B(P1_ADDR_REG_8__SCAN_IN), .ZN(n14483) );
  NAND2_X1 U16282 ( .A1(n14518), .A2(n14517), .ZN(n14461) );
  XOR2_X1 U16283 ( .A(P3_ADDR_REG_10__SCAN_IN), .B(P1_ADDR_REG_10__SCAN_IN), 
        .Z(n14481) );
  XNOR2_X1 U16284 ( .A(n14466), .B(P1_ADDR_REG_11__SCAN_IN), .ZN(n14522) );
  NAND2_X1 U16285 ( .A1(n14528), .A2(n14527), .ZN(n14467) );
  INV_X1 U16286 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n14469) );
  NAND2_X1 U16287 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(n14469), .ZN(n14470) );
  AOI22_X1 U16288 ( .A1(P3_ADDR_REG_13__SCAN_IN), .A2(n14471), .B1(n14529), 
        .B2(n14470), .ZN(n14532) );
  INV_X1 U16289 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n14472) );
  XNOR2_X1 U16290 ( .A(n14472), .B(P1_ADDR_REG_14__SCAN_IN), .ZN(n14533) );
  NOR2_X1 U16291 ( .A1(n14532), .A2(n14533), .ZN(n14473) );
  AOI21_X1 U16292 ( .B1(P3_ADDR_REG_14__SCAN_IN), .B2(n14474), .A(n14473), 
        .ZN(n14534) );
  INV_X1 U16293 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n14754) );
  NOR2_X1 U16294 ( .A1(P3_ADDR_REG_15__SCAN_IN), .A2(n14754), .ZN(n14476) );
  OAI22_X1 U16295 ( .A1(n14534), .A2(n14476), .B1(P1_ADDR_REG_15__SCAN_IN), 
        .B2(n14475), .ZN(n14538) );
  NAND2_X1 U16296 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(n14537), .ZN(n14536) );
  OAI21_X1 U16297 ( .B1(n14477), .B2(n14538), .A(n14536), .ZN(n14478) );
  NOR2_X1 U16298 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(n14478), .ZN(n14480) );
  XOR2_X1 U16299 ( .A(P1_ADDR_REG_17__SCAN_IN), .B(n14478), .Z(n14543) );
  AND2_X1 U16300 ( .A1(P3_ADDR_REG_17__SCAN_IN), .A2(n14543), .ZN(n14479) );
  XOR2_X1 U16301 ( .A(P3_ADDR_REG_18__SCAN_IN), .B(P1_ADDR_REG_18__SCAN_IN), 
        .Z(n14568) );
  XOR2_X1 U16302 ( .A(n14567), .B(n14568), .Z(n14548) );
  INV_X1 U16303 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n14891) );
  INV_X1 U16304 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n14868) );
  XOR2_X1 U16305 ( .A(n14482), .B(n14481), .Z(n14561) );
  XOR2_X1 U16306 ( .A(n14484), .B(n14483), .Z(n14515) );
  XNOR2_X1 U16307 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(n14485), .ZN(n14486) );
  NAND2_X1 U16308 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(n14486), .ZN(n14500) );
  INV_X1 U16309 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n14841) );
  XNOR2_X1 U16310 ( .A(n14486), .B(n14841), .ZN(n15521) );
  XNOR2_X1 U16311 ( .A(n14488), .B(n14487), .ZN(n14553) );
  XOR2_X1 U16312 ( .A(n14490), .B(n14489), .Z(n14491) );
  NAND2_X1 U16313 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n14491), .ZN(n14493) );
  AOI21_X1 U16314 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(n15027), .A(n14490), .ZN(
        n15524) );
  INV_X1 U16315 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n15523) );
  NOR2_X1 U16316 ( .A1(n15524), .A2(n15523), .ZN(n15532) );
  NAND2_X1 U16317 ( .A1(n14493), .A2(n14492), .ZN(n14554) );
  NAND2_X1 U16318 ( .A1(n14553), .A2(n14554), .ZN(n14494) );
  NOR2_X1 U16319 ( .A1(n14553), .A2(n14554), .ZN(n14552) );
  XNOR2_X1 U16320 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(n14495), .ZN(n14497) );
  NOR2_X1 U16321 ( .A1(n14496), .A2(n14497), .ZN(n15527) );
  NOR2_X1 U16322 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(n15528), .ZN(n14498) );
  NAND2_X1 U16323 ( .A1(n15521), .A2(n15520), .ZN(n14499) );
  NAND2_X1 U16324 ( .A1(n14500), .A2(n14499), .ZN(n14503) );
  NOR2_X1 U16325 ( .A1(n14503), .A2(n14502), .ZN(n14505) );
  XNOR2_X1 U16326 ( .A(n14503), .B(n14502), .ZN(n15522) );
  NOR2_X1 U16327 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n15522), .ZN(n14504) );
  NAND2_X1 U16328 ( .A1(n14506), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n14509) );
  XNOR2_X1 U16329 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(P3_ADDR_REG_6__SCAN_IN), 
        .ZN(n14508) );
  XOR2_X1 U16330 ( .A(n14508), .B(n14507), .Z(n14556) );
  NAND2_X1 U16331 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n14511), .ZN(n14513) );
  XNOR2_X1 U16332 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n14510), .ZN(n15526) );
  NAND2_X1 U16333 ( .A1(n15526), .A2(n15525), .ZN(n14512) );
  NOR2_X1 U16334 ( .A1(n14515), .A2(n14514), .ZN(n14516) );
  XNOR2_X1 U16335 ( .A(n14518), .B(n14517), .ZN(n14520) );
  NAND2_X1 U16336 ( .A1(n14519), .A2(n14520), .ZN(n14521) );
  XOR2_X1 U16337 ( .A(n14523), .B(n14522), .Z(n14524) );
  NOR2_X1 U16338 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(n14692), .ZN(n14526) );
  XNOR2_X1 U16339 ( .A(n14528), .B(n14527), .ZN(n14696) );
  XNOR2_X1 U16340 ( .A(P3_ADDR_REG_13__SCAN_IN), .B(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n14530) );
  XNOR2_X1 U16341 ( .A(n14530), .B(n14529), .ZN(n14700) );
  INV_X1 U16342 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n15464) );
  NAND2_X1 U16343 ( .A1(n14701), .A2(n14700), .ZN(n14699) );
  OAI21_X2 U16344 ( .B1(n14531), .B2(n15464), .A(n14699), .ZN(n14703) );
  XNOR2_X1 U16345 ( .A(n14533), .B(n14532), .ZN(n14704) );
  XNOR2_X1 U16346 ( .A(P1_ADDR_REG_15__SCAN_IN), .B(P3_ADDR_REG_15__SCAN_IN), 
        .ZN(n14535) );
  XOR2_X1 U16347 ( .A(n14535), .B(n14534), .Z(n14708) );
  OAI21_X1 U16348 ( .B1(n14537), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n14536), 
        .ZN(n14539) );
  XOR2_X1 U16349 ( .A(n14539), .B(n14538), .Z(n14540) );
  NOR2_X1 U16350 ( .A1(n14541), .A2(n14540), .ZN(n14711) );
  NOR2_X1 U16351 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(n14710), .ZN(n14542) );
  XNOR2_X1 U16352 ( .A(P3_ADDR_REG_17__SCAN_IN), .B(n14543), .ZN(n14545) );
  NOR2_X1 U16353 ( .A1(n14544), .A2(n14545), .ZN(n14565) );
  NOR2_X1 U16354 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(n14564), .ZN(n14546) );
  NOR2_X1 U16355 ( .A1(n14548), .A2(n14547), .ZN(n14574) );
  NOR2_X1 U16356 ( .A1(n14574), .A2(n14573), .ZN(n14549) );
  XOR2_X1 U16357 ( .A(P2_ADDR_REG_18__SCAN_IN), .B(n14549), .Z(SUB_1596_U62)
         );
  AOI21_X1 U16358 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n14550) );
  OAI21_X1 U16359 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n14550), 
        .ZN(U28) );
  AOI21_X1 U16360 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        P3_RD_REG_SCAN_IN), .ZN(n14551) );
  OAI21_X1 U16361 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(n14551), 
        .ZN(U29) );
  AOI21_X1 U16362 ( .B1(n14554), .B2(n14553), .A(n14552), .ZN(n14555) );
  XNOR2_X1 U16363 ( .A(n14555), .B(n9907), .ZN(SUB_1596_U61) );
  XOR2_X1 U16364 ( .A(n14557), .B(n14556), .Z(SUB_1596_U57) );
  XNOR2_X1 U16365 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n14558), .ZN(SUB_1596_U55)
         );
  XOR2_X1 U16366 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n14559), .Z(SUB_1596_U54) );
  AOI21_X1 U16367 ( .B1(n14561), .B2(n14560), .A(n6661), .ZN(n14563) );
  XNOR2_X1 U16368 ( .A(n14563), .B(n14562), .ZN(SUB_1596_U70) );
  NOR2_X1 U16369 ( .A1(n14565), .A2(n14564), .ZN(n14566) );
  XOR2_X1 U16370 ( .A(P2_ADDR_REG_17__SCAN_IN), .B(n14566), .Z(SUB_1596_U63)
         );
  INV_X1 U16371 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n15449) );
  NOR2_X1 U16372 ( .A1(n14568), .A2(n14567), .ZN(n14569) );
  AOI21_X1 U16373 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n15449), .A(n14569), 
        .ZN(n14570) );
  XOR2_X1 U16374 ( .A(n14570), .B(P3_ADDR_REG_19__SCAN_IN), .Z(n14572) );
  XNOR2_X1 U16375 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n14571) );
  XNOR2_X1 U16376 ( .A(n14572), .B(n14571), .ZN(n14575) );
  AOI21_X1 U16377 ( .B1(n8824), .B2(n14577), .A(n14576), .ZN(n14591) );
  OAI21_X1 U16378 ( .B1(n14579), .B2(P3_REG1_REG_17__SCAN_IN), .A(n14578), 
        .ZN(n14589) );
  INV_X1 U16379 ( .A(P3_ADDR_REG_17__SCAN_IN), .ZN(n14583) );
  NAND2_X1 U16380 ( .A1(n15031), .A2(n14580), .ZN(n14582) );
  OAI211_X1 U16381 ( .C1(n14583), .C2(n15028), .A(n14582), .B(n14581), .ZN(
        n14588) );
  AOI211_X1 U16382 ( .C1(n14586), .C2(n14585), .A(n15102), .B(n14584), .ZN(
        n14587) );
  AOI211_X1 U16383 ( .C1(n15109), .C2(n14589), .A(n14588), .B(n14587), .ZN(
        n14590) );
  OAI21_X1 U16384 ( .B1(n14591), .B2(n15113), .A(n14590), .ZN(P3_U3199) );
  AOI22_X1 U16385 ( .A1(n15031), .A2(n14592), .B1(n15106), .B2(
        P3_ADDR_REG_18__SCAN_IN), .ZN(n14608) );
  XNOR2_X1 U16386 ( .A(n14594), .B(n14593), .ZN(n14600) );
  AOI21_X1 U16387 ( .B1(n14597), .B2(n14596), .A(n14595), .ZN(n14598) );
  NOR2_X1 U16388 ( .A1(n14598), .A2(n15102), .ZN(n14599) );
  AOI21_X1 U16389 ( .B1(n15109), .B2(n14600), .A(n14599), .ZN(n14607) );
  INV_X1 U16390 ( .A(n14601), .ZN(n14604) );
  OAI221_X1 U16391 ( .B1(n14604), .B2(n14603), .C1(n14604), .C2(n14602), .A(
        n15023), .ZN(n14605) );
  NOR2_X1 U16392 ( .A1(n14610), .A2(n14609), .ZN(n14622) );
  AOI22_X1 U16393 ( .A1(n15150), .A2(n14611), .B1(n14622), .B2(n15132), .ZN(
        n14619) );
  OAI22_X1 U16394 ( .A1(n14614), .A2(n14613), .B1(n15132), .B2(n14612), .ZN(
        n14615) );
  INV_X1 U16395 ( .A(n14615), .ZN(n14616) );
  NAND2_X1 U16396 ( .A1(n14619), .A2(n14616), .ZN(P3_U3202) );
  AOI22_X1 U16397 ( .A1(n14623), .A2(n14617), .B1(P3_REG2_REG_30__SCAN_IN), 
        .B2(n13074), .ZN(n14618) );
  NAND2_X1 U16398 ( .A1(n14619), .A2(n14618), .ZN(P3_U3203) );
  AOI21_X1 U16399 ( .B1(n14620), .B2(n14638), .A(n14622), .ZN(n14639) );
  INV_X1 U16400 ( .A(P3_REG1_REG_31__SCAN_IN), .ZN(n14621) );
  AOI22_X1 U16401 ( .A1(n15222), .A2(n14639), .B1(n14621), .B2(n9126), .ZN(
        P3_U3490) );
  AOI21_X1 U16402 ( .B1(n14623), .B2(n14638), .A(n14622), .ZN(n14641) );
  INV_X1 U16403 ( .A(P3_REG1_REG_30__SCAN_IN), .ZN(n14624) );
  AOI22_X1 U16404 ( .A1(n15222), .A2(n14641), .B1(n14624), .B2(n9126), .ZN(
        P3_U3489) );
  OAI22_X1 U16405 ( .A1(n14626), .A2(n15201), .B1(n15200), .B2(n14625), .ZN(
        n14627) );
  NOR2_X1 U16406 ( .A1(n14628), .A2(n14627), .ZN(n14643) );
  INV_X1 U16407 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n14629) );
  AOI22_X1 U16408 ( .A1(n15222), .A2(n14643), .B1(n14629), .B2(n9126), .ZN(
        P3_U3472) );
  NOR2_X1 U16409 ( .A1(n14630), .A2(n15201), .ZN(n14632) );
  AOI211_X1 U16410 ( .C1(n14638), .C2(n14633), .A(n14632), .B(n14631), .ZN(
        n14645) );
  AOI22_X1 U16411 ( .A1(n15222), .A2(n14645), .B1(n11493), .B2(n9126), .ZN(
        P3_U3471) );
  NOR2_X1 U16412 ( .A1(n14634), .A2(n15201), .ZN(n14636) );
  AOI211_X1 U16413 ( .C1(n14638), .C2(n14637), .A(n14636), .B(n14635), .ZN(
        n14647) );
  INV_X1 U16414 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n15355) );
  AOI22_X1 U16415 ( .A1(n15222), .A2(n14647), .B1(n15355), .B2(n9126), .ZN(
        P3_U3470) );
  INV_X1 U16416 ( .A(P3_REG0_REG_31__SCAN_IN), .ZN(n14640) );
  AOI22_X1 U16417 ( .A1(n15206), .A2(n14640), .B1(n14639), .B2(n15205), .ZN(
        P3_U3458) );
  INV_X1 U16418 ( .A(P3_REG0_REG_30__SCAN_IN), .ZN(n14642) );
  AOI22_X1 U16419 ( .A1(n15206), .A2(n14642), .B1(n14641), .B2(n15205), .ZN(
        P3_U3457) );
  INV_X1 U16420 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n14644) );
  AOI22_X1 U16421 ( .A1(n15206), .A2(n14644), .B1(n14643), .B2(n15205), .ZN(
        P3_U3429) );
  INV_X1 U16422 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n14646) );
  AOI22_X1 U16423 ( .A1(n15206), .A2(n14646), .B1(n14645), .B2(n15205), .ZN(
        P3_U3426) );
  INV_X1 U16424 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n14648) );
  AOI22_X1 U16425 ( .A1(n15206), .A2(n14648), .B1(n14647), .B2(n15205), .ZN(
        P3_U3423) );
  OAI21_X1 U16426 ( .B1(n14650), .B2(n14999), .A(n14649), .ZN(n14653) );
  INV_X1 U16427 ( .A(n14651), .ZN(n14652) );
  AOI211_X1 U16428 ( .C1(n14654), .C2(n14983), .A(n14653), .B(n14652), .ZN(
        n14662) );
  AOI22_X1 U16429 ( .A1(n15019), .A2(n14662), .B1(n9341), .B2(n15017), .ZN(
        P2_U3513) );
  INV_X1 U16430 ( .A(n14655), .ZN(n14660) );
  OAI21_X1 U16431 ( .B1(n14657), .B2(n14999), .A(n14656), .ZN(n14659) );
  AOI211_X1 U16432 ( .C1(n15004), .C2(n14660), .A(n14659), .B(n14658), .ZN(
        n14664) );
  AOI22_X1 U16433 ( .A1(n15019), .A2(n14664), .B1(n11093), .B2(n15017), .ZN(
        P2_U3511) );
  INV_X1 U16434 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n14661) );
  AOI22_X1 U16435 ( .A1(n15007), .A2(n14662), .B1(n14661), .B2(n15005), .ZN(
        P2_U3472) );
  INV_X1 U16436 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n14663) );
  AOI22_X1 U16437 ( .A1(n15007), .A2(n14664), .B1(n14663), .B2(n15005), .ZN(
        P2_U3466) );
  INV_X1 U16438 ( .A(n14665), .ZN(n14667) );
  OAI22_X1 U16439 ( .A1(n14669), .A2(n14668), .B1(n14667), .B2(n14666), .ZN(
        n14678) );
  NAND2_X1 U16440 ( .A1(n14671), .A2(n14670), .ZN(n14673) );
  NAND2_X1 U16441 ( .A1(n14673), .A2(n14672), .ZN(n14675) );
  AOI21_X1 U16442 ( .B1(n14676), .B2(n14675), .A(n14674), .ZN(n14677) );
  AOI211_X1 U16443 ( .C1(n14680), .C2(n14679), .A(n14678), .B(n14677), .ZN(
        n14682) );
  OAI211_X1 U16444 ( .C1(n14684), .C2(n14683), .A(n14682), .B(n14681), .ZN(
        P1_U3215) );
  OAI21_X1 U16445 ( .B1(n14686), .B2(n14798), .A(n14685), .ZN(n14688) );
  AOI211_X1 U16446 ( .C1(n14803), .C2(n14689), .A(n14688), .B(n14687), .ZN(
        n14691) );
  AOI22_X1 U16447 ( .A1(n14811), .A2(n14691), .B1(n10399), .B2(n14809), .ZN(
        P1_U3539) );
  INV_X1 U16448 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n14690) );
  AOI22_X1 U16449 ( .A1(n14806), .A2(n14691), .B1(n14690), .B2(n14804), .ZN(
        P1_U3492) );
  NOR2_X1 U16450 ( .A1(n14693), .A2(n14692), .ZN(n14694) );
  XOR2_X1 U16451 ( .A(P2_ADDR_REG_11__SCAN_IN), .B(n14694), .Z(SUB_1596_U69)
         );
  AOI21_X1 U16452 ( .B1(n14697), .B2(n14696), .A(n14695), .ZN(n14698) );
  XNOR2_X1 U16453 ( .A(n14698), .B(n14868), .ZN(SUB_1596_U68) );
  OAI21_X1 U16454 ( .B1(n14701), .B2(n14700), .A(n14699), .ZN(n14702) );
  XNOR2_X1 U16455 ( .A(n14702), .B(P2_ADDR_REG_13__SCAN_IN), .ZN(SUB_1596_U67)
         );
  AOI21_X1 U16456 ( .B1(n14704), .B2(n14703), .A(n6655), .ZN(n14705) );
  XNOR2_X1 U16457 ( .A(n14705), .B(n11103), .ZN(SUB_1596_U66) );
  AOI21_X1 U16458 ( .B1(n14708), .B2(n14707), .A(n14706), .ZN(n14709) );
  XNOR2_X1 U16459 ( .A(n14709), .B(n14891), .ZN(SUB_1596_U65) );
  NOR2_X1 U16460 ( .A1(n14711), .A2(n14710), .ZN(n14712) );
  XOR2_X1 U16461 ( .A(P2_ADDR_REG_16__SCAN_IN), .B(n14712), .Z(SUB_1596_U64)
         );
  OAI21_X1 U16462 ( .B1(n14714), .B2(P1_REG1_REG_0__SCAN_IN), .A(n14713), .ZN(
        n14715) );
  XOR2_X1 U16463 ( .A(P1_IR_REG_0__SCAN_IN), .B(n14715), .Z(n14718) );
  AOI22_X1 U16464 ( .A1(n14719), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n14716) );
  OAI21_X1 U16465 ( .B1(n14718), .B2(n14717), .A(n14716), .ZN(P1_U3243) );
  AOI22_X1 U16466 ( .A1(n14719), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n14738) );
  INV_X1 U16467 ( .A(n14727), .ZN(n14734) );
  INV_X1 U16468 ( .A(n14720), .ZN(n14723) );
  NAND3_X1 U16469 ( .A1(n14723), .A2(n14722), .A3(n14721), .ZN(n14724) );
  AND3_X1 U16470 ( .A1(n14749), .A2(n14725), .A3(n14724), .ZN(n14733) );
  INV_X1 U16471 ( .A(n14726), .ZN(n14731) );
  MUX2_X1 U16472 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n15433), .S(n14727), .Z(
        n14730) );
  INV_X1 U16473 ( .A(n14728), .ZN(n14729) );
  AOI211_X1 U16474 ( .C1(n14731), .C2(n14730), .A(n14729), .B(n14746), .ZN(
        n14732) );
  AOI211_X1 U16475 ( .C1(n14735), .C2(n14734), .A(n14733), .B(n14732), .ZN(
        n14737) );
  NAND3_X1 U16476 ( .A1(n14738), .A2(n14737), .A3(n14736), .ZN(P1_U3245) );
  OAI21_X1 U16477 ( .B1(n14741), .B2(n14740), .A(n14739), .ZN(n14750) );
  AOI21_X1 U16478 ( .B1(n14743), .B2(P1_REG2_REG_15__SCAN_IN), .A(n14742), 
        .ZN(n14747) );
  OAI22_X1 U16479 ( .A1(n14747), .A2(n14746), .B1(n14745), .B2(n14744), .ZN(
        n14748) );
  AOI21_X1 U16480 ( .B1(n14750), .B2(n14749), .A(n14748), .ZN(n14752) );
  OAI211_X1 U16481 ( .C1(n14754), .C2(n14753), .A(n14752), .B(n14751), .ZN(
        P1_U3258) );
  NOR2_X1 U16482 ( .A1(n14755), .A2(n14760), .ZN(n14756) );
  MUX2_X1 U16483 ( .A(n14783), .B(n14756), .S(n8434), .Z(n14758) );
  NOR2_X1 U16484 ( .A1(n14758), .A2(n14757), .ZN(n14765) );
  OAI21_X1 U16485 ( .B1(n14760), .B2(n14792), .A(n14759), .ZN(n14794) );
  XNOR2_X1 U16486 ( .A(n14794), .B(n10352), .ZN(n14762) );
  OR2_X1 U16487 ( .A1(n14762), .A2(n14761), .ZN(n14764) );
  MUX2_X1 U16488 ( .A(n14765), .B(n14764), .S(n14763), .Z(n14769) );
  INV_X1 U16489 ( .A(n14766), .ZN(n14767) );
  NAND2_X1 U16490 ( .A1(n14767), .A2(n14803), .ZN(n14768) );
  OAI211_X1 U16491 ( .C1(n14771), .C2(n14770), .A(n14769), .B(n14768), .ZN(
        n14796) );
  OAI22_X1 U16492 ( .A1(n14794), .A2(n10823), .B1(n14792), .B2(n14772), .ZN(
        n14773) );
  NOR2_X1 U16493 ( .A1(n14796), .A2(n14773), .ZN(n14774) );
  MUX2_X1 U16494 ( .A(n14774), .B(n9935), .S(n14281), .Z(n14775) );
  OAI21_X1 U16495 ( .B1(n14777), .B2(n14776), .A(n14775), .ZN(P1_U3292) );
  INV_X1 U16496 ( .A(n14778), .ZN(n14784) );
  AOI21_X1 U16497 ( .B1(n14780), .B2(n8153), .A(n14779), .ZN(n14790) );
  INV_X1 U16498 ( .A(n14781), .ZN(n14782) );
  OAI21_X1 U16499 ( .B1(n14803), .B2(n14783), .A(n14782), .ZN(n14791) );
  OAI21_X1 U16500 ( .B1(n14784), .B2(n14790), .A(n14791), .ZN(n14785) );
  AOI22_X1 U16501 ( .A1(n14786), .A2(P1_REG3_REG_0__SCAN_IN), .B1(n14256), 
        .B2(n14785), .ZN(n14787) );
  OAI21_X1 U16502 ( .B1(n15326), .B2(n14256), .A(n14787), .ZN(P1_U3293) );
  INV_X1 U16503 ( .A(n14789), .ZN(n14788) );
  NOR2_X1 U16504 ( .A1(n14788), .A2(n15418), .ZN(P1_U3294) );
  AND2_X1 U16505 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n14789), .ZN(P1_U3295) );
  AND2_X1 U16506 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n14789), .ZN(P1_U3296) );
  INV_X1 U16507 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n15392) );
  NOR2_X1 U16508 ( .A1(n14788), .A2(n15392), .ZN(P1_U3297) );
  AND2_X1 U16509 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n14789), .ZN(P1_U3298) );
  AND2_X1 U16510 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n14789), .ZN(P1_U3299) );
  AND2_X1 U16511 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n14789), .ZN(P1_U3300) );
  AND2_X1 U16512 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n14789), .ZN(P1_U3301) );
  NOR2_X1 U16513 ( .A1(n14788), .A2(n15389), .ZN(P1_U3302) );
  AND2_X1 U16514 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n14789), .ZN(P1_U3303) );
  AND2_X1 U16515 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n14789), .ZN(P1_U3304) );
  AND2_X1 U16516 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n14789), .ZN(P1_U3305) );
  AND2_X1 U16517 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n14789), .ZN(P1_U3306) );
  AND2_X1 U16518 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n14789), .ZN(P1_U3307) );
  AND2_X1 U16519 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n14789), .ZN(P1_U3308) );
  AND2_X1 U16520 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n14789), .ZN(P1_U3309) );
  AND2_X1 U16521 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n14789), .ZN(P1_U3310) );
  AND2_X1 U16522 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n14789), .ZN(P1_U3311) );
  NOR2_X1 U16523 ( .A1(n14788), .A2(n15240), .ZN(P1_U3312) );
  AND2_X1 U16524 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n14789), .ZN(P1_U3313) );
  AND2_X1 U16525 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n14789), .ZN(P1_U3314) );
  AND2_X1 U16526 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n14789), .ZN(P1_U3315) );
  AND2_X1 U16527 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n14789), .ZN(P1_U3316) );
  AND2_X1 U16528 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n14789), .ZN(P1_U3317) );
  AND2_X1 U16529 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n14789), .ZN(P1_U3318) );
  AND2_X1 U16530 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n14789), .ZN(P1_U3319) );
  NOR2_X1 U16531 ( .A1(n14788), .A2(n15356), .ZN(P1_U3320) );
  AND2_X1 U16532 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n14789), .ZN(P1_U3321) );
  AND2_X1 U16533 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n14789), .ZN(P1_U3322) );
  AND2_X1 U16534 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n14789), .ZN(P1_U3323) );
  AND2_X1 U16535 ( .A1(n14791), .A2(n14790), .ZN(n14807) );
  AOI22_X1 U16536 ( .A1(n14806), .A2(n14807), .B1(n7692), .B2(n14804), .ZN(
        P1_U3459) );
  OAI22_X1 U16537 ( .A1(n14794), .A2(n14793), .B1(n14792), .B2(n14798), .ZN(
        n14795) );
  NOR2_X1 U16538 ( .A1(n14796), .A2(n14795), .ZN(n14808) );
  AOI22_X1 U16539 ( .A1(n14806), .A2(n14808), .B1(n7676), .B2(n14804), .ZN(
        P1_U3462) );
  OAI21_X1 U16540 ( .B1(n14799), .B2(n14798), .A(n14797), .ZN(n14801) );
  AOI211_X1 U16541 ( .C1(n14803), .C2(n14802), .A(n14801), .B(n14800), .ZN(
        n14810) );
  INV_X1 U16542 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n14805) );
  AOI22_X1 U16543 ( .A1(n14806), .A2(n14810), .B1(n14805), .B2(n14804), .ZN(
        P1_U3486) );
  AOI22_X1 U16544 ( .A1(n14811), .A2(n14807), .B1(n7691), .B2(n14809), .ZN(
        P1_U3528) );
  AOI22_X1 U16545 ( .A1(n14811), .A2(n14808), .B1(n15442), .B2(n14809), .ZN(
        P1_U3529) );
  AOI22_X1 U16546 ( .A1(n14811), .A2(n14810), .B1(n10160), .B2(n14809), .ZN(
        P1_U3537) );
  NOR2_X1 U16547 ( .A1(n14813), .A2(P2_U3947), .ZN(P2_U3087) );
  AOI22_X1 U16548 ( .A1(P2_REG1_REG_0__SCAN_IN), .A2(n14846), .B1(n14929), 
        .B2(P2_REG2_REG_0__SCAN_IN), .ZN(n14816) );
  OAI22_X1 U16549 ( .A1(P2_REG2_REG_0__SCAN_IN), .A2(n14907), .B1(n14922), 
        .B2(P2_REG1_REG_0__SCAN_IN), .ZN(n14812) );
  NOR2_X1 U16550 ( .A1(n14914), .A2(n14812), .ZN(n14815) );
  AOI22_X1 U16551 ( .A1(n14813), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3088), .ZN(n14814) );
  OAI221_X1 U16552 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n14816), .C1(n9160), .C2(
        n14815), .A(n14814), .ZN(P2_U3214) );
  INV_X1 U16553 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n15529) );
  OAI211_X1 U16554 ( .C1(n14819), .C2(n14818), .A(n14929), .B(n14817), .ZN(
        n14824) );
  OAI211_X1 U16555 ( .C1(n14822), .C2(n14821), .A(n14846), .B(n14820), .ZN(
        n14823) );
  OAI211_X1 U16556 ( .C1(n14921), .C2(n14825), .A(n14824), .B(n14823), .ZN(
        n14826) );
  INV_X1 U16557 ( .A(n14826), .ZN(n14828) );
  NAND2_X1 U16558 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_U3088), .ZN(n14827) );
  OAI211_X1 U16559 ( .C1(n14932), .C2(n15529), .A(n14828), .B(n14827), .ZN(
        P2_U3217) );
  OAI211_X1 U16560 ( .C1(n14831), .C2(n14830), .A(n14929), .B(n14829), .ZN(
        n14836) );
  OAI211_X1 U16561 ( .C1(n14834), .C2(n14833), .A(n14846), .B(n14832), .ZN(
        n14835) );
  OAI211_X1 U16562 ( .C1(n14921), .C2(n14837), .A(n14836), .B(n14835), .ZN(
        n14838) );
  INV_X1 U16563 ( .A(n14838), .ZN(n14840) );
  OAI211_X1 U16564 ( .C1(n14932), .C2(n14841), .A(n14840), .B(n14839), .ZN(
        P2_U3218) );
  INV_X1 U16565 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n14855) );
  OAI211_X1 U16566 ( .C1(n14844), .C2(n14843), .A(n14842), .B(n14929), .ZN(
        n14850) );
  OAI211_X1 U16567 ( .C1(n14848), .C2(n14847), .A(n14846), .B(n14845), .ZN(
        n14849) );
  OAI211_X1 U16568 ( .C1(n14921), .C2(n14851), .A(n14850), .B(n14849), .ZN(
        n14852) );
  INV_X1 U16569 ( .A(n14852), .ZN(n14854) );
  OAI211_X1 U16570 ( .C1(n14855), .C2(n14932), .A(n14854), .B(n14853), .ZN(
        P2_U3222) );
  AOI21_X1 U16571 ( .B1(n14914), .B2(n14857), .A(n14856), .ZN(n14867) );
  XNOR2_X1 U16572 ( .A(n14859), .B(n14858), .ZN(n14865) );
  NAND2_X1 U16573 ( .A1(n14861), .A2(n14860), .ZN(n14862) );
  AOI21_X1 U16574 ( .B1(n14863), .B2(n14862), .A(n14922), .ZN(n14864) );
  AOI21_X1 U16575 ( .B1(n14865), .B2(n14929), .A(n14864), .ZN(n14866) );
  OAI211_X1 U16576 ( .C1(n14868), .C2(n14932), .A(n14867), .B(n14866), .ZN(
        P2_U3226) );
  INV_X1 U16577 ( .A(n14869), .ZN(n14870) );
  AOI211_X1 U16578 ( .C1(n14872), .C2(n14871), .A(n14922), .B(n14870), .ZN(
        n14877) );
  AOI211_X1 U16579 ( .C1(n14875), .C2(n14874), .A(n14907), .B(n14873), .ZN(
        n14876) );
  AOI211_X1 U16580 ( .C1(n14914), .C2(n14878), .A(n14877), .B(n14876), .ZN(
        n14880) );
  NAND2_X1 U16581 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_U3088), .ZN(n14879)
         );
  OAI211_X1 U16582 ( .C1(n15464), .C2(n14932), .A(n14880), .B(n14879), .ZN(
        P2_U3227) );
  AOI211_X1 U16583 ( .C1(n14882), .C2(n9357), .A(n14881), .B(n14907), .ZN(
        n14887) );
  AOI211_X1 U16584 ( .C1(n14885), .C2(n14884), .A(n14883), .B(n14922), .ZN(
        n14886) );
  AOI211_X1 U16585 ( .C1(n14914), .C2(n14888), .A(n14887), .B(n14886), .ZN(
        n14890) );
  NAND2_X1 U16586 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(P2_U3088), .ZN(n14889)
         );
  OAI211_X1 U16587 ( .C1(n14891), .C2(n14932), .A(n14890), .B(n14889), .ZN(
        P2_U3229) );
  INV_X1 U16588 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n14903) );
  AOI211_X1 U16589 ( .C1(n14894), .C2(n14893), .A(n14892), .B(n14907), .ZN(
        n14899) );
  AOI211_X1 U16590 ( .C1(n14897), .C2(n14896), .A(n14895), .B(n14922), .ZN(
        n14898) );
  AOI211_X1 U16591 ( .C1(n14914), .C2(n14900), .A(n14899), .B(n14898), .ZN(
        n14902) );
  OAI211_X1 U16592 ( .C1(n14903), .C2(n14932), .A(n14902), .B(n14901), .ZN(
        P2_U3230) );
  INV_X1 U16593 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n14917) );
  AOI211_X1 U16594 ( .C1(n14906), .C2(n14905), .A(n14904), .B(n14922), .ZN(
        n14912) );
  AOI211_X1 U16595 ( .C1(n14910), .C2(n14909), .A(n14908), .B(n14907), .ZN(
        n14911) );
  AOI211_X1 U16596 ( .C1(n14914), .C2(n14913), .A(n14912), .B(n14911), .ZN(
        n14916) );
  OAI211_X1 U16597 ( .C1(n14917), .C2(n14932), .A(n14916), .B(n14915), .ZN(
        P2_U3231) );
  INV_X1 U16598 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n14933) );
  OAI21_X1 U16599 ( .B1(n14919), .B2(n9395), .A(n14918), .ZN(n14928) );
  NOR2_X1 U16600 ( .A1(n14921), .A2(n14920), .ZN(n14927) );
  AOI211_X1 U16601 ( .C1(n14925), .C2(n14924), .A(n14923), .B(n14922), .ZN(
        n14926) );
  AOI211_X1 U16602 ( .C1(n14929), .C2(n14928), .A(n14927), .B(n14926), .ZN(
        n14931) );
  OAI211_X1 U16603 ( .C1(n14933), .C2(n14932), .A(n14931), .B(n14930), .ZN(
        P2_U3232) );
  NAND2_X1 U16604 ( .A1(n14935), .A2(n14934), .ZN(n14938) );
  AOI22_X1 U16605 ( .A1(n14947), .A2(P2_REG2_REG_1__SCAN_IN), .B1(n14936), 
        .B2(P2_REG3_REG_1__SCAN_IN), .ZN(n14937) );
  OAI211_X1 U16606 ( .C1(n14940), .C2(n14939), .A(n14938), .B(n14937), .ZN(
        n14944) );
  NOR2_X1 U16607 ( .A1(n14942), .A2(n14941), .ZN(n14943) );
  NOR2_X1 U16608 ( .A1(n14944), .A2(n14943), .ZN(n14945) );
  OAI21_X1 U16609 ( .B1(n14947), .B2(n14946), .A(n14945), .ZN(P2_U3264) );
  NOR2_X1 U16610 ( .A1(n14956), .A2(n14948), .ZN(n14949) );
  AND2_X1 U16611 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n14950), .ZN(P2_U3266) );
  AND2_X1 U16612 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n14950), .ZN(P2_U3267) );
  AND2_X1 U16613 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n14950), .ZN(P2_U3268) );
  AND2_X1 U16614 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n14950), .ZN(P2_U3269) );
  AND2_X1 U16615 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n14950), .ZN(P2_U3270) );
  AND2_X1 U16616 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n14950), .ZN(P2_U3271) );
  INV_X1 U16617 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n15303) );
  NOR2_X1 U16618 ( .A1(n14949), .A2(n15303), .ZN(P2_U3272) );
  AND2_X1 U16619 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n14950), .ZN(P2_U3273) );
  AND2_X1 U16620 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n14950), .ZN(P2_U3274) );
  AND2_X1 U16621 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n14950), .ZN(P2_U3275) );
  AND2_X1 U16622 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n14950), .ZN(P2_U3276) );
  INV_X1 U16623 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n15227) );
  NOR2_X1 U16624 ( .A1(n14949), .A2(n15227), .ZN(P2_U3277) );
  AND2_X1 U16625 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n14950), .ZN(P2_U3278) );
  AND2_X1 U16626 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n14950), .ZN(P2_U3279) );
  AND2_X1 U16627 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n14950), .ZN(P2_U3280) );
  AND2_X1 U16628 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n14950), .ZN(P2_U3281) );
  AND2_X1 U16629 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n14950), .ZN(P2_U3282) );
  AND2_X1 U16630 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n14950), .ZN(P2_U3283) );
  AND2_X1 U16631 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n14950), .ZN(P2_U3284) );
  AND2_X1 U16632 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n14950), .ZN(P2_U3285) );
  AND2_X1 U16633 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n14950), .ZN(P2_U3286) );
  AND2_X1 U16634 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n14950), .ZN(P2_U3287) );
  INV_X1 U16635 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n15278) );
  NOR2_X1 U16636 ( .A1(n14949), .A2(n15278), .ZN(P2_U3288) );
  INV_X1 U16637 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n15249) );
  NOR2_X1 U16638 ( .A1(n14949), .A2(n15249), .ZN(P2_U3289) );
  AND2_X1 U16639 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n14950), .ZN(P2_U3290) );
  AND2_X1 U16640 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n14950), .ZN(P2_U3291) );
  AND2_X1 U16641 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n14950), .ZN(P2_U3292) );
  INV_X1 U16642 ( .A(P2_D_REG_4__SCAN_IN), .ZN(n15402) );
  NOR2_X1 U16643 ( .A1(n14949), .A2(n15402), .ZN(P2_U3293) );
  AND2_X1 U16644 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n14950), .ZN(P2_U3294) );
  AND2_X1 U16645 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n14950), .ZN(P2_U3295) );
  AOI22_X1 U16646 ( .A1(n14953), .A2(n14952), .B1(n14951), .B2(n14956), .ZN(
        P2_U3416) );
  INV_X1 U16647 ( .A(n14954), .ZN(n14955) );
  AOI21_X1 U16648 ( .B1(n14957), .B2(n14956), .A(n14955), .ZN(P2_U3417) );
  OAI211_X1 U16649 ( .C1(n14970), .C2(n14960), .A(n14959), .B(n14958), .ZN(
        n14961) );
  INV_X1 U16650 ( .A(n14961), .ZN(n15009) );
  AOI22_X1 U16651 ( .A1(n15007), .A2(n15009), .B1(n9162), .B2(n15005), .ZN(
        P2_U3430) );
  INV_X1 U16652 ( .A(n14967), .ZN(n14969) );
  AOI211_X1 U16653 ( .C1(n14965), .C2(n6721), .A(n14963), .B(n14962), .ZN(
        n14966) );
  OAI21_X1 U16654 ( .B1(n14970), .B2(n14967), .A(n14966), .ZN(n14968) );
  AOI21_X1 U16655 ( .B1(n14978), .B2(n14969), .A(n14968), .ZN(n15010) );
  AOI22_X1 U16656 ( .A1(n15007), .A2(n15010), .B1(n9218), .B2(n15005), .ZN(
        P2_U3445) );
  NOR2_X1 U16657 ( .A1(n14971), .A2(n14970), .ZN(n14976) );
  OAI211_X1 U16658 ( .C1(n14974), .C2(n14999), .A(n14973), .B(n14972), .ZN(
        n14975) );
  AOI211_X1 U16659 ( .C1(n14978), .C2(n14977), .A(n14976), .B(n14975), .ZN(
        n15012) );
  AOI22_X1 U16660 ( .A1(n15007), .A2(n15012), .B1(n9231), .B2(n15005), .ZN(
        P2_U3448) );
  OAI211_X1 U16661 ( .C1(n14981), .C2(n14999), .A(n14980), .B(n14979), .ZN(
        n14982) );
  AOI21_X1 U16662 ( .B1(n14984), .B2(n14983), .A(n14982), .ZN(n15014) );
  AOI22_X1 U16663 ( .A1(n15007), .A2(n15014), .B1(n9246), .B2(n15005), .ZN(
        P2_U3451) );
  INV_X1 U16664 ( .A(n14985), .ZN(n14989) );
  OAI21_X1 U16665 ( .B1(n7191), .B2(n14999), .A(n14986), .ZN(n14988) );
  AOI211_X1 U16666 ( .C1(n15004), .C2(n14989), .A(n14988), .B(n14987), .ZN(
        n15015) );
  INV_X1 U16667 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n14990) );
  AOI22_X1 U16668 ( .A1(n15007), .A2(n15015), .B1(n14990), .B2(n15005), .ZN(
        P2_U3454) );
  INV_X1 U16669 ( .A(n14991), .ZN(n14995) );
  OAI21_X1 U16670 ( .B1(n6979), .B2(n14999), .A(n14992), .ZN(n14994) );
  AOI211_X1 U16671 ( .C1(n15004), .C2(n14995), .A(n14994), .B(n14993), .ZN(
        n15016) );
  INV_X1 U16672 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n14996) );
  AOI22_X1 U16673 ( .A1(n15007), .A2(n15016), .B1(n14996), .B2(n15005), .ZN(
        P2_U3457) );
  INV_X1 U16674 ( .A(n14997), .ZN(n15003) );
  OAI21_X1 U16675 ( .B1(n15000), .B2(n14999), .A(n14998), .ZN(n15002) );
  AOI211_X1 U16676 ( .C1(n15004), .C2(n15003), .A(n15002), .B(n15001), .ZN(
        n15018) );
  INV_X1 U16677 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n15006) );
  AOI22_X1 U16678 ( .A1(n15007), .A2(n15018), .B1(n15006), .B2(n15005), .ZN(
        P2_U3460) );
  INV_X1 U16679 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n15008) );
  AOI22_X1 U16680 ( .A1(n15019), .A2(n15009), .B1(n15008), .B2(n15017), .ZN(
        P2_U3499) );
  AOI22_X1 U16681 ( .A1(n15019), .A2(n15010), .B1(n9219), .B2(n15017), .ZN(
        P2_U3504) );
  AOI22_X1 U16682 ( .A1(n15019), .A2(n15012), .B1(n15011), .B2(n15017), .ZN(
        P2_U3505) );
  AOI22_X1 U16683 ( .A1(n15019), .A2(n15014), .B1(n15013), .B2(n15017), .ZN(
        P2_U3506) );
  AOI22_X1 U16684 ( .A1(n15019), .A2(n15015), .B1(n9261), .B2(n15017), .ZN(
        P2_U3507) );
  AOI22_X1 U16685 ( .A1(n15019), .A2(n15016), .B1(n9273), .B2(n15017), .ZN(
        P2_U3508) );
  AOI22_X1 U16686 ( .A1(n15019), .A2(n15018), .B1(n10109), .B2(n15017), .ZN(
        P2_U3509) );
  NOR2_X1 U16687 ( .A1(P3_U3897), .A2(n15106), .ZN(P3_U3150) );
  NOR3_X1 U16688 ( .A1(n15023), .A2(n15109), .A3(n15085), .ZN(n15035) );
  INV_X1 U16689 ( .A(n15020), .ZN(n15021) );
  AOI22_X1 U16690 ( .A1(n15023), .A2(n15022), .B1(n15109), .B2(n15021), .ZN(
        n15033) );
  NAND2_X1 U16691 ( .A1(n15085), .A2(n8550), .ZN(n15026) );
  INV_X1 U16692 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n15024) );
  OAI22_X1 U16693 ( .A1(n15026), .A2(n15025), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n15024), .ZN(n15030) );
  NOR2_X1 U16694 ( .A1(n15028), .A2(n15027), .ZN(n15029) );
  AOI211_X1 U16695 ( .C1(n15031), .C2(n15507), .A(n15030), .B(n15029), .ZN(
        n15032) );
  OAI211_X1 U16696 ( .C1(n15035), .C2(n15034), .A(n15033), .B(n15032), .ZN(
        P3_U3182) );
  AOI21_X1 U16697 ( .B1(n10869), .B2(n15037), .A(n15036), .ZN(n15052) );
  NAND2_X1 U16698 ( .A1(n15039), .A2(n15038), .ZN(n15041) );
  OAI21_X1 U16699 ( .B1(n15042), .B2(n15041), .A(n15040), .ZN(n15047) );
  AOI21_X1 U16700 ( .B1(n15106), .B2(P3_ADDR_REG_3__SCAN_IN), .A(n15043), .ZN(
        n15044) );
  OAI21_X1 U16701 ( .B1(n15100), .B2(n15045), .A(n15044), .ZN(n15046) );
  AOI21_X1 U16702 ( .B1(n15047), .B2(n15085), .A(n15046), .ZN(n15051) );
  XNOR2_X1 U16703 ( .A(n15048), .B(P3_REG1_REG_3__SCAN_IN), .ZN(n15049) );
  NAND2_X1 U16704 ( .A1(n15109), .A2(n15049), .ZN(n15050) );
  OAI211_X1 U16705 ( .C1(n15052), .C2(n15113), .A(n15051), .B(n15050), .ZN(
        P3_U3185) );
  AOI21_X1 U16706 ( .B1(n15055), .B2(n15054), .A(n15053), .ZN(n15072) );
  OAI21_X1 U16707 ( .B1(n15058), .B2(n15057), .A(n15056), .ZN(n15063) );
  AOI21_X1 U16708 ( .B1(n15106), .B2(P3_ADDR_REG_4__SCAN_IN), .A(n15059), .ZN(
        n15060) );
  OAI21_X1 U16709 ( .B1(n15100), .B2(n15061), .A(n15060), .ZN(n15062) );
  AOI21_X1 U16710 ( .B1(n15063), .B2(n15085), .A(n15062), .ZN(n15071) );
  INV_X1 U16711 ( .A(n15064), .ZN(n15065) );
  AOI21_X1 U16712 ( .B1(n15067), .B2(n15066), .A(n15065), .ZN(n15068) );
  OR2_X1 U16713 ( .A1(n15069), .A2(n15068), .ZN(n15070) );
  OAI211_X1 U16714 ( .C1(n15072), .C2(n15113), .A(n15071), .B(n15070), .ZN(
        P3_U3186) );
  INV_X1 U16715 ( .A(n15073), .ZN(n15074) );
  AOI21_X1 U16716 ( .B1(n8603), .B2(n15075), .A(n15074), .ZN(n15091) );
  INV_X1 U16717 ( .A(n15076), .ZN(n15077) );
  NOR2_X1 U16718 ( .A1(n15078), .A2(n15077), .ZN(n15079) );
  XNOR2_X1 U16719 ( .A(n15080), .B(n15079), .ZN(n15086) );
  AOI21_X1 U16720 ( .B1(n15106), .B2(P3_ADDR_REG_5__SCAN_IN), .A(n15081), .ZN(
        n15082) );
  OAI21_X1 U16721 ( .B1(n15100), .B2(n15083), .A(n15082), .ZN(n15084) );
  AOI21_X1 U16722 ( .B1(n15086), .B2(n15085), .A(n15084), .ZN(n15090) );
  XNOR2_X1 U16723 ( .A(n15087), .B(P3_REG1_REG_5__SCAN_IN), .ZN(n15088) );
  NAND2_X1 U16724 ( .A1(n15109), .A2(n15088), .ZN(n15089) );
  OAI211_X1 U16725 ( .C1(n15091), .C2(n15113), .A(n15090), .B(n15089), .ZN(
        P3_U3187) );
  AOI21_X1 U16726 ( .B1(n15444), .B2(n15093), .A(n15092), .ZN(n15114) );
  INV_X1 U16727 ( .A(n15094), .ZN(n15099) );
  AOI21_X1 U16728 ( .B1(n15096), .B2(n15098), .A(n15095), .ZN(n15097) );
  AOI21_X1 U16729 ( .B1(n15099), .B2(n15098), .A(n15097), .ZN(n15103) );
  OAI22_X1 U16730 ( .A1(n15103), .A2(n15102), .B1(n15101), .B2(n15100), .ZN(
        n15104) );
  AOI211_X1 U16731 ( .C1(P3_ADDR_REG_9__SCAN_IN), .C2(n15106), .A(n15105), .B(
        n15104), .ZN(n15112) );
  OAI21_X1 U16732 ( .B1(P3_REG1_REG_9__SCAN_IN), .B2(n15108), .A(n15107), .ZN(
        n15110) );
  NAND2_X1 U16733 ( .A1(n15110), .A2(n15109), .ZN(n15111) );
  OAI211_X1 U16734 ( .C1(n15114), .C2(n15113), .A(n15112), .B(n15111), .ZN(
        P3_U3191) );
  XNOR2_X1 U16735 ( .A(n15116), .B(n15115), .ZN(n15129) );
  INV_X1 U16736 ( .A(n15129), .ZN(n15160) );
  NOR2_X1 U16737 ( .A1(n15117), .A2(n15200), .ZN(n15159) );
  INV_X1 U16738 ( .A(n15159), .ZN(n15119) );
  OAI22_X1 U16739 ( .A1(n15119), .A2(n15134), .B1(n10418), .B2(n15118), .ZN(
        n15130) );
  AOI22_X1 U16740 ( .A1(n15139), .A2(n15121), .B1(n15120), .B2(n15136), .ZN(
        n15128) );
  INV_X1 U16741 ( .A(n15122), .ZN(n15126) );
  AND3_X1 U16742 ( .A1(n15140), .A2(n15124), .A3(n15123), .ZN(n15125) );
  OAI21_X1 U16743 ( .B1(n15126), .B2(n15125), .A(n15143), .ZN(n15127) );
  OAI211_X1 U16744 ( .C1(n15129), .C2(n15147), .A(n15128), .B(n15127), .ZN(
        n15158) );
  AOI211_X1 U16745 ( .C1(n15131), .C2(n15160), .A(n15130), .B(n15158), .ZN(
        n15133) );
  AOI22_X1 U16746 ( .A1(n13074), .A2(n10859), .B1(n15133), .B2(n15132), .ZN(
        P3_U3231) );
  NOR2_X1 U16747 ( .A1(n8551), .A2(n15200), .ZN(n15155) );
  INV_X1 U16748 ( .A(n15134), .ZN(n15148) );
  XNOR2_X1 U16749 ( .A(n15135), .B(n15142), .ZN(n15149) );
  AOI22_X1 U16750 ( .A1(n15139), .A2(n15138), .B1(n15137), .B2(n15136), .ZN(
        n15146) );
  OAI21_X1 U16751 ( .B1(n15142), .B2(n15141), .A(n15140), .ZN(n15144) );
  NAND2_X1 U16752 ( .A1(n15144), .A2(n15143), .ZN(n15145) );
  OAI211_X1 U16753 ( .C1(n15149), .C2(n15147), .A(n15146), .B(n15145), .ZN(
        n15154) );
  AOI21_X1 U16754 ( .B1(n15155), .B2(n15148), .A(n15154), .ZN(n15153) );
  INV_X1 U16755 ( .A(n15149), .ZN(n15156) );
  AOI22_X1 U16756 ( .A1(n15156), .A2(n15151), .B1(P3_REG3_REG_1__SCAN_IN), 
        .B2(n15150), .ZN(n15152) );
  OAI221_X1 U16757 ( .B1(n13074), .B2(n15153), .C1(n15132), .C2(n10219), .A(
        n15152), .ZN(P3_U3232) );
  INV_X1 U16758 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n15157) );
  AOI211_X1 U16759 ( .C1(n15165), .C2(n15156), .A(n15155), .B(n15154), .ZN(
        n15207) );
  AOI22_X1 U16760 ( .A1(n15206), .A2(n15157), .B1(n15207), .B2(n15205), .ZN(
        P3_U3393) );
  INV_X1 U16761 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n15404) );
  AOI211_X1 U16762 ( .C1(n15160), .C2(n15165), .A(n15159), .B(n15158), .ZN(
        n15208) );
  AOI22_X1 U16763 ( .A1(n15206), .A2(n15404), .B1(n15208), .B2(n15205), .ZN(
        P3_U3396) );
  INV_X1 U16764 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n15166) );
  NOR2_X1 U16765 ( .A1(n15161), .A2(n15200), .ZN(n15163) );
  AOI211_X1 U16766 ( .C1(n15165), .C2(n15164), .A(n15163), .B(n15162), .ZN(
        n15209) );
  AOI22_X1 U16767 ( .A1(n15206), .A2(n15166), .B1(n15209), .B2(n15205), .ZN(
        P3_U3399) );
  INV_X1 U16768 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n15172) );
  INV_X1 U16769 ( .A(n15167), .ZN(n15169) );
  OAI22_X1 U16770 ( .A1(n15169), .A2(n15194), .B1(n15200), .B2(n15168), .ZN(
        n15170) );
  NOR2_X1 U16771 ( .A1(n15171), .A2(n15170), .ZN(n15211) );
  AOI22_X1 U16772 ( .A1(n15206), .A2(n15172), .B1(n15211), .B2(n15205), .ZN(
        P3_U3402) );
  INV_X1 U16773 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n15177) );
  OAI22_X1 U16774 ( .A1(n15174), .A2(n15194), .B1(n15200), .B2(n15173), .ZN(
        n15176) );
  NOR2_X1 U16775 ( .A1(n15176), .A2(n15175), .ZN(n15212) );
  AOI22_X1 U16776 ( .A1(n15206), .A2(n15177), .B1(n15212), .B2(n15205), .ZN(
        P3_U3405) );
  INV_X1 U16777 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n15182) );
  OAI22_X1 U16778 ( .A1(n15179), .A2(n15194), .B1(n15178), .B2(n15200), .ZN(
        n15181) );
  NOR2_X1 U16779 ( .A1(n15181), .A2(n15180), .ZN(n15214) );
  AOI22_X1 U16780 ( .A1(n15206), .A2(n15182), .B1(n15214), .B2(n15205), .ZN(
        P3_U3408) );
  INV_X1 U16781 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n15187) );
  OAI22_X1 U16782 ( .A1(n15184), .A2(n15194), .B1(n15200), .B2(n15183), .ZN(
        n15186) );
  NOR2_X1 U16783 ( .A1(n15186), .A2(n15185), .ZN(n15216) );
  AOI22_X1 U16784 ( .A1(n15206), .A2(n15187), .B1(n15216), .B2(n15205), .ZN(
        P3_U3411) );
  INV_X1 U16785 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n15192) );
  OAI22_X1 U16786 ( .A1(n15189), .A2(n15194), .B1(n15188), .B2(n15200), .ZN(
        n15190) );
  NOR2_X1 U16787 ( .A1(n15191), .A2(n15190), .ZN(n15218) );
  AOI22_X1 U16788 ( .A1(n15206), .A2(n15192), .B1(n15218), .B2(n15205), .ZN(
        P3_U3414) );
  INV_X1 U16789 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n15198) );
  OAI22_X1 U16790 ( .A1(n15195), .A2(n15194), .B1(n15200), .B2(n15193), .ZN(
        n15196) );
  NOR2_X1 U16791 ( .A1(n15197), .A2(n15196), .ZN(n15220) );
  AOI22_X1 U16792 ( .A1(n15206), .A2(n15198), .B1(n15220), .B2(n15205), .ZN(
        P3_U3417) );
  INV_X1 U16793 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n15453) );
  OAI22_X1 U16794 ( .A1(n15202), .A2(n15201), .B1(n15200), .B2(n15199), .ZN(
        n15203) );
  NOR2_X1 U16795 ( .A1(n15204), .A2(n15203), .ZN(n15221) );
  AOI22_X1 U16796 ( .A1(n15206), .A2(n15453), .B1(n15221), .B2(n15205), .ZN(
        P3_U3420) );
  AOI22_X1 U16797 ( .A1(n15222), .A2(n15207), .B1(n10331), .B2(n9126), .ZN(
        P3_U3460) );
  AOI22_X1 U16798 ( .A1(n15222), .A2(n15208), .B1(n10225), .B2(n9126), .ZN(
        P3_U3461) );
  AOI22_X1 U16799 ( .A1(n15222), .A2(n15209), .B1(n10868), .B2(n9126), .ZN(
        P3_U3462) );
  AOI22_X1 U16800 ( .A1(n15222), .A2(n15211), .B1(n15210), .B2(n9126), .ZN(
        P3_U3463) );
  AOI22_X1 U16801 ( .A1(n15222), .A2(n15212), .B1(n6740), .B2(n9126), .ZN(
        P3_U3464) );
  AOI22_X1 U16802 ( .A1(n15222), .A2(n15214), .B1(n15213), .B2(n9126), .ZN(
        P3_U3465) );
  INV_X1 U16803 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n15215) );
  AOI22_X1 U16804 ( .A1(n15222), .A2(n15216), .B1(n15215), .B2(n9126), .ZN(
        P3_U3466) );
  AOI22_X1 U16805 ( .A1(n15222), .A2(n15218), .B1(n15217), .B2(n9126), .ZN(
        P3_U3467) );
  INV_X1 U16806 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n15219) );
  AOI22_X1 U16807 ( .A1(n15222), .A2(n15220), .B1(n15219), .B2(n9126), .ZN(
        P3_U3468) );
  AOI22_X1 U16808 ( .A1(n15222), .A2(n15221), .B1(n10885), .B2(n9126), .ZN(
        P3_U3469) );
  NAND2_X1 U16809 ( .A1(n15223), .A2(P3_U3897), .ZN(n15224) );
  OAI21_X1 U16810 ( .B1(P3_U3897), .B2(P3_DATAO_REG_28__SCAN_IN), .A(n15224), 
        .ZN(n15432) );
  AOI22_X1 U16811 ( .A1(n15485), .A2(keyinput46), .B1(keyinput70), .B2(n15226), 
        .ZN(n15225) );
  OAI221_X1 U16812 ( .B1(n15485), .B2(keyinput46), .C1(n15226), .C2(keyinput70), .A(n15225), .ZN(n15236) );
  XNOR2_X1 U16813 ( .A(n15227), .B(keyinput6), .ZN(n15235) );
  XNOR2_X1 U16814 ( .A(n15228), .B(keyinput44), .ZN(n15234) );
  XOR2_X1 U16815 ( .A(n9206), .B(keyinput11), .Z(n15232) );
  XNOR2_X1 U16816 ( .A(P2_RD_REG_SCAN_IN), .B(keyinput109), .ZN(n15231) );
  XNOR2_X1 U16817 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput7), .ZN(n15230) );
  XNOR2_X1 U16818 ( .A(P1_IR_REG_29__SCAN_IN), .B(keyinput21), .ZN(n15229) );
  NAND4_X1 U16819 ( .A1(n15232), .A2(n15231), .A3(n15230), .A4(n15229), .ZN(
        n15233) );
  NOR4_X1 U16820 ( .A1(n15236), .A2(n15235), .A3(n15234), .A4(n15233), .ZN(
        n15276) );
  INV_X1 U16821 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n15238) );
  AOI22_X1 U16822 ( .A1(n15470), .A2(keyinput101), .B1(n15238), .B2(keyinput32), .ZN(n15237) );
  OAI221_X1 U16823 ( .B1(n15470), .B2(keyinput101), .C1(n15238), .C2(
        keyinput32), .A(n15237), .ZN(n15247) );
  AOI22_X1 U16824 ( .A1(n9273), .A2(keyinput95), .B1(keyinput17), .B2(n15240), 
        .ZN(n15239) );
  OAI221_X1 U16825 ( .B1(n9273), .B2(keyinput95), .C1(n15240), .C2(keyinput17), 
        .A(n15239), .ZN(n15246) );
  AOI22_X1 U16826 ( .A1(n15486), .A2(keyinput123), .B1(keyinput86), .B2(n15242), .ZN(n15241) );
  OAI221_X1 U16827 ( .B1(n15486), .B2(keyinput123), .C1(n15242), .C2(
        keyinput86), .A(n15241), .ZN(n15245) );
  AOI22_X1 U16828 ( .A1(n15464), .A2(keyinput50), .B1(n13541), .B2(keyinput53), 
        .ZN(n15243) );
  OAI221_X1 U16829 ( .B1(n15464), .B2(keyinput50), .C1(n13541), .C2(keyinput53), .A(n15243), .ZN(n15244) );
  NOR4_X1 U16830 ( .A1(n15247), .A2(n15246), .A3(n15245), .A4(n15244), .ZN(
        n15275) );
  AOI22_X1 U16831 ( .A1(n6740), .A2(keyinput103), .B1(keyinput27), .B2(n15249), 
        .ZN(n15248) );
  OAI221_X1 U16832 ( .B1(n6740), .B2(keyinput103), .C1(n15249), .C2(keyinput27), .A(n15248), .ZN(n15260) );
  AOI22_X1 U16833 ( .A1(n15252), .A2(keyinput68), .B1(keyinput98), .B2(n15251), 
        .ZN(n15250) );
  OAI221_X1 U16834 ( .B1(n15252), .B2(keyinput68), .C1(n15251), .C2(keyinput98), .A(n15250), .ZN(n15259) );
  AOI22_X1 U16835 ( .A1(n9395), .A2(keyinput91), .B1(n15254), .B2(keyinput59), 
        .ZN(n15253) );
  OAI221_X1 U16836 ( .B1(n9395), .B2(keyinput91), .C1(n15254), .C2(keyinput59), 
        .A(n15253), .ZN(n15258) );
  INV_X1 U16837 ( .A(P3_REG3_REG_26__SCAN_IN), .ZN(n15256) );
  AOI22_X1 U16838 ( .A1(n15256), .A2(keyinput56), .B1(keyinput45), .B2(n10027), 
        .ZN(n15255) );
  OAI221_X1 U16839 ( .B1(n15256), .B2(keyinput56), .C1(n10027), .C2(keyinput45), .A(n15255), .ZN(n15257) );
  NOR4_X1 U16840 ( .A1(n15260), .A2(n15259), .A3(n15258), .A4(n15257), .ZN(
        n15274) );
  AOI22_X1 U16841 ( .A1(n15262), .A2(keyinput114), .B1(keyinput66), .B2(n15442), .ZN(n15261) );
  OAI221_X1 U16842 ( .B1(n15262), .B2(keyinput114), .C1(n15442), .C2(
        keyinput66), .A(n15261), .ZN(n15272) );
  AOI22_X1 U16843 ( .A1(n15265), .A2(keyinput39), .B1(keyinput61), .B2(n15264), 
        .ZN(n15263) );
  OAI221_X1 U16844 ( .B1(n15265), .B2(keyinput39), .C1(n15264), .C2(keyinput61), .A(n15263), .ZN(n15271) );
  XOR2_X1 U16845 ( .A(n9150), .B(keyinput87), .Z(n15269) );
  XNOR2_X1 U16846 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(keyinput67), .ZN(n15268)
         );
  XNOR2_X1 U16847 ( .A(P2_REG3_REG_20__SCAN_IN), .B(keyinput78), .ZN(n15267)
         );
  XNOR2_X1 U16848 ( .A(P3_IR_REG_10__SCAN_IN), .B(keyinput124), .ZN(n15266) );
  NAND4_X1 U16849 ( .A1(n15269), .A2(n15268), .A3(n15267), .A4(n15266), .ZN(
        n15270) );
  NOR3_X1 U16850 ( .A1(n15272), .A2(n15271), .A3(n15270), .ZN(n15273) );
  NAND4_X1 U16851 ( .A1(n15276), .A2(n15275), .A3(n15274), .A4(n15273), .ZN(
        n15430) );
  AOI22_X1 U16852 ( .A1(n15469), .A2(keyinput72), .B1(n15278), .B2(keyinput107), .ZN(n15277) );
  OAI221_X1 U16853 ( .B1(n15469), .B2(keyinput72), .C1(n15278), .C2(
        keyinput107), .A(n15277), .ZN(n15288) );
  AOI22_X1 U16854 ( .A1(n15281), .A2(keyinput75), .B1(keyinput84), .B2(n15280), 
        .ZN(n15279) );
  OAI221_X1 U16855 ( .B1(n15281), .B2(keyinput75), .C1(n15280), .C2(keyinput84), .A(n15279), .ZN(n15287) );
  AOI22_X1 U16856 ( .A1(n15492), .A2(keyinput64), .B1(keyinput85), .B2(n13390), 
        .ZN(n15282) );
  OAI221_X1 U16857 ( .B1(n15492), .B2(keyinput64), .C1(n13390), .C2(keyinput85), .A(n15282), .ZN(n15286) );
  AOI22_X1 U16858 ( .A1(n7763), .A2(keyinput12), .B1(n15284), .B2(keyinput35), 
        .ZN(n15283) );
  OAI221_X1 U16859 ( .B1(n7763), .B2(keyinput12), .C1(n15284), .C2(keyinput35), 
        .A(n15283), .ZN(n15285) );
  NOR4_X1 U16860 ( .A1(n15288), .A2(n15287), .A3(n15286), .A4(n15285), .ZN(
        n15324) );
  AOI22_X1 U16861 ( .A1(n8524), .A2(keyinput126), .B1(keyinput92), .B2(n15523), 
        .ZN(n15289) );
  OAI221_X1 U16862 ( .B1(n8524), .B2(keyinput126), .C1(n15523), .C2(keyinput92), .A(n15289), .ZN(n15300) );
  AOI22_X1 U16863 ( .A1(n9173), .A2(keyinput76), .B1(n13767), .B2(keyinput111), 
        .ZN(n15290) );
  OAI221_X1 U16864 ( .B1(n9173), .B2(keyinput76), .C1(n13767), .C2(keyinput111), .A(n15290), .ZN(n15299) );
  AOI22_X1 U16865 ( .A1(n15293), .A2(keyinput73), .B1(n15292), .B2(keyinput79), 
        .ZN(n15291) );
  OAI221_X1 U16866 ( .B1(n15293), .B2(keyinput73), .C1(n15292), .C2(keyinput79), .A(n15291), .ZN(n15298) );
  XOR2_X1 U16867 ( .A(n15294), .B(keyinput99), .Z(n15296) );
  XNOR2_X1 U16868 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(keyinput41), .ZN(n15295)
         );
  NAND2_X1 U16869 ( .A1(n15296), .A2(n15295), .ZN(n15297) );
  NOR4_X1 U16870 ( .A1(n15300), .A2(n15299), .A3(n15298), .A4(n15297), .ZN(
        n15323) );
  AOI22_X1 U16871 ( .A1(n15461), .A2(keyinput88), .B1(keyinput22), .B2(n15460), 
        .ZN(n15301) );
  OAI221_X1 U16872 ( .B1(n15461), .B2(keyinput88), .C1(n15460), .C2(keyinput22), .A(n15301), .ZN(n15310) );
  AOI22_X1 U16873 ( .A1(n9526), .A2(keyinput113), .B1(n15303), .B2(keyinput117), .ZN(n15302) );
  OAI221_X1 U16874 ( .B1(n9526), .B2(keyinput113), .C1(n15303), .C2(
        keyinput117), .A(n15302), .ZN(n15309) );
  INV_X1 U16875 ( .A(P3_REG2_REG_20__SCAN_IN), .ZN(n15489) );
  AOI22_X1 U16876 ( .A1(n12197), .A2(keyinput31), .B1(n15489), .B2(keyinput23), 
        .ZN(n15304) );
  OAI221_X1 U16877 ( .B1(n12197), .B2(keyinput31), .C1(n15489), .C2(keyinput23), .A(n15304), .ZN(n15308) );
  XOR2_X1 U16878 ( .A(n9922), .B(keyinput120), .Z(n15306) );
  XNOR2_X1 U16879 ( .A(P1_IR_REG_25__SCAN_IN), .B(keyinput71), .ZN(n15305) );
  NAND2_X1 U16880 ( .A1(n15306), .A2(n15305), .ZN(n15307) );
  NOR4_X1 U16881 ( .A1(n15310), .A2(n15309), .A3(n15308), .A4(n15307), .ZN(
        n15322) );
  AOI22_X1 U16882 ( .A1(n15312), .A2(keyinput30), .B1(keyinput2), .B2(n15495), 
        .ZN(n15311) );
  OAI221_X1 U16883 ( .B1(n15312), .B2(keyinput30), .C1(n15495), .C2(keyinput2), 
        .A(n15311), .ZN(n15320) );
  AOI22_X1 U16884 ( .A1(n8925), .A2(keyinput42), .B1(keyinput58), .B2(n9159), 
        .ZN(n15313) );
  OAI221_X1 U16885 ( .B1(n8925), .B2(keyinput42), .C1(n9159), .C2(keyinput58), 
        .A(n15313), .ZN(n15319) );
  AOI22_X1 U16886 ( .A1(n15473), .A2(keyinput100), .B1(n11010), .B2(keyinput81), .ZN(n15314) );
  OAI221_X1 U16887 ( .B1(n15473), .B2(keyinput100), .C1(n11010), .C2(
        keyinput81), .A(n15314), .ZN(n15318) );
  XNOR2_X1 U16888 ( .A(P2_IR_REG_15__SCAN_IN), .B(keyinput28), .ZN(n15316) );
  XNOR2_X1 U16889 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(keyinput1), .ZN(n15315)
         );
  NAND2_X1 U16890 ( .A1(n15316), .A2(n15315), .ZN(n15317) );
  NOR4_X1 U16891 ( .A1(n15320), .A2(n15319), .A3(n15318), .A4(n15317), .ZN(
        n15321) );
  NAND4_X1 U16892 ( .A1(n15324), .A2(n15323), .A3(n15322), .A4(n15321), .ZN(
        n15429) );
  AOI22_X1 U16893 ( .A1(n15327), .A2(keyinput9), .B1(keyinput119), .B2(n15326), 
        .ZN(n15325) );
  OAI221_X1 U16894 ( .B1(n15327), .B2(keyinput9), .C1(n15326), .C2(keyinput119), .A(n15325), .ZN(n15337) );
  AOI22_X1 U16895 ( .A1(n15329), .A2(keyinput108), .B1(n15459), .B2(keyinput60), .ZN(n15328) );
  OAI221_X1 U16896 ( .B1(n15329), .B2(keyinput108), .C1(n15459), .C2(
        keyinput60), .A(n15328), .ZN(n15336) );
  INV_X1 U16897 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n15451) );
  AOI22_X1 U16898 ( .A1(n15488), .A2(keyinput63), .B1(n15451), .B2(keyinput13), 
        .ZN(n15330) );
  OAI221_X1 U16899 ( .B1(n15488), .B2(keyinput63), .C1(n15451), .C2(keyinput13), .A(n15330), .ZN(n15335) );
  AOI22_X1 U16900 ( .A1(n15333), .A2(keyinput24), .B1(n15332), .B2(keyinput4), 
        .ZN(n15331) );
  OAI221_X1 U16901 ( .B1(n15333), .B2(keyinput24), .C1(n15332), .C2(keyinput4), 
        .A(n15331), .ZN(n15334) );
  NOR4_X1 U16902 ( .A1(n15337), .A2(n15336), .A3(n15335), .A4(n15334), .ZN(
        n15375) );
  AOI22_X1 U16903 ( .A1(n10986), .A2(keyinput0), .B1(n8955), .B2(keyinput16), 
        .ZN(n15338) );
  OAI221_X1 U16904 ( .B1(n10986), .B2(keyinput0), .C1(n8955), .C2(keyinput16), 
        .A(n15338), .ZN(n15346) );
  AOI22_X1 U16905 ( .A1(n15449), .A2(keyinput105), .B1(n11722), .B2(keyinput43), .ZN(n15339) );
  OAI221_X1 U16906 ( .B1(n15449), .B2(keyinput105), .C1(n11722), .C2(
        keyinput43), .A(n15339), .ZN(n15345) );
  AOI22_X1 U16907 ( .A1(n15450), .A2(keyinput104), .B1(keyinput37), .B2(n15453), .ZN(n15340) );
  OAI221_X1 U16908 ( .B1(n15450), .B2(keyinput104), .C1(n15453), .C2(
        keyinput37), .A(n15340), .ZN(n15344) );
  INV_X1 U16909 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n15342) );
  AOI22_X1 U16910 ( .A1(n15342), .A2(keyinput52), .B1(keyinput26), .B2(n15454), 
        .ZN(n15341) );
  OAI221_X1 U16911 ( .B1(n15342), .B2(keyinput52), .C1(n15454), .C2(keyinput26), .A(n15341), .ZN(n15343) );
  NOR4_X1 U16912 ( .A1(n15346), .A2(n15345), .A3(n15344), .A4(n15343), .ZN(
        n15374) );
  INV_X1 U16913 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n15348) );
  AOI22_X1 U16914 ( .A1(n15348), .A2(keyinput36), .B1(keyinput40), .B2(n14164), 
        .ZN(n15347) );
  OAI221_X1 U16915 ( .B1(n15348), .B2(keyinput36), .C1(n14164), .C2(keyinput40), .A(n15347), .ZN(n15353) );
  AOI22_X1 U16916 ( .A1(n15452), .A2(keyinput93), .B1(keyinput29), .B2(n13732), 
        .ZN(n15349) );
  OAI221_X1 U16917 ( .B1(n15452), .B2(keyinput93), .C1(n13732), .C2(keyinput29), .A(n15349), .ZN(n15352) );
  XNOR2_X1 U16918 ( .A(n15350), .B(keyinput82), .ZN(n15351) );
  OR3_X1 U16919 ( .A1(n15353), .A2(n15352), .A3(n15351), .ZN(n15359) );
  AOI22_X1 U16920 ( .A1(n15355), .A2(keyinput62), .B1(n11493), .B2(keyinput115), .ZN(n15354) );
  OAI221_X1 U16921 ( .B1(n15355), .B2(keyinput62), .C1(n11493), .C2(
        keyinput115), .A(n15354), .ZN(n15358) );
  XNOR2_X1 U16922 ( .A(n15356), .B(keyinput112), .ZN(n15357) );
  NOR3_X1 U16923 ( .A1(n15359), .A2(n15358), .A3(n15357), .ZN(n15373) );
  INV_X1 U16924 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n15361) );
  AOI22_X1 U16925 ( .A1(n15444), .A2(keyinput97), .B1(keyinput69), .B2(n15361), 
        .ZN(n15360) );
  OAI221_X1 U16926 ( .B1(n15444), .B2(keyinput97), .C1(n15361), .C2(keyinput69), .A(n15360), .ZN(n15371) );
  AOI22_X1 U16927 ( .A1(n15462), .A2(keyinput125), .B1(keyinput122), .B2(
        n15363), .ZN(n15362) );
  OAI221_X1 U16928 ( .B1(n15462), .B2(keyinput125), .C1(n15363), .C2(
        keyinput122), .A(n15362), .ZN(n15370) );
  AOI22_X1 U16929 ( .A1(n8550), .A2(keyinput89), .B1(keyinput77), .B2(n8938), 
        .ZN(n15364) );
  OAI221_X1 U16930 ( .B1(n8550), .B2(keyinput89), .C1(n8938), .C2(keyinput77), 
        .A(n15364), .ZN(n15369) );
  XOR2_X1 U16931 ( .A(n15365), .B(keyinput33), .Z(n15367) );
  XNOR2_X1 U16932 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput57), .ZN(n15366) );
  NAND2_X1 U16933 ( .A1(n15367), .A2(n15366), .ZN(n15368) );
  NOR4_X1 U16934 ( .A1(n15371), .A2(n15370), .A3(n15369), .A4(n15368), .ZN(
        n15372) );
  NAND4_X1 U16935 ( .A1(n15375), .A2(n15374), .A3(n15373), .A4(n15372), .ZN(
        n15428) );
  INV_X1 U16936 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n15508) );
  AOI22_X1 U16937 ( .A1(n15508), .A2(keyinput74), .B1(keyinput18), .B2(n7851), 
        .ZN(n15376) );
  OAI221_X1 U16938 ( .B1(n15508), .B2(keyinput74), .C1(n7851), .C2(keyinput18), 
        .A(n15376), .ZN(n15384) );
  AOI22_X1 U16939 ( .A1(n9329), .A2(keyinput51), .B1(n15435), .B2(keyinput54), 
        .ZN(n15377) );
  OAI221_X1 U16940 ( .B1(n9329), .B2(keyinput51), .C1(n15435), .C2(keyinput54), 
        .A(n15377), .ZN(n15383) );
  AOI22_X1 U16941 ( .A1(n11188), .A2(keyinput110), .B1(n15379), .B2(
        keyinput118), .ZN(n15378) );
  OAI221_X1 U16942 ( .B1(n11188), .B2(keyinput110), .C1(n15379), .C2(
        keyinput118), .A(n15378), .ZN(n15382) );
  AOI22_X1 U16943 ( .A1(n7389), .A2(keyinput55), .B1(keyinput10), .B2(n15434), 
        .ZN(n15380) );
  OAI221_X1 U16944 ( .B1(n7389), .B2(keyinput55), .C1(n15434), .C2(keyinput10), 
        .A(n15380), .ZN(n15381) );
  NOR4_X1 U16945 ( .A1(n15384), .A2(n15383), .A3(n15382), .A4(n15381), .ZN(
        n15426) );
  AOI22_X1 U16946 ( .A1(n15386), .A2(keyinput90), .B1(n7870), .B2(keyinput127), 
        .ZN(n15385) );
  OAI221_X1 U16947 ( .B1(n15386), .B2(keyinput90), .C1(n7870), .C2(keyinput127), .A(n15385), .ZN(n15398) );
  AOI22_X1 U16948 ( .A1(n15389), .A2(keyinput116), .B1(n15388), .B2(keyinput20), .ZN(n15387) );
  OAI221_X1 U16949 ( .B1(n15389), .B2(keyinput116), .C1(n15388), .C2(
        keyinput20), .A(n15387), .ZN(n15397) );
  AOI22_X1 U16950 ( .A1(n15433), .A2(keyinput102), .B1(n15391), .B2(keyinput34), .ZN(n15390) );
  OAI221_X1 U16951 ( .B1(n15433), .B2(keyinput102), .C1(n15391), .C2(
        keyinput34), .A(n15390), .ZN(n15396) );
  XOR2_X1 U16952 ( .A(n15392), .B(keyinput65), .Z(n15394) );
  XNOR2_X1 U16953 ( .A(P2_REG3_REG_6__SCAN_IN), .B(keyinput38), .ZN(n15393) );
  NAND2_X1 U16954 ( .A1(n15394), .A2(n15393), .ZN(n15395) );
  NOR4_X1 U16955 ( .A1(n15398), .A2(n15397), .A3(n15396), .A4(n15395), .ZN(
        n15425) );
  AOI22_X1 U16956 ( .A1(n9341), .A2(keyinput5), .B1(n15400), .B2(keyinput3), 
        .ZN(n15399) );
  OAI221_X1 U16957 ( .B1(n9341), .B2(keyinput5), .C1(n15400), .C2(keyinput3), 
        .A(n15399), .ZN(n15410) );
  AOI22_X1 U16958 ( .A1(n15402), .A2(keyinput80), .B1(keyinput19), .B2(n10922), 
        .ZN(n15401) );
  OAI221_X1 U16959 ( .B1(n15402), .B2(keyinput80), .C1(n10922), .C2(keyinput19), .A(n15401), .ZN(n15409) );
  AOI22_X1 U16960 ( .A1(n15404), .A2(keyinput106), .B1(keyinput121), .B2(
        n15465), .ZN(n15403) );
  OAI221_X1 U16961 ( .B1(n15404), .B2(keyinput106), .C1(n15465), .C2(
        keyinput121), .A(n15403), .ZN(n15408) );
  XNOR2_X1 U16962 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(keyinput96), .ZN(n15406)
         );
  XNOR2_X1 U16963 ( .A(P3_B_REG_SCAN_IN), .B(keyinput49), .ZN(n15405) );
  NAND2_X1 U16964 ( .A1(n15406), .A2(n15405), .ZN(n15407) );
  NOR4_X1 U16965 ( .A1(n15410), .A2(n15409), .A3(n15408), .A4(n15407), .ZN(
        n15424) );
  AOI22_X1 U16966 ( .A1(n15437), .A2(keyinput83), .B1(keyinput48), .B2(n10267), 
        .ZN(n15411) );
  OAI221_X1 U16967 ( .B1(n15437), .B2(keyinput83), .C1(n10267), .C2(keyinput48), .A(n15411), .ZN(n15422) );
  AOI22_X1 U16968 ( .A1(n15436), .A2(keyinput47), .B1(n15413), .B2(keyinput15), 
        .ZN(n15412) );
  OAI221_X1 U16969 ( .B1(n15436), .B2(keyinput47), .C1(n15413), .C2(keyinput15), .A(n15412), .ZN(n15421) );
  AOI22_X1 U16970 ( .A1(n15416), .A2(keyinput8), .B1(n15415), .B2(keyinput94), 
        .ZN(n15414) );
  OAI221_X1 U16971 ( .B1(n15416), .B2(keyinput8), .C1(n15415), .C2(keyinput94), 
        .A(n15414), .ZN(n15420) );
  AOI22_X1 U16972 ( .A1(n15418), .A2(keyinput14), .B1(n11991), .B2(keyinput25), 
        .ZN(n15417) );
  OAI221_X1 U16973 ( .B1(n15418), .B2(keyinput14), .C1(n11991), .C2(keyinput25), .A(n15417), .ZN(n15419) );
  NOR4_X1 U16974 ( .A1(n15422), .A2(n15421), .A3(n15420), .A4(n15419), .ZN(
        n15423) );
  NAND4_X1 U16975 ( .A1(n15426), .A2(n15425), .A3(n15424), .A4(n15423), .ZN(
        n15427) );
  NOR4_X1 U16976 ( .A1(n15430), .A2(n15429), .A3(n15428), .A4(n15427), .ZN(
        n15431) );
  XNOR2_X1 U16977 ( .A(n15432), .B(n15431), .ZN(n15519) );
  NOR4_X1 U16978 ( .A1(P1_REG3_REG_25__SCAN_IN), .A2(P1_REG3_REG_12__SCAN_IN), 
        .A3(n15434), .A4(n15433), .ZN(n15441) );
  NOR4_X1 U16979 ( .A1(P3_D_REG_9__SCAN_IN), .A2(n7389), .A3(n15435), .A4(
        n11188), .ZN(n15440) );
  NOR4_X1 U16980 ( .A1(SI_21_), .A2(P3_REG2_REG_29__SCAN_IN), .A3(
        P1_REG0_REG_18__SCAN_IN), .A4(n15436), .ZN(n15439) );
  NOR4_X1 U16981 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .A3(n15437), .A4(n9341), .ZN(n15438) );
  AND4_X1 U16982 ( .A1(n15441), .A2(n15440), .A3(n15439), .A4(n15438), .ZN(
        n15448) );
  NAND4_X1 U16983 ( .A1(P2_REG0_REG_1__SCAN_IN), .A2(P2_REG3_REG_20__SCAN_IN), 
        .A3(P3_DATAO_REG_11__SCAN_IN), .A4(n15442), .ZN(n15443) );
  NOR3_X1 U16984 ( .A1(P3_D_REG_14__SCAN_IN), .A2(P2_REG3_REG_1__SCAN_IN), 
        .A3(n15443), .ZN(n15447) );
  NAND4_X1 U16985 ( .A1(P3_REG2_REG_24__SCAN_IN), .A2(P3_REG0_REG_0__SCAN_IN), 
        .A3(P3_DATAO_REG_26__SCAN_IN), .A4(n15444), .ZN(n15445) );
  NOR3_X1 U16986 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(n9329), .A3(n15445), .ZN(
        n15446) );
  AND3_X1 U16987 ( .A1(n15448), .A2(n15447), .A3(n15446), .ZN(n15517) );
  NAND4_X1 U16988 ( .A1(P3_REG2_REG_25__SCAN_IN), .A2(n15450), .A3(n11722), 
        .A4(n15449), .ZN(n15458) );
  NAND4_X1 U16989 ( .A1(P2_REG2_REG_7__SCAN_IN), .A2(P1_DATAO_REG_29__SCAN_IN), 
        .A3(P1_REG1_REG_29__SCAN_IN), .A4(n15451), .ZN(n15457) );
  NAND4_X1 U16990 ( .A1(P3_REG1_REG_11__SCAN_IN), .A2(n15452), .A3(n11493), 
        .A4(n13732), .ZN(n15456) );
  NAND4_X1 U16991 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P1_REG2_REG_23__SCAN_IN), 
        .A3(n15454), .A4(n15453), .ZN(n15455) );
  NOR4_X1 U16992 ( .A1(n15458), .A2(n15457), .A3(n15456), .A4(n15455), .ZN(
        n15516) );
  NAND4_X1 U16993 ( .A1(n15462), .A2(n15461), .A3(n15460), .A4(n15459), .ZN(
        n15463) );
  NOR3_X1 U16994 ( .A1(P2_D_REG_20__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .A3(
        n15463), .ZN(n15515) );
  NAND4_X1 U16995 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P3_REG1_REG_5__SCAN_IN), 
        .A3(n13541), .A4(n15464), .ZN(n15467) );
  NAND4_X1 U16996 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P3_REG0_REG_2__SCAN_IN), 
        .A3(n15465), .A4(n10922), .ZN(n15466) );
  NOR3_X1 U16997 ( .A1(n15468), .A2(n15467), .A3(n15466), .ZN(n15513) );
  NAND4_X1 U16998 ( .A1(P2_D_REG_9__SCAN_IN), .A2(P2_DATAO_REG_10__SCAN_IN), 
        .A3(P1_REG1_REG_17__SCAN_IN), .A4(n15469), .ZN(n15472) );
  NAND4_X1 U16999 ( .A1(P1_IR_REG_29__SCAN_IN), .A2(P2_REG1_REG_4__SCAN_IN), 
        .A3(P3_DATAO_REG_17__SCAN_IN), .A4(n15470), .ZN(n15471) );
  NOR2_X1 U17000 ( .A1(n15472), .A2(n15471), .ZN(n15477) );
  NAND4_X1 U17001 ( .A1(P2_D_REG_25__SCAN_IN), .A2(SI_2_), .A3(
        P2_REG3_REG_3__SCAN_IN), .A4(n9526), .ZN(n15475) );
  NAND4_X1 U17002 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(n8925), .A3(n11010), .A4(
        n15473), .ZN(n15474) );
  NOR2_X1 U17003 ( .A1(n15475), .A2(n15474), .ZN(n15476) );
  AND2_X1 U17004 ( .A1(n15477), .A2(n15476), .ZN(n15512) );
  NAND4_X1 U17005 ( .A1(n15481), .A2(n15480), .A3(n15479), .A4(n15478), .ZN(
        n15483) );
  NAND4_X1 U17006 ( .A1(n7155), .A2(P1_DATAO_REG_25__SCAN_IN), .A3(
        P2_REG3_REG_6__SCAN_IN), .A4(P1_DATAO_REG_22__SCAN_IN), .ZN(n15482) );
  NOR2_X1 U17007 ( .A1(n15483), .A2(n15482), .ZN(n15506) );
  NAND4_X1 U17008 ( .A1(n15485), .A2(n15484), .A3(P3_IR_REG_8__SCAN_IN), .A4(
        P3_IR_REG_11__SCAN_IN), .ZN(n15500) );
  AND4_X1 U17009 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_REG1_REG_30__SCAN_IN), 
        .A3(n15486), .A4(n9273), .ZN(n15487) );
  AND2_X1 U17010 ( .A1(n15487), .A2(n13767), .ZN(n15496) );
  NAND4_X1 U17011 ( .A1(P2_REG1_REG_30__SCAN_IN), .A2(P2_REG1_REG_23__SCAN_IN), 
        .A3(P1_REG2_REG_0__SCAN_IN), .A4(n15488), .ZN(n15491) );
  NAND4_X1 U17012 ( .A1(P2_REG2_REG_30__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), 
        .A3(P1_REG1_REG_4__SCAN_IN), .A4(n15489), .ZN(n15490) );
  NOR2_X1 U17013 ( .A1(n15491), .A2(n15490), .ZN(n15494) );
  AND4_X1 U17014 ( .A1(P3_REG0_REG_21__SCAN_IN), .A2(P2_REG2_REG_17__SCAN_IN), 
        .A3(n15492), .A4(n7763), .ZN(n15493) );
  AND4_X1 U17015 ( .A1(n15496), .A2(n15495), .A3(n15494), .A4(n15493), .ZN(
        n15497) );
  NAND3_X1 U17016 ( .A1(n15498), .A2(P3_DATAO_REG_31__SCAN_IN), .A3(n15497), 
        .ZN(n15499) );
  NOR2_X1 U17017 ( .A1(n15500), .A2(n15499), .ZN(n15505) );
  NAND4_X1 U17018 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_REG0_REG_17__SCAN_IN), 
        .A3(P2_REG0_REG_2__SCAN_IN), .A4(P2_ADDR_REG_0__SCAN_IN), .ZN(n15502)
         );
  NAND4_X1 U17019 ( .A1(P3_ADDR_REG_1__SCAN_IN), .A2(P3_D_REG_7__SCAN_IN), 
        .A3(P3_D_REG_26__SCAN_IN), .A4(P1_D_REG_28__SCAN_IN), .ZN(n15501) );
  NOR2_X1 U17020 ( .A1(n15502), .A2(n15501), .ZN(n15504) );
  AND4_X1 U17021 ( .A1(P3_D_REG_28__SCAN_IN), .A2(P1_DATAO_REG_23__SCAN_IN), 
        .A3(P2_DATAO_REG_20__SCAN_IN), .A4(P2_REG2_REG_18__SCAN_IN), .ZN(
        n15503) );
  AND4_X1 U17022 ( .A1(n15506), .A2(n15505), .A3(n15504), .A4(n15503), .ZN(
        n15511) );
  NOR4_X1 U17023 ( .A1(n15507), .A2(P3_REG3_REG_14__SCAN_IN), .A3(
        P3_REG3_REG_11__SCAN_IN), .A4(P3_IR_REG_30__SCAN_IN), .ZN(n15509) );
  AND3_X1 U17024 ( .A1(P3_REG3_REG_26__SCAN_IN), .A2(n15509), .A3(n15508), 
        .ZN(n15510) );
  AND4_X1 U17025 ( .A1(n15513), .A2(n15512), .A3(n15511), .A4(n15510), .ZN(
        n15514) );
  NAND4_X1 U17026 ( .A1(n15517), .A2(n15516), .A3(n15515), .A4(n15514), .ZN(
        n15518) );
  XNOR2_X1 U17027 ( .A(n15519), .B(n15518), .ZN(P3_U3519) );
  XOR2_X1 U17028 ( .A(n15521), .B(n15520), .Z(SUB_1596_U59) );
  XNOR2_X1 U17029 ( .A(P2_ADDR_REG_5__SCAN_IN), .B(n15522), .ZN(SUB_1596_U58)
         );
  AOI21_X1 U17030 ( .B1(n15524), .B2(n15523), .A(n15532), .ZN(SUB_1596_U53) );
  XOR2_X1 U17031 ( .A(n15525), .B(n15526), .Z(SUB_1596_U56) );
  NOR2_X1 U17032 ( .A1(n15528), .A2(n15527), .ZN(n15530) );
  XNOR2_X1 U17033 ( .A(n15530), .B(n15529), .ZN(SUB_1596_U60) );
  XOR2_X1 U17034 ( .A(n15532), .B(n15531), .Z(SUB_1596_U5) );
  CLKBUF_X2 U7297 ( .A(n12153), .Z(n12214) );
  CLKBUF_X1 U7304 ( .A(n12153), .Z(n12203) );
  NOR2_X1 U7344 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n7641) );
  CLKBUF_X2 U7345 ( .A(n8594), .Z(n12363) );
  CLKBUF_X1 U7954 ( .A(n14964), .Z(n6721) );
  CLKBUF_X1 U7987 ( .A(n9201), .Z(n9310) );
  CLKBUF_X1 U8460 ( .A(n7938), .Z(n6690) );
  NAND2_X1 U10781 ( .A1(n9049), .A2(n12478), .ZN(n11717) );
  NAND2_X1 U11709 ( .A1(n9340), .A2(n9339), .ZN(n12105) );
  CLKBUF_X3 U14519 ( .A(n7703), .Z(n8134) );
endmodule

